* NGSPICE file created from LSBs_magic_TG_flat.ext - technology: gf180mcuC

.subckt pex_LSBs_magic_TG VDD VSS B1 B2 B3 B4 B5 B6 ITAIL OUT+ OUT- OUT1 OUT2 OUT3 OUT4 OUT5 OUT6 SEL_L C32_D C32_U
X0 TG_0.IN TG_0.IN TG_0.IN VSS.t179 nfet_03v3 ad=64.3p pd=0.44m as=0.156p ps=1.12u w=0.6u l=0.5u
X1 OUT+ SEL_L.t0 TG_0.IN VSS.t19 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 Balance_Inverter_5.Inverter_0.OUT B6.t0 VDD.t208 VDD.t207 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X3 TG_1.IN a_n2280_5855.t12 OUT-.t59 VDD.t279 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 SD3_1 SDn_2.t24 VSS.t508 VSS.t15 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 TG_1.IN.t235 b6.t2 TG_1.IN.t235 VSS.t3 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X6 TG_0.IN TG_0.IN TG_0.IN VSS.t363 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X7 OUT+ SEL_L.t1 TG_0.IN VSS.t428 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X8 OUT6 IT.t24 SD3_1.t44 VSS.t310 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 TG_0.IN b6b.t2 TG_0.IN VSS.t84 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X10 TG_0.IN b2.t2 OUT2.t5 VSS.t153 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 TG_0.IN TG_0.IN TG_0.IN VSS.t172 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X12 OUT+ a_n2265_3941.t12 TG_0.IN VDD.t301 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X13 SD3_1 IT.t25 OUT6.t40 VSS.t311 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X14 TG_1.IN b5b.t2 OUT5.t47 VSS.t152 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 Gc_2 Gc_1.t94 Gc_1.t95 VDD.t0 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X16 VSS G2.t3 SD2_5.t15 VSS.t266 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 TG_1.IN SEL_L.t2 OUT-.t19 VSS.t431 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X18 SDc_2 Gc_2.t96 VDD.t1 VDD.t0 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X19 TG_0.IN a_n2265_3941.t13 OUT+.t68 VDD.t302 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X20 SD3_1 SDn_2.t25 VSS.t509 VSS.t303 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X21 TG_1.IN b4b.t2 OUT4.t7 VSS.t126 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X22 TG_0.IN b5.t2 OUT5.t22 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X23 TG_0.IN TG_0.IN TG_0.IN VSS.t168 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X24 OUT6 IT.t26 SD3_1.t46 VSS.t312 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X25 SDc_2 Gc_1.t96 C32_U.t95 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 OUT6 b6b.t3 TG_1.IN.t93 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X27 VDD SEL_L.t3 a_n2280_5855.t7 VDD.t193 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X28 TG_0.IN b5b.t3 TG_0.IN VSS.t150 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X29 OUT6 b6.t3 TG_0.IN VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X30 TG_1.IN b2b.t2 OUT2.t2 VSS.t315 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 SDc_1 SDn_2.t26 VSS.t511 VSS.t510 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X32 SDc_1 SDn_2.t27 VSS.t512 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X33 TG_0.IN SEL_L.t4 OUT+.t46 VSS.t339 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X34 SD3_1 IT.t27 OUT6.t38 VSS.t313 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X35 OUT- SEL_L.t5 TG_1.IN.t181 VSS.t340 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X36 TG_1.IN SEL_L.t6 OUT-.t18 VSS.t332 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X37 TG_0.IN SEL_L.t7 OUT+.t45 VSS.t333 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X38 TG_1.IN.t92 TG_1.IN.t91 TG_1.IN.t92 VSS.t321 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X39 SD2_5 ITAIL.t2 OUT4.t15 VSS.t328 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X40 b1b B1.t0 VSS.t320 VSS.t319 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X41 VDD Gc_2.t97 SDc_2.t30 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X42 SDc_1 IT.t28 Gc_1.t30 VSS.t314 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X43 VDD Gc_2.t98 SDc_2.t29 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X44 TG_0.IN TG_0.IN TG_0.IN VSS.t361 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X45 TG_1.IN b6b.t4 OUT6.t2 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X46 TG_0.IN SEL_L.t8 OUT+.t44 VSS.t103 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X47 VSS Balance_Inverter_5.Inverter_0.OUT b6.t1 VSS.t582 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X48 SDn_1 IT.t29 OUT5.t12 VSS.t495 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X49 SDn_2 SDn_2.t14 VSS.t507 VSS.t365 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X50 OUT+ a_n2265_3941.t14 TG_0.IN VDD.t303 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X51 OUT5 b5.t3 TG_0.IN VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X52 SDc_2 Gc_2.t99 VDD.t9 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X53 TG_0.IN b3.t2 OUT3.t9 VSS.t89 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X54 VSS SDn_2.t29 SD3_1.t38 VSS.t481 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X55 SDc_2 Gc_2.t100 VDD.t11 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X56 TG_0.IN b6.t4 OUT6.t72 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X57 TG_1.IN.t90 TG_1.IN.t89 TG_1.IN.t90 VSS.t180 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X58 b2b b2.t3 VDD.t79 VDD.t78 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X59 TG_1.IN a_n2280_5855.t13 OUT-.t58 VDD.t280 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X60 OUT6 IT.t30 SD3_1.t55 VSS.t241 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X61 OUT- SEL_L.t11 TG_1.IN.t179 VSS.t79 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X62 SD3_1 IT.t31 OUT6.t36 VSS.t524 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X63 TG_1.IN b6b.t5 OUT6.t3 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X64 TG_1.IN a_n2280_5855.t14 OUT-.t57 VDD.t281 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X65 OUT+ a_n2265_3941.t15 TG_0.IN VDD.t304 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X66 TG_0.IN a_n2265_3941.t16 OUT+.t71 VDD.t305 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X67 Gc_1 IT.t32 SDc_1.t30 VSS.t513 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X68 VDD Gc_2.t62 Gc_2.t63 VDD.t27 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X69 TG_0.IN TG_0.IN TG_0.IN VSS.t362 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X70 C32_U Gc_1.t97 SDc_2.t63 VDD.t98 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X71 TG_1.IN.t88 TG_1.IN.t87 TG_1.IN.t88 VSS.t178 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X72 TG_1.IN.t86 TG_1.IN.t85 TG_1.IN.t86 VSS.t173 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X73 OUT+ a_n2265_3941.t17 TG_0.IN VDD.t306 pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X74 OUT4 b4.t2 TG_0.IN VSS.t160 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X75 Gc_1 Gc_1.t44 Gc_2.t94 VDD.t12 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X76 SD3_1 IT.t33 OUT6.t35 VSS.t247 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X77 TG_1.IN.t84 TG_1.IN.t83 TG_1.IN.t84 VSS.t175 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X78 SD3_1 IT.t34 OUT6.t34 VSS.t533 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X79 SD2_1 G2.t4 VSS.t351 VSS.t269 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X80 VDD Gc_2.t101 SDc_2.t26 VDD.t12 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X81 OUT6 b6.t5 TG_0.IN VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X82 TG_1.IN.t117 b4.t3 TG_1.IN.t117 VSS.t133 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X83 OUT- a_n2280_5855.t15 TG_1.IN.t219 VDD.t282 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X84 OUT+ SEL_L.t13 TG_0.IN VSS.t393 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X85 OUT6 IT.t35 SD3_1.t59 VSS.t535 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X86 SDc_1 IT.t36 Gc_1.t29 VSS.t503 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X87 SDc_1 SDn_2.t30 VSS.t484 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X88 SDn_2 IT.t14 IT.t15 VSS.t371 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X89 TG_1.IN.t118 b4.t4 TG_1.IN.t118 VSS.t161 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X90 SDc_1 SDn_2.t31 VSS.t485 VSS.t377 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X91 TG_1.IN b6b.t6 OUT6.t4 VSS.t67 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X92 TG_0.IN SEL_L.t14 OUT+.t42 VSS.t380 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X93 OUT+ SEL_L.t15 TG_0.IN VSS.t381 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X94 IT G1_2.t24 SD1_1.t13 VDD.t213 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X95 OUT- a_n2280_5855.t16 TG_1.IN.t218 VDD.t314 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X96 SDc_1 IT.t37 Gc_1.t28 VSS.t466 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X97 SDc_1 SDn_2.t32 VSS.t486 VSS.t304 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X98 TG_1.IN.t115 b2.t4 TG_1.IN.t115 VSS.t154 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X99 VSS G2.t5 SD2_4.t7 VSS.t282 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X100 TG_1.IN b6b.t7 OUT6.t5 VSS.t67 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X101 TG_0.IN TG_0.IN TG_0.IN VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X102 OUT6 b6.t6 TG_0.IN VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X103 OUT6 IT.t38 SD3_1.t60 VSS.t249 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X104 TG_0.IN TG_0.IN TG_0.IN VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X105 TG_0.IN a_n2265_3941.t18 OUT+.t73 VDD.t307 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X106 VSS SDn_2.t33 SDn_1.t31 VSS.t376 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X107 G1_1 G1_2.t16 G1_2.t17 VDD.t224 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X108 TG_1.IN.t123 b5.t4 TG_1.IN.t123 VSS.t98 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X109 Gc_2 Gc_2.t60 VDD.t103 VDD.t80 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X110 OUT4 ITAIL.t3 SD2_5.t7 VSS.t124 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X111 C32_U C32_U.t28 C32_D.t95 VSS.t164 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X112 TG_0.IN TG_0.IN TG_0.IN VSS.t173 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X113 SDc_2 Gc_1.t99 C32_U.t93 VDD.t80 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X114 TG_1.IN.t82 TG_1.IN.t81 TG_1.IN.t82 VSS.t173 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X115 TG_1.IN.t80 TG_1.IN.t79 TG_1.IN.t80 VSS.t172 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X116 OUT6 b6b.t8 TG_1.IN.t8 VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X117 TG_1.IN SEL_L.t16 OUT-.t17 VSS.t448 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X118 OUT+ SEL_L.t17 TG_0.IN VSS.t449 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X119 TG_0.IN b6b.t9 TG_0.IN VSS.t69 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X120 OUT6 b6.t7 TG_0.IN VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X121 TG_0.IN SEL_L.t18 OUT+.t39 VSS.t410 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X122 SD2_1 ITAIL.t4 G1_2.t7 VSS.t119 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X123 C32_D C32_D.t62 VSS.t141 VSS.t140 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X124 Gc_2 Gc_2.t58 VDD.t102 VDD.t101 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X125 SDc_1 IT.t39 Gc_1.t27 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X126 VSS C32_D.t60 C32_D.t61 VSS.t164 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X127 TG_1.IN SEL_L.t19 OUT-.t16 VSS.t411 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X128 VDD SEL_L.t20 a_n2265_3941.t6 VDD.t186 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X129 VSS SDn_2.t34 SD3_1.t37 VSS.t373 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X130 G1_2 G1_2.t22 G1_1.t22 VDD.t227 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X131 Balance_Inverter_1.Inverter_0.OUT B3.t0 VDD.t313 VDD.t312 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X132 TG_0.IN b4b.t3 TG_0.IN VSS.t432 nfet_03v3 ad=0.16p pd=1.64u as=0 ps=0 w=0.3u l=0.5u
X133 SDc_1 SDn_2.t35 VSS.t491 VSS.t314 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X134 TG_0.IN b6.t8 OUT6.t68 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X135 TG_1.IN a_n2280_5855.t17 OUT-.t56 VDD.t315 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X136 TG_0.IN b4.t5 OUT4.t17 VSS.t443 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X137 Gc_2 Gc_1.t92 Gc_1.t93 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X138 TG_0.IN SEL_L.t21 OUT+.t38 VSS.t447 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X139 TG_1.IN.t125 b6.t9 TG_1.IN.t125 VSS.t279 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X140 TG_0.IN TG_0.IN TG_0.IN VSS.t172 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X141 TG_0.IN TG_0.IN TG_0.IN VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X142 SDc_2 Gc_2.t104 VDD.t16 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X143 TG_1.IN b6b.t10 OUT6.t7 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X144 OUT5 b5b.t4 TG_1.IN.t98 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X145 Gc_1 Gc_1.t42 Gc_2.t92 VDD.t30 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X146 C32_D C32_U.t60 C32_U.t61 VSS.t140 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X147 C32_U C32_U.t12 C32_D.t93 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X148 VSS SDn_2.t36 SD3_1.t36 VSS.t492 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X149 G1_2 ITAIL.t5 SD2_1.t7 VSS.t122 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X150 OUT6 IT.t40 SD3_1.t0 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X151 SD1_1 G1_2.t26 IT.t17 VDD.t214 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X152 TG_1.IN.t109 b5.t5 TG_1.IN.t109 VSS.t139 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X153 SDn_1 SDn_2.t37 VSS.t496 VSS.t495 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X154 OUT5 b5.t6 TG_0.IN VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X155 OUT- SEL_L.t23 TG_1.IN.t176 VSS.t408 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X156 VDD G1_1.t24 SD1_1.t2 VDD.t218 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X157 OUT- SEL_L.t24 TG_1.IN.t175 VSS.t433 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X158 SD3_1 IT.t41 OUT6.t30 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X159 VSS SDn_2.t38 SDn_1.t29 VSS.t497 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X160 TG_1.IN.t78 TG_1.IN.t77 TG_1.IN.t78 VSS.t171 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X161 TG_1.IN.t76 TG_1.IN.t75 TG_1.IN.t76 VSS.t170 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X162 OUT5 b5b.t5 TG_1.IN.t253 VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X163 Gc_1 Gc_1.t40 Gc_2.t91 VDD.t29 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X164 TG_0.IN a_n2265_3941.t19 OUT+.t49 VDD.t283 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X165 TG_1.IN.t136 b5.t7 TG_1.IN.t136 VSS.t128 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X166 OUT- SEL_L.t25 TG_1.IN.t174 VSS.t434 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X167 TG_0.IN b6.t10 OUT6.t67 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X168 OUT6 IT.t42 SD3_1.t2 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X169 SDn_1 IT.t43 OUT5.t11 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X170 VSS C32_D.t58 C32_D.t59 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X171 TG_0.IN a_n2265_3941.t20 OUT+.t50 VDD.t284 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X172 G1_2 G1_2.t20 G1_1.t21 VDD.t226 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X173 OUT- a_n2280_5855.t18 TG_1.IN.t216 VDD.t316 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X174 VDD Gc_2.t56 Gc_2.t57 VDD.t98 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X175 Gc_1 Gc_1.t38 Gc_2.t90 VDD.t28 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X176 TG_0.IN b6.t11 OUT6.t66 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X177 OUT- SEL_L.t27 TG_1.IN.t173 VSS.t383 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X178 OUT+ SEL_L.t28 TG_0.IN VSS.t394 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X179 TG_0.IN b6b.t11 TG_0.IN VSS.t70 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X180 TG_0.IN TG_0.IN TG_0.IN VSS.t325 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X181 VDD Gc_2.t54 Gc_2.t55 VDD.t124 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X182 VSS G2.t6 SD2_5.t14 VSS.t111 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X183 VDD b3b.t2 b3.t1 VDD.t343 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X184 VSS Balance_Inverter_0.Inverter_0.OUT b4.t1 VSS.t593 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X185 OUT6 b6b.t12 TG_1.IN.t10 VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X186 OUT- SEL_L.t29 TG_1.IN.t172 VSS.t395 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X187 TG_0.IN TG_0.IN TG_0.IN VSS.t167 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X188 OUT6 IT.t44 SD3_1.t3 VSS.t14 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X189 VSS G2.t7 SD2_5.t13 VSS.t266 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X190 Gc_1 Gc_1.t36 Gc_2.t89 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X191 TG_0.IN TG_0.IN TG_0.IN VSS.t180 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X192 SD3_1 IT.t45 OUT6.t27 VSS.t15 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X193 VSS SDn_2.t39 SDn_1.t28 VSS.t307 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X194 VDD G1_1.t14 G1_1.t15 VDD.t142 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X195 OUT5 b5b.t6 TG_1.IN.t252 VSS.t96 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X196 TG_0.IN TG_0.IN TG_0.IN VSS.t180 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X197 TG_1.IN SEL_L.t30 OUT-.t15 VSS.t337 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X198 SDc_1 SDn_2.t40 VSS.t502 VSS.t308 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X199 TG_1.IN b1b.t2 OUT1.t1 VSS.t372 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X200 SDc_1 SDn_2.t41 VSS.t504 VSS.t503 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X201 OUT+ a_n2265_3941.t21 TG_0.IN VDD.t285 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X202 SD3_1 SDn_2.t42 VSS.t464 VSS.t311 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X203 SDc_1 IT.t46 Gc_1.t26 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X204 OUT- a_n2280_5855.t19 TG_1.IN.t215 VDD.t317 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X205 OUT3 ITAIL.t6 SD2_4.t3 VSS.t123 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X206 OUT6 b6b.t13 TG_1.IN.t239 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X207 SDn_1 IT.t47 OUT5.t10 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X208 SDc_1 SDn_2.t43 VSS.t465 VSS.t309 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X209 SDc_1 IT.t48 Gc_1.t25 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X210 TG_1.IN.t126 b6.t12 TG_1.IN.t126 VSS.t69 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X211 SDc_2 Gc_2.t105 VDD.t18 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X212 SDc_1 SDn_2.t44 VSS.t467 VSS.t466 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X213 SDc_1 IT.t49 Gc_1.t24 VSS.t304 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X214 SD3_1 IT.t50 OUT6.t26 VSS.t305 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X215 TG_1.IN.t137 b5.t8 TG_1.IN.t137 VSS.t318 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X216 SDc_1 SDn_2.t45 VSS.t469 VSS.t468 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X217 VSS SDn_2.t46 SD3_1.t34 VSS.t312 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X218 SDn_1 IT.t51 OUT5.t9 VSS.t306 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X219 SDc_1 IT.t52 Gc_1.t23 VSS.t254 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X220 OUT+ a_n2265_3941.t22 TG_0.IN VDD.t286 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X221 SD1_1 G1_1.t25 VDD.t116 VDD.t115 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X222 SDc_2 Gc_1.t104 C32_U.t92 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X223 TG_1.IN SEL_L.t31 OUT-.t14 VSS.t338 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X224 SD3_1 SDn_2.t47 VSS.t472 VSS.t313 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X225 TG_0.IN b3b.t3 TG_0.IN VSS.t58 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X226 OUT5 b5b.t7 TG_1.IN.t251 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X227 TG_1.IN SEL_L.t32 OUT-.t13 VSS.t198 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X228 TG_0.IN TG_0.IN TG_0.IN VSS.t326 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X229 VSS SDn_2.t48 SDn_1.t27 VSS.t302 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X230 OUT5 b5.t9 TG_0.IN VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X231 Gc_1 Gc_1.t34 Gc_2.t88 VDD.t27 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X232 VDD Gc_2.t106 SDc_2.t23 VDD.t27 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X233 OUT6 b6.t13 TG_0.IN VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X234 TG_1.IN a_n2280_5855.t20 OUT-.t55 VDD.t308 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X235 OUT6 b6b.t14 TG_1.IN.t240 VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X236 SD3_1 SDn_2.t49 VSS.t475 VSS.t385 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X237 TG_0.IN b4b.t4 TG_0.IN VSS.t589 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X238 C32_D C32_D.t56 VSS.t422 VSS.t322 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X239 Gc_2 Gc_1.t90 Gc_1.t91 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X240 VSS SDn_2.t50 SDn_1.t26 VSS.t476 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X241 TG_1.IN.t127 b6.t14 TG_1.IN.t127 VSS.t8 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X242 TG_1.IN b5b.t8 OUT5.t42 VSS.t127 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X243 Gc_2 Gc_2.t52 VDD.t332 VDD.t46 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X244 Gc_1 IT.t53 SDc_1.t22 VSS.t259 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X245 OUT- a_n2280_5855.t21 TG_1.IN.t213 VDD.t309 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X246 TG_0.IN a_n2265_3941.t23 OUT+.t53 VDD.t287 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X247 SDn_1 SDn_2.t51 VSS.t480 VSS.t479 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X248 TG_1.IN.t256 b4.t6 TG_1.IN.t256 VSS.t591 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X249 VSS SDn_2.t52 SD3_1.t31 VSS.t241 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X250 G1_1 G1_1.t12 VDD.t148 VDD.t147 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X251 TG_0.IN TG_0.IN TG_0.IN VSS.t325 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X252 TG_1.IN.t128 b6.t15 TG_1.IN.t128 VSS.t70 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X253 TG_0.IN SEL_L.t33 OUT+.t36 VSS.t199 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X254 TG_0.IN b6b.t15 TG_0.IN VSS.t3 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X255 TG_0.IN b5.t10 OUT5.t28 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X256 C32_D C32_U.t58 C32_U.t59 VSS.t322 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X257 OUT- SEL_L.t34 TG_1.IN.t168 VSS.t341 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X258 SD2_1 G2.t8 VSS.t270 VSS.t269 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X259 SD2_5 G2.t9 VSS.t271 VSS.t72 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X260 VSS C32_D.t54 C32_D.t55 VSS.t116 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X261 SDn_2 SDn_2.t12 VSS.t506 VSS.t369 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X262 TG_1.IN.t130 b6.t16 TG_1.IN.t130 VSS.t84 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X263 TG_1.IN.t131 b6.t17 TG_1.IN.t131 VSS.t4 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X264 TG_0.IN a_n2265_3941.t24 OUT+.t54 VDD.t288 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X265 TG_1.IN.t74 TG_1.IN.t73 TG_1.IN.t74 VSS.t169 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X266 VSS Balance_Inverter_2.Inverter_0.OUT b2.t1 VSS.t456 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X267 OUT5 b5b.t9 TG_1.IN.t249 VSS.t96 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X268 Balance_Inverter_3.Inverter_0.OUT B1.t1 VSS.t78 VSS.t77 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X269 VSS SDn_2.t54 SD3_1.t30 VSS.t244 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X270 VSS G2.t10 SD2_1.t13 VSS.t74 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X271 SD3_1 SDn_2.t55 VSS.t248 VSS.t247 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X272 TG_1.IN.t72 TG_1.IN.t71 TG_1.IN.t72 VSS.t168 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X273 C32_U C32_U.t62 C32_D.t91 VSS.t116 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X274 TG_1.IN.t132 b6.t18 TG_1.IN.t132 VSS.t7 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X275 OUT5 IT.t54 SDn_1.t11 VSS.t307 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X276 TG_1.IN b6b.t16 OUT6.t92 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X277 VSS G2.t11 SD2_4.t6 VSS.t282 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X278 SD2_3 G2.t12 VSS.t285 VSS.t182 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X279 OUT+ SEL_L.t35 TG_0.IN VSS.t342 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X280 TG_1.IN SEL_L.t36 OUT-.t12 VSS.t343 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X281 OUT+ SEL_L.t37 TG_0.IN VSS.t344 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X282 Gc_1 Gc_1.t32 Gc_2.t86 VDD.t26 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X283 TG_1.IN b6b.t17 OUT6.t93 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X284 SDn_2 SDn_2.t10 VSS.t505 VSS.t371 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X285 TG_1.IN a_n2280_5855.t22 OUT-.t54 VDD.t310 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X286 TG_1.IN.t99 b3.t3 TG_1.IN.t99 VSS.t94 nfet_03v3 ad=0.16p pd=1.64u as=0 ps=0 w=0.3u l=0.5u
X287 OUT4 b4b.t5 TG_1.IN.t255 VSS.t590 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X288 TG_0.IN b6.t19 OUT6.t64 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X289 OUT+ SEL_L.t38 TG_0.IN VSS.t345 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X290 SDc_2 Gc_1.t107 C32_U.t91 VDD.t0 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X291 TG_1.IN.t70 TG_1.IN.t69 TG_1.IN.t70 VSS.t167 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X292 TG_0.IN b6.t20 OUT6.t63 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X293 OUT6 b6b.t18 TG_1.IN.t243 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X294 OUT6 b6b.t19 TG_1.IN.t244 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X295 OUT+ a_n2265_3941.t25 TG_0.IN VDD.t295 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X296 SDn_2 IT.t12 IT.t13 VSS.t370 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X297 Gc_2 Gc_1.t88 Gc_1.t89 VDD.t101 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X298 TG_0.IN TG_0.IN TG_0.IN VSS.t177 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X299 OUT4 ITAIL.t7 SD2_5.t0 VSS.t124 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X300 G2 ITAIL.t0 ITAIL.t1 VSS.t183 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X301 VSS SDn_2.t57 SD3_1.t28 VSS.t249 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X302 SDc_2 Gc_2.t108 VDD.t253 VDD.t101 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X303 VDD SEL_L.t39 a_n2280_5855.t5 VDD.t181 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X304 C32_U Gc_1.t108 SDc_2.t62 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X305 VDD b1b.t3 b1.t0 VDD.t34 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X306 C32_U Gc_1.t109 SDc_2.t61 VDD.t124 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X307 VDD Gc_2.t109 SDc_2.t21 VDD.t26 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X308 SDc_1 IT.t55 Gc_1.t22 VSS.t308 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X309 TG_0.IN b4b.t6 TG_0.IN VSS.t440 nfet_03v3 ad=0.16p pd=1.64u as=0 ps=0 w=0.3u l=0.5u
X310 VDD SEL_L.t40 a_n2280_5855.t4 VDD.t178 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X311 VDD Gc_2.t50 Gc_2.t51 VDD.t30 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X312 VDD Gc_2.t48 Gc_2.t49 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X313 OUT- a_n2280_5855.t23 TG_1.IN.t211 VDD.t149 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X314 SDn_1 SDn_2.t58 VSS.t252 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X315 TG_0.IN SEL_L.t41 OUT+.t32 VSS.t35 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X316 SDc_1 IT.t56 Gc_1.t21 VSS.t309 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X317 SDc_1 SDn_2.t59 VSS.t253 VSS.t18 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X318 SD1_1 G1_2.t28 IT.t18 VDD.t215 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X319 C32_U Gc_1.t110 SDc_2.t60 VDD.t30 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X320 TG_1.IN SEL_L.t42 OUT-.t11 VSS.t401 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X321 TG_0.IN b4b.t7 TG_0.IN VSS.t441 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X322 SDc_2 Gc_2.t110 VDD.t256 VDD.t68 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X323 Gc_1 Gc_1.t62 Gc_2.t84 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X324 TG_0.IN a_n2265_3941.t26 OUT+.t62 VDD.t296 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X325 OUT+ a_n2265_3941.t27 TG_0.IN VDD.t297 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X326 SDc_1 IT.t57 Gc_1.t20 VSS.t468 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X327 b5b b5.t11 VDD.t244 VDD.t243 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X328 SDc_2 Gc_1.t112 C32_U.t87 VDD.t70 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X329 G1_1 G1_1.t10 VDD.t146 VDD.t145 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X330 SDn_1 IT.t58 OUT5.t8 VSS.t479 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X331 VDD Gc_2.t46 Gc_2.t47 VDD.t29 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X332 SDc_1 SDn_2.t60 VSS.t255 VSS.t254 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X333 VSS G2.t13 SD2_3.t2 VSS.t106 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X334 TG_0.IN b6.t21 OUT6.t62 VSS.t67 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X335 OUT- SEL_L.t43 TG_1.IN.t165 VSS.t402 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X336 C32_U Gc_1.t113 SDc_2.t59 VDD.t29 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X337 TG_0.IN b6b.t20 TG_0.IN VSS.t4 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X338 G1_2 ITAIL.t8 SD2_1.t6 VSS.t122 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X339 SD2_5 ITAIL.t9 OUT4.t9 VSS.t125 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X340 C32_U Gc_1.t114 SDc_2.t58 VDD.t27 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X341 Gc_1 Gc_1.t60 Gc_2.t83 VDD.t98 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X342 VDD Gc_2.t44 Gc_2.t45 VDD.t28 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X343 TG_1.IN.t68 TG_1.IN.t67 TG_1.IN.t68 VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X344 TG_1.IN a_n2280_5855.t24 OUT-.t53 VDD.t150 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X345 TG_0.IN SEL_L.t44 OUT+.t31 VSS.t200 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X346 SD3_1 SDn_2.t61 VSS.t256 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X347 VDD Gc_2.t111 SDc_2.t19 VDD.t98 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X348 C32_U Gc_1.t116 SDc_2.t57 VDD.t28 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X349 VDD Gc_2.t112 SDc_2.t18 VDD.t29 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X350 OUT5 b5.t12 TG_0.IN VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X351 Gc_1 Gc_1.t58 Gc_2.t82 VDD.t124 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X352 SD2_5 G2.t14 VSS.t110 VSS.t109 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X353 TG_1.IN a_n2280_5855.t25 OUT-.t52 VDD.t151 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X354 VDD Gc_2.t113 SDc_2.t17 VDD.t124 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X355 Gc_2 Gc_1.t86 Gc_1.t87 VDD.t87 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X356 VDD G1_1.t8 G1_1.t9 VDD.t112 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X357 OUT5 b5b.t10 TG_1.IN.t250 VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X358 VDD Gc_2.t42 Gc_2.t43 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X359 TG_0.IN b6b.t21 TG_0.IN VSS.t7 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X360 TG_1.IN a_n2280_5855.t26 OUT-.t51 VDD.t318 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X361 OUT+ a_n2265_3941.t28 TG_0.IN VDD.t298 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X362 OUT6 IT.t59 SD3_1.t54 VSS.t492 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X363 VSS SDn_2.t62 SD3_1.t26 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X364 b5b B5.t0 VSS.t130 VSS.t129 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X365 TG_0.IN a_n2265_3941.t29 OUT+.t65 VDD.t299 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X366 TG_0.IN b4b.t8 TG_0.IN VSS.t442 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X367 TG_0.IN b5b.t11 TG_0.IN VSS.t151 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X368 SDc_2 Gc_1.t118 C32_U.t83 VDD.t82 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X369 C32_U Gc_1.t119 SDc_2.t56 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X370 VSS SDn_2.t63 SDc_1.t50 VSS.t259 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X371 SD3_1 SDn_2.t64 VSS.t556 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X372 VSS SDn_2.t8 SDn_2.t9 VSS.t364 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X373 VSS G2.t15 SD2_5.t10 VSS.t111 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X374 VDD Gc_2.t40 Gc_2.t41 VDD.t54 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X375 TG_1.IN SEL_L.t46 OUT-.t10 VSS.t451 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X376 b3b b3.t4 VDD.t38 VDD.t37 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X377 SD1_1 G1_1.t28 VDD.t118 VDD.t117 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X378 TG_0.IN b5b.t12 TG_0.IN VSS.t463 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X379 TG_0.IN b5b.t13 TG_0.IN VSS.t93 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X380 OUT+ SEL_L.t47 TG_0.IN VSS.t452 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X381 VSS SDn_2.t6 SDn_2.t7 VSS.t367 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X382 TG_1.IN.t257 b4.t7 TG_1.IN.t257 VSS.t222 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X383 TG_1.IN.t66 TG_1.IN.t65 TG_1.IN.t66 VSS.t325 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X384 SD3_1 SDn_2.t65 VSS.t557 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X385 TG_1.IN b6b.t22 OUT6.t74 VSS.t67 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X386 VDD b4b.t9 b4.t0 VDD.t248 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X387 VDD G1_1.t29 SD1_1.t14 VDD.t270 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X388 TG_0.IN b6.t22 OUT6.t61 VSS.t67 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X389 Balance_Inverter_0.Inverter_0.OUT B4.t0 VSS.t186 VSS.t185 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X390 TG_1.IN.t64 TG_1.IN.t63 TG_1.IN.t64 VSS.t167 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X391 OUT4 b4.t8 TG_0.IN VSS.t137 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X392 TG_0.IN SEL_L.t48 OUT+.t29 VSS.t453 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X393 SD1_1 G1_2.t29 IT.t19 VDD.t216 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X394 OUT3 ITAIL.t10 SD2_4.t2 VSS.t123 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X395 OUT5 b5.t13 TG_0.IN VSS.t96 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X396 TG_0.IN TG_0.IN TG_0.IN VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X397 VSS SDn_2.t66 SD3_1.t23 VSS.t14 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X398 TG_1.IN.t62 TG_1.IN.t61 TG_1.IN.t62 VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X399 OUT- a_n2280_5855.t27 TG_1.IN.t207 VDD.t319 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X400 OUT- a_n2280_5855.t28 TG_1.IN.t206 VDD.t320 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X401 TG_0.IN b5b.t14 TG_0.IN VSS.t150 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X402 SD1_1 G1_1.t30 VDD.t274 VDD.t273 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X403 TG_0.IN TG_0.IN TG_0.IN VSS.t173 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X404 OUT4 b4b.t10 TG_1.IN.t245 VSS.t160 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X405 OUT6 b6.t23 TG_0.IN VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X406 OUT- a_n2280_5855.t29 TG_1.IN.t205 VDD.t95 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X407 TG_0.IN b2b.t3 TG_0.IN VSS.t316 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X408 OUT6 b6b.t23 TG_1.IN.t120 VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X409 Gc_2 Gc_2.t38 VDD.t327 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X410 TG_0.IN TG_0.IN TG_0.IN VSS.t361 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X411 C32_D C32_U.t56 C32_U.t57 VSS.t174 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X412 SD3_1 SDn_2.t67 VSS.t560 VSS.t305 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X413 G1_2 ITAIL.t11 SD2_1.t5 VSS.t181 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X414 VDD G1_1.t6 G1_1.t7 VDD.t41 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X415 TG_1.IN b4b.t11 OUT4.t4 VSS.t443 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X416 SDc_2 Gc_1.t120 C32_U.t81 VDD.t17 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X417 Gc_2 Gc_1.t84 Gc_1.t85 VDD.t46 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X418 TG_1.IN b6b.t24 OUT6.t76 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X419 b4b B4.t1 VSS.t188 VSS.t187 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X420 SDn_1 SDn_2.t68 VSS.t561 VSS.t306 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X421 G1_1 G1_1.t4 VDD.t40 VDD.t39 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X422 TG_0.IN b4.t9 OUT4.t19 VSS.t138 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X423 SDc_2 Gc_2.t115 VDD.t47 VDD.t46 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X424 OUT5 IT.t60 SDn_1.t9 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X425 OUT+ SEL_L.t49 TG_0.IN VSS.t80 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X426 SDn_1 SDn_2.t69 VSS.t562 VSS.t387 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X427 VDD SEL_L.t50 a_n2265_3941.t4 VDD.t173 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X428 TG_1.IN.t100 b3.t5 TG_1.IN.t100 VSS.t90 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X429 OUT1 b1.t2 TG_0.IN VSS.t295 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X430 TG_1.IN.t60 TG_1.IN.t59 TG_1.IN.t60 VSS.t324 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X431 TG_1.IN a_n2280_5855.t30 OUT-.t50 VDD.t96 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X432 C32_D C32_D.t52 VSS.t212 VSS.t174 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X433 VSS SDn_2.t70 SDc_1.t49 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X434 OUT5 IT.t61 SDn_1.t8 VSS.t497 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X435 OUT5 IT.t62 SDn_1.t7 VSS.t476 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X436 VDD b5b.t15 b5.t1 VDD.t75 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X437 TG_1.IN.t58 TG_1.IN.t57 TG_1.IN.t58 VSS.t180 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X438 TG_1.IN SEL_L.t51 OUT-.t9 VSS.t81 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X439 VDD SEL_L.t52 a_n2265_3941.t3 VDD.t170 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X440 OUT5 IT.t63 SDn_1.t6 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X441 TG_1.IN.t258 b4.t10 TG_1.IN.t258 VSS.t592 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X442 Gc_1 IT.t64 SDc_1.t18 VSS.t549 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X443 OUT6 b6.t24 TG_0.IN VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X444 OUT+ a_n2265_3941.t30 TG_0.IN VDD.t300 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X445 VSS SDn_2.t71 SD3_1.t21 VSS.t56 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X446 TG_1.IN b5b.t16 OUT5.t39 VSS.t152 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X447 TG_1.IN a_n2280_5855.t31 OUT-.t49 VDD.t97 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X448 Gc_1 IT.t65 SDc_1.t17 VSS.t384 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X449 OUT6 b6.t25 TG_0.IN VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X450 TG_1.IN SEL_L.t53 OUT-.t8 VSS.t429 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X451 OUT+ SEL_L.t54 TG_0.IN VSS.t430 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X452 SD3_1 IT.t66 OUT6.t24 VSS.t385 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X453 SD1_1 G1_2.t30 IT.t20 VDD.t217 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X454 TG_0.IN SEL_L.t55 OUT+.t26 VSS.t329 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X455 SD2_5 G2.t16 VSS.t73 VSS.t72 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X456 TG_0.IN TG_0.IN TG_0.IN VSS.t170 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X457 TG_0.IN b5.t14 OUT5.t2 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X458 OUT6 IT.t67 SD3_1.t51 VSS.t26 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X459 TG_1.IN.t260 b4.t11 TG_1.IN.t260 VSS.t596 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X460 SDn_2 IT.t10 IT.t11 VSS.t369 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X461 TG_0.IN TG_0.IN TG_0.IN VSS.t360 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X462 TG_0.IN TG_0.IN TG_0.IN VSS.t359 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X463 OUT+ SEL_L.t56 TG_0.IN VSS.t330 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X464 VDD Gc_2.t36 Gc_2.t37 VDD.t26 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X465 OUT3 b3.t6 TG_0.IN VSS.t95 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X466 C32_U Gc_1.t121 SDc_2.t55 VDD.t26 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X467 SD3_1 IT.t68 OUT6.t22 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X468 VSS G2.t17 SD2_1.t12 VSS.t74 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X469 OUT- SEL_L.t57 TG_1.IN.t161 VSS.t331 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X470 TG_0.IN b6.t26 OUT6.t57 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X471 TG_0.IN a_n2265_3941.t31 OUT+.t0 VDD.t106 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X472 Balance_Inverter_2.Inverter_0.OUT B2.t0 VSS.t265 VSS.t264 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X473 TG_1.IN b6b.t25 OUT6.t77 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X474 SDn_1 SDn_2.t72 VSS.t567 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X475 SD2_3 ITAIL.t12 OUT2.t0 VSS.t182 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X476 TG_0.IN b6b.t26 TG_0.IN VSS.t69 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X477 TG_0.IN b6b.t27 TG_0.IN VSS.t279 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X478 TG_0.IN a_n2265_3941.t32 OUT+.t1 VDD.t107 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X479 OUT- SEL_L.t59 TG_1.IN.t160 VSS.t418 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X480 OUT6 IT.t69 SD3_1.t53 VSS.t244 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X481 SDn_1 IT.t70 OUT5.t7 VSS.t386 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X482 TG_1.IN.t56 TG_1.IN.t55 TG_1.IN.t56 VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X483 C32_U C32_U.t0 C32_D.t89 VSS.t207 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X484 Gc_1 Gc_1.t56 Gc_2.t79 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X485 TG_0.IN TG_0.IN TG_0.IN VSS.t180 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X486 C32_U Gc_1.t123 SDc_2.t54 VDD.t54 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X487 VDD Gc_2.t116 SDc_2.t15 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X488 TG_1.IN.t54 TG_1.IN.t53 TG_1.IN.t54 VSS.t180 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X489 TG_0.IN b6b.t28 TG_0.IN VSS.t8 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X490 TG_0.IN SEL_L.t60 OUT+.t24 VSS.t419 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X491 IT IT.t8 SDn_2.t20 VSS.t368 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X492 SD2_2 ITAIL.t13 OUT1.t0 VSS.t183 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X493 VDD Gc_2.t34 Gc_2.t35 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X494 IT IT.t6 SDn_2.t19 VSS.t367 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X495 SDn_1 IT.t73 OUT5.t6 VSS.t387 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X496 C32_D C32_D.t50 VSS.t211 VSS.t210 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X497 OUT- a_n2280_5855.t32 TG_1.IN.t202 VDD.t204 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X498 TG_1.IN.t52 TG_1.IN.t51 TG_1.IN.t52 VSS.t323 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X499 OUT4 ITAIL.t14 SD2_5.t2 VSS.t184 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X500 C32_U Gc_1.t124 SDc_2.t53 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X501 Balance_Inverter_4.Inverter_0.OUT B5.t1 VSS.t132 VSS.t131 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X502 TG_0.IN b3b.t4 TG_0.IN VSS.t61 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X503 TG_1.IN.t102 b5.t15 TG_1.IN.t102 VSS.t98 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X504 b2b B2.t1 VSS.t263 VSS.t262 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X505 OUT6 b6.t27 TG_0.IN VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X506 TG_0.IN b4b.t12 TG_0.IN VSS.t133 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X507 b1b b1.t3 VDD.t141 VDD.t140 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X508 C32_D C32_U.t54 C32_U.t55 VSS.t145 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X509 VSS C32_D.t48 C32_D.t49 VSS.t207 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X510 SDn_1 SDn_2.t73 VSS.t568 VSS.t374 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X511 TG_1.IN.t129 b6.t28 TG_1.IN.t129 VSS.t3 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X512 SDc_2 Gc_2.t117 VDD.t51 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X513 OUT- a_n2280_5855.t33 TG_1.IN.t201 VDD.t205 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X514 SD3_1 SDn_2.t74 VSS.t538 VSS.t301 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X515 TG_0.IN b6b.t29 TG_0.IN VSS.t84 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X516 TG_1.IN.t50 TG_1.IN.t49 TG_1.IN.t50 VSS.t178 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X517 TG_1.IN.t48 TG_1.IN.t47 TG_1.IN.t48 VSS.t173 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X518 SDn_1 SDn_2.t75 VSS.t539 VSS.t386 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X519 VSS C32_D.t46 C32_D.t47 VSS.t204 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X520 TG_1.IN.t46 TG_1.IN.t45 TG_1.IN.t46 VSS.t177 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X521 C32_U C32_U.t26 C32_D.t87 VSS.t102 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X522 C32_D C32_U.t52 C32_U.t53 VSS.t210 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X523 Gc_2 Gc_2.t32 VDD.t322 VDD.t82 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X524 OUT6 b6.t29 TG_0.IN VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X525 VDD Gc_2.t119 SDc_2.t13 VDD.t30 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X526 VSS C32_D.t44 C32_D.t45 VSS.t147 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X527 C32_D C32_D.t42 VSS.t146 VSS.t145 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X528 OUT+ a_n2265_3941.t33 TG_0.IN VDD.t108 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X529 OUT6 b6.t30 TG_0.IN VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X530 OUT+ a_n2265_3941.t34 TG_0.IN VDD.t109 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X531 TG_1.IN b4b.t13 OUT4.t3 VSS.t134 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X532 TG_0.IN TG_0.IN TG_0.IN VSS.t168 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X533 TG_0.IN TG_0.IN TG_0.IN VSS.t170 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X534 C32_D C32_U.t50 C32_U.t51 VSS.t225 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X535 Gc_2 Gc_2.t30 VDD.t321 VDD.t87 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X536 OUT2 ITAIL.t15 SD2_3.t0 VSS.t106 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X537 TG_1.IN SEL_L.t61 OUT-.t7 VSS.t196 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X538 TG_0.IN b6b.t30 TG_0.IN VSS.t70 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X539 SDc_2 Gc_1.t125 C32_U.t77 VDD.t87 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X540 OUT+ a_n2265_3941.t35 TG_0.IN VDD.t110 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X541 TG_0.IN TG_0.IN TG_0.IN VSS.t172 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X542 C32_D C32_D.t40 VSS.t144 VSS.t115 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X543 C32_U C32_U.t24 C32_D.t84 VSS.t204 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X544 TG_0.IN b6.t31 OUT6.t53 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X545 SD2_5 ITAIL.t16 OUT4.t12 VSS.t125 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X546 TG_0.IN b5.t16 OUT5.t19 VSS.t127 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X547 VSS C32_D.t38 C32_D.t39 VSS.t102 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X548 Gc_2 Gc_1.t82 Gc_1.t83 VDD.t68 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X549 TG_0.IN TG_0.IN TG_0.IN VSS.t167 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X550 C32_D C32_D.t36 VSS.t230 VSS.t114 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X551 VSS C32_D.t34 C32_D.t35 VSS.t227 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X552 TG_1.IN b6b.t31 OUT6.t78 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X553 TG_0.IN TG_0.IN TG_0.IN VSS.t167 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X554 Balance_Inverter_3.Inverter_0.OUT B1.t2 VDD.t126 VDD.t125 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X555 C32_U C32_U.t22 C32_D.t83 VSS.t147 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X556 TG_1.IN a_n2280_5855.t34 OUT-.t48 VDD.t206 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X557 SD2_5 G2.t18 VSS.t585 VSS.t109 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X558 TG_1.IN b5b.t17 OUT5.t38 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X559 Gc_1 Gc_1.t54 Gc_2.t77 VDD.t54 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X560 Gc_1 IT.t74 SDc_1.t16 VSS.t29 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X561 VSS SDn_2.t76 SD3_1.t19 VSS.t540 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X562 C32_U C32_U.t20 C32_D.t82 VSS.t292 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X563 C32_D C32_D.t32 VSS.t226 VSS.t225 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X564 SD2_4 G2.t19 VSS.t586 VSS.t274 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X565 VDD Gc_2.t121 SDc_2.t12 VDD.t54 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X566 VSS SDn_2.t77 SDc_1.t48 VSS.t296 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X567 Gc_1 IT.t75 SDc_1.t15 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X568 C32_D C32_U.t48 C32_U.t49 VSS.t115 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X569 SD3_1 IT.t76 OUT6.t20 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X570 TG_1.IN.t104 b5.t17 TG_1.IN.t104 VSS.t128 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X571 TG_0.IN a_n2265_3941.t36 OUT+.t5 VDD.t111 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X572 TG_0.IN SEL_L.t62 OUT+.t23 VSS.t197 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X573 C32_D C32_U.t46 C32_U.t47 VSS.t114 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X574 VSS SDn_2.t78 SDc_1.t47 VSS.t297 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X575 VSS SDn_2.t79 SDc_1.t46 VSS.t298 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X576 VSS SDn_2.t80 SDc_1.t45 VSS.t549 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X577 TG_1.IN.t139 b6.t32 TG_1.IN.t139 VSS.t279 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X578 C32_U C32_U.t18 C32_D.t79 VSS.t227 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X579 OUT- a_n2280_5855.t35 TG_1.IN.t199 VDD.t200 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X580 TG_1.IN a_n2280_5855.t36 OUT-.t47 VDD.t201 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X581 TG_0.IN a_n2265_3941.t37 OUT+.t74 VDD.t335 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X582 TG_0.IN TG_0.IN TG_0.IN VSS.t358 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X583 C32_D C32_U.t44 C32_U.t45 VSS.t290 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X584 VSS SDn_2.t81 SDc_1.t44 VSS.t384 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X585 TG_0.IN TG_0.IN TG_0.IN VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X586 OUT- SEL_L.t63 TG_1.IN.t158 VSS.t335 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X587 TG_0.IN SEL_L.t64 OUT+.t22 VSS.t336 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X588 TG_1.IN.t44 TG_1.IN.t43 TG_1.IN.t44 VSS.t172 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X589 C32_D C32_D.t30 VSS.t224 VSS.t223 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X590 VSS C32_D.t28 C32_D.t29 VSS.t292 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X591 Gc_1 IT.t77 SDc_1.t14 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X592 TG_0.IN a_n2265_3941.t38 OUT+.t75 VDD.t336 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X593 TG_1.IN b3b.t5 OUT3.t11 VSS.t60 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X594 TG_1.IN.t42 TG_1.IN.t41 TG_1.IN.t42 VSS.t176 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X595 SD3_1 IT.t78 OUT6.t19 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X596 VSS Balance_Inverter_4.Inverter_0.OUT b5.t0 VSS.t99 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X597 b4b b4.t12 VDD.t342 VDD.t341 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X598 C32_D C32_D.t26 VSS.t291 VSS.t290 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X599 VSS C32_D.t24 C32_D.t25 VSS.t86 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X600 TG_1.IN b6b.t32 OUT6.t79 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X601 TG_0.IN b6.t33 OUT6.t52 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X602 C32_D C32_U.t42 C32_U.t43 VSS.t223 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X603 C32_U Gc_1.t127 SDc_2.t52 VDD.t72 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X604 VDD Gc_2.t122 SDc_2.t11 VDD.t22 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X605 TG_0.IN b6.t34 OUT6.t51 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X606 OUT+ SEL_L.t66 TG_0.IN VSS.t334 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X607 TG_0.IN TG_0.IN TG_0.IN VSS.t176 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X608 TG_1.IN b6b.t33 OUT6.t80 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X609 OUT- SEL_L.t67 TG_1.IN.t157 VSS.t201 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X610 SD3_1 IT.t79 OUT6.t18 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X611 VDD Gc_2.t123 SDc_2.t10 VDD.t28 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X612 VSS SDn_2.t82 SDc_1.t43 VSS.t300 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X613 OUT- a_n2280_5855.t37 TG_1.IN.t197 VDD.t202 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X614 VDD Gc_2.t28 Gc_2.t29 VDD.t72 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X615 TG_0.IN b3b.t6 TG_0.IN VSS.t58 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X616 VSS G2.t20 SD2_1.t11 VSS.t276 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X617 SDn_2 SDn_2.t4 VSS.t573 VSS.t370 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X618 C32_U C32_U.t16 C32_D.t76 VSS.t86 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X619 Gc_1 IT.t80 SDc_1.t13 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X620 VSS SDn_2.t84 SDn_1.t18 VSS.t20 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X621 Gc_1 Gc_1.t52 Gc_2.t76 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X622 TG_0.IN b4b.t14 TG_0.IN VSS.t135 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X623 TG_1.IN.t40 TG_1.IN.t39 TG_1.IN.t40 VSS.t173 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X624 G1_2 ITAIL.t17 SD2_1.t4 VSS.t181 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X625 VDD SEL_L.t68 a_n2280_5855.t1 VDD.t163 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X626 OUT+ SEL_L.t69 TG_0.IN VSS.t346 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X627 G1_1 G1_2.t14 G1_2.t15 VDD.t240 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X628 TG_0.IN b5.t18 OUT5.t20 VSS.t127 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X629 IT G1_2.t31 SD1_1.t8 VDD.t236 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X630 OUT5 b5b.t18 TG_1.IN.t95 VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X631 OUT6 b6.t35 TG_0.IN VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X632 SDc_2 Gc_2.t124 VDD.t62 VDD.t61 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X633 OUT4 b4.t13 TG_0.IN VSS.t590 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X634 OUT4 b4b.t15 TG_1.IN.t106 VSS.t136 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X635 TG_1.IN.t140 b6.t36 TG_1.IN.t140 VSS.t4 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X636 TG_1.IN b5b.t19 OUT5.t36 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X637 Balance_Inverter_0.Inverter_0.OUT B4.t2 VDD.t123 VDD.t122 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X638 SD2_1 ITAIL.t18 G1_2.t2 VSS.t117 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X639 OUT+ a_n2265_3941.t39 TG_0.IN VDD.t337 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X640 TG_1.IN.t38 TG_1.IN.t37 TG_1.IN.t38 VSS.t175 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X641 TG_0.IN TG_0.IN TG_0.IN VSS.t356 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X642 TG_0.IN TG_0.IN TG_0.IN VSS.t324 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X643 TG_1.IN SEL_L.t70 OUT-.t6 VSS.t347 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X644 SD2_1 G2.t21 VSS.t273 VSS.t272 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X645 TG_0.IN a_n2265_3941.t40 OUT+.t77 VDD.t338 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X646 OUT+ a_n2265_3941.t41 TG_0.IN VDD.t339 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X647 TG_1.IN.t141 b6.t37 TG_1.IN.t141 VSS.t7 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X648 Gc_2 Gc_1.t80 Gc_1.t81 VDD.t61 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X649 OUT6 b6b.t34 TG_1.IN.t226 VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X650 VSS SDn_2.t85 SD3_1.t18 VSS.t23 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X651 VSS Balance_Inverter_1.Inverter_0.OUT b3.t0 VSS.t157 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X652 b6b B6.t1 VSS.t83 VSS.t82 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X653 Gc_2 Gc_2.t26 VDD.t71 VDD.t70 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X654 TG_0.IN b2b.t4 TG_0.IN VSS.t92 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X655 OUT- SEL_L.t71 TG_1.IN.t155 VSS.t202 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X656 OUT6 b6b.t35 TG_1.IN.t227 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X657 TG_0.IN SEL_L.t72 OUT+.t19 VSS.t203 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X658 OUT6 IT.t81 SD3_1.t8 VSS.t56 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X659 G1_1 G1_2.t12 G1_2.t13 VDD.t239 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X660 Gc_2 Gc_1.t78 Gc_1.t79 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X661 OUT6 b6b.t36 TG_1.IN.t228 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X662 TG_1.IN.t36 TG_1.IN.t35 TG_1.IN.t36 VSS.t170 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X663 TG_0.IN SEL_L.t73 OUT+.t18 VSS.t120 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X664 TG_1.IN.t34 TG_1.IN.t33 TG_1.IN.t34 VSS.t327 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X665 VSS G2.t1 G2.t2 VSS.t435 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X666 VSS SDn_2.t86 SD3_1.t17 VSS.t26 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X667 VSS SDn_2.t87 SDc_1.t42 VSS.t29 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X668 VSS SDn_2.t88 SDn_1.t17 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X669 SD3_1 SDn_2.t89 VSS.t36 VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X670 Gc_1 IT.t82 SDc_1.t12 VSS.t57 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X671 TG_1.IN.t261 b4.t14 TG_1.IN.t261 VSS.t589 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X672 TG_1.IN a_n2280_5855.t38 OUT-.t46 VDD.t203 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X673 OUT+ a_n2265_3941.t42 TG_0.IN VDD.t340 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X674 TG_0.IN a_n2265_3941.t43 OUT+.t55 VDD.t289 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X675 Gc_1 IT.t83 SDc_1.t11 VSS.t296 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X676 TG_1.IN.t101 b3.t7 TG_1.IN.t101 VSS.t94 nfet_03v3 ad=0.16p pd=1.64u as=0 ps=0 w=0.3u l=0.5u
X677 VSS SDn_2.t90 SDc_1.t41 VSS.t37 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X678 VSS SDn_2.t91 SDc_1.t40 VSS.t40 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X679 SD3_1 SDn_2.t92 VSS.t44 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X680 SD2_4 ITAIL.t19 OUT3.t3 VSS.t118 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X681 SDc_2 Gc_2.t126 VDD.t81 VDD.t80 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X682 Gc_1 IT.t84 SDc_1.t10 VSS.t297 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X683 Gc_1 IT.t85 SDc_1.t9 VSS.t298 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X684 TG_1.IN b6b.t37 OUT6.t84 VSS.t67 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X685 OUT3 b3b.t7 TG_1.IN.t2 VSS.t59 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X686 TG_1.IN a_n2280_5855.t39 OUT-.t45 VDD.t275 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X687 Gc_2 Gc_1.t76 Gc_1.t77 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X688 Gc_1 IT.t86 SDc_1.t8 VSS.t299 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X689 IT G1_2.t32 SD1_1.t7 VDD.t237 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X690 TG_1.IN SEL_L.t74 OUT-.t5 VSS.t121 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X691 VSS SDn_2.t93 SDc_1.t39 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X692 TG_0.IN TG_0.IN TG_0.IN VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X693 TG_0.IN a_n2265_3941.t44 OUT+.t56 VDD.t290 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X694 OUT4 ITAIL.t20 SD2_5.t4 VSS.t184 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X695 Gc_2 Gc_1.t74 Gc_1.t75 VDD.t82 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X696 Balance_Inverter_5.Inverter_0.OUT B6.t2 VSS.t462 VSS.t461 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X697 OUT+ SEL_L.t75 TG_0.IN VSS.t578 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X698 OUT3 b3.t8 TG_0.IN VSS.t95 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X699 OUT6 b6b.t38 TG_1.IN.t230 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X700 TG_0.IN b1b.t4 TG_0.IN VSS.t316 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X701 SDc_2 Gc_2.t127 VDD.t83 VDD.t82 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X702 VSS SEL_L.t76 a_n2280_5855.t10 VSS.t579 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X703 OUT- a_n2280_5855.t40 TG_1.IN.t194 VDD.t276 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X704 TG_1.IN.t133 b5.t19 TG_1.IN.t133 VSS.t139 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X705 OUT- a_n2280_5855.t41 TG_1.IN.t193 VDD.t277 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X706 Gc_2 Gc_2.t24 VDD.t69 VDD.t68 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X707 VSS SEL_L.t78 a_n2280_5855.t9 VSS.t348 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X708 SDc_2 Gc_1.t129 C32_U.t75 VDD.t68 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X709 VDD Gc_2.t22 Gc_2.t23 VDD.t31 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X710 OUT- SEL_L.t79 TG_1.IN.t153 VSS.t382 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X711 Gc_1 IT.t87 SDc_1.t7 VSS.t300 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X712 OUT- a_n2280_5855.t42 TG_1.IN.t192 VDD.t278 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X713 SD3_1 IT.t88 OUT6.t16 VSS.t301 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X714 VSS SDn_2.t94 SDn_1.t16 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X715 TG_0.IN SEL_L.t80 OUT+.t16 VSS.t371 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X716 VSS SDn_2.t95 SD3_1.t14 VSS.t310 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X717 TG_1.IN.t116 b2.t5 TG_1.IN.t116 VSS.t155 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X718 Gc_1 Gc_1.t50 Gc_2.t71 VDD.t22 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X719 OUT- a_n2280_5855.t43 TG_1.IN.t191 VDD.t196 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X720 OUT+ SEL_L.t81 TG_0.IN VSS.t409 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X721 VSS Balance_Inverter_3.Inverter_0.OUT b1.t1 VSS.t388 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X722 VSS SDn_2.t96 SDc_1.t38 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X723 OUT+ a_n2265_3941.t45 TG_0.IN VDD.t291 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X724 Gc_2 Gc_2.t20 VDD.t65 VDD.t64 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X725 TG_1.IN.t142 b6.t38 TG_1.IN.t142 VSS.t69 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X726 Balance_Inverter_4.Inverter_0.OUT B5.t2 VDD.t45 VDD.t44 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X727 OUT6 b6b.t39 TG_1.IN.t231 VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X728 TG_0.IN b4.t15 OUT4.t22 VSS.t134 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X729 Gc_2 Gc_1.t72 Gc_1.t73 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X730 OUT- a_n2280_5855.t44 TG_1.IN.t190 VDD.t197 pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.28u
X731 TG_0.IN b5.t20 OUT5.t25 VSS.t152 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X732 OUT5 IT.t89 SDn_1.t3 VSS.t302 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X733 TG_1.IN.t32 TG_1.IN.t31 TG_1.IN.t32 VSS.t326 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X734 SD3_1 IT.t90 OUT6.t15 VSS.t303 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X735 TG_0.IN TG_0.IN TG_0.IN VSS.t92 nfet_03v3 ad=0 pd=0 as=94.8f ps=0.92u w=0.3u l=0.5u
X736 VDD SEL_L.t82 a_n2265_3941.t0 VDD.t158 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X737 Gc_2 Gc_2.t18 VDD.t63 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X738 TG_1.IN SEL_L.t83 OUT-.t4 VSS.t398 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X739 TG_1.IN b5b.t20 OUT5.t35 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X740 TG_1.IN b5b.t21 OUT5.t34 VSS.t127 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X741 OUT6 b6.t39 TG_0.IN VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X742 TG_1.IN a_n2280_5855.t45 OUT-.t44 VDD.t198 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X743 SD2_4 G2.t22 VSS.t275 VSS.t274 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X744 OUT6 b6b.t40 TG_1.IN.t232 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X745 Balance_Inverter_2.Inverter_0.OUT B2.t2 VDD.t128 VDD.t127 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X746 TG_1.IN SEL_L.t85 OUT-.t3 VSS.t391 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X747 TG_0.IN b3.t9 OUT3.t6 VSS.t89 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X748 C32_D C32_U.t40 C32_U.t41 VSS.t218 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X749 TG_0.IN b5.t21 OUT5.t26 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X750 TG_0.IN b4.t16 OUT4.t23 VSS.t126 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X751 TG_0.IN TG_0.IN TG_0.IN VSS.t173 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X752 TG_1.IN SEL_L.t86 OUT-.t2 VSS.t392 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X753 TG_0.IN b5b.t22 TG_0.IN VSS.t151 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X754 OUT+ SEL_L.t87 TG_0.IN VSS.t459 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X755 TG_0.IN SEL_L.t88 OUT+.t13 VSS.t460 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X756 OUT6 IT.t91 SD3_1.t61 VSS.t540 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X757 TG_1.IN.t247 b5.t22 TG_1.IN.t247 VSS.t318 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X758 TG_0.IN TG_0.IN TG_0.IN VSS.t173 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X759 TG_0.IN b6.t40 OUT6.t48 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X760 OUT6 b6b.t41 TG_1.IN.t233 VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X761 VSS C32_D.t22 C32_D.t23 VSS.t163 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X762 C32_U C32_U.t14 C32_D.t74 VSS.t215 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X763 Gc_2 Gc_2.t16 VDD.t269 VDD.t0 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X764 OUT6 b6b.t42 TG_1.IN.t234 VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X765 SD2_5 ITAIL.t21 OUT4.t14 VSS.t328 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X766 TG_1.IN a_n2280_5855.t46 OUT-.t43 VDD.t199 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X767 IT IT.t4 SDn_2.t18 VSS.t366 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X768 VSS C32_D.t20 C32_D.t21 VSS.t162 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X769 C32_D C32_D.t18 VSS.t219 VSS.t218 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X770 Gc_1 Gc_1.t48 Gc_2.t69 VDD.t72 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X771 TG_1.IN a_n2280_5855.t47 OUT-.t42 VDD.t152 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X772 TG_0.IN TG_0.IN TG_0.IN VSS.t357 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X773 TG_0.IN b5b.t23 TG_0.IN VSS.t463 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X774 OUT6 IT.t93 SD3_1.t62 VSS.t481 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X775 TG_0.IN b5b.t24 TG_0.IN VSS.t93 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X776 VDD Gc_2.t132 SDc_2.t6 VDD.t72 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X777 OUT4 b4.t17 TG_0.IN VSS.t136 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X778 VDD Gc_2.t14 Gc_2.t15 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X779 VSS SDn_2.t2 SDn_2.t3 VSS.t368 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X780 TG_1.IN.t236 b6.t41 TG_1.IN.t236 VSS.t70 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X781 TG_0.IN TG_0.IN TG_0.IN VSS.t180 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X782 SD3_1 SDn_2.t97 VSS.t525 VSS.t524 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X783 SD3_1 SDn_2.t98 VSS.t526 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X784 OUT4 b4b.t16 TG_1.IN.t107 VSS.t137 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X785 C32_D C32_U.t38 C32_U.t39 VSS.t213 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X786 C32_U Gc_1.t132 SDc_2.t51 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X787 SDc_1 SDn_2.t99 VSS.t527 VSS.t375 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X788 VSS SDn_2.t100 SDc_1.t36 VSS.t57 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X789 C32_D C32_U.t36 C32_U.t37 VSS.t236 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X790 C32_U C32_U.t10 C32_D.t71 VSS.t163 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X791 VSS C32_D.t16 C32_D.t17 VSS.t215 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X792 TG_0.IN b6.t42 OUT6.t47 VSS.t67 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X793 TG_1.IN.t30 TG_1.IN.t29 TG_1.IN.t30 VSS.t167 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X794 C32_U C32_U.t8 C32_D.t70 VSS.t162 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X795 OUT- SEL_L.t89 TG_1.IN.t149 VSS.t396 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X796 SDc_1 IT.t94 Gc_1.t19 VSS.t518 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X797 Gc_1 IT.t95 SDc_1.t5 VSS.t37 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X798 Gc_1 IT.t96 SDc_1.t4 VSS.t40 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X799 OUT- SEL_L.t90 TG_1.IN.t148 VSS.t397 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X800 TG_1.IN.t28 TG_1.IN.t27 TG_1.IN.t28 VSS.t321 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X801 VDD G1_1.t2 G1_1.t3 VDD.t119 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X802 VDD b2b.t5 b2.t0 VDD.t245 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X803 TG_1.IN.t26 TG_1.IN.t25 TG_1.IN.t26 VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X804 VSS G2.t23 SD2_1.t9 VSS.t276 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X805 SDc_2 Gc_1.t133 C32_U.t73 VDD.t64 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X806 SDc_1 SDn_2.t101 VSS.t530 VSS.t378 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X807 VSS SDn_2.t102 SDc_1.t34 VSS.t299 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X808 SD3_1 SDn_2.t103 VSS.t534 VSS.t533 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X809 TG_0.IN TG_0.IN TG_0.IN VSS.t178 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X810 OUT5 b5.t23 TG_0.IN VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X811 OUT- SEL_L.t91 TG_1.IN.t147 VSS.t192 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X812 TG_1.IN b3b.t8 OUT3.t1 VSS.t60 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X813 VDD G1_1.t32 SD1_1.t3 VDD.t228 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X814 C32_D C32_D.t14 VSS.t214 VSS.t213 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X815 TG_0.IN a_n2265_3941.t46 OUT+.t58 VDD.t292 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X816 TG_0.IN b5.t24 OUT5.t31 VSS.t152 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X817 VSS C32_D.t12 C32_D.t13 VSS.t238 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X818 C32_D C32_D.t10 VSS.t237 VSS.t236 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X819 Gc_2 Gc_2.t12 VDD.t266 VDD.t61 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X820 OUT- a_n2280_5855.t48 TG_1.IN.t186 VDD.t153 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X821 OUT5 b5b.t25 TG_1.IN.t248 VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X822 VSS SDn_2.t104 SD3_1.t10 VSS.t535 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X823 C32_U C32_U.t6 C32_D.t69 VSS.t231 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X824 TG_1.IN.t97 b3.t10 TG_1.IN.t97 VSS.t90 nfet_03v3 ad=94.8f pd=0.92u as=0 ps=0 w=0.3u l=0.5u
X825 G1_2 G1_2.t18 G1_1.t18 VDD.t225 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X826 SDc_2 Gc_1.t134 C32_U.t72 VDD.t61 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X827 TG_1.IN b5b.t26 OUT5.t32 VSS.t97 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X828 C32_D C32_D.t8 VSS.t235 VSS.t234 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X829 SD2_1 ITAIL.t22 G1_2.t1 VSS.t117 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X830 Gc_2 Gc_1.t70 Gc_1.t71 VDD.t70 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X831 SDc_2 Gc_2.t134 VDD.t86 VDD.t70 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X832 G1_1 G1_2.t10 G1_2.t11 VDD.t210 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X833 OUT2 b2b.t6 TG_1.IN.t135 VSS.t317 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X834 SD2_1 G2.t24 VSS.t444 VSS.t272 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X835 Gc_2 Gc_2.t10 VDD.t265 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X836 VSS SEL_L.t92 a_n2265_3941.t10 VSS.t193 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X837 TG_1.IN.t259 b4.t18 TG_1.IN.t259 VSS.t440 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X838 C32_D C32_U.t34 C32_U.t35 VSS.t426 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X839 C32_U C32_U.t4 C32_D.t67 VSS.t238 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X840 SDc_2 Gc_1.t135 C32_U.t71 VDD.t10 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X841 VDD b6b.t43 b6.t0 VDD.t221 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X842 TG_1.IN SEL_L.t93 OUT-.t1 VSS.t414 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X843 C32_U C32_U.t2 C32_D.t66 VSS.t189 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X844 VSS C32_D.t6 C32_D.t7 VSS.t231 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X845 OUT+ a_n2265_3941.t47 TG_0.IN VDD.t293 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X846 TG_1.IN.t237 b6.t43 TG_1.IN.t237 VSS.t8 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X847 SDn_2 IT.t2 IT.t3 VSS.t365 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X848 C32_D C32_U.t32 C32_U.t33 VSS.t234 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X849 SDc_1 IT.t97 Gc_1.t18 VSS.t510 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X850 TG_1.IN a_n2280_5855.t49 OUT-.t41 VDD.t154 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X851 OUT+ a_n2265_3941.t48 TG_0.IN VDD.t294 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X852 VSS SEL_L.t94 a_n2265_3941.t9 VSS.t415 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.28u
X853 TG_0.IN b6b.t44 TG_0.IN VSS.t279 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X854 TG_1.IN.t24 TG_1.IN.t23 TG_1.IN.t24 VSS.t325 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X855 VDD Gc_2.t8 Gc_2.t9 VDD.t12 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X856 TG_0.IN TG_0.IN TG_0.IN VSS.t167 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X857 OUT+ SEL_L.t95 TG_0.IN VSS.t454 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X858 G1_1 G1_1.t0 VDD.t212 VDD.t211 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X859 TG_1.IN.t22 TG_1.IN.t21 TG_1.IN.t22 VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X860 TG_1.IN.t20 TG_1.IN.t19 TG_1.IN.t20 VSS.t167 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X861 TG_1.IN SEL_L.t96 OUT-.t0 VSS.t455 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X862 OUT+ a_n2265_3941.t49 TG_0.IN VDD.t137 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X863 OUT5 b5.t25 TG_0.IN VSS.t96 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X864 C32_U Gc_1.t136 SDc_2.t50 VDD.t12 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X865 TG_0.IN b6b.t45 TG_0.IN VSS.t3 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X866 C32_D C32_D.t4 VSS.t427 VSS.t426 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X867 b6b b6.t44 VDD.t242 VDD.t241 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X868 OUT6 IT.t98 SD3_1.t63 VSS.t23 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X869 Balance_Inverter_1.Inverter_0.OUT B3.t1 VSS.t63 VSS.t62 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X870 TG_1.IN.t238 b6.t45 TG_1.IN.t238 VSS.t84 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X871 C32_D C32_D.t2 VSS.t425 VSS.t165 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X872 VSS C32_D.t0 C32_D.t1 VSS.t189 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X873 VSS G2.t25 SD2_2.t1 VSS.t435 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X874 Gc_2 Gc_2.t6 VDD.t25 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X875 TG_1.IN b4b.t17 OUT4.t0 VSS.t138 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X876 TG_0.IN TG_0.IN TG_0.IN VSS.t172 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X877 SDc_2 Gc_1.t137 C32_U.t69 VDD.t8 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X878 SDc_2 Gc_1.t138 C32_U.t68 VDD.t46 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X879 TG_0.IN TG_0.IN TG_0.IN VSS.t356 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X880 IT IT.t0 SDn_2.t16 VSS.t364 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X881 TG_1.IN.t124 b1.t4 TG_1.IN.t124 VSS.t154 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X882 SDc_2 Gc_2.t137 VDD.t88 VDD.t87 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X883 TG_1.IN.t18 TG_1.IN.t17 TG_1.IN.t18 VSS.t168 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X884 TG_0.IN SEL_L.t97 OUT+.t11 VSS.t403 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X885 OUT6 IT.t100 SD3_1.t48 VSS.t373 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X886 TG_0.IN b6b.t46 TG_0.IN VSS.t4 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X887 TG_0.IN a_n2265_3941.t50 OUT+.t7 VDD.t138 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X888 SDn_1 IT.t101 OUT5.t5 VSS.t374 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X889 SD1_1 G1_1.t34 VDD.t232 VDD.t231 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X890 SD2_4 ITAIL.t23 OUT3.t2 VSS.t118 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X891 TG_1.IN b6b.t47 OUT6.t0 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X892 TG_1.IN a_n2280_5855.t50 OUT-.t40 VDD.t155 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X893 C32_D C32_U.t30 C32_U.t31 VSS.t165 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X894 IT G1_2.t34 SD1_1.t6 VDD.t238 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X895 TG_0.IN SEL_L.t99 OUT+.t10 VSS.t379 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X896 TG_0.IN TG_0.IN TG_0.IN VSS.t178 nfet_03v3 ad=0.156p pd=1.12u as=0 ps=0 w=0.6u l=0.5u
X897 VDD Gc_2.t138 SDc_2.t3 VDD.t89 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X898 TG_1.IN b6b.t48 OUT6.t1 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X899 SD3_1 IT.t102 OUT6.t10 VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X900 SD2_1 ITAIL.t24 G1_2.t0 VSS.t119 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X901 OUT6 b6.t46 TG_0.IN VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X902 C32_U Gc_1.t139 SDc_2.t49 VDD.t31 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X903 VSS SDn_2.t105 SDc_1.t33 VSS.t513 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X904 OUT2 b2.t6 TG_0.IN VSS.t156 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X905 b3b B3.t2 VSS.t65 VSS.t64 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X906 Gc_2 Gc_1.t68 Gc_1.t69 VDD.t80 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X907 OUT6 b6.t47 TG_0.IN VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X908 TG_0.IN b3b.t9 TG_0.IN VSS.t61 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X909 TG_0.IN b6b.t49 TG_0.IN VSS.t7 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X910 TG_0.IN b6.t48 OUT6.t44 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X911 TG_0.IN b6.t49 OUT6.t43 VSS.t67 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X912 Gc_1 Gc_1.t46 Gc_2.t66 VDD.t31 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X913 OUT- a_n2280_5855.t51 TG_1.IN.t183 VDD.t311 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X914 VDD Gc_2.t139 SDc_2.t2 VDD.t31 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X915 TG_1.IN.t16 TG_1.IN.t15 TG_1.IN.t16 VSS.t180 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X916 TG_1.IN.t14 TG_1.IN.t13 TG_1.IN.t14 VSS.t166 nfet_03v3 ad=0 pd=0 as=0.264p ps=2.08u w=0.6u l=0.5u
X917 VDD Gc_2.t4 Gc_2.t5 VDD.t22 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X918 OUT- SEL_L.t101 TG_1.IN.t144 VSS.t412 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X919 OUT5 IT.t103 SDn_1.t1 VSS.t20 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X920 SDc_2 Gc_1.t141 C32_U.t66 VDD.t101 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X921 Gc_2 Gc_1.t66 Gc_1.t67 VDD.t64 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X922 TG_0.IN a_n2265_3941.t51 OUT+.t8 VDD.t139 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X923 TG_0.IN b4b.t18 TG_0.IN VSS.t222 nfet_03v3 ad=0 pd=0 as=0.16p ps=1.64u w=0.3u l=0.5u
X924 TG_1.IN.t12 TG_1.IN.t11 TG_1.IN.t12 VSS.t179 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X925 C32_U Gc_1.t142 SDc_2.t48 VDD.t22 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X926 SDc_2 Gc_2.t140 VDD.t94 VDD.t64 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X927 OUT6 b6.t50 TG_0.IN VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X928 VSS SDn_2.t106 SD3_1.t9 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X929 OUT5 b5.t26 TG_0.IN VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X930 Gc_2 Gc_2.t2 VDD.t21 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X931 SDc_1 IT.t104 Gc_1.t17 VSS.t375 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X932 OUT- SEL_L.t102 TG_1.IN.t143 VSS.t413 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X933 OUT5 IT.t105 SDn_1.t0 VSS.t376 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X934 G1_2 G1_2.t8 G1_1.t16 VDD.t209 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X935 SDc_2 Gc_1.t143 C32_U.t64 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X936 VDD G1_1.t35 SD1_1.t5 VDD.t233 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X937 Gc_2 Gc_2.t0 VDD.t19 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X938 SDc_1 IT.t106 Gc_1.t16 VSS.t377 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X939 SDc_1 SDn_2.t107 VSS.t519 VSS.t518 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X940 OUT3 b3b.t10 TG_1.IN.t262 VSS.t59 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X941 Gc_2 Gc_1.t64 Gc_1.t65 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X942 TG_0.IN b6b.t50 TG_0.IN VSS.t8 nfet_03v3 ad=0 pd=0 as=0.156p ps=1.12u w=0.6u l=0.5u
X943 SDc_2 Gc_2.t143 VDD.t33 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X944 SDc_1 IT.t107 Gc_1.t15 VSS.t378 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X945 OUT+ SEL_L.t103 TG_0.IN VSS.t450 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X946 VSS SDn_2.t0 SDn_2.t1 VSS.t366 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
R0 VSS.t262 VSS.n1639 2045.19
R1 VSS.t64 VSS.n1641 2003.92
R2 VSS.t319 VSS.n1645 2003.92
R3 VSS.n1711 VSS.n1565 1938.34
R4 VSS.n1711 VSS 1757.65
R5 VSS VSS.n1711 1677.99
R6 VSS.n1711 VSS 1677.99
R7 VSS.n1563 VSS.t456 1561.78
R8 VSS.n1565 VSS.t157 1530.27
R9 VSS.n1562 VSS.t388 1530.27
R10 VSS.n426 VSS.n425 1447.46
R11 VSS.n1564 VSS.n1563 1436.69
R12 VSS.n1564 VSS.n1562 1407.7
R13 VSS.n1646 VSS.t262 1070.94
R14 VSS.n1646 VSS.t64 1049.33
R15 VSS.n1646 VSS.t319 1049.33
R16 VSS.n469 VSS.t412 335.526
R17 VSS.n478 VSS.t455 322.368
R18 VSS.n535 VSS.t418 319.079
R19 VSS.n511 VSS.t343 289.474
R20 VSS.n523 VSS.t402 289.474
R21 VSS.n490 VSS.t337 286.185
R22 VSS.n502 VSS.t434 286.185
R23 VSS.n457 VSS.t201 273.026
R24 VSS.n1711 VSS.n1564 268.024
R25 VSS.n457 VSS.t401 253.29
R26 VSS.n434 VSS.t579 252.085
R27 VSS.n490 VSS.t331 240.132
R28 VSS.n502 VSS.t81 240.132
R29 VSS.n511 VSS.t408 236.843
R30 VSS.n523 VSS.t451 236.843
R31 VSS.n535 VSS.t429 207.238
R32 VSS.n1432 VSS.t322 205.987
R33 VSS.n478 VSS.t335 203.947
R34 VSS.n1407 VSS.t207 198.357
R35 VSS.n1418 VSS.t164 198.357
R36 VSS.n469 VSS.t198 190.79
R37 VSS.n481 VSS.t397 190.79
R38 VSS.n1407 VSS.t236 190.728
R39 VSS.n1418 VSS.t140 190.728
R40 VSS.n532 VSS.t392 187.5
R41 VSS.n544 VSS.t395 187.5
R42 VSS.n1432 VSS.t227 183.1
R43 VSS.n434 VSS.t399 181.611
R44 VSS.n514 VSS.t340 157.895
R45 VSS.n526 VSS.t448 157.895
R46 VSS.n1429 VSS.t231 156.398
R47 VSS.n499 VSS.t411 154.606
R48 VSS.n1130 VSS.t99 148.899
R49 VSS.n1408 VSS.t210 148.768
R50 VSS.n1417 VSS.t174 148.768
R51 VSS.n1306 VSS.t582 146.244
R52 VSS.n438 VSS.t104 143.661
R53 VSS.n1128 VSS.n1127 143.173
R54 VSS.n1139 VSS.t254 143.173
R55 VSS.n460 VSS.t347 141.447
R56 VSS.n1406 VSS.t162 141.139
R57 VSS.n1421 VSS.t163 141.139
R58 VSS.t297 VSS.n1519 140.565
R59 VSS.n1143 VSS.n1142 138.877
R60 VSS.n1122 VSS.t51 137.446
R61 VSS.n1144 VSS.t593 137.446
R62 VSS.n1555 VSS.n1554 136.013
R63 VSS.n1433 VSS.t225 133.51
R64 VSS.n1509 VSS.t37 124.677
R65 VSS.n454 VSS.t79 121.712
R66 VSS.n466 VSS.t431 121.712
R67 VSS.n1440 VSS.t292 114.438
R68 VSS.n1300 VSS.t16 110.291
R69 VSS.n493 VSS.t398 108.553
R70 VSS.n505 VSS.t382 108.553
R71 VSS.t299 VSS.n1558 107.379
R72 VSS.n1428 VSS.t426 106.808
R73 VSS.n1530 VSS.t549 105.948
R74 VSS.n1138 VSS.t300 105.948
R75 VSS.n520 VSS.t202 105.263
R76 VSS.n1120 VSS.t375 100.221
R77 VSS.n1546 VSS.t468 100.221
R78 VSS.n1411 VSS.t204 99.1789
R79 VSS.n1416 VSS.t86 99.1789
R80 VSS.n1403 VSS.t115 91.5498
R81 VSS.n1422 VSS.t213 91.5498
R82 VSS.t55 VSS.n1135 87.3353
R83 VSS.n1434 VSS.t189 83.9207
R84 VSS.t129 VSS.t518 83.0401
R85 VSS.n1299 VSS.t57 79.1226
R86 VSS.n538 VSS.t383 75.6584
R87 VSS.n1656 VSS.n1655 73.6511
R88 VSS.n432 VSS.t348 73.1865
R89 VSS.n475 VSS.t196 72.3689
R90 VSS.n487 VSS.t433 72.3689
R91 VSS.n1544 VSS.t187 71.5864
R92 VSS.n1448 VSS.t165 70.5698
R93 VSS.n1532 VSS.t378 68.723
R94 VSS.n1137 VSS.t9 68.723
R95 VSS.n1439 VSS.t290 64.8479
R96 VSS.n1660 VSS.t106 64.2774
R97 VSS.n1118 VSS.t259 62.9961
R98 VSS.n1549 VSS.t298 62.9961
R99 VSS.n1512 VSS.t82 61.0534
R100 VSS.n1528 VSS.t129 60.1327
R101 VSS.n472 VSS.t341 59.211
R102 VSS.n484 VSS.t414 59.211
R103 VSS.n1427 VSS.t147 57.2188
R104 VSS.t11 VSS.t365 56.0954
R105 VSS.n541 VSS.t338 55.9216
R106 VSS.n1647 VSS.n1646 55.0085
R107 VSS.n699 VSS.t177 52.9321
R108 VSS.n888 VSS.n887 52.1759
R109 VSS.n1105 VSS.t384 51.1145
R110 VSS.n690 VSS.t409 50.6636
R111 VSS.t82 VSS.t466 49.6947
R112 VSS.n1412 VSS.t218 49.5897
R113 VSS.n1413 VSS.t223 49.5897
R114 VSS.n335 VSS.t103 49.207
R115 VSS.n363 VSS.t10 49.0836
R116 VSS.n1296 VSS.t377 47.9533
R117 VSS.n657 VSS.t596 47.6389
R118 VSS.n398 VSS.t303 47.4036
R119 VSS.n41 VSS.t80 47.3306
R120 VSS.n319 VSS.t578 46.8828
R121 VSS.n1672 VSS.t74 46.6512
R122 VSS.n93 VSS.t386 45.0912
R123 VSS.n1667 VSS.t109 43.7093
R124 VSS.n1984 VSS.t15 42.7789
R125 VSS.n358 VSS.t336 42.0717
R126 VSS.n372 VSS.t481 42.0717
R127 VSS.t346 VSS.t52 42.0717
R128 VSS.n1667 VSS.t124 42.0282
R129 VSS.n1402 VSS.t102 41.9606
R130 VSS.n1423 VSS.t0 41.9606
R131 VSS.t495 VSS.t311 41.6227
R132 VSS.t302 VSS.t26 41.6227
R133 VSS.n294 VSS.t94 41.5896
R134 VSS.n80 VSS.t492 40.4665
R135 VSS.n1675 VSS.n1674 40.3471
R136 VSS.n297 VSS.t89 40.0773
R137 VSS.t58 VSS.t171 40.0773
R138 VSS.n1672 VSS.t272 39.0862
R139 VSS.t12 VSS.t334 38.5658
R140 VSS.n1010 VSS.t69 38.1825
R141 VSS.n628 VSS.t156 37.8088
R142 VSS.n1516 VSS.t309 36.9162
R143 VSS.n1959 VSS.t535 36.8128
R144 VSS.n678 VSS.t323 36.2965
R145 VSS.n1631 VSS.t328 36.241
R146 VSS.n90 VSS.t48 35.8418
R147 VSS.n1673 VSS.t117 35.724
R148 VSS.n1017 VSS.t85 35.5939
R149 VSS.n1851 VSS.t325 35.5939
R150 VSS.n991 VSS.t589 34.9467
R151 VSS.n1435 VSS.t234 34.3315
R152 VSS.n1911 VSS.t72 34.2996
R153 VSS.n38 VSS.t476 34.1833
R154 VSS.n982 VSS.t173 33.6524
R155 VSS.n1711 VSS.t304 33.6226
R156 VSS.n1655 VSS.t183 33.478
R157 VSS.n384 VSS.t364 33.3069
R158 VSS.t357 VSS.t134 33.2718
R159 VSS.n1883 VSS.t269 33.0053
R160 VSS.n1668 VSS.t266 32.7821
R161 VSS.n625 VSS.t460 32.5156
R162 VSS.n1023 VSS.t443 32.3581
R163 VSS.n622 VSS.t359 31.7595
R164 VSS.n1891 VSS.t128 31.711
R165 VSS.n1535 VSS.t513 31.4983
R166 VSS.n1136 VSS.t55 31.4983
R167 VSS.n1032 VSS.t166 31.0638
R168 VSS.n116 VSS.n115 31.0638
R169 VSS.n663 VSS.t175 31.0033
R170 VSS.n120 VSS.n119 30.4167
R171 VSS.n681 VSS.t92 30.2471
R172 VSS.n75 VSS.t54 30.061
R173 VSS.n1613 VSS.t435 29.4607
R174 VSS.n597 VSS.t403 28.9244
R175 VSS.n985 VSS.t133 28.4752
R176 VSS.n1647 VSS.n1635 28.4752
R177 VSS.n397 VSS.n396 28.3267
R178 VSS.n1671 VSS.t122 28.159
R179 VSS.n631 VSS.t394 27.9786
R180 VSS.n390 VSS.t56 27.7486
R181 VSS.t259 VSS.n1108 27.0903
R182 VSS.n87 VSS.t479 26.5925
R183 VSS.n1878 VSS.t88 26.5338
R184 VSS.n517 VSS.t121 26.3163
R185 VSS.n529 VSS.t396 26.3163
R186 VSS.n365 VSS.t524 26.295
R187 VSS.n1949 VSS.t344 26.295
R188 VSS.n1856 VSS.t98 25.8866
R189 VSS.n1894 VSS.t318 25.8866
R190 VSS.n1568 VSS.t18 25.7714
R191 VSS.n1115 VSS.t510 25.5575
R192 VSS.n1326 VSS.t238 24.7951
R193 VSS.t368 VSS.t453 24.542
R194 VSS.n1907 VSS.t184 23.298
R195 VSS.n496 VSS.t192 23.0268
R196 VSS.n508 VSS.t391 23.0268
R197 VSS.n1961 VSS.t53 22.7891
R198 VSS.n1663 VSS.t282 22.6954
R199 VSS.t222 VSS.t6 22.6508
R200 VSS.t181 VSS.t87 22.0037
R201 VSS.n702 VSS.t410 21.9293
R202 VSS.n1574 VSS.t40 21.8549
R203 VSS.n1669 VSS.t125 21.8549
R204 VSS.n1020 VSS.t179 21.3565
R205 VSS.t53 VSS.t380 21.0361
R206 VSS.n1014 VSS.n1013 20.7094
R207 VSS.n1646 VSS.t274 20.5066
R208 VSS.n36 VSS.t17 20.1596
R209 VSS.n558 VSS.t430 20.1596
R210 VSS.n1003 VSS.t4 20.0622
R211 VSS.n684 VSS.t126 19.6608
R212 VSS.n343 VSS.t14 19.2831
R213 VSS.n603 VSS.t342 19.2831
R214 VSS.n361 VSS.t454 19.2831
R215 VSS.n370 VSS.t247 19.2831
R216 VSS.n58 VSS.t370 19.2831
R217 VSS.t549 VSS.n1109 18.6128
R218 VSS.n687 VSS.t372 18.1485
R219 VSS.n1020 VSS.t67 18.1208
R220 VSS.n122 VSS.t97 18.1208
R221 VSS.n1635 VSS.t123 18.1208
R222 VSS.n1578 VSS.t503 17.6521
R223 VSS.n85 VSS.t302 17.3431
R224 VSS.n393 VSS.t301 17.3431
R225 VSS.n1035 VSS.t138 16.8265
R226 VSS.n640 VSS.t155 16.6361
R227 VSS.n643 VSS.t432 15.88
R228 VSS.n606 VSS.t339 15.7772
R229 VSS.n352 VSS.t12 15.7772
R230 VSS.n370 VSS.t19 15.7772
R231 VSS.n1241 VSS.n1240 15.5852
R232 VSS.t167 VSS.t168 15.5322
R233 VSS.t7 VSS.t180 15.5322
R234 VSS.t5 VSS.t70 15.5322
R235 VSS.n994 VSS.t68 15.5322
R236 VSS.t463 VSS.t170 15.5322
R237 VSS.t127 VSS.t139 15.5322
R238 VSS.n1886 VSS.t276 15.5322
R239 VSS.n1438 VSS.t116 15.2587
R240 VSS.n435 VSS.n433 14.975
R241 VSS.n555 VSS.t419 14.9007
R242 VSS.n1711 VSS.t264 14.7111
R243 VSS.n1711 VSS.t62 14.4262
R244 VSS.n1711 VSS.t77 14.4262
R245 VSS.t385 VSS.t345 14.0242
R246 VSS.n672 VSS.t362 13.6115
R247 VSS.n684 VSS.t315 13.6115
R248 VSS.n615 VSS.t452 13.6115
R249 VSS.n1003 VSS.t71 13.5907
R250 VSS.n1017 VSS.t279 13.5907
R251 VSS.n241 VSS.n239 13.5907
R252 VSS.n1844 VSS.t463 12.9436
R253 VSS.n660 VSS.t404 12.8553
R254 VSS.t590 VSS.t329 12.8553
R255 VSS.n391 VSS.t305 12.7184
R256 VSS.n245 VSS.t172 12.2964
R257 VSS.n48 VSS.t333 12.2713
R258 VSS.n379 VSS.t366 12.2713
R259 VSS.n68 VSS.t330 12.2713
R260 VSS.t95 VSS.t415 12.0991
R261 VSS.n1665 VSS.t118 11.7682
R262 VSS.n72 VSS.n71 11.5622
R263 VSS.n1554 VSS.n1139 11.4542
R264 VSS.n310 VSS.t60 11.343
R265 VSS.n666 VSS.t406 11.343
R266 VSS.t84 VSS.t222 11.0021
R267 VSS.n1010 VSS.t66 11.0021
R268 VSS.n1867 VSS.t96 11.0021
R269 VSS.t304 VSS.n1710 10.9277
R270 VSS.n381 VSS.t371 10.5183
R271 VSS.n1859 VSS.t127 10.3549
R272 VSS.n451 VSS.t332 9.86892
R273 VSS.n463 VSS.t413 9.86892
R274 VSS.n705 VSS.t393 9.83065
R275 VSS.n1836 VSS.t178 9.70779
R276 VSS.t32 VSS.t385 9.64182
R277 VSS.t17 VSS.t310 9.64182
R278 VSS.t476 VSS.t313 9.64182
R279 VSS.t524 VSS.t497 9.64182
R280 VSS.t540 VSS.t374 9.64182
R281 VSS.n1638 VSS.t263 9.48597
R282 VSS.n1640 VSS.t65 9.48597
R283 VSS.n1644 VSS.t320 9.48597
R284 VSS.n1149 VSS.t188 9.33385
R285 VSS.n1734 VSS.t83 9.33385
R286 VSS.n1729 VSS.t130 9.33385
R287 VSS.n1637 VSS.n1636 9.32914
R288 VSS.n1561 VSS.n1560 9.32914
R289 VSS.n1557 VSS.n1147 9.32914
R290 VSS.n1732 VSS.n1106 9.32914
R291 VSS.n1727 VSS.n1110 9.32914
R292 VSS.n1643 VSS.n1642 9.32914
R293 VSS.n675 VSS.t169 9.07449
R294 VSS.n699 VSS.t321 9.07449
R295 VSS.n104 VSS.t120 9.07449
R296 VSS.n976 VSS.t7 9.06064
R297 VSS.n979 VSS.t326 9.06064
R298 VSS.n988 VSS.t5 9.06064
R299 VSS.n1870 VSS.t150 9.06064
R300 VSS.n1566 VSS.t265 8.96939
R301 VSS.n1712 VSS.t63 8.96939
R302 VSS.n1730 VSS.t462 8.96939
R303 VSS.n1148 VSS.t132 8.96939
R304 VSS.n1714 VSS.t186 8.96939
R305 VSS.n1567 VSS.t78 8.96939
R306 VSS.n1935 VSS.t199 8.76533
R307 VSS.n1955 VSS.t367 8.76533
R308 VSS.n1957 VSS.t346 8.76533
R309 VSS.n1964 VSS.t249 8.76533
R310 VSS.n303 VSS.t442 8.31832
R311 VSS.n656 VSS.t95 8.31832
R312 VSS.t193 VSS.t441 8.31832
R313 VSS.n1013 VSS.t360 8.31832
R314 VSS.n82 VSS.t495 8.09371
R315 VSS.n1933 VSS.t20 7.88885
R316 VSS.n1029 VSS.t136 7.76633
R317 VSS.n1994 VSS.t509 7.64137
R318 VSS.n1401 VSS.t145 7.62961
R319 VSS.n1424 VSS.t114 7.62961
R320 VSS.t404 VSS.t90 7.56216
R321 VSS.t323 VSS.t176 7.56216
R322 VSS.t126 VSS.t327 7.56216
R323 VSS.t315 VSS.t316 7.56216
R324 VSS.t372 VSS.t590 7.56216
R325 VSS.t134 VSS.t295 7.56216
R326 VSS.n696 VSS.t160 7.56216
R327 VSS VSS.n1108 7.19973
R328 VSS.n1170 VSS.n1169 7.19342
R329 VSS.n240 VSS.t111 7.11918
R330 VSS.n1601 VSS.n1600 7.09117
R331 VSS.n349 VSS.t35 7.01237
R332 VSS.n567 VSS.t449 7.01237
R333 VSS.n73 VSS.n72 6.93753
R334 VSS.n1985 VSS.n1984 6.93753
R335 VSS.n27 VSS.n26 6.51634
R336 VSS.n1026 VSS.t8 6.47203
R337 VSS.n1604 VSS.t586 6.41395
R338 VSS.n1971 VSS.t507 6.41267
R339 VSS.n1932 VSS.n103 6.41267
R340 VSS.n1951 VSS.t568 6.41267
R341 VSS.n1954 VSS.n100 6.41267
R342 VSS.n1972 VSS.n97 6.41267
R343 VSS.n1993 VSS.t539 6.41267
R344 VSS.n1391 VSS.n1390 6.37382
R345 VSS.n1168 VSS.n1167 6.36926
R346 VSS.n1973 VSS.t376 6.35945
R347 VSS.n1443 VSS.t425 6.35593
R348 VSS.n1595 VSS.t504 6.35232
R349 VSS.n1601 VSS.t285 6.26682
R350 VSS.n594 VSS.t428 6.13588
R351 VSS.n1935 VSS.t387 6.13588
R352 VSS.n34 VSS.t32 6.13588
R353 VSS.n1928 VSS.n111 5.89743
R354 VSS.n1628 VSS.n1627 5.8805
R355 VSS.n1630 VSS.n1629 5.8805
R356 VSS.n1602 VSS.n1599 5.8805
R357 VSS.n1603 VSS.n1598 5.8805
R358 VSS.n1604 VSS.t275 5.8805
R359 VSS.n1875 VSS.t181 5.82487
R360 VSS.n1132 VSS.t314 5.72737
R361 VSS.n1651 VSS.t182 5.35691
R362 VSS.n300 VSS.t59 5.29366
R363 VSS.n651 VSS.t356 5.29366
R364 VSS.n38 VSS.t379 5.2594
R365 VSS.n1957 VSS.t369 5.2594
R366 VSS.n56 VSS.t368 5.2594
R367 VSS.n61 VSS.t459 5.2594
R368 VSS.n1966 VSS.t533 5.2594
R369 VSS.n66 VSS.t23 5.2594
R370 VSS.n1639 VSS.n1638 5.2005
R371 VSS.n1641 VSS.n1640 5.2005
R372 VSS.n1513 VSS.n1512 5.2005
R373 VSS.n1515 VSS.n1514 5.2005
R374 VSS.n1517 VSS.n1516 5.2005
R375 VSS.n1520 VSS.t297 5.2005
R376 VSS.n1522 VSS.n1521 5.2005
R377 VSS.n1733 VSS.n1105 5.2005
R378 VSS.n1116 VSS.n1115 5.2005
R379 VSS.n1307 VSS.n1306 5.2005
R380 VSS.n1308 VSS.n1305 5.2005
R381 VSS.n1309 VSS.n1304 5.2005
R382 VSS.n1311 VSS.n1301 5.2005
R383 VSS.n1645 VSS.n1644 5.2005
R384 VSS.n1614 VSS.n1613 5.2005
R385 VSS.n1135 VSS 5.2005
R386 VSS VSS.n1558 5.2005
R387 VSS.n1556 VSS.n1555 5.2005
R388 VSS.n1728 VSS.n1109 5.2005
R389 VSS.n1589 VSS.t299 5.2005
R390 VSS.n1146 VSS.n1145 5.2005
R391 VSS.n1717 VSS.n1144 5.2005
R392 VSS.n1718 VSS.n1143 5.2005
R393 VSS VSS.n1139 5.2005
R394 VSS.n1720 VSS.n1138 5.2005
R395 VSS.n1721 VSS.n1137 5.2005
R396 VSS.n1722 VSS.n1136 5.2005
R397 VSS.n1724 VSS.n1132 5.2005
R398 VSS.n1131 VSS.n1130 5.2005
R399 VSS.n1129 VSS.n1128 5.2005
R400 VSS.n1126 VSS.n1125 5.2005
R401 VSS.n1123 VSS.n1122 5.2005
R402 VSS.n1121 VSS.n1120 5.2005
R403 VSS.n1119 VSS.n1118 5.2005
R404 VSS.n1524 VSS.n1523 5.2005
R405 VSS.n1526 VSS.n1525 5.2005
R406 VSS.n1529 VSS.n1528 5.2005
R407 VSS.n1531 VSS.n1530 5.2005
R408 VSS.n1533 VSS.n1532 5.2005
R409 VSS.n1536 VSS.n1535 5.2005
R410 VSS.n1538 VSS.n1537 5.2005
R411 VSS.n1540 VSS.n1539 5.2005
R412 VSS.n1542 VSS.n1541 5.2005
R413 VSS.n1545 VSS.n1544 5.2005
R414 VSS.n1554 VSS.n1553 5.2005
R415 VSS.n1552 VSS.n1546 5.2005
R416 VSS.n1550 VSS.n1549 5.2005
R417 VSS.n1569 VSS.n1568 5.2005
R418 VSS.n1571 VSS.n1570 5.2005
R419 VSS.n1702 VSS.n1700 5.2005
R420 VSS.n1709 VSS.n1708 5.2005
R421 VSS.n1706 VSS.n1575 5.2005
R422 VSS.n1702 VSS.n1579 5.2005
R423 VSS.n1597 VSS.n1596 5.2005
R424 VSS.n1327 VSS.n1326 5.2005
R425 VSS.n1349 VSS.n1347 5.2005
R426 VSS.n1451 VSS.n1449 5.2005
R427 VSS.n1400 VSS.n1398 5.2005
R428 VSS.n1400 VSS.n1397 5.2005
R429 VSS.n1486 VSS.n1401 5.2005
R430 VSS.n1485 VSS.n1402 5.2005
R431 VSS.n1484 VSS.n1403 5.2005
R432 VSS.n1482 VSS.n1406 5.2005
R433 VSS.n1481 VSS.n1407 5.2005
R434 VSS.n1480 VSS.n1408 5.2005
R435 VSS.n1478 VSS.n1411 5.2005
R436 VSS.n1477 VSS.n1412 5.2005
R437 VSS.n1476 VSS.t215 5.2005
R438 VSS.n1475 VSS.n1413 5.2005
R439 VSS.n1473 VSS.n1416 5.2005
R440 VSS.n1472 VSS.n1417 5.2005
R441 VSS.n1471 VSS.n1418 5.2005
R442 VSS.n1469 VSS.n1421 5.2005
R443 VSS.n1468 VSS.n1422 5.2005
R444 VSS.n1467 VSS.n1423 5.2005
R445 VSS.n1466 VSS.n1424 5.2005
R446 VSS.n1464 VSS.n1427 5.2005
R447 VSS.n1463 VSS.n1428 5.2005
R448 VSS.n1462 VSS.n1429 5.2005
R449 VSS.n1460 VSS.n1432 5.2005
R450 VSS.n1459 VSS.n1433 5.2005
R451 VSS.n1458 VSS.n1434 5.2005
R452 VSS.n1457 VSS.n1435 5.2005
R453 VSS.n1455 VSS.n1438 5.2005
R454 VSS.n1454 VSS.n1439 5.2005
R455 VSS.n1453 VSS.n1440 5.2005
R456 VSS.n1451 VSS.n1448 5.2005
R457 VSS.n1349 VSS.n1348 5.2005
R458 VSS.n1327 VSS.n1325 5.2005
R459 VSS.n1312 VSS.n1300 5.2005
R460 VSS.n1313 VSS.n1299 5.2005
R461 VSS.n1315 VSS.n1296 5.2005
R462 VSS.n1316 VSS.n1295 5.2005
R463 VSS.n1318 VSS.n1172 5.2005
R464 VSS.n1166 VSS.n1164 5.2005
R465 VSS.n1494 VSS.n1493 5.2005
R466 VSS.n1494 VSS.n1492 5.2005
R467 VSS.n1166 VSS.n1163 5.2005
R468 VSS.n1501 VSS.n1500 5.2005
R469 VSS.n1504 VSS.n1503 5.2005
R470 VSS.n1506 VSS.n1505 5.2005
R471 VSS.n1508 VSS.n1507 5.2005
R472 VSS.n1510 VSS.n1509 5.2005
R473 VSS.n29 VSS.n28 5.2005
R474 VSS.n32 VSS.n31 5.2005
R475 VSS.n35 VSS.n34 5.2005
R476 VSS.n37 VSS.n36 5.2005
R477 VSS.n39 VSS.n38 5.2005
R478 VSS.n42 VSS.n41 5.2005
R479 VSS.n47 VSS.n46 5.2005
R480 VSS.n49 VSS.n48 5.2005
R481 VSS.n52 VSS.n51 5.2005
R482 VSS.n54 VSS.n53 5.2005
R483 VSS.n57 VSS.n56 5.2005
R484 VSS.n59 VSS.n58 5.2005
R485 VSS.n62 VSS.n61 5.2005
R486 VSS.n64 VSS.n63 5.2005
R487 VSS.n67 VSS.n66 5.2005
R488 VSS.n69 VSS.n68 5.2005
R489 VSS.n74 VSS.n73 5.2005
R490 VSS.n77 VSS.n76 5.2005
R491 VSS.n81 VSS.n80 5.2005
R492 VSS.n83 VSS.n82 5.2005
R493 VSS.n86 VSS.n85 5.2005
R494 VSS.n88 VSS.n87 5.2005
R495 VSS.n91 VSS.n90 5.2005
R496 VSS.n94 VSS.n93 5.2005
R497 VSS.n1934 VSS.n1933 5.2005
R498 VSS.n1936 VSS.n1935 5.2005
R499 VSS.n1938 VSS.n1937 5.2005
R500 VSS.n1940 VSS.n1939 5.2005
R501 VSS.n1944 VSS.n1943 5.2005
R502 VSS.n1948 VSS.n1947 5.2005
R503 VSS.n1950 VSS.n1949 5.2005
R504 VSS.n1953 VSS.n1952 5.2005
R505 VSS.n1956 VSS.n1955 5.2005
R506 VSS.n1958 VSS.n1957 5.2005
R507 VSS.n1960 VSS.n1959 5.2005
R508 VSS.n1962 VSS.n1961 5.2005
R509 VSS.n1965 VSS.n1964 5.2005
R510 VSS.n1967 VSS.n1966 5.2005
R511 VSS.n1969 VSS.n1968 5.2005
R512 VSS.n1971 VSS.n1970 5.2005
R513 VSS.n1975 VSS.n1974 5.2005
R514 VSS.n1977 VSS.n1976 5.2005
R515 VSS.n1979 VSS.n1978 5.2005
R516 VSS.n1982 VSS.n1981 5.2005
R517 VSS.n1986 VSS.n1985 5.2005
R518 VSS.n1988 VSS.n1987 5.2005
R519 VSS.n1990 VSS.n1989 5.2005
R520 VSS.n1992 VSS.n1991 5.2005
R521 VSS.n404 VSS.n399 5.2005
R522 VSS.n405 VSS.n398 5.2005
R523 VSS.n406 VSS.n397 5.2005
R524 VSS.n408 VSS.n393 5.2005
R525 VSS.n409 VSS.n392 5.2005
R526 VSS.n410 VSS.n391 5.2005
R527 VSS.n411 VSS.n390 5.2005
R528 VSS.n419 VSS.t11 5.2005
R529 VSS.n385 VSS.n384 5.2005
R530 VSS.n382 VSS.n381 5.2005
R531 VSS.n380 VSS.n379 5.2005
R532 VSS.n378 VSS.n377 5.2005
R533 VSS.n375 VSS.n374 5.2005
R534 VSS.n373 VSS.n372 5.2005
R535 VSS.n371 VSS.n370 5.2005
R536 VSS.n369 VSS.n368 5.2005
R537 VSS.n366 VSS.n365 5.2005
R538 VSS.n364 VSS.n363 5.2005
R539 VSS.n362 VSS.n361 5.2005
R540 VSS.n359 VSS.n358 5.2005
R541 VSS.n357 VSS.n356 5.2005
R542 VSS.n355 VSS.n354 5.2005
R543 VSS.n353 VSS.n352 5.2005
R544 VSS.n350 VSS.n349 5.2005
R545 VSS.n338 VSS.n337 5.2005
R546 VSS.n336 VSS.n335 5.2005
R547 VSS.n334 VSS.n333 5.2005
R548 VSS.n345 VSS.n343 5.2005
R549 VSS.n1684 VSS.n1683 5.2005
R550 VSS.n1682 VSS.n1681 5.2005
R551 VSS.n401 VSS.n400 5.2005
R552 VSS.n1686 VSS.n1679 5.2005
R553 VSS.n1687 VSS.n1678 5.2005
R554 VSS.n1688 VSS.n1677 5.2005
R555 VSS.n1689 VSS.n1676 5.2005
R556 VSS.n1690 VSS.n1675 5.2005
R557 VSS.n1691 VSS.n1673 5.2005
R558 VSS.n1692 VSS.n1672 5.2005
R559 VSS.n1693 VSS.n1671 5.2005
R560 VSS.n1694 VSS.n1670 5.2005
R561 VSS.n1695 VSS.n1669 5.2005
R562 VSS.n1696 VSS.n1668 5.2005
R563 VSS.n1697 VSS.n1667 5.2005
R564 VSS.n1699 VSS.n1698 5.2005
R565 VSS.n1666 VSS.n1665 5.2005
R566 VSS.n1664 VSS.n1663 5.2005
R567 VSS.n1661 VSS.n1660 5.2005
R568 VSS.n1659 VSS.n1658 5.2005
R569 VSS.n1657 VSS.n1656 5.2005
R570 VSS.n1654 VSS.n1653 5.2005
R571 VSS.n1652 VSS.n1651 5.2005
R572 VSS.n1650 VSS.n1649 5.2005
R573 VSS.n1648 VSS.n1647 5.2005
R574 VSS.n1634 VSS.n1633 5.2005
R575 VSS.n1632 VSS.n1631 5.2005
R576 VSS.n125 VSS.n124 5.2005
R577 VSS.n1917 VSS.n123 5.2005
R578 VSS.n1918 VSS.n122 5.2005
R579 VSS.n1919 VSS.n121 5.2005
R580 VSS.n1920 VSS.n120 5.2005
R581 VSS.n1921 VSS.n118 5.2005
R582 VSS.n1922 VSS.n117 5.2005
R583 VSS.n1923 VSS.n116 5.2005
R584 VSS.n1924 VSS.n113 5.2005
R585 VSS.n1925 VSS.n112 5.2005
R586 VSS.n1915 VSS 4.8968
R587 VSS.n1500 VSS.t308 4.79578
R588 VSS.n313 VSS.n312 4.62254
R589 VSS.n429 VSS.n426 4.62185
R590 VSS.n657 VSS.n656 4.53749
R591 VSS.t360 VSS.t153 4.53749
R592 VSS.n693 VSS.t357 4.53749
R593 VSS.n997 VSS.t84 4.53057
R594 VSS.n1887 VSS.t152 4.53057
R595 VSS.n1702 VSS.n1701 4.5005
R596 VSS.n1400 VSS.n1399 4.5005
R597 VSS.n1451 VSS.n1450 4.5005
R598 VSS.n1349 VSS.n1345 4.5005
R599 VSS.n1166 VSS.n1165 4.5005
R600 VSS.n345 VSS.n344 4.5005
R601 VSS.n314 VSS.n309 4.48602
R602 VSS.n646 VSS.t407 4.48602
R603 VSS.n430 VSS.n424 4.48602
R604 VSS.n441 VSS.t105 4.48602
R605 VSS.n1135 VSS.t131 4.29565
R606 VSS.n1558 VSS.t185 4.29565
R607 VSS.n1974 VSS.n1973 4.0471
R608 VSS.n396 VSS.t244 4.0471
R609 VSS.n1096 VSS.t137 3.88342
R610 VSS.n1835 VSS.t361 3.88342
R611 VSS.n1624 VSS.n1623 3.78833
R612 VSS.n110 VSS.n109 3.78833
R613 VSS.n1700 VSS.n1597 3.78299
R614 VSS.t66 VSS.n1009 3.78299
R615 VSS.n1489 VSS.n1389 3.77011
R616 VSS.n89 VSS.n3 3.7355
R617 VSS.n78 VSS.n7 3.7355
R618 VSS.n65 VSS.n11 3.7355
R619 VSS.n55 VSS.n15 3.7355
R620 VSS.n43 VSS.n19 3.7355
R621 VSS.n33 VSS.n23 3.7355
R622 VSS.n1490 VSS.n1321 3.72662
R623 VSS.n1609 VSS.n1608 3.71473
R624 VSS.n30 VSS.n25 3.7042
R625 VSS.n40 VSS.n21 3.7042
R626 VSS.n50 VSS.n17 3.7042
R627 VSS.n60 VSS.n13 3.7042
R628 VSS.n70 VSS.n9 3.7042
R629 VSS.n84 VSS.n5 3.7042
R630 VSS.n92 VSS.n1 3.7042
R631 VSS.n1941 VSS.n102 3.68267
R632 VSS.n1963 VSS.n99 3.68267
R633 VSS.n1983 VSS.n96 3.68267
R634 VSS.n1619 VSS.n1618 3.67443
R635 VSS.n650 VSS.n316 3.66702
R636 VSS.n437 VSS.n423 3.66702
R637 VSS.n1502 VSS.n1161 3.65528
R638 VSS.n1511 VSS.n1159 3.65528
R639 VSS.n1518 VSS.n1157 3.65528
R640 VSS.n1527 VSS.n1155 3.65528
R641 VSS.n1534 VSS.n1153 3.65528
R642 VSS.n1543 VSS.n1151 3.65528
R643 VSS.n1551 VSS.n1548 3.65528
R644 VSS.n1707 VSS.n1573 3.65528
R645 VSS.n1567 VSS.n1559 3.65208
R646 VSS.n407 VSS.n395 3.64941
R647 VSS.n412 VSS.n389 3.64941
R648 VSS.n416 VSS.n387 3.64941
R649 VSS.n383 VSS.n323 3.64941
R650 VSS.n376 VSS.n325 3.64941
R651 VSS.n367 VSS.n327 3.64941
R652 VSS.n360 VSS.n329 3.64941
R653 VSS.n351 VSS.n331 3.64941
R654 VSS.n1714 VSS.n1713 3.64802
R655 VSS.n1386 VSS.n1329 3.6318
R656 VSS.n1381 VSS.n1331 3.6318
R657 VSS.n1377 VSS.n1333 3.6318
R658 VSS.n1372 VSS.n1335 3.6318
R659 VSS.n1368 VSS.n1337 3.6318
R660 VSS.n1363 VSS.n1339 3.6318
R661 VSS.n1359 VSS.n1341 3.6318
R662 VSS.n1354 VSS.n1343 3.6318
R663 VSS.n1456 VSS.n1437 3.62593
R664 VSS.n1461 VSS.n1431 3.62593
R665 VSS.n1465 VSS.n1426 3.62593
R666 VSS.n1470 VSS.n1420 3.62593
R667 VSS.n1474 VSS.n1415 3.62593
R668 VSS.n1479 VSS.n1410 3.62593
R669 VSS.n1483 VSS.n1405 3.62593
R670 VSS.n1588 VSS.n1587 3.61811
R671 VSS.n1719 VSS.n1141 3.61811
R672 VSS.n1723 VSS.n1134 3.61811
R673 VSS.n1124 VSS.n1112 3.61811
R674 VSS.n1117 VSS.n1114 3.61811
R675 VSS.n1310 VSS.n1303 3.61811
R676 VSS.n1314 VSS.n1298 3.61811
R677 VSS.n337 VSS.t450 3.50643
R678 VSS.n368 VSS.t540 3.50643
R679 VSS.t481 VSS.t203 3.50643
R680 VSS.t307 VSS.n79 3.46902
R681 VSS.n1710 VSS.n1709 3.36271
R682 VSS.n1575 VSS.n1574 3.36271
R683 VSS.n1579 VSS.n1578 3.36271
R684 VSS.n1582 VSS.n1580 3.36271
R685 VSS.n1490 VSS.n1489 3.26287
R686 VSS.n1624 VSS.n1621 3.1505
R687 VSS.n1619 VSS.n1616 3.1505
R688 VSS.n110 VSS.n107 3.1505
R689 VSS.n1609 VSS.n1606 3.1505
R690 VSS.t295 VSS.t154 3.02516
R691 VSS.t321 VSS.t358 3.02516
R692 VSS.n395 VSS.t538 2.7305
R693 VSS.n395 VSS.n394 2.7305
R694 VSS.n389 VSS.t508 2.7305
R695 VSS.n389 VSS.n388 2.7305
R696 VSS.n387 VSS.t557 2.7305
R697 VSS.n387 VSS.n386 2.7305
R698 VSS.n323 VSS.t534 2.7305
R699 VSS.n323 VSS.n322 2.7305
R700 VSS.n325 VSS.t256 2.7305
R701 VSS.n325 VSS.n324 2.7305
R702 VSS.n327 VSS.t525 2.7305
R703 VSS.n327 VSS.n326 2.7305
R704 VSS.n329 VSS.t475 2.7305
R705 VSS.n329 VSS.n328 2.7305
R706 VSS.n331 VSS.t36 2.7305
R707 VSS.n331 VSS.n330 2.7305
R708 VSS.n1621 VSS.t444 2.7305
R709 VSS.n1621 VSS.n1620 2.7305
R710 VSS.n1623 VSS.t273 2.7305
R711 VSS.n1623 VSS.n1622 2.7305
R712 VSS.n1618 VSS.t110 2.7305
R713 VSS.n1618 VSS.n1617 2.7305
R714 VSS.n1616 VSS.t585 2.7305
R715 VSS.n1616 VSS.n1615 2.7305
R716 VSS.n107 VSS.t270 2.7305
R717 VSS.n107 VSS.n106 2.7305
R718 VSS.n109 VSS.t351 2.7305
R719 VSS.n109 VSS.n108 2.7305
R720 VSS.n1608 VSS.t271 2.7305
R721 VSS.n1608 VSS.n1607 2.7305
R722 VSS.n1606 VSS.t73 2.7305
R723 VSS.n1606 VSS.n1605 2.7305
R724 VSS.n1437 VSS.t235 2.7305
R725 VSS.n1437 VSS.n1436 2.7305
R726 VSS.n1431 VSS.t422 2.7305
R727 VSS.n1431 VSS.n1430 2.7305
R728 VSS.n1426 VSS.t230 2.7305
R729 VSS.n1426 VSS.n1425 2.7305
R730 VSS.n1420 VSS.t141 2.7305
R731 VSS.n1420 VSS.n1419 2.7305
R732 VSS.n1415 VSS.t224 2.7305
R733 VSS.n1415 VSS.n1414 2.7305
R734 VSS.n1410 VSS.t211 2.7305
R735 VSS.n1410 VSS.n1409 2.7305
R736 VSS.n1405 VSS.t144 2.7305
R737 VSS.n1405 VSS.n1404 2.7305
R738 VSS.n1329 VSS.t146 2.7305
R739 VSS.n1329 VSS.n1328 2.7305
R740 VSS.n1331 VSS.t237 2.7305
R741 VSS.n1331 VSS.n1330 2.7305
R742 VSS.n1333 VSS.t219 2.7305
R743 VSS.n1333 VSS.n1332 2.7305
R744 VSS.n1335 VSS.t212 2.7305
R745 VSS.n1335 VSS.n1334 2.7305
R746 VSS.n1337 VSS.t214 2.7305
R747 VSS.n1337 VSS.n1336 2.7305
R748 VSS.n1339 VSS.t427 2.7305
R749 VSS.n1339 VSS.n1338 2.7305
R750 VSS.n1341 VSS.t226 2.7305
R751 VSS.n1341 VSS.n1340 2.7305
R752 VSS.n1343 VSS.t291 2.7305
R753 VSS.n1343 VSS.n1342 2.7305
R754 VSS.n1161 VSS.t502 2.7305
R755 VSS.n1161 VSS.n1160 2.7305
R756 VSS.n1159 VSS.t484 2.7305
R757 VSS.n1159 VSS.n1158 2.7305
R758 VSS.n1157 VSS.t465 2.7305
R759 VSS.n1157 VSS.n1156 2.7305
R760 VSS.n1155 VSS.t527 2.7305
R761 VSS.n1155 VSS.n1154 2.7305
R762 VSS.n1153 VSS.t530 2.7305
R763 VSS.n1153 VSS.n1152 2.7305
R764 VSS.n1151 VSS.t512 2.7305
R765 VSS.n1151 VSS.n1150 2.7305
R766 VSS.n1548 VSS.t469 2.7305
R767 VSS.n1548 VSS.n1547 2.7305
R768 VSS.n1573 VSS.t486 2.7305
R769 VSS.n1573 VSS.n1572 2.7305
R770 VSS.n1587 VSS.t253 2.7305
R771 VSS.n1587 VSS.n1586 2.7305
R772 VSS.n1141 VSS.t255 2.7305
R773 VSS.n1141 VSS.n1140 2.7305
R774 VSS.n1134 VSS.t491 2.7305
R775 VSS.n1134 VSS.n1133 2.7305
R776 VSS.n1112 VSS.t519 2.7305
R777 VSS.n1112 VSS.n1111 2.7305
R778 VSS.n1114 VSS.t511 2.7305
R779 VSS.n1114 VSS.n1113 2.7305
R780 VSS.n1303 VSS.t467 2.7305
R781 VSS.n1303 VSS.n1302 2.7305
R782 VSS.n1298 VSS.t485 2.7305
R783 VSS.n1298 VSS.n1297 2.7305
R784 VSS.n25 VSS.t44 2.7305
R785 VSS.n25 VSS.n24 2.7305
R786 VSS.n21 VSS.t472 2.7305
R787 VSS.n21 VSS.n20 2.7305
R788 VSS.n17 VSS.t248 2.7305
R789 VSS.n17 VSS.n16 2.7305
R790 VSS.n13 VSS.t526 2.7305
R791 VSS.n13 VSS.n12 2.7305
R792 VSS.n9 VSS.t556 2.7305
R793 VSS.n9 VSS.n8 2.7305
R794 VSS.n5 VSS.t464 2.7305
R795 VSS.n5 VSS.n4 2.7305
R796 VSS.n1 VSS.t560 2.7305
R797 VSS.n1 VSS.n0 2.7305
R798 VSS.n3 VSS.t480 2.7305
R799 VSS.n3 VSS.n2 2.7305
R800 VSS.n7 VSS.t561 2.7305
R801 VSS.n7 VSS.n6 2.7305
R802 VSS.n11 VSS.t505 2.7305
R803 VSS.n11 VSS.n10 2.7305
R804 VSS.n15 VSS.t506 2.7305
R805 VSS.n15 VSS.n14 2.7305
R806 VSS.n19 VSS.t567 2.7305
R807 VSS.n19 VSS.n18 2.7305
R808 VSS.n23 VSS.t562 2.7305
R809 VSS.n23 VSS.n22 2.7305
R810 VSS.n102 VSS.t252 2.7305
R811 VSS.n102 VSS.n101 2.7305
R812 VSS.n99 VSS.t573 2.7305
R813 VSS.n99 VSS.n98 2.7305
R814 VSS.n96 VSS.t496 2.7305
R815 VSS.n96 VSS.n95 2.7305
R816 VSS.n927 VSS.n926 2.63579
R817 VSS.n1943 VSS.n1942 2.62995
R818 VSS.n886 VSS.n814 2.6255
R819 VSS.n885 VSS.n816 2.60377
R820 VSS.n1826 VSS.n250 2.60285
R821 VSS.n346 VSS.n341 2.60175
R822 VSS.n1583 VSS.n1582 2.60175
R823 VSS.n1497 VSS.n1496 2.60175
R824 VSS.n1171 VSS.n1170 2.60175
R825 VSS.n1442 VSS.n1441 2.60175
R826 VSS.n1394 VSS.n1393 2.60175
R827 VSS.n1351 VSS.n1344 2.60175
R828 VSS.n1324 VSS.n1323 2.60175
R829 VSS.n1444 VSS.n1442 2.601
R830 VSS.n1498 VSS.n1497 2.601
R831 VSS.n347 VSS.n346 2.601
R832 VSS.n1320 VSS.n1171 2.601
R833 VSS.n1395 VSS.n1394 2.601
R834 VSS.n546 VSS.n545 2.6005
R835 VSS.n545 VSS.n544 2.6005
R836 VSS.n516 VSS.n515 2.6005
R837 VSS.n515 VSS.n514 2.6005
R838 VSS.n519 VSS.n518 2.6005
R839 VSS.n518 VSS.n517 2.6005
R840 VSS.n522 VSS.n521 2.6005
R841 VSS.n521 VSS.n520 2.6005
R842 VSS.n525 VSS.n524 2.6005
R843 VSS.n524 VSS.n523 2.6005
R844 VSS.n528 VSS.n527 2.6005
R845 VSS.n527 VSS.n526 2.6005
R846 VSS.n531 VSS.n530 2.6005
R847 VSS.n530 VSS.n529 2.6005
R848 VSS.n534 VSS.n533 2.6005
R849 VSS.n533 VSS.n532 2.6005
R850 VSS.n537 VSS.n536 2.6005
R851 VSS.n536 VSS.n535 2.6005
R852 VSS.n540 VSS.n539 2.6005
R853 VSS.n539 VSS.n538 2.6005
R854 VSS.n543 VSS.n542 2.6005
R855 VSS.n542 VSS.n541 2.6005
R856 VSS.n513 VSS.n512 2.6005
R857 VSS.n512 VSS.n511 2.6005
R858 VSS.n510 VSS.n509 2.6005
R859 VSS.n509 VSS.n508 2.6005
R860 VSS.n495 VSS.n494 2.6005
R861 VSS.n494 VSS.n493 2.6005
R862 VSS.n498 VSS.n497 2.6005
R863 VSS.n497 VSS.n496 2.6005
R864 VSS.n501 VSS.n500 2.6005
R865 VSS.n500 VSS.n499 2.6005
R866 VSS.n504 VSS.n503 2.6005
R867 VSS.n503 VSS.n502 2.6005
R868 VSS.n507 VSS.n506 2.6005
R869 VSS.n506 VSS.n505 2.6005
R870 VSS.n492 VSS.n491 2.6005
R871 VSS.n491 VSS.n490 2.6005
R872 VSS.n489 VSS.n488 2.6005
R873 VSS.n488 VSS.n487 2.6005
R874 VSS.n474 VSS.n473 2.6005
R875 VSS.n473 VSS.n472 2.6005
R876 VSS.n477 VSS.n476 2.6005
R877 VSS.n476 VSS.n475 2.6005
R878 VSS.n480 VSS.n479 2.6005
R879 VSS.n479 VSS.n478 2.6005
R880 VSS.n483 VSS.n482 2.6005
R881 VSS.n482 VSS.n481 2.6005
R882 VSS.n486 VSS.n485 2.6005
R883 VSS.n485 VSS.n484 2.6005
R884 VSS.n471 VSS.n470 2.6005
R885 VSS.n470 VSS.n469 2.6005
R886 VSS.n468 VSS.n467 2.6005
R887 VSS.n467 VSS.n466 2.6005
R888 VSS.n453 VSS.n452 2.6005
R889 VSS.n452 VSS.n451 2.6005
R890 VSS.n456 VSS.n455 2.6005
R891 VSS.n455 VSS.n454 2.6005
R892 VSS.n459 VSS.n458 2.6005
R893 VSS.n458 VSS.n457 2.6005
R894 VSS.n462 VSS.n461 2.6005
R895 VSS.n461 VSS.n460 2.6005
R896 VSS.n465 VSS.n464 2.6005
R897 VSS.n464 VSS.n463 2.6005
R898 VSS.n450 VSS.n449 2.6005
R899 VSS.n449 VSS.n448 2.6005
R900 VSS.n447 VSS.n446 2.6005
R901 VSS.n446 VSS.n445 2.6005
R902 VSS.n428 VSS.n427 2.6005
R903 VSS.n433 VSS.n431 2.6005
R904 VSS.n433 VSS.n432 2.6005
R905 VSS.n436 VSS.n435 2.6005
R906 VSS.n435 VSS.n434 2.6005
R907 VSS.n440 VSS.n439 2.6005
R908 VSS.n439 VSS.n438 2.6005
R909 VSS.n444 VSS.n443 2.6005
R910 VSS.n443 VSS.n442 2.6005
R911 VSS.n549 VSS.n548 2.6005
R912 VSS.n548 VSS.n547 2.6005
R913 VSS.n550 VSS.n421 2.6005
R914 VSS.n1750 VSS.n1102 2.6005
R915 VSS.n1221 VSS.n1220 2.6005
R916 VSS.n1224 VSS.n1223 2.6005
R917 VSS.n1223 VSS.n1222 2.6005
R918 VSS.n1227 VSS.n1226 2.6005
R919 VSS.n1226 VSS.n1225 2.6005
R920 VSS.n1230 VSS.n1229 2.6005
R921 VSS.n1229 VSS.n1228 2.6005
R922 VSS.n1233 VSS.n1232 2.6005
R923 VSS.n1232 VSS.n1231 2.6005
R924 VSS.n1236 VSS.n1235 2.6005
R925 VSS.n1235 VSS.n1234 2.6005
R926 VSS.n1239 VSS.n1238 2.6005
R927 VSS.n1238 VSS.n1237 2.6005
R928 VSS.n1243 VSS.n1242 2.6005
R929 VSS.n1242 VSS.n1241 2.6005
R930 VSS.n1246 VSS.n1245 2.6005
R931 VSS.n1245 VSS.n1244 2.6005
R932 VSS.n1249 VSS.n1248 2.6005
R933 VSS.n1248 VSS.n1247 2.6005
R934 VSS.n1252 VSS.n1251 2.6005
R935 VSS.n1251 VSS.n1250 2.6005
R936 VSS.n1255 VSS.n1254 2.6005
R937 VSS.n1254 VSS.n1253 2.6005
R938 VSS.n1258 VSS.n1257 2.6005
R939 VSS.n1257 VSS.n1256 2.6005
R940 VSS.n1261 VSS.n1260 2.6005
R941 VSS.n1260 VSS.n1259 2.6005
R942 VSS.n1264 VSS.n1263 2.6005
R943 VSS.n1263 VSS.n1262 2.6005
R944 VSS.n1267 VSS.n1266 2.6005
R945 VSS.n1266 VSS.n1265 2.6005
R946 VSS.n1270 VSS.n1269 2.6005
R947 VSS.n1269 VSS.n1268 2.6005
R948 VSS.n1273 VSS.n1272 2.6005
R949 VSS.n1272 VSS.n1271 2.6005
R950 VSS.n1276 VSS.n1275 2.6005
R951 VSS.n1275 VSS.n1274 2.6005
R952 VSS.n1279 VSS.n1278 2.6005
R953 VSS.n1278 VSS.n1277 2.6005
R954 VSS.n1282 VSS.n1281 2.6005
R955 VSS.n1281 VSS.n1280 2.6005
R956 VSS.n1285 VSS.n1284 2.6005
R957 VSS.n1284 VSS.n1283 2.6005
R958 VSS.n1738 VSS.n1737 2.6005
R959 VSS.n1740 VSS.n1739 2.6005
R960 VSS.n1743 VSS.n1742 2.6005
R961 VSS.n1746 VSS.n1745 2.6005
R962 VSS.n1749 VSS.n1748 2.6005
R963 VSS.n1291 VSS.n1290 2.6005
R964 VSS.n1293 VSS.n1292 2.6005
R965 VSS.n1192 VSS.n1191 2.6005
R966 VSS.n1195 VSS.n1194 2.6005
R967 VSS.n1197 VSS.n1196 2.6005
R968 VSS.n1200 VSS.n1199 2.6005
R969 VSS.n1202 VSS.n1201 2.6005
R970 VSS.n1205 VSS.n1204 2.6005
R971 VSS.n1207 VSS.n1206 2.6005
R972 VSS.n1210 VSS.n1209 2.6005
R973 VSS.n1212 VSS.n1211 2.6005
R974 VSS.n1216 VSS.n1215 2.6005
R975 VSS.n1288 VSS.n1287 2.6005
R976 VSS.n1287 VSS.n1286 2.6005
R977 VSS.n1104 VSS.n1103 2.6005
R978 VSS.n1219 VSS.n1218 2.6005
R979 VSS.n1218 VSS.n1217 2.6005
R980 VSS.n1901 VSS.n1900 2.6005
R981 VSS.n1900 VSS.n1899 2.6005
R982 VSS.n250 VSS.n249 2.6005
R983 VSS.n133 VSS.n132 2.6005
R984 VSS.n135 VSS.n134 2.6005
R985 VSS.n137 VSS.n136 2.6005
R986 VSS.n139 VSS.n138 2.6005
R987 VSS.n141 VSS.n140 2.6005
R988 VSS.n143 VSS.n142 2.6005
R989 VSS.n254 VSS.n253 2.6005
R990 VSS.n230 VSS.n229 2.6005
R991 VSS.n228 VSS.n227 2.6005
R992 VSS.n226 VSS.n225 2.6005
R993 VSS.n221 VSS.n220 2.6005
R994 VSS.n219 VSS.n218 2.6005
R995 VSS.n217 VSS.n216 2.6005
R996 VSS.n216 VSS.n215 2.6005
R997 VSS.n214 VSS.n213 2.6005
R998 VSS.n211 VSS.n210 2.6005
R999 VSS.n209 VSS.n208 2.6005
R1000 VSS.n207 VSS.n206 2.6005
R1001 VSS.n204 VSS.n203 2.6005
R1002 VSS.n202 VSS.n201 2.6005
R1003 VSS.n201 VSS.n200 2.6005
R1004 VSS.n199 VSS.n198 2.6005
R1005 VSS.n195 VSS.n194 2.6005
R1006 VSS.n193 VSS.n192 2.6005
R1007 VSS.n192 VSS.n191 2.6005
R1008 VSS.n190 VSS.n189 2.6005
R1009 VSS.n187 VSS.n186 2.6005
R1010 VSS.n185 VSS.n184 2.6005
R1011 VSS.n183 VSS.n182 2.6005
R1012 VSS.n180 VSS.n179 2.6005
R1013 VSS.n178 VSS.n177 2.6005
R1014 VSS.n176 VSS.n175 2.6005
R1015 VSS.n174 VSS.n173 2.6005
R1016 VSS.n171 VSS.n170 2.6005
R1017 VSS.n233 VSS.n232 2.6005
R1018 VSS.n232 VSS.n231 2.6005
R1019 VSS.n1830 VSS.n1829 2.6005
R1020 VSS.n1829 VSS.n1828 2.6005
R1021 VSS.n247 VSS.n246 2.6005
R1022 VSS.n246 VSS.n245 2.6005
R1023 VSS.n238 VSS.n237 2.6005
R1024 VSS.n237 VSS.n236 2.6005
R1025 VSS.n243 VSS.n242 2.6005
R1026 VSS.n242 VSS.n241 2.6005
R1027 VSS.n1905 VSS.n1904 2.6005
R1028 VSS.n1904 VSS.n1903 2.6005
R1029 VSS.n1909 VSS.n1908 2.6005
R1030 VSS.n1908 VSS.n1907 2.6005
R1031 VSS.n1838 VSS.n1837 2.6005
R1032 VSS.n1837 VSS.n1836 2.6005
R1033 VSS.n1842 VSS.n1841 2.6005
R1034 VSS.n1841 VSS.n1840 2.6005
R1035 VSS.n1846 VSS.n1845 2.6005
R1036 VSS.n1845 VSS.n1844 2.6005
R1037 VSS.n1850 VSS.n1849 2.6005
R1038 VSS.n1849 VSS.n1848 2.6005
R1039 VSS.n1881 VSS.n1880 2.6005
R1040 VSS.n1880 VSS.n1879 2.6005
R1041 VSS.n1834 VSS.n1833 2.6005
R1042 VSS.n1833 VSS.n1832 2.6005
R1043 VSS.n1854 VSS.n1853 2.6005
R1044 VSS.n1853 VSS.n1852 2.6005
R1045 VSS.n1858 VSS.n1857 2.6005
R1046 VSS.n1857 VSS.n1856 2.6005
R1047 VSS.n1862 VSS.n1861 2.6005
R1048 VSS.n1861 VSS.n1860 2.6005
R1049 VSS.n1865 VSS.n1864 2.6005
R1050 VSS.n1864 VSS.n1863 2.6005
R1051 VSS.n1869 VSS.n1868 2.6005
R1052 VSS.n1868 VSS.n1867 2.6005
R1053 VSS.n1873 VSS.n1872 2.6005
R1054 VSS.n1872 VSS.n1871 2.6005
R1055 VSS.n1877 VSS.n1876 2.6005
R1056 VSS.n1876 VSS.n1875 2.6005
R1057 VSS.n1885 VSS.n1884 2.6005
R1058 VSS.n1884 VSS.n1883 2.6005
R1059 VSS.n1889 VSS.n1888 2.6005
R1060 VSS.n1888 VSS.n1887 2.6005
R1061 VSS.n1893 VSS.n1892 2.6005
R1062 VSS.n1892 VSS.n1891 2.6005
R1063 VSS.n1897 VSS.n1896 2.6005
R1064 VSS.n1896 VSS.n1895 2.6005
R1065 VSS.n1825 VSS.n1824 2.6005
R1066 VSS.n1824 VSS.n1823 2.6005
R1067 VSS.n1822 VSS.n1821 2.6005
R1068 VSS.n1820 VSS.n1819 2.6005
R1069 VSS.n1818 VSS.n1817 2.6005
R1070 VSS.n1814 VSS.n1813 2.6005
R1071 VSS.n1812 VSS.n1811 2.6005
R1072 VSS.n1811 VSS.n1810 2.6005
R1073 VSS.n1809 VSS.n1808 2.6005
R1074 VSS.n1808 VSS.n1807 2.6005
R1075 VSS.n1806 VSS.n1805 2.6005
R1076 VSS.n1803 VSS.n1802 2.6005
R1077 VSS.n1801 VSS.n1800 2.6005
R1078 VSS.n1799 VSS.n1798 2.6005
R1079 VSS.n293 VSS.n292 2.6005
R1080 VSS.n291 VSS.n290 2.6005
R1081 VSS.n290 VSS.n289 2.6005
R1082 VSS.n288 VSS.n287 2.6005
R1083 VSS.n284 VSS.n283 2.6005
R1084 VSS.n282 VSS.n281 2.6005
R1085 VSS.n281 VSS.n280 2.6005
R1086 VSS.n279 VSS.n278 2.6005
R1087 VSS.n276 VSS.n275 2.6005
R1088 VSS.n274 VSS.n273 2.6005
R1089 VSS.n272 VSS.n271 2.6005
R1090 VSS.n269 VSS.n268 2.6005
R1091 VSS.n267 VSS.n266 2.6005
R1092 VSS.n265 VSS.n264 2.6005
R1093 VSS.n263 VSS.n262 2.6005
R1094 VSS.n260 VSS.n259 2.6005
R1095 VSS.n157 VSS.n156 2.6005
R1096 VSS.n165 VSS.n164 2.6005
R1097 VSS.n159 VSS.n158 2.6005
R1098 VSS.n155 VSS.n154 2.6005
R1099 VSS.n153 VSS.n152 2.6005
R1100 VSS.n151 VSS.n150 2.6005
R1101 VSS.n149 VSS.n148 2.6005
R1102 VSS.n147 VSS.n146 2.6005
R1103 VSS.n145 VSS.n144 2.6005
R1104 VSS.n258 VSS.n257 2.6005
R1105 VSS.n256 VSS.n255 2.6005
R1106 VSS.n252 VSS.n251 2.6005
R1107 VSS.n127 VSS.n126 2.6005
R1108 VSS.n129 VSS.n128 2.6005
R1109 VSS.n131 VSS.n130 2.6005
R1110 VSS.n161 VSS.n160 2.6005
R1111 VSS.n163 VSS.n162 2.6005
R1112 VSS.n167 VSS.n166 2.6005
R1113 VSS.n169 VSS.n168 2.6005
R1114 VSS.n1753 VSS.n1752 2.6005
R1115 VSS.n1755 VSS.n1754 2.6005
R1116 VSS.n1758 VSS.n1757 2.6005
R1117 VSS.n1761 VSS.n1760 2.6005
R1118 VSS.n1764 VSS.n1763 2.6005
R1119 VSS.n1767 VSS.n1766 2.6005
R1120 VSS.n1770 VSS.n1769 2.6005
R1121 VSS.n1773 VSS.n1772 2.6005
R1122 VSS.n1776 VSS.n1775 2.6005
R1123 VSS.n1779 VSS.n1778 2.6005
R1124 VSS.n1782 VSS.n1781 2.6005
R1125 VSS.n1785 VSS.n1784 2.6005
R1126 VSS.n1788 VSS.n1787 2.6005
R1127 VSS.n1791 VSS.n1790 2.6005
R1128 VSS.n1794 VSS.n1793 2.6005
R1129 VSS.n1091 VSS.n1090 2.6005
R1130 VSS.n1088 VSS.n1087 2.6005
R1131 VSS.n1085 VSS.n1084 2.6005
R1132 VSS.n1082 VSS.n1081 2.6005
R1133 VSS.n1079 VSS.n1078 2.6005
R1134 VSS.n1076 VSS.n1075 2.6005
R1135 VSS.n1073 VSS.n1072 2.6005
R1136 VSS.n1070 VSS.n1069 2.6005
R1137 VSS.n1067 VSS.n1066 2.6005
R1138 VSS.n1064 VSS.n1063 2.6005
R1139 VSS.n1061 VSS.n1060 2.6005
R1140 VSS.n1058 VSS.n1057 2.6005
R1141 VSS.n1055 VSS.n1054 2.6005
R1142 VSS.n1052 VSS.n1051 2.6005
R1143 VSS.n1050 VSS.n1049 2.6005
R1144 VSS.n1048 VSS.n1047 2.6005
R1145 VSS.n1046 VSS.n1045 2.6005
R1146 VSS.n811 VSS.n810 2.6005
R1147 VSS.n810 VSS.n809 2.6005
R1148 VSS.n808 VSS.n807 2.6005
R1149 VSS.n807 VSS.n806 2.6005
R1150 VSS.n805 VSS.n804 2.6005
R1151 VSS.n804 VSS.n803 2.6005
R1152 VSS.n801 VSS.n800 2.6005
R1153 VSS.n800 VSS.n799 2.6005
R1154 VSS.n798 VSS.n797 2.6005
R1155 VSS.n797 VSS.n796 2.6005
R1156 VSS.n795 VSS.n794 2.6005
R1157 VSS.n791 VSS.n790 2.6005
R1158 VSS.n788 VSS.n787 2.6005
R1159 VSS.n785 VSS.n784 2.6005
R1160 VSS.n782 VSS.n781 2.6005
R1161 VSS.n779 VSS.n778 2.6005
R1162 VSS.n776 VSS.n775 2.6005
R1163 VSS.n773 VSS.n772 2.6005
R1164 VSS.n771 VSS.n770 2.6005
R1165 VSS.n945 VSS.n944 2.6005
R1166 VSS.n947 VSS.n946 2.6005
R1167 VSS.n950 VSS.n949 2.6005
R1168 VSS.n952 VSS.n951 2.6005
R1169 VSS.n955 VSS.n954 2.6005
R1170 VSS.n957 VSS.n956 2.6005
R1171 VSS.n960 VSS.n959 2.6005
R1172 VSS.n962 VSS.n961 2.6005
R1173 VSS.n966 VSS.n965 2.6005
R1174 VSS.n1042 VSS.n1041 2.6005
R1175 VSS.n1041 VSS.n1040 2.6005
R1176 VSS.n1037 VSS.n1036 2.6005
R1177 VSS.n1036 VSS.n1035 2.6005
R1178 VSS.n1034 VSS.n1033 2.6005
R1179 VSS.n1033 VSS.n1032 2.6005
R1180 VSS.n1031 VSS.n1030 2.6005
R1181 VSS.n1030 VSS.n1029 2.6005
R1182 VSS.n1028 VSS.n1027 2.6005
R1183 VSS.n1027 VSS.n1026 2.6005
R1184 VSS.n1025 VSS.n1024 2.6005
R1185 VSS.n1024 VSS.n1023 2.6005
R1186 VSS.n1022 VSS.n1021 2.6005
R1187 VSS.n1021 VSS.n1020 2.6005
R1188 VSS.n1019 VSS.n1018 2.6005
R1189 VSS.n1018 VSS.n1017 2.6005
R1190 VSS.n1016 VSS.n1015 2.6005
R1191 VSS.n1015 VSS.n1014 2.6005
R1192 VSS.n1012 VSS.n1011 2.6005
R1193 VSS.n1011 VSS.n1010 2.6005
R1194 VSS.n1008 VSS.n1007 2.6005
R1195 VSS.n1007 VSS.n1006 2.6005
R1196 VSS.n1005 VSS.n1004 2.6005
R1197 VSS.n1004 VSS.n1003 2.6005
R1198 VSS.n1002 VSS.n1001 2.6005
R1199 VSS.n1001 VSS.n1000 2.6005
R1200 VSS.n999 VSS.n998 2.6005
R1201 VSS.n998 VSS.n997 2.6005
R1202 VSS.n996 VSS.n995 2.6005
R1203 VSS.n995 VSS.n994 2.6005
R1204 VSS.n993 VSS.n992 2.6005
R1205 VSS.n992 VSS.n991 2.6005
R1206 VSS.n990 VSS.n989 2.6005
R1207 VSS.n989 VSS.n988 2.6005
R1208 VSS.n987 VSS.n986 2.6005
R1209 VSS.n986 VSS.n985 2.6005
R1210 VSS.n984 VSS.n983 2.6005
R1211 VSS.n983 VSS.n982 2.6005
R1212 VSS.n981 VSS.n980 2.6005
R1213 VSS.n980 VSS.n979 2.6005
R1214 VSS.n978 VSS.n977 2.6005
R1215 VSS.n977 VSS.n976 2.6005
R1216 VSS.n975 VSS.n974 2.6005
R1217 VSS.n974 VSS.n973 2.6005
R1218 VSS.n972 VSS.n971 2.6005
R1219 VSS.n971 VSS.t167 2.6005
R1220 VSS.n970 VSS.n969 2.6005
R1221 VSS.n969 VSS.n968 2.6005
R1222 VSS.n814 VSS.n813 2.6005
R1223 VSS.n884 VSS.n883 2.6005
R1224 VSS.n882 VSS.n881 2.6005
R1225 VSS.n868 VSS.n867 2.6005
R1226 VSS.n866 VSS.n865 2.6005
R1227 VSS.n863 VSS.n862 2.6005
R1228 VSS.n860 VSS.n859 2.6005
R1229 VSS.n858 VSS.n857 2.6005
R1230 VSS.n855 VSS.n854 2.6005
R1231 VSS.n853 VSS.n852 2.6005
R1232 VSS.n850 VSS.n849 2.6005
R1233 VSS.n848 VSS.n847 2.6005
R1234 VSS.n845 VSS.n844 2.6005
R1235 VSS.n843 VSS.n842 2.6005
R1236 VSS.n840 VSS.n839 2.6005
R1237 VSS.n838 VSS.n837 2.6005
R1238 VSS.n836 VSS.n835 2.6005
R1239 VSS.n834 VSS.n833 2.6005
R1240 VSS.n832 VSS.n831 2.6005
R1241 VSS.n830 VSS.n829 2.6005
R1242 VSS.n828 VSS.n827 2.6005
R1243 VSS.n826 VSS.n825 2.6005
R1244 VSS.n824 VSS.n823 2.6005
R1245 VSS.n822 VSS.n821 2.6005
R1246 VSS.n820 VSS.n819 2.6005
R1247 VSS.n818 VSS.n817 2.6005
R1248 VSS.n1174 VSS.n1173 2.6005
R1249 VSS.n1176 VSS.n1175 2.6005
R1250 VSS.n1178 VSS.n1177 2.6005
R1251 VSS.n1180 VSS.n1179 2.6005
R1252 VSS.n1182 VSS.n1181 2.6005
R1253 VSS.n1184 VSS.n1183 2.6005
R1254 VSS.n1186 VSS.n1185 2.6005
R1255 VSS.n1188 VSS.n1187 2.6005
R1256 VSS.n1190 VSS.n1189 2.6005
R1257 VSS.n1093 VSS.n1092 2.6005
R1258 VSS.n1099 VSS.n1098 2.6005
R1259 VSS.n311 VSS.n310 2.6005
R1260 VSS.n655 VSS.n654 2.6005
R1261 VSS.n656 VSS.n655 2.6005
R1262 VSS.n653 VSS.n652 2.6005
R1263 VSS.n652 VSS.n651 2.6005
R1264 VSS.n649 VSS.n648 2.6005
R1265 VSS.n648 VSS.n647 2.6005
R1266 VSS.n645 VSS.n644 2.6005
R1267 VSS.n644 VSS.n643 2.6005
R1268 VSS.n642 VSS.n641 2.6005
R1269 VSS.n641 VSS.n640 2.6005
R1270 VSS.n612 VSS.n320 2.6005
R1271 VSS.n320 VSS.n319 2.6005
R1272 VSS.n617 VSS.n616 2.6005
R1273 VSS.n616 VSS.n615 2.6005
R1274 VSS.n614 VSS.n613 2.6005
R1275 VSS.n620 VSS.n619 2.6005
R1276 VSS.n619 VSS.n618 2.6005
R1277 VSS.n621 VSS.n318 2.6005
R1278 VSS.n318 VSS.n317 2.6005
R1279 VSS.n636 VSS.n635 2.6005
R1280 VSS.n635 VSS.n634 2.6005
R1281 VSS.n633 VSS.n632 2.6005
R1282 VSS.n632 VSS.n631 2.6005
R1283 VSS.n630 VSS.n629 2.6005
R1284 VSS.n629 VSS.n628 2.6005
R1285 VSS.n627 VSS.n626 2.6005
R1286 VSS.n626 VSS.n625 2.6005
R1287 VSS.n624 VSS.n623 2.6005
R1288 VSS.n623 VSS.n622 2.6005
R1289 VSS.n639 VSS.n638 2.6005
R1290 VSS.n638 VSS.n637 2.6005
R1291 VSS.n768 VSS.n767 2.6005
R1292 VSS.n762 VSS.n761 2.6005
R1293 VSS.n759 VSS.n758 2.6005
R1294 VSS.n756 VSS.n755 2.6005
R1295 VSS.n753 VSS.n752 2.6005
R1296 VSS.n750 VSS.n749 2.6005
R1297 VSS.n747 VSS.n746 2.6005
R1298 VSS.n744 VSS.n743 2.6005
R1299 VSS.n741 VSS.n740 2.6005
R1300 VSS.n738 VSS.n737 2.6005
R1301 VSS.n735 VSS.n734 2.6005
R1302 VSS.n732 VSS.n731 2.6005
R1303 VSS.n729 VSS.n728 2.6005
R1304 VSS.n726 VSS.n725 2.6005
R1305 VSS.n723 VSS.n722 2.6005
R1306 VSS.n720 VSS.n719 2.6005
R1307 VSS.n718 VSS.n717 2.6005
R1308 VSS.n716 VSS.n715 2.6005
R1309 VSS.n714 VSS.n713 2.6005
R1310 VSS.n893 VSS.n892 2.6005
R1311 VSS.n892 VSS.n891 2.6005
R1312 VSS.n890 VSS.n889 2.6005
R1313 VSS.n889 VSS.n888 2.6005
R1314 VSS.n296 VSS.n295 2.6005
R1315 VSS.n295 VSS.n294 2.6005
R1316 VSS.n299 VSS.n298 2.6005
R1317 VSS.n298 VSS.n297 2.6005
R1318 VSS.n302 VSS.n301 2.6005
R1319 VSS.n301 VSS.n300 2.6005
R1320 VSS.n305 VSS.n304 2.6005
R1321 VSS.n304 VSS.n303 2.6005
R1322 VSS.n308 VSS.n307 2.6005
R1323 VSS.n307 VSS.n306 2.6005
R1324 VSS.n659 VSS.n658 2.6005
R1325 VSS.n658 VSS.n657 2.6005
R1326 VSS.n662 VSS.n661 2.6005
R1327 VSS.n661 VSS.n660 2.6005
R1328 VSS.n665 VSS.n664 2.6005
R1329 VSS.n664 VSS.n663 2.6005
R1330 VSS.n668 VSS.n667 2.6005
R1331 VSS.n667 VSS.n666 2.6005
R1332 VSS.n671 VSS.n670 2.6005
R1333 VSS.n670 VSS.n669 2.6005
R1334 VSS.n674 VSS.n673 2.6005
R1335 VSS.n673 VSS.n672 2.6005
R1336 VSS.n677 VSS.n676 2.6005
R1337 VSS.n676 VSS.n675 2.6005
R1338 VSS.n680 VSS.n679 2.6005
R1339 VSS.n679 VSS.n678 2.6005
R1340 VSS.n683 VSS.n682 2.6005
R1341 VSS.n682 VSS.n681 2.6005
R1342 VSS.n686 VSS.n685 2.6005
R1343 VSS.n685 VSS.n684 2.6005
R1344 VSS.n689 VSS.n688 2.6005
R1345 VSS.n688 VSS.n687 2.6005
R1346 VSS.n692 VSS.n691 2.6005
R1347 VSS.n691 VSS.n690 2.6005
R1348 VSS.n695 VSS.n694 2.6005
R1349 VSS.n694 VSS.n693 2.6005
R1350 VSS.n698 VSS.n697 2.6005
R1351 VSS.n697 VSS.n696 2.6005
R1352 VSS.n701 VSS.n700 2.6005
R1353 VSS.n700 VSS.n699 2.6005
R1354 VSS.n704 VSS.n703 2.6005
R1355 VSS.n703 VSS.n702 2.6005
R1356 VSS.n707 VSS.n706 2.6005
R1357 VSS.n706 VSS.n705 2.6005
R1358 VSS.n711 VSS.n710 2.6005
R1359 VSS.n710 VSS.n709 2.6005
R1360 VSS.n895 VSS.n894 2.6005
R1361 VSS.n897 VSS.n896 2.6005
R1362 VSS.n899 VSS.n898 2.6005
R1363 VSS.n901 VSS.n900 2.6005
R1364 VSS.n903 VSS.n902 2.6005
R1365 VSS.n905 VSS.n904 2.6005
R1366 VSS.n907 VSS.n906 2.6005
R1367 VSS.n910 VSS.n909 2.6005
R1368 VSS.n912 VSS.n911 2.6005
R1369 VSS.n915 VSS.n914 2.6005
R1370 VSS.n917 VSS.n916 2.6005
R1371 VSS.n920 VSS.n919 2.6005
R1372 VSS.n922 VSS.n921 2.6005
R1373 VSS.n925 VSS.n924 2.6005
R1374 VSS.n928 VSS.n927 2.6005
R1375 VSS.n930 VSS.n929 2.6005
R1376 VSS.n933 VSS.n932 2.6005
R1377 VSS.n935 VSS.n934 2.6005
R1378 VSS.n942 VSS.n941 2.6005
R1379 VSS.n45 VSS.n44 2.6005
R1380 VSS.n581 VSS.n580 2.6005
R1381 VSS.n580 VSS.n579 2.6005
R1382 VSS.n578 VSS.n577 2.6005
R1383 VSS.n577 VSS.n576 2.6005
R1384 VSS.n575 VSS.n574 2.6005
R1385 VSS.n574 VSS.n573 2.6005
R1386 VSS.n572 VSS.n571 2.6005
R1387 VSS.n571 VSS.n570 2.6005
R1388 VSS.n569 VSS.n568 2.6005
R1389 VSS.n568 VSS.n567 2.6005
R1390 VSS.n566 VSS.n565 2.6005
R1391 VSS.n565 VSS.n564 2.6005
R1392 VSS.n563 VSS.n562 2.6005
R1393 VSS.n562 VSS.n561 2.6005
R1394 VSS.n560 VSS.n559 2.6005
R1395 VSS.n559 VSS.n558 2.6005
R1396 VSS.n557 VSS.n556 2.6005
R1397 VSS.n556 VSS.n555 2.6005
R1398 VSS.n553 VSS.n552 2.6005
R1399 VSS.n552 VSS.n551 2.6005
R1400 VSS.n1946 VSS.n1945 2.6005
R1401 VSS.n584 VSS.n321 2.6005
R1402 VSS.n599 VSS.n598 2.6005
R1403 VSS.n598 VSS.n597 2.6005
R1404 VSS.n596 VSS.n595 2.6005
R1405 VSS.n595 VSS.n594 2.6005
R1406 VSS.n593 VSS.n592 2.6005
R1407 VSS.n592 VSS.n591 2.6005
R1408 VSS.n590 VSS.n589 2.6005
R1409 VSS.n589 VSS.n588 2.6005
R1410 VSS.n587 VSS.n586 2.6005
R1411 VSS.n586 VSS.n585 2.6005
R1412 VSS.n602 VSS.n601 2.6005
R1413 VSS.n601 VSS.n600 2.6005
R1414 VSS.n611 VSS.n610 2.6005
R1415 VSS.n610 VSS.n609 2.6005
R1416 VSS.n608 VSS.n607 2.6005
R1417 VSS.n607 VSS.n606 2.6005
R1418 VSS.n605 VSS.n604 2.6005
R1419 VSS.n604 VSS.n603 2.6005
R1420 VSS.n1914 VSS.n1913 2.6005
R1421 VSS.n1913 VSS.n1912 2.6005
R1422 VSS.n806 VSS.t324 2.58911
R1423 VSS.n1703 VSS.n1576 2.55463
R1424 VSS.n1713 VSS.n1712 2.50665
R1425 VSS.n1566 VSS.n1559 2.50664
R1426 VSS.n1350 VSS.n1349 2.41907
R1427 VSS.n1495 VSS.n1494 2.41795
R1428 VSS.n1703 VSS.n1702 2.41733
R1429 VSS.n1596 VSS.n1595 2.41463
R1430 VSS.n1452 VSS.n1451 2.40822
R1431 VSS.n1168 VSS.n1166 2.40807
R1432 VSS.n1487 VSS.n1400 2.4075
R1433 VSS.n1388 VSS.n1327 2.40736
R1434 VSS.n1100 VSS.t296 2.39814
R1435 VSS.n722 VSS.n721 2.33733
R1436 VSS.n725 VSS.n724 2.33733
R1437 VSS.n728 VSS.n727 2.33733
R1438 VSS.n731 VSS.n730 2.33733
R1439 VSS.n734 VSS.n733 2.33733
R1440 VSS.n737 VSS.n736 2.33733
R1441 VSS.n740 VSS.n739 2.33733
R1442 VSS.n743 VSS.n742 2.33733
R1443 VSS.n746 VSS.n745 2.33733
R1444 VSS.n749 VSS.n748 2.33733
R1445 VSS.n752 VSS.n751 2.33733
R1446 VSS.n755 VSS.n754 2.33733
R1447 VSS.n758 VSS.n757 2.33733
R1448 VSS.n761 VSS.n760 2.33733
R1449 VSS.n775 VSS.n774 2.33733
R1450 VSS.n778 VSS.n777 2.33733
R1451 VSS.n781 VSS.n780 2.33733
R1452 VSS.n784 VSS.n783 2.33733
R1453 VSS.n787 VSS.n786 2.33733
R1454 VSS.n790 VSS.n789 2.33733
R1455 VSS.n1054 VSS.n1053 2.31748
R1456 VSS.n1057 VSS.n1056 2.31748
R1457 VSS.n1060 VSS.n1059 2.31748
R1458 VSS.n1063 VSS.n1062 2.31748
R1459 VSS.n1066 VSS.n1065 2.31748
R1460 VSS.n1069 VSS.n1068 2.31748
R1461 VSS.n1072 VSS.n1071 2.31748
R1462 VSS.n1075 VSS.n1074 2.31748
R1463 VSS.n1078 VSS.n1077 2.31748
R1464 VSS.n1081 VSS.n1080 2.31748
R1465 VSS.n1084 VSS.n1083 2.31748
R1466 VSS.n1087 VSS.n1086 2.31748
R1467 VSS.n1745 VSS.n1744 2.31748
R1468 VSS.n1742 VSS.n1741 2.31748
R1469 VSS.n1748 VSS.n1747 2.31748
R1470 VSS.n1793 VSS.n1792 2.31748
R1471 VSS.n1790 VSS.n1789 2.31748
R1472 VSS.n1787 VSS.n1786 2.31748
R1473 VSS.n1784 VSS.n1783 2.31748
R1474 VSS.n1781 VSS.n1780 2.31748
R1475 VSS.n1778 VSS.n1777 2.31748
R1476 VSS.n1775 VSS.n1774 2.31748
R1477 VSS.n1772 VSS.n1771 2.31748
R1478 VSS.n1769 VSS.n1768 2.31748
R1479 VSS.n1766 VSS.n1765 2.31748
R1480 VSS.n1763 VSS.n1762 2.31748
R1481 VSS.n1760 VSS.n1759 2.31748
R1482 VSS.n1757 VSS.n1756 2.31748
R1483 VSS.n392 VSS.t241 2.31284
R1484 VSS.n300 VSS.t58 2.269
R1485 VSS.n634 VSS.t447 2.269
R1486 VSS.n622 VSS.t381 2.269
R1487 VSS.n709 VSS.t200 2.269
R1488 VSS.n1495 VSS.n1490 2.26028
R1489 VSS.n1446 VSS.n1445 2.25438
R1490 VSS.n1489 VSS.n1488 2.25101
R1491 VSS.n1324 VSS.n1322 2.21822
R1492 VSS.n345 VSS.n342 2.15773
R1493 VSS.n1108 VSS.t461 2.13963
R1494 VSS.n71 VSS.t373 2.09053
R1495 VSS.n249 VSS.n248 1.94196
R1496 VSS.n1828 VSS.n1827 1.94196
R1497 VSS.n1832 VSS.n1831 1.94196
R1498 VSS.n1836 VSS.n1835 1.94196
R1499 VSS.n1840 VSS.n1839 1.94196
R1500 VSS.n1844 VSS.n1843 1.94196
R1501 VSS.n1848 VSS.n1847 1.94196
R1502 VSS.n1852 VSS.n1851 1.94196
R1503 VSS.n1856 VSS.n1855 1.94196
R1504 VSS.n1860 VSS.n1859 1.94196
R1505 VSS.n1867 VSS.n1866 1.94196
R1506 VSS.n1871 VSS.n1870 1.94196
R1507 VSS.n1875 VSS.n1874 1.94196
R1508 VSS.n1879 VSS.n1878 1.94196
R1509 VSS.n1883 VSS.n1882 1.94196
R1510 VSS.n1887 VSS.n1886 1.94196
R1511 VSS.n1891 VSS.n1890 1.94196
R1512 VSS.n1899 VSS.n1898 1.94196
R1513 VSS.n1903 VSS.n1902 1.94196
R1514 VSS.n1907 VSS.n1906 1.94196
R1515 VSS.n1906 VSS.t93 1.94196
R1516 VSS.n1912 VSS.n1911 1.94196
R1517 VSS.n245 VSS.n244 1.94196
R1518 VSS.n241 VSS.n240 1.94196
R1519 VSS.n236 VSS.n235 1.94196
R1520 VSS.n1349 VSS.n1346 1.9177
R1521 VSS.n313 VSS.n311 1.91746
R1522 VSS.n429 VSS.n428 1.91738
R1523 VSS.n1393 VSS.n1392 1.90778
R1524 VSS.n550 VSS.n549 1.90092
R1525 VSS.n1451 VSS.n1447 1.87311
R1526 VSS.n1400 VSS.n1396 1.82853
R1527 VSS.n1702 VSS.n1577 1.78394
R1528 VSS.n1933 VSS.t43 1.75347
R1529 VSS.n31 VSS.t312 1.75347
R1530 VSS.n1947 VSS.n1946 1.75347
R1531 VSS.n365 VSS.t197 1.75347
R1532 VSS.n46 VSS.n45 1.75347
R1533 VSS.n1494 VSS.n1491 1.73935
R1534 VSS.n1817 VSS.n1816 1.72162
R1535 VSS.n804 VSS.n802 1.7198
R1536 VSS.n909 VSS.n908 1.70459
R1537 VSS.n914 VSS.n913 1.70459
R1538 VSS.n919 VSS.n918 1.70459
R1539 VSS.n924 VSS.n923 1.70459
R1540 VSS.n932 VSS.n931 1.70459
R1541 VSS.n941 VSS.n940 1.70459
R1542 VSS.n954 VSS.n953 1.70459
R1543 VSS.n959 VSS.n958 1.70459
R1544 VSS.n965 VSS.n964 1.70459
R1545 VSS.n1582 VSS.n1581 1.68161
R1546 VSS.n225 VSS.n224 1.66913
R1547 VSS.n1805 VSS.n1804 1.61162
R1548 VSS.n1798 VSS.n1797 1.61162
R1549 VSS.n287 VSS.n286 1.61162
R1550 VSS.n278 VSS.n277 1.61162
R1551 VSS.n271 VSS.n270 1.61162
R1552 VSS.n262 VSS.n261 1.61162
R1553 VSS.n1166 VSS.n1162 1.6056
R1554 VSS.n1194 VSS.n1193 1.60368
R1555 VSS.n1199 VSS.n1198 1.60357
R1556 VSS.n1204 VSS.n1203 1.60357
R1557 VSS.n1209 VSS.n1208 1.60357
R1558 VSS.n1215 VSS.n1214 1.60357
R1559 VSS.n1290 VSS.n1289 1.60357
R1560 VSS.n862 VSS.n861 1.60357
R1561 VSS.n857 VSS.n856 1.60357
R1562 VSS.n852 VSS.n851 1.60357
R1563 VSS.n847 VSS.n846 1.60357
R1564 VSS.n842 VSS.n841 1.60357
R1565 VSS.n816 VSS.n815 1.58772
R1566 VSS.n1596 VSS.n1584 1.56101
R1567 VSS.n206 VSS.n205 1.55723
R1568 VSS.n189 VSS.n188 1.55723
R1569 VSS.n213 VSS.n212 1.55656
R1570 VSS.n198 VSS.n197 1.55656
R1571 VSS.n182 VSS.n181 1.55656
R1572 VSS.n173 VSS.n172 1.55656
R1573 VSS.t60 VSS.t61 1.51283
R1574 VSS.t92 VSS.t317 1.51283
R1575 VSS.n333 VSS.n332 1.51283
R1576 VSS.n1735 VSS.n1734 1.49543
R1577 VSS.n944 VSS.n943 1.45409
R1578 VSS.n949 VSS.n948 1.45409
R1579 VSS.n1096 VSS.n1094 1.44276
R1580 VSS.n1096 VSS.n1095 1.44276
R1581 VSS.n1994 VSS.n1993 1.43392
R1582 VSS.n765 VSS.n763 1.43284
R1583 VSS.n765 VSS.n764 1.43284
R1584 VSS.n1555 VSS.t45 1.43222
R1585 VSS.n1041 VSS.n1039 1.38322
R1586 VSS.n770 VSS.n769 1.35581
R1587 VSS.n713 VSS.n712 1.35581
R1588 VSS.n767 VSS.n766 1.35567
R1589 VSS.n794 VSS.n793 1.35567
R1590 VSS.n1045 VSS.n1044 1.34579
R1591 VSS.n1098 VSS.n1097 1.34579
R1592 VSS.n881 VSS.n880 1.34565
R1593 VSS.n865 VSS.n864 1.34565
R1594 VSS.n1090 VSS.n1089 1.34565
R1595 VSS.n1752 VSS.n1751 1.34565
R1596 VSS.n1102 VSS.n1101 1.34565
R1597 VSS.n1737 VSS.n1736 1.34565
R1598 VSS.n1932 VSS.n1931 1.34093
R1599 VSS.n118 VSS.t151 1.29481
R1600 VSS.n121 VSS.t91 1.29481
R1601 VSS.t119 VSS.n1894 1.29481
R1602 VSS.n1039 VSS.n1038 1.28007
R1603 VSS.n1927 VSS.n1926 1.22876
R1604 VSS.n1163 VSS.t29 1.19932
R1605 VSS.n76 VSS.n75 1.15667
R1606 VSS.n1976 VSS.t306 1.15667
R1607 VSS.n80 VSS.t307 1.15667
R1608 VSS.n1981 VSS.n1980 1.15667
R1609 VSS.n1713 VSS.n1559 1.11085
R1610 VSS.n1596 VSS.n1585 1.0212
R1611 VSS.n1625 VSS.n1624 0.96262
R1612 VSS.n1685 VSS.n1680 0.950708
R1613 VSS.t80 VSS.t13 0.876983
R1614 VSS.n1700 VSS.n1699 0.841053
R1615 VSS.n1097 VSS.n1096 0.838098
R1616 VSS.n1101 VSS.n1100 0.837901
R1617 VSS.n880 VSS.n879 0.837901
R1618 VSS.n793 VSS.n792 0.83122
R1619 VSS.n766 VSS.n765 0.83122
R1620 VSS.n316 VSS.t405 0.8195
R1621 VSS.n316 VSS.n315 0.8195
R1622 VSS.n423 VSS.t400 0.8195
R1623 VSS.n423 VSS.n422 0.8195
R1624 VSS.t171 VSS.t363 0.756666
R1625 VSS.t442 VSS.t592 0.756666
R1626 VSS.t596 VSS.t135 0.756666
R1627 VSS.t441 VSS.t161 0.756666
R1628 VSS.n663 VSS.t193 0.756666
R1629 VSS.t432 VSS.t591 0.756666
R1630 VSS.n1662 VSS.n1630 0.7259
R1631 VSS.n1149 VSS.n1148 0.702093
R1632 VSS.n1730 VSS.n1729 0.687093
R1633 VSS.n29 VSS.n27 0.661796
R1634 VSS.t133 VSS.t3 0.647653
R1635 VSS.n1006 VSS.t440 0.647653
R1636 VSS.n116 VSS.n114 0.647653
R1637 VSS.n1895 VSS.t119 0.647653
R1638 VSS.n223 VSS.n222 0.647653
R1639 VSS.n1702 VSS.n1583 0.645288
R1640 VSS.n404 VSS.n403 0.644436
R1641 VSS.n1796 VSS.n1795 0.619447
R1642 VSS.n403 VSS.n401 0.609948
R1643 VSS.n1630 VSS.n1628 0.5873
R1644 VSS.n334 VSS.n105 0.572793
R1645 VSS.n1731 VSS.n1107 0.546075
R1646 VSS.n1726 VSS.n1725 0.546075
R1647 VSS.n1716 VSS.n1715 0.546075
R1648 VSS.n197 VSS.n196 0.523222
R1649 VSS.n1603 VSS.n1602 0.506362
R1650 VSS.n1214 VSS.n1213 0.499715
R1651 VSS.n879 VSS.n878 0.499715
R1652 VSS.n879 VSS.n877 0.499715
R1653 VSS.n879 VSS.n876 0.499715
R1654 VSS.n879 VSS.n875 0.499715
R1655 VSS.n879 VSS.n874 0.499715
R1656 VSS.n879 VSS.n873 0.499715
R1657 VSS.n879 VSS.n872 0.499715
R1658 VSS.n879 VSS.n871 0.499715
R1659 VSS.n879 VSS.n870 0.499715
R1660 VSS.n879 VSS.n869 0.499715
R1661 VSS.n286 VSS.n285 0.49569
R1662 VSS.n111 VSS.n110 0.491587
R1663 VSS.n224 VSS.n223 0.466933
R1664 VSS.n1611 VSS.n1610 0.4638
R1665 VSS.n1626 VSS.n1625 0.46349
R1666 VSS.n1628 VSS.n1626 0.4559
R1667 VSS.n1637 VSS 0.451296
R1668 VSS VSS.n1561 0.451296
R1669 VSS.n1643 VSS 0.451296
R1670 VSS.n939 VSS.n938 0.449449
R1671 VSS.n964 VSS.n963 0.449206
R1672 VSS.n939 VSS.n937 0.449206
R1673 VSS.n939 VSS.n936 0.449206
R1674 VSS.n940 VSS.n939 0.449206
R1675 VSS.n1816 VSS.n1815 0.440691
R1676 VSS.n1610 VSS.n1609 0.438385
R1677 VSS.n105 VSS.n104 0.43314
R1678 VSS.n346 VSS.n345 0.426384
R1679 VSS.n710 VSS.n708 0.424742
R1680 VSS.n1931 VSS.n105 0.419588
R1681 VSS.n314 VSS.n313 0.418027
R1682 VSS.n430 VSS.n429 0.417783
R1683 VSS.n1611 VSS.n1604 0.4145
R1684 VSS.n1625 VSS.n1619 0.407107
R1685 VSS.n1927 VSS.n1925 0.406886
R1686 VSS.n1612 VSS.n1603 0.393086
R1687 VSS.n1686 VSS.n1685 0.381896
R1688 VSS.n1626 VSS.n1614 0.36591
R1689 VSS.n1219 VSS.n1216 0.358535
R1690 VSS.n1685 VSS.n1684 0.35163
R1691 VSS.n403 VSS.n402 0.312204
R1692 VSS.n1930 VSS.n1929 0.300993
R1693 VSS.n1928 VSS.n1927 0.296642
R1694 VSS.n1317 VSS.n1294 0.274667
R1695 VSS.n1715 VSS.n1557 0.274482
R1696 VSS.n1727 VSS.n1726 0.250589
R1697 VSS.n405 VSS.n404 0.242079
R1698 VSS.n1931 VSS.n1930 0.236806
R1699 VSS.n1602 VSS.n1601 0.230155
R1700 VSS.n1731 VSS 0.229881
R1701 VSS.n1612 VSS.n1611 0.225254
R1702 VSS.n1732 VSS.n1731 0.221916
R1703 VSS.n1726 VSS 0.201208
R1704 VSS.n554 VSS.n420 0.195703
R1705 VSS.n1915 VSS.n1914 0.183525
R1706 VSS VSS.n1994 0.183461
R1707 VSS.n1916 VSS.n1915 0.181256
R1708 VSS.n1715 VSS 0.177314
R1709 VSS.n621 VSS.n620 0.167855
R1710 VSS.n605 VSS.n602 0.167855
R1711 VSS.n584 VSS.n583 0.167855
R1712 VSS.n569 VSS.n566 0.167855
R1713 VSS.n471 VSS.n468 0.167855
R1714 VSS.n492 VSS.n489 0.167855
R1715 VSS.n513 VSS.n510 0.167855
R1716 VSS.n534 VSS.n531 0.167855
R1717 VSS.n1046 VSS.n1043 0.1605
R1718 VSS.n886 VSS.n885 0.159151
R1719 VSS.n1294 VSS.n1293 0.156333
R1720 VSS.n1734 VSS.n1733 0.152624
R1721 VSS.n1729 VSS.n1728 0.152624
R1722 VSS.n1556 VSS.n1149 0.152624
R1723 VSS.n642 VSS.n639 0.150091
R1724 VSS.n450 VSS.n447 0.150091
R1725 VSS.n639 VSS.n636 0.14926
R1726 VSS.n636 VSS.n633 0.14926
R1727 VSS.n633 VSS.n630 0.14926
R1728 VSS.n630 VSS.n627 0.14926
R1729 VSS.n627 VSS.n624 0.14926
R1730 VSS.n624 VSS.n621 0.14926
R1731 VSS.n620 VSS.n617 0.14926
R1732 VSS.n617 VSS.n614 0.14926
R1733 VSS.n614 VSS.n612 0.14926
R1734 VSS.n612 VSS.n611 0.14926
R1735 VSS.n611 VSS.n608 0.14926
R1736 VSS.n608 VSS.n605 0.14926
R1737 VSS.n602 VSS.n599 0.14926
R1738 VSS.n599 VSS.n596 0.14926
R1739 VSS.n596 VSS.n593 0.14926
R1740 VSS.n593 VSS.n590 0.14926
R1741 VSS.n590 VSS.n587 0.14926
R1742 VSS.n587 VSS.n584 0.14926
R1743 VSS.n583 VSS.n582 0.14926
R1744 VSS.n582 VSS.n581 0.14926
R1745 VSS.n581 VSS.n578 0.14926
R1746 VSS.n578 VSS.n575 0.14926
R1747 VSS.n575 VSS.n572 0.14926
R1748 VSS.n572 VSS.n569 0.14926
R1749 VSS.n566 VSS.n563 0.14926
R1750 VSS.n563 VSS.n560 0.14926
R1751 VSS.n453 VSS.n450 0.14926
R1752 VSS.n456 VSS.n453 0.14926
R1753 VSS.n459 VSS.n456 0.14926
R1754 VSS.n462 VSS.n459 0.14926
R1755 VSS.n465 VSS.n462 0.14926
R1756 VSS.n468 VSS.n465 0.14926
R1757 VSS.n474 VSS.n471 0.14926
R1758 VSS.n477 VSS.n474 0.14926
R1759 VSS.n480 VSS.n477 0.14926
R1760 VSS.n483 VSS.n480 0.14926
R1761 VSS.n486 VSS.n483 0.14926
R1762 VSS.n489 VSS.n486 0.14926
R1763 VSS.n495 VSS.n492 0.14926
R1764 VSS.n498 VSS.n495 0.14926
R1765 VSS.n501 VSS.n498 0.14926
R1766 VSS.n504 VSS.n501 0.14926
R1767 VSS.n507 VSS.n504 0.14926
R1768 VSS.n510 VSS.n507 0.14926
R1769 VSS.n516 VSS.n513 0.14926
R1770 VSS.n519 VSS.n516 0.14926
R1771 VSS.n522 VSS.n519 0.14926
R1772 VSS.n525 VSS.n522 0.14926
R1773 VSS.n528 VSS.n525 0.14926
R1774 VSS.n531 VSS.n528 0.14926
R1775 VSS.n537 VSS.n534 0.14926
R1776 VSS.n540 VSS.n537 0.14926
R1777 VSS.n543 VSS.n540 0.14926
R1778 VSS.n546 VSS.n543 0.14926
R1779 VSS VSS.n1637 0.139881
R1780 VSS VSS.n1561 0.139881
R1781 VSS VSS.n1732 0.139881
R1782 VSS VSS.n1727 0.139881
R1783 VSS.n1557 VSS 0.139881
R1784 VSS VSS.n1643 0.139881
R1785 VSS.n560 VSS.n557 0.138103
R1786 VSS.n1486 VSS.n1485 0.133192
R1787 VSS.n1485 VSS.n1484 0.133192
R1788 VSS.n1482 VSS.n1481 0.133192
R1789 VSS.n1481 VSS.n1480 0.133192
R1790 VSS.n1478 VSS.n1477 0.133192
R1791 VSS.n1477 VSS.n1476 0.133192
R1792 VSS.n1476 VSS.n1475 0.133192
R1793 VSS.n1473 VSS.n1472 0.133192
R1794 VSS.n1472 VSS.n1471 0.133192
R1795 VSS.n1469 VSS.n1468 0.133192
R1796 VSS.n1468 VSS.n1467 0.133192
R1797 VSS.n1467 VSS.n1466 0.133192
R1798 VSS.n1464 VSS.n1463 0.133192
R1799 VSS.n1463 VSS.n1462 0.133192
R1800 VSS.n1460 VSS.n1459 0.133192
R1801 VSS.n1459 VSS.n1458 0.133192
R1802 VSS.n1458 VSS.n1457 0.133192
R1803 VSS.n1455 VSS.n1454 0.133192
R1804 VSS.n1454 VSS.n1453 0.133192
R1805 VSS.n1385 VSS.n1384 0.133192
R1806 VSS.n1384 VSS.n1383 0.133192
R1807 VSS.n1383 VSS.n1382 0.133192
R1808 VSS.n1380 VSS.n1379 0.133192
R1809 VSS.n1379 VSS.n1378 0.133192
R1810 VSS.n1376 VSS.n1375 0.133192
R1811 VSS.n1375 VSS.n1374 0.133192
R1812 VSS.n1374 VSS.n1373 0.133192
R1813 VSS.n1371 VSS.n1370 0.133192
R1814 VSS.n1370 VSS.n1369 0.133192
R1815 VSS.n1367 VSS.n1366 0.133192
R1816 VSS.n1366 VSS.n1365 0.133192
R1817 VSS.n1365 VSS.n1364 0.133192
R1818 VSS.n1362 VSS.n1361 0.133192
R1819 VSS.n1361 VSS.n1360 0.133192
R1820 VSS.n1358 VSS.n1357 0.133192
R1821 VSS.n1357 VSS.n1356 0.133192
R1822 VSS.n1356 VSS.n1355 0.133192
R1823 VSS.n1506 VSS.n1504 0.133192
R1824 VSS.n1508 VSS.n1506 0.133192
R1825 VSS.n1510 VSS.n1508 0.133192
R1826 VSS.n1515 VSS.n1513 0.133192
R1827 VSS.n1517 VSS.n1515 0.133192
R1828 VSS.n1522 VSS.n1520 0.133192
R1829 VSS.n1524 VSS.n1522 0.133192
R1830 VSS.n1526 VSS.n1524 0.133192
R1831 VSS.n1531 VSS.n1529 0.133192
R1832 VSS.n1533 VSS.n1531 0.133192
R1833 VSS.n1538 VSS.n1536 0.133192
R1834 VSS.n1540 VSS.n1538 0.133192
R1835 VSS.n1542 VSS.n1540 0.133192
R1836 VSS.n1553 VSS.n1545 0.133192
R1837 VSS.n1553 VSS.n1552 0.133192
R1838 VSS.n1571 VSS.n1569 0.133192
R1839 VSS.n1708 VSS.n1571 0.133192
R1840 VSS.n1316 VSS.n1315 0.133192
R1841 VSS.n1313 VSS.n1312 0.133192
R1842 VSS.n1312 VSS.n1311 0.133192
R1843 VSS.n1309 VSS.n1308 0.133192
R1844 VSS.n1308 VSS.n1307 0.133192
R1845 VSS.n1121 VSS.n1119 0.133192
R1846 VSS.n1123 VSS.n1121 0.133192
R1847 VSS.n1129 VSS.n1126 0.133192
R1848 VSS.n1131 VSS.n1129 0.133192
R1849 VSS.n1722 VSS.n1721 0.133192
R1850 VSS.n1721 VSS.n1720 0.133192
R1851 VSS.n1720 VSS 0.133192
R1852 VSS.n1718 VSS.n1717 0.133192
R1853 VSS.n1590 VSS.n1589 0.133192
R1854 VSS.n1591 VSS.n1590 0.133192
R1855 VSS.n650 VSS.n649 0.13302
R1856 VSS.n440 VSS.n437 0.13302
R1857 VSS.n1381 VSS.n1380 0.132038
R1858 VSS.n1513 VSS.n1511 0.132038
R1859 VSS.n1719 VSS.n1718 0.132038
R1860 VSS.n1462 VSS.n1461 0.129731
R1861 VSS.n972 VSS.n970 0.127128
R1862 VSS.n975 VSS.n972 0.127128
R1863 VSS.n978 VSS.n975 0.127128
R1864 VSS.n981 VSS.n978 0.127128
R1865 VSS.n984 VSS.n981 0.127128
R1866 VSS.n987 VSS.n984 0.127128
R1867 VSS.n990 VSS.n987 0.127128
R1868 VSS.n993 VSS.n990 0.127128
R1869 VSS.n996 VSS.n993 0.127128
R1870 VSS.n999 VSS.n996 0.127128
R1871 VSS.n1002 VSS.n999 0.127128
R1872 VSS.n1005 VSS.n1002 0.127128
R1873 VSS.n1008 VSS.n1005 0.127128
R1874 VSS.n1012 VSS.n1008 0.127128
R1875 VSS.n1016 VSS.n1012 0.127128
R1876 VSS.n1019 VSS.n1016 0.127128
R1877 VSS.n1022 VSS.n1019 0.127128
R1878 VSS.n1025 VSS.n1022 0.127128
R1879 VSS.n1028 VSS.n1025 0.127128
R1880 VSS.n1031 VSS.n1028 0.127128
R1881 VSS.n1034 VSS.n1031 0.127128
R1882 VSS.n1037 VSS.n1034 0.127128
R1883 VSS.n1042 VSS.n1037 0.127128
R1884 VSS.n1221 VSS.n1219 0.127128
R1885 VSS.n1224 VSS.n1221 0.127128
R1886 VSS.n1227 VSS.n1224 0.127128
R1887 VSS.n1230 VSS.n1227 0.127128
R1888 VSS.n1233 VSS.n1230 0.127128
R1889 VSS.n1236 VSS.n1233 0.127128
R1890 VSS.n1239 VSS.n1236 0.127128
R1891 VSS.n1243 VSS.n1239 0.127128
R1892 VSS.n1246 VSS.n1243 0.127128
R1893 VSS.n1249 VSS.n1246 0.127128
R1894 VSS.n1252 VSS.n1249 0.127128
R1895 VSS.n1255 VSS.n1252 0.127128
R1896 VSS.n1258 VSS.n1255 0.127128
R1897 VSS.n1261 VSS.n1258 0.127128
R1898 VSS.n1264 VSS.n1261 0.127128
R1899 VSS.n1267 VSS.n1264 0.127128
R1900 VSS.n1270 VSS.n1267 0.127128
R1901 VSS.n1273 VSS.n1270 0.127128
R1902 VSS.n1276 VSS.n1273 0.127128
R1903 VSS.n1279 VSS.n1276 0.127128
R1904 VSS.n1282 VSS.n1279 0.127128
R1905 VSS.n1285 VSS.n1282 0.127128
R1906 VSS.n1288 VSS.n1285 0.127128
R1907 VSS.n1318 VSS.n1317 0.124538
R1908 VSS.n1388 VSS.n1387 0.121842
R1909 VSS.n1124 VSS.n1123 0.121654
R1910 VSS.n336 VSS.n334 0.121553
R1911 VSS.n338 VSS.n336 0.121553
R1912 VSS.n355 VSS.n353 0.121553
R1913 VSS.n357 VSS.n355 0.121553
R1914 VSS.n359 VSS.n357 0.121553
R1915 VSS.n364 VSS.n362 0.121553
R1916 VSS.n366 VSS.n364 0.121553
R1917 VSS.n371 VSS.n369 0.121553
R1918 VSS.n373 VSS.n371 0.121553
R1919 VSS.n375 VSS.n373 0.121553
R1920 VSS.n380 VSS.n378 0.121553
R1921 VSS.n382 VSS.n380 0.121553
R1922 VSS.n419 VSS.n418 0.121553
R1923 VSS.n418 VSS.n417 0.121553
R1924 VSS.n415 VSS.n414 0.121553
R1925 VSS.n414 VSS.n413 0.121553
R1926 VSS.n411 VSS.n410 0.121553
R1927 VSS.n410 VSS.n409 0.121553
R1928 VSS.n409 VSS.n408 0.121553
R1929 VSS.n406 VSS.n405 0.121553
R1930 VSS.n1684 VSS.n1682 0.121553
R1931 VSS.n1925 VSS.n1924 0.121553
R1932 VSS.n1924 VSS.n1923 0.121553
R1933 VSS.n1923 VSS.n1922 0.121553
R1934 VSS.n1922 VSS.n1921 0.121553
R1935 VSS.n1921 VSS.n1920 0.121553
R1936 VSS.n1920 VSS.n1919 0.121553
R1937 VSS.n1919 VSS.n1918 0.121553
R1938 VSS.n1918 VSS.n1917 0.121553
R1939 VSS.n1632 VSS.n125 0.121553
R1940 VSS.n1634 VSS.n1632 0.121553
R1941 VSS.n1648 VSS.n1634 0.121553
R1942 VSS.n1650 VSS.n1648 0.121553
R1943 VSS.n1652 VSS.n1650 0.121553
R1944 VSS.n1654 VSS.n1652 0.121553
R1945 VSS.n1657 VSS.n1654 0.121553
R1946 VSS.n1659 VSS.n1657 0.121553
R1947 VSS.n1661 VSS.n1659 0.121553
R1948 VSS.n1666 VSS.n1664 0.121553
R1949 VSS.n1698 VSS.n1666 0.121553
R1950 VSS.n1698 VSS.n1697 0.121553
R1951 VSS.n1697 VSS.n1696 0.121553
R1952 VSS.n1696 VSS.n1695 0.121553
R1953 VSS.n1695 VSS.n1694 0.121553
R1954 VSS.n1694 VSS.n1693 0.121553
R1955 VSS.n1693 VSS.n1692 0.121553
R1956 VSS.n1692 VSS.n1691 0.121553
R1957 VSS.n1691 VSS.n1690 0.121553
R1958 VSS.n1690 VSS.n1689 0.121553
R1959 VSS.n1689 VSS.n1688 0.121553
R1960 VSS.n1688 VSS.n1687 0.121553
R1961 VSS.n1687 VSS.n1686 0.121553
R1962 VSS.n1487 VSS.n1486 0.120957
R1963 VSS.n1372 VSS.n1371 0.119346
R1964 VSS.n1529 VSS.n1527 0.119346
R1965 VSS.n362 VSS.n360 0.118395
R1966 VSS.n549 VSS.n546 0.118174
R1967 VSS.n811 VSS.n808 0.117688
R1968 VSS.n808 VSS.n805 0.117688
R1969 VSS.n805 VSS.n801 0.117688
R1970 VSS.n553 VSS.n550 0.117383
R1971 VSS.n1471 VSS.n1470 0.117038
R1972 VSS.n1453 VSS.n1452 0.116533
R1973 VSS.n37 VSS.n35 0.116289
R1974 VSS.n39 VSS.n37 0.116289
R1975 VSS.n49 VSS.n47 0.116289
R1976 VSS.n54 VSS.n52 0.116289
R1977 VSS.n59 VSS.n57 0.116289
R1978 VSS.n64 VSS.n62 0.116289
R1979 VSS.n69 VSS.n67 0.116289
R1980 VSS.n77 VSS.n74 0.116289
R1981 VSS.n83 VSS.n81 0.116289
R1982 VSS.n88 VSS.n86 0.116289
R1983 VSS.n1936 VSS.n1934 0.116289
R1984 VSS.n1938 VSS.n1936 0.116289
R1985 VSS.n1940 VSS.n1938 0.116289
R1986 VSS.n1948 VSS.n1944 0.116289
R1987 VSS.n1950 VSS.n1948 0.116289
R1988 VSS.n1958 VSS.n1956 0.116289
R1989 VSS.n1960 VSS.n1958 0.116289
R1990 VSS.n1962 VSS.n1960 0.116289
R1991 VSS.n1967 VSS.n1965 0.116289
R1992 VSS.n1969 VSS.n1967 0.116289
R1993 VSS.n1971 VSS.n1969 0.116289
R1994 VSS.n1977 VSS.n1975 0.116289
R1995 VSS.n1979 VSS.n1977 0.116289
R1996 VSS.n1982 VSS.n1979 0.116289
R1997 VSS.n1988 VSS.n1986 0.116289
R1998 VSS.n1990 VSS.n1988 0.116289
R1999 VSS.n1992 VSS.n1990 0.116289
R2000 VSS.n1951 VSS.n1950 0.115763
R2001 VSS.n645 VSS.n642 0.115458
R2002 VSS.n447 VSS.n444 0.115458
R2003 VSS.n350 VSS.n348 0.115237
R2004 VSS.n554 VSS.n553 0.115045
R2005 VSS.n1706 VSS.n1705 0.112423
R2006 VSS.n1592 VSS.n1591 0.112423
R2007 VSS.n798 VSS.n795 0.11207
R2008 VSS.n1319 VSS.n1318 0.111846
R2009 VSS.n50 VSS.n49 0.109974
R2010 VSS.n1501 VSS.n1499 0.109538
R2011 VSS.n1353 VSS.n1352 0.108962
R2012 VSS.n1311 VSS.n1310 0.108962
R2013 VSS.n86 VSS.n84 0.107868
R2014 VSS.n893 VSS.n890 0.107607
R2015 VSS.n299 VSS.n296 0.107607
R2016 VSS.n302 VSS.n299 0.107607
R2017 VSS.n305 VSS.n302 0.107607
R2018 VSS.n308 VSS.n305 0.107607
R2019 VSS.n659 VSS.n308 0.107607
R2020 VSS.n662 VSS.n659 0.107607
R2021 VSS.n665 VSS.n662 0.107607
R2022 VSS.n668 VSS.n665 0.107607
R2023 VSS.n671 VSS.n668 0.107607
R2024 VSS.n674 VSS.n671 0.107607
R2025 VSS.n677 VSS.n674 0.107607
R2026 VSS.n680 VSS.n677 0.107607
R2027 VSS.n683 VSS.n680 0.107607
R2028 VSS.n686 VSS.n683 0.107607
R2029 VSS.n689 VSS.n686 0.107607
R2030 VSS.n692 VSS.n689 0.107607
R2031 VSS.n695 VSS.n692 0.107607
R2032 VSS.n698 VSS.n695 0.107607
R2033 VSS.n701 VSS.n698 0.107607
R2034 VSS.n704 VSS.n701 0.107607
R2035 VSS.n707 VSS.n704 0.107607
R2036 VSS.n711 VSS.n707 0.107607
R2037 VSS.n378 VSS.n376 0.106816
R2038 VSS.n1363 VSS.n1362 0.106654
R2039 VSS.n1545 VSS.n1543 0.106654
R2040 VSS.n260 VSS.n258 0.10537
R2041 VSS.n1480 VSS.n1479 0.104346
R2042 VSS.n247 VSS.n243 0.104161
R2043 VSS.n149 VSS.n147 0.104161
R2044 VSS.n159 VSS.n157 0.104161
R2045 VSS.n167 VSS.n165 0.104161
R2046 VSS.n1885 VSS.n1881 0.104161
R2047 VSS.n1905 VSS.n1901 0.104161
R2048 VSS.n243 VSS.n238 0.103357
R2049 VSS.n169 VSS.n167 0.103357
R2050 VSS.n226 VSS.n221 0.102773
R2051 VSS.n1483 VSS.n1482 0.102038
R2052 VSS.n151 VSS.n149 0.10175
R2053 VSS.n1889 VSS.n1885 0.10175
R2054 VSS.n1360 VSS.n1359 0.0997308
R2055 VSS.n1552 VSS.n1551 0.0997308
R2056 VSS.n141 VSS.n139 0.0993393
R2057 VSS.n161 VSS.n159 0.0993393
R2058 VSS.n1869 VSS.n1865 0.0993393
R2059 VSS.n1909 VSS.n1905 0.0993393
R2060 VSS.n135 VSS.n133 0.0985357
R2061 VSS.n1858 VSS.n1854 0.0985357
R2062 VSS.n1818 VSS.n1814 0.0983261
R2063 VSS.n137 VSS.n135 0.0977321
R2064 VSS.n1842 VSS.n1838 0.0977321
R2065 VSS.n1862 VSS.n1858 0.0977321
R2066 VSS.n1314 VSS.n1313 0.0974231
R2067 VSS.n895 VSS.n893 0.0963383
R2068 VSS.n254 VSS.n252 0.096125
R2069 VSS.n131 VSS.n129 0.096125
R2070 VSS.n1838 VSS.n1834 0.096125
R2071 VSS.n1850 VSS.n1846 0.096125
R2072 VSS.n1662 VSS.n1661 0.0957632
R2073 VSS.n970 VSS.n967 0.0957326
R2074 VSS.n143 VSS.n141 0.0953214
R2075 VSS.n153 VSS.n151 0.0953214
R2076 VSS.n1873 VSS.n1869 0.0953214
R2077 VSS.n1893 VSS.n1889 0.0953214
R2078 VSS.n416 VSS.n415 0.0952368
R2079 VSS.n649 VSS.n646 0.094752
R2080 VSS.n441 VSS.n440 0.094752
R2081 VSS.n1717 VSS.n1716 0.0945385
R2082 VSS.n139 VSS.n137 0.0945179
R2083 VSS.n147 VSS.n145 0.0945179
R2084 VSS.n157 VSS.n155 0.0945179
R2085 VSS.n165 VSS.n163 0.0945179
R2086 VSS.n1865 VSS.n1862 0.0945179
R2087 VSS.n1881 VSS.n1877 0.0945179
R2088 VSS.n1901 VSS.n1897 0.0945179
R2089 VSS.n1354 VSS.n1353 0.0939615
R2090 VSS.n1707 VSS.n1706 0.0939615
R2091 VSS.n221 VSS.n219 0.0937727
R2092 VSS.n413 VSS.n412 0.0931316
R2093 VSS.n882 VSS.n868 0.093
R2094 VSS.n868 VSS.n866 0.093
R2095 VSS.n866 VSS.n863 0.093
R2096 VSS.n863 VSS.n860 0.093
R2097 VSS.n860 VSS.n858 0.093
R2098 VSS.n858 VSS.n855 0.093
R2099 VSS.n855 VSS.n853 0.093
R2100 VSS.n853 VSS.n850 0.093
R2101 VSS.n850 VSS.n848 0.093
R2102 VSS.n848 VSS.n845 0.093
R2103 VSS.n845 VSS.n843 0.093
R2104 VSS.n843 VSS.n840 0.093
R2105 VSS.n840 VSS.n838 0.093
R2106 VSS.n838 VSS.n836 0.093
R2107 VSS.n836 VSS.n834 0.093
R2108 VSS.n834 VSS.n832 0.093
R2109 VSS.n832 VSS.n830 0.093
R2110 VSS.n830 VSS.n828 0.093
R2111 VSS.n828 VSS.n826 0.093
R2112 VSS.n826 VSS.n824 0.093
R2113 VSS.n824 VSS.n822 0.093
R2114 VSS.n822 VSS.n820 0.093
R2115 VSS.n820 VSS.n818 0.093
R2116 VSS.n1176 VSS.n1174 0.093
R2117 VSS.n1178 VSS.n1176 0.093
R2118 VSS.n1180 VSS.n1178 0.093
R2119 VSS.n1182 VSS.n1180 0.093
R2120 VSS.n1184 VSS.n1182 0.093
R2121 VSS.n1186 VSS.n1184 0.093
R2122 VSS.n1188 VSS.n1186 0.093
R2123 VSS.n1190 VSS.n1188 0.093
R2124 VSS.n1192 VSS.n1190 0.093
R2125 VSS.n1195 VSS.n1192 0.093
R2126 VSS.n1197 VSS.n1195 0.093
R2127 VSS.n1200 VSS.n1197 0.093
R2128 VSS.n1202 VSS.n1200 0.093
R2129 VSS.n1205 VSS.n1202 0.093
R2130 VSS.n1207 VSS.n1205 0.093
R2131 VSS.n1210 VSS.n1207 0.093
R2132 VSS.n1212 VSS.n1210 0.093
R2133 VSS.n1216 VSS.n1212 0.093
R2134 VSS.n1048 VSS.n1046 0.093
R2135 VSS.n1050 VSS.n1048 0.093
R2136 VSS.n1052 VSS.n1050 0.093
R2137 VSS.n1055 VSS.n1052 0.093
R2138 VSS.n1058 VSS.n1055 0.093
R2139 VSS.n1061 VSS.n1058 0.093
R2140 VSS.n1064 VSS.n1061 0.093
R2141 VSS.n1067 VSS.n1064 0.093
R2142 VSS.n1070 VSS.n1067 0.093
R2143 VSS.n1073 VSS.n1070 0.093
R2144 VSS.n1076 VSS.n1073 0.093
R2145 VSS.n1079 VSS.n1076 0.093
R2146 VSS.n1082 VSS.n1079 0.093
R2147 VSS.n1085 VSS.n1082 0.093
R2148 VSS.n1088 VSS.n1085 0.093
R2149 VSS.n1091 VSS.n1088 0.093
R2150 VSS.n1093 VSS.n1091 0.093
R2151 VSS.n1099 VSS.n1093 0.093
R2152 VSS.n1794 VSS.n1791 0.093
R2153 VSS.n1791 VSS.n1788 0.093
R2154 VSS.n1788 VSS.n1785 0.093
R2155 VSS.n1785 VSS.n1782 0.093
R2156 VSS.n1782 VSS.n1779 0.093
R2157 VSS.n1779 VSS.n1776 0.093
R2158 VSS.n1776 VSS.n1773 0.093
R2159 VSS.n1773 VSS.n1770 0.093
R2160 VSS.n1770 VSS.n1767 0.093
R2161 VSS.n1767 VSS.n1764 0.093
R2162 VSS.n1764 VSS.n1761 0.093
R2163 VSS.n1761 VSS.n1758 0.093
R2164 VSS.n1758 VSS.n1755 0.093
R2165 VSS.n1755 VSS.n1753 0.093
R2166 VSS.n1753 VSS.n1750 0.093
R2167 VSS.n1750 VSS.n1749 0.093
R2168 VSS.n1749 VSS.n1746 0.093
R2169 VSS.n1746 VSS.n1743 0.093
R2170 VSS.n1743 VSS.n1740 0.093
R2171 VSS.n1740 VSS.n1738 0.093
R2172 VSS.n1291 VSS.n1104 0.093
R2173 VSS.n1293 VSS.n1291 0.093
R2174 VSS.n256 VSS.n254 0.0929107
R2175 VSS.n1834 VSS.n1830 0.0929107
R2176 VSS.n339 VSS.n338 0.0926987
R2177 VSS.n219 VSS.n217 0.0921364
R2178 VSS.n47 VSS.n43 0.0915526
R2179 VSS.n67 VSS.n65 0.0910263
R2180 VSS.n92 VSS.n91 0.0910263
R2181 VSS.n202 VSS.n199 0.0905
R2182 VSS.n185 VSS.n183 0.0905
R2183 VSS.n176 VSS.n174 0.0905
R2184 VSS.n129 VSS.n127 0.0905
R2185 VSS.n145 VSS.n143 0.0905
R2186 VSS.n155 VSS.n153 0.0905
R2187 VSS.n163 VSS.n161 0.0905
R2188 VSS.n1846 VSS.n1842 0.0905
R2189 VSS.n1877 VSS.n1873 0.0905
R2190 VSS.n1897 VSS.n1893 0.0905
R2191 VSS.n716 VSS.n714 0.0897562
R2192 VSS.n718 VSS.n716 0.0897562
R2193 VSS.n720 VSS.n718 0.0897562
R2194 VSS.n723 VSS.n720 0.0897562
R2195 VSS.n726 VSS.n723 0.0897562
R2196 VSS.n729 VSS.n726 0.0897562
R2197 VSS.n732 VSS.n729 0.0897562
R2198 VSS.n735 VSS.n732 0.0897562
R2199 VSS.n738 VSS.n735 0.0897562
R2200 VSS.n741 VSS.n738 0.0897562
R2201 VSS.n744 VSS.n741 0.0897562
R2202 VSS.n747 VSS.n744 0.0897562
R2203 VSS.n750 VSS.n747 0.0897562
R2204 VSS.n753 VSS.n750 0.0897562
R2205 VSS.n756 VSS.n753 0.0897562
R2206 VSS.n759 VSS.n756 0.0897562
R2207 VSS.n762 VSS.n759 0.0897562
R2208 VSS.n768 VSS.n762 0.0897562
R2209 VSS.n771 VSS.n768 0.0897562
R2210 VSS.n773 VSS.n771 0.0897562
R2211 VSS.n776 VSS.n773 0.0897562
R2212 VSS.n779 VSS.n776 0.0897562
R2213 VSS.n782 VSS.n779 0.0897562
R2214 VSS.n785 VSS.n782 0.0897562
R2215 VSS.n788 VSS.n785 0.0897562
R2216 VSS.n791 VSS.n788 0.0897562
R2217 VSS.n795 VSS.n791 0.0897562
R2218 VSS.n1814 VSS.n1812 0.0897174
R2219 VSS.n133 VSS.n131 0.0896964
R2220 VSS.n1854 VSS.n1850 0.0896964
R2221 VSS.n209 VSS.n207 0.0896818
R2222 VSS.n1474 VSS.n1473 0.0893462
R2223 VSS.n42 VSS.n40 0.0889211
R2224 VSS.n228 VSS.n226 0.0888636
R2225 VSS.n1738 VSS.n1735 0.0888333
R2226 VSS.n1812 VSS.n1809 0.0881522
R2227 VSS.n1916 VSS.n125 0.0873421
R2228 VSS.n1369 VSS.n1368 0.0870385
R2229 VSS.n1534 VSS.n1533 0.0870385
R2230 VSS.n91 VSS.n89 0.0868158
R2231 VSS.n291 VSS.n288 0.086587
R2232 VSS.n274 VSS.n272 0.086587
R2233 VSS.n265 VSS.n263 0.086587
R2234 VSS.n1801 VSS.n1799 0.0858043
R2235 VSS.n217 VSS.n214 0.0855909
R2236 VSS.n214 VSS.n211 0.0855909
R2237 VSS.n207 VSS.n204 0.0855909
R2238 VSS.n199 VSS.n195 0.0855909
R2239 VSS.n190 VSS.n187 0.0855909
R2240 VSS.n183 VSS.n180 0.0855909
R2241 VSS.n178 VSS.n176 0.0855909
R2242 VSS.n174 VSS.n171 0.0855909
R2243 VSS.n1820 VSS.n1818 0.0850217
R2244 VSS.n1119 VSS.n1117 0.0847308
R2245 VSS.n884 VSS.n882 0.0838333
R2246 VSS.n407 VSS.n406 0.0836579
R2247 VSS.n233 VSS.n230 0.0831364
R2248 VSS.n193 VSS.n190 0.0831364
R2249 VSS.n1944 VSS.n1941 0.0831316
R2250 VSS.n1795 VSS.n1794 0.083
R2251 VSS.n814 VSS.n812 0.0828529
R2252 VSS.n1965 VSS.n1963 0.0826053
R2253 VSS.n967 VSS.n966 0.0824863
R2254 VSS.n1809 VSS.n1806 0.0818913
R2255 VSS.n1806 VSS.n1803 0.0818913
R2256 VSS.n288 VSS.n284 0.0818913
R2257 VSS.n279 VSS.n276 0.0818913
R2258 VSS.n272 VSS.n269 0.0818913
R2259 VSS.n267 VSS.n265 0.0818913
R2260 VSS.n263 VSS.n260 0.0818913
R2261 VSS.n383 VSS.n382 0.0815526
R2262 VSS.n1116 VSS.n1107 0.0812692
R2263 VSS.n230 VSS.n228 0.0798636
R2264 VSS.n1825 VSS.n1822 0.0795435
R2265 VSS.n282 VSS.n279 0.0795435
R2266 VSS.n1986 VSS.n1983 0.0783947
R2267 VSS.n211 VSS.n209 0.0782273
R2268 VSS.n204 VSS.n202 0.0782273
R2269 VSS.n195 VSS.n193 0.0782273
R2270 VSS.n187 VSS.n185 0.0782273
R2271 VSS.n180 VSS.n178 0.0782273
R2272 VSS.n1465 VSS.n1464 0.0766538
R2273 VSS.n1822 VSS.n1820 0.076413
R2274 VSS.n654 VSS.n314 0.0763268
R2275 VSS.n431 VSS.n430 0.0763268
R2276 VSS.n60 VSS.n59 0.0762895
R2277 VSS.n1826 VSS.n1825 0.0756304
R2278 VSS.n237 VSS.n234 0.0749681
R2279 VSS VSS.n653 0.0749094
R2280 VSS.n436 VSS 0.0749094
R2281 VSS.n1803 VSS.n1801 0.0748478
R2282 VSS.n293 VSS.n291 0.0748478
R2283 VSS.n284 VSS.n282 0.0748478
R2284 VSS.n276 VSS.n274 0.0748478
R2285 VSS.n269 VSS.n267 0.0748478
R2286 VSS.n897 VSS.n895 0.0744726
R2287 VSS.n899 VSS.n897 0.0744726
R2288 VSS.n901 VSS.n899 0.0744726
R2289 VSS.n903 VSS.n901 0.0744726
R2290 VSS.n905 VSS.n903 0.0744726
R2291 VSS.n907 VSS.n905 0.0744726
R2292 VSS.n910 VSS.n907 0.0744726
R2293 VSS.n912 VSS.n910 0.0744726
R2294 VSS.n915 VSS.n912 0.0744726
R2295 VSS.n917 VSS.n915 0.0744726
R2296 VSS.n920 VSS.n917 0.0744726
R2297 VSS.n922 VSS.n920 0.0744726
R2298 VSS.n925 VSS.n922 0.0744726
R2299 VSS.n928 VSS.n925 0.0744726
R2300 VSS.n930 VSS.n928 0.0744726
R2301 VSS.n933 VSS.n930 0.0744726
R2302 VSS.n935 VSS.n933 0.0744726
R2303 VSS.n942 VSS.n935 0.0744726
R2304 VSS.n945 VSS.n942 0.0744726
R2305 VSS.n947 VSS.n945 0.0744726
R2306 VSS.n950 VSS.n947 0.0744726
R2307 VSS.n952 VSS.n950 0.0744726
R2308 VSS.n955 VSS.n952 0.0744726
R2309 VSS.n957 VSS.n955 0.0744726
R2310 VSS.n960 VSS.n957 0.0744726
R2311 VSS.n962 VSS.n960 0.0744726
R2312 VSS.n966 VSS.n962 0.0744726
R2313 VSS.n1378 VSS.n1377 0.0743462
R2314 VSS.n1518 VSS.n1517 0.0743462
R2315 VSS.n1588 VSS.n1146 0.0743462
R2316 VSS.n74 VSS.n70 0.0741842
R2317 VSS.n1725 VSS.n1131 0.0726154
R2318 VSS.n1972 VSS.n1971 0.0720789
R2319 VSS.n1386 VSS.n1385 0.0720385
R2320 VSS.n1504 VSS.n1502 0.0720385
R2321 VSS.n1723 VSS.n1722 0.0720385
R2322 VSS.n885 VSS.n884 0.0713333
R2323 VSS.n367 VSS.n366 0.0699737
R2324 VSS.n1457 VSS.n1456 0.0697308
R2325 VSS.n420 VSS.n419 0.0694474
R2326 VSS VSS.n1566 0.0689956
R2327 VSS.n1712 VSS 0.0689956
R2328 VSS VSS.n1730 0.0689956
R2329 VSS.n1148 VSS 0.0689956
R2330 VSS VSS.n1714 0.0689956
R2331 VSS VSS.n1567 0.0689956
R2332 VSS.n171 VSS.n169 0.0689789
R2333 VSS.n714 VSS.n711 0.068186
R2334 VSS.n1954 VSS.n1953 0.0678684
R2335 VSS.n654 VSS 0.0678228
R2336 VSS.n431 VSS 0.0678228
R2337 VSS.n801 VSS.n798 0.0648001
R2338 VSS.n1456 VSS.n1455 0.0639615
R2339 VSS.n78 VSS.n77 0.0636579
R2340 VSS.n353 VSS.n351 0.0636579
R2341 VSS.n1614 VSS.n1612 0.062959
R2342 VSS.n1929 VSS.n1928 0.0624089
R2343 VSS.n1387 VSS.n1386 0.0616538
R2344 VSS.n1502 VSS.n1501 0.0616538
R2345 VSS.n1724 VSS.n1723 0.0616538
R2346 VSS.n30 VSS.n29 0.0615526
R2347 VSS.n1725 VSS.n1724 0.0610769
R2348 VSS.n238 VSS.n233 0.0607533
R2349 VSS.n55 VSS.n54 0.0594474
R2350 VSS.n1377 VSS.n1376 0.0593462
R2351 VSS.n1520 VSS.n1518 0.0593462
R2352 VSS.n1589 VSS.n1588 0.0593462
R2353 VSS.n33 VSS.n32 0.058921
R2354 VSS.n351 VSS.n350 0.0583947
R2355 VSS.n35 VSS.n33 0.0578684
R2356 VSS.n57 VSS.n55 0.0573421
R2357 VSS.n1466 VSS.n1465 0.0570385
R2358 VSS.n32 VSS.n30 0.0552368
R2359 VSS.n258 VSS.n256 0.05508
R2360 VSS.n81 VSS.n78 0.0531316
R2361 VSS.n1910 VSS.n1909 0.0527321
R2362 VSS.n420 VSS.n385 0.0526053
R2363 VSS.n1307 VSS.n1107 0.0524231
R2364 VSS.n369 VSS.n367 0.052079
R2365 VSS.n1830 VSS.n1826 0.0503214
R2366 VSS.n1934 VSS.n1932 0.0494474
R2367 VSS.n1117 VSS.n1116 0.0489615
R2368 VSS.n1956 VSS.n1954 0.0489211
R2369 VSS.n646 VSS.n645 0.0479803
R2370 VSS.n444 VSS.n441 0.0479803
R2371 VSS.n1368 VSS.n1367 0.0466538
R2372 VSS.n1536 VSS.n1534 0.0466538
R2373 VSS.n1975 VSS.n1972 0.0447105
R2374 VSS.n1475 VSS.n1474 0.0443462
R2375 VSS.n70 VSS.n69 0.0426053
R2376 VSS.n1799 VSS.n1796 0.0411957
R2377 VSS.n1796 VSS.n293 0.0411957
R2378 VSS.n62 VSS.n60 0.0405
R2379 VSS.n385 VSS.n383 0.0405
R2380 VSS.n1355 VSS.n1354 0.0397308
R2381 VSS.n1708 VSS.n1707 0.0397308
R2382 VSS.n1716 VSS.n1146 0.0391538
R2383 VSS.n1983 VSS.n1982 0.0383947
R2384 VSS.n408 VSS.n407 0.0383947
R2385 VSS.n1910 VSS.n247 0.0366607
R2386 VSS.n1315 VSS.n1314 0.0362692
R2387 VSS.n1917 VSS.n1916 0.0347105
R2388 VSS.n1963 VSS.n1962 0.0341842
R2389 VSS.n1359 VSS.n1358 0.0339615
R2390 VSS.n1551 VSS.n1550 0.0339615
R2391 VSS.n1941 VSS.n1940 0.0336579
R2392 VSS.n1484 VSS.n1483 0.0316538
R2393 VSS.n89 VSS.n88 0.0299737
R2394 VSS.n1479 VSS.n1478 0.0293462
R2395 VSS.n412 VSS.n411 0.0289211
R2396 VSS.n40 VSS.n39 0.0278684
R2397 VSS.n1364 VSS.n1363 0.0270385
R2398 VSS.n1543 VSS.n1542 0.0270385
R2399 VSS.n417 VSS.n416 0.0268158
R2400 VSS.n1664 VSS.n1662 0.0262895
R2401 VSS.n65 VSS.n64 0.0257632
R2402 VSS.n94 VSS.n92 0.0257632
R2403 VSS.n967 VSS.n886 0.0257083
R2404 VSS.n43 VSS.n42 0.0252368
R2405 VSS.n1352 VSS.n1351 0.0247308
R2406 VSS.n1310 VSS.n1309 0.0247308
R2407 VSS.n1395 VSS.n1391 0.0241538
R2408 VSS.n1499 VSS.n1498 0.0241538
R2409 VSS.n347 VSS.n340 0.0231316
R2410 VSS.n1320 VSS.n1319 0.0218462
R2411 VSS.n1705 VSS.n1704 0.0212692
R2412 VSS.n1593 VSS.n1592 0.0212692
R2413 VSS.n1470 VSS.n1469 0.0166538
R2414 VSS.n376 VSS.n375 0.0152368
R2415 VSS.n1043 VSS.n1042 0.0151318
R2416 VSS.n1373 VSS.n1372 0.0143462
R2417 VSS.n1527 VSS.n1526 0.0143462
R2418 VSS.n1043 VSS.n811 0.013625
R2419 VSS.n340 VSS.n339 0.0128813
R2420 VSS.n1389 VSS.n1388 0.0122131
R2421 VSS.n1126 VSS.n1124 0.0120385
R2422 VSS.n1488 VSS.n1487 0.0119467
R2423 VSS.n1294 VSS.n1288 0.0109651
R2424 VSS.n1321 VSS.n1168 0.0108811
R2425 VSS.n1452 VSS.n1446 0.0106146
R2426 VSS.n1795 VSS.n1099 0.0105
R2427 VSS.n1444 VSS.n1443 0.00973077
R2428 VSS.n653 VSS.n650 0.0097126
R2429 VSS.n437 VSS.n436 0.0097126
R2430 VSS.n1317 VSS.n1316 0.00915385
R2431 VSS.n84 VSS.n83 0.00892105
R2432 VSS VSS.n94 0.00892105
R2433 VSS.n1446 VSS.n1444 0.008
R2434 VSS.n1704 VSS.n1703 0.008
R2435 VSS.n1594 VSS.n1593 0.00742308
R2436 VSS.n1321 VSS.n1320 0.00684615
R2437 VSS.n52 VSS.n50 0.00681579
R2438 VSS.n348 VSS.n347 0.00681579
R2439 VSS.n1993 VSS.n1992 0.00471053
R2440 VSS.n1735 VSS.n1104 0.00466667
R2441 VSS.n1595 VSS.n1594 0.00420487
R2442 VSS.n1461 VSS.n1460 0.00396154
R2443 VSS.n360 VSS.n359 0.00365789
R2444 VSS.n557 VSS.n554 0.00283766
R2445 VSS.n1914 VSS.n1910 0.00276891
R2446 VSS.n1488 VSS.n1395 0.00223077
R2447 VSS.n1382 VSS.n1381 0.00165385
R2448 VSS.n1351 VSS.n1350 0.00165385
R2449 VSS.n1498 VSS.n1495 0.00165385
R2450 VSS.n1511 VSS.n1510 0.00165385
R2451 VSS VSS.n1719 0.00165385
R2452 VSS.n1638 VSS 0.00129646
R2453 VSS.n1640 VSS 0.00129646
R2454 VSS.n1733 VSS 0.00129646
R2455 VSS.n1728 VSS 0.00129646
R2456 VSS VSS.n1556 0.00129646
R2457 VSS.n1644 VSS 0.00129646
R2458 VSS.n1389 VSS.n1324 0.00107692
R2459 VSS.n1953 VSS.n1951 0.00102632
R2460 SEL_L.n46 SEL_L.n45 59.4622
R2461 SEL_L.n94 SEL_L.n93 58.2146
R2462 SEL_L.n0 SEL_L.t100 51.4916
R2463 SEL_L.n48 SEL_L.t12 51.4916
R2464 SEL_L.n7 SEL_L.t29 48.0881
R2465 SEL_L.n55 SEL_L.t56 48.0881
R2466 SEL_L.n4 SEL_L.t78 43.2791
R2467 SEL_L.n3 SEL_L.t84 43.2791
R2468 SEL_L.n2 SEL_L.t76 43.2791
R2469 SEL_L.n1 SEL_L.t9 43.2791
R2470 SEL_L.n52 SEL_L.t94 43.2791
R2471 SEL_L.n51 SEL_L.t98 43.2791
R2472 SEL_L.n50 SEL_L.t92 43.2791
R2473 SEL_L.n49 SEL_L.t22 43.2791
R2474 SEL_L.n7 SEL_L.t31 34.2844
R2475 SEL_L.n8 SEL_L.t27 34.2844
R2476 SEL_L.n9 SEL_L.t53 34.2844
R2477 SEL_L.n10 SEL_L.t59 34.2844
R2478 SEL_L.n11 SEL_L.t86 34.2844
R2479 SEL_L.n12 SEL_L.t89 34.2844
R2480 SEL_L.n13 SEL_L.t16 34.2844
R2481 SEL_L.n14 SEL_L.t43 34.2844
R2482 SEL_L.n15 SEL_L.t46 34.2844
R2483 SEL_L.n16 SEL_L.t71 34.2844
R2484 SEL_L.n17 SEL_L.t74 34.2844
R2485 SEL_L.n18 SEL_L.t5 34.2844
R2486 SEL_L.n19 SEL_L.t36 34.2844
R2487 SEL_L.n20 SEL_L.t23 34.2844
R2488 SEL_L.n21 SEL_L.t85 34.2844
R2489 SEL_L.n22 SEL_L.t79 34.2844
R2490 SEL_L.n23 SEL_L.t51 34.2844
R2491 SEL_L.n24 SEL_L.t25 34.2844
R2492 SEL_L.n25 SEL_L.t19 34.2844
R2493 SEL_L.n26 SEL_L.t91 34.2844
R2494 SEL_L.n27 SEL_L.t83 34.2844
R2495 SEL_L.n28 SEL_L.t57 34.2844
R2496 SEL_L.n29 SEL_L.t30 34.2844
R2497 SEL_L.n30 SEL_L.t24 34.2844
R2498 SEL_L.n31 SEL_L.t93 34.2844
R2499 SEL_L.n32 SEL_L.t90 34.2844
R2500 SEL_L.n33 SEL_L.t96 34.2844
R2501 SEL_L.n34 SEL_L.t63 34.2844
R2502 SEL_L.n35 SEL_L.t61 34.2844
R2503 SEL_L.n36 SEL_L.t34 34.2844
R2504 SEL_L.n37 SEL_L.t32 34.2844
R2505 SEL_L.n38 SEL_L.t101 34.2844
R2506 SEL_L.n39 SEL_L.t2 34.2844
R2507 SEL_L.n40 SEL_L.t102 34.2844
R2508 SEL_L.n41 SEL_L.t70 34.2844
R2509 SEL_L.n42 SEL_L.t67 34.2844
R2510 SEL_L.n43 SEL_L.t42 34.2844
R2511 SEL_L.n44 SEL_L.t11 34.2844
R2512 SEL_L.n55 SEL_L.t60 34.2844
R2513 SEL_L.n56 SEL_L.t54 34.2844
R2514 SEL_L.n57 SEL_L.t80 34.2844
R2515 SEL_L.n58 SEL_L.t87 34.2844
R2516 SEL_L.n59 SEL_L.t14 34.2844
R2517 SEL_L.n60 SEL_L.t17 34.2844
R2518 SEL_L.n61 SEL_L.t48 34.2844
R2519 SEL_L.n62 SEL_L.t69 34.2844
R2520 SEL_L.n63 SEL_L.t72 34.2844
R2521 SEL_L.n64 SEL_L.t0 34.2844
R2522 SEL_L.n65 SEL_L.t7 34.2844
R2523 SEL_L.n66 SEL_L.t37 34.2844
R2524 SEL_L.n67 SEL_L.t62 34.2844
R2525 SEL_L.n68 SEL_L.t49 34.2844
R2526 SEL_L.n69 SEL_L.t99 34.2844
R2527 SEL_L.n70 SEL_L.t95 34.2844
R2528 SEL_L.n71 SEL_L.t64 34.2844
R2529 SEL_L.n72 SEL_L.t38 34.2844
R2530 SEL_L.n73 SEL_L.t33 34.2844
R2531 SEL_L.n74 SEL_L.t1 34.2844
R2532 SEL_L.n75 SEL_L.t97 34.2844
R2533 SEL_L.n76 SEL_L.t66 34.2844
R2534 SEL_L.n77 SEL_L.t41 34.2844
R2535 SEL_L.n78 SEL_L.t35 34.2844
R2536 SEL_L.n79 SEL_L.t4 34.2844
R2537 SEL_L.n80 SEL_L.t103 34.2844
R2538 SEL_L.n81 SEL_L.t8 34.2844
R2539 SEL_L.n82 SEL_L.t75 34.2844
R2540 SEL_L.n83 SEL_L.t73 34.2844
R2541 SEL_L.n84 SEL_L.t47 34.2844
R2542 SEL_L.n85 SEL_L.t44 34.2844
R2543 SEL_L.n86 SEL_L.t13 34.2844
R2544 SEL_L.n87 SEL_L.t18 34.2844
R2545 SEL_L.n88 SEL_L.t15 34.2844
R2546 SEL_L.n89 SEL_L.t88 34.2844
R2547 SEL_L.n90 SEL_L.t81 34.2844
R2548 SEL_L.n91 SEL_L.t55 34.2844
R2549 SEL_L.n92 SEL_L.t28 34.2844
R2550 SEL_L.n6 SEL_L.t3 30.6344
R2551 SEL_L.n5 SEL_L.t10 30.6344
R2552 SEL_L.n4 SEL_L.t40 30.6344
R2553 SEL_L.n3 SEL_L.t45 30.6344
R2554 SEL_L.n2 SEL_L.t39 30.6344
R2555 SEL_L.n1 SEL_L.t65 30.6344
R2556 SEL_L.n0 SEL_L.t68 30.6344
R2557 SEL_L.n54 SEL_L.t20 30.6344
R2558 SEL_L.n53 SEL_L.t26 30.6344
R2559 SEL_L.n52 SEL_L.t52 30.6344
R2560 SEL_L.n51 SEL_L.t58 30.6344
R2561 SEL_L.n50 SEL_L.t50 30.6344
R2562 SEL_L.n49 SEL_L.t77 30.6344
R2563 SEL_L.n48 SEL_L.t82 30.6344
R2564 SEL_L.n45 SEL_L.t6 30.5041
R2565 SEL_L.n93 SEL_L.t21 30.5041
R2566 SEL_L.n46 SEL_L.n6 23.6891
R2567 SEL_L.n94 SEL_L.n54 23.6891
R2568 SEL_L.n6 SEL_L.n5 20.8576
R2569 SEL_L.n5 SEL_L.n4 20.8576
R2570 SEL_L.n4 SEL_L.n3 20.8576
R2571 SEL_L.n3 SEL_L.n2 20.8576
R2572 SEL_L.n2 SEL_L.n1 20.8576
R2573 SEL_L.n1 SEL_L.n0 20.8576
R2574 SEL_L.n54 SEL_L.n53 20.8576
R2575 SEL_L.n53 SEL_L.n52 20.8576
R2576 SEL_L.n52 SEL_L.n51 20.8576
R2577 SEL_L.n51 SEL_L.n50 20.8576
R2578 SEL_L.n50 SEL_L.n49 20.8576
R2579 SEL_L.n49 SEL_L.n48 20.8576
R2580 SEL_L.n45 SEL_L.n44 17.4541
R2581 SEL_L.n93 SEL_L.n92 17.4541
R2582 SEL_L.n8 SEL_L.n7 13.8041
R2583 SEL_L.n9 SEL_L.n8 13.8041
R2584 SEL_L.n10 SEL_L.n9 13.8041
R2585 SEL_L.n11 SEL_L.n10 13.8041
R2586 SEL_L.n12 SEL_L.n11 13.8041
R2587 SEL_L.n13 SEL_L.n12 13.8041
R2588 SEL_L.n14 SEL_L.n13 13.8041
R2589 SEL_L.n15 SEL_L.n14 13.8041
R2590 SEL_L.n16 SEL_L.n15 13.8041
R2591 SEL_L.n17 SEL_L.n16 13.8041
R2592 SEL_L.n18 SEL_L.n17 13.8041
R2593 SEL_L.n19 SEL_L.n18 13.8041
R2594 SEL_L.n20 SEL_L.n19 13.8041
R2595 SEL_L.n21 SEL_L.n20 13.8041
R2596 SEL_L.n22 SEL_L.n21 13.8041
R2597 SEL_L.n23 SEL_L.n22 13.8041
R2598 SEL_L.n24 SEL_L.n23 13.8041
R2599 SEL_L.n25 SEL_L.n24 13.8041
R2600 SEL_L.n26 SEL_L.n25 13.8041
R2601 SEL_L.n27 SEL_L.n26 13.8041
R2602 SEL_L.n28 SEL_L.n27 13.8041
R2603 SEL_L.n29 SEL_L.n28 13.8041
R2604 SEL_L.n30 SEL_L.n29 13.8041
R2605 SEL_L.n31 SEL_L.n30 13.8041
R2606 SEL_L.n32 SEL_L.n31 13.8041
R2607 SEL_L.n33 SEL_L.n32 13.8041
R2608 SEL_L.n34 SEL_L.n33 13.8041
R2609 SEL_L.n35 SEL_L.n34 13.8041
R2610 SEL_L.n36 SEL_L.n35 13.8041
R2611 SEL_L.n37 SEL_L.n36 13.8041
R2612 SEL_L.n38 SEL_L.n37 13.8041
R2613 SEL_L.n39 SEL_L.n38 13.8041
R2614 SEL_L.n40 SEL_L.n39 13.8041
R2615 SEL_L.n41 SEL_L.n40 13.8041
R2616 SEL_L.n42 SEL_L.n41 13.8041
R2617 SEL_L.n43 SEL_L.n42 13.8041
R2618 SEL_L.n44 SEL_L.n43 13.8041
R2619 SEL_L.n56 SEL_L.n55 13.8041
R2620 SEL_L.n57 SEL_L.n56 13.8041
R2621 SEL_L.n58 SEL_L.n57 13.8041
R2622 SEL_L.n59 SEL_L.n58 13.8041
R2623 SEL_L.n60 SEL_L.n59 13.8041
R2624 SEL_L.n61 SEL_L.n60 13.8041
R2625 SEL_L.n62 SEL_L.n61 13.8041
R2626 SEL_L.n63 SEL_L.n62 13.8041
R2627 SEL_L.n64 SEL_L.n63 13.8041
R2628 SEL_L.n65 SEL_L.n64 13.8041
R2629 SEL_L.n66 SEL_L.n65 13.8041
R2630 SEL_L.n67 SEL_L.n66 13.8041
R2631 SEL_L.n68 SEL_L.n67 13.8041
R2632 SEL_L.n69 SEL_L.n68 13.8041
R2633 SEL_L.n70 SEL_L.n69 13.8041
R2634 SEL_L.n71 SEL_L.n70 13.8041
R2635 SEL_L.n72 SEL_L.n71 13.8041
R2636 SEL_L.n73 SEL_L.n72 13.8041
R2637 SEL_L.n74 SEL_L.n73 13.8041
R2638 SEL_L.n75 SEL_L.n74 13.8041
R2639 SEL_L.n76 SEL_L.n75 13.8041
R2640 SEL_L.n77 SEL_L.n76 13.8041
R2641 SEL_L.n78 SEL_L.n77 13.8041
R2642 SEL_L.n79 SEL_L.n78 13.8041
R2643 SEL_L.n80 SEL_L.n79 13.8041
R2644 SEL_L.n81 SEL_L.n80 13.8041
R2645 SEL_L.n82 SEL_L.n81 13.8041
R2646 SEL_L.n83 SEL_L.n82 13.8041
R2647 SEL_L.n84 SEL_L.n83 13.8041
R2648 SEL_L.n85 SEL_L.n84 13.8041
R2649 SEL_L.n86 SEL_L.n85 13.8041
R2650 SEL_L.n87 SEL_L.n86 13.8041
R2651 SEL_L.n88 SEL_L.n87 13.8041
R2652 SEL_L.n89 SEL_L.n88 13.8041
R2653 SEL_L.n90 SEL_L.n89 13.8041
R2654 SEL_L.n91 SEL_L.n90 13.8041
R2655 SEL_L.n92 SEL_L.n91 13.8041
R2656 SEL_L SEL_L.n47 3.33134
R2657 SEL_L.n47 SEL_L 2.52957
R2658 SEL_L.n47 SEL_L 2.05983
R2659 SEL_L SEL_L.n46 0.00592169
R2660 SEL_L SEL_L.n94 0.00495545
R2661 OUT+.n99 OUT+.n96 3.81941
R2662 OUT+.n94 OUT+.n91 3.81941
R2663 OUT+.n89 OUT+.n86 3.81941
R2664 OUT+.n84 OUT+.n81 3.81941
R2665 OUT+.n79 OUT+.n76 3.81941
R2666 OUT+.n74 OUT+.n71 3.81941
R2667 OUT+.n69 OUT+.n66 3.81941
R2668 OUT+.n64 OUT+.n61 3.81941
R2669 OUT+.n59 OUT+.n56 3.81941
R2670 OUT+.n54 OUT+.n51 3.81941
R2671 OUT+.n49 OUT+.n46 3.81941
R2672 OUT+.n44 OUT+.n41 3.81941
R2673 OUT+.n39 OUT+.n36 3.81941
R2674 OUT+.n34 OUT+.n31 3.81941
R2675 OUT+.n29 OUT+.n26 3.81941
R2676 OUT+.n24 OUT+.n21 3.81941
R2677 OUT+.n19 OUT+.n16 3.81941
R2678 OUT+.n14 OUT+.n11 3.81941
R2679 OUT+.n9 OUT+.n6 3.81941
R2680 OUT+.n4 OUT+.n1 3.81941
R2681 OUT+.n99 OUT+.n98 3.1505
R2682 OUT+.n94 OUT+.n93 3.1505
R2683 OUT+.n89 OUT+.n88 3.1505
R2684 OUT+.n84 OUT+.n83 3.1505
R2685 OUT+.n79 OUT+.n78 3.1505
R2686 OUT+.n74 OUT+.n73 3.1505
R2687 OUT+.n69 OUT+.n68 3.1505
R2688 OUT+.n64 OUT+.n63 3.1505
R2689 OUT+.n59 OUT+.n58 3.1505
R2690 OUT+.n54 OUT+.n53 3.1505
R2691 OUT+.n49 OUT+.n48 3.1505
R2692 OUT+.n44 OUT+.n43 3.1505
R2693 OUT+.n39 OUT+.n38 3.1505
R2694 OUT+.n34 OUT+.n33 3.1505
R2695 OUT+.n29 OUT+.n28 3.1505
R2696 OUT+.n24 OUT+.n23 3.1505
R2697 OUT+.n19 OUT+.n18 3.1505
R2698 OUT+.n14 OUT+.n13 3.1505
R2699 OUT+.n9 OUT+.n8 3.1505
R2700 OUT+.n4 OUT+.n3 3.1505
R2701 OUT+.n96 OUT+.t56 0.9105
R2702 OUT+.n96 OUT+.n95 0.9105
R2703 OUT+.n91 OUT+.t71 0.9105
R2704 OUT+.n91 OUT+.n90 0.9105
R2705 OUT+.n86 OUT+.t65 0.9105
R2706 OUT+.n86 OUT+.n85 0.9105
R2707 OUT+.n81 OUT+.t55 0.9105
R2708 OUT+.n81 OUT+.n80 0.9105
R2709 OUT+.n76 OUT+.t8 0.9105
R2710 OUT+.n76 OUT+.n75 0.9105
R2711 OUT+.n71 OUT+.t54 0.9105
R2712 OUT+.n71 OUT+.n70 0.9105
R2713 OUT+.n66 OUT+.t75 0.9105
R2714 OUT+.n66 OUT+.n65 0.9105
R2715 OUT+.n61 OUT+.t5 0.9105
R2716 OUT+.n61 OUT+.n60 0.9105
R2717 OUT+.n56 OUT+.t7 0.9105
R2718 OUT+.n56 OUT+.n55 0.9105
R2719 OUT+.n51 OUT+.t0 0.9105
R2720 OUT+.n51 OUT+.n50 0.9105
R2721 OUT+.n46 OUT+.t58 0.9105
R2722 OUT+.n46 OUT+.n45 0.9105
R2723 OUT+.n41 OUT+.t50 0.9105
R2724 OUT+.n41 OUT+.n40 0.9105
R2725 OUT+.n36 OUT+.t1 0.9105
R2726 OUT+.n36 OUT+.n35 0.9105
R2727 OUT+.n31 OUT+.t49 0.9105
R2728 OUT+.n31 OUT+.n30 0.9105
R2729 OUT+.n26 OUT+.t74 0.9105
R2730 OUT+.n26 OUT+.n25 0.9105
R2731 OUT+.n21 OUT+.t53 0.9105
R2732 OUT+.n21 OUT+.n20 0.9105
R2733 OUT+.n16 OUT+.t68 0.9105
R2734 OUT+.n16 OUT+.n15 0.9105
R2735 OUT+.n11 OUT+.t77 0.9105
R2736 OUT+.n11 OUT+.n10 0.9105
R2737 OUT+.n6 OUT+.t62 0.9105
R2738 OUT+.n6 OUT+.n5 0.9105
R2739 OUT+.n1 OUT+.t73 0.9105
R2740 OUT+.n1 OUT+.n0 0.9105
R2741 OUT+.n98 OUT+.t38 0.8195
R2742 OUT+.n98 OUT+.n97 0.8195
R2743 OUT+.n93 OUT+.t26 0.8195
R2744 OUT+.n93 OUT+.n92 0.8195
R2745 OUT+.n88 OUT+.t13 0.8195
R2746 OUT+.n88 OUT+.n87 0.8195
R2747 OUT+.n83 OUT+.t39 0.8195
R2748 OUT+.n83 OUT+.n82 0.8195
R2749 OUT+.n78 OUT+.t31 0.8195
R2750 OUT+.n78 OUT+.n77 0.8195
R2751 OUT+.n73 OUT+.t18 0.8195
R2752 OUT+.n73 OUT+.n72 0.8195
R2753 OUT+.n68 OUT+.t44 0.8195
R2754 OUT+.n68 OUT+.n67 0.8195
R2755 OUT+.n63 OUT+.t46 0.8195
R2756 OUT+.n63 OUT+.n62 0.8195
R2757 OUT+.n58 OUT+.t32 0.8195
R2758 OUT+.n58 OUT+.n57 0.8195
R2759 OUT+.n53 OUT+.t11 0.8195
R2760 OUT+.n53 OUT+.n52 0.8195
R2761 OUT+.n48 OUT+.t36 0.8195
R2762 OUT+.n48 OUT+.n47 0.8195
R2763 OUT+.n43 OUT+.t22 0.8195
R2764 OUT+.n43 OUT+.n42 0.8195
R2765 OUT+.n38 OUT+.t10 0.8195
R2766 OUT+.n38 OUT+.n37 0.8195
R2767 OUT+.n33 OUT+.t23 0.8195
R2768 OUT+.n33 OUT+.n32 0.8195
R2769 OUT+.n28 OUT+.t45 0.8195
R2770 OUT+.n28 OUT+.n27 0.8195
R2771 OUT+.n23 OUT+.t19 0.8195
R2772 OUT+.n23 OUT+.n22 0.8195
R2773 OUT+.n18 OUT+.t29 0.8195
R2774 OUT+.n18 OUT+.n17 0.8195
R2775 OUT+.n13 OUT+.t42 0.8195
R2776 OUT+.n13 OUT+.n12 0.8195
R2777 OUT+.n8 OUT+.t16 0.8195
R2778 OUT+.n8 OUT+.n7 0.8195
R2779 OUT+.n3 OUT+.t24 0.8195
R2780 OUT+.n3 OUT+.n2 0.8195
R2781 OUT+.n100 OUT+.n99 0.730098
R2782 OUT+.n100 OUT+.n94 0.503326
R2783 OUT+.n101 OUT+.n89 0.503326
R2784 OUT+.n102 OUT+.n84 0.503326
R2785 OUT+.n103 OUT+.n79 0.503326
R2786 OUT+.n104 OUT+.n74 0.503326
R2787 OUT+.n105 OUT+.n69 0.503326
R2788 OUT+.n106 OUT+.n64 0.503326
R2789 OUT+.n107 OUT+.n59 0.503326
R2790 OUT+.n108 OUT+.n54 0.503326
R2791 OUT+.n109 OUT+.n49 0.503326
R2792 OUT+.n110 OUT+.n44 0.503326
R2793 OUT+.n111 OUT+.n39 0.503326
R2794 OUT+.n112 OUT+.n34 0.503326
R2795 OUT+.n113 OUT+.n29 0.503326
R2796 OUT+.n114 OUT+.n24 0.503326
R2797 OUT+.n115 OUT+.n19 0.503326
R2798 OUT+.n116 OUT+.n14 0.503326
R2799 OUT+.n117 OUT+.n9 0.503326
R2800 OUT+.n118 OUT+.n4 0.503326
R2801 OUT+ OUT+.n118 0.267665
R2802 OUT+.n101 OUT+.n100 0.227272
R2803 OUT+.n102 OUT+.n101 0.227272
R2804 OUT+.n103 OUT+.n102 0.227272
R2805 OUT+.n104 OUT+.n103 0.227272
R2806 OUT+.n105 OUT+.n104 0.227272
R2807 OUT+.n106 OUT+.n105 0.227272
R2808 OUT+.n107 OUT+.n106 0.227272
R2809 OUT+.n108 OUT+.n107 0.227272
R2810 OUT+.n109 OUT+.n108 0.227272
R2811 OUT+.n110 OUT+.n109 0.227272
R2812 OUT+.n111 OUT+.n110 0.227272
R2813 OUT+.n112 OUT+.n111 0.227272
R2814 OUT+.n113 OUT+.n112 0.227272
R2815 OUT+.n114 OUT+.n113 0.227272
R2816 OUT+.n115 OUT+.n114 0.227272
R2817 OUT+.n116 OUT+.n115 0.227272
R2818 OUT+.n117 OUT+.n116 0.227272
R2819 OUT+.n118 OUT+.n117 0.227272
R2820 B6.n2 B6.t1 48.4147
R2821 B6.n0 B6.t2 19.0247
R2822 B6.n0 B6.t0 17.3935
R2823 B6.n2 B6 10.8029
R2824 B6.n1 B6.n0 4.12942
R2825 B6 B6.n1 2.25699
R2826 B6 B6.n2 0.233179
R2827 B6.n1 B6 0.0067069
R2828 VDD.n411 VDD.t245 490.522
R2829 VDD.n416 VDD.t343 490.522
R2830 VDD.n433 VDD.t248 490.522
R2831 VDD.n428 VDD.t75 490.522
R2832 VDD.n423 VDD.t221 490.522
R2833 VDD.n406 VDD.t34 490.522
R2834 VDD.n411 VDD.t78 485.783
R2835 VDD.n416 VDD.t37 485.783
R2836 VDD.n433 VDD.t341 485.783
R2837 VDD.n428 VDD.t243 485.783
R2838 VDD.n423 VDD.t241 485.783
R2839 VDD.n406 VDD.t140 485.783
R2840 VDD VDD.t127 432.043
R2841 VDD VDD.t312 432.043
R2842 VDD VDD.t207 432.043
R2843 VDD VDD.t44 432.043
R2844 VDD VDD.t122 432.043
R2845 VDD VDD.t125 432.043
R2846 VDD.n78 VDD.t239 166.102
R2847 VDD.n95 VDD.t228 161.018
R2848 VDD.n64 VDD.t209 159.322
R2849 VDD.n80 VDD.t226 155.933
R2850 VDD.n96 VDD.t215 150.847
R2851 VDD.n62 VDD.t210 149.154
R2852 VDD.n82 VDD.t147 145.763
R2853 VDD.n97 VDD.t213 140.679
R2854 VDD.n60 VDD.t112 138.983
R2855 VDD.n3 VDD.t218 135.114
R2856 VDD.n123 VDD.t193 132.868
R2857 VDD.n138 VDD.t166 132.868
R2858 VDD.n272 VDD.t186 132.868
R2859 VDD.n287 VDD.t161 132.868
R2860 VDD.n98 VDD.t231 130.508
R2861 VDD.n75 VDD.t142 118.865
R2862 VDD.n4 VDD.t216 118.644
R2863 VDD.n46 VDD.t227 118.644
R2864 VDD.n73 VDD.t39 111.865
R2865 VDD.n755 VDD.t214 110.169
R2866 VDD.n6 VDD.t238 108.475
R2867 VDD.n44 VDD.t240 108.475
R2868 VDD.n160 VDD.t308 107.992
R2869 VDD.n309 VDD.t299 107.992
R2870 VDD.n214 VDD.t200 102.593
R2871 VDD.n226 VDD.t203 102.593
R2872 VDD.n363 VDD.t294 102.593
R2873 VDD.n375 VDD.t302 102.593
R2874 VDD.n750 VDD.t236 100.001
R2875 VDD.n8 VDD.t273 98.3056
R2876 VDD.n42 VDD.t119 98.3056
R2877 VDD.n51 VDD.t211 98.3056
R2878 VDD.n190 VDD.t150 97.1927
R2879 VDD.n202 VDD.t149 97.1927
R2880 VDD.n339 VDD.t106 97.1927
R2881 VDD.n351 VDD.t300 97.1927
R2882 VDD.n169 VDD.t152 91.7932
R2883 VDD.n181 VDD.t320 91.7932
R2884 VDD.n318 VDD.t139 91.7932
R2885 VDD.n330 VDD.t108 91.7932
R2886 VDD.n123 VDD.t191 90.9096
R2887 VDD.n138 VDD.t163 90.9096
R2888 VDD.n272 VDD.t184 90.9096
R2889 VDD.n287 VDD.t158 90.9096
R2890 VDD.n751 VDD.t117 89.831
R2891 VDD.n11 VDD.t233 88.1361
R2892 VDD.n235 VDD.t281 86.3936
R2893 VDD.n235 VDD.t196 86.3936
R2894 VDD.n169 VDD.t153 80.994
R2895 VDD.n181 VDD.t96 80.994
R2896 VDD.n318 VDD.t301 80.994
R2897 VDD.n330 VDD.t111 80.994
R2898 VDD.n13 VDD.t217 77.9666
R2899 VDD.n28 VDD.t225 77.9666
R2900 VDD.n134 VDD.t181 76.9236
R2901 VDD.n283 VDD.t173 76.9236
R2902 VDD.n190 VDD.t282 75.5945
R2903 VDD.n202 VDD.t280 75.5945
R2904 VDD.n339 VDD.t285 75.5945
R2905 VDD.n351 VDD.t284 75.5945
R2906 VDD.n390 VDD.t304 75.5945
R2907 VDD.n214 VDD.t310 70.1949
R2908 VDD.n226 VDD.t319 70.1949
R2909 VDD.n363 VDD.t335 70.1949
R2910 VDD.n375 VDD.t340 70.1949
R2911 VDD.n15 VDD.t237 67.7971
R2912 VDD.n26 VDD.t224 67.7971
R2913 VDD.n33 VDD.t145 67.7971
R2914 VDD.n148 VDD.t201 64.7953
R2915 VDD.n157 VDD.t317 64.7953
R2916 VDD.n160 VDD.t205 64.7953
R2917 VDD.n297 VDD.t290 64.7953
R2918 VDD.n306 VDD.t297 64.7953
R2919 VDD.n309 VDD.t339 64.7953
R2920 VDD.n386 VDD.t296 62.6355
R2921 VDD.n211 VDD.t154 59.3957
R2922 VDD.n223 VDD.t311 59.3957
R2923 VDD.n360 VDD.t283 59.3957
R2924 VDD.n372 VDD.t286 59.3957
R2925 VDD.n17 VDD.t115 57.6276
R2926 VDD.n24 VDD.t41 57.6276
R2927 VDD.n193 VDD.t95 53.9962
R2928 VDD.n205 VDD.t151 53.9962
R2929 VDD.n342 VDD.t110 53.9962
R2930 VDD.n354 VDD.t107 53.9962
R2931 VDD.n102 VDD.t270 52.5429
R2932 VDD.n166 VDD.t204 48.5966
R2933 VDD.n178 VDD.t97 48.5966
R2934 VDD.n315 VDD.t337 48.5966
R2935 VDD.n327 VDD.t336 48.5966
R2936 VDD.n231 VDD.t314 43.197
R2937 VDD.n240 VDD.t199 43.197
R2938 VDD.n380 VDD.t298 43.197
R2939 VDD.n395 VDD.t307 43.197
R2940 VDD.n502 VDD.t80 42.5052
R2941 VDD.n620 VDD.t54 40.9872
R2942 VDD.n600 VDD.t70 39.4692
R2943 VDD.n600 VDD.t27 37.9512
R2944 VDD.n172 VDD.t315 37.7975
R2945 VDD.n184 VDD.t277 37.7975
R2946 VDD.n321 VDD.t288 37.7975
R2947 VDD.n333 VDD.t293 37.7975
R2948 VDD.n620 VDD.t20 36.4331
R2949 VDD.n128 VDD.t178 34.9655
R2950 VDD.n141 VDD.t156 34.9655
R2951 VDD.n277 VDD.t170 34.9655
R2952 VDD.n290 VDD.t189 34.9655
R2953 VDD.n502 VDD.t89 34.9151
R2954 VDD.n638 VDD.t48 32.6381
R2955 VDD.n187 VDD.t198 32.3979
R2956 VDD.n199 VDD.t278 32.3979
R2957 VDD.n336 VDD.t138 32.3979
R2958 VDD.n348 VDD.t137 32.3979
R2959 VDD.n617 VDD.t64 31.12
R2960 VDD.n597 VDD.t26 29.602
R2961 VDD.n602 VDD.t10 28.084
R2962 VDD.n217 VDD.t309 26.9983
R2963 VDD.n366 VDD.t109 26.9983
R2964 VDD.n623 VDD.t30 26.566
R2965 VDD.n503 VDD.t46 25.0479
R2966 VDD.n635 VDD.t15 22.7709
R2967 VDD.n151 VDD.t202 21.5988
R2968 VDD.n154 VDD.t155 21.5988
R2969 VDD.n163 VDD.t206 21.5988
R2970 VDD.n300 VDD.t291 21.5988
R2971 VDD.n303 VDD.t305 21.5988
R2972 VDD.n312 VDD.t289 21.5988
R2973 VDD.n615 VDD.t5 21.2529
R2974 VDD.n130 VDD.t176 20.9795
R2975 VDD.n279 VDD.t168 20.9795
R2976 VDD.n594 VDD.t61 19.7348
R2977 VDD.n605 VDD.t28 18.2168
R2978 VDD.n625 VDD.t32 16.6988
R2979 VDD.n208 VDD.t276 16.1992
R2980 VDD.n220 VDD.t279 16.1992
R2981 VDD.n357 VDD.t303 16.1992
R2982 VDD.n369 VDD.t287 16.1992
R2983 VDD.n453 VDD.t31 15.9398
R2984 VDD.n131 VDD.n129 14.3187
R2985 VDD.n280 VDD.n278 14.3187
R2986 VDD.n633 VDD.t2 12.9037
R2987 VDD.n612 VDD.t68 11.3857
R2988 VDD.n196 VDD.t275 10.7996
R2989 VDD.n345 VDD.t292 10.7996
R2990 VDD.n719 VDD.t87 10.6267
R2991 VDD.n592 VDD.t98 9.86767
R2992 VDD.n412 VDD.t79 9.56883
R2993 VDD.n417 VDD.t38 9.56883
R2994 VDD.n424 VDD.t242 9.56883
R2995 VDD.n407 VDD.t141 9.56883
R2996 VDD.n413 VDD.n410 9.47246
R2997 VDD.n418 VDD.n415 9.47246
R2998 VDD.n425 VDD.n422 9.47246
R2999 VDD.n430 VDD.n421 9.47246
R3000 VDD.n427 VDD.t244 9.47246
R3001 VDD.n435 VDD.n420 9.47246
R3002 VDD.n432 VDD.t342 9.47246
R3003 VDD.n408 VDD.n405 9.47246
R3004 VDD.n607 VDD.t0 8.34965
R3005 VDD.n23 VDD.n22 8.30127
R3006 VDD.n743 VDD.n742 8.09245
R3007 VDD.n84 VDD.t148 7.67003
R3008 VDD.n628 VDD.t72 6.83162
R3009 VDD.n414 VDD.t128 6.40636
R3010 VDD.n419 VDD.t313 6.40636
R3011 VDD.n426 VDD.t208 6.40636
R3012 VDD.n431 VDD.t45 6.40636
R3013 VDD.n436 VDD.t123 6.40636
R3014 VDD.n409 VDD.t126 6.40636
R3015 VDD.n726 VDD.n725 6.37537
R3016 VDD.n412 VDD.n411 6.3005
R3017 VDD.n417 VDD.n416 6.3005
R3018 VDD.n424 VDD.n423 6.3005
R3019 VDD.n429 VDD.n428 6.3005
R3020 VDD.n434 VDD.n433 6.3005
R3021 VDD.n720 VDD.n719 6.3005
R3022 VDD.n579 VDD.t29 6.3005
R3023 VDD.n590 VDD.t82 6.3005
R3024 VDD.n593 VDD.n592 6.3005
R3025 VDD.n595 VDD.n594 6.3005
R3026 VDD.n598 VDD.n597 6.3005
R3027 VDD.n601 VDD.n600 6.3005
R3028 VDD.n603 VDD.n602 6.3005
R3029 VDD.n606 VDD.n605 6.3005
R3030 VDD.n608 VDD.n607 6.3005
R3031 VDD.n611 VDD.n610 6.3005
R3032 VDD.n613 VDD.n612 6.3005
R3033 VDD.n616 VDD.n615 6.3005
R3034 VDD.n618 VDD.n617 6.3005
R3035 VDD.n621 VDD.n620 6.3005
R3036 VDD.n624 VDD.n623 6.3005
R3037 VDD.n626 VDD.n625 6.3005
R3038 VDD.n629 VDD.n628 6.3005
R3039 VDD.n631 VDD.n630 6.3005
R3040 VDD.n634 VDD.n633 6.3005
R3041 VDD.n636 VDD.n635 6.3005
R3042 VDD.n639 VDD.n638 6.3005
R3043 VDD.n733 VDD.n732 6.3005
R3044 VDD.n521 VDD.n520 6.3005
R3045 VDD.n532 VDD.n531 6.3005
R3046 VDD.n584 VDD.n583 6.3005
R3047 VDD.n457 VDD.n454 6.3005
R3048 VDD.n539 VDD.n502 6.3005
R3049 VDD.n538 VDD.n503 6.3005
R3050 VDD.n407 VDD.n406 6.3005
R3051 VDD.n246 VDD.n245 6.3005
R3052 VDD.n245 VDD.n244 6.3005
R3053 VDD.n385 VDD.n384 6.3005
R3054 VDD.n392 VDD.n391 6.3005
R3055 VDD.n391 VDD.n390 6.3005
R3056 VDD.n103 VDD.n102 6.3005
R3057 VDD.n753 VDD.n750 6.3005
R3058 VDD.n752 VDD.n751 6.3005
R3059 VDD.n89 VDD.n86 6.3005
R3060 VDD.n76 VDD.n73 6.3005
R3061 VDD.n52 VDD.n51 6.3005
R3062 VDD.n34 VDD.n33 6.3005
R3063 VDD.n5 VDD.n4 6.3005
R3064 VDD.n7 VDD.n6 6.3005
R3065 VDD.n9 VDD.n8 6.3005
R3066 VDD.n12 VDD.n11 6.3005
R3067 VDD.n14 VDD.n13 6.3005
R3068 VDD.n16 VDD.n15 6.3005
R3069 VDD.n18 VDD.n17 6.3005
R3070 VDD.n21 VDD.n20 6.3005
R3071 VDD.n25 VDD.n24 6.3005
R3072 VDD.n27 VDD.n26 6.3005
R3073 VDD.n29 VDD.n28 6.3005
R3074 VDD.n43 VDD.n42 6.3005
R3075 VDD.n45 VDD.n44 6.3005
R3076 VDD.n47 VDD.n46 6.3005
R3077 VDD.n61 VDD.n60 6.3005
R3078 VDD.n63 VDD.n62 6.3005
R3079 VDD.n65 VDD.n64 6.3005
R3080 VDD.n79 VDD.n78 6.3005
R3081 VDD.n81 VDD.n80 6.3005
R3082 VDD.n83 VDD.n82 6.3005
R3083 VDD.n767 VDD.n95 6.3005
R3084 VDD.n766 VDD.n96 6.3005
R3085 VDD.n765 VDD.n97 6.3005
R3086 VDD.n764 VDD.n98 6.3005
R3087 VDD.n752 VDD.t118 6.18063
R3088 VDD.n574 VDD.n489 6.13519
R3089 VDD.n671 VDD.n670 6.12312
R3090 VDD.n653 VDD.t321 6.12266
R3091 VDD.n714 VDD.t88 6.11709
R3092 VDD.n3 VDD.n2 6.10984
R3093 VDD.n768 VDD.n94 6.09557
R3094 VDD.n19 VDD.t116 6.09557
R3095 VDD.n175 VDD.t316 5.40007
R3096 VDD.n324 VDD.t295 5.40007
R3097 VDD.n250 VDD.n249 5.35463
R3098 VDD.n522 VDD.t17 5.31359
R3099 VDD.n72 VDD.n71 4.98502
R3100 VDD.n717 VDD.n716 4.86789
R3101 VDD.n249 VDD.t197 4.69594
R3102 VDD.n573 VDD.n568 4.68801
R3103 VDD.n579 VDD.n578 4.5005
R3104 VDD.n722 VDD.n721 4.5005
R3105 VDD.n457 VDD.n456 4.5005
R3106 VDD.n519 VDD.n518 4.5005
R3107 VDD.n518 VDD.n517 4.5005
R3108 VDD.n530 VDD.n529 4.5005
R3109 VDD.n529 VDD.n528 4.5005
R3110 VDD.n512 VDD.n511 4.5005
R3111 VDD.n511 VDD.n510 4.5005
R3112 VDD.n739 VDD.n738 4.5005
R3113 VDD.n738 VDD.n737 4.5005
R3114 VDD.n388 VDD.n387 4.5005
R3115 VDD.n387 VDD.n386 4.5005
R3116 VDD.n89 VDD.n88 4.5005
R3117 VDD.n52 VDD.n50 4.5005
R3118 VDD.n34 VDD.n32 4.5005
R3119 VDD.n103 VDD.n101 4.5005
R3120 VDD.n59 VDD.n58 4.26092
R3121 VDD.n41 VDD.n40 4.24066
R3122 VDD.n726 VDD.n718 4.2252
R3123 VDD.n507 VDD.t22 4.17507
R3124 VDD.n144 VDD.t157 4.00385
R3125 VDD.n293 VDD.t190 4.00385
R3126 VDD.n122 VDD.n120 3.98789
R3127 VDD.n271 VDD.n269 3.98789
R3128 VDD.n737 VDD.t101 3.79557
R3129 VDD.n756 VDD.n755 3.70875
R3130 VDD.n748 VDD.n747 3.62297
R3131 VDD.n58 VDD.n57 3.2271
R3132 VDD.n40 VDD.n39 3.20234
R3133 VDD.n744 VDD.n743 3.19795
R3134 VDD.n71 VDD.n70 3.17695
R3135 VDD.n746 VDD.n745 3.16881
R3136 VDD.n122 VDD.n121 3.16646
R3137 VDD.n271 VDD.n270 3.16646
R3138 VDD.n748 VDD.n404 3.15399
R3139 VDD.n649 VDD.n460 3.15224
R3140 VDD.n643 VDD.n464 3.15224
R3141 VDD.n637 VDD.n468 3.15224
R3142 VDD.n627 VDD.n472 3.15224
R3143 VDD.n619 VDD.n476 3.15224
R3144 VDD.n609 VDD.n480 3.15224
R3145 VDD.n599 VDD.n484 3.15224
R3146 VDD.n591 VDD.n488 3.15224
R3147 VDD.n588 VDD.n587 3.15175
R3148 VDD.n677 VDD.n676 3.15175
R3149 VDD.n54 VDD.n53 3.15175
R3150 VDD.n92 VDD.n91 3.15175
R3151 VDD.n458 VDD.n451 3.15175
R3152 VDD.n36 VDD.n35 3.15175
R3153 VDD.n69 VDD.n68 3.15175
R3154 VDD.n759 VDD.n105 3.15175
R3155 VDD.n587 VDD.n586 3.151
R3156 VDD.n728 VDD.n458 3.151
R3157 VDD.n91 VDD.n90 3.151
R3158 VDD.n105 VDD.n104 3.151
R3159 VDD.n37 VDD.n36 3.151
R3160 VDD.n451 VDD.n450 3.151
R3161 VDD.n68 VDD.n67 3.151
R3162 VDD.n55 VDD.n54 3.151
R3163 VDD.n513 VDD.n509 3.1505
R3164 VDD.n509 VDD.n508 3.1505
R3165 VDD.n534 VDD.n533 3.1505
R3166 VDD.n535 VDD.n534 3.1505
R3167 VDD.n523 VDD.n522 3.1505
R3168 VDD.n524 VDD.n523 3.1505
R3169 VDD.n736 VDD.n735 3.1505
R3170 VDD.n735 VDD.n734 3.1505
R3171 VDD.n143 VDD.n142 3.1505
R3172 VDD.n142 VDD.n141 3.1505
R3173 VDD.n125 VDD.n124 3.1505
R3174 VDD.n124 VDD.n123 3.1505
R3175 VDD.n129 VDD.n127 3.1505
R3176 VDD.n129 VDD.n128 3.1505
R3177 VDD.n132 VDD.n131 3.1505
R3178 VDD.n131 VDD.n130 3.1505
R3179 VDD.n136 VDD.n135 3.1505
R3180 VDD.n135 VDD.n134 3.1505
R3181 VDD.n140 VDD.n139 3.1505
R3182 VDD.n139 VDD.n138 3.1505
R3183 VDD.n147 VDD.n146 3.1505
R3184 VDD.n146 VDD.n145 3.1505
R3185 VDD.n150 VDD.n149 3.1505
R3186 VDD.n149 VDD.n148 3.1505
R3187 VDD.n153 VDD.n152 3.1505
R3188 VDD.n152 VDD.n151 3.1505
R3189 VDD.n156 VDD.n155 3.1505
R3190 VDD.n155 VDD.n154 3.1505
R3191 VDD.n159 VDD.n158 3.1505
R3192 VDD.n158 VDD.n157 3.1505
R3193 VDD.n162 VDD.n161 3.1505
R3194 VDD.n161 VDD.n160 3.1505
R3195 VDD.n165 VDD.n164 3.1505
R3196 VDD.n164 VDD.n163 3.1505
R3197 VDD.n168 VDD.n167 3.1505
R3198 VDD.n167 VDD.n166 3.1505
R3199 VDD.n171 VDD.n170 3.1505
R3200 VDD.n170 VDD.n169 3.1505
R3201 VDD.n174 VDD.n173 3.1505
R3202 VDD.n173 VDD.n172 3.1505
R3203 VDD.n177 VDD.n176 3.1505
R3204 VDD.n176 VDD.n175 3.1505
R3205 VDD.n180 VDD.n179 3.1505
R3206 VDD.n179 VDD.n178 3.1505
R3207 VDD.n183 VDD.n182 3.1505
R3208 VDD.n182 VDD.n181 3.1505
R3209 VDD.n186 VDD.n185 3.1505
R3210 VDD.n185 VDD.n184 3.1505
R3211 VDD.n189 VDD.n188 3.1505
R3212 VDD.n188 VDD.n187 3.1505
R3213 VDD.n192 VDD.n191 3.1505
R3214 VDD.n191 VDD.n190 3.1505
R3215 VDD.n195 VDD.n194 3.1505
R3216 VDD.n194 VDD.n193 3.1505
R3217 VDD.n198 VDD.n197 3.1505
R3218 VDD.n197 VDD.n196 3.1505
R3219 VDD.n201 VDD.n200 3.1505
R3220 VDD.n200 VDD.n199 3.1505
R3221 VDD.n204 VDD.n203 3.1505
R3222 VDD.n203 VDD.n202 3.1505
R3223 VDD.n207 VDD.n206 3.1505
R3224 VDD.n206 VDD.n205 3.1505
R3225 VDD.n210 VDD.n209 3.1505
R3226 VDD.n209 VDD.n208 3.1505
R3227 VDD.n213 VDD.n212 3.1505
R3228 VDD.n212 VDD.n211 3.1505
R3229 VDD.n216 VDD.n215 3.1505
R3230 VDD.n215 VDD.n214 3.1505
R3231 VDD.n219 VDD.n218 3.1505
R3232 VDD.n218 VDD.n217 3.1505
R3233 VDD.n222 VDD.n221 3.1505
R3234 VDD.n221 VDD.n220 3.1505
R3235 VDD.n225 VDD.n224 3.1505
R3236 VDD.n224 VDD.n223 3.1505
R3237 VDD.n228 VDD.n227 3.1505
R3238 VDD.n227 VDD.n226 3.1505
R3239 VDD.n230 VDD.n229 3.1505
R3240 VDD.n229 VDD.t318 3.1505
R3241 VDD.n233 VDD.n232 3.1505
R3242 VDD.n232 VDD.n231 3.1505
R3243 VDD.n237 VDD.n236 3.1505
R3244 VDD.n236 VDD.n235 3.1505
R3245 VDD.n292 VDD.n291 3.1505
R3246 VDD.n291 VDD.n290 3.1505
R3247 VDD.n274 VDD.n273 3.1505
R3248 VDD.n273 VDD.n272 3.1505
R3249 VDD.n278 VDD.n276 3.1505
R3250 VDD.n278 VDD.n277 3.1505
R3251 VDD.n281 VDD.n280 3.1505
R3252 VDD.n280 VDD.n279 3.1505
R3253 VDD.n285 VDD.n284 3.1505
R3254 VDD.n284 VDD.n283 3.1505
R3255 VDD.n289 VDD.n288 3.1505
R3256 VDD.n288 VDD.n287 3.1505
R3257 VDD.n296 VDD.n295 3.1505
R3258 VDD.n295 VDD.n294 3.1505
R3259 VDD.n299 VDD.n298 3.1505
R3260 VDD.n298 VDD.n297 3.1505
R3261 VDD.n302 VDD.n301 3.1505
R3262 VDD.n301 VDD.n300 3.1505
R3263 VDD.n305 VDD.n304 3.1505
R3264 VDD.n304 VDD.n303 3.1505
R3265 VDD.n308 VDD.n307 3.1505
R3266 VDD.n307 VDD.n306 3.1505
R3267 VDD.n311 VDD.n310 3.1505
R3268 VDD.n310 VDD.n309 3.1505
R3269 VDD.n314 VDD.n313 3.1505
R3270 VDD.n313 VDD.n312 3.1505
R3271 VDD.n317 VDD.n316 3.1505
R3272 VDD.n316 VDD.n315 3.1505
R3273 VDD.n320 VDD.n319 3.1505
R3274 VDD.n319 VDD.n318 3.1505
R3275 VDD.n323 VDD.n322 3.1505
R3276 VDD.n322 VDD.n321 3.1505
R3277 VDD.n326 VDD.n325 3.1505
R3278 VDD.n325 VDD.n324 3.1505
R3279 VDD.n329 VDD.n328 3.1505
R3280 VDD.n328 VDD.n327 3.1505
R3281 VDD.n332 VDD.n331 3.1505
R3282 VDD.n331 VDD.n330 3.1505
R3283 VDD.n335 VDD.n334 3.1505
R3284 VDD.n334 VDD.n333 3.1505
R3285 VDD.n338 VDD.n337 3.1505
R3286 VDD.n337 VDD.n336 3.1505
R3287 VDD.n341 VDD.n340 3.1505
R3288 VDD.n340 VDD.n339 3.1505
R3289 VDD.n344 VDD.n343 3.1505
R3290 VDD.n343 VDD.n342 3.1505
R3291 VDD.n347 VDD.n346 3.1505
R3292 VDD.n346 VDD.n345 3.1505
R3293 VDD.n350 VDD.n349 3.1505
R3294 VDD.n349 VDD.n348 3.1505
R3295 VDD.n353 VDD.n352 3.1505
R3296 VDD.n352 VDD.n351 3.1505
R3297 VDD.n356 VDD.n355 3.1505
R3298 VDD.n355 VDD.n354 3.1505
R3299 VDD.n359 VDD.n358 3.1505
R3300 VDD.n358 VDD.n357 3.1505
R3301 VDD.n362 VDD.n361 3.1505
R3302 VDD.n361 VDD.n360 3.1505
R3303 VDD.n365 VDD.n364 3.1505
R3304 VDD.n364 VDD.n363 3.1505
R3305 VDD.n368 VDD.n367 3.1505
R3306 VDD.n367 VDD.n366 3.1505
R3307 VDD.n371 VDD.n370 3.1505
R3308 VDD.n370 VDD.n369 3.1505
R3309 VDD.n374 VDD.n373 3.1505
R3310 VDD.n373 VDD.n372 3.1505
R3311 VDD.n377 VDD.n376 3.1505
R3312 VDD.n376 VDD.n375 3.1505
R3313 VDD.n379 VDD.n378 3.1505
R3314 VDD.n378 VDD.t338 3.1505
R3315 VDD.n382 VDD.n381 3.1505
R3316 VDD.n381 VDD.n380 3.1505
R3317 VDD.n596 VDD.n486 3.08376
R3318 VDD.n604 VDD.n482 3.08376
R3319 VDD.n614 VDD.n478 3.08376
R3320 VDD.n622 VDD.n474 3.08376
R3321 VDD.n632 VDD.n470 3.08376
R3322 VDD.n640 VDD.n466 3.08376
R3323 VDD.n646 VDD.n462 3.08376
R3324 VDD.n682 VDD.n669 3.08376
R3325 VDD.n686 VDD.n667 3.08376
R3326 VDD.n691 VDD.n665 3.08376
R3327 VDD.n695 VDD.n663 3.08376
R3328 VDD.n700 VDD.n661 3.08376
R3329 VDD.n704 VDD.n659 3.08376
R3330 VDD.n709 VDD.n657 3.08376
R3331 VDD.n137 VDD.n115 3.07789
R3332 VDD.n133 VDD.n117 3.07789
R3333 VDD.n126 VDD.n119 3.07789
R3334 VDD.n286 VDD.n264 3.07789
R3335 VDD.n282 VDD.n266 3.07789
R3336 VDD.n275 VDD.n268 3.07789
R3337 VDD.n762 VDD.n100 3.06224
R3338 VDD.n10 VDD.n1 3.06224
R3339 VDD.n730 VDD.n447 3.05441
R3340 VDD.n537 VDD.n505 3.05441
R3341 VDD.n541 VDD.n501 3.05441
R3342 VDD.n546 VDD.n499 3.05441
R3343 VDD.n550 VDD.n497 3.05441
R3344 VDD.n555 VDD.n495 3.05441
R3345 VDD.n560 VDD.n493 3.05441
R3346 VDD.n564 VDD.n491 3.05441
R3347 VDD.n630 VDD.t8 3.03655
R3348 VDD.n486 VDD.t266 3.03383
R3349 VDD.n486 VDD.n485 3.03383
R3350 VDD.n482 VDD.t265 3.03383
R3351 VDD.n482 VDD.n481 3.03383
R3352 VDD.n478 VDD.t69 3.03383
R3353 VDD.n478 VDD.n477 3.03383
R3354 VDD.n474 VDD.t21 3.03383
R3355 VDD.n474 VDD.n473 3.03383
R3356 VDD.n470 VDD.t25 3.03383
R3357 VDD.n470 VDD.n469 3.03383
R3358 VDD.n466 VDD.t103 3.03383
R3359 VDD.n466 VDD.n465 3.03383
R3360 VDD.n462 VDD.t327 3.03383
R3361 VDD.n462 VDD.n461 3.03383
R3362 VDD.n460 VDD.t253 3.03383
R3363 VDD.n460 VDD.n459 3.03383
R3364 VDD.n464 VDD.t47 3.03383
R3365 VDD.n464 VDD.n463 3.03383
R3366 VDD.n468 VDD.t16 3.03383
R3367 VDD.n468 VDD.n467 3.03383
R3368 VDD.n472 VDD.t33 3.03383
R3369 VDD.n472 VDD.n471 3.03383
R3370 VDD.n476 VDD.t94 3.03383
R3371 VDD.n476 VDD.n475 3.03383
R3372 VDD.n480 VDD.t1 3.03383
R3373 VDD.n480 VDD.n479 3.03383
R3374 VDD.n484 VDD.t86 3.03383
R3375 VDD.n484 VDD.n483 3.03383
R3376 VDD.n488 VDD.t83 3.03383
R3377 VDD.n488 VDD.n487 3.03383
R3378 VDD.n669 VDD.t62 3.03383
R3379 VDD.n669 VDD.n668 3.03383
R3380 VDD.n667 VDD.t11 3.03383
R3381 VDD.n667 VDD.n666 3.03383
R3382 VDD.n665 VDD.t256 3.03383
R3383 VDD.n665 VDD.n664 3.03383
R3384 VDD.n663 VDD.t51 3.03383
R3385 VDD.n663 VDD.n662 3.03383
R3386 VDD.n661 VDD.t9 3.03383
R3387 VDD.n661 VDD.n660 3.03383
R3388 VDD.n659 VDD.t81 3.03383
R3389 VDD.n659 VDD.n658 3.03383
R3390 VDD.n657 VDD.t18 3.03383
R3391 VDD.n657 VDD.n656 3.03383
R3392 VDD.n447 VDD.t102 3.03383
R3393 VDD.n447 VDD.n446 3.03383
R3394 VDD.n505 VDD.t332 3.03383
R3395 VDD.n505 VDD.n504 3.03383
R3396 VDD.n501 VDD.t19 3.03383
R3397 VDD.n501 VDD.n500 3.03383
R3398 VDD.n499 VDD.t63 3.03383
R3399 VDD.n499 VDD.n498 3.03383
R3400 VDD.n497 VDD.t65 3.03383
R3401 VDD.n497 VDD.n496 3.03383
R3402 VDD.n495 VDD.t269 3.03383
R3403 VDD.n495 VDD.n494 3.03383
R3404 VDD.n493 VDD.t71 3.03383
R3405 VDD.n493 VDD.n492 3.03383
R3406 VDD.n491 VDD.t322 3.03383
R3407 VDD.n491 VDD.n490 3.03383
R3408 VDD.n100 VDD.t232 3.03383
R3409 VDD.n100 VDD.n99 3.03383
R3410 VDD.n1 VDD.t274 3.03383
R3411 VDD.n1 VDD.n0 3.03383
R3412 VDD.n71 VDD.t40 2.69573
R3413 VDD.n40 VDD.t146 2.66058
R3414 VDD.n744 VDD.n419 2.63002
R3415 VDD.n745 VDD.n414 2.62915
R3416 VDD.n242 VDD.n241 2.6255
R3417 VDD.n241 VDD.n240 2.6255
R3418 VDD.n401 VDD.n400 2.6255
R3419 VDD.n400 VDD.t306 2.6255
R3420 VDD.n397 VDD.n396 2.6255
R3421 VDD.n396 VDD.n395 2.6255
R3422 VDD.n58 VDD.t212 2.62483
R3423 VDD.n77 VDD.n76 2.62147
R3424 VDD.n404 VDD.n254 2.61247
R3425 VDD.n573 VDD.n572 2.46941
R3426 VDD.n749 VDD.n748 2.31907
R3427 VDD.n454 VDD.n453 2.27754
R3428 VDD.n456 VDD.n455 2.27754
R3429 VDD.n254 VDD.n253 2.25578
R3430 VDD.n718 VDD.n655 2.25504
R3431 VDD.n403 VDD.n402 2.25132
R3432 VDD.n574 VDD.n573 2.2505
R3433 VDD.n742 VDD.n741 2.2505
R3434 VDD.n113 VDD.n112 2.2505
R3435 VDD.n586 VDD.n585 2.1005
R3436 VDD.n34 VDD.n31 1.88512
R3437 VDD.n76 VDD.n74 1.83127
R3438 VDD.n89 VDD.n87 1.77742
R3439 VDD.n725 VDD.n724 1.7738
R3440 VDD.n585 VDD.n584 1.62266
R3441 VDD.n387 VDD.n385 1.5755
R3442 VDD.n52 VDD.n49 1.56204
R3443 VDD.n610 VDD.t124 1.51853
R3444 VDD.n741 VDD.n740 1.49894
R3445 VDD.n754 VDD.n749 1.49872
R3446 VDD.n579 VDD.n576 1.463
R3447 VDD.n404 VDD.n403 1.44464
R3448 VDD.n449 VDD.n448 1.3505
R3449 VDD.n675 VDD.n674 1.313
R3450 VDD.n723 VDD.n722 1.24541
R3451 VDD.n457 VDD.n452 1.2005
R3452 VDD.n747 VDD 1.19267
R3453 VDD.n458 VDD.n457 1.19071
R3454 VDD.n747 VDD.n746 1.17203
R3455 VDD.n586 VDD.n580 1.13902
R3456 VDD.n54 VDD.n52 1.12174
R3457 VDD.n722 VDD.n720 1.09451
R3458 VDD.n676 VDD.n675 0.985261
R3459 VDD.n450 VDD.n449 0.916649
R3460 VDD.n253 VDD.n250 0.912795
R3461 VDD.n745 VDD.n744 0.911065
R3462 VDD.n115 VDD.t167 0.9105
R3463 VDD.n115 VDD.n114 0.9105
R3464 VDD.n117 VDD.t177 0.9105
R3465 VDD.n117 VDD.n116 0.9105
R3466 VDD.n119 VDD.t192 0.9105
R3467 VDD.n119 VDD.n118 0.9105
R3468 VDD.n264 VDD.t162 0.9105
R3469 VDD.n264 VDD.n263 0.9105
R3470 VDD.n266 VDD.t169 0.9105
R3471 VDD.n266 VDD.n265 0.9105
R3472 VDD.n268 VDD.t185 0.9105
R3473 VDD.n268 VDD.n267 0.9105
R3474 VDD.n402 VDD.n401 0.903728
R3475 VDD.n523 VDD.n521 0.792716
R3476 VDD.n578 VDD.n577 0.759513
R3477 VDD.n528 VDD.t12 0.759513
R3478 VDD.n534 VDD.n532 0.754991
R3479 VDD.n587 VDD.n579 0.747944
R3480 VDD.n432 VDD.n431 0.742062
R3481 VDD.n427 VDD.n426 0.727335
R3482 VDD.n91 VDD.n89 0.724621
R3483 VDD.n105 VDD.n103 0.59316
R3484 VDD.n582 VDD.n581 0.587761
R3485 VDD.n735 VDD.n733 0.528644
R3486 VDD.n36 VDD.n34 0.525399
R3487 VDD VDD.n413 0.510235
R3488 VDD VDD.n418 0.510235
R3489 VDD VDD.n425 0.510235
R3490 VDD VDD.n430 0.510235
R3491 VDD VDD.n435 0.510235
R3492 VDD VDD.n408 0.510235
R3493 VDD.n743 VDD.n436 0.429578
R3494 VDD.n76 VDD.n75 0.415309
R3495 VDD.n746 VDD.n409 0.394447
R3496 VDD.t29 VDD.n575 0.380007
R3497 VDD.n508 VDD.n507 0.380007
R3498 VDD.n249 VDD.n248 0.247932
R3499 VDD.n168 VDD.n165 0.144117
R3500 VDD.n189 VDD.n186 0.144117
R3501 VDD.n210 VDD.n207 0.144117
R3502 VDD.n230 VDD.n228 0.144117
R3503 VDD.n317 VDD.n314 0.144117
R3504 VDD.n338 VDD.n335 0.144117
R3505 VDD.n359 VDD.n356 0.144117
R3506 VDD.n379 VDD.n377 0.144117
R3507 VDD.n742 VDD.n437 0.137788
R3508 VDD.n254 VDD.n113 0.135259
R3509 VDD.n143 VDD.n140 0.12816
R3510 VDD.n150 VDD.n147 0.12816
R3511 VDD.n153 VDD.n150 0.12816
R3512 VDD.n156 VDD.n153 0.12816
R3513 VDD.n159 VDD.n156 0.12816
R3514 VDD.n162 VDD.n159 0.12816
R3515 VDD.n165 VDD.n162 0.12816
R3516 VDD.n171 VDD.n168 0.12816
R3517 VDD.n174 VDD.n171 0.12816
R3518 VDD.n177 VDD.n174 0.12816
R3519 VDD.n180 VDD.n177 0.12816
R3520 VDD.n183 VDD.n180 0.12816
R3521 VDD.n186 VDD.n183 0.12816
R3522 VDD.n192 VDD.n189 0.12816
R3523 VDD.n195 VDD.n192 0.12816
R3524 VDD.n198 VDD.n195 0.12816
R3525 VDD.n201 VDD.n198 0.12816
R3526 VDD.n204 VDD.n201 0.12816
R3527 VDD.n207 VDD.n204 0.12816
R3528 VDD.n213 VDD.n210 0.12816
R3529 VDD.n216 VDD.n213 0.12816
R3530 VDD.n219 VDD.n216 0.12816
R3531 VDD.n222 VDD.n219 0.12816
R3532 VDD.n225 VDD.n222 0.12816
R3533 VDD.n228 VDD.n225 0.12816
R3534 VDD.n233 VDD.n230 0.12816
R3535 VDD.n292 VDD.n289 0.12816
R3536 VDD.n299 VDD.n296 0.12816
R3537 VDD.n302 VDD.n299 0.12816
R3538 VDD.n305 VDD.n302 0.12816
R3539 VDD.n308 VDD.n305 0.12816
R3540 VDD.n311 VDD.n308 0.12816
R3541 VDD.n314 VDD.n311 0.12816
R3542 VDD.n320 VDD.n317 0.12816
R3543 VDD.n323 VDD.n320 0.12816
R3544 VDD.n326 VDD.n323 0.12816
R3545 VDD.n329 VDD.n326 0.12816
R3546 VDD.n332 VDD.n329 0.12816
R3547 VDD.n335 VDD.n332 0.12816
R3548 VDD.n341 VDD.n338 0.12816
R3549 VDD.n344 VDD.n341 0.12816
R3550 VDD.n347 VDD.n344 0.12816
R3551 VDD.n350 VDD.n347 0.12816
R3552 VDD.n353 VDD.n350 0.12816
R3553 VDD.n356 VDD.n353 0.12816
R3554 VDD.n362 VDD.n359 0.12816
R3555 VDD.n365 VDD.n362 0.12816
R3556 VDD.n368 VDD.n365 0.12816
R3557 VDD.n371 VDD.n368 0.12816
R3558 VDD.n374 VDD.n371 0.12816
R3559 VDD.n377 VDD.n374 0.12816
R3560 VDD.n382 VDD.n379 0.12816
R3561 VDD.n147 VDD.n144 0.122257
R3562 VDD.n296 VDD.n293 0.122257
R3563 VDD.n403 VDD.n255 0.119602
R3564 VDD.n137 VDD.n136 0.118585
R3565 VDD.n286 VDD.n285 0.118585
R3566 VDD.n111 VDD.n110 0.118414
R3567 VDD.n5 VDD.n3 0.115744
R3568 VDD.n7 VDD.n5 0.115744
R3569 VDD.n9 VDD.n7 0.115744
R3570 VDD.n14 VDD.n12 0.115744
R3571 VDD.n16 VDD.n14 0.115744
R3572 VDD.n18 VDD.n16 0.115744
R3573 VDD.n27 VDD.n25 0.115744
R3574 VDD.n29 VDD.n27 0.115744
R3575 VDD.n45 VDD.n43 0.115744
R3576 VDD.n47 VDD.n45 0.115744
R3577 VDD.n63 VDD.n61 0.115744
R3578 VDD.n65 VDD.n63 0.115744
R3579 VDD.n81 VDD.n79 0.115744
R3580 VDD.n83 VDD.n81 0.115744
R3581 VDD.n767 VDD.n766 0.115744
R3582 VDD.n766 VDD.n765 0.115744
R3583 VDD.n765 VDD.n764 0.115744
R3584 VDD.n753 VDD.n752 0.115744
R3585 VDD.n585 VDD.n582 0.113674
R3586 VDD.n724 VDD.n723 0.113071
R3587 VDD.n125 VDD.n122 0.112202
R3588 VDD.n274 VDD.n271 0.112202
R3589 VDD.n30 VDD.n29 0.109159
R3590 VDD.n754 VDD.n753 0.108104
R3591 VDD.n595 VDD.n593 0.107201
R3592 VDD.n603 VDD.n601 0.107201
R3593 VDD.n608 VDD.n606 0.107201
R3594 VDD.n613 VDD.n611 0.107201
R3595 VDD.n618 VDD.n616 0.107201
R3596 VDD.n626 VDD.n624 0.107201
R3597 VDD.n631 VDD.n629 0.107201
R3598 VDD.n636 VDD.n634 0.107201
R3599 VDD.n642 VDD.n641 0.107201
R3600 VDD.n645 VDD.n644 0.107201
R3601 VDD.n648 VDD.n647 0.107201
R3602 VDD.n680 VDD.n679 0.107201
R3603 VDD.n681 VDD.n680 0.107201
R3604 VDD.n684 VDD.n683 0.107201
R3605 VDD.n685 VDD.n684 0.107201
R3606 VDD.n688 VDD.n687 0.107201
R3607 VDD.n689 VDD.n688 0.107201
R3608 VDD.n690 VDD.n689 0.107201
R3609 VDD.n693 VDD.n692 0.107201
R3610 VDD.n694 VDD.n693 0.107201
R3611 VDD.n697 VDD.n696 0.107201
R3612 VDD.n698 VDD.n697 0.107201
R3613 VDD.n699 VDD.n698 0.107201
R3614 VDD.n702 VDD.n701 0.107201
R3615 VDD.n703 VDD.n702 0.107201
R3616 VDD.n706 VDD.n705 0.107201
R3617 VDD.n707 VDD.n706 0.107201
R3618 VDD.n708 VDD.n707 0.107201
R3619 VDD.n711 VDD.n710 0.107201
R3620 VDD.n712 VDD.n711 0.107201
R3621 VDD.n79 VDD.n77 0.106804
R3622 VDD.n599 VDD.n598 0.106273
R3623 VDD.n48 VDD.n47 0.105866
R3624 VDD.n108 VDD.n107 0.104678
R3625 VDD.n253 VDD.n252 0.104412
R3626 VDD.n640 VDD.n639 0.102562
R3627 VDD.n704 VDD.n703 0.102562
R3628 VDD.n563 VDD.n562 0.0995431
R3629 VDD.n562 VDD.n561 0.0995431
R3630 VDD.n559 VDD.n558 0.0995431
R3631 VDD.n558 VDD.n557 0.0995431
R3632 VDD.n557 VDD.n556 0.0995431
R3633 VDD.n554 VDD.n553 0.0995431
R3634 VDD.n553 VDD.n552 0.0995431
R3635 VDD.n552 VDD.n551 0.0995431
R3636 VDD.n549 VDD.n548 0.0995431
R3637 VDD.n548 VDD.n547 0.0995431
R3638 VDD.n545 VDD.n544 0.0995431
R3639 VDD.n544 VDD.n543 0.0995431
R3640 VDD.n543 VDD.n542 0.0995431
R3641 VDD.n539 VDD.n538 0.0995431
R3642 VDD.n561 VDD.n560 0.0986818
R3643 VDD.n621 VDD.n619 0.0979227
R3644 VDD.n66 VDD.n65 0.0970854
R3645 VDD.n429 VDD.n427 0.0968717
R3646 VDD.n434 VDD.n432 0.0968717
R3647 VDD VDD.n768 0.0959878
R3648 VDD.n61 VDD.n59 0.0957073
R3649 VDD.n84 VDD.n83 0.0953491
R3650 VDD.n590 VDD.n589 0.0951392
R3651 VDD.n679 VDD.n678 0.0946753
R3652 VDD.n443 VDD.n442 0.0935509
R3653 VDD.n126 VDD.n125 0.0930532
R3654 VDD.n275 VDD.n274 0.0930532
R3655 VDD.n622 VDD.n621 0.0923557
R3656 VDD.n695 VDD.n694 0.0923557
R3657 VDD.n540 VDD 0.0917919
R3658 VDD.n43 VDD.n41 0.0913202
R3659 VDD.n550 VDD.n549 0.0909306
R3660 VDD.n258 VDD.n257 0.0894222
R3661 VDD.n10 VDD.n9 0.0883049
R3662 VDD.n639 VDD.n637 0.0877165
R3663 VDD.n136 VDD.n133 0.0866702
R3664 VDD.n285 VDD.n282 0.0866702
R3665 VDD.n413 VDD 0.0857212
R3666 VDD.n418 VDD 0.0857212
R3667 VDD.n425 VDD 0.0857212
R3668 VDD.n430 VDD 0.0857212
R3669 VDD.n435 VDD 0.0857212
R3670 VDD.n408 VDD 0.0857212
R3671 VDD.n764 VDD.n763 0.085561
R3672 VDD.n598 VDD.n596 0.0840052
R3673 VDD.n683 VDD.n682 0.0840052
R3674 VDD.n440 VDD.n439 0.0828729
R3675 VDD.n604 VDD.n603 0.0821495
R3676 VDD.n686 VDD.n685 0.0821495
R3677 VDD.n541 VDD.n540 0.0814569
R3678 VDD.n566 VDD.n565 0.0810263
R3679 VDD.n25 VDD.n23 0.0789756
R3680 VDD.n643 VDD.n642 0.0784381
R3681 VDD.n713 VDD.n712 0.0784381
R3682 VDD.n654 VDD.n653 0.0765825
R3683 VDD.n19 VDD.n18 0.0751341
R3684 VDD.n616 VDD.n614 0.073799
R3685 VDD.n692 VDD.n691 0.073799
R3686 VDD.n538 VDD.n537 0.0728445
R3687 VDD.n23 VDD.n21 0.0723902
R3688 VDD.n393 VDD.n392 0.07175
R3689 VDD.n383 VDD.n382 0.0706323
R3690 VDD.n238 VDD.n237 0.0698048
R3691 VDD.n246 VDD.n243 0.0698048
R3692 VDD.n132 VDD 0.0694362
R3693 VDD.n281 VDD 0.0694362
R3694 VDD.n758 VDD.n757 0.0690976
R3695 VDD.n627 VDD.n626 0.068232
R3696 VDD.n650 VDD.n649 0.0673041
R3697 VDD.n730 VDD.n729 0.0650933
R3698 VDD.n634 VDD.n632 0.0635928
R3699 VDD.n701 VDD.n700 0.0635928
R3700 VDD.n547 VDD.n546 0.0633708
R3701 VDD.n262 VDD.n261 0.0619371
R3702 VDD.n399 VDD.n398 0.0615714
R3703 VDD.n593 VDD.n591 0.0598814
R3704 VDD.n414 VDD 0.0594381
R3705 VDD.n419 VDD 0.0594381
R3706 VDD.n426 VDD 0.0594381
R3707 VDD.n431 VDD 0.0594381
R3708 VDD.n436 VDD 0.0594381
R3709 VDD.n409 VDD 0.0594381
R3710 VDD.n127 VDD 0.0592234
R3711 VDD.n276 VDD 0.0592234
R3712 VDD.n609 VDD.n608 0.0580258
R3713 VDD.n564 VDD.n563 0.0556196
R3714 VDD.n646 VDD.n645 0.0543144
R3715 VDD.n709 VDD.n708 0.0543144
R3716 VDD.n556 VDD.n555 0.0538971
R3717 VDD.n647 VDD.n646 0.0533866
R3718 VDD.n710 VDD.n709 0.0533866
R3719 VDD.n515 VDD.n514 0.0521746
R3720 VDD.n144 VDD.n143 0.0515638
R3721 VDD.n293 VDD.n292 0.0515638
R3722 VDD.n234 VDD.n233 0.0509733
R3723 VDD.n611 VDD.n609 0.0496753
R3724 VDD.n237 VDD.n234 0.0491096
R3725 VDD.n591 VDD.n590 0.0478196
R3726 VDD.n555 VDD.n554 0.0461459
R3727 VDD.n565 VDD.n564 0.0444234
R3728 VDD.n632 VDD.n631 0.0441082
R3729 VDD.n700 VDD.n699 0.0441082
R3730 VDD.n526 VDD.n525 0.0431316
R3731 VDD.n133 VDD.n132 0.0419894
R3732 VDD.n282 VDD.n281 0.0419894
R3733 VDD.n21 VDD.n19 0.0411098
R3734 VDD.n629 VDD.n627 0.0394691
R3735 VDD.n509 VDD.n506 0.0382246
R3736 VDD.n546 VDD.n545 0.0366722
R3737 VDD.n127 VDD.n126 0.0356064
R3738 VDD.n276 VDD.n275 0.0356064
R3739 VDD.n614 VDD.n613 0.0339021
R3740 VDD.n691 VDD.n690 0.0339021
R3741 VDD.n571 VDD.n570 0.0333378
R3742 VDD.n388 VDD.n383 0.031515
R3743 VDD.n649 VDD.n648 0.0301907
R3744 VDD.n257 VDD.n256 0.0296018
R3745 VDD.n644 VDD.n643 0.0292629
R3746 VDD.n109 VDD.n108 0.0282397
R3747 VDD.n12 VDD.n10 0.027939
R3748 VDD.n402 VDD.n262 0.0276213
R3749 VDD.n444 VDD.n443 0.0274492
R3750 VDD.n513 VDD.n512 0.0271986
R3751 VDD.n401 VDD.n399 0.0256786
R3752 VDD.n606 VDD.n604 0.0255515
R3753 VDD.n687 VDD.n686 0.0255515
R3754 VDD.n757 VDD.n756 0.0251951
R3755 VDD.n441 VDD.n440 0.0243983
R3756 VDD.n596 VDD.n595 0.0236959
R3757 VDD.n682 VDD.n681 0.0236959
R3758 VDD.n512 VDD.n445 0.023323
R3759 VDD.n759 VDD.n758 0.0224512
R3760 VDD.n731 VDD.n730 0.0220311
R3761 VDD.n718 VDD.n717 0.021875
R3762 VDD.n259 VDD.n258 0.021518
R3763 VDD.n261 VDD.n260 0.021518
R3764 VDD.n394 VDD.n393 0.0213929
R3765 VDD.n398 VDD.n397 0.0213929
R3766 VDD.n739 VDD.n736 0.0211699
R3767 VDD.n519 VDD.n516 0.0207392
R3768 VDD.n728 VDD.n727 0.0203086
R3769 VDD.n239 VDD.n238 0.0202326
R3770 VDD.n112 VDD.n111 0.0202326
R3771 VDD.n637 VDD.n636 0.0199845
R3772 VDD.n243 VDD.n242 0.0197513
R3773 VDD.n252 VDD.n251 0.0197513
R3774 VDD.n69 VDD.n66 0.0191585
R3775 VDD.n652 VDD.n651 0.0190567
R3776 VDD.n567 VDD.n566 0.0190167
R3777 VDD.n542 VDD.n541 0.0185861
R3778 VDD.n537 VDD.n536 0.0185861
R3779 VDD.n535 VDD.n530 0.0185861
R3780 VDD.n524 VDD.n519 0.0185861
R3781 VDD.n38 VDD.n37 0.018061
R3782 VDD.n588 VDD.n574 0.0176649
R3783 VDD.n527 VDD.n526 0.0167884
R3784 VDD.n677 VDD.n673 0.0167371
R3785 VDD.n740 VDD.n739 0.0161944
R3786 VDD.n716 VDD.n715 0.0158093
R3787 VDD.n530 VDD.n527 0.0154295
R3788 VDD.n624 VDD.n622 0.0153454
R3789 VDD.n696 VDD.n695 0.0153454
R3790 VDD.n92 VDD.n85 0.0153171
R3791 VDD.n56 VDD.n55 0.0147683
R3792 VDD.n740 VDD.n445 0.0145807
R3793 VDD VDD.n412 0.0140398
R3794 VDD VDD.n417 0.0140398
R3795 VDD VDD.n424 0.0140398
R3796 VDD VDD.n429 0.0140398
R3797 VDD VDD.n434 0.0140398
R3798 VDD VDD.n407 0.0140398
R3799 VDD.n716 VDD.n713 0.0139536
R3800 VDD.n763 VDD.n762 0.0136707
R3801 VDD VDD.n93 0.013122
R3802 VDD.n672 VDD.n671 0.0130258
R3803 VDD.n678 VDD.n677 0.0130258
R3804 VDD.n589 VDD.n588 0.0125619
R3805 VDD.n389 VDD.n388 0.0122857
R3806 VDD.n655 VDD.n654 0.0121334
R3807 VDD.n651 VDD.n650 0.0107062
R3808 VDD.n439 VDD.n438 0.0106695
R3809 VDD.n442 VDD.n441 0.0106695
R3810 VDD.n55 VDD.n48 0.010378
R3811 VDD.n572 VDD.n571 0.0102297
R3812 VDD.n260 VDD.n259 0.0102006
R3813 VDD.n397 VDD.n394 0.0101429
R3814 VDD.n140 VDD.n137 0.0100745
R3815 VDD.n289 VDD.n286 0.0100745
R3816 VDD.n756 VDD.n754 0.0100485
R3817 VDD.n93 VDD.n92 0.00982927
R3818 VDD.n619 VDD.n618 0.00977835
R3819 VDD.n525 VDD.n524 0.00954306
R3820 VDD.n41 VDD.n38 0.00933668
R3821 VDD.n762 VDD.n761 0.00928049
R3822 VDD.n551 VDD.n550 0.00911244
R3823 VDD.n536 VDD.n535 0.00911244
R3824 VDD.n516 VDD.n515 0.00911244
R3825 VDD.n77 VDD.n72 0.00876098
R3826 VDD VDD.n539 0.0082512
R3827 VDD.n59 VDD.n56 0.00824116
R3828 VDD.n247 VDD.n246 0.00820054
R3829 VDD.n250 VDD.n247 0.00820054
R3830 VDD.n85 VDD.n84 0.00805275
R3831 VDD.n242 VDD.n239 0.00771925
R3832 VDD.n741 VDD.n444 0.00761864
R3833 VDD.n729 VDD.n728 0.00738995
R3834 VDD.n107 VDD.n106 0.00728082
R3835 VDD.n37 VDD.n30 0.00708537
R3836 VDD.n727 VDD.n726 0.00684905
R3837 VDD.n761 VDD.n760 0.00653659
R3838 VDD.n736 VDD.n731 0.00652871
R3839 VDD.n715 VDD.n714 0.00606701
R3840 VDD.n392 VDD.n389 0.00585714
R3841 VDD.n641 VDD.n640 0.00513918
R3842 VDD.n705 VDD.n704 0.00513918
R3843 VDD.n768 VDD.n767 0.00434146
R3844 VDD.n760 VDD.n759 0.00269512
R3845 VDD.n72 VDD.n69 0.00214634
R3846 VDD.n655 VDD.n652 0.00192811
R3847 VDD.n568 VDD.n567 0.00179187
R3848 VDD.n570 VDD.n569 0.00171622
R3849 VDD.n601 VDD.n599 0.00142783
R3850 VDD.n560 VDD.n559 0.00136124
R3851 VDD.n749 VDD.n109 0.00111644
R3852 VDD.n673 VDD.n672 0.000963918
R3853 VDD.n514 VDD.n513 0.000930622
R3854 a_n2280_5855.n48 a_n2280_5855.t36 102.981
R3855 a_n2280_5855.n10 a_n2280_5855.t44 49.5689
R3856 a_n2280_5855.t36 a_n2280_5855.n47 49.5689
R3857 a_n2280_5855.n10 a_n2280_5855.t46 26.0719
R3858 a_n2280_5855.n11 a_n2280_5855.t43 26.0719
R3859 a_n2280_5855.n12 a_n2280_5855.t14 26.0719
R3860 a_n2280_5855.n13 a_n2280_5855.t16 26.0719
R3861 a_n2280_5855.n14 a_n2280_5855.t26 26.0719
R3862 a_n2280_5855.n15 a_n2280_5855.t27 26.0719
R3863 a_n2280_5855.n16 a_n2280_5855.t38 26.0719
R3864 a_n2280_5855.n17 a_n2280_5855.t51 26.0719
R3865 a_n2280_5855.n18 a_n2280_5855.t12 26.0719
R3866 a_n2280_5855.n19 a_n2280_5855.t21 26.0719
R3867 a_n2280_5855.n20 a_n2280_5855.t22 26.0719
R3868 a_n2280_5855.n21 a_n2280_5855.t35 26.0719
R3869 a_n2280_5855.n22 a_n2280_5855.t49 26.0719
R3870 a_n2280_5855.n23 a_n2280_5855.t40 26.0719
R3871 a_n2280_5855.n24 a_n2280_5855.t25 26.0719
R3872 a_n2280_5855.n25 a_n2280_5855.t23 26.0719
R3873 a_n2280_5855.n26 a_n2280_5855.t13 26.0719
R3874 a_n2280_5855.n27 a_n2280_5855.t42 26.0719
R3875 a_n2280_5855.n28 a_n2280_5855.t39 26.0719
R3876 a_n2280_5855.n29 a_n2280_5855.t29 26.0719
R3877 a_n2280_5855.n30 a_n2280_5855.t24 26.0719
R3878 a_n2280_5855.n31 a_n2280_5855.t15 26.0719
R3879 a_n2280_5855.n32 a_n2280_5855.t45 26.0719
R3880 a_n2280_5855.n33 a_n2280_5855.t41 26.0719
R3881 a_n2280_5855.n34 a_n2280_5855.t30 26.0719
R3882 a_n2280_5855.n35 a_n2280_5855.t28 26.0719
R3883 a_n2280_5855.n36 a_n2280_5855.t31 26.0719
R3884 a_n2280_5855.n37 a_n2280_5855.t18 26.0719
R3885 a_n2280_5855.n38 a_n2280_5855.t17 26.0719
R3886 a_n2280_5855.n39 a_n2280_5855.t48 26.0719
R3887 a_n2280_5855.n40 a_n2280_5855.t47 26.0719
R3888 a_n2280_5855.n41 a_n2280_5855.t32 26.0719
R3889 a_n2280_5855.n42 a_n2280_5855.t34 26.0719
R3890 a_n2280_5855.n43 a_n2280_5855.t33 26.0719
R3891 a_n2280_5855.n44 a_n2280_5855.t20 26.0719
R3892 a_n2280_5855.n45 a_n2280_5855.t19 26.0719
R3893 a_n2280_5855.n46 a_n2280_5855.t50 26.0719
R3894 a_n2280_5855.n47 a_n2280_5855.t37 26.0719
R3895 a_n2280_5855.n11 a_n2280_5855.n10 19.6341
R3896 a_n2280_5855.n12 a_n2280_5855.n11 19.6341
R3897 a_n2280_5855.n13 a_n2280_5855.n12 19.6341
R3898 a_n2280_5855.n14 a_n2280_5855.n13 19.6341
R3899 a_n2280_5855.n15 a_n2280_5855.n14 19.6341
R3900 a_n2280_5855.n16 a_n2280_5855.n15 19.6341
R3901 a_n2280_5855.n17 a_n2280_5855.n16 19.6341
R3902 a_n2280_5855.n18 a_n2280_5855.n17 19.6341
R3903 a_n2280_5855.n19 a_n2280_5855.n18 19.6341
R3904 a_n2280_5855.n20 a_n2280_5855.n19 19.6341
R3905 a_n2280_5855.n21 a_n2280_5855.n20 19.6341
R3906 a_n2280_5855.n22 a_n2280_5855.n21 19.6341
R3907 a_n2280_5855.n23 a_n2280_5855.n22 19.6341
R3908 a_n2280_5855.n24 a_n2280_5855.n23 19.6341
R3909 a_n2280_5855.n25 a_n2280_5855.n24 19.6341
R3910 a_n2280_5855.n26 a_n2280_5855.n25 19.6341
R3911 a_n2280_5855.n27 a_n2280_5855.n26 19.6341
R3912 a_n2280_5855.n28 a_n2280_5855.n27 19.6341
R3913 a_n2280_5855.n29 a_n2280_5855.n28 19.6341
R3914 a_n2280_5855.n30 a_n2280_5855.n29 19.6341
R3915 a_n2280_5855.n31 a_n2280_5855.n30 19.6341
R3916 a_n2280_5855.n32 a_n2280_5855.n31 19.6341
R3917 a_n2280_5855.n33 a_n2280_5855.n32 19.6341
R3918 a_n2280_5855.n34 a_n2280_5855.n33 19.6341
R3919 a_n2280_5855.n35 a_n2280_5855.n34 19.6341
R3920 a_n2280_5855.n36 a_n2280_5855.n35 19.6341
R3921 a_n2280_5855.n37 a_n2280_5855.n36 19.6341
R3922 a_n2280_5855.n38 a_n2280_5855.n37 19.6341
R3923 a_n2280_5855.n39 a_n2280_5855.n38 19.6341
R3924 a_n2280_5855.n40 a_n2280_5855.n39 19.6341
R3925 a_n2280_5855.n41 a_n2280_5855.n40 19.6341
R3926 a_n2280_5855.n42 a_n2280_5855.n41 19.6341
R3927 a_n2280_5855.n43 a_n2280_5855.n42 19.6341
R3928 a_n2280_5855.n44 a_n2280_5855.n43 19.6341
R3929 a_n2280_5855.n45 a_n2280_5855.n44 19.6341
R3930 a_n2280_5855.n46 a_n2280_5855.n45 19.6341
R3931 a_n2280_5855.n47 a_n2280_5855.n46 19.6341
R3932 a_n2280_5855.n50 a_n2280_5855.n3 3.7805
R3933 a_n2280_5855.n49 a_n2280_5855.n7 3.7805
R3934 a_n2280_5855.n52 a_n2280_5855.n50 3.7255
R3935 a_n2280_5855.n48 a_n2280_5855.n9 3.13775
R3936 a_n2280_5855.n50 a_n2280_5855.n1 3.09941
R3937 a_n2280_5855.n49 a_n2280_5855.n5 3.09941
R3938 a_n2280_5855.n9 a_n2280_5855.t1 0.9105
R3939 a_n2280_5855.n9 a_n2280_5855.n8 0.9105
R3940 a_n2280_5855.n1 a_n2280_5855.t4 0.9105
R3941 a_n2280_5855.n1 a_n2280_5855.n0 0.9105
R3942 a_n2280_5855.n5 a_n2280_5855.t5 0.9105
R3943 a_n2280_5855.n5 a_n2280_5855.n4 0.9105
R3944 a_n2280_5855.t7 a_n2280_5855.n52 0.9105
R3945 a_n2280_5855.n52 a_n2280_5855.n51 0.9105
R3946 a_n2280_5855.n3 a_n2280_5855.t9 0.8195
R3947 a_n2280_5855.n3 a_n2280_5855.n2 0.8195
R3948 a_n2280_5855.n7 a_n2280_5855.t10 0.8195
R3949 a_n2280_5855.n7 a_n2280_5855.n6 0.8195
R3950 a_n2280_5855.n50 a_n2280_5855.n49 0.626587
R3951 a_n2280_5855.n49 a_n2280_5855.n48 0.565935
R3952 OUT-.n99 OUT-.n96 3.81941
R3953 OUT-.n94 OUT-.n91 3.81941
R3954 OUT-.n89 OUT-.n86 3.81941
R3955 OUT-.n84 OUT-.n81 3.81941
R3956 OUT-.n79 OUT-.n76 3.81941
R3957 OUT-.n74 OUT-.n71 3.81941
R3958 OUT-.n69 OUT-.n66 3.81941
R3959 OUT-.n64 OUT-.n61 3.81941
R3960 OUT-.n59 OUT-.n56 3.81941
R3961 OUT-.n54 OUT-.n51 3.81941
R3962 OUT-.n49 OUT-.n46 3.81941
R3963 OUT-.n44 OUT-.n41 3.81941
R3964 OUT-.n39 OUT-.n36 3.81941
R3965 OUT-.n34 OUT-.n31 3.81941
R3966 OUT-.n29 OUT-.n26 3.81941
R3967 OUT-.n24 OUT-.n21 3.81941
R3968 OUT-.n19 OUT-.n16 3.81941
R3969 OUT-.n14 OUT-.n11 3.81941
R3970 OUT-.n9 OUT-.n6 3.81941
R3971 OUT-.n4 OUT-.n1 3.81941
R3972 OUT-.n99 OUT-.n98 3.1505
R3973 OUT-.n94 OUT-.n93 3.1505
R3974 OUT-.n89 OUT-.n88 3.1505
R3975 OUT-.n84 OUT-.n83 3.1505
R3976 OUT-.n79 OUT-.n78 3.1505
R3977 OUT-.n74 OUT-.n73 3.1505
R3978 OUT-.n69 OUT-.n68 3.1505
R3979 OUT-.n64 OUT-.n63 3.1505
R3980 OUT-.n59 OUT-.n58 3.1505
R3981 OUT-.n54 OUT-.n53 3.1505
R3982 OUT-.n49 OUT-.n48 3.1505
R3983 OUT-.n44 OUT-.n43 3.1505
R3984 OUT-.n39 OUT-.n38 3.1505
R3985 OUT-.n34 OUT-.n33 3.1505
R3986 OUT-.n29 OUT-.n28 3.1505
R3987 OUT-.n24 OUT-.n23 3.1505
R3988 OUT-.n19 OUT-.n18 3.1505
R3989 OUT-.n14 OUT-.n13 3.1505
R3990 OUT-.n9 OUT-.n8 3.1505
R3991 OUT-.n4 OUT-.n3 3.1505
R3992 OUT-.n96 OUT-.t47 0.9105
R3993 OUT-.n96 OUT-.n95 0.9105
R3994 OUT-.n91 OUT-.t40 0.9105
R3995 OUT-.n91 OUT-.n90 0.9105
R3996 OUT-.n86 OUT-.t55 0.9105
R3997 OUT-.n86 OUT-.n85 0.9105
R3998 OUT-.n81 OUT-.t48 0.9105
R3999 OUT-.n81 OUT-.n80 0.9105
R4000 OUT-.n76 OUT-.t42 0.9105
R4001 OUT-.n76 OUT-.n75 0.9105
R4002 OUT-.n71 OUT-.t56 0.9105
R4003 OUT-.n71 OUT-.n70 0.9105
R4004 OUT-.n66 OUT-.t49 0.9105
R4005 OUT-.n66 OUT-.n65 0.9105
R4006 OUT-.n61 OUT-.t50 0.9105
R4007 OUT-.n61 OUT-.n60 0.9105
R4008 OUT-.n56 OUT-.t44 0.9105
R4009 OUT-.n56 OUT-.n55 0.9105
R4010 OUT-.n51 OUT-.t53 0.9105
R4011 OUT-.n51 OUT-.n50 0.9105
R4012 OUT-.n46 OUT-.t45 0.9105
R4013 OUT-.n46 OUT-.n45 0.9105
R4014 OUT-.n41 OUT-.t58 0.9105
R4015 OUT-.n41 OUT-.n40 0.9105
R4016 OUT-.n36 OUT-.t52 0.9105
R4017 OUT-.n36 OUT-.n35 0.9105
R4018 OUT-.n31 OUT-.t41 0.9105
R4019 OUT-.n31 OUT-.n30 0.9105
R4020 OUT-.n26 OUT-.t54 0.9105
R4021 OUT-.n26 OUT-.n25 0.9105
R4022 OUT-.n21 OUT-.t59 0.9105
R4023 OUT-.n21 OUT-.n20 0.9105
R4024 OUT-.n16 OUT-.t46 0.9105
R4025 OUT-.n16 OUT-.n15 0.9105
R4026 OUT-.n11 OUT-.t51 0.9105
R4027 OUT-.n11 OUT-.n10 0.9105
R4028 OUT-.n6 OUT-.t57 0.9105
R4029 OUT-.n6 OUT-.n5 0.9105
R4030 OUT-.n1 OUT-.t43 0.9105
R4031 OUT-.n1 OUT-.n0 0.9105
R4032 OUT-.n98 OUT-.t18 0.8195
R4033 OUT-.n98 OUT-.n97 0.8195
R4034 OUT-.n93 OUT-.t11 0.8195
R4035 OUT-.n93 OUT-.n92 0.8195
R4036 OUT-.n88 OUT-.t6 0.8195
R4037 OUT-.n88 OUT-.n87 0.8195
R4038 OUT-.n83 OUT-.t19 0.8195
R4039 OUT-.n83 OUT-.n82 0.8195
R4040 OUT-.n78 OUT-.t13 0.8195
R4041 OUT-.n78 OUT-.n77 0.8195
R4042 OUT-.n73 OUT-.t7 0.8195
R4043 OUT-.n73 OUT-.n72 0.8195
R4044 OUT-.n68 OUT-.t0 0.8195
R4045 OUT-.n68 OUT-.n67 0.8195
R4046 OUT-.n63 OUT-.t1 0.8195
R4047 OUT-.n63 OUT-.n62 0.8195
R4048 OUT-.n58 OUT-.t15 0.8195
R4049 OUT-.n58 OUT-.n57 0.8195
R4050 OUT-.n53 OUT-.t4 0.8195
R4051 OUT-.n53 OUT-.n52 0.8195
R4052 OUT-.n48 OUT-.t16 0.8195
R4053 OUT-.n48 OUT-.n47 0.8195
R4054 OUT-.n43 OUT-.t9 0.8195
R4055 OUT-.n43 OUT-.n42 0.8195
R4056 OUT-.n38 OUT-.t3 0.8195
R4057 OUT-.n38 OUT-.n37 0.8195
R4058 OUT-.n33 OUT-.t12 0.8195
R4059 OUT-.n33 OUT-.n32 0.8195
R4060 OUT-.n28 OUT-.t5 0.8195
R4061 OUT-.n28 OUT-.n27 0.8195
R4062 OUT-.n23 OUT-.t10 0.8195
R4063 OUT-.n23 OUT-.n22 0.8195
R4064 OUT-.n18 OUT-.t17 0.8195
R4065 OUT-.n18 OUT-.n17 0.8195
R4066 OUT-.n13 OUT-.t2 0.8195
R4067 OUT-.n13 OUT-.n12 0.8195
R4068 OUT-.n8 OUT-.t8 0.8195
R4069 OUT-.n8 OUT-.n7 0.8195
R4070 OUT-.n3 OUT-.t14 0.8195
R4071 OUT-.n3 OUT-.n2 0.8195
R4072 OUT-.n100 OUT-.n99 0.730098
R4073 OUT-.n100 OUT-.n94 0.503326
R4074 OUT-.n101 OUT-.n89 0.503326
R4075 OUT-.n102 OUT-.n84 0.503326
R4076 OUT-.n103 OUT-.n79 0.503326
R4077 OUT-.n104 OUT-.n74 0.503326
R4078 OUT-.n105 OUT-.n69 0.503326
R4079 OUT-.n106 OUT-.n64 0.503326
R4080 OUT-.n107 OUT-.n59 0.503326
R4081 OUT-.n108 OUT-.n54 0.503326
R4082 OUT-.n109 OUT-.n49 0.503326
R4083 OUT-.n110 OUT-.n44 0.503326
R4084 OUT-.n111 OUT-.n39 0.503326
R4085 OUT-.n112 OUT-.n34 0.503326
R4086 OUT-.n113 OUT-.n29 0.503326
R4087 OUT-.n114 OUT-.n24 0.503326
R4088 OUT-.n115 OUT-.n19 0.503326
R4089 OUT-.n116 OUT-.n14 0.503326
R4090 OUT-.n117 OUT-.n9 0.503326
R4091 OUT-.n118 OUT-.n4 0.503326
R4092 OUT- OUT-.n118 0.267665
R4093 OUT-.n101 OUT-.n100 0.227272
R4094 OUT-.n102 OUT-.n101 0.227272
R4095 OUT-.n103 OUT-.n102 0.227272
R4096 OUT-.n104 OUT-.n103 0.227272
R4097 OUT-.n105 OUT-.n104 0.227272
R4098 OUT-.n106 OUT-.n105 0.227272
R4099 OUT-.n107 OUT-.n106 0.227272
R4100 OUT-.n108 OUT-.n107 0.227272
R4101 OUT-.n109 OUT-.n108 0.227272
R4102 OUT-.n110 OUT-.n109 0.227272
R4103 OUT-.n111 OUT-.n110 0.227272
R4104 OUT-.n112 OUT-.n111 0.227272
R4105 OUT-.n113 OUT-.n112 0.227272
R4106 OUT-.n114 OUT-.n113 0.227272
R4107 OUT-.n115 OUT-.n114 0.227272
R4108 OUT-.n116 OUT-.n115 0.227272
R4109 OUT-.n117 OUT-.n116 0.227272
R4110 OUT-.n118 OUT-.n117 0.227272
R4111 TG_1.IN.n260 TG_1.IN.t73 27.5082
R4112 TG_1.IN.n161 TG_1.IN.t15 18.6921
R4113 TG_1.IN.n87 TG_1.IN.t79 18.1625
R4114 TG_1.IN.n33 TG_1.IN.t59 17.9053
R4115 TG_1.IN.n23 TG_1.IN.t41 17.7975
R4116 TG_1.IN.n31 TG_1.IN.t11 17.7975
R4117 TG_1.IN.n108 TG_1.IN.t63 17.3759
R4118 TG_1.IN.n52 TG_1.IN.t65 17.0653
R4119 TG_1.IN.n193 TG_1.IN.t13 16.8013
R4120 TG_1.IN.n47 TG_1.IN.t87 16.6295
R4121 TG_1.IN.n49 TG_1.IN.t35 16.6295
R4122 TG_1.IN.n63 TG_1.IN.t43 16.5565
R4123 TG_1.IN.n34 TG_1.IN.t45 16.0963
R4124 TG_1.IN.n163 TG_1.IN.t47 15.9834
R4125 TG_1.IN.n261 TG_1.IN.t33 15.5061
R4126 TG_1.IN.n267 TG_1.IN.t91 14.8228
R4127 TG_1.IN.n66 TG_1.IN.t49 14.5125
R4128 TG_1.IN.n255 TG_1.IN.t27 14.3746
R4129 TG_1.IN.n68 TG_1.IN.t75 14.3665
R4130 TG_1.IN.n71 TG_1.IN.t23 14.3665
R4131 TG_1.IN.n112 TG_1.IN.t39 14.3665
R4132 TG_1.IN.n172 TG_1.IN.t25 13.5635
R4133 TG_1.IN.n120 TG_1.IN.t29 12.7025
R4134 TG_1.IN.n131 TG_1.IN.t85 12.5565
R4135 TG_1.IN.n126 TG_1.IN.t57 12.4105
R4136 TG_1.IN.n144 TG_1.IN.t67 12.3279
R4137 TG_1.IN.n207 TG_1.IN.t17 12.1185
R4138 TG_1.IN.n144 TG_1.IN.t61 11.6643
R4139 TG_1.IN.n394 TG_1.IN.n274 11.4676
R4140 TG_1.IN.n126 TG_1.IN.t53 11.4615
R4141 TG_1.IN.n131 TG_1.IN.t81 11.3155
R4142 TG_1.IN.n120 TG_1.IN.t19 11.1695
R4143 TG_1.IN.n226 TG_1.IN.t55 10.6585
R4144 TG_1.IN.n11 TG_1.IN.t31 10.5855
R4145 TG_1.IN.n226 TG_1.IN.t21 10.5125
R4146 TG_1.IN.n108 TG_1.IN.t89 10.2935
R4147 TG_1.IN.n250 TG_1.IN.t83 9.9285
R4148 TG_1.IN.n161 TG_1.IN.t69 9.9285
R4149 TG_1.IN.n100 TG_1.IN.n99 9.56292
R4150 TG_1.IN.n38 TG_1.IN.n36 9.14299
R4151 TG_1.IN.n207 TG_1.IN.t71 9.0525
R4152 TG_1.IN.n244 TG_1.IN.t101 8.54636
R4153 TG_1.IN.n238 TG_1.IN.t261 8.54439
R4154 TG_1.IN.n244 TG_1.IN.t99 8.50912
R4155 TG_1.IN.n274 TG_1.IN.t38 8.4005
R4156 TG_1.IN.n272 TG_1.IN.t84 8.4005
R4157 TG_1.IN.n250 TG_1.IN.t37 7.7385
R4158 TG_1.IN.n11 TG_1.IN.t77 7.6655
R4159 TG_1.IN.n261 TG_1.IN.n260 7.06268
R4160 TG_1.IN.n27 TG_1.IN.n26 6.58106
R4161 TG_1.IN.n128 TG_1.IN.t58 6.17646
R4162 TG_1.IN.n129 TG_1.IN.t54 6.14704
R4163 TG_1.IN.n0 TG_1.IN.t132 6.12938
R4164 TG_1.IN.n264 TG_1.IN.t74 6.1271
R4165 TG_1.IN.n50 TG_1.IN.t36 6.12579
R4166 TG_1.IN.n0 TG_1.IN.t141 6.11154
R4167 TG_1.IN.n223 TG_1.IN.t127 6.07519
R4168 TG_1.IN.n69 TG_1.IN.t76 6.07285
R4169 TG_1.IN.n223 TG_1.IN.t237 6.07152
R4170 TG_1.IN.n199 TG_1.IN.t126 6.03932
R4171 TG_1.IN.n178 TG_1.IN.n175 6.02244
R4172 TG_1.IN.n222 TG_1.IN.t125 6.00521
R4173 TG_1.IN.n247 TG_1.IN.n246 5.9303
R4174 TG_1.IN.n219 TG_1.IN.t140 5.8805
R4175 TG_1.IN.n200 TG_1.IN.t131 5.8805
R4176 TG_1.IN.n212 TG_1.IN.t236 5.8805
R4177 TG_1.IN.n210 TG_1.IN.n0 5.74421
R4178 TG_1.IN.n257 TG_1.IN.n256 5.5964
R4179 TG_1.IN.n8 TG_1.IN.t257 5.2505
R4180 TG_1.IN.n16 TG_1.IN.t117 5.2505
R4181 TG_1.IN.n16 TG_1.IN.t32 5.2505
R4182 TG_1.IN.n13 TG_1.IN.t258 5.2505
R4183 TG_1.IN.n13 TG_1.IN.t78 5.2505
R4184 TG_1.IN.n2 TG_1.IN.t100 5.2505
R4185 TG_1.IN.n1 TG_1.IN.t97 5.2505
R4186 TG_1.IN.n365 TG_1.IN.t172 5.18841
R4187 TG_1.IN.n196 TG_1.IN.n195 5.06613
R4188 TG_1.IN.n260 TG_1.IN.t51 4.3805
R4189 TG_1.IN.n364 TG_1.IN.n363 4.36941
R4190 TG_1.IN.n359 TG_1.IN.n358 4.36941
R4191 TG_1.IN.n354 TG_1.IN.n353 4.36941
R4192 TG_1.IN.n349 TG_1.IN.n348 4.36941
R4193 TG_1.IN.n344 TG_1.IN.n343 4.36941
R4194 TG_1.IN.n339 TG_1.IN.n338 4.36941
R4195 TG_1.IN.n334 TG_1.IN.n333 4.36941
R4196 TG_1.IN.n329 TG_1.IN.n328 4.36941
R4197 TG_1.IN.n324 TG_1.IN.n323 4.36941
R4198 TG_1.IN.n319 TG_1.IN.n318 4.36941
R4199 TG_1.IN.n314 TG_1.IN.n313 4.36941
R4200 TG_1.IN.n309 TG_1.IN.n308 4.36941
R4201 TG_1.IN.n304 TG_1.IN.n303 4.36941
R4202 TG_1.IN.n299 TG_1.IN.n298 4.36941
R4203 TG_1.IN.n294 TG_1.IN.n293 4.36941
R4204 TG_1.IN.n289 TG_1.IN.n288 4.36941
R4205 TG_1.IN.n284 TG_1.IN.n283 4.36941
R4206 TG_1.IN.n279 TG_1.IN.n278 4.36941
R4207 TG_1.IN.n374 TG_1.IN.n371 4.36941
R4208 TG_1.IN.n233 TG_1.IN.t256 4.36508
R4209 TG_1.IN.n255 TG_1.IN.t28 4.29173
R4210 TG_1.IN.n267 TG_1.IN.t92 4.22806
R4211 TG_1.IN.n268 TG_1.IN.t115 4.20189
R4212 TG_1.IN.n233 TG_1.IN.t259 4.201
R4213 TG_1.IN.n270 TG_1.IN.t116 4.15013
R4214 TG_1.IN.n256 TG_1.IN.t124 4.1302
R4215 TG_1.IN.n393 TG_1.IN.n392 4.08655
R4216 TG_1.IN.n121 TG_1.IN.n120 4.0005
R4217 TG_1.IN.n127 TG_1.IN.n126 4.0005
R4218 TG_1.IN.n132 TG_1.IN.n131 4.0005
R4219 TG_1.IN.n146 TG_1.IN.n144 4.0005
R4220 TG_1.IN.n162 TG_1.IN.n161 4.0005
R4221 TG_1.IN.n109 TG_1.IN.n108 4.0005
R4222 TG_1.IN.n208 TG_1.IN.n207 4.0005
R4223 TG_1.IN.n228 TG_1.IN.n226 4.0005
R4224 TG_1.IN.n12 TG_1.IN.n11 4.0005
R4225 TG_1.IN.n251 TG_1.IN.n250 4.0005
R4226 TG_1.IN.n262 TG_1.IN.n261 4.0005
R4227 TG_1.IN.n188 TG_1.IN.n187 3.74421
R4228 TG_1.IN.n142 TG_1.IN.n139 3.71646
R4229 TG_1.IN.n22 TG_1.IN.n19 3.6527
R4230 TG_1.IN.n154 TG_1.IN.n153 3.65144
R4231 TG_1.IN.n190 TG_1.IN.n189 3.64267
R4232 TG_1.IN.n76 TG_1.IN.n75 3.62822
R4233 TG_1.IN.n232 TG_1.IN.n101 3.57702
R4234 TG_1.IN.n269 TG_1.IN.n266 3.57312
R4235 TG_1.IN.n188 TG_1.IN.n182 3.55437
R4236 TG_1.IN.n191 TG_1.IN.n104 3.53697
R4237 TG_1.IN.n174 TG_1.IN.n170 3.51226
R4238 TG_1.IN.n365 TG_1.IN.t190 3.5105
R4239 TG_1.IN.n391 TG_1.IN.n390 3.5105
R4240 TG_1.IN.n168 TG_1.IN.n160 3.50854
R4241 TG_1.IN.n118 TG_1.IN.n117 3.47247
R4242 TG_1.IN.n231 TG_1.IN.n230 3.47027
R4243 TG_1.IN.n107 TG_1.IN.t90 3.46533
R4244 TG_1.IN.n88 TG_1.IN.n86 3.45237
R4245 TG_1.IN.n125 TG_1.IN.n124 3.44226
R4246 TG_1.IN.n187 TG_1.IN.n184 3.42242
R4247 TG_1.IN.n53 TG_1.IN.n45 3.41785
R4248 TG_1.IN.n123 TG_1.IN.n122 3.41123
R4249 TG_1.IN.n64 TG_1.IN.n62 3.40581
R4250 TG_1.IN.n135 TG_1.IN.n134 3.40419
R4251 TG_1.IN.n83 TG_1.IN.n82 3.40162
R4252 TG_1.IN.n48 TG_1.IN.n46 3.39579
R4253 TG_1.IN.n178 TG_1.IN.n177 3.39116
R4254 TG_1.IN.n239 TG_1.IN.n7 3.38977
R4255 TG_1.IN.n118 TG_1.IN.n115 3.38766
R4256 TG_1.IN.n217 TG_1.IN.n201 3.3856
R4257 TG_1.IN.n209 TG_1.IN.n205 3.38009
R4258 TG_1.IN.n99 TG_1.IN.n42 3.37847
R4259 TG_1.IN.n83 TG_1.IN.n80 3.36743
R4260 TG_1.IN.n263 TG_1.IN.n252 3.3665
R4261 TG_1.IN.n147 TG_1.IN.n143 3.36165
R4262 TG_1.IN.n217 TG_1.IN.n202 3.35805
R4263 TG_1.IN.n229 TG_1.IN.n225 3.35805
R4264 TG_1.IN.n7 TG_1.IN.t118 3.35317
R4265 TG_1.IN.n229 TG_1.IN.n224 3.35254
R4266 TG_1.IN.n187 TG_1.IN.n186 3.34851
R4267 TG_1.IN.n67 TG_1.IN.n65 3.34285
R4268 TG_1.IN.n113 TG_1.IN.n106 3.34109
R4269 TG_1.IN.n239 TG_1.IN.n238 3.33961
R4270 TG_1.IN.n14 TG_1.IN.n13 3.33223
R4271 TG_1.IN.n92 TG_1.IN.n89 3.32708
R4272 TG_1.IN.n72 TG_1.IN.n64 3.31948
R4273 TG_1.IN.n259 TG_1.IN.n258 3.31879
R4274 TG_1.IN.n173 TG_1.IN.n171 3.31638
R4275 TG_1.IN.n209 TG_1.IN.n204 3.31581
R4276 TG_1.IN.n198 TG_1.IN.n197 3.3125
R4277 TG_1.IN.n270 TG_1.IN.n269 3.29517
R4278 TG_1.IN.n249 TG_1.IN.n1 3.29336
R4279 TG_1.IN.n211 TG_1.IN.n203 3.2909
R4280 TG_1.IN.n221 TG_1.IN.n102 3.2783
R4281 TG_1.IN.n84 TG_1.IN.n83 3.27278
R4282 TG_1.IN.n257 TG_1.IN.n254 3.26657
R4283 TG_1.IN.n248 TG_1.IN.n2 3.23175
R4284 TG_1.IN.n394 TG_1.IN.n393 3.22511
R4285 TG_1.IN.n7 TG_1.IN.t260 3.20968
R4286 TG_1.IN.n234 TG_1.IN.n232 3.20101
R4287 TG_1.IN.n94 TG_1.IN.n93 3.1505
R4288 TG_1.IN.n77 TG_1.IN.n59 3.1505
R4289 TG_1.IN.n78 TG_1.IN.n57 3.1505
R4290 TG_1.IN.n85 TG_1.IN.n55 3.1505
R4291 TG_1.IN.n98 TG_1.IN.n43 3.1505
R4292 TG_1.IN.n36 TG_1.IN.n35 3.1505
R4293 TG_1.IN.n38 TG_1.IN.n37 3.1505
R4294 TG_1.IN.n22 TG_1.IN.n21 3.1505
R4295 TG_1.IN.n26 TG_1.IN.n25 3.1505
R4296 TG_1.IN.n30 TG_1.IN.n29 3.1505
R4297 TG_1.IN.n194 TG_1.IN.n192 3.1505
R4298 TG_1.IN.n149 TG_1.IN.n148 3.1505
R4299 TG_1.IN.n154 TG_1.IN.n151 3.1505
R4300 TG_1.IN.n142 TG_1.IN.n141 3.1505
R4301 TG_1.IN.n167 TG_1.IN.n166 3.1505
R4302 TG_1.IN.n179 TG_1.IN.n158 3.1505
R4303 TG_1.IN.n181 TG_1.IN.n137 3.1505
R4304 TG_1.IN.n17 TG_1.IN.n16 3.1505
R4305 TG_1.IN.n237 TG_1.IN.n8 3.1505
R4306 TG_1.IN.n241 TG_1.IN.n4 3.1505
R4307 TG_1.IN.n27 TG_1.IN.n22 3.14562
R4308 TG_1.IN.n84 TG_1.IN.n78 2.93789
R4309 TG_1.IN.n240 TG_1.IN.n239 2.82033
R4310 TG_1.IN.n85 TG_1.IN.n84 2.75648
R4311 TG_1.IN.n4 TG_1.IN.t2 2.7305
R4312 TG_1.IN.n4 TG_1.IN.n3 2.7305
R4313 TG_1.IN.n42 TG_1.IN.t102 2.7305
R4314 TG_1.IN.n42 TG_1.IN.t109 2.7305
R4315 TG_1.IN.n43 TG_1.IN.t123 2.7305
R4316 TG_1.IN.n43 TG_1.IN.t133 2.7305
R4317 TG_1.IN.n86 TG_1.IN.t250 2.7305
R4318 TG_1.IN.n86 TG_1.IN.t80 2.7305
R4319 TG_1.IN.n93 TG_1.IN.t136 2.7305
R4320 TG_1.IN.n93 TG_1.IN.t247 2.7305
R4321 TG_1.IN.n89 TG_1.IN.t104 2.7305
R4322 TG_1.IN.n89 TG_1.IN.t137 2.7305
R4323 TG_1.IN.n55 TG_1.IN.t253 2.7305
R4324 TG_1.IN.n55 TG_1.IN.n54 2.7305
R4325 TG_1.IN.n80 TG_1.IN.t98 2.7305
R4326 TG_1.IN.n80 TG_1.IN.n79 2.7305
R4327 TG_1.IN.n82 TG_1.IN.t251 2.7305
R4328 TG_1.IN.n82 TG_1.IN.n81 2.7305
R4329 TG_1.IN.n57 TG_1.IN.t252 2.7305
R4330 TG_1.IN.n57 TG_1.IN.n56 2.7305
R4331 TG_1.IN.n59 TG_1.IN.t249 2.7305
R4332 TG_1.IN.n59 TG_1.IN.n58 2.7305
R4333 TG_1.IN.n75 TG_1.IN.t95 2.7305
R4334 TG_1.IN.n75 TG_1.IN.n74 2.7305
R4335 TG_1.IN.n61 TG_1.IN.t24 2.7305
R4336 TG_1.IN.n61 TG_1.IN.n60 2.7305
R4337 TG_1.IN.n62 TG_1.IN.t248 2.7305
R4338 TG_1.IN.n62 TG_1.IN.t44 2.7305
R4339 TG_1.IN.n65 TG_1.IN.t50 2.7305
R4340 TG_1.IN.n45 TG_1.IN.t66 2.7305
R4341 TG_1.IN.n45 TG_1.IN.n44 2.7305
R4342 TG_1.IN.n46 TG_1.IN.t88 2.7305
R4343 TG_1.IN.n37 TG_1.IN.t107 2.7305
R4344 TG_1.IN.n37 TG_1.IN.t60 2.7305
R4345 TG_1.IN.n35 TG_1.IN.t245 2.7305
R4346 TG_1.IN.n35 TG_1.IN.t46 2.7305
R4347 TG_1.IN.n29 TG_1.IN.t12 2.7305
R4348 TG_1.IN.n29 TG_1.IN.n28 2.7305
R4349 TG_1.IN.n19 TG_1.IN.t255 2.7305
R4350 TG_1.IN.n19 TG_1.IN.n18 2.7305
R4351 TG_1.IN.n21 TG_1.IN.t106 2.7305
R4352 TG_1.IN.n21 TG_1.IN.n20 2.7305
R4353 TG_1.IN.n25 TG_1.IN.t42 2.7305
R4354 TG_1.IN.n25 TG_1.IN.n24 2.7305
R4355 TG_1.IN.n192 TG_1.IN.t244 2.7305
R4356 TG_1.IN.n192 TG_1.IN.t14 2.7305
R4357 TG_1.IN.n115 TG_1.IN.t120 2.7305
R4358 TG_1.IN.n115 TG_1.IN.n114 2.7305
R4359 TG_1.IN.n117 TG_1.IN.t234 2.7305
R4360 TG_1.IN.n117 TG_1.IN.n116 2.7305
R4361 TG_1.IN.n184 TG_1.IN.t243 2.7305
R4362 TG_1.IN.n184 TG_1.IN.n183 2.7305
R4363 TG_1.IN.n186 TG_1.IN.t228 2.7305
R4364 TG_1.IN.n186 TG_1.IN.n185 2.7305
R4365 TG_1.IN.n122 TG_1.IN.t20 2.7305
R4366 TG_1.IN.n124 TG_1.IN.t30 2.7305
R4367 TG_1.IN.n134 TG_1.IN.t82 2.7305
R4368 TG_1.IN.n134 TG_1.IN.n133 2.7305
R4369 TG_1.IN.n137 TG_1.IN.t86 2.7305
R4370 TG_1.IN.n137 TG_1.IN.n136 2.7305
R4371 TG_1.IN.n148 TG_1.IN.t230 2.7305
R4372 TG_1.IN.n148 TG_1.IN.t68 2.7305
R4373 TG_1.IN.n143 TG_1.IN.t232 2.7305
R4374 TG_1.IN.n143 TG_1.IN.t62 2.7305
R4375 TG_1.IN.n153 TG_1.IN.t93 2.7305
R4376 TG_1.IN.n153 TG_1.IN.n152 2.7305
R4377 TG_1.IN.n151 TG_1.IN.t227 2.7305
R4378 TG_1.IN.n151 TG_1.IN.n150 2.7305
R4379 TG_1.IN.n139 TG_1.IN.t240 2.7305
R4380 TG_1.IN.n139 TG_1.IN.n138 2.7305
R4381 TG_1.IN.n141 TG_1.IN.t10 2.7305
R4382 TG_1.IN.n141 TG_1.IN.n140 2.7305
R4383 TG_1.IN.n158 TG_1.IN.t233 2.7305
R4384 TG_1.IN.n158 TG_1.IN.n157 2.7305
R4385 TG_1.IN.n170 TG_1.IN.t226 2.7305
R4386 TG_1.IN.n170 TG_1.IN.n169 2.7305
R4387 TG_1.IN.n171 TG_1.IN.t239 2.7305
R4388 TG_1.IN.n171 TG_1.IN.t26 2.7305
R4389 TG_1.IN.n166 TG_1.IN.t70 2.7305
R4390 TG_1.IN.n166 TG_1.IN.t16 2.7305
R4391 TG_1.IN.n160 TG_1.IN.t48 2.7305
R4392 TG_1.IN.n160 TG_1.IN.n159 2.7305
R4393 TG_1.IN.n177 TG_1.IN.t8 2.7305
R4394 TG_1.IN.n177 TG_1.IN.n176 2.7305
R4395 TG_1.IN.n106 TG_1.IN.t40 2.7305
R4396 TG_1.IN.n106 TG_1.IN.n105 2.7305
R4397 TG_1.IN.n104 TG_1.IN.t231 2.7305
R4398 TG_1.IN.n104 TG_1.IN.n103 2.7305
R4399 TG_1.IN.n197 TG_1.IN.t139 2.7305
R4400 TG_1.IN.n205 TG_1.IN.t18 2.7305
R4401 TG_1.IN.n204 TG_1.IN.t72 2.7305
R4402 TG_1.IN.n203 TG_1.IN.t129 2.7305
R4403 TG_1.IN.n202 TG_1.IN.t238 2.7305
R4404 TG_1.IN.n201 TG_1.IN.t130 2.7305
R4405 TG_1.IN.n102 TG_1.IN.t142 2.7305
R4406 TG_1.IN.n225 TG_1.IN.t56 2.7305
R4407 TG_1.IN.n224 TG_1.IN.t22 2.7305
R4408 TG_1.IN.n6 TG_1.IN.t262 2.7305
R4409 TG_1.IN.n6 TG_1.IN.n5 2.7305
R4410 TG_1.IN.n254 TG_1.IN.n253 2.7305
R4411 TG_1.IN.n258 TG_1.IN.t34 2.7305
R4412 TG_1.IN.n252 TG_1.IN.t52 2.7305
R4413 TG_1.IN.n266 TG_1.IN.t135 2.7305
R4414 TG_1.IN.n266 TG_1.IN.n265 2.7305
R4415 TG_1.IN.n364 TG_1.IN.n361 2.6005
R4416 TG_1.IN.n359 TG_1.IN.n356 2.6005
R4417 TG_1.IN.n354 TG_1.IN.n351 2.6005
R4418 TG_1.IN.n349 TG_1.IN.n346 2.6005
R4419 TG_1.IN.n344 TG_1.IN.n341 2.6005
R4420 TG_1.IN.n339 TG_1.IN.n336 2.6005
R4421 TG_1.IN.n334 TG_1.IN.n331 2.6005
R4422 TG_1.IN.n329 TG_1.IN.n326 2.6005
R4423 TG_1.IN.n324 TG_1.IN.n321 2.6005
R4424 TG_1.IN.n319 TG_1.IN.n316 2.6005
R4425 TG_1.IN.n314 TG_1.IN.n311 2.6005
R4426 TG_1.IN.n309 TG_1.IN.n306 2.6005
R4427 TG_1.IN.n304 TG_1.IN.n301 2.6005
R4428 TG_1.IN.n299 TG_1.IN.n296 2.6005
R4429 TG_1.IN.n294 TG_1.IN.n291 2.6005
R4430 TG_1.IN.n289 TG_1.IN.n286 2.6005
R4431 TG_1.IN.n284 TG_1.IN.n281 2.6005
R4432 TG_1.IN.n279 TG_1.IN.n276 2.6005
R4433 TG_1.IN.n374 TG_1.IN.n373 2.6005
R4434 TG_1.IN.n30 TG_1.IN.n27 2.56342
R4435 TG_1.IN.n77 TG_1.IN.n76 2.52272
R4436 TG_1.IN.n269 TG_1.IN.n268 2.48586
R4437 TG_1.IN.n189 TG_1.IN.n118 2.2505
R4438 TG_1.IN.n231 TG_1.IN.n222 2.2505
R4439 TG_1.IN.n214 TG_1.IN.t235 2.05255
R4440 TG_1.IN.n76 TG_1.IN.n73 2.04187
R4441 TG_1.IN.n215 TG_1.IN.n214 1.94696
R4442 TG_1.IN.n232 TG_1.IN.n231 1.93866
R4443 TG_1.IN.n109 TG_1.IN.n107 1.85121
R4444 TG_1.IN.n214 TG_1.IN.t128 1.76935
R4445 TG_1.IN.n168 TG_1.IN.n167 1.59579
R4446 TG_1.IN.n101 TG_1.IN.n100 1.54309
R4447 TG_1.IN.n174 TG_1.IN.n173 1.50579
R4448 TG_1.IN.n240 TG_1.IN.n6 1.43159
R4449 TG_1.IN.n73 TG_1.IN.n61 1.42496
R4450 TG_1.IN.n107 TG_1.IN.t64 1.39688
R4451 TG_1.IN.n97 TG_1.IN.n96 1.35988
R4452 TG_1.IN.n235 TG_1.IN.n17 1.25562
R4453 TG_1.IN.n95 TG_1.IN.n88 1.04863
R4454 TG_1.IN.n271 TG_1.IN.n270 1.04839
R4455 TG_1.IN.n242 TG_1.IN.n241 1.04638
R4456 TG_1.IN.n155 TG_1.IN.n149 1.02685
R4457 TG_1.IN.n181 TG_1.IN.n180 1.02681
R4458 TG_1.IN.n191 TG_1.IN.n190 0.955153
R4459 TG_1.IN.n195 TG_1.IN.n194 0.945859
R4460 TG_1.IN.n361 TG_1.IN.t191 0.9105
R4461 TG_1.IN.n361 TG_1.IN.n360 0.9105
R4462 TG_1.IN.n356 TG_1.IN.t218 0.9105
R4463 TG_1.IN.n356 TG_1.IN.n355 0.9105
R4464 TG_1.IN.n351 TG_1.IN.t207 0.9105
R4465 TG_1.IN.n351 TG_1.IN.n350 0.9105
R4466 TG_1.IN.n346 TG_1.IN.t183 0.9105
R4467 TG_1.IN.n346 TG_1.IN.n345 0.9105
R4468 TG_1.IN.n341 TG_1.IN.t199 0.9105
R4469 TG_1.IN.n341 TG_1.IN.n340 0.9105
R4470 TG_1.IN.n336 TG_1.IN.t194 0.9105
R4471 TG_1.IN.n336 TG_1.IN.n335 0.9105
R4472 TG_1.IN.n331 TG_1.IN.t211 0.9105
R4473 TG_1.IN.n331 TG_1.IN.n330 0.9105
R4474 TG_1.IN.n326 TG_1.IN.t192 0.9105
R4475 TG_1.IN.n326 TG_1.IN.n325 0.9105
R4476 TG_1.IN.n321 TG_1.IN.t205 0.9105
R4477 TG_1.IN.n321 TG_1.IN.n320 0.9105
R4478 TG_1.IN.n316 TG_1.IN.t219 0.9105
R4479 TG_1.IN.n316 TG_1.IN.n315 0.9105
R4480 TG_1.IN.n311 TG_1.IN.t193 0.9105
R4481 TG_1.IN.n311 TG_1.IN.n310 0.9105
R4482 TG_1.IN.n306 TG_1.IN.t206 0.9105
R4483 TG_1.IN.n306 TG_1.IN.n305 0.9105
R4484 TG_1.IN.n301 TG_1.IN.t216 0.9105
R4485 TG_1.IN.n301 TG_1.IN.n300 0.9105
R4486 TG_1.IN.n296 TG_1.IN.t186 0.9105
R4487 TG_1.IN.n296 TG_1.IN.n295 0.9105
R4488 TG_1.IN.n291 TG_1.IN.t202 0.9105
R4489 TG_1.IN.n291 TG_1.IN.n290 0.9105
R4490 TG_1.IN.n286 TG_1.IN.t201 0.9105
R4491 TG_1.IN.n286 TG_1.IN.n285 0.9105
R4492 TG_1.IN.n281 TG_1.IN.t215 0.9105
R4493 TG_1.IN.n281 TG_1.IN.n280 0.9105
R4494 TG_1.IN.n276 TG_1.IN.t197 0.9105
R4495 TG_1.IN.n276 TG_1.IN.n275 0.9105
R4496 TG_1.IN.n373 TG_1.IN.t213 0.9105
R4497 TG_1.IN.n373 TG_1.IN.n372 0.9105
R4498 TG_1.IN.n220 TG_1.IN.n219 0.84268
R4499 TG_1.IN.n213 TG_1.IN.n212 0.840053
R4500 TG_1.IN.n195 TG_1.IN.n191 0.823637
R4501 TG_1.IN.n371 TG_1.IN.t155 0.8195
R4502 TG_1.IN.n371 TG_1.IN.n370 0.8195
R4503 TG_1.IN.n363 TG_1.IN.t173 0.8195
R4504 TG_1.IN.n363 TG_1.IN.n362 0.8195
R4505 TG_1.IN.n358 TG_1.IN.t160 0.8195
R4506 TG_1.IN.n358 TG_1.IN.n357 0.8195
R4507 TG_1.IN.n353 TG_1.IN.t149 0.8195
R4508 TG_1.IN.n353 TG_1.IN.n352 0.8195
R4509 TG_1.IN.n348 TG_1.IN.t165 0.8195
R4510 TG_1.IN.n348 TG_1.IN.n347 0.8195
R4511 TG_1.IN.n343 TG_1.IN.t181 0.8195
R4512 TG_1.IN.n343 TG_1.IN.n342 0.8195
R4513 TG_1.IN.n338 TG_1.IN.t176 0.8195
R4514 TG_1.IN.n338 TG_1.IN.n337 0.8195
R4515 TG_1.IN.n333 TG_1.IN.t153 0.8195
R4516 TG_1.IN.n333 TG_1.IN.n332 0.8195
R4517 TG_1.IN.n328 TG_1.IN.t174 0.8195
R4518 TG_1.IN.n328 TG_1.IN.n327 0.8195
R4519 TG_1.IN.n323 TG_1.IN.t147 0.8195
R4520 TG_1.IN.n323 TG_1.IN.n322 0.8195
R4521 TG_1.IN.n318 TG_1.IN.t161 0.8195
R4522 TG_1.IN.n318 TG_1.IN.n317 0.8195
R4523 TG_1.IN.n313 TG_1.IN.t175 0.8195
R4524 TG_1.IN.n313 TG_1.IN.n312 0.8195
R4525 TG_1.IN.n308 TG_1.IN.t148 0.8195
R4526 TG_1.IN.n308 TG_1.IN.n307 0.8195
R4527 TG_1.IN.n303 TG_1.IN.t158 0.8195
R4528 TG_1.IN.n303 TG_1.IN.n302 0.8195
R4529 TG_1.IN.n298 TG_1.IN.t168 0.8195
R4530 TG_1.IN.n298 TG_1.IN.n297 0.8195
R4531 TG_1.IN.n293 TG_1.IN.t144 0.8195
R4532 TG_1.IN.n293 TG_1.IN.n292 0.8195
R4533 TG_1.IN.n288 TG_1.IN.t143 0.8195
R4534 TG_1.IN.n288 TG_1.IN.n287 0.8195
R4535 TG_1.IN.n283 TG_1.IN.t157 0.8195
R4536 TG_1.IN.n283 TG_1.IN.n282 0.8195
R4537 TG_1.IN.n278 TG_1.IN.t179 0.8195
R4538 TG_1.IN.n278 TG_1.IN.n277 0.8195
R4539 TG_1.IN.n366 TG_1.IN.n365 0.688999
R4540 TG_1.IN.n175 TG_1.IN.n168 0.68553
R4541 TG_1.IN.n175 TG_1.IN.n174 0.681061
R4542 TG_1.IN.n200 TG_1.IN.n199 0.672487
R4543 TG_1.IN.n180 TG_1.IN.n156 0.661654
R4544 TG_1.IN.n156 TG_1.IN.n155 0.658192
R4545 TG_1.IN.n96 TG_1.IN.n95 0.61175
R4546 TG_1.IN.n96 TG_1.IN.n85 0.563
R4547 TG_1.IN.n78 TG_1.IN.n77 0.549186
R4548 TG_1.IN.n190 TG_1.IN.n113 0.532045
R4549 TG_1.IN.n212 TG_1.IN.n211 0.505815
R4550 TG_1.IN.n221 TG_1.IN.n220 0.4919
R4551 TG_1.IN.n256 TG_1.IN.n255 0.482612
R4552 TG_1.IN.n366 TG_1.IN.n364 0.481804
R4553 TG_1.IN.n367 TG_1.IN.n359 0.481804
R4554 TG_1.IN.n368 TG_1.IN.n354 0.481804
R4555 TG_1.IN.n369 TG_1.IN.n349 0.481804
R4556 TG_1.IN.n376 TG_1.IN.n344 0.481804
R4557 TG_1.IN.n377 TG_1.IN.n339 0.481804
R4558 TG_1.IN.n378 TG_1.IN.n334 0.481804
R4559 TG_1.IN.n379 TG_1.IN.n329 0.481804
R4560 TG_1.IN.n380 TG_1.IN.n324 0.481804
R4561 TG_1.IN.n381 TG_1.IN.n319 0.481804
R4562 TG_1.IN.n382 TG_1.IN.n314 0.481804
R4563 TG_1.IN.n383 TG_1.IN.n309 0.481804
R4564 TG_1.IN.n384 TG_1.IN.n304 0.481804
R4565 TG_1.IN.n385 TG_1.IN.n299 0.481804
R4566 TG_1.IN.n386 TG_1.IN.n294 0.481804
R4567 TG_1.IN.n387 TG_1.IN.n289 0.481804
R4568 TG_1.IN.n388 TG_1.IN.n284 0.481804
R4569 TG_1.IN.n389 TG_1.IN.n279 0.481804
R4570 TG_1.IN.n375 TG_1.IN.n374 0.481804
R4571 TG_1.IN.n241 TG_1.IN.n240 0.481551
R4572 TG_1.IN.n268 TG_1.IN.n267 0.460088
R4573 TG_1.IN.n271 TG_1.IN.n264 0.4595
R4574 TG_1.IN.n198 TG_1.IN.n196 0.44352
R4575 TG_1.IN.n391 TG_1.IN.n389 0.437328
R4576 TG_1.IN.n393 TG_1.IN.n391 0.434305
R4577 TG_1.IN.n26 TG_1.IN.n23 0.421942
R4578 TG_1.IN.n234 TG_1.IN.n233 0.420112
R4579 TG_1.IN.n218 TG_1.IN.n217 0.380704
R4580 TG_1.IN.n95 TG_1.IN.n94 0.377076
R4581 TG_1.IN.n194 TG_1.IN.n193 0.374377
R4582 TG_1.IN.n217 TG_1.IN.n216 0.369684
R4583 TG_1.IN.n156 TG_1.IN.n142 0.365692
R4584 TG_1.IN.n36 TG_1.IN.n34 0.364915
R4585 TG_1.IN.n98 TG_1.IN.n97 0.358735
R4586 TG_1.IN.n235 TG_1.IN.n234 0.355045
R4587 TG_1.IN.n39 TG_1.IN.n38 0.344664
R4588 TG_1.IN.n263 TG_1.IN.n262 0.332093
R4589 TG_1.IN.n92 TG_1.IN.n90 0.3305
R4590 TG_1.IN.n264 TG_1.IN.n263 0.3299
R4591 TG_1.IN.n222 TG_1.IN.n221 0.326814
R4592 TG_1.IN.n15 TG_1.IN.n9 0.324154
R4593 TG_1.IN.n92 TG_1.IN.n91 0.321026
R4594 TG_1.IN.n259 TG_1.IN.n257 0.3083
R4595 TG_1.IN.n99 TG_1.IN.n41 0.2905
R4596 TG_1.IN.n199 TG_1.IN.n198 0.287031
R4597 TG_1.IN.n189 TG_1.IN.n188 0.280143
R4598 TG_1.IN.n99 TG_1.IN.n40 0.272167
R4599 TG_1.IN.n211 TG_1.IN.n210 0.266717
R4600 TG_1.IN.n182 TG_1.IN.n181 0.266607
R4601 TG_1.IN.n32 TG_1.IN.n31 0.265864
R4602 TG_1.IN.n0 TG_1.IN.n209 0.265586
R4603 TG_1.IN.n165 TG_1.IN.n164 0.259092
R4604 TG_1.IN.n155 TG_1.IN.n154 0.258613
R4605 TG_1.IN.n180 TG_1.IN.n179 0.258613
R4606 TG_1.IN.n230 TG_1.IN.n229 0.255409
R4607 TG_1.IN.n216 TG_1.IN.n213 0.233471
R4608 TG_1.IN.n219 TG_1.IN.n218 0.233471
R4609 TG_1.IN.n149 TG_1.IN.n147 0.227231
R4610 TG_1.IN.n99 TG_1.IN.n98 0.226104
R4611 TG_1.IN.n179 TG_1.IN.n178 0.223476
R4612 TG_1.IN.n17 TG_1.IN.n15 0.221668
R4613 TG_1.IN.n389 TG_1.IN.n388 0.207694
R4614 TG_1.IN.n388 TG_1.IN.n387 0.207694
R4615 TG_1.IN.n387 TG_1.IN.n386 0.207694
R4616 TG_1.IN.n386 TG_1.IN.n385 0.207694
R4617 TG_1.IN.n385 TG_1.IN.n384 0.207694
R4618 TG_1.IN.n384 TG_1.IN.n383 0.207694
R4619 TG_1.IN.n383 TG_1.IN.n382 0.207694
R4620 TG_1.IN.n382 TG_1.IN.n381 0.207694
R4621 TG_1.IN.n381 TG_1.IN.n380 0.207694
R4622 TG_1.IN.n380 TG_1.IN.n379 0.207694
R4623 TG_1.IN.n379 TG_1.IN.n378 0.207694
R4624 TG_1.IN.n378 TG_1.IN.n377 0.207694
R4625 TG_1.IN.n377 TG_1.IN.n376 0.207694
R4626 TG_1.IN.n376 TG_1.IN.n375 0.207694
R4627 TG_1.IN.n375 TG_1.IN.n369 0.207694
R4628 TG_1.IN.n369 TG_1.IN.n368 0.207694
R4629 TG_1.IN.n368 TG_1.IN.n367 0.207694
R4630 TG_1.IN.n367 TG_1.IN.n366 0.207694
R4631 TG_1.IN.n218 TG_1.IN.n200 0.20592
R4632 TG_1.IN.n216 TG_1.IN.n215 0.20592
R4633 TG_1.IN.n94 TG_1.IN.n92 0.198742
R4634 TG_1.IN.n273 TG_1.IN.n272 0.194429
R4635 TG_1.IN.n32 TG_1.IN.n30 0.193426
R4636 TG_1.IN.n236 TG_1.IN.n235 0.185594
R4637 TG_1.IN.n272 TG_1.IN.n271 0.185121
R4638 TG_1.IN.n238 TG_1.IN.n237 0.183725
R4639 TG_1.IN.n97 TG_1.IN.n53 0.182375
R4640 TG_1.IN.n167 TG_1.IN.n165 0.1805
R4641 TG_1.IN.n73 TG_1.IN.n72 0.180219
R4642 TG_1.IN.n70 TG_1.IN.n69 0.177731
R4643 TG_1.IN.n111 TG_1.IN.n110 0.172572
R4644 TG_1.IN.n274 TG_1.IN.n273 0.1505
R4645 TG_1.IN.n12 TG_1.IN.n10 0.145885
R4646 TG_1.IN.n243 TG_1.IN.n242 0.143357
R4647 TG_1.IN.n68 TG_1.IN.n67 0.143115
R4648 TG_1.IN.n69 TG_1.IN.n68 0.143115
R4649 TG_1.IN.n64 TG_1.IN.n63 0.141731
R4650 TG_1.IN.n237 TG_1.IN.n236 0.141474
R4651 TG_1.IN.n71 TG_1.IN.n70 0.140346
R4652 TG_1.IN.n72 TG_1.IN.n71 0.140346
R4653 TG_1.IN.n121 TG_1.IN.n119 0.140346
R4654 TG_1.IN.n246 TG_1.IN.n245 0.138962
R4655 TG_1.IN.n228 TG_1.IN.n227 0.138858
R4656 TG_1.IN.n88 TG_1.IN.n87 0.138227
R4657 TG_1.IN.n48 TG_1.IN.n47 0.137515
R4658 TG_1.IN.n49 TG_1.IN.n48 0.137515
R4659 TG_1.IN.n50 TG_1.IN.n49 0.137515
R4660 TG_1.IN.n229 TG_1.IN.n228 0.137515
R4661 TG_1.IN.n67 TG_1.IN.n66 0.136734
R4662 TG_1.IN.n51 TG_1.IN.n50 0.136172
R4663 TG_1.IN.n110 TG_1.IN.n109 0.135487
R4664 TG_1.IN.n53 TG_1.IN.n52 0.134808
R4665 TG_1.IN.n113 TG_1.IN.n112 0.134176
R4666 TG_1.IN.n130 TG_1.IN.n129 0.132929
R4667 TG_1.IN.n112 TG_1.IN.n111 0.131529
R4668 TG_1.IN.n165 TG_1.IN.n162 0.131063
R4669 TG_1.IN.n164 TG_1.IN.n163 0.131063
R4670 TG_1.IN.n251 TG_1.IN.n249 0.129461
R4671 TG_1.IN.n132 TG_1.IN.n130 0.129071
R4672 TG_1.IN.n247 TG_1.IN.n243 0.127903
R4673 TG_1.IN.n173 TG_1.IN.n172 0.126253
R4674 TG_1.IN.n209 TG_1.IN.n208 0.1253
R4675 TG_1.IN.n147 TG_1.IN.n146 0.124554
R4676 TG_1.IN.n146 TG_1.IN.n145 0.122122
R4677 TG_1.IN.n208 TG_1.IN.n206 0.1217
R4678 TG_1.IN.n52 TG_1.IN.n51 0.120473
R4679 TG_1.IN.n101 TG_1.IN.n32 0.119848
R4680 TG_1.IN.n248 TG_1.IN.n247 0.118552
R4681 TG_1.IN.n14 TG_1.IN.n12 0.109885
R4682 TG_1.IN.n273 TG_1.IN.n251 0.108227
R4683 TG_1.IN.n246 TG_1.IN.n244 0.106654
R4684 TG_1.IN.n123 TG_1.IN.n121 0.101577
R4685 TG_1.IN.n128 TG_1.IN.n127 0.100935
R4686 TG_1.IN.n127 TG_1.IN.n125 0.0983261
R4687 TG_1.IN.n262 TG_1.IN.n259 0.0860738
R4688 TG_1.IN.n100 TG_1.IN.n39 0.0846936
R4689 TG_1.IN.n135 TG_1.IN.n132 0.0815
R4690 TG_1.IN.n39 TG_1.IN.n33 0.0527857
R4691 TG_1.IN.n230 TG_1.IN.n223 0.046625
R4692 TG_1.IN.n15 TG_1.IN.n14 0.0264615
R4693 TG_1.IN.n182 TG_1.IN.n135 0.0141364
R4694 TG_1.IN TG_1.IN.n394 0.00772628
R4695 TG_1.IN.n249 TG_1.IN.n248 0.00634416
R4696 TG_1.IN.n125 TG_1.IN.n123 0.00532143
R4697 TG_1.IN.n129 TG_1.IN.n128 0.00396154
R4698 SDn_2.n66 SDn_2.n65 83.0274
R4699 SDn_2 SDn_2.n64 57.7204
R4700 SDn_2.n65 SDn_2.n33 50.5649
R4701 SDn_2.n74 SDn_2.n73 48.6672
R4702 SDn_2.n101 SDn_2.n100 47.4505
R4703 SDn_2.n3 SDn_2.t66 35.1054
R4704 SDn_2.n94 SDn_2.t84 34.0104
R4705 SDn_2.n34 SDn_2.t87 33.7184
R4706 SDn_2.n104 SDn_2.n103 21.2922
R4707 SDn_2.n95 SDn_2.n94 21.0894
R4708 SDn_2.n96 SDn_2.n95 21.0894
R4709 SDn_2.n97 SDn_2.n96 21.0894
R4710 SDn_2.n98 SDn_2.n97 21.0894
R4711 SDn_2.n99 SDn_2.n98 21.0894
R4712 SDn_2.n100 SDn_2.n99 21.0894
R4713 SDn_2.n102 SDn_2.n101 21.0894
R4714 SDn_2.n104 SDn_2.n102 21.0894
R4715 SDn_2.n76 SDn_2.n75 21.0894
R4716 SDn_2.n4 SDn_2.n3 21.0894
R4717 SDn_2.n5 SDn_2.n4 21.0894
R4718 SDn_2.n6 SDn_2.n5 21.0894
R4719 SDn_2.n7 SDn_2.n6 21.0894
R4720 SDn_2.n8 SDn_2.n7 21.0894
R4721 SDn_2.n9 SDn_2.n8 21.0894
R4722 SDn_2.n10 SDn_2.n9 21.0894
R4723 SDn_2.n11 SDn_2.n10 21.0894
R4724 SDn_2.n12 SDn_2.n11 21.0894
R4725 SDn_2.n13 SDn_2.n12 21.0894
R4726 SDn_2.n14 SDn_2.n13 21.0894
R4727 SDn_2.n15 SDn_2.n14 21.0894
R4728 SDn_2.n16 SDn_2.n15 21.0894
R4729 SDn_2.n17 SDn_2.n16 21.0894
R4730 SDn_2.n18 SDn_2.n17 21.0894
R4731 SDn_2.n19 SDn_2.n18 21.0894
R4732 SDn_2.n20 SDn_2.n19 21.0894
R4733 SDn_2.n21 SDn_2.n20 21.0894
R4734 SDn_2.n22 SDn_2.n21 21.0894
R4735 SDn_2.n23 SDn_2.n22 21.0894
R4736 SDn_2.n24 SDn_2.n23 21.0894
R4737 SDn_2.n25 SDn_2.n24 21.0894
R4738 SDn_2.n26 SDn_2.n25 21.0894
R4739 SDn_2.n27 SDn_2.n26 21.0894
R4740 SDn_2.n28 SDn_2.n27 21.0894
R4741 SDn_2.n29 SDn_2.n28 21.0894
R4742 SDn_2.n30 SDn_2.n29 21.0894
R4743 SDn_2.n31 SDn_2.n30 21.0894
R4744 SDn_2.n32 SDn_2.n31 21.0894
R4745 SDn_2.n33 SDn_2.n32 21.0894
R4746 SDn_2.n35 SDn_2.n34 21.0894
R4747 SDn_2.n36 SDn_2.n35 21.0894
R4748 SDn_2.n37 SDn_2.n36 21.0894
R4749 SDn_2.n38 SDn_2.n37 21.0894
R4750 SDn_2.n39 SDn_2.n38 21.0894
R4751 SDn_2.n40 SDn_2.n39 21.0894
R4752 SDn_2.n41 SDn_2.n40 21.0894
R4753 SDn_2.n42 SDn_2.n41 21.0894
R4754 SDn_2.n43 SDn_2.n42 21.0894
R4755 SDn_2.n44 SDn_2.n43 21.0894
R4756 SDn_2.n45 SDn_2.n44 21.0894
R4757 SDn_2.n46 SDn_2.n45 21.0894
R4758 SDn_2.n47 SDn_2.n46 21.0894
R4759 SDn_2.n48 SDn_2.n47 21.0894
R4760 SDn_2.n49 SDn_2.n48 21.0894
R4761 SDn_2.n50 SDn_2.n49 21.0894
R4762 SDn_2.n51 SDn_2.n50 21.0894
R4763 SDn_2.n52 SDn_2.n51 21.0894
R4764 SDn_2.n53 SDn_2.n52 21.0894
R4765 SDn_2.n54 SDn_2.n53 21.0894
R4766 SDn_2.n55 SDn_2.n54 21.0894
R4767 SDn_2.n56 SDn_2.n55 21.0894
R4768 SDn_2.n57 SDn_2.n56 21.0894
R4769 SDn_2.n58 SDn_2.n57 21.0894
R4770 SDn_2.n59 SDn_2.n58 21.0894
R4771 SDn_2.n60 SDn_2.n59 21.0894
R4772 SDn_2.n61 SDn_2.n60 21.0894
R4773 SDn_2.n62 SDn_2.n61 21.0894
R4774 SDn_2.n63 SDn_2.n62 21.0894
R4775 SDn_2.n64 SDn_2.n63 21.0894
R4776 SDn_2.n67 SDn_2.n66 21.0894
R4777 SDn_2.n68 SDn_2.n67 21.0894
R4778 SDn_2.n69 SDn_2.n68 21.0894
R4779 SDn_2.n70 SDn_2.n69 21.0894
R4780 SDn_2.n71 SDn_2.n70 21.0894
R4781 SDn_2.n72 SDn_2.n71 21.0894
R4782 SDn_2.n73 SDn_2.n72 21.0894
R4783 SDn_2.n77 SDn_2.n74 21.0894
R4784 SDn_2.n77 SDn_2.n76 21.0894
R4785 SDn_2.n65 SDn_2 14.9729
R4786 SDn_2.n3 SDn_2.t89 14.7465
R4787 SDn_2.n4 SDn_2.t106 14.7465
R4788 SDn_2.n7 SDn_2.t49 14.7465
R4789 SDn_2.n8 SDn_2.t95 14.7465
R4790 SDn_2.n11 SDn_2.t97 14.7465
R4791 SDn_2.n12 SDn_2.t76 14.7465
R4792 SDn_2.n15 SDn_2.t61 14.7465
R4793 SDn_2.n16 SDn_2.t104 14.7465
R4794 SDn_2.n19 SDn_2.t103 14.7465
R4795 SDn_2.n20 SDn_2.t85 14.7465
R4796 SDn_2.n23 SDn_2.t65 14.7465
R4797 SDn_2.n24 SDn_2.t36 14.7465
R4798 SDn_2.n27 SDn_2.t24 14.7465
R4799 SDn_2.n28 SDn_2.t71 14.7465
R4800 SDn_2.n31 SDn_2.t74 14.7465
R4801 SDn_2.n32 SDn_2.t54 14.7465
R4802 SDn_2.n94 SDn_2.t69 14.3815
R4803 SDn_2.n95 SDn_2.t88 14.3815
R4804 SDn_2.n98 SDn_2.t72 14.3815
R4805 SDn_2.n99 SDn_2.t38 14.3815
R4806 SDn_2.n102 SDn_2.t12 14.3815
R4807 SDn_2.n76 SDn_2.t10 14.3815
R4808 SDn_2.n67 SDn_2.t94 14.3815
R4809 SDn_2.n68 SDn_2.t51 14.3815
R4810 SDn_2.n71 SDn_2.t39 14.3815
R4811 SDn_2.n72 SDn_2.t68 14.3815
R4812 SDn_2.n5 SDn_2.t92 14.0165
R4813 SDn_2.n6 SDn_2.t46 14.0165
R4814 SDn_2.n9 SDn_2.t47 14.0165
R4815 SDn_2.n10 SDn_2.t62 14.0165
R4816 SDn_2.n13 SDn_2.t55 14.0165
R4817 SDn_2.n14 SDn_2.t29 14.0165
R4818 SDn_2.n17 SDn_2.t98 14.0165
R4819 SDn_2.n18 SDn_2.t57 14.0165
R4820 SDn_2.n21 SDn_2.t64 14.0165
R4821 SDn_2.n22 SDn_2.t34 14.0165
R4822 SDn_2.n25 SDn_2.t42 14.0165
R4823 SDn_2.n26 SDn_2.t86 14.0165
R4824 SDn_2.n29 SDn_2.t67 14.0165
R4825 SDn_2.n30 SDn_2.t52 14.0165
R4826 SDn_2.n33 SDn_2.t25 14.0165
R4827 SDn_2.n34 SDn_2.t40 13.3595
R4828 SDn_2.n35 SDn_2.t77 13.3595
R4829 SDn_2.n38 SDn_2.t30 13.3595
R4830 SDn_2.n39 SDn_2.t90 13.3595
R4831 SDn_2.n42 SDn_2.t43 13.3595
R4832 SDn_2.n43 SDn_2.t78 13.3595
R4833 SDn_2.n46 SDn_2.t99 13.3595
R4834 SDn_2.n47 SDn_2.t70 13.3595
R4835 SDn_2.n50 SDn_2.t101 13.3595
R4836 SDn_2.n51 SDn_2.t105 13.3595
R4837 SDn_2.n54 SDn_2.t27 13.3595
R4838 SDn_2.n55 SDn_2.t82 13.3595
R4839 SDn_2.n58 SDn_2.t45 13.3595
R4840 SDn_2.n59 SDn_2.t79 13.3595
R4841 SDn_2.n62 SDn_2.t32 13.3595
R4842 SDn_2.n63 SDn_2.t91 13.3595
R4843 SDn_2.n101 SDn_2.t6 12.9916
R4844 SDn_2.n103 SDn_2.t4 12.9916
R4845 SDn_2.n75 SDn_2.t0 12.9916
R4846 SDn_2.n96 SDn_2.t58 12.9215
R4847 SDn_2.n97 SDn_2.t50 12.9215
R4848 SDn_2.n100 SDn_2.t73 12.9215
R4849 SDn_2.n66 SDn_2.t75 12.9215
R4850 SDn_2.n69 SDn_2.t48 12.9215
R4851 SDn_2.n70 SDn_2.t37 12.9215
R4852 SDn_2.n73 SDn_2.t33 12.9215
R4853 SDn_2.n74 SDn_2.t14 12.9215
R4854 SDn_2.n36 SDn_2.t31 12.6295
R4855 SDn_2.n37 SDn_2.t100 12.6295
R4856 SDn_2.n40 SDn_2.t44 12.6295
R4857 SDn_2.n41 SDn_2.t81 12.6295
R4858 SDn_2.n44 SDn_2.t26 12.6295
R4859 SDn_2.n45 SDn_2.t63 12.6295
R4860 SDn_2.n48 SDn_2.t107 12.6295
R4861 SDn_2.n49 SDn_2.t80 12.6295
R4862 SDn_2.n52 SDn_2.t35 12.6295
R4863 SDn_2.n53 SDn_2.t96 12.6295
R4864 SDn_2.n56 SDn_2.t60 12.6295
R4865 SDn_2.n57 SDn_2.t93 12.6295
R4866 SDn_2.n60 SDn_2.t59 12.6295
R4867 SDn_2.n61 SDn_2.t102 12.6295
R4868 SDn_2.n64 SDn_2.t41 12.6295
R4869 SDn_2.n106 SDn_2.t2 10.7743
R4870 SDn_2.n79 SDn_2.t8 10.7743
R4871 SDn_2.n107 SDn_2.n105 3.54502
R4872 SDn_2.n80 SDn_2.n78 3.54477
R4873 SDn_2.n107 SDn_2.n106 3.50535
R4874 SDn_2.n80 SDn_2.n79 3.50535
R4875 SDn_2.n91 SDn_2.n88 3.07598
R4876 SDn_2.n117 SDn_2.n84 3.01065
R4877 SDn_2.n86 SDn_2.n85 2.90221
R4878 SDn_2.n114 SDn_2.n113 2.90214
R4879 SDn_2.n109 SDn_2.n108 2.88451
R4880 SDn_2.n81 SDn_2.n2 2.88438
R4881 SDn_2.n93 SDn_2.n92 2.87834
R4882 SDn_2.n88 SDn_2.n87 2.87828
R4883 SDn_2.n90 SDn_2.n89 2.87828
R4884 SDn_2.n84 SDn_2.n83 2.82902
R4885 SDn_2.n82 SDn_2.n1 2.76772
R4886 SDn_2.n110 SDn_2.n93 2.75462
R4887 SDn_2.n1 SDn_2.t16 2.7305
R4888 SDn_2.n1 SDn_2.n0 2.7305
R4889 SDn_2.n122 SDn_2.t9 2.7305
R4890 SDn_2.n122 SDn_2.n121 2.7305
R4891 SDn_2.n91 SDn_2.n90 2.50797
R4892 SDn_2.n112 SDn_2.n86 2.50522
R4893 SDn_2.n84 SDn_2.t1 2.49942
R4894 SDn_2.n90 SDn_2.t19 2.43824
R4895 SDn_2.n88 SDn_2.t7 2.43824
R4896 SDn_2.n93 SDn_2.t20 2.4382
R4897 SDn_2.n114 SDn_2.t18 2.40701
R4898 SDn_2.n86 SDn_2.t3 2.40696
R4899 SDn_2.n110 SDn_2.n109 2.35277
R4900 SDn_2.n82 SDn_2.n81 2.3515
R4901 SDn_2.n116 SDn_2.n115 2.24989
R4902 SDn_2.n125 SDn_2.n124 1.50283
R4903 SDn_2.n123 SDn_2.n122 1.42666
R4904 SDn_2.n115 SDn_2.n114 1.0106
R4905 SDn_2.n78 SDn_2.n77 0.967483
R4906 SDn_2.n105 SDn_2.n104 0.96743
R4907 SDn_2.n116 SDn_2.n112 0.610728
R4908 SDn_2.n111 SDn_2.n91 0.564953
R4909 SDn_2.n119 SDn_2.n118 0.560976
R4910 SDn_2.n111 SDn_2.n110 0.141929
R4911 SDn_2.n123 SDn_2 0.140162
R4912 SDn_2.n120 SDn_2.n82 0.119429
R4913 SDn_2.n120 SDn_2.n119 0.0205
R4914 SDn_2.n118 SDn_2.n117 0.0171667
R4915 SDn_2.n124 SDn_2.n123 0.0135282
R4916 SDn_2.n112 SDn_2.n111 0.013514
R4917 SDn_2.n117 SDn_2.n116 0.0109989
R4918 SDn_2.n125 SDn_2.n120 0.00943873
R4919 SDn_2.n81 SDn_2.n80 0.0045
R4920 SDn_2 SDn_2.n125 0.00355856
R4921 SDn_2.n109 SDn_2.n107 0.0025
R4922 SD3_1.n97 SD3_1.n7 3.48971
R4923 SD3_1.n109 SD3_1.n3 3.48281
R4924 SD3_1.n56 SD3_1.n55 3.07792
R4925 SD3_1.n85 SD3_1.n27 3.07726
R4926 SD3_1.n88 SD3_1.n22 3.07632
R4927 SD3_1.n120 SD3_1.n117 3.07564
R4928 SD3_1.n76 SD3_1.n42 3.0732
R4929 SD3_1.n82 SD3_1.n32 3.07118
R4930 SD3_1.n79 SD3_1.n37 3.06982
R4931 SD3_1.n70 SD3_1.n44 3.06866
R4932 SD3_1.n91 SD3_1.n17 3.06533
R4933 SD3_1.n64 SD3_1.n49 3.06484
R4934 SD3_1 SD3_1.n1 3.06384
R4935 SD3_1.n58 SD3_1.n51 3.05987
R4936 SD3_1.n100 SD3_1.n5 3.05915
R4937 SD3_1.n94 SD3_1.n12 3.05307
R4938 SD3_1.n12 SD3_1.n11 2.90211
R4939 SD3_1.n102 SD3_1.n101 2.90208
R4940 SD3_1.n119 SD3_1.t30 2.7305
R4941 SD3_1.n119 SD3_1.n118 2.7305
R4942 SD3_1.n117 SD3_1.t53 2.7305
R4943 SD3_1.n117 SD3_1.n116 2.7305
R4944 SD3_1.n106 SD3_1.t21 2.7305
R4945 SD3_1.n106 SD3_1.n105 2.7305
R4946 SD3_1.n9 SD3_1.t36 2.7305
R4947 SD3_1.n9 SD3_1.n8 2.7305
R4948 SD3_1.n14 SD3_1.t48 2.7305
R4949 SD3_1.n14 SD3_1.n13 2.7305
R4950 SD3_1.n19 SD3_1.t18 2.7305
R4951 SD3_1.n19 SD3_1.n18 2.7305
R4952 SD3_1.n24 SD3_1.t60 2.7305
R4953 SD3_1.n24 SD3_1.n23 2.7305
R4954 SD3_1.n29 SD3_1.t10 2.7305
R4955 SD3_1.n29 SD3_1.n28 2.7305
R4956 SD3_1.n34 SD3_1.t62 2.7305
R4957 SD3_1.n34 SD3_1.n33 2.7305
R4958 SD3_1.n39 SD3_1.t19 2.7305
R4959 SD3_1.n39 SD3_1.n38 2.7305
R4960 SD3_1.n73 SD3_1.t0 2.7305
R4961 SD3_1.n73 SD3_1.n72 2.7305
R4962 SD3_1.n46 SD3_1.t14 2.7305
R4963 SD3_1.n46 SD3_1.n45 2.7305
R4964 SD3_1.n66 SD3_1.t46 2.7305
R4965 SD3_1.n66 SD3_1.n65 2.7305
R4966 SD3_1.n60 SD3_1.t9 2.7305
R4967 SD3_1.n60 SD3_1.n59 2.7305
R4968 SD3_1.n53 SD3_1.t3 2.7305
R4969 SD3_1.n53 SD3_1.n52 2.7305
R4970 SD3_1.n55 SD3_1.t23 2.7305
R4971 SD3_1.n55 SD3_1.n54 2.7305
R4972 SD3_1.n51 SD3_1.t2 2.7305
R4973 SD3_1.n51 SD3_1.n50 2.7305
R4974 SD3_1.n49 SD3_1.t34 2.7305
R4975 SD3_1.n49 SD3_1.n48 2.7305
R4976 SD3_1.n44 SD3_1.t44 2.7305
R4977 SD3_1.n44 SD3_1.n43 2.7305
R4978 SD3_1.n42 SD3_1.t26 2.7305
R4979 SD3_1.n42 SD3_1.n41 2.7305
R4980 SD3_1.n37 SD3_1.t61 2.7305
R4981 SD3_1.n37 SD3_1.n36 2.7305
R4982 SD3_1.n32 SD3_1.t38 2.7305
R4983 SD3_1.n32 SD3_1.n31 2.7305
R4984 SD3_1.n27 SD3_1.t59 2.7305
R4985 SD3_1.n27 SD3_1.n26 2.7305
R4986 SD3_1.n22 SD3_1.t28 2.7305
R4987 SD3_1.n22 SD3_1.n21 2.7305
R4988 SD3_1.n17 SD3_1.t63 2.7305
R4989 SD3_1.n17 SD3_1.n16 2.7305
R4990 SD3_1.n7 SD3_1.t54 2.7305
R4991 SD3_1.n7 SD3_1.n6 2.7305
R4992 SD3_1.n5 SD3_1.t17 2.7305
R4993 SD3_1.n5 SD3_1.n4 2.7305
R4994 SD3_1.n3 SD3_1.t8 2.7305
R4995 SD3_1.n3 SD3_1.n2 2.7305
R4996 SD3_1.n1 SD3_1.t31 2.7305
R4997 SD3_1.n1 SD3_1.n0 2.7305
R4998 SD3_1.n112 SD3_1.t55 2.7305
R4999 SD3_1.n112 SD3_1.n111 2.7305
R5000 SD3_1.n56 SD3_1.n53 2.5571
R5001 SD3_1.n120 SD3_1.n119 2.55706
R5002 SD3_1.n102 SD3_1.t51 2.40707
R5003 SD3_1.n12 SD3_1.t37 2.40704
R5004 SD3_1.n108 SD3_1.n107 2.24937
R5005 SD3_1.n104 SD3_1.n103 2.24505
R5006 SD3_1.n62 SD3_1.n61 2.24478
R5007 SD3_1.n68 SD3_1.n67 2.24478
R5008 SD3_1.n75 SD3_1.n74 1.49476
R5009 SD3_1.n87 SD3_1.n25 1.49463
R5010 SD3_1.n115 SD3_1.n114 1.49463
R5011 SD3_1.n81 SD3_1.n35 1.49463
R5012 SD3_1.n90 SD3_1.n20 1.49463
R5013 SD3_1.n69 SD3_1.n47 1.49439
R5014 SD3_1.n84 SD3_1.n30 1.49439
R5015 SD3_1.n78 SD3_1.n40 1.49439
R5016 SD3_1.n93 SD3_1.n15 1.49439
R5017 SD3_1.n96 SD3_1.n10 1.49439
R5018 SD3_1.n40 SD3_1.n39 1.43788
R5019 SD3_1.n74 SD3_1.n73 1.43788
R5020 SD3_1.n10 SD3_1.n9 1.43741
R5021 SD3_1.n25 SD3_1.n24 1.43741
R5022 SD3_1.n30 SD3_1.n29 1.43741
R5023 SD3_1.n47 SD3_1.n46 1.43741
R5024 SD3_1.n20 SD3_1.n19 1.43705
R5025 SD3_1.n107 SD3_1.n106 1.43694
R5026 SD3_1.n35 SD3_1.n34 1.43694
R5027 SD3_1.n67 SD3_1.n66 1.43694
R5028 SD3_1.n15 SD3_1.n14 1.43673
R5029 SD3_1.n61 SD3_1.n60 1.43673
R5030 SD3_1.n113 SD3_1.n112 1.42872
R5031 SD3_1.n103 SD3_1.n102 1.01023
R5032 SD3_1.n108 SD3_1.n104 0.593824
R5033 SD3_1.n57 SD3_1.n56 0.593282
R5034 SD3_1.n69 SD3_1.n68 0.586829
R5035 SD3_1.n99 SD3_1.n98 0.583544
R5036 SD3_1.n63 SD3_1.n62 0.581823
R5037 SD3_1.n78 SD3_1.n77 0.579925
R5038 SD3_1.n121 SD3_1.n120 0.577695
R5039 SD3_1.n93 SD3_1.n92 0.577272
R5040 SD3_1.n84 SD3_1.n83 0.576023
R5041 SD3_1.n90 SD3_1.n89 0.575664
R5042 SD3_1.n96 SD3_1.n95 0.575142
R5043 SD3_1.n81 SD3_1.n80 0.573011
R5044 SD3_1.n87 SD3_1.n86 0.572285
R5045 SD3_1.n115 SD3_1.n110 0.571741
R5046 SD3_1.n75 SD3_1.n71 0.569825
R5047 SD3_1.n113 SD3_1 0.0644679
R5048 SD3_1.n71 SD3_1.n70 0.0254398
R5049 SD3_1.n92 SD3_1.n91 0.0254398
R5050 SD3_1 SD3_1.n121 0.0243554
R5051 SD3_1.n80 SD3_1.n79 0.0232711
R5052 SD3_1.n98 SD3_1.n97 0.0232711
R5053 SD3_1.n110 SD3_1.n109 0.0232711
R5054 SD3_1.n88 SD3_1.n87 0.0218667
R5055 SD3_1.n86 SD3_1.n85 0.0211024
R5056 SD3_1.n95 SD3_1.n94 0.0211024
R5057 SD3_1.n82 SD3_1.n81 0.0200598
R5058 SD3_1.n77 SD3_1.n76 0.0200181
R5059 SD3_1.n76 SD3_1.n75 0.0190332
R5060 SD3_1.n83 SD3_1.n82 0.0189337
R5061 SD3_1.n85 SD3_1.n84 0.0186111
R5062 SD3_1.n94 SD3_1.n93 0.0178882
R5063 SD3_1.n89 SD3_1.n88 0.0178494
R5064 SD3_1.n58 SD3_1.n57 0.0166884
R5065 SD3_1.n68 SD3_1.n64 0.0166884
R5066 SD3_1.n79 SD3_1.n78 0.0157195
R5067 SD3_1.n97 SD3_1.n96 0.0157195
R5068 SD3_1.n62 SD3_1.n58 0.0156041
R5069 SD3_1.n64 SD3_1.n63 0.0156041
R5070 SD3_1.n104 SD3_1.n100 0.0150649
R5071 SD3_1 SD3_1.n115 0.0143027
R5072 SD3_1.n70 SD3_1.n69 0.0142737
R5073 SD3_1.n91 SD3_1.n90 0.0135538
R5074 SD3_1.n114 SD3_1.n113 0.00977503
R5075 SD3_1.n109 SD3_1.n108 0.00641934
R5076 SD3_1.n100 SD3_1.n99 0.00592169
R5077 b6.n8 b6.n7 64.4419
R5078 b6.n31 b6.n24 51.1109
R5079 b6.n25 b6.t44 50.6807
R5080 b6.n23 b6.n22 49.8352
R5081 b6.n35 b6.t24 47.9333
R5082 b6.n5 b6.t14 40.2611
R5083 b6.n0 b6.t37 39.8961
R5084 b6.n43 b6.n42 33.0652
R5085 b6.n44 b6.n43 31.6402
R5086 b6.n20 b6.n19 30.5682
R5087 b6.n4 b6.n3 26.0261
R5088 b6.n2 b6.n1 25.6611
R5089 b6.n11 b6.t6 24.8545
R5090 b6.n22 b6.t42 24.5042
R5091 b6.n7 b6.t2 23.0349
R5092 b6.t24 b6.t39 21.6159
R5093 b6.t10 b6.t26 21.5355
R5094 b6.t6 b6.t25 21.5355
R5095 b6.t40 b6.t11 21.5355
R5096 b6.t14 b6.t43 21.1705
R5097 b6.t37 b6.t18 21.1705
R5098 b6.t16 b6.t45 21.1705
R5099 b6.t36 b6.t17 21.1705
R5100 b6.n9 b6.t32 18.5039
R5101 b6.n36 b6.t19 14.6735
R5102 b6.n39 b6.t46 14.6735
R5103 b6.n43 b6.t10 14.6735
R5104 b6.n13 b6.t48 14.4545
R5105 b6.n16 b6.t30 14.4545
R5106 b6.n19 b6.t40 14.4545
R5107 b6.n22 b6.t23 14.3815
R5108 b6.n23 b6.t4 14.3815
R5109 b6.n24 b6.t29 14.3815
R5110 b6.n7 b6.t15 14.3085
R5111 b6.n8 b6.t12 14.3085
R5112 b6.n2 b6.t16 14.2355
R5113 b6.n3 b6.t36 14.2355
R5114 b6.n11 b6.t49 13.9435
R5115 b6.n12 b6.t27 13.9435
R5116 b6.n17 b6.t8 13.9435
R5117 b6.n18 b6.t35 13.9435
R5118 b6.n0 b6.t28 13.7975
R5119 b6.n1 b6.t41 13.7975
R5120 b6.n35 b6.t50 13.7245
R5121 b6.n42 b6.t31 13.7245
R5122 b6.n5 b6.t9 13.4325
R5123 b6.n4 b6.t38 13.4325
R5124 b6.n33 b6.t22 12.1915
R5125 b6.n34 b6.t3 12.1915
R5126 b6.n40 b6.t5 12.0455
R5127 b6.t31 b6.n41 12.0455
R5128 b6.n40 b6.t7 11.8265
R5129 b6.n41 b6.t33 11.8265
R5130 b6.n33 b6.t21 11.6805
R5131 b6.t50 b6.n34 11.6805
R5132 b6.n27 b6.t0 11.6029
R5133 b6.n1 b6.n0 11.5035
R5134 b6.n3 b6.n2 11.5035
R5135 b6.n36 b6.n35 11.1652
R5136 b6.n39 b6.n36 11.1652
R5137 b6.n42 b6.n39 11.1652
R5138 b6.t46 b6.n38 11.0965
R5139 b6.n14 b6.t20 10.8045
R5140 b6.n15 b6.t47 10.8045
R5141 b6.t30 b6.n15 10.7315
R5142 b6.n37 b6.t34 10.4395
R5143 b6.n38 b6.t13 10.4395
R5144 b6.n38 b6.n37 10.4005
R5145 b6.n12 b6.n11 10.4005
R5146 b6.n13 b6.n12 10.4005
R5147 b6.n16 b6.n13 10.4005
R5148 b6.n17 b6.n16 10.4005
R5149 b6.n18 b6.n17 10.4005
R5150 b6.n19 b6.n18 10.4005
R5151 b6.n24 b6.n23 10.1232
R5152 b6.n27 b6.t1 9.49371
R5153 b6.n15 b6.n14 8.93226
R5154 b6.n41 b6.n40 8.53084
R5155 b6.n34 b6.n33 7.66919
R5156 b6.n31 b6.n30 6.19053
R5157 b6.n6 b6.n5 5.28339
R5158 b6.n10 b6.n6 5.02841
R5159 b6.n9 b6.n8 4.53153
R5160 b6.n29 b6.n28 4.5305
R5161 b6.n10 b6.n9 3.85224
R5162 b6.n6 b6.n4 3.74655
R5163 b6.n28 b6.n27 3.63044
R5164 b6.n20 b6.n10 2.50672
R5165 b6.n29 b6.n26 2.2505
R5166 b6.n21 b6.n20 1.74245
R5167 b6.n46 b6.n45 1.50779
R5168 b6.n46 b6.n31 1.35684
R5169 b6.n28 b6 0.0263621
R5170 b6 b6.n21 0.0166901
R5171 b6 b6.n26 0.00567241
R5172 b6.n26 b6.n25 0.00360345
R5173 b6.n45 b6.n32 0.00355446
R5174 b6.n30 b6.n29 0.0035
R5175 b6.n45 b6.n44 0.00227316
R5176 b6 b6.n46 0.00137379
R5177 IT.n117 IT.n116 132.385
R5178 IT.n111 IT.n110 131.189
R5179 IT.n0 IT.t74 117.912
R5180 IT.n36 IT.t44 117.838
R5181 IT.n91 IT.n90 108.54
R5182 IT.n96 IT.n95 106.138
R5183 IT.n14 IT.n13 105.665
R5184 IT.n85 IT.n84 105.632
R5185 IT.n50 IT.n49 105.126
R5186 IT.n145 IT.n144 104.26
R5187 IT.n74 IT.n73 103.823
R5188 IT.n109 IT.n108 103.823
R5189 IT.n38 IT.n37 103.823
R5190 IT.n40 IT.n39 103.823
R5191 IT.n42 IT.n41 103.823
R5192 IT.n44 IT.n43 103.823
R5193 IT.n46 IT.n45 103.823
R5194 IT.n48 IT.n47 103.823
R5195 IT.n17 IT.n16 103.823
R5196 IT.n19 IT.n18 103.823
R5197 IT.n21 IT.n20 103.823
R5198 IT.n23 IT.n22 103.823
R5199 IT.n25 IT.n24 103.823
R5200 IT.n27 IT.n26 103.823
R5201 IT.n29 IT.n28 103.823
R5202 IT.n2 IT.n1 103.823
R5203 IT.n4 IT.n3 103.823
R5204 IT.n6 IT.n5 103.823
R5205 IT.n8 IT.n7 103.823
R5206 IT.n10 IT.n9 103.823
R5207 IT.n12 IT.n11 103.823
R5208 IT.n67 IT.n66 103.823
R5209 IT.n65 IT.n64 103.823
R5210 IT.n63 IT.n62 103.823
R5211 IT.n61 IT.n60 103.823
R5212 IT.n59 IT.n58 103.823
R5213 IT.n78 IT.n77 103.823
R5214 IT.n87 IT.n86 103.823
R5215 IT.n100 IT.n99 36.3254
R5216 IT.n108 IT.t73 34.7404
R5217 IT.n16 IT.t55 33.7914
R5218 IT.n89 IT.n87 33.2561
R5219 IT.n30 IT.n29 22.1542
R5220 IT.n79 IT.n78 22.0563
R5221 IT.n75 IT.n74 21.6519
R5222 IT.n110 IT.n109 21.0894
R5223 IT.n144 IT.n143 21.0894
R5224 IT.n37 IT.n36 21.0894
R5225 IT.n39 IT.n38 21.0894
R5226 IT.n41 IT.n40 21.0894
R5227 IT.n43 IT.n42 21.0894
R5228 IT.n45 IT.n44 21.0894
R5229 IT.n47 IT.n46 21.0894
R5230 IT.n49 IT.n48 21.0894
R5231 IT.n18 IT.n17 21.0894
R5232 IT.n20 IT.n19 21.0894
R5233 IT.n22 IT.n21 21.0894
R5234 IT.n24 IT.n23 21.0894
R5235 IT.n26 IT.n25 21.0894
R5236 IT.n28 IT.n27 21.0894
R5237 IT.n1 IT.n0 21.0894
R5238 IT.n3 IT.n2 21.0894
R5239 IT.n5 IT.n4 21.0894
R5240 IT.n7 IT.n6 21.0894
R5241 IT.n9 IT.n8 21.0894
R5242 IT.n11 IT.n10 21.0894
R5243 IT.n13 IT.n12 21.0894
R5244 IT.n68 IT.n67 21.0894
R5245 IT.n66 IT.n65 21.0894
R5246 IT.n64 IT.n63 21.0894
R5247 IT.n62 IT.n61 21.0894
R5248 IT.n60 IT.n59 21.0894
R5249 IT.n58 IT.n57 21.0894
R5250 IT.n77 IT.n76 21.0894
R5251 IT.n86 IT.n85 21.0894
R5252 IT.n0 IT.t106 14.0895
R5253 IT.n1 IT.t82 14.0895
R5254 IT.n2 IT.t37 14.0895
R5255 IT.n3 IT.t65 14.0895
R5256 IT.n4 IT.t97 14.0895
R5257 IT.n5 IT.t53 14.0895
R5258 IT.n6 IT.t94 14.0895
R5259 IT.n7 IT.t64 14.0895
R5260 IT.n8 IT.t28 14.0895
R5261 IT.n9 IT.t80 14.0895
R5262 IT.n10 IT.t52 14.0895
R5263 IT.n11 IT.t77 14.0895
R5264 IT.n12 IT.t48 14.0895
R5265 IT.n13 IT.t86 14.0895
R5266 IT.n36 IT.t68 14.0165
R5267 IT.n37 IT.t26 14.0165
R5268 IT.n38 IT.t27 14.0165
R5269 IT.n39 IT.t40 14.0165
R5270 IT.n40 IT.t33 14.0165
R5271 IT.n41 IT.t93 14.0165
R5272 IT.n42 IT.t78 14.0165
R5273 IT.n43 IT.t38 14.0165
R5274 IT.n44 IT.t41 14.0165
R5275 IT.n45 IT.t100 14.0165
R5276 IT.n46 IT.t25 14.0165
R5277 IT.n47 IT.t67 14.0165
R5278 IT.n48 IT.t50 14.0165
R5279 IT.n49 IT.t30 14.0165
R5280 IT.n67 IT.t88 14.0165
R5281 IT.n66 IT.t81 14.0165
R5282 IT.n65 IT.t45 14.0165
R5283 IT.n64 IT.t59 14.0165
R5284 IT.n63 IT.t79 14.0165
R5285 IT.n62 IT.t98 14.0165
R5286 IT.n61 IT.t34 14.0165
R5287 IT.n60 IT.t35 14.0165
R5288 IT.n59 IT.t76 14.0165
R5289 IT.n58 IT.t91 14.0165
R5290 IT.n57 IT.t31 14.0165
R5291 IT.n76 IT.t24 14.0165
R5292 IT.n77 IT.t66 14.0165
R5293 IT.n78 IT.t42 14.0165
R5294 IT.n144 IT.t89 13.7245
R5295 IT.n143 IT.t29 13.7245
R5296 IT.n99 IT.t105 13.7245
R5297 IT.n85 IT.t47 13.7245
R5298 IT.n86 IT.t62 13.7245
R5299 IT.n87 IT.t101 13.7245
R5300 IT.n74 IT.t58 13.6515
R5301 IT.n73 IT.t54 13.6515
R5302 IT.n116 IT.t51 13.6515
R5303 IT.n108 IT.t60 13.6515
R5304 IT.n109 IT.t43 13.6515
R5305 IT.n110 IT.t61 13.6515
R5306 IT.n145 IT.t70 13.2848
R5307 IT.n75 IT.t63 13.0378
R5308 IT.n16 IT.t83 12.7025
R5309 IT.n17 IT.t46 12.7025
R5310 IT.n18 IT.t95 12.7025
R5311 IT.n19 IT.t56 12.7025
R5312 IT.n20 IT.t84 12.7025
R5313 IT.n21 IT.t104 12.7025
R5314 IT.n22 IT.t75 12.7025
R5315 IT.n23 IT.t107 12.7025
R5316 IT.n24 IT.t32 12.7025
R5317 IT.n25 IT.t39 12.7025
R5318 IT.n26 IT.t87 12.7025
R5319 IT.n27 IT.t57 12.7025
R5320 IT.n28 IT.t85 12.7025
R5321 IT.n29 IT.t49 12.7025
R5322 IT.n118 IT.t14 12.6295
R5323 IT.n117 IT.t0 12.6295
R5324 IT.n91 IT.t12 12.5565
R5325 IT.n95 IT.t4 12.5565
R5326 IT.n112 IT.t8 12.3375
R5327 IT.n111 IT.t10 12.3375
R5328 IT.n96 IT.t2 12.1915
R5329 IT.n14 IT.t36 11.1683
R5330 IT.n84 IT.t103 10.8639
R5331 IT.n80 IT.t102 10.4542
R5332 IT.n56 IT.t69 10.4093
R5333 IT.n89 IT.n88 10.1427
R5334 IT.n72 IT.n35 9.76656
R5335 IT.n52 IT.t90 9.3445
R5336 IT.n15 IT.t96 8.94772
R5337 IT.n90 IT.t6 7.7385
R5338 IT.n94 IT.n93 7.45611
R5339 IT.n137 IT.n136 7.24501
R5340 IT.n90 IT.n89 6.3515
R5341 IT.n101 IT.t3 6.33405
R5342 IT.n84 IT.n83 6.07308
R5343 IT.n119 IT.n117 4.63315
R5344 IT.n104 IT.n100 4.5005
R5345 IT.n94 IT.n91 4.33237
R5346 IT.n34 IT.n14 4.33006
R5347 IT.n113 IT.n111 4.19412
R5348 IT.n119 IT.n118 4.03194
R5349 IT.n95 IT.n94 4.01149
R5350 IT.n113 IT.n112 3.88348
R5351 IT.n136 IT.n133 3.67213
R5352 IT.n127 IT.n75 3.64368
R5353 IT.n81 IT.n79 3.54502
R5354 IT.n81 IT.n80 3.51942
R5355 IT.n31 IT.n15 3.51248
R5356 IT.n31 IT.n30 3.50535
R5357 IT.n123 IT.n122 3.43549
R5358 IT.n114 IT.n107 3.41085
R5359 IT.n71 IT.n54 3.14528
R5360 IT.n133 IT.t19 3.03383
R5361 IT.n133 IT.n132 3.03383
R5362 IT.n135 IT.t20 3.03383
R5363 IT.n135 IT.n134 3.03383
R5364 IT.n131 IT.t18 3.03383
R5365 IT.n131 IT.n130 3.03383
R5366 IT.n129 IT.t17 3.03383
R5367 IT.n129 IT.n128 3.03383
R5368 IT.n54 IT.n53 2.88564
R5369 IT.n83 IT.n82 2.88451
R5370 IT.n33 IT.n32 2.88425
R5371 IT.n146 IT.n145 2.8819
R5372 IT.n137 IT.n131 2.82159
R5373 IT.n138 IT.n129 2.82159
R5374 IT.n136 IT.n135 2.81922
R5375 IT.n122 IT.t15 2.7305
R5376 IT.n122 IT.n121 2.7305
R5377 IT.n107 IT.t11 2.7305
R5378 IT.n107 IT.n106 2.7305
R5379 IT.n93 IT.t13 2.7305
R5380 IT.n93 IT.n92 2.7305
R5381 IT.n53 IT.n52 2.3365
R5382 IT.n71 IT.n70 2.25242
R5383 IT.n34 IT.n33 2.25102
R5384 IT.n124 IT.n123 2.24675
R5385 IT.n51 IT.n50 2.23635
R5386 IT.n70 IT.n69 2.12238
R5387 IT.n114 IT.n113 2.11998
R5388 IT.n69 IT.n68 2.1175
R5389 IT.n98 IT.n97 1.90845
R5390 IT.n139 IT.n138 1.44061
R5391 IT.n115 IT.n114 1.3863
R5392 IT.n120 IT.n119 1.32705
R5393 IT.n69 IT.n56 1.21129
R5394 IT.n105 IT.n104 1.13148
R5395 IT.n127 IT.n126 1.01644
R5396 IT.n147 IT.n141 0.927254
R5397 IT.n97 IT.n96 0.747091
R5398 IT.n100 IT.n98 0.581182
R5399 IT.n138 IT.n137 0.525071
R5400 IT.n140 IT.n139 0.400171
R5401 IT.n72 IT.n71 0.350424
R5402 IT.n140 IT.n72 0.31999
R5403 IT.n126 IT.n105 0.286359
R5404 IT.n126 IT.n125 0.166826
R5405 IT.n139 IT.n127 0.0964132
R5406 IT.n142 IT 0.0795
R5407 IT.n146 IT.n142 0.0275
R5408 IT.n102 IT.n101 0.0250455
R5409 IT.n123 IT.n120 0.0151731
R5410 IT.n141 IT.n140 0.0133571
R5411 IT.n125 IT.n124 0.00905634
R5412 IT.n70 IT.n55 0.00457413
R5413 IT.n33 IT.n31 0.0045
R5414 IT.n35 IT.n34 0.00399501
R5415 IT.n104 IT.n103 0.00356818
R5416 IT.n103 IT.n102 0.00356818
R5417 IT IT.n147 0.00340389
R5418 IT.n83 IT.n81 0.0025
R5419 IT.n147 IT.n146 0.00159453
R5420 IT.n54 IT.n51 0.0015
R5421 IT.n35 IT 0.00102252
R5422 IT.n124 IT.n115 0.000816901
R5423 OUT6 OUT6.n94 18.695
R5424 OUT6.n126 OUT6.t15 6.52669
R5425 OUT6.n141 OUT6.n95 6.10941
R5426 OUT6.n72 OUT6.n71 4.24612
R5427 OUT6.n50 OUT6.n49 4.22703
R5428 OUT6.n93 OUT6.n92 4.04138
R5429 OUT6.n28 OUT6.n1 3.99956
R5430 OUT6.n83 OUT6.n80 3.71646
R5431 OUT6.n16 OUT6.n13 3.70904
R5432 OUT6.n23 OUT6.n20 3.66108
R5433 OUT6.n39 OUT6.n36 3.66108
R5434 OUT6.n67 OUT6.n64 3.65144
R5435 OUT6.n55 OUT6.n52 3.65144
R5436 OUT6.n126 OUT6.n125 3.52028
R5437 OUT6.n128 OUT6.n121 3.52028
R5438 OUT6.n130 OUT6.n117 3.52028
R5439 OUT6.n132 OUT6.n113 3.52028
R5440 OUT6.n134 OUT6.n109 3.52028
R5441 OUT6.n136 OUT6.n105 3.52028
R5442 OUT6.n138 OUT6.n101 3.52028
R5443 OUT6.n140 OUT6.n97 3.52028
R5444 OUT6.n58 OUT6.n43 3.40302
R5445 OUT6.n75 OUT6.n60 3.40023
R5446 OUT6.n139 OUT6.n99 3.37941
R5447 OUT6.n137 OUT6.n103 3.37941
R5448 OUT6.n135 OUT6.n107 3.37941
R5449 OUT6.n133 OUT6.n111 3.37941
R5450 OUT6.n131 OUT6.n115 3.37941
R5451 OUT6.n129 OUT6.n119 3.37941
R5452 OUT6.n127 OUT6.n123 3.37941
R5453 OUT6.n85 OUT6.n76 3.32729
R5454 OUT6.n16 OUT6.n15 3.1505
R5455 OUT6.n17 OUT6.n11 3.1505
R5456 OUT6.n18 OUT6.n9 3.1505
R5457 OUT6.n23 OUT6.n22 3.1505
R5458 OUT6.n26 OUT6.n5 3.1505
R5459 OUT6.n25 OUT6.n7 3.1505
R5460 OUT6.n27 OUT6.n3 3.1505
R5461 OUT6.n39 OUT6.n38 3.1505
R5462 OUT6.n67 OUT6.n66 3.1505
R5463 OUT6.n72 OUT6.n69 3.1505
R5464 OUT6.n74 OUT6.n62 3.1505
R5465 OUT6.n50 OUT6.n47 3.1505
R5466 OUT6.n55 OUT6.n54 3.1505
R5467 OUT6.n57 OUT6.n45 3.1505
R5468 OUT6.n83 OUT6.n82 3.1505
R5469 OUT6.n84 OUT6.n78 3.1505
R5470 OUT6.n86 OUT6.n41 3.1505
R5471 OUT6.n89 OUT6.n32 3.1505
R5472 OUT6.n88 OUT6.n34 3.1505
R5473 OUT6.n90 OUT6.n30 3.1505
R5474 OUT6.n76 OUT6.n58 2.88513
R5475 OUT6.n94 OUT6.n93 2.83512
R5476 OUT6.n1 OUT6.t2 2.7305
R5477 OUT6.n1 OUT6.n0 2.7305
R5478 OUT6.n3 OUT6.t68 2.7305
R5479 OUT6.n3 OUT6.n2 2.7305
R5480 OUT6.n7 OUT6.t93 2.7305
R5481 OUT6.n7 OUT6.n6 2.7305
R5482 OUT6.n5 OUT6.t1 2.7305
R5483 OUT6.n5 OUT6.n4 2.7305
R5484 OUT6.n9 OUT6.t52 2.7305
R5485 OUT6.n9 OUT6.n8 2.7305
R5486 OUT6.n11 OUT6.t53 2.7305
R5487 OUT6.n11 OUT6.n10 2.7305
R5488 OUT6.n15 OUT6.t76 2.7305
R5489 OUT6.n15 OUT6.n14 2.7305
R5490 OUT6.n13 OUT6.t77 2.7305
R5491 OUT6.n13 OUT6.n12 2.7305
R5492 OUT6.n20 OUT6.t48 2.7305
R5493 OUT6.n20 OUT6.n19 2.7305
R5494 OUT6.n22 OUT6.t66 2.7305
R5495 OUT6.n22 OUT6.n21 2.7305
R5496 OUT6.n30 OUT6.t7 2.7305
R5497 OUT6.n30 OUT6.n29 2.7305
R5498 OUT6.n34 OUT6.t63 2.7305
R5499 OUT6.n34 OUT6.n33 2.7305
R5500 OUT6.n32 OUT6.t44 2.7305
R5501 OUT6.n32 OUT6.n31 2.7305
R5502 OUT6.n36 OUT6.t84 2.7305
R5503 OUT6.n36 OUT6.n35 2.7305
R5504 OUT6.n38 OUT6.t5 2.7305
R5505 OUT6.n38 OUT6.n37 2.7305
R5506 OUT6.n41 OUT6.t80 2.7305
R5507 OUT6.n41 OUT6.n40 2.7305
R5508 OUT6.n60 OUT6.t64 2.7305
R5509 OUT6.n60 OUT6.n59 2.7305
R5510 OUT6.n62 OUT6.t51 2.7305
R5511 OUT6.n62 OUT6.n61 2.7305
R5512 OUT6.n64 OUT6.t4 2.7305
R5513 OUT6.n64 OUT6.n63 2.7305
R5514 OUT6.n66 OUT6.t74 2.7305
R5515 OUT6.n66 OUT6.n65 2.7305
R5516 OUT6.n69 OUT6.t3 2.7305
R5517 OUT6.n69 OUT6.n68 2.7305
R5518 OUT6.n71 OUT6.t47 2.7305
R5519 OUT6.n71 OUT6.n70 2.7305
R5520 OUT6.n43 OUT6.t92 2.7305
R5521 OUT6.n43 OUT6.n42 2.7305
R5522 OUT6.n45 OUT6.t79 2.7305
R5523 OUT6.n45 OUT6.n44 2.7305
R5524 OUT6.n47 OUT6.t72 2.7305
R5525 OUT6.n47 OUT6.n46 2.7305
R5526 OUT6.n49 OUT6.t0 2.7305
R5527 OUT6.n49 OUT6.n48 2.7305
R5528 OUT6.n52 OUT6.t67 2.7305
R5529 OUT6.n52 OUT6.n51 2.7305
R5530 OUT6.n54 OUT6.t57 2.7305
R5531 OUT6.n54 OUT6.n53 2.7305
R5532 OUT6.n78 OUT6.t78 2.7305
R5533 OUT6.n78 OUT6.n77 2.7305
R5534 OUT6.n80 OUT6.t61 2.7305
R5535 OUT6.n80 OUT6.n79 2.7305
R5536 OUT6.n82 OUT6.t62 2.7305
R5537 OUT6.n82 OUT6.n81 2.7305
R5538 OUT6.n92 OUT6.t43 2.7305
R5539 OUT6.n92 OUT6.n91 2.7305
R5540 OUT6.n99 OUT6.t22 2.7305
R5541 OUT6.n99 OUT6.n98 2.7305
R5542 OUT6.n103 OUT6.t38 2.7305
R5543 OUT6.n103 OUT6.n102 2.7305
R5544 OUT6.n107 OUT6.t35 2.7305
R5545 OUT6.n107 OUT6.n106 2.7305
R5546 OUT6.n111 OUT6.t19 2.7305
R5547 OUT6.n111 OUT6.n110 2.7305
R5548 OUT6.n115 OUT6.t30 2.7305
R5549 OUT6.n115 OUT6.n114 2.7305
R5550 OUT6.n119 OUT6.t40 2.7305
R5551 OUT6.n119 OUT6.n118 2.7305
R5552 OUT6.n123 OUT6.t26 2.7305
R5553 OUT6.n123 OUT6.n122 2.7305
R5554 OUT6.n125 OUT6.t16 2.7305
R5555 OUT6.n125 OUT6.n124 2.7305
R5556 OUT6.n121 OUT6.t27 2.7305
R5557 OUT6.n121 OUT6.n120 2.7305
R5558 OUT6.n117 OUT6.t18 2.7305
R5559 OUT6.n117 OUT6.n116 2.7305
R5560 OUT6.n113 OUT6.t34 2.7305
R5561 OUT6.n113 OUT6.n112 2.7305
R5562 OUT6.n109 OUT6.t20 2.7305
R5563 OUT6.n109 OUT6.n108 2.7305
R5564 OUT6.n105 OUT6.t36 2.7305
R5565 OUT6.n105 OUT6.n104 2.7305
R5566 OUT6.n101 OUT6.t24 2.7305
R5567 OUT6.n101 OUT6.n100 2.7305
R5568 OUT6.n97 OUT6.t10 2.7305
R5569 OUT6.n97 OUT6.n96 2.7305
R5570 OUT6.n76 OUT6.n75 2.2505
R5571 OUT6.n94 OUT6.n28 2.2505
R5572 OUT6.n17 OUT6.n16 1.08037
R5573 OUT6.n84 OUT6.n83 1.06999
R5574 OUT6.n24 OUT6.n23 0.890115
R5575 OUT6.n56 OUT6.n55 0.87333
R5576 OUT6.n87 OUT6.n39 0.853769
R5577 OUT6.n73 OUT6.n67 0.827481
R5578 OUT6.n27 OUT6.n26 0.682695
R5579 OUT6.n90 OUT6.n89 0.681139
R5580 OUT6.n18 OUT6.n17 0.564306
R5581 OUT6.n26 OUT6.n25 0.511077
R5582 OUT6.n89 OUT6.n88 0.501443
R5583 OUT6.n73 OUT6.n72 0.438262
R5584 OUT6.n141 OUT6.n140 0.417773
R5585 OUT6.n140 OUT6.n139 0.417773
R5586 OUT6.n139 OUT6.n138 0.417773
R5587 OUT6.n138 OUT6.n137 0.417773
R5588 OUT6.n137 OUT6.n136 0.417773
R5589 OUT6.n136 OUT6.n135 0.417773
R5590 OUT6.n135 OUT6.n134 0.417773
R5591 OUT6.n134 OUT6.n133 0.417773
R5592 OUT6.n133 OUT6.n132 0.417773
R5593 OUT6.n132 OUT6.n131 0.417773
R5594 OUT6.n131 OUT6.n130 0.417773
R5595 OUT6.n130 OUT6.n129 0.417773
R5596 OUT6.n129 OUT6.n128 0.417773
R5597 OUT6.n128 OUT6.n127 0.417773
R5598 OUT6.n127 OUT6.n126 0.417773
R5599 OUT6.n87 OUT6.n86 0.416349
R5600 OUT6.n24 OUT6.n18 0.389629
R5601 OUT6.n56 OUT6.n50 0.380241
R5602 OUT6.n85 OUT6.n84 0.257226
R5603 OUT6.n86 OUT6.n85 0.253149
R5604 OUT6.n88 OUT6.n87 0.236538
R5605 OUT6.n74 OUT6.n73 0.220379
R5606 OUT6.n58 OUT6.n57 0.213967
R5607 OUT6.n75 OUT6.n74 0.208465
R5608 OUT6.n28 OUT6.n27 0.207865
R5609 OUT6.n25 OUT6.n24 0.185692
R5610 OUT6.n57 OUT6.n56 0.178802
R5611 OUT6.n93 OUT6.n90 0.164923
R5612 OUT6 OUT6.n141 0.133455
R5613 b6b.n0 b6b.t49 84.0965
R5614 b6b.n17 b6b.t4 74.5586
R5615 b6b.n2 b6b.n1 70.0805
R5616 b6b.n19 b6b.n18 61.2726
R5617 b6b.n7 b6b.t21 58.8447
R5618 b6b.n40 b6b.t47 54.2651
R5619 b6b.n23 b6b.t25 47.5922
R5620 b6b.n13 b6b.n12 45.3788
R5621 b6b.n46 b6b.n45 39.4461
R5622 b6b.n47 b6b.n46 37.6576
R5623 b6b.n31 b6b.n30 33.0652
R5624 b6b.n32 b6b.n31 32.8101
R5625 b6b.n12 b6b.n9 26.5717
R5626 b6b.t40 b6b.t38 23.9755
R5627 b6b.t25 b6b.t24 23.8715
R5628 b6b.n8 b6b.n7 23.854
R5629 b6b.n20 b6b.n19 22.5861
R5630 b6b b6b.t43 19.4018
R5631 b6b.n41 b6b.t34 14.8195
R5632 b6b.n42 b6b.t5 14.8195
R5633 b6b.n46 b6b.t13 14.8195
R5634 b6b.n24 b6b.t14 14.5275
R5635 b6b.n27 b6b.t33 14.5275
R5636 b6b.n31 b6b.t40 14.5275
R5637 b6b.n7 b6b.t11 14.0165
R5638 b6b.n12 b6b.t9 14.0165
R5639 b6b.n0 b6b.t29 14.0165
R5640 b6b.n1 b6b.t46 14.0165
R5641 b6b.n2 b6b.t28 14.0165
R5642 b6b.n8 b6b.t2 13.9428
R5643 b6b.n23 b6b.t17 13.5785
R5644 b6b.n30 b6b.t36 13.5785
R5645 b6b.n13 b6b.t50 13.4138
R5646 b6b.n9 b6b.n8 13.3558
R5647 b6b.n41 b6b.n40 13.3198
R5648 b6b.n42 b6b.n41 13.3198
R5649 b6b.n45 b6b.n42 13.3198
R5650 b6b.n40 b6b.t32 13.2865
R5651 b6b.n45 b6b.t3 13.2865
R5652 b6b.n17 b6b.t39 13.2865
R5653 b6b.n18 b6b.t10 13.2865
R5654 b6b.n19 b6b.t19 13.2865
R5655 b6b.n25 b6b.t12 12.7025
R5656 b6b.n26 b6b.t31 12.7025
R5657 b6b.n18 b6b.n17 12.4464
R5658 b6b.n43 b6b.t22 11.6075
R5659 b6b.t3 b6b.n44 11.6075
R5660 b6b.t33 b6b.n26 11.1695
R5661 b6b.n27 b6b.n24 11.1652
R5662 b6b.n24 b6b.n23 11.1652
R5663 b6b.n30 b6b.n27 11.1652
R5664 b6b.n38 b6b.t41 11.0235
R5665 b6b.n39 b6b.t16 11.0235
R5666 b6b.n5 b6b.t45 11.0235
R5667 b6b.t11 b6b.n6 11.0235
R5668 b6b.n10 b6b.t27 11.0235
R5669 b6b.t9 b6b.n11 11.0235
R5670 b6b.n21 b6b.t23 10.8775
R5671 b6b.n22 b6b.t48 10.8775
R5672 b6b.n28 b6b.t7 10.8045
R5673 b6b.t36 b6b.n29 10.8045
R5674 b6b.n28 b6b.t37 10.7315
R5675 b6b.n29 b6b.t18 10.7315
R5676 b6b.n21 b6b.t42 10.6585
R5677 b6b.t17 b6b.n22 10.6585
R5678 b6b.n38 b6b.t8 10.5125
R5679 b6b.t32 b6b.n39 10.5125
R5680 b6b.n44 b6b.n43 10.26
R5681 b6b.n5 b6b.t15 10.1475
R5682 b6b.n6 b6b.t30 10.1475
R5683 b6b.n10 b6b.t44 10.1475
R5684 b6b.n11 b6b.t26 10.1475
R5685 b6b.n6 b6b.n5 10.1232
R5686 b6b.n43 b6b.t6 9.9285
R5687 b6b.n44 b6b.t35 9.9285
R5688 b6b.n11 b6b.n10 9.73383
R5689 b6b.n36 b6b.n34 9.49418
R5690 b6b.n1 b6b.n0 9.4905
R5691 b6b.n29 b6b.n28 9.4905
R5692 b6b.n36 b6b.n35 9.40022
R5693 b6b.n39 b6b.n38 9.37334
R5694 b6b.n22 b6b.n21 9.0386
R5695 b6b.n26 b6b.n25 8.16394
R5696 b6b.n3 b6b.n2 7.52054
R5697 b6b.n9 b6b.t20 7.0085
R5698 b6b.n49 b6b.n48 4.53085
R5699 b6b.n37 b6b.n36 2.2505
R5700 b6b.n14 b6b.n13 2.13621
R5701 b6b.n33 b6b.n32 2.04965
R5702 b6b.n15 b6b.n14 1.5034
R5703 b6b.n32 b6b.n20 1.40687
R5704 b6b.n49 b6b.n37 1.33542
R5705 b6b.n47 b6b.n33 1.12144
R5706 b6b.n20 b6b.n16 1.00188
R5707 b6b b6b.n49 0.0343961
R5708 b6b.n15 b6b.n3 0.0197857
R5709 b6b.n16 b6b.n15 0.0191429
R5710 b6b b6b.n33 0.0120079
R5711 b6b.n14 b6b.n4 0.00265339
R5712 b6b.n48 b6b.n47 0.00259302
R5713 b6b.n37 b6b 0.00192857
R5714 b2.n0 b2.t3 49.5502
R5715 b2.n10 b2.n9 44.2287
R5716 b2.n9 b2.t2 22.1139
R5717 b2.n12 b2.n10 21.2987
R5718 b2.n6 b2.t6 19.8669
R5719 b2.n11 b2.t1 9.49371
R5720 b2.n11 b2.t0 9.3756
R5721 b2.n4 b2.t4 7.0085
R5722 b2.n10 b2.n8 4.66598
R5723 b2.n8 b2.n7 4.5005
R5724 b2.n12 b2.n11 2.53871
R5725 b2 b2.n0 2.25981
R5726 b2.n9 b2.t5 2.1905
R5727 b2 b2.n12 1.11809
R5728 b2.n5 b2.n4 0.8035
R5729 b2.n6 b2.n5 0.8035
R5730 b2.n7 b2.n6 0.2195
R5731 b2.n0 b2 0.14127
R5732 b2.n3 b2.n2 0.0340106
R5733 b2.n8 b2.n1 0.00371429
R5734 b2.n8 b2.n3 0.00145745
R5735 OUT2.n6 OUT2.n5 17.8839
R5736 OUT2 OUT2.t0 6.00764
R5737 OUT2.n7 OUT2.n0 5.8805
R5738 OUT2.n5 OUT2.n2 4.04862
R5739 OUT2.n7 OUT2.n6 3.51222
R5740 OUT2.n5 OUT2.n4 3.38961
R5741 OUT2.n2 OUT2.t5 2.7305
R5742 OUT2.n2 OUT2.n1 2.7305
R5743 OUT2.n4 OUT2.t2 2.7305
R5744 OUT2.n4 OUT2.n3 2.7305
R5745 OUT2.n6 OUT2 2.31942
R5746 OUT2 OUT2.n7 0.068
R5747 a_n2265_3941.n50 a_n2265_3941.t44 102.981
R5748 a_n2265_3941.n12 a_n2265_3941.t17 49.5689
R5749 a_n2265_3941.t44 a_n2265_3941.n49 49.5689
R5750 a_n2265_3941.n12 a_n2265_3941.t18 26.0719
R5751 a_n2265_3941.n13 a_n2265_3941.t15 26.0719
R5752 a_n2265_3941.n14 a_n2265_3941.t26 26.0719
R5753 a_n2265_3941.n15 a_n2265_3941.t28 26.0719
R5754 a_n2265_3941.n16 a_n2265_3941.t40 26.0719
R5755 a_n2265_3941.n17 a_n2265_3941.t42 26.0719
R5756 a_n2265_3941.n18 a_n2265_3941.t13 26.0719
R5757 a_n2265_3941.n19 a_n2265_3941.t22 26.0719
R5758 a_n2265_3941.n20 a_n2265_3941.t23 26.0719
R5759 a_n2265_3941.n21 a_n2265_3941.t34 26.0719
R5760 a_n2265_3941.n22 a_n2265_3941.t37 26.0719
R5761 a_n2265_3941.n23 a_n2265_3941.t48 26.0719
R5762 a_n2265_3941.n24 a_n2265_3941.t19 26.0719
R5763 a_n2265_3941.n25 a_n2265_3941.t14 26.0719
R5764 a_n2265_3941.n26 a_n2265_3941.t32 26.0719
R5765 a_n2265_3941.n27 a_n2265_3941.t30 26.0719
R5766 a_n2265_3941.n28 a_n2265_3941.t20 26.0719
R5767 a_n2265_3941.n29 a_n2265_3941.t49 26.0719
R5768 a_n2265_3941.n30 a_n2265_3941.t46 26.0719
R5769 a_n2265_3941.n31 a_n2265_3941.t35 26.0719
R5770 a_n2265_3941.n32 a_n2265_3941.t31 26.0719
R5771 a_n2265_3941.n33 a_n2265_3941.t21 26.0719
R5772 a_n2265_3941.n34 a_n2265_3941.t50 26.0719
R5773 a_n2265_3941.n35 a_n2265_3941.t47 26.0719
R5774 a_n2265_3941.n36 a_n2265_3941.t36 26.0719
R5775 a_n2265_3941.n37 a_n2265_3941.t33 26.0719
R5776 a_n2265_3941.n38 a_n2265_3941.t38 26.0719
R5777 a_n2265_3941.n39 a_n2265_3941.t25 26.0719
R5778 a_n2265_3941.n40 a_n2265_3941.t24 26.0719
R5779 a_n2265_3941.n41 a_n2265_3941.t12 26.0719
R5780 a_n2265_3941.n42 a_n2265_3941.t51 26.0719
R5781 a_n2265_3941.n43 a_n2265_3941.t39 26.0719
R5782 a_n2265_3941.n44 a_n2265_3941.t43 26.0719
R5783 a_n2265_3941.n45 a_n2265_3941.t41 26.0719
R5784 a_n2265_3941.n46 a_n2265_3941.t29 26.0719
R5785 a_n2265_3941.n47 a_n2265_3941.t27 26.0719
R5786 a_n2265_3941.n48 a_n2265_3941.t16 26.0719
R5787 a_n2265_3941.n49 a_n2265_3941.t45 26.0719
R5788 a_n2265_3941.n13 a_n2265_3941.n12 19.6341
R5789 a_n2265_3941.n14 a_n2265_3941.n13 19.6341
R5790 a_n2265_3941.n15 a_n2265_3941.n14 19.6341
R5791 a_n2265_3941.n16 a_n2265_3941.n15 19.6341
R5792 a_n2265_3941.n17 a_n2265_3941.n16 19.6341
R5793 a_n2265_3941.n18 a_n2265_3941.n17 19.6341
R5794 a_n2265_3941.n19 a_n2265_3941.n18 19.6341
R5795 a_n2265_3941.n20 a_n2265_3941.n19 19.6341
R5796 a_n2265_3941.n21 a_n2265_3941.n20 19.6341
R5797 a_n2265_3941.n22 a_n2265_3941.n21 19.6341
R5798 a_n2265_3941.n23 a_n2265_3941.n22 19.6341
R5799 a_n2265_3941.n24 a_n2265_3941.n23 19.6341
R5800 a_n2265_3941.n25 a_n2265_3941.n24 19.6341
R5801 a_n2265_3941.n26 a_n2265_3941.n25 19.6341
R5802 a_n2265_3941.n27 a_n2265_3941.n26 19.6341
R5803 a_n2265_3941.n28 a_n2265_3941.n27 19.6341
R5804 a_n2265_3941.n29 a_n2265_3941.n28 19.6341
R5805 a_n2265_3941.n30 a_n2265_3941.n29 19.6341
R5806 a_n2265_3941.n31 a_n2265_3941.n30 19.6341
R5807 a_n2265_3941.n32 a_n2265_3941.n31 19.6341
R5808 a_n2265_3941.n33 a_n2265_3941.n32 19.6341
R5809 a_n2265_3941.n34 a_n2265_3941.n33 19.6341
R5810 a_n2265_3941.n35 a_n2265_3941.n34 19.6341
R5811 a_n2265_3941.n36 a_n2265_3941.n35 19.6341
R5812 a_n2265_3941.n37 a_n2265_3941.n36 19.6341
R5813 a_n2265_3941.n38 a_n2265_3941.n37 19.6341
R5814 a_n2265_3941.n39 a_n2265_3941.n38 19.6341
R5815 a_n2265_3941.n40 a_n2265_3941.n39 19.6341
R5816 a_n2265_3941.n41 a_n2265_3941.n40 19.6341
R5817 a_n2265_3941.n42 a_n2265_3941.n41 19.6341
R5818 a_n2265_3941.n43 a_n2265_3941.n42 19.6341
R5819 a_n2265_3941.n44 a_n2265_3941.n43 19.6341
R5820 a_n2265_3941.n45 a_n2265_3941.n44 19.6341
R5821 a_n2265_3941.n46 a_n2265_3941.n45 19.6341
R5822 a_n2265_3941.n47 a_n2265_3941.n46 19.6341
R5823 a_n2265_3941.n48 a_n2265_3941.n47 19.6341
R5824 a_n2265_3941.n49 a_n2265_3941.n48 19.6341
R5825 a_n2265_3941.n10 a_n2265_3941.n7 3.7805
R5826 a_n2265_3941.n11 a_n2265_3941.n3 3.7805
R5827 a_n2265_3941.n10 a_n2265_3941.n9 3.7255
R5828 a_n2265_3941.n51 a_n2265_3941.n50 3.13775
R5829 a_n2265_3941.n10 a_n2265_3941.n5 3.09941
R5830 a_n2265_3941.n11 a_n2265_3941.n1 3.09941
R5831 a_n2265_3941.n9 a_n2265_3941.t6 0.9105
R5832 a_n2265_3941.n9 a_n2265_3941.n8 0.9105
R5833 a_n2265_3941.n5 a_n2265_3941.t3 0.9105
R5834 a_n2265_3941.n5 a_n2265_3941.n4 0.9105
R5835 a_n2265_3941.n1 a_n2265_3941.t4 0.9105
R5836 a_n2265_3941.n1 a_n2265_3941.n0 0.9105
R5837 a_n2265_3941.n51 a_n2265_3941.t0 0.9105
R5838 a_n2265_3941.n52 a_n2265_3941.n51 0.9105
R5839 a_n2265_3941.n7 a_n2265_3941.t9 0.8195
R5840 a_n2265_3941.n7 a_n2265_3941.n6 0.8195
R5841 a_n2265_3941.n3 a_n2265_3941.t10 0.8195
R5842 a_n2265_3941.n3 a_n2265_3941.n2 0.8195
R5843 a_n2265_3941.n11 a_n2265_3941.n10 0.626587
R5844 a_n2265_3941.n50 a_n2265_3941.n11 0.565935
R5845 b5b.t24 b5b.n11 75.0723
R5846 b5b.n10 b5b.t23 72.0525
R5847 b5b.n13 b5b.t21 62.2995
R5848 b5b.n14 b5b.n12 47.9184
R5849 b5b.n7 b5b.t8 47.5922
R5850 b5b.n18 b5b.n17 36.7152
R5851 b5b.n12 b5b.t13 24.4555
R5852 b5b.t13 b5b.t24 21.0034
R5853 b5b.t22 b5b.t11 20.7325
R5854 b5b.t14 b5b.t3 20.7325
R5855 b5b.t23 b5b.t12 20.7325
R5856 b5b.n19 b5b.t15 19.1982
R5857 b5b.n11 b5b.n10 14.8925
R5858 b5b.n8 b5b.t18 14.5275
R5859 b5b.n19 b5b.n18 14.5057
R5860 b5b.n13 b5b.t5 14.3815
R5861 b5b.n12 b5b.t10 14.3815
R5862 b5b.n14 b5b.t2 14.3815
R5863 b5b.n15 b5b.t16 14.2355
R5864 b5b.n7 b5b.t19 13.5785
R5865 b5b.n17 b5b.t7 13.5785
R5866 b5b.n11 b5b.t22 11.6075
R5867 b5b.n10 b5b.t14 11.6075
R5868 b5b.n8 b5b.n7 11.1652
R5869 b5b.n17 b5b.n16 11.1652
R5870 b5b.n16 b5b.n8 11.1652
R5871 b5b.n3 b5b.t20 11.0235
R5872 b5b.n4 b5b.t4 11.0235
R5873 b5b.n5 b5b.t9 10.9505
R5874 b5b.t19 b5b.n6 10.9505
R5875 b5b.n5 b5b.t6 10.5855
R5876 b5b.n6 b5b.t17 10.5855
R5877 b5b.n3 b5b.t26 10.5125
R5878 b5b.t7 b5b.n4 10.5125
R5879 b5b.n14 b5b.n13 9.73383
R5880 b5b.n18 b5b.t25 9.7095
R5881 b5b.n2 b5b.n0 9.49418
R5882 b5b.n2 b5b.n1 9.40022
R5883 b5b.n6 b5b.n5 9.37334
R5884 b5b.n4 b5b.n3 9.14749
R5885 b5b b5b.n14 6.02162
R5886 b5b.n15 b5b 4.0055
R5887 b5b b5b.n2 2.25319
R5888 b5b.n16 b5b.n15 0.2925
R5889 b5b b5b.n19 0.224828
R5890 b5b.n16 b5b.n9 0.0735
R5891 OUT5.n65 OUT5.n64 11.1462
R5892 OUT5 OUT5.n46 9.06769
R5893 OUT5.n57 OUT5.n56 6.90515
R5894 OUT5.n62 OUT5.t7 6.48993
R5895 OUT5.n65 OUT5.t5 6.12071
R5896 OUT5.n69 OUT5.n47 6.11137
R5897 OUT5.n42 OUT5.n41 3.88773
R5898 OUT5.n8 OUT5.n7 3.88773
R5899 OUT5.n19 OUT5.n18 3.88773
R5900 OUT5.n31 OUT5.n30 3.80786
R5901 OUT5.n57 OUT5.n55 3.54767
R5902 OUT5.n62 OUT5.n61 3.46159
R5903 OUT5.n66 OUT5.n53 3.46159
R5904 OUT5.n68 OUT5.n49 3.46159
R5905 OUT5.n63 OUT5.n59 3.38137
R5906 OUT5.n67 OUT5.n51 3.38137
R5907 OUT5.n42 OUT5.n39 3.1505
R5908 OUT5.n43 OUT5.n37 3.1505
R5909 OUT5.n44 OUT5.n35 3.1505
R5910 OUT5.n31 OUT5.n28 3.1505
R5911 OUT5.n32 OUT5.n26 3.1505
R5912 OUT5.n33 OUT5.n24 3.1505
R5913 OUT5.n8 OUT5.n5 3.1505
R5914 OUT5.n9 OUT5.n3 3.1505
R5915 OUT5.n10 OUT5.n1 3.1505
R5916 OUT5.n20 OUT5.n14 3.1505
R5917 OUT5.n19 OUT5.n16 3.1505
R5918 OUT5.n21 OUT5.n12 3.1505
R5919 OUT5.n46 OUT5.n22 3.00524
R5920 OUT5.n59 OUT5.t12 2.7305
R5921 OUT5.n59 OUT5.n58 2.7305
R5922 OUT5.n61 OUT5.t8 2.7305
R5923 OUT5.n61 OUT5.n60 2.7305
R5924 OUT5.n55 OUT5.t9 2.7305
R5925 OUT5.n55 OUT5.n54 2.7305
R5926 OUT5.n35 OUT5.t22 2.7305
R5927 OUT5.n35 OUT5.n34 2.7305
R5928 OUT5.n37 OUT5.t35 2.7305
R5929 OUT5.n37 OUT5.n36 2.7305
R5930 OUT5.n39 OUT5.t32 2.7305
R5931 OUT5.n39 OUT5.n38 2.7305
R5932 OUT5.n41 OUT5.t2 2.7305
R5933 OUT5.n41 OUT5.n40 2.7305
R5934 OUT5.n24 OUT5.t47 2.7305
R5935 OUT5.n24 OUT5.n23 2.7305
R5936 OUT5.n26 OUT5.t25 2.7305
R5937 OUT5.n26 OUT5.n25 2.7305
R5938 OUT5.n28 OUT5.t31 2.7305
R5939 OUT5.n28 OUT5.n27 2.7305
R5940 OUT5.n30 OUT5.t39 2.7305
R5941 OUT5.n30 OUT5.n29 2.7305
R5942 OUT5.n1 OUT5.t34 2.7305
R5943 OUT5.n1 OUT5.n0 2.7305
R5944 OUT5.n3 OUT5.t19 2.7305
R5945 OUT5.n3 OUT5.n2 2.7305
R5946 OUT5.n5 OUT5.t20 2.7305
R5947 OUT5.n5 OUT5.n4 2.7305
R5948 OUT5.n7 OUT5.t42 2.7305
R5949 OUT5.n7 OUT5.n6 2.7305
R5950 OUT5.n12 OUT5.t26 2.7305
R5951 OUT5.n12 OUT5.n11 2.7305
R5952 OUT5.n18 OUT5.t28 2.7305
R5953 OUT5.n18 OUT5.n17 2.7305
R5954 OUT5.n16 OUT5.t36 2.7305
R5955 OUT5.n16 OUT5.n15 2.7305
R5956 OUT5.n14 OUT5.t38 2.7305
R5957 OUT5.n14 OUT5.n13 2.7305
R5958 OUT5.n51 OUT5.t10 2.7305
R5959 OUT5.n51 OUT5.n50 2.7305
R5960 OUT5.n53 OUT5.t11 2.7305
R5961 OUT5.n53 OUT5.n52 2.7305
R5962 OUT5.n49 OUT5.t6 2.7305
R5963 OUT5.n49 OUT5.n48 2.7305
R5964 OUT5.n46 OUT5.n45 2.2555
R5965 OUT5.n22 OUT5.n10 0.916077
R5966 OUT5.n44 OUT5.n43 0.826683
R5967 OUT5.n33 OUT5.n32 0.74308
R5968 OUT5.n21 OUT5.n20 0.73453
R5969 OUT5.n10 OUT5.n9 0.733978
R5970 OUT5.n45 OUT5.n44 0.698412
R5971 OUT5.n43 OUT5.n42 0.565394
R5972 OUT5.n32 OUT5.n31 0.565394
R5973 OUT5.n9 OUT5.n8 0.565394
R5974 OUT5.n20 OUT5.n19 0.565394
R5975 OUT5.n64 OUT5.n63 0.379057
R5976 OUT5.n63 OUT5.n62 0.379057
R5977 OUT5.n69 OUT5.n68 0.379057
R5978 OUT5.n68 OUT5.n67 0.379057
R5979 OUT5.n67 OUT5.n66 0.379057
R5980 OUT5.n45 OUT5.n33 0.376378
R5981 OUT5.n66 OUT5.n65 0.370706
R5982 OUT5.n22 OUT5.n21 0.304973
R5983 OUT5 OUT5.n69 0.136892
R5984 OUT5.n64 OUT5.n57 0.00235567
R5985 Gc_1.n160 Gc_1.n48 31.7026
R5986 Gc_1.n194 Gc_1.n193 28.879
R5987 Gc_1.n192 Gc_1.t139 24.4555
R5988 Gc_1.n191 Gc_1.t141 24.4555
R5989 Gc_1.n188 Gc_1.t136 24.4555
R5990 Gc_1.n187 Gc_1.t138 24.4555
R5991 Gc_1.n184 Gc_1.t108 24.4555
R5992 Gc_1.n183 Gc_1.t96 24.4555
R5993 Gc_1.n180 Gc_1.t127 24.4555
R5994 Gc_1.n179 Gc_1.t104 24.4555
R5995 Gc_1.n34 Gc_1.t123 24.4555
R5996 Gc_1.n35 Gc_1.t133 24.4555
R5997 Gc_1.n38 Gc_1.t109 24.4555
R5998 Gc_1.n39 Gc_1.t107 24.4555
R5999 Gc_1.n42 Gc_1.t114 24.4555
R6000 Gc_1.n43 Gc_1.t112 24.4555
R6001 Gc_1.n46 Gc_1.t97 24.4555
R6002 Gc_1.n47 Gc_1.t118 24.4555
R6003 Gc_1.n104 Gc_1.t86 23.86
R6004 Gc_1.n149 Gc_1.t40 23.86
R6005 Gc_1.n104 Gc_1.t46 23.1415
R6006 Gc_1.n105 Gc_1.t88 23.1415
R6007 Gc_1.n149 Gc_1.t74 23.1415
R6008 Gc_1.n150 Gc_1.t60 23.1415
R6009 Gc_1.n152 Gc_1.t70 23.1415
R6010 Gc_1.n56 Gc_1.t34 23.1415
R6011 Gc_1.n58 Gc_1.t94 23.1415
R6012 Gc_1.n67 Gc_1.t58 23.1415
R6013 Gc_1.n69 Gc_1.t66 23.1415
R6014 Gc_1.n78 Gc_1.t54 23.1415
R6015 Gc_1.n80 Gc_1.t64 23.1415
R6016 Gc_1.n89 Gc_1.t48 23.1415
R6017 Gc_1.n91 Gc_1.t92 23.1415
R6018 Gc_1.n121 Gc_1.t56 23.1415
R6019 Gc_1.n123 Gc_1.t84 23.1415
R6020 Gc_1.n102 Gc_1.t44 23.1415
R6021 Gc_1.n106 Gc_1.t50 13.8705
R6022 Gc_1.n151 Gc_1.t80 13.8705
R6023 Gc_1.n153 Gc_1.t32 13.8705
R6024 Gc_1.n57 Gc_1.t78 13.8705
R6025 Gc_1.n59 Gc_1.t38 13.8705
R6026 Gc_1.n68 Gc_1.t82 13.8705
R6027 Gc_1.n70 Gc_1.t36 13.8705
R6028 Gc_1.n79 Gc_1.t72 13.8705
R6029 Gc_1.n81 Gc_1.t42 13.8705
R6030 Gc_1.n90 Gc_1.t76 13.8705
R6031 Gc_1.n92 Gc_1.t62 13.8705
R6032 Gc_1.n122 Gc_1.t68 13.8705
R6033 Gc_1.n124 Gc_1.t52 13.8705
R6034 Gc_1.n103 Gc_1.t90 13.8705
R6035 Gc_1.n193 Gc_1.t125 13.7245
R6036 Gc_1.n190 Gc_1.t142 13.7245
R6037 Gc_1.n189 Gc_1.t120 13.7245
R6038 Gc_1.n186 Gc_1.t132 13.7245
R6039 Gc_1.n185 Gc_1.t99 13.7245
R6040 Gc_1.n182 Gc_1.t124 13.7245
R6041 Gc_1.n181 Gc_1.t137 13.7245
R6042 Gc_1.n178 Gc_1.t110 13.7245
R6043 Gc_1.n33 Gc_1.t143 13.7245
R6044 Gc_1.n36 Gc_1.t119 13.7245
R6045 Gc_1.n37 Gc_1.t129 13.7245
R6046 Gc_1.n40 Gc_1.t116 13.7245
R6047 Gc_1.n41 Gc_1.t135 13.7245
R6048 Gc_1.n44 Gc_1.t121 13.7245
R6049 Gc_1.n45 Gc_1.t134 13.7245
R6050 Gc_1.n48 Gc_1.t113 13.7245
R6051 Gc_1.n193 Gc_1.n192 10.6935
R6052 Gc_1.n192 Gc_1.n191 10.6935
R6053 Gc_1.n191 Gc_1.n190 10.6935
R6054 Gc_1.n190 Gc_1.n189 10.6935
R6055 Gc_1.n189 Gc_1.n188 10.6935
R6056 Gc_1.n188 Gc_1.n187 10.6935
R6057 Gc_1.n187 Gc_1.n186 10.6935
R6058 Gc_1.n186 Gc_1.n185 10.6935
R6059 Gc_1.n185 Gc_1.n184 10.6935
R6060 Gc_1.n184 Gc_1.n183 10.6935
R6061 Gc_1.n183 Gc_1.n182 10.6935
R6062 Gc_1.n182 Gc_1.n181 10.6935
R6063 Gc_1.n181 Gc_1.n180 10.6935
R6064 Gc_1.n180 Gc_1.n179 10.6935
R6065 Gc_1.n179 Gc_1.n178 10.6935
R6066 Gc_1.n34 Gc_1.n33 10.6935
R6067 Gc_1.n35 Gc_1.n34 10.6935
R6068 Gc_1.n36 Gc_1.n35 10.6935
R6069 Gc_1.n37 Gc_1.n36 10.6935
R6070 Gc_1.n38 Gc_1.n37 10.6935
R6071 Gc_1.n39 Gc_1.n38 10.6935
R6072 Gc_1.n40 Gc_1.n39 10.6935
R6073 Gc_1.n41 Gc_1.n40 10.6935
R6074 Gc_1.n42 Gc_1.n41 10.6935
R6075 Gc_1.n43 Gc_1.n42 10.6935
R6076 Gc_1.n44 Gc_1.n43 10.6935
R6077 Gc_1.n45 Gc_1.n44 10.6935
R6078 Gc_1.n46 Gc_1.n45 10.6935
R6079 Gc_1.n47 Gc_1.n46 10.6935
R6080 Gc_1.n48 Gc_1.n47 10.6935
R6081 Gc_1.n105 Gc_1.n104 9.98997
R6082 Gc_1.n106 Gc_1.n105 9.98997
R6083 Gc_1.n150 Gc_1.n149 9.98997
R6084 Gc_1.n151 Gc_1.n150 9.98997
R6085 Gc_1.n153 Gc_1.n152 9.98997
R6086 Gc_1.n57 Gc_1.n56 9.98997
R6087 Gc_1.n59 Gc_1.n58 9.98997
R6088 Gc_1.n68 Gc_1.n67 9.98997
R6089 Gc_1.n70 Gc_1.n69 9.98997
R6090 Gc_1.n79 Gc_1.n78 9.98997
R6091 Gc_1.n81 Gc_1.n80 9.98997
R6092 Gc_1.n90 Gc_1.n89 9.98997
R6093 Gc_1.n92 Gc_1.n91 9.98997
R6094 Gc_1.n122 Gc_1.n121 9.98997
R6095 Gc_1.n124 Gc_1.n123 9.98997
R6096 Gc_1.n103 Gc_1.n102 9.98997
R6097 Gc_1.n154 Gc_1.n151 6.72418
R6098 Gc_1.n177 Gc_1.t29 6.14854
R6099 Gc_1.n161 Gc_1.n32 6.14854
R6100 Gc_1.n60 Gc_1.n57 5.85971
R6101 Gc_1.n125 Gc_1.n122 5.85971
R6102 Gc_1.n82 Gc_1.n79 5.37945
R6103 Gc_1.n71 Gc_1.n70 5.18734
R6104 Gc_1.n93 Gc_1.n90 5.18734
R6105 Gc_1.n107 Gc_1.n106 5.18734
R6106 Gc_1.n71 Gc_1.n68 4.80313
R6107 Gc_1.n93 Gc_1.n92 4.80313
R6108 Gc_1.n107 Gc_1.n103 4.80313
R6109 Gc_1.n82 Gc_1.n81 4.61103
R6110 Gc_1.n159 Gc_1.n49 4.29033
R6111 Gc_1.n60 Gc_1.n59 4.13076
R6112 Gc_1.n125 Gc_1.n124 4.13076
R6113 Gc_1.n162 Gc_1.n31 3.44202
R6114 Gc_1.n164 Gc_1.n27 3.44202
R6115 Gc_1.n166 Gc_1.n23 3.44202
R6116 Gc_1.n168 Gc_1.n19 3.44202
R6117 Gc_1.n170 Gc_1.n15 3.44202
R6118 Gc_1.n172 Gc_1.n11 3.44202
R6119 Gc_1.n174 Gc_1.n7 3.44202
R6120 Gc_1.n176 Gc_1.n3 3.44202
R6121 Gc_1.n175 Gc_1.n5 3.41854
R6122 Gc_1.n173 Gc_1.n9 3.41854
R6123 Gc_1.n171 Gc_1.n13 3.41854
R6124 Gc_1.n169 Gc_1.n17 3.41854
R6125 Gc_1.n167 Gc_1.n21 3.41854
R6126 Gc_1.n165 Gc_1.n25 3.41854
R6127 Gc_1.n163 Gc_1.n29 3.41854
R6128 Gc_1.n154 Gc_1.n153 3.26629
R6129 Gc_1.n119 Gc_1.t69 3.03383
R6130 Gc_1.n119 Gc_1.n118 3.03383
R6131 Gc_1.n88 Gc_1.t77 3.03383
R6132 Gc_1.n88 Gc_1.n87 3.03383
R6133 Gc_1.n77 Gc_1.t73 3.03383
R6134 Gc_1.n77 Gc_1.n76 3.03383
R6135 Gc_1.n66 Gc_1.t83 3.03383
R6136 Gc_1.n66 Gc_1.n65 3.03383
R6137 Gc_1.n55 Gc_1.t79 3.03383
R6138 Gc_1.n55 Gc_1.n54 3.03383
R6139 Gc_1.n147 Gc_1.t81 3.03383
R6140 Gc_1.n147 Gc_1.n146 3.03383
R6141 Gc_1.n101 Gc_1.t91 3.03383
R6142 Gc_1.n101 Gc_1.n100 3.03383
R6143 Gc_1.n1 Gc_1.t87 3.03383
R6144 Gc_1.n111 Gc_1.t89 3.03383
R6145 Gc_1.n111 Gc_1.n110 3.03383
R6146 Gc_1.n99 Gc_1.t85 3.03383
R6147 Gc_1.n99 Gc_1.n98 3.03383
R6148 Gc_1.n97 Gc_1.t93 3.03383
R6149 Gc_1.n97 Gc_1.n96 3.03383
R6150 Gc_1.n86 Gc_1.t65 3.03383
R6151 Gc_1.n86 Gc_1.n85 3.03383
R6152 Gc_1.n75 Gc_1.t67 3.03383
R6153 Gc_1.n75 Gc_1.n74 3.03383
R6154 Gc_1.n64 Gc_1.t95 3.03383
R6155 Gc_1.n64 Gc_1.n63 3.03383
R6156 Gc_1.n53 Gc_1.t71 3.03383
R6157 Gc_1.n53 Gc_1.n52 3.03383
R6158 Gc_1.n51 Gc_1.t75 3.03383
R6159 Gc_1.n51 Gc_1.n50 3.03383
R6160 Gc_1.n73 Gc_1.n66 2.92153
R6161 Gc_1.n95 Gc_1.n88 2.91939
R6162 Gc_1.n62 Gc_1.n55 2.91939
R6163 Gc_1.n84 Gc_1.n77 2.91724
R6164 Gc_1.n109 Gc_1.n101 2.91616
R6165 Gc_1.n120 Gc_1.n119 2.88224
R6166 Gc_1.n155 Gc_1.n154 2.8805
R6167 Gc_1.n61 Gc_1.n60 2.8805
R6168 Gc_1.n72 Gc_1.n71 2.8805
R6169 Gc_1.n83 Gc_1.n82 2.8805
R6170 Gc_1.n94 Gc_1.n93 2.8805
R6171 Gc_1.n126 Gc_1.n125 2.8805
R6172 Gc_1.n108 Gc_1.n107 2.8805
R6173 Gc_1.n148 Gc_1.n147 2.87637
R6174 Gc_1.n117 Gc_1.n99 2.79692
R6175 Gc_1.n133 Gc_1.n86 2.79126
R6176 Gc_1.n158 Gc_1.n51 2.7872
R6177 Gc_1.n141 Gc_1.n64 2.78604
R6178 Gc_1.n113 Gc_1.n111 2.78592
R6179 Gc_1.n145 Gc_1.n53 2.78535
R6180 Gc_1.n129 Gc_1.n97 2.78113
R6181 Gc_1.n137 Gc_1.n75 2.78104
R6182 Gc_1.n31 Gc_1.t22 2.7305
R6183 Gc_1.n31 Gc_1.n30 2.7305
R6184 Gc_1.n27 Gc_1.t26 2.7305
R6185 Gc_1.n27 Gc_1.n26 2.7305
R6186 Gc_1.n23 Gc_1.t21 2.7305
R6187 Gc_1.n23 Gc_1.n22 2.7305
R6188 Gc_1.n19 Gc_1.t17 2.7305
R6189 Gc_1.n19 Gc_1.n18 2.7305
R6190 Gc_1.n15 Gc_1.t15 2.7305
R6191 Gc_1.n15 Gc_1.n14 2.7305
R6192 Gc_1.n11 Gc_1.t27 2.7305
R6193 Gc_1.n11 Gc_1.n10 2.7305
R6194 Gc_1.n7 Gc_1.t20 2.7305
R6195 Gc_1.n7 Gc_1.n6 2.7305
R6196 Gc_1.n3 Gc_1.t24 2.7305
R6197 Gc_1.n3 Gc_1.n2 2.7305
R6198 Gc_1.n5 Gc_1.t25 2.7305
R6199 Gc_1.n5 Gc_1.n4 2.7305
R6200 Gc_1.n9 Gc_1.t23 2.7305
R6201 Gc_1.n9 Gc_1.n8 2.7305
R6202 Gc_1.n13 Gc_1.t30 2.7305
R6203 Gc_1.n13 Gc_1.n12 2.7305
R6204 Gc_1.n17 Gc_1.t19 2.7305
R6205 Gc_1.n17 Gc_1.n16 2.7305
R6206 Gc_1.n21 Gc_1.t18 2.7305
R6207 Gc_1.n21 Gc_1.n20 2.7305
R6208 Gc_1.n25 Gc_1.t28 2.7305
R6209 Gc_1.n25 Gc_1.n24 2.7305
R6210 Gc_1.n29 Gc_1.t16 2.7305
R6211 Gc_1.n29 Gc_1.n28 2.7305
R6212 Gc_1.n198 Gc_1.n197 2.25044
R6213 Gc_1.n159 Gc_1.n158 1.80304
R6214 Gc_1.n194 Gc_1.n177 1.70664
R6215 Gc_1.n195 Gc_1.n1 1.65036
R6216 Gc_1.n161 Gc_1.n160 1.58193
R6217 Gc_1.n131 Gc_1.n95 1.12294
R6218 Gc_1.n135 Gc_1.n84 1.12294
R6219 Gc_1.n139 Gc_1.n73 1.12294
R6220 Gc_1.n143 Gc_1.n62 1.12294
R6221 Gc_1.n115 Gc_1.n109 1.12294
R6222 Gc_1.n129 Gc_1.n128 0.897847
R6223 Gc_1.n156 Gc_1.n155 0.897706
R6224 Gc_1.n127 Gc_1.n126 0.897685
R6225 Gc_1.n158 Gc_1.n157 0.815997
R6226 Gc_1.n113 Gc_1.n112 0.568009
R6227 Gc_1.n162 Gc_1.n161 0.525071
R6228 Gc_1.n163 Gc_1.n162 0.525071
R6229 Gc_1.n164 Gc_1.n163 0.525071
R6230 Gc_1.n165 Gc_1.n164 0.525071
R6231 Gc_1.n166 Gc_1.n165 0.525071
R6232 Gc_1.n167 Gc_1.n166 0.525071
R6233 Gc_1.n168 Gc_1.n167 0.525071
R6234 Gc_1.n169 Gc_1.n168 0.525071
R6235 Gc_1.n170 Gc_1.n169 0.525071
R6236 Gc_1.n171 Gc_1.n170 0.525071
R6237 Gc_1.n172 Gc_1.n171 0.525071
R6238 Gc_1.n173 Gc_1.n172 0.525071
R6239 Gc_1.n174 Gc_1.n173 0.525071
R6240 Gc_1.n175 Gc_1.n174 0.525071
R6241 Gc_1.n176 Gc_1.n175 0.525071
R6242 Gc_1.n177 Gc_1.n176 0.525071
R6243 Gc_1.n127 Gc_1.n117 0.463101
R6244 Gc_1.n114 Gc_1.n113 0.454175
R6245 Gc_1.n156 Gc_1.n145 0.450577
R6246 Gc_1.n138 Gc_1.n137 0.450366
R6247 Gc_1.n134 Gc_1.n133 0.449023
R6248 Gc_1.n145 Gc_1.n144 0.444603
R6249 Gc_1.n130 Gc_1.n129 0.44182
R6250 Gc_1.n137 Gc_1.n136 0.440282
R6251 Gc_1.n142 Gc_1.n141 0.437596
R6252 Gc_1.n133 Gc_1.n132 0.434458
R6253 Gc_1.n141 Gc_1.n140 0.434202
R6254 Gc_1.n117 Gc_1.n116 0.430393
R6255 Gc_1.n160 Gc_1.n159 0.306942
R6256 Gc_1.n195 Gc_1 0.234679
R6257 Gc_1.n112 Gc_1.n0 0.103625
R6258 Gc_1 Gc_1.n194 0.0866429
R6259 Gc_1.n157 Gc_1.n156 0.0335786
R6260 Gc_1.n128 Gc_1.n127 0.0335252
R6261 Gc_1.n115 Gc_1.n114 0.0292629
R6262 Gc_1.n131 Gc_1.n130 0.0292629
R6263 Gc_1.n135 Gc_1.n134 0.0292629
R6264 Gc_1.n139 Gc_1.n138 0.0292629
R6265 Gc_1.n143 Gc_1.n142 0.0292629
R6266 Gc_1.n116 Gc_1.n115 0.0283351
R6267 Gc_1.n132 Gc_1.n131 0.0283351
R6268 Gc_1.n136 Gc_1.n135 0.0283351
R6269 Gc_1.n140 Gc_1.n139 0.0283351
R6270 Gc_1.n144 Gc_1.n143 0.0283351
R6271 Gc_1 Gc_1.n199 0.017375
R6272 Gc_1.n155 Gc_1.n148 0.0163824
R6273 Gc_1 Gc_1.n198 0.00887472
R6274 Gc_1.n126 Gc_1.n120 0.0086
R6275 Gc_1.n95 Gc_1.n94 0.00797279
R6276 Gc_1.n84 Gc_1.n83 0.00797279
R6277 Gc_1.n73 Gc_1.n72 0.00797279
R6278 Gc_1.n62 Gc_1.n61 0.00797279
R6279 Gc_1.n109 Gc_1.n108 0.00797279
R6280 Gc_1.n197 Gc_1.n195 0.00615724
R6281 Gc_1.n198 Gc_1.n0 0.00324972
R6282 Gc_1.n197 Gc_1.n196 0.00192857
R6283 Gc_2.n161 Gc_2.t112 110.841
R6284 Gc_2.n190 Gc_2.n189 104.686
R6285 Gc_2.n112 Gc_2.t46 104.368
R6286 Gc_2.n163 Gc_2.n162 98.3584
R6287 Gc_2.n165 Gc_2.n164 98.3584
R6288 Gc_2.n167 Gc_2.n166 98.3584
R6289 Gc_2.n169 Gc_2.n168 98.3584
R6290 Gc_2.n171 Gc_2.n170 98.3584
R6291 Gc_2.n173 Gc_2.n172 98.3584
R6292 Gc_2.n159 Gc_2.n158 98.3584
R6293 Gc_2.n157 Gc_2.n156 98.3584
R6294 Gc_2.n155 Gc_2.n154 98.3584
R6295 Gc_2.n121 Gc_2.n120 98.3584
R6296 Gc_2.n123 Gc_2.n122 98.3584
R6297 Gc_2.n125 Gc_2.n124 98.3584
R6298 Gc_2.n200 Gc_2.n199 93.5628
R6299 Gc_2.n103 Gc_2.n101 92.4117
R6300 Gc_2.n175 Gc_2.n174 91.8697
R6301 Gc_2.n115 Gc_2.n114 39.19
R6302 Gc_2.n92 Gc_2.n91 39.19
R6303 Gc_2.n72 Gc_2.n71 39.19
R6304 Gc_2.n52 Gc_2.n51 39.19
R6305 Gc_2.n32 Gc_2.n31 39.19
R6306 Gc_2.n12 Gc_2.n11 39.19
R6307 Gc_2.n200 Gc_2.t22 34.2144
R6308 Gc_2.n101 Gc_2.t32 32.4624
R6309 Gc_2.n103 Gc_2.n102 21.8774
R6310 Gc_2.n82 Gc_2.n81 21.8774
R6311 Gc_2.n62 Gc_2.n61 21.8044
R6312 Gc_2.n42 Gc_2.n41 21.8044
R6313 Gc_2.n22 Gc_2.n21 21.8044
R6314 Gc_2.n199 Gc_2.n198 21.7314
R6315 Gc_2.n126 Gc_2.n125 21.2596
R6316 Gc_2.n160 Gc_2.n159 20.792
R6317 Gc_2.n162 Gc_2.n161 19.9794
R6318 Gc_2.n164 Gc_2.n163 19.9794
R6319 Gc_2.n166 Gc_2.n165 19.9794
R6320 Gc_2.n168 Gc_2.n167 19.9794
R6321 Gc_2.n170 Gc_2.n169 19.9794
R6322 Gc_2.n172 Gc_2.n171 19.9794
R6323 Gc_2.n174 Gc_2.n173 19.9794
R6324 Gc_2.n158 Gc_2.n157 19.9794
R6325 Gc_2.n156 Gc_2.n155 19.9794
R6326 Gc_2.n154 Gc_2.n153 19.9794
R6327 Gc_2.n120 Gc_2.n119 19.9794
R6328 Gc_2.n122 Gc_2.n121 19.9794
R6329 Gc_2.n124 Gc_2.n123 19.9794
R6330 Gc_2.n101 Gc_2.t56 12.4835
R6331 Gc_2.n102 Gc_2.t62 12.4835
R6332 Gc_2.n81 Gc_2.t54 12.4835
R6333 Gc_2.n61 Gc_2.t40 12.4835
R6334 Gc_2.n41 Gc_2.t28 12.4835
R6335 Gc_2.n21 Gc_2.t48 12.4835
R6336 Gc_2.n199 Gc_2.t8 12.4835
R6337 Gc_2.n161 Gc_2.t124 12.4835
R6338 Gc_2.n162 Gc_2.t109 12.4835
R6339 Gc_2.n163 Gc_2.t100 12.4835
R6340 Gc_2.n164 Gc_2.t123 12.4835
R6341 Gc_2.n165 Gc_2.t110 12.4835
R6342 Gc_2.n166 Gc_2.t98 12.4835
R6343 Gc_2.n167 Gc_2.t117 12.4835
R6344 Gc_2.n168 Gc_2.t119 12.4835
R6345 Gc_2.n169 Gc_2.t99 12.4835
R6346 Gc_2.n170 Gc_2.t97 12.4835
R6347 Gc_2.n171 Gc_2.t126 12.4835
R6348 Gc_2.n172 Gc_2.t138 12.4835
R6349 Gc_2.n173 Gc_2.t105 12.4835
R6350 Gc_2.n174 Gc_2.t122 12.4835
R6351 Gc_2.n159 Gc_2.t108 12.4835
R6352 Gc_2.n158 Gc_2.t101 12.4835
R6353 Gc_2.n157 Gc_2.t115 12.4835
R6354 Gc_2.n156 Gc_2.t116 12.4835
R6355 Gc_2.n155 Gc_2.t104 12.4835
R6356 Gc_2.n154 Gc_2.t132 12.4835
R6357 Gc_2.n153 Gc_2.t143 12.4835
R6358 Gc_2.n119 Gc_2.t121 12.4835
R6359 Gc_2.n120 Gc_2.t140 12.4835
R6360 Gc_2.n121 Gc_2.t113 12.4835
R6361 Gc_2.n122 Gc_2.t96 12.4835
R6362 Gc_2.n123 Gc_2.t106 12.4835
R6363 Gc_2.n124 Gc_2.t134 12.4835
R6364 Gc_2.n125 Gc_2.t111 12.4835
R6365 Gc_2.n175 Gc_2.t137 12.0283
R6366 Gc_2.n160 Gc_2.t139 11.589
R6367 Gc_2.n190 Gc_2.t30 11.5215
R6368 Gc_2.n189 Gc_2.t4 11.0965
R6369 Gc_2.n11 Gc_2.t14 11.0965
R6370 Gc_2.n31 Gc_2.t34 11.0965
R6371 Gc_2.n51 Gc_2.t50 11.0965
R6372 Gc_2.n71 Gc_2.t42 11.0965
R6373 Gc_2.n91 Gc_2.t44 11.0965
R6374 Gc_2.n114 Gc_2.t36 11.0965
R6375 Gc_2.n126 Gc_2.t127 11.079
R6376 Gc_2.n197 Gc_2.t52 10.6585
R6377 Gc_2.n201 Gc_2.t58 10.6585
R6378 Gc_2.n23 Gc_2.t0 10.5125
R6379 Gc_2.n63 Gc_2.t20 10.4395
R6380 Gc_2.n43 Gc_2.t18 10.4395
R6381 Gc_2.n104 Gc_2.t26 10.2935
R6382 Gc_2.n83 Gc_2.t16 10.2935
R6383 Gc_2.n150 Gc_2.t38 9.8555
R6384 Gc_2.n117 Gc_2.t12 9.7825
R6385 Gc_2.n33 Gc_2.t6 9.7095
R6386 Gc_2.n13 Gc_2.t60 9.6365
R6387 Gc_2.n53 Gc_2.t2 9.6365
R6388 Gc_2.n73 Gc_2.t24 9.6365
R6389 Gc_2.n93 Gc_2.t10 9.6365
R6390 Gc_2.n152 Gc_2.n149 8.1312
R6391 Gc_2.n118 Gc_2.n117 8.0005
R6392 Gc_2.n151 Gc_2.n150 6.87221
R6393 Gc_2.n127 Gc_2.n126 6.39299
R6394 Gc_2.n176 Gc_2.n160 6.3739
R6395 Gc_2.n191 Gc_2.n190 5.29995
R6396 Gc_2.n176 Gc_2.n175 5.26022
R6397 Gc_2.n26 Gc_2.n23 5.13129
R6398 Gc_2.n66 Gc_2.n63 4.86057
R6399 Gc_2.n86 Gc_2.n83 4.85692
R6400 Gc_2.n197 Gc_2.n196 4.77724
R6401 Gc_2.n46 Gc_2.n43 4.77137
R6402 Gc_2.n107 Gc_2.n104 4.67773
R6403 Gc_2.n78 Gc_2.n77 4.52348
R6404 Gc_2.n38 Gc_2.n37 4.43803
R6405 Gc_2.n18 Gc_2.n17 4.43412
R6406 Gc_2.n98 Gc_2.n97 4.36026
R6407 Gc_2.n58 Gc_2.n57 4.27334
R6408 Gc_2.n202 Gc_2.n201 4.0005
R6409 Gc_2.n133 Gc_2.n130 3.1855
R6410 Gc_2.n134 Gc_2.n109 3.1855
R6411 Gc_2.n136 Gc_2.n88 3.1855
R6412 Gc_2.n138 Gc_2.n68 3.1855
R6413 Gc_2.n140 Gc_2.n48 3.1855
R6414 Gc_2.n142 Gc_2.n28 3.1855
R6415 Gc_2.n144 Gc_2.n8 3.1855
R6416 Gc_2.n194 Gc_2.n146 3.1855
R6417 Gc_2.n192 Gc_2.n186 3.1855
R6418 Gc_2.n118 Gc_2.n113 3.05635
R6419 Gc_2.n132 Gc_2.t47 3.03383
R6420 Gc_2.n132 Gc_2.n131 3.03383
R6421 Gc_2.n130 Gc_2.t91 3.03383
R6422 Gc_2.n130 Gc_2.n129 3.03383
R6423 Gc_2.n109 Gc_2.t57 3.03383
R6424 Gc_2.n109 Gc_2.n108 3.03383
R6425 Gc_2.n100 Gc_2.t37 3.03383
R6426 Gc_2.n100 Gc_2.n99 3.03383
R6427 Gc_2.n88 Gc_2.t63 3.03383
R6428 Gc_2.n88 Gc_2.n87 3.03383
R6429 Gc_2.n80 Gc_2.t45 3.03383
R6430 Gc_2.n80 Gc_2.n79 3.03383
R6431 Gc_2.n68 Gc_2.t55 3.03383
R6432 Gc_2.n68 Gc_2.n67 3.03383
R6433 Gc_2.n60 Gc_2.t43 3.03383
R6434 Gc_2.n60 Gc_2.n59 3.03383
R6435 Gc_2.n48 Gc_2.t41 3.03383
R6436 Gc_2.n48 Gc_2.n47 3.03383
R6437 Gc_2.n40 Gc_2.t51 3.03383
R6438 Gc_2.n40 Gc_2.n39 3.03383
R6439 Gc_2.n28 Gc_2.t29 3.03383
R6440 Gc_2.n28 Gc_2.n27 3.03383
R6441 Gc_2.n20 Gc_2.t35 3.03383
R6442 Gc_2.n20 Gc_2.n19 3.03383
R6443 Gc_2.n8 Gc_2.t49 3.03383
R6444 Gc_2.n8 Gc_2.n7 3.03383
R6445 Gc_2.n6 Gc_2.t15 3.03383
R6446 Gc_2.n6 Gc_2.n5 3.03383
R6447 Gc_2.n146 Gc_2.t9 3.03383
R6448 Gc_2.n146 Gc_2.n145 3.03383
R6449 Gc_2.n184 Gc_2.t5 3.03383
R6450 Gc_2.n184 Gc_2.n183 3.03383
R6451 Gc_2.n1 Gc_2.t71 3.03383
R6452 Gc_2.n1 Gc_2.n0 3.03383
R6453 Gc_2.n4 Gc_2.t76 3.03383
R6454 Gc_2.n4 Gc_2.n3 3.03383
R6455 Gc_2.n25 Gc_2.t84 3.03383
R6456 Gc_2.n25 Gc_2.n24 3.03383
R6457 Gc_2.n45 Gc_2.t92 3.03383
R6458 Gc_2.n45 Gc_2.n44 3.03383
R6459 Gc_2.n65 Gc_2.t89 3.03383
R6460 Gc_2.n65 Gc_2.n64 3.03383
R6461 Gc_2.n85 Gc_2.t90 3.03383
R6462 Gc_2.n85 Gc_2.n84 3.03383
R6463 Gc_2.n106 Gc_2.t86 3.03383
R6464 Gc_2.n106 Gc_2.n105 3.03383
R6465 Gc_2.n188 Gc_2.t66 3.03383
R6466 Gc_2.n188 Gc_2.n187 3.03383
R6467 Gc_2.n10 Gc_2.t79 3.03383
R6468 Gc_2.n10 Gc_2.n9 3.03383
R6469 Gc_2.n30 Gc_2.t69 3.03383
R6470 Gc_2.n30 Gc_2.n29 3.03383
R6471 Gc_2.n50 Gc_2.t77 3.03383
R6472 Gc_2.n50 Gc_2.n49 3.03383
R6473 Gc_2.n70 Gc_2.t82 3.03383
R6474 Gc_2.n70 Gc_2.n69 3.03383
R6475 Gc_2.n90 Gc_2.t88 3.03383
R6476 Gc_2.n90 Gc_2.n89 3.03383
R6477 Gc_2.n111 Gc_2.t83 3.03383
R6478 Gc_2.n111 Gc_2.n110 3.03383
R6479 Gc_2.n148 Gc_2.t94 3.03383
R6480 Gc_2.n148 Gc_2.n147 3.03383
R6481 Gc_2.n186 Gc_2.t23 3.03383
R6482 Gc_2.n186 Gc_2.n185 3.03383
R6483 Gc_2.n179 Gc_2.n152 3.00506
R6484 Gc_2.n74 Gc_2.n73 2.88655
R6485 Gc_2.n77 Gc_2.n76 2.88655
R6486 Gc_2.n133 Gc_2.n132 2.84507
R6487 Gc_2.n135 Gc_2.n100 2.84507
R6488 Gc_2.n137 Gc_2.n80 2.84507
R6489 Gc_2.n139 Gc_2.n60 2.84507
R6490 Gc_2.n141 Gc_2.n40 2.84507
R6491 Gc_2.n143 Gc_2.n20 2.84507
R6492 Gc_2.n195 Gc_2.n6 2.84507
R6493 Gc_2.n193 Gc_2.n184 2.84507
R6494 Gc_2.n34 Gc_2.n33 2.75828
R6495 Gc_2.n14 Gc_2.n13 2.75828
R6496 Gc_2.n17 Gc_2.n16 2.75828
R6497 Gc_2.n196 Gc_2.n4 2.6005
R6498 Gc_2.n26 Gc_2.n25 2.6005
R6499 Gc_2.n46 Gc_2.n45 2.6005
R6500 Gc_2.n66 Gc_2.n65 2.6005
R6501 Gc_2.n86 Gc_2.n85 2.6005
R6502 Gc_2.n107 Gc_2.n106 2.6005
R6503 Gc_2.n2 Gc_2.n1 2.6005
R6504 Gc_2.n18 Gc_2.n10 2.6005
R6505 Gc_2.n38 Gc_2.n30 2.6005
R6506 Gc_2.n58 Gc_2.n50 2.6005
R6507 Gc_2.n78 Gc_2.n70 2.6005
R6508 Gc_2.n98 Gc_2.n90 2.6005
R6509 Gc_2.n128 Gc_2.n111 2.6005
R6510 Gc_2.n182 Gc_2.n148 2.6005
R6511 Gc_2.n191 Gc_2.n188 2.6005
R6512 Gc_2.n54 Gc_2.n53 2.58592
R6513 Gc_2.n57 Gc_2.n56 2.58592
R6514 Gc_2.n96 Gc_2.n95 2.49787
R6515 Gc_2.n76 Gc_2.n75 2.49787
R6516 Gc_2.n56 Gc_2.n55 2.49787
R6517 Gc_2.n36 Gc_2.n35 2.49787
R6518 Gc_2.n16 Gc_2.n15 2.49787
R6519 Gc_2.n94 Gc_2.n93 2.4825
R6520 Gc_2.n97 Gc_2.n96 2.4825
R6521 Gc_2.n37 Gc_2.n36 2.43383
R6522 Gc_2.n177 Gc_2.n176 1.65162
R6523 Gc_2.n13 Gc_2.n12 1.4605
R6524 Gc_2.n53 Gc_2.n52 1.4605
R6525 Gc_2.n73 Gc_2.n72 1.4605
R6526 Gc_2.n93 Gc_2.n92 1.4605
R6527 Gc_2.n113 Gc_2.n112 1.44187
R6528 Gc_2.n33 Gc_2.n32 1.3875
R6529 Gc_2.n116 Gc_2.n115 1.2415
R6530 Gc_2.n179 Gc_2.n178 1.13001
R6531 Gc_2.n128 Gc_2.n127 1.01243
R6532 Gc_2.n202 Gc_2.n2 1.00561
R6533 Gc_2.n37 Gc_2.n34 0.973833
R6534 Gc_2.n152 Gc_2.n151 0.893792
R6535 Gc_2.n77 Gc_2.n74 0.849337
R6536 Gc_2.n17 Gc_2.n14 0.811611
R6537 Gc_2.n182 Gc_2.n181 0.804097
R6538 Gc_2.n57 Gc_2.n54 0.760917
R6539 Gc_2.n97 Gc_2.n94 0.7305
R6540 Gc_2.n196 Gc_2.n195 0.5855
R6541 Gc_2.n143 Gc_2.n26 0.5855
R6542 Gc_2.n141 Gc_2.n46 0.5855
R6543 Gc_2.n139 Gc_2.n66 0.5855
R6544 Gc_2.n137 Gc_2.n86 0.5855
R6545 Gc_2.n135 Gc_2.n107 0.5855
R6546 Gc_2.n193 Gc_2.n2 0.5855
R6547 Gc_2.n134 Gc_2.n133 0.44291
R6548 Gc_2.n135 Gc_2.n134 0.44291
R6549 Gc_2.n136 Gc_2.n135 0.44291
R6550 Gc_2.n137 Gc_2.n136 0.44291
R6551 Gc_2.n138 Gc_2.n137 0.44291
R6552 Gc_2.n139 Gc_2.n138 0.44291
R6553 Gc_2.n140 Gc_2.n139 0.44291
R6554 Gc_2.n141 Gc_2.n140 0.44291
R6555 Gc_2.n142 Gc_2.n141 0.44291
R6556 Gc_2.n143 Gc_2.n142 0.44291
R6557 Gc_2.n144 Gc_2.n143 0.44291
R6558 Gc_2.n195 Gc_2.n144 0.44291
R6559 Gc_2.n195 Gc_2.n194 0.44291
R6560 Gc_2.n193 Gc_2.n192 0.44291
R6561 Gc_2.n104 Gc_2.n103 0.2925
R6562 Gc_2.n83 Gc_2.n82 0.2925
R6563 Gc_2.n144 Gc_2.n18 0.245065
R6564 Gc_2.n142 Gc_2.n38 0.245065
R6565 Gc_2.n140 Gc_2.n58 0.245065
R6566 Gc_2.n138 Gc_2.n78 0.245065
R6567 Gc_2.n136 Gc_2.n98 0.245065
R6568 Gc_2.n134 Gc_2.n128 0.245065
R6569 Gc_2.n194 Gc_2.n182 0.245065
R6570 Gc_2.n192 Gc_2.n191 0.245065
R6571 Gc_2.n194 Gc_2 0.236886
R6572 Gc_2.n63 Gc_2.n62 0.2195
R6573 Gc_2.n43 Gc_2.n42 0.2195
R6574 Gc_2 Gc_2.n193 0.206524
R6575 Gc_2.n23 Gc_2.n22 0.1465
R6576 Gc_2.n198 Gc_2.n197 0.0735
R6577 Gc_2.n201 Gc_2.n200 0.0735
R6578 Gc_2.n117 Gc_2.n116 0.0735
R6579 Gc_2.n178 Gc_2.n177 0.0332273
R6580 Gc_2.n180 Gc_2.n179 0.0241252
R6581 Gc_2.n181 Gc_2.n180 0.0141364
R6582 Gc_2.n127 Gc_2.n118 0.0133843
R6583 Gc_2 Gc_2.n202 0.0123033
R6584 G2.n1 G2.n0 102.993
R6585 G2.n3 G2.n2 101.566
R6586 G2.n6 G2.n5 99.4048
R6587 G2.n8 G2.n7 99.4048
R6588 G2.n10 G2.n4 70.7294
R6589 G2.n9 G2.n8 39.5325
R6590 G2.n10 G2.n9 39.4595
R6591 G2.n4 G2.n3 37.7091
R6592 G2.n0 G2.t10 29.4988
R6593 G2.n5 G2.t4 29.1477
R6594 G2.t10 G2.t17 23.7985
R6595 G2.t21 G2.t24 23.7985
R6596 G2.t3 G2.t7 23.7985
R6597 G2.t14 G2.t18 23.7985
R6598 G2.t5 G2.t11 23.7985
R6599 G2.t4 G2.t8 23.7985
R6600 G2.t20 G2.t23 23.7985
R6601 G2.t9 G2.t16 23.7985
R6602 G2.t6 G2.t15 23.7985
R6603 G2.t19 G2.t22 23.7985
R6604 G2.n2 G2.n1 16.5048
R6605 G2.n7 G2.n6 16.1537
R6606 G2.n9 G2.t12 13.1405
R6607 G2.n4 G2.t13 13.0675
R6608 G2.t1 G2.n10 13.0675
R6609 G2.n0 G2.t21 12.9945
R6610 G2.n1 G2.t3 12.9945
R6611 G2.n2 G2.t14 12.9945
R6612 G2.n3 G2.t5 12.9945
R6613 G2.n5 G2.t20 12.9945
R6614 G2.n6 G2.t9 12.9945
R6615 G2.n7 G2.t6 12.9945
R6616 G2.n8 G2.t19 12.9945
R6617 G2.n11 G2.t25 12.6295
R6618 G2.n11 G2.t1 11.1695
R6619 G2.n14 G2.n11 4.0005
R6620 G2 G2.n13 3.34309
R6621 G2.n13 G2.t2 2.7305
R6622 G2.n13 G2.n12 2.7305
R6623 G2.n14 G2 0.0935
R6624 G2 G2.n14 0.0065
R6625 SD2_5 SD2_5.n10 4.78409
R6626 SD2_5.n4 SD2_5.n3 3.44212
R6627 SD2_5.n9 SD2_5.n8 3.43911
R6628 SD2_5.n15 SD2_5.n12 3.41246
R6629 SD2_5.n20 SD2_5.n19 3.38757
R6630 SD2_5.n15 SD2_5.n14 3.38387
R6631 SD2_5.n4 SD2_5.n1 3.38278
R6632 SD2_5.n9 SD2_5.n6 3.38274
R6633 SD2_5 SD2_5.n17 3.29941
R6634 SD2_5.n10 SD2_5.n4 2.87871
R6635 SD2_5.n21 SD2_5.n15 2.87758
R6636 SD2_5.n17 SD2_5.t0 2.7305
R6637 SD2_5.n17 SD2_5.n16 2.7305
R6638 SD2_5.n12 SD2_5.t13 2.7305
R6639 SD2_5.n12 SD2_5.n11 2.7305
R6640 SD2_5.n14 SD2_5.t15 2.7305
R6641 SD2_5.n14 SD2_5.n13 2.7305
R6642 SD2_5.n6 SD2_5.t10 2.7305
R6643 SD2_5.n6 SD2_5.n5 2.7305
R6644 SD2_5.n8 SD2_5.t14 2.7305
R6645 SD2_5.n8 SD2_5.n7 2.7305
R6646 SD2_5.n1 SD2_5.t4 2.7305
R6647 SD2_5.n1 SD2_5.n0 2.7305
R6648 SD2_5.n3 SD2_5.t2 2.7305
R6649 SD2_5.n3 SD2_5.n2 2.7305
R6650 SD2_5.n19 SD2_5.t7 2.7305
R6651 SD2_5.n19 SD2_5.n18 2.7305
R6652 SD2_5.n10 SD2_5.n9 2.2505
R6653 SD2_5.n21 SD2_5.n20 2.2505
R6654 SD2_5.n20 SD2_5 0.116906
R6655 SD2_5 SD2_5.n21 0.00283766
R6656 SDc_2.n59 SDc_2.n58 3.51171
R6657 SDc_2.n75 SDc_2.n38 3.49726
R6658 SDc_2.n103 SDc_2.n6 3.49243
R6659 SDc_2.n114 SDc_2.n110 3.0975
R6660 SDc_2 SDc_2.n1 3.08791
R6661 SDc_2.n69 SDc_2.n40 3.08362
R6662 SDc_2.n66 SDc_2.n45 3.08133
R6663 SDc_2.n87 SDc_2.n26 3.07918
R6664 SDc_2.n81 SDc_2.n36 3.07654
R6665 SDc_2.n60 SDc_2.n54 3.07634
R6666 SDc_2.n92 SDc_2.n24 3.07504
R6667 SDc_2.n94 SDc_2.n20 3.0749
R6668 SDc_2.n63 SDc_2.n50 3.07479
R6669 SDc_2.n84 SDc_2.n31 3.07402
R6670 SDc_2.n100 SDc_2.n11 3.0734
R6671 SDc_2.n97 SDc_2.n16 3.07148
R6672 SDc_2.n112 SDc_2.t2 3.03383
R6673 SDc_2.n112 SDc_2.n111 3.03383
R6674 SDc_2.n3 SDc_2.t48 3.03383
R6675 SDc_2.n3 SDc_2.n2 3.03383
R6676 SDc_2.n105 SDc_2.t26 3.03383
R6677 SDc_2.n105 SDc_2.n104 3.03383
R6678 SDc_2.n8 SDc_2.t51 3.03383
R6679 SDc_2.n8 SDc_2.n7 3.03383
R6680 SDc_2.n13 SDc_2.t15 3.03383
R6681 SDc_2.n13 SDc_2.n12 3.03383
R6682 SDc_2.n18 SDc_2.t53 3.03383
R6683 SDc_2.n18 SDc_2.n17 3.03383
R6684 SDc_2.n22 SDc_2.t6 3.03383
R6685 SDc_2.n22 SDc_2.n21 3.03383
R6686 SDc_2.n89 SDc_2.t60 3.03383
R6687 SDc_2.n89 SDc_2.n88 3.03383
R6688 SDc_2.n28 SDc_2.t12 3.03383
R6689 SDc_2.n28 SDc_2.n27 3.03383
R6690 SDc_2.n33 SDc_2.t56 3.03383
R6691 SDc_2.n33 SDc_2.n32 3.03383
R6692 SDc_2.n38 SDc_2.t61 3.03383
R6693 SDc_2.n38 SDc_2.n37 3.03383
R6694 SDc_2.n77 SDc_2.t17 3.03383
R6695 SDc_2.n77 SDc_2.n76 3.03383
R6696 SDc_2.n40 SDc_2.t10 3.03383
R6697 SDc_2.n40 SDc_2.n39 3.03383
R6698 SDc_2.n71 SDc_2.t57 3.03383
R6699 SDc_2.n71 SDc_2.n70 3.03383
R6700 SDc_2.n42 SDc_2.t23 3.03383
R6701 SDc_2.n42 SDc_2.n41 3.03383
R6702 SDc_2.n47 SDc_2.t55 3.03383
R6703 SDc_2.n47 SDc_2.n46 3.03383
R6704 SDc_2.n52 SDc_2.t19 3.03383
R6705 SDc_2.n52 SDc_2.n51 3.03383
R6706 SDc_2.n56 SDc_2.t59 3.03383
R6707 SDc_2.n56 SDc_2.n55 3.03383
R6708 SDc_2.n58 SDc_2.t18 3.03383
R6709 SDc_2.n58 SDc_2.n57 3.03383
R6710 SDc_2.n54 SDc_2.t63 3.03383
R6711 SDc_2.n54 SDc_2.n53 3.03383
R6712 SDc_2.n50 SDc_2.t21 3.03383
R6713 SDc_2.n50 SDc_2.n49 3.03383
R6714 SDc_2.n45 SDc_2.t58 3.03383
R6715 SDc_2.n45 SDc_2.n44 3.03383
R6716 SDc_2.n36 SDc_2.t29 3.03383
R6717 SDc_2.n36 SDc_2.n35 3.03383
R6718 SDc_2.n31 SDc_2.t54 3.03383
R6719 SDc_2.n31 SDc_2.n30 3.03383
R6720 SDc_2.n26 SDc_2.t13 3.03383
R6721 SDc_2.n26 SDc_2.n25 3.03383
R6722 SDc_2.n24 SDc_2.t52 3.03383
R6723 SDc_2.n24 SDc_2.n23 3.03383
R6724 SDc_2.n20 SDc_2.t30 3.03383
R6725 SDc_2.n20 SDc_2.n19 3.03383
R6726 SDc_2.n16 SDc_2.t62 3.03383
R6727 SDc_2.n16 SDc_2.n15 3.03383
R6728 SDc_2.n11 SDc_2.t3 3.03383
R6729 SDc_2.n11 SDc_2.n10 3.03383
R6730 SDc_2.n6 SDc_2.t50 3.03383
R6731 SDc_2.n6 SDc_2.n5 3.03383
R6732 SDc_2.n1 SDc_2.t11 3.03383
R6733 SDc_2.n1 SDc_2.n0 3.03383
R6734 SDc_2.n110 SDc_2.t49 3.03383
R6735 SDc_2.n110 SDc_2.n109 3.03383
R6736 SDc_2.n95 SDc_2.n18 2.75468
R6737 SDc_2.n61 SDc_2.n52 2.75468
R6738 SDc_2.n93 SDc_2.n22 2.75423
R6739 SDc_2.n59 SDc_2.n56 2.38139
R6740 SDc_2.n107 SDc_2.n106 2.24447
R6741 SDc_2.n73 SDc_2.n72 2.24419
R6742 SDc_2.n79 SDc_2.n78 2.24419
R6743 SDc_2.n108 SDc_2.n4 1.49481
R6744 SDc_2.n91 SDc_2.n90 1.4947
R6745 SDc_2.n82 SDc_2.n34 1.49456
R6746 SDc_2.n101 SDc_2.n9 1.49456
R6747 SDc_2.n64 SDc_2.n48 1.49431
R6748 SDc_2.n67 SDc_2.n43 1.49431
R6749 SDc_2.n85 SDc_2.n29 1.49431
R6750 SDc_2.n98 SDc_2.n14 1.49431
R6751 SDc_2.n9 SDc_2.n8 1.26132
R6752 SDc_2.n14 SDc_2.n13 1.26101
R6753 SDc_2.n48 SDc_2.n47 1.26087
R6754 SDc_2.n106 SDc_2.n105 1.26056
R6755 SDc_2.n29 SDc_2.n28 1.26056
R6756 SDc_2.n34 SDc_2.n33 1.26043
R6757 SDc_2.n4 SDc_2.n3 1.25998
R6758 SDc_2.n90 SDc_2.n89 1.25998
R6759 SDc_2.n78 SDc_2.n77 1.25998
R6760 SDc_2.n72 SDc_2.n71 1.25998
R6761 SDc_2.n43 SDc_2.n42 1.25966
R6762 SDc_2.n113 SDc_2.n112 1.24434
R6763 SDc_2.n114 SDc_2.n113 1.14086
R6764 SDc_2.n60 SDc_2.n59 0.612813
R6765 SDc_2.n102 SDc_2.n101 0.611577
R6766 SDc_2.n92 SDc_2.n91 0.610706
R6767 SDc_2.n94 SDc_2.n93 0.608363
R6768 SDc_2.n68 SDc_2.n67 0.596198
R6769 SDc_2.n108 SDc_2.n107 0.59153
R6770 SDc_2.n74 SDc_2.n73 0.591483
R6771 SDc_2.n115 SDc_2.n114 0.585814
R6772 SDc_2.n83 SDc_2.n82 0.584906
R6773 SDc_2.n65 SDc_2.n64 0.583676
R6774 SDc_2.n62 SDc_2.n61 0.582832
R6775 SDc_2.n96 SDc_2.n95 0.582832
R6776 SDc_2.n99 SDc_2.n98 0.582069
R6777 SDc_2.n86 SDc_2.n85 0.579994
R6778 SDc_2.n80 SDc_2.n79 0.577353
R6779 SDc_2.n113 SDc_2 0.0774668
R6780 SDc_2 SDc_2.n115 0.0278418
R6781 SDc_2.n66 SDc_2.n65 0.0244241
R6782 SDc_2.n87 SDc_2.n86 0.0244241
R6783 SDc_2.n97 SDc_2.n96 0.0244241
R6784 SDc_2.n100 SDc_2.n99 0.0232848
R6785 SDc_2.n81 SDc_2.n80 0.0221456
R6786 SDc_2.n84 SDc_2.n83 0.0221456
R6787 SDc_2.n63 SDc_2.n62 0.0210063
R6788 SDc_2.n64 SDc_2.n63 0.0183749
R6789 SDc_2.n82 SDc_2.n81 0.0176185
R6790 SDc_2.n85 SDc_2.n84 0.0172357
R6791 SDc_2.n69 SDc_2.n68 0.016908
R6792 SDc_2.n79 SDc_2.n75 0.016908
R6793 SDc_2.n101 SDc_2.n100 0.0164793
R6794 SDc_2.n107 SDc_2.n103 0.0163417
R6795 SDc_2.n61 SDc_2.n60 0.015337
R6796 SDc_2.n93 SDc_2.n92 0.015337
R6797 SDc_2.n91 SDc_2.n87 0.0150107
R6798 SDc_2.n67 SDc_2.n66 0.0149572
R6799 SDc_2.n98 SDc_2.n97 0.0149572
R6800 SDc_2.n73 SDc_2.n69 0.0146295
R6801 SDc_2.n75 SDc_2.n74 0.0146295
R6802 SDc_2.n95 SDc_2.n94 0.0141978
R6803 SDc_2 SDc_2.n108 0.0126401
R6804 SDc_2.n103 SDc_2.n102 0.00277848
R6805 b4b.n3 b4b.t8 135.346
R6806 b4b.n6 b4b.t12 122.275
R6807 b4b.n7 b4b.t16 87.2463
R6808 b4b.n2 b4b.t10 86.6191
R6809 b4b.n3 b4b.n2 75.3342
R6810 b4b.t12 b4b.t4 68.4445
R6811 b4b.t7 b4b.t3 56.6204
R6812 b4b.n8 b4b.n6 52.2803
R6813 b4b.t10 b4b.t13 41.8693
R6814 b4b.n9 b4b.n8 32.8633
R6815 b4b b4b.t9 19.4226
R6816 b4b.t3 b4b.n3 18.8389
R6817 b4b.n2 b4b.t2 18.7955
R6818 b4b.n6 b4b.t6 18.4057
R6819 b4b.n7 b4b.t11 18.0315
R6820 b4b.n5 b4b.n4 16.0319
R6821 b4b.n1 b4b.n0 15.4944
R6822 b4b.n0 b4b.t15 10.7315
R6823 b4b.n1 b4b.t17 10.7315
R6824 b4b.n0 b4b.t5 9.6365
R6825 b4b.t13 b4b.n1 9.6365
R6826 b4b.n18 b4b.n13 9.49418
R6827 b4b.n17 b4b.n16 9.39762
R6828 b4b.n4 b4b.t18 9.3445
R6829 b4b.n4 b4b.t7 8.9065
R6830 b4b.n5 b4b.t14 8.9065
R6831 b4b.t4 b4b.n5 7.1545
R6832 b4b.n12 b4b.n11 4.5005
R6833 b4b.n8 b4b.n7 3.6505
R6834 b4b.n17 b4b.n15 2.37493
R6835 b4b.n19 b4b.n18 2.2505
R6836 b4b.n19 b4b.n12 0.113387
R6837 b4b.n14 b4b.n12 0.0210063
R6838 b4b.n15 b4b.n14 0.0118924
R6839 b4b.n11 b4b.n9 0.0112067
R6840 b4b b4b.n19 0.00318657
R6841 b4b.n18 b4b.n17 0.0031087
R6842 b4b.n11 b4b.n10 0.0021391
R6843 b4b.n10 b4b 0.00213881
R6844 OUT4.n31 OUT4.n30 15.3782
R6845 OUT4.n32 OUT4.n31 8.93169
R6846 OUT4.n5 OUT4.t15 6.44473
R6847 OUT4.n2 OUT4.n0 6.42383
R6848 OUT4.n2 OUT4.n1 5.8805
R6849 OUT4.n33 OUT4.t9 5.8805
R6850 OUT4.n32 OUT4.t12 5.8805
R6851 OUT4.n6 OUT4.n4 5.8805
R6852 OUT4.n7 OUT4.n3 5.8805
R6853 OUT4.n5 OUT4.t14 5.8805
R6854 OUT4.n27 OUT4.n26 3.85309
R6855 OUT4.n16 OUT4.n15 3.82489
R6856 OUT4.n17 OUT4.n11 3.1505
R6857 OUT4.n16 OUT4.n13 3.1505
R6858 OUT4.n18 OUT4.n9 3.1505
R6859 OUT4.n28 OUT4.n22 3.1505
R6860 OUT4.n27 OUT4.n24 3.1505
R6861 OUT4.n29 OUT4.n20 3.1505
R6862 OUT4.n9 OUT4.t7 2.7305
R6863 OUT4.n9 OUT4.n8 2.7305
R6864 OUT4.n13 OUT4.t17 2.7305
R6865 OUT4.n13 OUT4.n12 2.7305
R6866 OUT4.n11 OUT4.t23 2.7305
R6867 OUT4.n11 OUT4.n10 2.7305
R6868 OUT4.n15 OUT4.t4 2.7305
R6869 OUT4.n15 OUT4.n14 2.7305
R6870 OUT4.n20 OUT4.t22 2.7305
R6871 OUT4.n20 OUT4.n19 2.7305
R6872 OUT4.n24 OUT4.t0 2.7305
R6873 OUT4.n24 OUT4.n23 2.7305
R6874 OUT4.n22 OUT4.t3 2.7305
R6875 OUT4.n22 OUT4.n21 2.7305
R6876 OUT4.n26 OUT4.t19 2.7305
R6877 OUT4.n26 OUT4.n25 2.7305
R6878 OUT4.n31 OUT4.n7 2.72598
R6879 OUT4.n6 OUT4.n5 1.79955
R6880 OUT4 OUT4.n33 1.70642
R6881 OUT4.n30 OUT4.n18 1.02158
R6882 OUT4.n29 OUT4.n28 0.689162
R6883 OUT4.n18 OUT4.n17 0.669768
R6884 OUT4.n33 OUT4.n32 0.599276
R6885 OUT4.n7 OUT4.n6 0.575794
R6886 OUT4.n28 OUT4.n27 0.483385
R6887 OUT4.n17 OUT4.n16 0.474274
R6888 OUT4.n30 OUT4.n29 0.132857
R6889 OUT4 OUT4.n2 0.0205
R6890 b5.t19 b5.t7 109.68
R6891 b5 b5.t11 51.8095
R6892 b5.n14 b5.n13 48.5408
R6893 b5.n11 b5.t6 28.2458
R6894 b5.n4 b5.t16 25.4465
R6895 b5.t6 b5.t9 21.5355
R6896 b5.t16 b5.t18 21.5355
R6897 b5.n16 b5.t4 20.3746
R6898 b5.n4 b5.t13 14.4545
R6899 b5.n5 b5.t21 14.4545
R6900 b5.n10 b5.t12 14.4545
R6901 b5.n11 b5.n10 14.398
R6902 b5.n13 b5.t23 14.1625
R6903 b5.n14 b5.t10 14.1625
R6904 b5.t26 b5.n6 13.9435
R6905 b5.n9 b5.t20 13.9435
R6906 b5.n12 b5.n11 13.9116
R6907 b5.n13 b5.n12 13.5102
R6908 b5.n15 b5.t25 13.2865
R6909 b5.n7 b5.t26 12.1185
R6910 b5.t20 b5.n8 12.1185
R6911 b5.n5 b5.n4 11.5035
R6912 b5.n9 b5.n6 11.5035
R6913 b5.n6 b5.n5 11.5035
R6914 b5.n10 b5.n9 11.5035
R6915 b5.n15 b5.n14 10.7362
R6916 b5.n0 b5.t22 10.4395
R6917 b5.t7 b5.n1 10.4395
R6918 b5.n2 b5.t19 10.4395
R6919 b5.t4 b5.n3 10.4395
R6920 b5.n2 b5.t5 10.2935
R6921 b5.n0 b5.t8 10.2935
R6922 b5.n1 b5.t17 10.2935
R6923 b5.n3 b5.t15 10.2935
R6924 b5.n12 b5.t14 9.6365
R6925 b5.n17 b5.t0 9.49371
R6926 b5.n1 b5.n0 9.4905
R6927 b5.n3 b5.n2 9.4905
R6928 b5.n7 b5.t3 9.4175
R6929 b5.n8 b5.t24 9.4175
R6930 b5.n17 b5.t1 9.3756
R6931 b5.n8 b5.n7 9.14749
R6932 b5.n18 b5.n16 5.49961
R6933 b5.n16 b5.n15 5.23946
R6934 b5.n11 b5.t2 4.3805
R6935 b5.n18 b5.n17 3.24728
R6936 b5 b5.n18 0.374557
R6937 C32_U.n103 C32_U.n102 107.18
R6938 C32_U.n127 C32_U.n123 107.18
R6939 C32_U.n13 C32_U.n12 103.823
R6940 C32_U.n18 C32_U.n17 103.823
R6941 C32_U.n23 C32_U.n22 103.823
R6942 C32_U.n28 C32_U.n27 103.823
R6943 C32_U.n146 C32_U.n145 103.823
R6944 C32_U.n144 C32_U.n143 103.823
R6945 C32_U.n55 C32_U.n54 103.823
R6946 C32_U.n53 C32_U.n52 103.823
R6947 C32_U.n51 C32_U.n50 103.823
R6948 C32_U.n130 C32_U.n128 103.823
R6949 C32_U.n12 C32_U.n11 23.4254
R6950 C32_U.n147 C32_U.n146 23.4254
R6951 C32_U.n17 C32_U.n13 21.0894
R6952 C32_U.n22 C32_U.n18 21.0894
R6953 C32_U.n27 C32_U.n23 21.0894
R6954 C32_U.n145 C32_U.n144 21.0894
R6955 C32_U.n143 C32_U.n142 21.0894
R6956 C32_U.n29 C32_U.n28 21.0894
R6957 C32_U.n54 C32_U.n53 21.0894
R6958 C32_U.n52 C32_U.n51 21.0894
R6959 C32_U.n50 C32_U.n49 21.0894
R6960 C32_U.n102 C32_U.n101 21.0894
R6961 C32_U.n128 C32_U.n127 21.0894
R6962 C32_U.n130 C32_U.n129 21.0894
R6963 C32_U.n56 C32_U.n55 21.0894
R6964 C32_U.n55 C32_U.t46 14.0895
R6965 C32_U.n53 C32_U.t60 14.0895
R6966 C32_U.n51 C32_U.t42 14.0895
R6967 C32_U.n49 C32_U.t52 14.0895
R6968 C32_U.n102 C32_U.t48 14.0895
R6969 C32_U.n128 C32_U.t32 14.0895
R6970 C32_U.n129 C32_U.t58 14.0895
R6971 C32_U.n12 C32_U.t26 12.7025
R6972 C32_U.n13 C32_U.t36 12.7025
R6973 C32_U.n18 C32_U.t40 12.7025
R6974 C32_U.n23 C32_U.t56 12.7025
R6975 C32_U.n28 C32_U.t38 12.7025
R6976 C32_U.n146 C32_U.t44 12.7025
R6977 C32_U.n144 C32_U.t50 12.7025
R6978 C32_U.n142 C32_U.t34 12.7025
R6979 C32_U.n42 C32_U.t10 10.7315
R6980 C32_U.n45 C32_U.t16 10.7315
R6981 C32_U.n48 C32_U.t24 10.7315
R6982 C32_U.n100 C32_U.t8 10.7315
R6983 C32_U.n103 C32_U.t4 10.7315
R6984 C32_U.n123 C32_U.t30 10.7315
R6985 C32_U.n126 C32_U.t62 10.7315
R6986 C32_U.n11 C32_U.t54 10.3665
R6987 C32_U.n16 C32_U.t0 10.3665
R6988 C32_U.n21 C32_U.t14 10.3665
R6989 C32_U.n26 C32_U.t28 10.3665
R6990 C32_U.n147 C32_U.t20 10.3665
R6991 C32_U.n4 C32_U.t2 10.3665
R6992 C32_U.n131 C32_U.t18 10.2068
R6993 C32_U.n139 C32_U.t6 9.14387
R6994 C32_U.n62 C32_U.t22 8.1765
R6995 C32_U.n36 C32_U.t12 7.8845
R6996 C32_U.n126 C32_U.n125 7.54963
R6997 C32_U.n42 C32_U.n41 7.51539
R6998 C32_U.n45 C32_U.n44 7.51309
R6999 C32_U.n100 C32_U.n99 7.50659
R7000 C32_U.n48 C32_U.n47 7.50213
R7001 C32_U.n11 C32_U.n10 7.49191
R7002 C32_U.n16 C32_U.n15 7.48719
R7003 C32_U.n21 C32_U.n20 7.48706
R7004 C32_U.n26 C32_U.n25 7.47354
R7005 C32_U.n4 C32_U.n3 7.4684
R7006 C32_U.n105 C32_U.n96 6.07641
R7007 C32_U.n121 C32_U.t77 6.07641
R7008 C32_U.n104 C32_U.n97 6.03311
R7009 C32_U.n122 C32_U.t31 6.01354
R7010 C32_U.n123 C32_U.n122 4.09071
R7011 C32_U.n104 C32_U.n103 4.07073
R7012 C32_U.n135 C32_U 4.0021
R7013 C32_U.n148 C32_U.n147 4.0005
R7014 C32_U.n134 C32_U.n133 3.57136
R7015 C32_U.n35 C32_U.n30 3.54754
R7016 C32_U.n61 C32_U.n57 3.54049
R7017 C32_U.n60 C32_U.n59 3.4968
R7018 C32_U.n148 C32_U.n1 3.49193
R7019 C32_U.n7 C32_U.n6 3.46025
R7020 C32_U.n33 C32_U.n32 3.43615
R7021 C32_U.n54 C32_U.n42 3.3585
R7022 C32_U.n52 C32_U.n45 3.3585
R7023 C32_U.n50 C32_U.n48 3.3585
R7024 C32_U.n101 C32_U.n100 3.3585
R7025 C32_U.n127 C32_U.n126 3.3585
R7026 C32_U.n93 C32_U.t72 3.03383
R7027 C32_U.n93 C32_U.n92 3.03383
R7028 C32_U.n89 C32_U.t71 3.03383
R7029 C32_U.n89 C32_U.n88 3.03383
R7030 C32_U.n85 C32_U.t75 3.03383
R7031 C32_U.n85 C32_U.n84 3.03383
R7032 C32_U.n81 C32_U.t64 3.03383
R7033 C32_U.n81 C32_U.n80 3.03383
R7034 C32_U.n77 C32_U.t69 3.03383
R7035 C32_U.n77 C32_U.n76 3.03383
R7036 C32_U.n73 C32_U.t93 3.03383
R7037 C32_U.n73 C32_U.n72 3.03383
R7038 C32_U.n69 C32_U.t81 3.03383
R7039 C32_U.n69 C32_U.n68 3.03383
R7040 C32_U.n67 C32_U.t66 3.03383
R7041 C32_U.n67 C32_U.n66 3.03383
R7042 C32_U.n71 C32_U.t68 3.03383
R7043 C32_U.n71 C32_U.n70 3.03383
R7044 C32_U.n75 C32_U.t95 3.03383
R7045 C32_U.n75 C32_U.n74 3.03383
R7046 C32_U.n79 C32_U.t92 3.03383
R7047 C32_U.n79 C32_U.n78 3.03383
R7048 C32_U.n83 C32_U.t73 3.03383
R7049 C32_U.n83 C32_U.n82 3.03383
R7050 C32_U.n87 C32_U.t91 3.03383
R7051 C32_U.n87 C32_U.n86 3.03383
R7052 C32_U.n91 C32_U.t87 3.03383
R7053 C32_U.n91 C32_U.n90 3.03383
R7054 C32_U.n95 C32_U.t83 3.03383
R7055 C32_U.n95 C32_U.n94 3.03383
R7056 C32_U.n120 C32_U.n67 3.00941
R7057 C32_U.n118 C32_U.n71 3.00941
R7058 C32_U.n116 C32_U.n75 3.00941
R7059 C32_U.n114 C32_U.n79 3.00941
R7060 C32_U.n112 C32_U.n83 3.00941
R7061 C32_U.n110 C32_U.n87 3.00941
R7062 C32_U.n108 C32_U.n91 3.00941
R7063 C32_U.n106 C32_U.n95 3.00941
R7064 C32_U.n107 C32_U.n93 2.99767
R7065 C32_U.n109 C32_U.n89 2.99767
R7066 C32_U.n111 C32_U.n85 2.99767
R7067 C32_U.n113 C32_U.n81 2.99767
R7068 C32_U.n115 C32_U.n77 2.99767
R7069 C32_U.n117 C32_U.n73 2.99767
R7070 C32_U.n119 C32_U.n69 2.99767
R7071 C32_U.n64 C32_U.n63 2.88757
R7072 C32_U.n38 C32_U.n37 2.88525
R7073 C32_U.n131 C32_U.n130 2.8333
R7074 C32_U.n10 C32_U.t55 2.7305
R7075 C32_U.n10 C32_U.n9 2.7305
R7076 C32_U.n15 C32_U.t37 2.7305
R7077 C32_U.n15 C32_U.n14 2.7305
R7078 C32_U.n20 C32_U.t41 2.7305
R7079 C32_U.n20 C32_U.n19 2.7305
R7080 C32_U.n25 C32_U.t57 2.7305
R7081 C32_U.n25 C32_U.n24 2.7305
R7082 C32_U.n1 C32_U.t45 2.7305
R7083 C32_U.n1 C32_U.n0 2.7305
R7084 C32_U.n3 C32_U.t51 2.7305
R7085 C32_U.n3 C32_U.n2 2.7305
R7086 C32_U.n6 C32_U.t35 2.7305
R7087 C32_U.n6 C32_U.n5 2.7305
R7088 C32_U.n32 C32_U.t39 2.7305
R7089 C32_U.n32 C32_U.n31 2.7305
R7090 C32_U.n41 C32_U.t61 2.7305
R7091 C32_U.n41 C32_U.n40 2.7305
R7092 C32_U.n44 C32_U.t43 2.7305
R7093 C32_U.n44 C32_U.n43 2.7305
R7094 C32_U.n47 C32_U.t53 2.7305
R7095 C32_U.n47 C32_U.n46 2.7305
R7096 C32_U.n99 C32_U.t49 2.7305
R7097 C32_U.n99 C32_U.n98 2.7305
R7098 C32_U.n125 C32_U.t33 2.7305
R7099 C32_U.n125 C32_U.n124 2.7305
R7100 C32_U.n133 C32_U.t59 2.7305
R7101 C32_U.n133 C32_U.n132 2.7305
R7102 C32_U.n59 C32_U.t47 2.7305
R7103 C32_U.n59 C32_U.n58 2.7305
R7104 C32_U.n17 C32_U.n16 2.3365
R7105 C32_U.n22 C32_U.n21 2.3365
R7106 C32_U.n27 C32_U.n26 2.3365
R7107 C32_U.n145 C32_U.n4 2.3365
R7108 C32_U.n65 C32_U.n64 2.2505
R7109 C32_U.n39 C32_U.n38 2.2505
R7110 C32_U.n138 C32_U.n137 2.2505
R7111 C32_U.n135 C32_U.n134 2.2505
R7112 C32_U.n57 C32_U.n56 2.17864
R7113 C32_U.n37 C32_U.n36 2.1175
R7114 C32_U.n63 C32_U.n62 2.1175
R7115 C32_U.n141 C32_U.n138 1.78472
R7116 C32_U.n105 C32_U.n104 1.74861
R7117 C32_U.n122 C32_U.n121 1.7405
R7118 C32_U.n143 C32_U.n141 1.31264
R7119 C32_U.n137 C32_U.n39 1.27751
R7120 C32_U.n140 C32_U.n139 1.18026
R7121 C32_U.n30 C32_U.n29 1.1585
R7122 C32_U.n137 C32_U.n136 0.952132
R7123 C32_U.n134 C32_U.n131 0.761354
R7124 C32_U.n136 C32_U.n65 0.640509
R7125 C32_U.n136 C32_U.n135 0.593536
R7126 C32_U.n141 C32_U.n140 0.465844
R7127 C32_U.n107 C32_U.n106 0.331311
R7128 C32_U.n108 C32_U.n107 0.331311
R7129 C32_U.n109 C32_U.n108 0.331311
R7130 C32_U.n110 C32_U.n109 0.331311
R7131 C32_U.n111 C32_U.n110 0.331311
R7132 C32_U.n112 C32_U.n111 0.331311
R7133 C32_U.n113 C32_U.n112 0.331311
R7134 C32_U.n114 C32_U.n113 0.331311
R7135 C32_U.n115 C32_U.n114 0.331311
R7136 C32_U.n116 C32_U.n115 0.331311
R7137 C32_U.n117 C32_U.n116 0.331311
R7138 C32_U.n118 C32_U.n117 0.331311
R7139 C32_U.n119 C32_U.n118 0.331311
R7140 C32_U.n120 C32_U.n119 0.331311
R7141 C32_U.n106 C32_U.n105 0.259959
R7142 C32_U.n121 C32_U.n120 0.259959
R7143 C32_U.n61 C32_U.n60 0.0533261
R7144 C32_U.n34 C32_U.n33 0.049413
R7145 C32_U.n8 C32_U.n7 0.0234787
R7146 C32_U.n64 C32_U.n61 0.0161522
R7147 C32_U.n35 C32_U.n34 0.0102826
R7148 C32_U C32_U.n148 0.0075
R7149 C32_U.n138 C32_U.n8 0.0060102
R7150 C32_U.n38 C32_U.n35 0.0045
R7151 b2b b2b.n2 33.3766
R7152 b2b b2b.t5 19.4226
R7153 b2b.n0 b2b.t6 13.1296
R7154 b2b.n1 b2b.t3 10.5977
R7155 b2b.n0 b2b.t4 10.5411
R7156 b2b.n5 b2b.n3 9.44853
R7157 b2b.n5 b2b.n4 9.35588
R7158 b2b.n2 b2b.t2 9.19699
R7159 b2b.n1 b2b.n0 8.57376
R7160 b2b.n6 b2b 3.36483
R7161 b2b b2b.n6 2.25319
R7162 b2b.n2 b2b.n1 0.226273
R7163 b2b.n6 b2b.n5 0.00180435
R7164 SDc_1.n104 SDc_1.n103 4.5005
R7165 SDc_1.n88 SDc_1.n5 3.42922
R7166 SDc_1.n73 SDc_1.n13 3.42426
R7167 SDc_1.n112 SDc_1.n111 3.14063
R7168 SDc_1.n37 SDc_1.n36 3.01875
R7169 SDc_1.n41 SDc_1.n28 3.00463
R7170 SDc_1.n94 SDc_1.n3 3.00249
R7171 SDc_1.n38 SDc_1.n32 3.00075
R7172 SDc_1.n47 SDc_1.n26 3.00075
R7173 SDc_1.n62 SDc_1.n17 3.00062
R7174 SDc_1.n71 SDc_1.n15 2.99808
R7175 SDc_1.n59 SDc_1.n19 2.99741
R7176 SDc_1.n100 SDc_1.n1 2.9958
R7177 SDc_1.n79 SDc_1.n9 2.995
R7178 SDc_1.n85 SDc_1.n7 2.99139
R7179 SDc_1.n50 SDc_1.n21 2.9875
R7180 SDc_1.n120 SDc_1.n106 2.9875
R7181 SDc_1.n39 SDc_1.n30 2.93157
R7182 SDc_1.n34 SDc_1.n33 2.9022
R7183 SDc_1.n36 SDc_1.n35 2.90217
R7184 SDc_1.n7 SDc_1.n6 2.90216
R7185 SDc_1.n68 SDc_1.n67 2.90215
R7186 SDc_1.n3 SDc_1.n2 2.90213
R7187 SDc_1.n76 SDc_1.n75 2.90213
R7188 SDc_1.n117 SDc_1.n116 2.90211
R7189 SDc_1.n82 SDc_1.n81 2.90211
R7190 SDc_1.n11 SDc_1.n10 2.90211
R7191 SDc_1.n108 SDc_1.n107 2.90211
R7192 SDc_1.n32 SDc_1.n31 2.90211
R7193 SDc_1.n26 SDc_1.n25 2.90211
R7194 SDc_1.n17 SDc_1.n16 2.90209
R7195 SDc_1.n19 SDc_1.n18 2.90209
R7196 SDc_1.n1 SDc_1.n0 2.90209
R7197 SDc_1.n114 SDc_1.n113 2.8968
R7198 SDc_1.n43 SDc_1.n42 2.87834
R7199 SDc_1.n21 SDc_1.n20 2.87834
R7200 SDc_1.n106 SDc_1.n105 2.87834
R7201 SDc_1.n96 SDc_1.n95 2.87826
R7202 SDc_1.n90 SDc_1.n89 2.87826
R7203 SDc_1.n9 SDc_1.n8 2.87826
R7204 SDc_1.n28 SDc_1.n27 2.87826
R7205 SDc_1.n102 SDc_1.n101 2.87824
R7206 SDc_1.n15 SDc_1.n14 2.87824
R7207 SDc_1.n64 SDc_1.t22 2.7305
R7208 SDc_1.n64 SDc_1.n63 2.7305
R7209 SDc_1.n56 SDc_1.t47 2.7305
R7210 SDc_1.n56 SDc_1.n55 2.7305
R7211 SDc_1.n52 SDc_1.t17 2.7305
R7212 SDc_1.n52 SDc_1.n51 2.7305
R7213 SDc_1.n23 SDc_1.t41 2.7305
R7214 SDc_1.n23 SDc_1.n22 2.7305
R7215 SDc_1.n30 SDc_1.t48 2.7305
R7216 SDc_1.n30 SDc_1.n29 2.7305
R7217 SDc_1.n13 SDc_1.t45 2.7305
R7218 SDc_1.n13 SDc_1.n12 2.7305
R7219 SDc_1.n5 SDc_1.t7 2.7305
R7220 SDc_1.n5 SDc_1.n4 2.7305
R7221 SDc_1.n110 SDc_1.n109 2.678
R7222 SDc_1.n115 SDc_1.n108 2.51419
R7223 SDc_1.n37 SDc_1.n34 2.50516
R7224 SDc_1.n74 SDc_1.n11 2.50487
R7225 SDc_1.n102 SDc_1.t46 2.43827
R7226 SDc_1.n15 SDc_1.t15 2.43827
R7227 SDc_1.n28 SDc_1.t36 2.43825
R7228 SDc_1.n96 SDc_1.t14 2.43825
R7229 SDc_1.n90 SDc_1.t43 2.43825
R7230 SDc_1.n9 SDc_1.t30 2.43825
R7231 SDc_1.n43 SDc_1.t12 2.43818
R7232 SDc_1.n21 SDc_1.t44 2.43818
R7233 SDc_1.n106 SDc_1.t34 2.43818
R7234 SDc_1.n17 SDc_1.t50 2.40706
R7235 SDc_1.n19 SDc_1.t10 2.40706
R7236 SDc_1.n1 SDc_1.t9 2.40706
R7237 SDc_1.n108 SDc_1.t40 2.40704
R7238 SDc_1.n32 SDc_1.t11 2.40704
R7239 SDc_1.n26 SDc_1.t5 2.40704
R7240 SDc_1.n117 SDc_1.t8 2.40704
R7241 SDc_1.n82 SDc_1.t13 2.40704
R7242 SDc_1.n11 SDc_1.t18 2.40704
R7243 SDc_1.n76 SDc_1.t33 2.40703
R7244 SDc_1.n3 SDc_1.t39 2.40702
R7245 SDc_1.n68 SDc_1.t49 2.40701
R7246 SDc_1.n36 SDc_1.t42 2.407
R7247 SDc_1.n7 SDc_1.t38 2.407
R7248 SDc_1.n34 SDc_1.t16 2.40696
R7249 SDc_1.n58 SDc_1.n57 2.24993
R7250 SDc_1.n70 SDc_1.n69 2.24993
R7251 SDc_1.n84 SDc_1.n83 2.24993
R7252 SDc_1.n78 SDc_1.n77 2.24966
R7253 SDc_1.n45 SDc_1.n44 2.24539
R7254 SDc_1.n92 SDc_1.n91 2.24539
R7255 SDc_1.n98 SDc_1.n97 2.24539
R7256 SDc_1.n119 SDc_1.n118 2.24512
R7257 SDc_1.n54 SDc_1.n53 2.24486
R7258 SDc_1.n66 SDc_1.n65 2.24459
R7259 SDc_1.n113 SDc_1.t4 2.10341
R7260 SDc_1.n115 SDc_1.n114 1.98438
R7261 SDc_1.n48 SDc_1.n24 1.49518
R7262 SDc_1.n65 SDc_1.n64 1.43771
R7263 SDc_1.n57 SDc_1.n56 1.43737
R7264 SDc_1.n53 SDc_1.n52 1.43737
R7265 SDc_1.n24 SDc_1.n23 1.43737
R7266 SDc_1.n69 SDc_1.n68 1.01063
R7267 SDc_1.n77 SDc_1.n76 1.01049
R7268 SDc_1.n83 SDc_1.n82 1.01042
R7269 SDc_1.n118 SDc_1.n117 1.01042
R7270 SDc_1.n44 SDc_1.n43 1.00841
R7271 SDc_1.n91 SDc_1.n90 1.00788
R7272 SDc_1.n97 SDc_1.n96 1.00788
R7273 SDc_1.n103 SDc_1.n102 1.00774
R7274 SDc_1.n40 SDc_1.n39 0.607669
R7275 SDc_1.n78 SDc_1.n74 0.607459
R7276 SDc_1.n70 SDc_1.n66 0.604141
R7277 SDc_1.n58 SDc_1.n54 0.601465
R7278 SDc_1.n119 SDc_1.n115 0.60093
R7279 SDc_1.n38 SDc_1.n37 0.598744
R7280 SDc_1.n99 SDc_1.n98 0.597758
R7281 SDc_1.n93 SDc_1.n92 0.595615
R7282 SDc_1.n49 SDc_1.n48 0.594387
R7283 SDc_1.n87 SDc_1.n86 0.588179
R7284 SDc_1.n84 SDc_1.n80 0.586535
R7285 SDc_1.n122 SDc_1.n121 0.58175
R7286 SDc_1.n73 SDc_1.n72 0.580143
R7287 SDc_1.n61 SDc_1.n60 0.570963
R7288 SDc_1.n46 SDc_1.n45 0.564543
R7289 SDc_1.n111 SDc_1.n110 0.053
R7290 SDc_1.n112 SDc_1 0.0505538
R7291 SDc_1.n47 SDc_1.n46 0.0251429
R7292 SDc_1.n60 SDc_1.n59 0.0240714
R7293 SDc_1.n72 SDc_1.n71 0.023
R7294 SDc_1.n80 SDc_1.n79 0.023
R7295 SDc_1.n86 SDc_1.n85 0.023
R7296 SDc_1.n114 SDc_1.n112 0.022869
R7297 SDc_1 SDc_1.n122 0.0219286
R7298 SDc_1.n74 SDc_1.n73 0.017366
R7299 SDc_1.n62 SDc_1.n61 0.0159634
R7300 SDc_1.n50 SDc_1.n49 0.0154306
R7301 SDc_1.n120 SDc_1.n119 0.0148978
R7302 SDc_1.n39 SDc_1.n38 0.0145059
R7303 SDc_1.n45 SDc_1.n41 0.0143648
R7304 SDc_1.n92 SDc_1.n88 0.0143648
R7305 SDc_1.n54 SDc_1.n50 0.0143592
R7306 SDc_1.n66 SDc_1.n62 0.0138205
R7307 SDc_1.n98 SDc_1.n94 0.0132934
R7308 SDc_1.n48 SDc_1.n47 0.011654
R7309 SDc_1.n100 SDc_1.n99 0.00585714
R7310 SDc_1.n41 SDc_1.n40 0.00478571
R7311 SDc_1.n88 SDc_1.n87 0.00478571
R7312 SDc_1.n94 SDc_1.n93 0.00478571
R7313 SDc_1.n79 SDc_1.n78 0.00474841
R7314 SDc_1.n59 SDc_1.n58 0.00421327
R7315 SDc_1.n71 SDc_1.n70 0.00421327
R7316 SDc_1.n85 SDc_1.n84 0.00421327
R7317 SDc_1.n121 SDc_1.n120 0.00264286
R7318 SDc_1.n104 SDc_1.n100 0.00157143
R7319 SDc_1 SDc_1.n104 0.00157143
R7320 ITAIL.n22 ITAIL.n6 333.663
R7321 ITAIL.n18 ITAIL.t22 116.817
R7322 ITAIL.n20 ITAIL.n19 103.823
R7323 ITAIL.n2 ITAIL.t17 97.648
R7324 ITAIL.n6 ITAIL.n5 90.8936
R7325 ITAIL.n22 ITAIL.n21 88.6306
R7326 ITAIL.n4 ITAIL.n3 84.9459
R7327 ITAIL.n19 ITAIL.n18 48.8699
R7328 ITAIL.n21 ITAIL.n20 47.0449
R7329 ITAIL.n3 ITAIL.n2 38.4914
R7330 ITAIL.n5 ITAIL.n4 38.4914
R7331 ITAIL.n17 ITAIL.n16 27.9195
R7332 ITAIL ITAIL.t15 27.414
R7333 ITAIL.t17 ITAIL.t11 23.7985
R7334 ITAIL.t4 ITAIL.t24 23.7985
R7335 ITAIL.t20 ITAIL.t14 23.7985
R7336 ITAIL.t2 ITAIL.t21 23.7985
R7337 ITAIL.t10 ITAIL.t6 23.7985
R7338 ITAIL.t23 ITAIL.t19 23.7985
R7339 ITAIL.t7 ITAIL.t3 23.7985
R7340 ITAIL.t16 ITAIL.t9 23.7985
R7341 ITAIL.t8 ITAIL.t5 23.7985
R7342 ITAIL.n21 ITAIL.t23 12.9945
R7343 ITAIL.n20 ITAIL.t7 12.9945
R7344 ITAIL.n19 ITAIL.t16 12.9945
R7345 ITAIL.n18 ITAIL.t8 12.9945
R7346 ITAIL.t15 ITAIL.n22 12.7755
R7347 ITAIL.n2 ITAIL.t4 12.7025
R7348 ITAIL.n3 ITAIL.t20 12.7025
R7349 ITAIL.n4 ITAIL.t2 12.7025
R7350 ITAIL.n5 ITAIL.t10 12.7025
R7351 ITAIL.n6 ITAIL.t12 10.8045
R7352 ITAIL.n1 ITAIL.t1 10.1411
R7353 ITAIL.n0 ITAIL.t0 8.6875
R7354 ITAIL.n17 ITAIL.t18 8.3955
R7355 ITAIL.t22 ITAIL.n17 8.1035
R7356 ITAIL.n0 ITAIL.t13 7.3735
R7357 ITAIL ITAIL.n1 4.95899
R7358 ITAIL.n1 ITAIL.n0 2.47975
R7359 ITAIL.n8 ITAIL 1.57458
R7360 ITAIL.n15 ITAIL.n14 0.656661
R7361 ITAIL.n16 ITAIL.n15 0.645581
R7362 ITAIL.n9 ITAIL.n8 0.642688
R7363 ITAIL.n11 ITAIL.n10 0.0405512
R7364 ITAIL.n14 ITAIL.n13 0.0405512
R7365 ITAIL.n15 ITAIL.n12 0.0121407
R7366 ITAIL.n10 ITAIL.n9 0.0117788
R7367 ITAIL.n16 ITAIL.n7 0.0103977
R7368 ITAIL.n12 ITAIL.n11 0.00211125
R7369 B1 B1.t0 48.6474
R7370 B1.n0 B1.t1 19.0247
R7371 B1.n0 B1.t2 17.3935
R7372 B1.n1 B1.n0 4.12942
R7373 B1.n1 B1 2.25699
R7374 B1 B1.n1 0.0067069
R7375 b1b b1b.n5 37.091
R7376 b1b.n3 b1b.t2 26.9594
R7377 b1b b1b.t3 19.4226
R7378 b1b.n5 b1b.n2 9.59479
R7379 b1b.n7 b1b.n0 9.49418
R7380 b1b.n6 b1b.n1 9.39109
R7381 b1b.n4 b1b.n3 7.55447
R7382 b1b.n3 b1b.n2 4.95899
R7383 b1b.n6 b1b 3.31968
R7384 b1b.t4 b1b.n2 2.79883
R7385 b1b b1b.n7 2.25319
R7386 b1b.n5 b1b.n4 1.68928
R7387 b1b.n4 b1b.t4 0.678302
R7388 b1b.n7 b1b.n6 0.00963044
R7389 SDn_1.n38 SDn_1.n35 4.73161
R7390 SDn_1.n34 SDn_1.n33 3.08659
R7391 SDn_1.n41 SDn_1.n40 3.04854
R7392 SDn_1.n25 SDn_1.n10 3.04726
R7393 SDn_1.n17 SDn_1.n16 3.04688
R7394 SDn_1.n52 SDn_1.n6 3.04375
R7395 SDn_1.n43 SDn_1.n8 3.04171
R7396 SDn_1.n19 SDn_1.n12 3.03541
R7397 SDn_1.n40 SDn_1.n39 2.9021
R7398 SDn_1.n4 SDn_1.t1 2.7305
R7399 SDn_1.n4 SDn_1.n3 2.7305
R7400 SDn_1.n49 SDn_1.t17 2.7305
R7401 SDn_1.n49 SDn_1.n48 2.7305
R7402 SDn_1.n45 SDn_1.t7 2.7305
R7403 SDn_1.n45 SDn_1.n44 2.7305
R7404 SDn_1.n37 SDn_1.t29 2.7305
R7405 SDn_1.n37 SDn_1.n36 2.7305
R7406 SDn_1.n31 SDn_1.t0 2.7305
R7407 SDn_1.n31 SDn_1.n30 2.7305
R7408 SDn_1.n27 SDn_1.t28 2.7305
R7409 SDn_1.n27 SDn_1.n26 2.7305
R7410 SDn_1.n21 SDn_1.t3 2.7305
R7411 SDn_1.n21 SDn_1.n20 2.7305
R7412 SDn_1.n14 SDn_1.t16 2.7305
R7413 SDn_1.n14 SDn_1.n13 2.7305
R7414 SDn_1.n16 SDn_1.t6 2.7305
R7415 SDn_1.n16 SDn_1.n15 2.7305
R7416 SDn_1.n12 SDn_1.t27 2.7305
R7417 SDn_1.n12 SDn_1.n11 2.7305
R7418 SDn_1.n10 SDn_1.t11 2.7305
R7419 SDn_1.n10 SDn_1.n9 2.7305
R7420 SDn_1.n33 SDn_1.t31 2.7305
R7421 SDn_1.n33 SDn_1.n32 2.7305
R7422 SDn_1.n8 SDn_1.t26 2.7305
R7423 SDn_1.n8 SDn_1.n7 2.7305
R7424 SDn_1.n6 SDn_1.t9 2.7305
R7425 SDn_1.n6 SDn_1.n5 2.7305
R7426 SDn_1.n1 SDn_1.t18 2.7305
R7427 SDn_1.n1 SDn_1.n0 2.7305
R7428 SDn_1.n17 SDn_1.n14 2.56247
R7429 SDn_1.n38 SDn_1.n37 2.56221
R7430 SDn_1.n34 SDn_1.n31 2.562
R7431 SDn_1.n54 SDn_1.n4 2.55991
R7432 SDn_1.n40 SDn_1.t8 2.40706
R7433 SDn_1.n51 SDn_1.n50 1.49447
R7434 SDn_1.n23 SDn_1.n22 1.49447
R7435 SDn_1.n29 SDn_1.n28 1.49423
R7436 SDn_1.n47 SDn_1.n46 1.49423
R7437 SDn_1.n50 SDn_1.n49 1.43787
R7438 SDn_1.n28 SDn_1.n27 1.43765
R7439 SDn_1.n46 SDn_1.n45 1.43732
R7440 SDn_1.n22 SDn_1.n21 1.437
R7441 SDn_1.n2 SDn_1.n1 1.4264
R7442 SDn_1.n55 SDn_1.n2 1.14083
R7443 SDn_1.n51 SDn_1.n47 0.58072
R7444 SDn_1.n18 SDn_1.n17 0.575838
R7445 SDn_1.n24 SDn_1.n23 0.574178
R7446 SDn_1.n54 SDn_1.n53 0.566624
R7447 SDn_1.n35 SDn_1.n29 0.554675
R7448 SDn_1.n42 SDn_1.n41 0.513212
R7449 SDn_1.n55 SDn_1.n54 0.482617
R7450 SDn_1.n2 SDn_1 0.157421
R7451 SDn_1.n19 SDn_1.n18 0.0271667
R7452 SDn_1.n53 SDn_1.n52 0.0249444
R7453 SDn_1.n47 SDn_1.n43 0.0212506
R7454 SDn_1.n25 SDn_1.n24 0.0205
R7455 SDn_1.n29 SDn_1.n25 0.0201395
R7456 SDn_1.n43 SDn_1.n42 0.0193889
R7457 SDn_1.n52 SDn_1.n51 0.0153623
R7458 SDn_1.n23 SDn_1.n19 0.0134755
R7459 SDn_1.n35 SDn_1.n34 0.0132059
R7460 SDn_1 SDn_1.n55 0.00682738
R7461 SDn_1.n41 SDn_1.n38 0.00579412
R7462 b3.t8 b3.t2 102.266
R7463 b3.n0 b3.t4 49.5502
R7464 b3 b3.t5 34.9792
R7465 b3.t9 b3.t7 28.703
R7466 b3.t10 b3.t6 26.4242
R7467 b3.t2 b3.t9 22.0465
R7468 b3.t6 b3.t8 22.0465
R7469 b3.t7 b3.t3 17.6665
R7470 b3.t5 b3.t10 17.6665
R7471 b3.n1 b3.t0 9.49371
R7472 b3.n1 b3.t1 9.3756
R7473 b3 b3.n1 3.6563
R7474 b3.n0 b3 3.36711
R7475 b3 b3.n0 2.25981
R7476 OUT3.n14 OUT3.n10 19.1949
R7477 OUT3.n13 OUT3.n11 6.45579
R7478 OUT3.n15 OUT3.n14 6.06989
R7479 OUT3.n13 OUT3.n12 5.8805
R7480 OUT3.n16 OUT3.t2 5.8805
R7481 OUT3.n15 OUT3.t3 5.8805
R7482 OUT3.n4 OUT3.n1 3.63586
R7483 OUT3.n9 OUT3.n6 3.63586
R7484 OUT3.n4 OUT3.n3 3.1505
R7485 OUT3.n9 OUT3.n8 3.1505
R7486 OUT3.n1 OUT3.t6 2.7305
R7487 OUT3.n1 OUT3.n0 2.7305
R7488 OUT3.n3 OUT3.t9 2.7305
R7489 OUT3.n3 OUT3.n2 2.7305
R7490 OUT3.n6 OUT3.t11 2.7305
R7491 OUT3.n6 OUT3.n5 2.7305
R7492 OUT3.n8 OUT3.t1 2.7305
R7493 OUT3.n8 OUT3.n7 2.7305
R7494 OUT3.n14 OUT3 2.39886
R7495 OUT3.n10 OUT3.n4 0.804767
R7496 OUT3.n16 OUT3.n15 0.564731
R7497 OUT3 OUT3.n13 0.199912
R7498 OUT3.n10 OUT3.n9 0.190191
R7499 OUT3 OUT3.n16 0.0558846
R7500 b4.n3 b4.n0 485.19
R7501 b4.n7 b4.n6 79.2611
R7502 b4.n1 b4.t10 65.6295
R7503 b4.n5 b4.t8 64.5576
R7504 b4.t13 b4.t15 62.9752
R7505 b4.t7 b4.n7 62.5658
R7506 b4.n10 b4.t12 51.8002
R7507 b4.t16 b4.t13 41.6538
R7508 b4.t17 b4.t9 32.3937
R7509 b4.t8 b4.t2 20.3675
R7510 b4.t5 b4.t16 20.3675
R7511 b4.n6 b4.n5 20.0889
R7512 b4.t18 b4.t6 18.2505
R7513 b4 b4.n9 17.3009
R7514 b4.t10 b4.t3 16.0605
R7515 b4.n8 b4.t14 15.7355
R7516 b4.n6 b4.t5 13.8705
R7517 b4.n4 b4.t4 13.2149
R7518 b4.n8 b4.t7 10.1176
R7519 b4.n5 b4.t17 10.0015
R7520 b4.n11 b4.t1 9.49371
R7521 b4.n11 b4.t0 9.3756
R7522 b4.n2 b4.n1 8.61736
R7523 b4.n4 b4.n3 8.26992
R7524 b4.n9 b4.n8 5.77524
R7525 b4.n7 b4.t18 5.4025
R7526 b4.n3 b4.n2 4.86717
R7527 b4.n9 b4.n4 4.43773
R7528 b4 b4.n11 3.6563
R7529 b4.n1 b4.n0 2.03842
R7530 b4.t11 b4.n0 1.91942
R7531 b4.n2 b4.t11 0.122167
R7532 b4 b4.n10 0.00981034
R7533 b4.n10 b4 0.00256897
R7534 SD2_1 SD2_1.n20 9.24575
R7535 SD2_1.n19 SD2_1.n18 3.45039
R7536 SD2_1.n14 SD2_1.n13 3.44985
R7537 SD2_1.n9 SD2_1.n8 3.44969
R7538 SD2_1.n4 SD2_1.n3 3.44925
R7539 SD2_1.n14 SD2_1.n11 3.4367
R7540 SD2_1.n19 SD2_1.n16 3.43615
R7541 SD2_1.n4 SD2_1.n1 3.43133
R7542 SD2_1 SD2_1.n6 3.3305
R7543 SD2_1.n20 SD2_1.n19 2.87896
R7544 SD2_1 SD2_1.n4 2.8298
R7545 SD2_1.n6 SD2_1.t6 2.7305
R7546 SD2_1.n6 SD2_1.n5 2.7305
R7547 SD2_1.n11 SD2_1.t9 2.7305
R7548 SD2_1.n11 SD2_1.n10 2.7305
R7549 SD2_1.n13 SD2_1.t11 2.7305
R7550 SD2_1.n13 SD2_1.n12 2.7305
R7551 SD2_1.n16 SD2_1.t4 2.7305
R7552 SD2_1.n16 SD2_1.n15 2.7305
R7553 SD2_1.n18 SD2_1.t5 2.7305
R7554 SD2_1.n18 SD2_1.n17 2.7305
R7555 SD2_1.n1 SD2_1.t12 2.7305
R7556 SD2_1.n1 SD2_1.n0 2.7305
R7557 SD2_1.n3 SD2_1.t13 2.7305
R7558 SD2_1.n3 SD2_1.n2 2.7305
R7559 SD2_1.n8 SD2_1.t7 2.7305
R7560 SD2_1.n8 SD2_1.n7 2.7305
R7561 SD2_1.n20 SD2_1.n14 2.25147
R7562 SD2_1 SD2_1.n9 2.2505
R7563 SD2_1.n9 SD2_1 0.100126
R7564 G1_2.n6 G1_2.n2 147.578
R7565 G1_2.n17 G1_2.n16 142.844
R7566 G1_2.n15 G1_2.n14 101.016
R7567 G1_2.n1 G1_2.n0 101.016
R7568 G1_2.n5 G1_2.n4 101.016
R7569 G1_2.n13 G1_2.n12 101.016
R7570 G1_2.n14 G1_2.t29 33.5864
R7571 G1_2.n0 G1_2.t31 33.5864
R7572 G1_2.n16 G1_2.n15 20.5194
R7573 G1_2.n2 G1_2.n1 20.5194
R7574 G1_2.n6 G1_2.n5 20.5194
R7575 G1_2.n4 G1_2.n3 20.5194
R7576 G1_2.n12 G1_2.n11 20.5194
R7577 G1_2.n17 G1_2.n13 20.5194
R7578 G1_2.n14 G1_2.t34 13.0675
R7579 G1_2.n15 G1_2.t30 13.0675
R7580 G1_2.n16 G1_2.t32 13.0675
R7581 G1_2.n0 G1_2.t26 13.0675
R7582 G1_2.n1 G1_2.t24 13.0675
R7583 G1_2.n2 G1_2.t28 13.0675
R7584 G1_2.n5 G1_2.t12 13.0675
R7585 G1_2.n4 G1_2.t8 13.0675
R7586 G1_2.n3 G1_2.t10 13.0675
R7587 G1_2.n11 G1_2.t22 13.0675
R7588 G1_2.n12 G1_2.t14 13.0675
R7589 G1_2.n13 G1_2.t18 13.0675
R7590 G1_2.n9 G1_2.t16 8.3225
R7591 G1_2.n47 G1_2.t20 8.1765
R7592 G1_2.n43 G1_2.n41 6.51833
R7593 G1_2.n37 G1_2.t7 6.51833
R7594 G1_2.n45 G1_2.t1 5.8805
R7595 G1_2.n44 G1_2.t2 5.8805
R7596 G1_2.n43 G1_2.n42 5.8805
R7597 G1_2.n39 G1_2.n35 5.8805
R7598 G1_2.n38 G1_2.n36 5.8805
R7599 G1_2.n37 G1_2.t0 5.8805
R7600 G1_2.n46 G1_2.n45 5.81863
R7601 G1_2.n40 G1_2.n39 5.52662
R7602 G1_2.n49 G1_2.n48 4.5005
R7603 G1_2.n46 G1_2.n40 4.28996
R7604 G1_2.n8 G1_2.n7 3.53359
R7605 G1_2.n33 G1_2.n18 3.50535
R7606 G1_2.n20 G1_2.t17 3.03383
R7607 G1_2.n20 G1_2.n19 3.03383
R7608 G1_2.n22 G1_2.t15 3.03383
R7609 G1_2.n22 G1_2.n21 3.03383
R7610 G1_2.n24 G1_2.t11 3.03383
R7611 G1_2.n24 G1_2.n23 3.03383
R7612 G1_2.n26 G1_2.t13 3.03383
R7613 G1_2.n26 G1_2.n25 3.03383
R7614 G1_2.n34 G1_2.n10 2.88425
R7615 G1_2.n30 G1_2.n22 2.8392
R7616 G1_2.n29 G1_2.n24 2.8392
R7617 G1_2.n31 G1_2.n20 2.80007
R7618 G1_2.n28 G1_2.n26 2.80007
R7619 G1_2.n40 G1_2.n34 2.5439
R7620 G1_2.n10 G1_2.n9 2.1905
R7621 G1_2.n44 G1_2.n43 2.07441
R7622 G1_2.n48 G1_2.n47 2.0445
R7623 G1_2.n38 G1_2.n37 2.0118
R7624 G1_2.n49 G1_2.n46 1.80063
R7625 G1_2.n30 G1_2.n29 1.59702
R7626 G1_2.n31 G1_2.n30 1.58339
R7627 G1_2.n29 G1_2.n28 1.58339
R7628 G1_2.n7 G1_2.n6 1.15481
R7629 G1_2.n18 G1_2.n17 1.06529
R7630 G1_2.n45 G1_2.n44 0.638326
R7631 G1_2.n39 G1_2.n38 0.638326
R7632 G1_2.n32 G1_2.n31 0.0932273
R7633 G1_2 G1_2.n27 0.0876818
R7634 G1_2.n33 G1_2.n32 0.0305
R7635 G1_2.n27 G1_2.n8 0.0265
R7636 G1_2.n28 G1_2 0.0100455
R7637 G1_2 G1_2.n8 0.0085
R7638 G1_2.n34 G1_2.n33 0.0055
R7639 G1_2 G1_2.n49 0.0025
R7640 SD1_1.n15 SD1_1.n14 7.78572
R7641 SD1_1.n9 SD1_1.n8 3.20235
R7642 SD1_1.n17 SD1_1.n16 3.17681
R7643 SD1_1.n1 SD1_1.t3 3.03383
R7644 SD1_1.n1 SD1_1.n0 3.03383
R7645 SD1_1.n22 SD1_1.t13 3.03383
R7646 SD1_1.n22 SD1_1.n21 3.03383
R7647 SD1_1.n19 SD1_1.t14 3.03383
R7648 SD1_1.n19 SD1_1.n18 3.03383
R7649 SD1_1.n13 SD1_1.t7 3.03383
R7650 SD1_1.n13 SD1_1.n12 3.03383
R7651 SD1_1.n5 SD1_1.t5 3.03383
R7652 SD1_1.n5 SD1_1.n4 3.03383
R7653 SD1_1.n7 SD1_1.t6 3.03383
R7654 SD1_1.n7 SD1_1.n6 3.03383
R7655 SD1_1.n20 SD1_1.n17 2.97146
R7656 SD1_1.n10 SD1_1.n9 2.94829
R7657 SD1_1.n10 SD1_1.n7 2.75112
R7658 SD1_1.n17 SD1_1.t8 2.69498
R7659 SD1_1.n9 SD1_1.t2 2.66057
R7660 SD1_1.n14 SD1_1.n13 2.38615
R7661 SD1_1.n23 SD1_1.n22 2.37424
R7662 SD1_1.n20 SD1_1.n19 2.37412
R7663 SD1_1.n11 SD1_1.n5 2.37207
R7664 SD1_1.n2 SD1_1.n1 1.63787
R7665 SD1_1.n15 SD1_1.n3 1.12886
R7666 SD1_1.n23 SD1_1.n20 0.626727
R7667 SD1_1.n11 SD1_1.n10 0.613463
R7668 SD1_1.n14 SD1_1.n11 0.609042
R7669 SD1_1.n24 SD1_1.n23 0.584266
R7670 SD1_1.n2 SD1_1 0.0568907
R7671 SD1_1 SD1_1.n24 0.0265
R7672 SD1_1.n3 SD1_1.n2 0.0213805
R7673 SD1_1 SD1_1.n15 0.00686644
R7674 SD2_4.n10 SD2_4.n4 5.11704
R7675 SD2_4.n4 SD2_4.n1 3.44424
R7676 SD2_4.n9 SD2_4.n8 3.37323
R7677 SD2_4.n4 SD2_4.n3 3.33687
R7678 SD2_4 SD2_4.n6 3.31692
R7679 SD2_4.n6 SD2_4.t6 2.7305
R7680 SD2_4.n6 SD2_4.n5 2.7305
R7681 SD2_4.n1 SD2_4.t2 2.7305
R7682 SD2_4.n1 SD2_4.n0 2.7305
R7683 SD2_4.n3 SD2_4.t3 2.7305
R7684 SD2_4.n3 SD2_4.n2 2.7305
R7685 SD2_4.n8 SD2_4.t7 2.7305
R7686 SD2_4.n8 SD2_4.n7 2.7305
R7687 SD2_4.n10 SD2_4.n9 2.2505
R7688 SD2_4.n9 SD2_4 0.116226
R7689 SD2_4 SD2_4.n10 0.00261765
R7690 G1_1.n27 G1_1.t24 113.573
R7691 G1_1.n17 G1_1.t28 113.573
R7692 G1_1.n29 G1_1.n28 101.016
R7693 G1_1.n19 G1_1.n18 101.016
R7694 G1_1.n21 G1_1.n20 101.016
R7695 G1_1.n23 G1_1.n22 101.016
R7696 G1_1.n25 G1_1.n24 101.016
R7697 G1_1.n30 G1_1.n26 101.016
R7698 G1_1.n20 G1_1.n19 67.0816
R7699 G1_1.n30 G1_1.n29 62.3464
R7700 G1_1.n28 G1_1.n27 20.5194
R7701 G1_1.n18 G1_1.n17 20.5194
R7702 G1_1.n22 G1_1.n21 20.5194
R7703 G1_1.n24 G1_1.n23 20.5194
R7704 G1_1.n26 G1_1.n25 20.5194
R7705 G1_1.n27 G1_1.t30 12.5565
R7706 G1_1.n28 G1_1.t35 12.5565
R7707 G1_1.n29 G1_1.t25 12.5565
R7708 G1_1.n17 G1_1.t29 12.5565
R7709 G1_1.n18 G1_1.t34 12.5565
R7710 G1_1.n19 G1_1.t32 12.5565
R7711 G1_1.n21 G1_1.t14 12.5565
R7712 G1_1.n22 G1_1.t4 12.5565
R7713 G1_1.n23 G1_1.t8 12.5565
R7714 G1_1.n24 G1_1.t0 12.5565
R7715 G1_1.n25 G1_1.t2 12.5565
R7716 G1_1.n26 G1_1.t10 12.5565
R7717 G1_1.n0 G1_1.t12 10.2935
R7718 G1_1.n31 G1_1.t6 10.2935
R7719 G1_1.n32 G1_1.n31 4.12693
R7720 G1_1 G1_1.n0 4.0015
R7721 G1_1.n2 G1_1.t21 3.03383
R7722 G1_1.n2 G1_1.n1 3.03383
R7723 G1_1.n16 G1_1.t7 3.03383
R7724 G1_1.n16 G1_1.n15 3.03383
R7725 G1_1.n4 G1_1.t15 3.03383
R7726 G1_1.n4 G1_1.n3 3.03383
R7727 G1_1.n6 G1_1.t16 3.03383
R7728 G1_1.n6 G1_1.n5 3.03383
R7729 G1_1.n8 G1_1.t9 3.03383
R7730 G1_1.n8 G1_1.n7 3.03383
R7731 G1_1.n10 G1_1.t22 3.03383
R7732 G1_1.n10 G1_1.n9 3.03383
R7733 G1_1.n12 G1_1.t3 3.03383
R7734 G1_1.n12 G1_1.n11 3.03383
R7735 G1_1.n14 G1_1.t18 3.03383
R7736 G1_1.n14 G1_1.n13 3.03383
R7737 G1_1.n38 G1_1.n4 2.82159
R7738 G1_1.n37 G1_1.n6 2.82159
R7739 G1_1.n36 G1_1.n8 2.82159
R7740 G1_1.n35 G1_1.n10 2.82159
R7741 G1_1.n34 G1_1.n12 2.82159
R7742 G1_1.n33 G1_1.n14 2.82159
R7743 G1_1.n39 G1_1.n2 2.78833
R7744 G1_1.n32 G1_1.n16 2.78833
R7745 G1_1.n20 G1_1.n0 2.2635
R7746 G1_1.n31 G1_1.n30 2.2635
R7747 G1_1.n34 G1_1.n33 0.798761
R7748 G1_1.n35 G1_1.n34 0.798761
R7749 G1_1.n36 G1_1.n35 0.798761
R7750 G1_1.n37 G1_1.n36 0.798761
R7751 G1_1.n38 G1_1.n37 0.798761
R7752 G1_1.n33 G1_1.n32 0.786618
R7753 G1_1 G1_1.n38 0.626587
R7754 G1_1.n39 G1_1 0.160531
R7755 G1_1 G1_1.n39 0.0949286
R7756 C32_D.n183 C32_D.t2 34.1564
R7757 C32_D.n184 C32_D.t28 12.0455
R7758 C32_D.n139 C32_D.t6 12.0455
R7759 C32_D.n136 C32_D.t4 12.0455
R7760 C32_D.n119 C32_D.t58 12.0455
R7761 C32_D.n116 C32_D.t14 12.0455
R7762 C32_D.n99 C32_D.t60 12.0455
R7763 C32_D.n96 C32_D.t52 12.0455
R7764 C32_D.n79 C32_D.t16 12.0455
R7765 C32_D.n76 C32_D.t18 12.0455
R7766 C32_D.n59 C32_D.t48 12.0455
R7767 C32_D.n56 C32_D.t10 12.0455
R7768 C32_D.n39 C32_D.t38 12.0455
R7769 C32_D.n36 C32_D.t42 12.0455
R7770 C32_D.n159 C32_D.t0 11.5345
R7771 C32_D.n156 C32_D.t32 10.8775
R7772 C32_D.n169 C32_D.t54 10.7315
R7773 C32_D.n166 C32_D.t8 10.7315
R7774 C32_D.n146 C32_D.t56 10.7315
R7775 C32_D.n129 C32_D.t44 10.7315
R7776 C32_D.n126 C32_D.t36 10.7315
R7777 C32_D.n109 C32_D.t22 10.7315
R7778 C32_D.n106 C32_D.t62 10.7315
R7779 C32_D.n89 C32_D.t24 10.7315
R7780 C32_D.n86 C32_D.t30 10.7315
R7781 C32_D.n69 C32_D.t46 10.7315
R7782 C32_D.n66 C32_D.t50 10.7315
R7783 C32_D.n49 C32_D.t20 10.7315
R7784 C32_D.n46 C32_D.t40 10.7315
R7785 C32_D.n28 C32_D.t12 10.7315
R7786 C32_D.n149 C32_D.t34 10.5125
R7787 C32_D.n180 C32_D.t26 9.5635
R7788 C32_D.n179 C32_D 5.27919
R7789 C32_D.n31 C32_D.n28 4.05396
R7790 C32_D.n185 C32_D.n184 4.0005
R7791 C32_D.n37 C32_D.n36 4.0005
R7792 C32_D.n40 C32_D.n39 4.0005
R7793 C32_D.n47 C32_D.n46 4.0005
R7794 C32_D.n50 C32_D.n49 4.0005
R7795 C32_D.n57 C32_D.n56 4.0005
R7796 C32_D.n60 C32_D.n59 4.0005
R7797 C32_D.n67 C32_D.n66 4.0005
R7798 C32_D.n70 C32_D.n69 4.0005
R7799 C32_D.n77 C32_D.n76 4.0005
R7800 C32_D.n80 C32_D.n79 4.0005
R7801 C32_D.n87 C32_D.n86 4.0005
R7802 C32_D.n90 C32_D.n89 4.0005
R7803 C32_D.n97 C32_D.n96 4.0005
R7804 C32_D.n100 C32_D.n99 4.0005
R7805 C32_D.n107 C32_D.n106 4.0005
R7806 C32_D.n110 C32_D.n109 4.0005
R7807 C32_D.n117 C32_D.n116 4.0005
R7808 C32_D.n120 C32_D.n119 4.0005
R7809 C32_D.n127 C32_D.n126 4.0005
R7810 C32_D.n130 C32_D.n129 4.0005
R7811 C32_D.n137 C32_D.n136 4.0005
R7812 C32_D.n140 C32_D.n139 4.0005
R7813 C32_D.n147 C32_D.n146 4.0005
R7814 C32_D.n150 C32_D.n149 4.0005
R7815 C32_D.n157 C32_D.n156 4.0005
R7816 C32_D.n160 C32_D.n159 4.0005
R7817 C32_D.n167 C32_D.n166 4.0005
R7818 C32_D.n170 C32_D.n169 4.0005
R7819 C32_D.n178 C32_D.n177 3.50928
R7820 C32_D.n156 C32_D.n155 3.5045
R7821 C32_D.n31 C32_D.n30 3.48115
R7822 C32_D.n190 C32_D.n187 3.47528
R7823 C32_D.n34 C32_D.n33 3.47333
R7824 C32_D.n43 C32_D.n42 3.40485
R7825 C32_D.n54 C32_D.n53 3.40485
R7826 C32_D.n63 C32_D.n62 3.40485
R7827 C32_D.n74 C32_D.n73 3.40485
R7828 C32_D.n83 C32_D.n82 3.40485
R7829 C32_D.n94 C32_D.n93 3.40485
R7830 C32_D.n103 C32_D.n102 3.40485
R7831 C32_D.n114 C32_D.n113 3.40485
R7832 C32_D.n123 C32_D.n122 3.40485
R7833 C32_D.n134 C32_D.n133 3.40485
R7834 C32_D.n143 C32_D.n142 3.40485
R7835 C32_D.n174 C32_D.n173 3.40485
R7836 C32_D.n163 C32_D.n162 3.39898
R7837 C32_D.n154 C32_D.n153 3.3892
R7838 C32_D.n190 C32_D.n189 3.38528
R7839 C32_D.n171 C32_D.n1 3.35007
R7840 C32_D.n131 C32_D.n9 3.35007
R7841 C32_D.n111 C32_D.n13 3.35007
R7842 C32_D.n91 C32_D.n17 3.35007
R7843 C32_D.n71 C32_D.n21 3.35007
R7844 C32_D.n51 C32_D.n25 3.35007
R7845 C32_D.n44 C32_D.n27 3.35007
R7846 C32_D.n64 C32_D.n23 3.35007
R7847 C32_D.n84 C32_D.n19 3.35007
R7848 C32_D.n104 C32_D.n15 3.35007
R7849 C32_D.n124 C32_D.n11 3.35007
R7850 C32_D.n144 C32_D.n7 3.35007
R7851 C32_D.n164 C32_D.n3 3.35007
R7852 C32_D.n151 C32_D.n5 3.3442
R7853 C32_D.n182 C32_D.n181 2.87342
R7854 C32_D.n159 C32_D.n158 2.8475
R7855 C32_D.n173 C32_D.t91 2.7305
R7856 C32_D.n173 C32_D.n172 2.7305
R7857 C32_D.n1 C32_D.t55 2.7305
R7858 C32_D.n1 C32_D.n0 2.7305
R7859 C32_D.n162 C32_D.t1 2.7305
R7860 C32_D.n162 C32_D.n161 2.7305
R7861 C32_D.n153 C32_D.t79 2.7305
R7862 C32_D.n153 C32_D.n152 2.7305
R7863 C32_D.n5 C32_D.t35 2.7305
R7864 C32_D.n5 C32_D.n4 2.7305
R7865 C32_D.n142 C32_D.t7 2.7305
R7866 C32_D.n142 C32_D.n141 2.7305
R7867 C32_D.n133 C32_D.t83 2.7305
R7868 C32_D.n133 C32_D.n132 2.7305
R7869 C32_D.n9 C32_D.t45 2.7305
R7870 C32_D.n9 C32_D.n8 2.7305
R7871 C32_D.n122 C32_D.t59 2.7305
R7872 C32_D.n122 C32_D.n121 2.7305
R7873 C32_D.n113 C32_D.t71 2.7305
R7874 C32_D.n113 C32_D.n112 2.7305
R7875 C32_D.n13 C32_D.t23 2.7305
R7876 C32_D.n13 C32_D.n12 2.7305
R7877 C32_D.n102 C32_D.t61 2.7305
R7878 C32_D.n102 C32_D.n101 2.7305
R7879 C32_D.n93 C32_D.t76 2.7305
R7880 C32_D.n93 C32_D.n92 2.7305
R7881 C32_D.n17 C32_D.t25 2.7305
R7882 C32_D.n17 C32_D.n16 2.7305
R7883 C32_D.n82 C32_D.t17 2.7305
R7884 C32_D.n82 C32_D.n81 2.7305
R7885 C32_D.n73 C32_D.t84 2.7305
R7886 C32_D.n73 C32_D.n72 2.7305
R7887 C32_D.n21 C32_D.t47 2.7305
R7888 C32_D.n21 C32_D.n20 2.7305
R7889 C32_D.n62 C32_D.t49 2.7305
R7890 C32_D.n62 C32_D.n61 2.7305
R7891 C32_D.n53 C32_D.t70 2.7305
R7892 C32_D.n53 C32_D.n52 2.7305
R7893 C32_D.n25 C32_D.t21 2.7305
R7894 C32_D.n25 C32_D.n24 2.7305
R7895 C32_D.n42 C32_D.t39 2.7305
R7896 C32_D.n42 C32_D.n41 2.7305
R7897 C32_D.n30 C32_D.t13 2.7305
R7898 C32_D.n30 C32_D.n29 2.7305
R7899 C32_D.n33 C32_D.t67 2.7305
R7900 C32_D.n33 C32_D.n32 2.7305
R7901 C32_D.n189 C32_D.t29 2.7305
R7902 C32_D.n189 C32_D.n188 2.7305
R7903 C32_D.n187 C32_D.t82 2.7305
R7904 C32_D.n187 C32_D.n186 2.7305
R7905 C32_D.n27 C32_D.t87 2.7305
R7906 C32_D.n27 C32_D.n26 2.7305
R7907 C32_D.n23 C32_D.t89 2.7305
R7908 C32_D.n23 C32_D.n22 2.7305
R7909 C32_D.n19 C32_D.t74 2.7305
R7910 C32_D.n19 C32_D.n18 2.7305
R7911 C32_D.n15 C32_D.t95 2.7305
R7912 C32_D.n15 C32_D.n14 2.7305
R7913 C32_D.n11 C32_D.t93 2.7305
R7914 C32_D.n11 C32_D.n10 2.7305
R7915 C32_D.n7 C32_D.t69 2.7305
R7916 C32_D.n7 C32_D.n6 2.7305
R7917 C32_D.n3 C32_D.t66 2.7305
R7918 C32_D.n3 C32_D.n2 2.7305
R7919 C32_D.n149 C32_D.n148 2.5555
R7920 C32_D.n181 C32_D.n180 2.4095
R7921 C32_D.n184 C32_D.n183 2.3365
R7922 C32_D.n169 C32_D.n168 2.3365
R7923 C32_D.n166 C32_D.n165 2.3365
R7924 C32_D.n146 C32_D.n145 2.3365
R7925 C32_D.n139 C32_D.n138 2.3365
R7926 C32_D.n136 C32_D.n135 2.3365
R7927 C32_D.n129 C32_D.n128 2.3365
R7928 C32_D.n126 C32_D.n125 2.3365
R7929 C32_D.n119 C32_D.n118 2.3365
R7930 C32_D.n116 C32_D.n115 2.3365
R7931 C32_D.n109 C32_D.n108 2.3365
R7932 C32_D.n106 C32_D.n105 2.3365
R7933 C32_D.n99 C32_D.n98 2.3365
R7934 C32_D.n96 C32_D.n95 2.3365
R7935 C32_D.n89 C32_D.n88 2.3365
R7936 C32_D.n86 C32_D.n85 2.3365
R7937 C32_D.n79 C32_D.n78 2.3365
R7938 C32_D.n76 C32_D.n75 2.3365
R7939 C32_D.n69 C32_D.n68 2.3365
R7940 C32_D.n66 C32_D.n65 2.3365
R7941 C32_D.n59 C32_D.n58 2.3365
R7942 C32_D.n56 C32_D.n55 2.3365
R7943 C32_D.n49 C32_D.n48 2.3365
R7944 C32_D.n46 C32_D.n45 2.3365
R7945 C32_D.n39 C32_D.n38 2.3365
R7946 C32_D.n36 C32_D.n35 2.3365
R7947 C32_D.n177 C32_D.n176 1.02542
R7948 C32_D.n40 C32_D.n37 0.313543
R7949 C32_D.n60 C32_D.n57 0.313543
R7950 C32_D.n80 C32_D.n77 0.313543
R7951 C32_D.n100 C32_D.n97 0.313543
R7952 C32_D.n120 C32_D.n117 0.313543
R7953 C32_D.n140 C32_D.n137 0.313543
R7954 C32_D.n160 C32_D.n157 0.313543
R7955 C32_D.n185 C32_D.n182 0.301108
R7956 C32_D.n50 C32_D.n47 0.284446
R7957 C32_D.n70 C32_D.n67 0.284446
R7958 C32_D.n90 C32_D.n87 0.284446
R7959 C32_D.n110 C32_D.n107 0.284446
R7960 C32_D.n130 C32_D.n127 0.284446
R7961 C32_D.n170 C32_D.n167 0.284446
R7962 C32_D.n150 C32_D.n147 0.283774
R7963 C32_D C32_D.n190 0.1015
R7964 C32_D.n34 C32_D.n31 0.0826739
R7965 C32_D.n37 C32_D.n34 0.0795
R7966 C32_D.n43 C32_D.n40 0.0795
R7967 C32_D.n57 C32_D.n54 0.0795
R7968 C32_D.n63 C32_D.n60 0.0795
R7969 C32_D.n77 C32_D.n74 0.0795
R7970 C32_D.n83 C32_D.n80 0.0795
R7971 C32_D.n97 C32_D.n94 0.0795
R7972 C32_D.n103 C32_D.n100 0.0795
R7973 C32_D.n117 C32_D.n114 0.0795
R7974 C32_D.n123 C32_D.n120 0.0795
R7975 C32_D.n137 C32_D.n134 0.0795
R7976 C32_D.n143 C32_D.n140 0.0795
R7977 C32_D.n157 C32_D.n154 0.0795
R7978 C32_D.n163 C32_D.n160 0.0795
R7979 C32_D.n47 C32_D.n44 0.0695226
R7980 C32_D.n51 C32_D.n50 0.0695226
R7981 C32_D.n67 C32_D.n64 0.0695226
R7982 C32_D.n71 C32_D.n70 0.0695226
R7983 C32_D.n87 C32_D.n84 0.0695226
R7984 C32_D.n91 C32_D.n90 0.0695226
R7985 C32_D.n107 C32_D.n104 0.0695226
R7986 C32_D.n111 C32_D.n110 0.0695226
R7987 C32_D.n127 C32_D.n124 0.0695226
R7988 C32_D.n131 C32_D.n130 0.0695226
R7989 C32_D.n147 C32_D.n144 0.0695226
R7990 C32_D.n167 C32_D.n164 0.0695226
R7991 C32_D.n171 C32_D.n170 0.0695226
R7992 C32_D.n151 C32_D.n150 0.068
R7993 C32_D.n175 C32_D.n174 0.0465
R7994 C32_D.n178 C32_D.n175 0.0335
R7995 C32_D.n182 C32_D.n179 0.0128487
R7996 C32_D.n154 C32_D.n151 0.011299
R7997 C32_D.n164 C32_D.n163 0.0104247
R7998 C32_D.n44 C32_D.n43 0.00953213
R7999 C32_D.n54 C32_D.n51 0.00953213
R8000 C32_D.n64 C32_D.n63 0.00953213
R8001 C32_D.n74 C32_D.n71 0.00953213
R8002 C32_D.n84 C32_D.n83 0.00953213
R8003 C32_D.n94 C32_D.n91 0.00953213
R8004 C32_D.n104 C32_D.n103 0.00953213
R8005 C32_D.n114 C32_D.n111 0.00953213
R8006 C32_D.n124 C32_D.n123 0.00953213
R8007 C32_D.n134 C32_D.n131 0.00953213
R8008 C32_D.n144 C32_D.n143 0.00953213
R8009 C32_D.n174 C32_D.n171 0.00953213
R8010 C32_D C32_D.n185 0.0015
R8011 C32_D.n179 C32_D.n178 0.0015
R8012 B3 B3.t2 48.6474
R8013 B3.n0 B3.t1 19.0247
R8014 B3.n0 B3.t0 17.3935
R8015 B3.n1 B3.n0 4.12942
R8016 B3.n1 B3 2.25699
R8017 B3 B3.n1 0.0067069
R8018 b3b.n6 b3b.t3 36.6929
R8019 b3b.t5 b3b.t8 22.0465
R8020 b3b.t7 b3b.t10 22.0465
R8021 b3b.n6 b3b.t2 18.6988
R8022 b3b.t9 b3b.t4 17.6665
R8023 b3b.t3 b3b.t6 17.6665
R8024 b3b.n4 b3b.t5 12.209
R8025 b3b.n5 b3b.t7 12.0202
R8026 b3b.t6 b3b.n5 11.1473
R8027 b3b.n4 b3b.t9 10.8684
R8028 b3b.n1 b3b.n0 9.49288
R8029 b3b.n3 b3b.n2 9.40022
R8030 b3b.n5 b3b.n4 8.7605
R8031 b3b b3b.n3 2.25319
R8032 b3b b3b.n6 0.681545
R8033 b3b.n1 b3b 0.177597
R8034 b3b.n3 b3b.n1 0.00180435
R8035 OUT1 OUT1.n1 24.2283
R8036 OUT1 OUT1.t0 5.96093
R8037 OUT1.n1 OUT1.t1 2.7305
R8038 OUT1.n1 OUT1.n0 2.7305
R8039 SD2_3.n3 SD2_3.n2 6.50095
R8040 SD2_3.n2 SD2_3.n0 6.4673
R8041 SD2_3 SD2_3.t0 6.08127
R8042 SD2_3.n3 SD2_3.t2 5.8805
R8043 SD2_3.n2 SD2_3.n1 5.8805
R8044 SD2_3 SD2_3.n3 0.291269
R8045 b1.n4 b1.t3 50.6785
R8046 b1.n1 b1.n0 41.4888
R8047 b1 b1.n3 33.4868
R8048 b1.n1 b1.t2 17.9739
R8049 b1.n5 b1.t1 9.49371
R8050 b1.n5 b1.t0 9.3756
R8051 b1.n3 b1.n0 6.4245
R8052 b1.t4 b1.n0 4.50217
R8053 b1 b1.n5 3.6563
R8054 b1.n3 b1.n2 2.47632
R8055 b1.n2 b1.n1 1.66454
R8056 b1.n4 b1 0.858629
R8057 b1.n2 b1.t4 0.254192
R8058 b1 b1.n4 0.0800215
R8059 B5.n2 B5.t0 48.3651
R8060 B5.n0 B5.t1 19.0247
R8061 B5.n0 B5.t2 17.3935
R8062 B5.n2 B5 9.03551
R8063 B5.n1 B5.n0 4.12942
R8064 B5 B5.n1 2.25699
R8065 B5 B5.n2 0.273499
R8066 B5.n1 B5 0.0067069
R8067 B4 B4.t1 48.6474
R8068 B4.n0 B4.t0 19.0247
R8069 B4.n0 B4.t2 17.3935
R8070 B4.n1 B4.n0 4.12942
R8071 B4.n1 B4 2.25699
R8072 B4 B4.n1 0.0067069
R8073 B2 B2.t1 48.6474
R8074 B2.n0 B2.t0 19.0247
R8075 B2.n0 B2.t2 17.3935
R8076 B2.n1 B2.n0 4.12942
R8077 B2.n1 B2 2.25699
R8078 B2 B2.n1 0.0067069
R8079 SD2_2 SD2_2.n1 3.20344
R8080 SD2_2.n1 SD2_2.t1 2.7305
R8081 SD2_2.n1 SD2_2.n0 2.7305
C0 VDD b2 0.819f
C1 OUT2 SD2_1 0.00162f
C2 b1b B1 0.26f
C3 G1_1 SD1_1 0.279f
C4 b2 SD2_3 1.08e-19
C5 OUT3 SD2_5 0.182f
C6 b3 b5 0.0494f
C7 b3b b5b 0.0105f
C8 G1_2 OUT4 2.09f
C9 b2b SD2_4 0.00446f
C10 SDn_2 b3b 0.0274f
C11 b4 Balance_Inverter_4.Inverter_0.OUT 0.00897f
C12 b4 Balance_Inverter_1.Inverter_0.OUT 0.00255f
C13 b2 B2 0.101f
C14 VDD SD2_1 0.127f
C15 G2 SD2_2 0.0436f
C16 SD2_1 SD2_3 8.03e-19
C17 SD2_5 SD2_4 0.31f
C18 VDD C32_U 3.44f
C19 b6 SDc_1 6.59e-19
C20 b6b Gc_1 8.32e-19
C21 b5b b5 1.92f
C22 TG_0.IN b1b 0.256f
C23 IT SD3_1 1.01f
C24 SDc_2 C32_D 0.0287f
C25 TG_0.IN G1_1 8.45e-19
C26 TG_1.IN b3b 0.25f
C27 OUT+ IT 0.0189f
C28 SEL_L b1 6.5e-19
C29 IT b4b 9.29e-19
C30 TG_0.IN b6 2.79f
C31 TG_1.IN OUT4 0.841f
C32 IT Balance_Inverter_5.Inverter_0.OUT 0.0034f
C33 IT Balance_Inverter_0.Inverter_0.OUT 0.0034f
C34 b1b OUT5 0.204f
C35 b1 SDn_1 0.129f
C36 OUT6 b2b 0.323f
C37 SD3_1 b2 0.167f
C38 TG_1.IN b5 2.15f
C39 OUT+ b2 0.00128f
C40 b3b OUT4 0.0472f
C41 b1b ITAIL 0.0195f
C42 OUT1 G1_2 0.0347f
C43 OUT5 G1_1 0.0268f
C44 b1 G2 0.0264f
C45 b2b OUT2 0.0772f
C46 b2 b4b 0.0522f
C47 b1b Balance_Inverter_3.Inverter_0.OUT 0.0252f
C48 VDD b2b 0.687f
C49 b3 SDc_1 0.0347f
C50 b3 B3 0.0954f
C51 b2 Balance_Inverter_2.Inverter_0.OUT 0.224f
C52 b3 B5 0.0927f
C53 G1_2 SD1_1 0.646f
C54 G1_1 ITAIL 0.00302f
C55 b2b SD2_3 0.00175f
C56 b3b b5 4.52e-19
C57 OUT3 SD2_4 0.373f
C58 OUT2 SD2_5 0.363f
C59 SDn_2 OUT1 4.33e-19
C60 b2b B2 0.376f
C61 VDD SD2_5 1.38e-19
C62 SD2_5 SD2_3 0.0442f
C63 SDn_2 SD1_1 0.0268f
C64 VDD SDc_2 3.06f
C65 b6 Gc_1 1.52e-19
C66 b5b B5 0.169f
C67 b5b B3 0.0015f
C68 TG_0.IN b3 0.534f
C69 b5b B1 0.0019f
C70 SDn_2 B5 0.0593f
C71 SDn_2 SDc_1 0.654f
C72 SDn_2 B1 0.0616f
C73 SDn_2 B3 0.0613f
C74 IT b1 0.2f
C75 TG_0.IN G1_2 3.98e-19
C76 SEL_L b1b 9.16e-19
C77 TG_1.IN OUT1 0.257f
C78 IT b4 6.09e-19
C79 TG_0.IN b5b 1.39f
C80 TG_0.IN SDn_2 9.86e-21
C81 IT b6b 0.00534f
C82 SD3_1 b2b 0.576f
C83 OUT6 OUT3 0.00428f
C84 b3 OUT5 3.51e-19
C85 b1 b2 0.0351f
C86 b1b SDn_1 0.132f
C87 TG_1.IN SDc_1 7.58e-19
C88 TG_1.IN B5 2.65e-20
C89 TG_1.IN B3 1.23e-19
C90 TG_1.IN B1 7.92e-19
C91 OUT+ b2b 3.55e-19
C92 b2b b4b 0.033f
C93 b1 SD2_1 0.0946f
C94 b2 b4 0.0116f
C95 b3b SD1_1 0.0957f
C96 OUT5 G1_2 0.0345f
C97 SDn_1 G1_1 0.00119f
C98 b1b G2 0.0134f
C99 OUT1 OUT4 1.78f
C100 OUT3 OUT2 0.265f
C101 b3 Balance_Inverter_4.Inverter_0.OUT 0.0057f
C102 b3 Balance_Inverter_1.Inverter_0.OUT 0.228f
C103 VDD OUT3 4.91e-20
C104 b3b B5 0.00227f
C105 b3 Gc_1 0.033f
C106 b2b Balance_Inverter_2.Inverter_0.OUT 0.0239f
C107 b3b B1 0.0288f
C108 OUT4 SD1_1 0.0013f
C109 G1_2 ITAIL 0.568f
C110 OUT5 b5b 1.6f
C111 OUT2 SD2_4 0.281f
C112 b3b B3 0.596f
C113 OUT3 SD2_3 0.401f
C114 SDn_2 OUT5 0.926f
C115 TG_1.IN TG_0.IN 16.2f
C116 VDD OUT- 0.519f
C117 SD2_4 SD2_3 0.461f
C118 SD2_5 SD2_2 0.0175f
C119 ITAIL b5b 9.45e-19
C120 SDn_2 ITAIL 0.178f
C121 b5b Balance_Inverter_4.Inverter_0.OUT 0.00753f
C122 VDD C32_D 0.0116f
C123 b5 B5 0.0874f
C124 TG_0.IN b3b 0.391f
C125 b5 B3 1.07e-19
C126 SDn_2 Gc_1 1.33f
C127 IT b1b 0.316f
C128 TG_0.IN OUT4 0.815f
C129 TG_1.IN OUT5 2.33f
C130 SEL_L b3 4.54e-20
C131 IT G1_1 0.375f
C132 TG_0.IN b5 1.33f
C133 TG_1.IN ITAIL 1.71e-20
C134 TG_1.IN Balance_Inverter_4.Inverter_0.OUT 0.00136f
C135 TG_1.IN Balance_Inverter_3.Inverter_0.OUT 4.26e-21
C136 IT b6 0.00122f
C137 b3b OUT5 0.0251f
C138 b1 b2b 0.0403f
C139 b1b b2 0.0845f
C140 TG_1.IN Gc_1 2.41e-21
C141 VDD OUT6 0.0408f
C142 b1b SD2_1 0.0398f
C143 OUT1 SD1_1 5.9e-19
C144 b1 SD2_5 0.0356f
C145 OUT3 b4b 0.0594f
C146 b2 G1_1 0.0077f
C147 SDn_1 G1_2 5.13e-19
C148 b2b b4 9.46e-20
C149 b3b ITAIL 0.02f
C150 OUT5 OUT4 0.0458f
C151 OUT- OUT+ 0.0182f
C152 b3b Balance_Inverter_1.Inverter_0.OUT 0.0887f
C153 OUT6 B6 2.15e-19
C154 VDD OUT2 0.0816f
C155 OUT5 b5 1.49f
C156 OUT4 ITAIL 0.346f
C157 OUT2 SD2_3 0.16f
C158 G1_2 G2 0.192f
C159 SDn_2 SDn_1 0.586f
C160 G2 b5b 0.00908f
C161 VDD B6 0.359f
C162 VDD B4 0.566f
C163 VDD B2 0.455f
C164 SDn_2 G2 4.62e-20
C165 b5 Balance_Inverter_4.Inverter_0.OUT 0.219f
C166 SEL_L TG_1.IN 1.3f
C167 VDD m1_n558_n5402# 0.0568f
C168 B4 B6 0.00236f
C169 B3 B5 0.00166f
C170 TG_0.IN OUT1 0.172f
C171 IT b3 0.0686f
C172 TG_0.IN SD1_1 5.17e-20
C173 SEL_L b3b 0.13f
C174 IT G1_2 2.95f
C175 OUT6 SD3_1 3.97f
C176 TG_0.IN B1 0.00379f
C177 TG_1.IN G2 2.86e-20
C178 OUT+ OUT6 0.0226f
C179 IT b5b 9.39e-19
C180 b1 OUT3 0.0392f
C181 OUT6 b4b 0.19f
C182 b3 b2 0.0682f
C183 OUT1 OUT5 0.551f
C184 b3b SDn_1 0.11f
C185 b1b b2b 1.03f
C186 IT SDn_2 8.51f
C187 VDD SD3_1 0.147f
C188 b1b SD2_5 0.0386f
C189 b2 G1_2 0.045f
C190 OUT1 ITAIL 0.168f
C191 OUT3 b4 0.1f
C192 b3b G2 0.0141f
C193 b1 SD2_4 0.0372f
C194 b2b G1_1 0.0281f
C195 OUT5 SD1_1 0.0778f
C196 OUT2 b4b 0.107f
C197 VDD OUT+ 0.496f
C198 VDD b4b 0.428f
C199 OUT4 G2 0.246f
C200 SD1_1 ITAIL 0.00106f
C201 OUT5 B1 3.74e-21
C202 G1_2 SD2_1 0.906f
C203 OUT3 b6b 3.6e-21
C204 OUT2 SD2_2 0.00234f
C205 SDn_2 b2 0.0229f
C206 b4b B6 5.71e-19
C207 b4b B4 0.2f
C208 VDD Balance_Inverter_5.Inverter_0.OUT 0.14f
C209 VDD Balance_Inverter_0.Inverter_0.OUT 0.14f
C210 VDD Balance_Inverter_2.Inverter_0.OUT 0.154f
C211 b4b m1_n558_n5402# 0.0175f
C212 TG_1.IN IT 9.14e-20
C213 SD2_1 b5b 0.00393f
C214 B6 Balance_Inverter_5.Inverter_0.OUT 0.158f
C215 Balance_Inverter_0.Inverter_0.OUT B6 5.16e-19
C216 B5 Balance_Inverter_4.Inverter_0.OUT 0.159f
C217 B4 Balance_Inverter_0.Inverter_0.OUT 0.158f
C218 B3 Balance_Inverter_1.Inverter_0.OUT 0.139f
C219 B2 Balance_Inverter_2.Inverter_0.OUT 0.158f
C220 B1 Balance_Inverter_3.Inverter_0.OUT 0.158f
C221 B5 Gc_1 3.67e-20
C222 SDc_1 Gc_1 3.86f
C223 TG_0.IN OUT5 1.49f
C224 IT b3b 0.272f
C225 TG_1.IN b2 0.562f
C226 TG_0.IN Balance_Inverter_4.Inverter_0.OUT 3.2e-20
C227 IT OUT4 0.00118f
C228 OUT6 b1 0.0167f
C229 TG_1.IN SD2_1 7.37e-19
C230 OUT+ SD3_1 0.0884f
C231 IT b5 5.73e-19
C232 OUT1 SDn_1 0.00609f
C233 b3b b2 3.71f
C234 OUT6 b4 0.282f
C235 b3 b2b 0.127f
C236 b1 OUT2 1.07f
C237 b1b OUT3 0.0345f
C238 VDD b1 0.944f
C239 b3b SD2_1 0.0885f
C240 OUT5 ITAIL 0.0132f
C241 b2 OUT4 0.0745f
C242 OUT2 b4 0.00657f
C243 OUT1 G2 0.0299f
C244 b1 SD2_3 0.0369f
C245 b2b G1_2 0.0676f
C246 b1b SD2_4 0.0374f
C247 OUT3 G1_1 5.54e-20
C248 SDn_1 SD1_1 0.0889f
C249 OUT6 b6b 1.29f
C250 VDD b4 1.22f
C251 b4b Balance_Inverter_5.Inverter_0.OUT 1.27e-19
C252 b4b Balance_Inverter_0.Inverter_0.OUT 0.00424f
C253 b2b b5b 4.11e-19
C254 G1_2 SD2_5 0.00259f
C255 OUT4 SD2_1 0.0612f
C256 b2 b5 0.00157f
C257 SDn_2 b2b 0.105f
C258 b4 B6 0.0528f
C259 b4 B4 0.0688f
C260 SEL_L TG_0.IN 1.15f
C261 VDD b6b 0.316f
C262 b4 m1_n558_n5402# 1.3e-19
C263 G2 B1 4.42e-19
C264 SD2_1 b5 0.0012f
C265 b6b B6 0.209f
C266 SDc_1 Gc_2 0.0472f
C267 IT OUT1 0.00193f
C268 TG_0.IN G2 0.00111f
C269 TG_1.IN b2b 0.406f
C270 IT SD1_1 2.13f
C271 OUT6 b1b 0.199f
C272 SD3_1 b1 0.00977f
C273 OUT+ b1 7.91e-20
C274 IT SDc_1 0.909f
C275 IT B5 0.0859f
C276 IT B3 0.0741f
C277 IT B1 0.0736f
C278 b1 b4b 5.58e-20
C279 OUT1 b2 0.0236f
C280 OUT5 SDn_1 2.14f
C281 b1b OUT2 0.0214f
C282 b3 OUT3 0.139f
C283 b3b b2b 0.132f
C284 VDD b1b 0.594f
C285 b1 SD2_2 0.00207f
C286 OUT5 G2 0.0135f
C287 b1b SD2_3 0.0345f
C288 OUT2 G1_1 0.0171f
C289 b2 SD1_1 0.0595f
C290 OUT3 G1_2 0.0268f
C291 b2b OUT4 0.056f
C292 b4b b4 4.11f
C293 OUT6 b6 1.42f
C294 OUT1 SD2_1 0.023f
C295 b3b SD2_5 0.00858f
C296 VDD G1_1 8.11f
C297 b4 Balance_Inverter_5.Inverter_0.OUT 0.00832f
C298 b4 Balance_Inverter_0.Inverter_0.OUT 0.219f
C299 TG_0.IN IT 6.56e-19
C300 b2 B3 7.24e-19
C301 G1_2 SD2_4 2.28e-19
C302 b2 B1 0.193f
C303 b2b b5 0.00104f
C304 OUT3 b5b 0.00986f
C305 OUT4 SD2_5 1.05f
C306 ITAIL G2 1.17f
C307 b4b b6b 0.235f
C308 G2 Balance_Inverter_3.Inverter_0.OUT 4.19e-20
C309 VDD b6 0.567f
C310 b6b Balance_Inverter_5.Inverter_0.OUT 0.00445f
C311 SD2_1 B1 0.00539f
C312 b6 B6 0.0742f
C313 Gc_1 Gc_2 10.9f
C314 TG_0.IN b2 0.792f
C315 IT OUT5 1.02f
C316 TG_0.IN SD2_1 0.00903f
C317 TG_1.IN OUT3 0.7f
C318 IT ITAIL 0.321f
C319 OUT6 b3 0.835f
C320 SD3_1 b1b 0.272f
C321 TG_1.IN OUT- 18.1f
C322 IT Balance_Inverter_4.Inverter_0.OUT 0.0034f
C323 OUT+ b1b 7.18e-20
C324 IT Gc_1 0.799f
C325 OUT5 b2 0.0264f
C326 b3 OUT2 4.2e-20
C327 b1 b4 1.1e-19
C328 OUT1 b2b 0.00657f
C329 b3b OUT3 0.111f
C330 b1b b4b 0.00121f
C331 VDD b3 0.766f
C332 OUT2 G1_2 0.273f
C333 b3b SD2_4 9.52e-20
C334 OUT5 SD2_1 0.0727f
C335 OUT3 OUT4 1.33f
C336 OUT1 SD2_5 0.548f
C337 b2 ITAIL 0.00993f
C338 b4b G1_1 5.38e-19
C339 b2b SD1_1 0.0397f
C340 SDn_2 OUT6 1.22f
C341 b3 B6 0.412f
C342 b3 B2 0.164f
C343 b2 Balance_Inverter_3.Inverter_0.OUT 0.00628f
C344 b3 B4 0.0628f
C345 VDD G1_2 3.63f
C346 b3 m1_n558_n5402# 0.00587f
C347 OUT4 SD2_4 0.00348f
C348 ITAIL SD2_1 0.192f
C349 OUT3 b5 0.00482f
C350 b4 b6b 0.286f
C351 b2b B1 0.102f
C352 b4b b6 0.213f
C353 G1_2 SD2_3 8.28e-20
C354 b2b B3 0.00608f
C355 SDn_2 OUT2 0.0016f
C356 SD2_1 Balance_Inverter_3.Inverter_0.OUT 5.32e-19
C357 VDD b5b 0.38f
C358 b6 Balance_Inverter_5.Inverter_0.OUT 0.22f
C359 SEL_L IT 0.0536f
C360 VDD SDn_2 0.382f
C361 b5b B6 0.0476f
C362 b5b B2 6.52e-21
C363 SDn_2 B4 0.0665f
C364 SDn_2 B6 0.0868f
C365 Gc_1 C32_U 2.33f
C366 SDn_2 B2 0.0657f
C367 b5b m1_n558_n5402# 2.68e-20
C368 TG_0.IN b2b 0.48f
C369 TG_1.IN OUT6 6.7f
C370 IT SDn_1 1.02f
C371 TG_1.IN OUT2 0.471f
C372 SEL_L b2 0.00243f
C373 IT G2 0.00271f
C374 b1 b1b 2.47f
C375 OUT6 b3b 0.215f
C376 VDD TG_1.IN 6.13f
C377 IT Gc_2 0.136f
C378 TG_1.IN B6 0.00132f
C379 TG_1.IN B2 1.01e-20
C380 OUT5 b2b 0.164f
C381 OUT1 OUT3 0.223f
C382 b1 G1_1 0.0912f
C383 b3 b4b 0.202f
C384 SDn_1 b2 0.0994f
C385 VDD b3b 1.31f
C386 b3 Balance_Inverter_5.Inverter_0.OUT 0.00505f
C387 b3 Balance_Inverter_0.Inverter_0.OUT 0.0157f
C388 b3 Balance_Inverter_2.Inverter_0.OUT 0.00384f
C389 OUT1 SD2_4 0.00368f
C390 OUT2 OUT4 1.26f
C391 b3b SD2_3 6.42e-20
C392 b2 G2 0.0209f
C393 OUT3 SD1_1 1.31e-19
C394 b2b ITAIL 0.0175f
C395 SDn_2 SD3_1 0.716f
C396 b2b Balance_Inverter_1.Inverter_0.OUT 0.00182f
C397 b3b B6 0.00179f
C398 b2b Balance_Inverter_3.Inverter_0.OUT 0.00219f
C399 b3b B4 0.0167f
C400 b3b B2 0.0616f
C401 VDD OUT4 0.00148f
C402 OUT+ SDn_2 0.00114f
C403 b3b m1_n558_n5402# 0.00129f
C404 b4 b6 0.783f
C405 ITAIL SD2_5 0.265f
C406 b4b b5b 0.11f
C407 G2 SD2_1 0.214f
C408 OUT3 B1 3.71e-20
C409 OUT4 SD2_3 0.00229f
C410 VDD b5 0.754f
C411 b5b Balance_Inverter_5.Inverter_0.OUT 0.0132f
C412 b6b b6 3.11f
C413 b5 B6 0.0144f
C414 b5 B2 4.82e-19
C415 Gc_1 SDc_2 1.14f
C416 Gc_2 C32_U 0.714f
C417 b5 m1_n558_n5402# 1.27e-20
C418 TG_0.IN OUT3 1.43f
C419 IT b2 0.161f
C420 TG_1.IN OUT+ 4.74e-20
C421 TG_1.IN b4b 1.34f
C422 SEL_L b2b 0.00167f
C423 IT SD2_1 0.0154f
C424 b1 b3 6.43e-19
C425 OUT6 OUT1 0.0634f
C426 SD3_1 b3b 0.159f
C427 TG_1.IN Balance_Inverter_5.Inverter_0.OUT 2.36e-19
C428 OUT+ b3b 0.245f
C429 SDn_1 b2b 0.111f
C430 OUT1 OUT2 0.352f
C431 b1 G1_2 0.25f
C432 b1b G1_1 0.0784f
C433 OUT5 OUT3 0.0882f
C434 b3b b4b 0.0222f
C435 b3 b4 0.304f
C436 VDD OUT1 0.0376f
C437 b3b Balance_Inverter_0.Inverter_0.OUT 0.00272f
C438 b3b Balance_Inverter_2.Inverter_0.OUT 0.00135f
C439 OUT3 ITAIL 0.128f
C440 b1 b5b 9.41e-19
C441 b2b G2 0.0203f
C442 b2 SD2_1 0.0523f
C443 b3 b6b 0.0399f
C444 OUT2 SD1_1 0.0494f
C445 b4b OUT4 0.224f
C446 OUT1 SD2_3 0.00462f
C447 SDn_2 b1 0.0286f
C448 VDD SD1_1 1.94f
C449 b4b b5 0.154f
C450 G2 SD2_5 0.248f
C451 b4 b5b 0.0441f
C452 ITAIL SD2_4 0.124f
C453 VDD B5 0.354f
C454 VDD SDc_1 0.236f
C455 VDD B1 1.2f
C456 VDD B3 0.624f
C457 b5 Balance_Inverter_5.Inverter_0.OUT 0.00537f
C458 TG_0.IN OUT6 5.41f
C459 b6b b5b 0.00479f
C460 SDn_2 b6b 0.00212f
C461 B5 B6 1.99f
C462 B6 SDc_1 0.207f
C463 B3 B6 3.58e-19
C464 B4 B5 0.704f
C465 B3 B4 0.123f
C466 B2 B3 0.214f
C467 B1 B2 0.233f
C468 Gc_2 SDc_2 1.43f
C469 Gc_1 C32_D 0.00118f
C470 TG_0.IN OUT2 0.798f
C471 TG_1.IN b1 0.294f
C472 IT b2b 0.267f
C473 VDD TG_0.IN 5.93f
C474 TG_1.IN b4 1.52f
C475 TG_0.IN B6 1.53e-19
C476 TG_0.IN B2 0.0069f
C477 b1b b3 3.65e-19
C478 OUT6 OUT5 0.0131f
C479 b1 b3b 1.42e-19
C480 SEL_L OUT- 1.33f
C481 TG_1.IN b6b 2.62f
C482 OUT5 OUT2 0.0703f
C483 b1b G1_2 0.0867f
C484 b3b b4 0.00815f
C485 b1 OUT4 0.103f
C486 OUT1 b4b 4.44e-19
C487 b2 b2b 4.83f
C488 VDD OUT5 0.165f
C489 b2 SD2_5 0.0557f
C490 b3 b6 0.638f
C491 OUT3 G2 0.131f
C492 b2b SD2_1 0.0528f
C493 OUT1 SD2_2 0.037f
C494 OUT2 ITAIL 0.148f
C495 b1b b5b 0.00116f
C496 b4 OUT4 0.286f
C497 b1 b5 7.09e-19
C498 G1_1 G1_2 2.47f
C499 SDn_2 b1b 0.0933f
C500 OUT5 B2 1.94e-19
C501 VDD ITAIL 0.105f
C502 b4b B5 0.101f
C503 OUT4 b6b 0.0011f
C504 ITAIL SD2_3 0.0655f
C505 b4 b5 0.473f
C506 SD2_1 SD2_5 0.0861f
C507 G2 SD2_4 0.162f
C508 b4b B3 0.0144f
C509 VDD Balance_Inverter_4.Inverter_0.OUT 0.14f
C510 VDD Balance_Inverter_1.Inverter_0.OUT 0.153f
C511 VDD Balance_Inverter_3.Inverter_0.OUT 0.154f
C512 SDn_2 G1_1 0.012f
C513 VDD Gc_1 18.6f
C514 Balance_Inverter_5.Inverter_0.OUT SDc_1 7.75e-20
C515 Balance_Inverter_4.Inverter_0.OUT B6 0.00172f
C516 B5 Balance_Inverter_5.Inverter_0.OUT 0.00101f
C517 Balance_Inverter_0.Inverter_0.OUT B5 0.00206f
C518 B4 Balance_Inverter_4.Inverter_0.OUT 9.91e-19
C519 Balance_Inverter_1.Inverter_0.OUT B4 5.37e-20
C520 B3 Balance_Inverter_0.Inverter_0.OUT 0.00299f
C521 B1 Balance_Inverter_2.Inverter_0.OUT 0.00299f
C522 Balance_Inverter_2.Inverter_0.OUT B3 5.45e-20
C523 B2 Balance_Inverter_1.Inverter_0.OUT 0.00207f
C524 Balance_Inverter_3.Inverter_0.OUT B2 5.37e-20
C525 TG_0.IN SD3_1 0.0139f
C526 b6 b5b 0.0019f
C527 b6b b5 0.0482f
C528 SDn_2 b6 5.16e-20
C529 B6 Gc_1 0.0129f
C530 B4 Gc_1 4.45e-21
C531 TG_0.IN OUT+ 18.2f
C532 Gc_2 C32_D 0.0107f
C533 C32_U SDc_2 3.46f
C534 TG_0.IN b4b 1.18f
C535 SEL_L OUT6 0.102f
C536 TG_1.IN b1b 0.131f
C537 IT OUT3 4.23e-20
C538 TG_0.IN Balance_Inverter_5.Inverter_0.OUT 3.93e-21
C539 TG_0.IN Balance_Inverter_2.Inverter_0.OUT 3.09e-21
C540 TG_1.IN G1_1 4.07e-20
C541 OUT6 SDn_1 0.0272f
C542 SD3_1 OUT5 0.0124f
C543 b1 OUT1 0.14f
C544 b1b b3b 1.73e-19
C545 VDD SEL_L 3.04f
C546 TG_1.IN b6 3.42f
C547 b1b OUT4 0.0382f
C548 b3b G1_1 0.00976f
C549 OUT5 b4b 0.00918f
C550 b1 SD1_1 0.136f
C551 SDn_1 OUT2 0.00105f
C552 OUT1 b4 5.52e-19
C553 b2 OUT3 0.0568f
C554 VDD SDn_1 0.0091f
C555 OUT5 Balance_Inverter_5.Inverter_0.OUT 7.09e-20
C556 G1_1 OUT4 2.54e-19
C557 b1 B1 0.0809f
C558 b2b SD2_5 0.0626f
C559 OUT3 SD2_1 1.08f
C560 b3 b5b 0.0546f
C561 b2 SD2_4 1.72e-19
C562 OUT2 G2 0.0518f
C563 b1b b5 5.92e-19
C564 SDn_2 b3 0.0353f
C565 b4b Balance_Inverter_4.Inverter_0.OUT 0.0129f
C566 b4b Balance_Inverter_1.Inverter_0.OUT 1.07e-19
C567 VDD G2 0.0272f
C568 b4 B3 0.138f
C569 b4 B5 0.0616f
C570 G1_2 b5b 2.13e-19
C571 G2 SD2_3 0.0979f
C572 SD2_1 SD2_4 0.00298f
C573 ITAIL SD2_2 0.00992f
C574 SDn_2 G1_2 9.11e-20
C575 Balance_Inverter_4.Inverter_0.OUT Balance_Inverter_5.Inverter_0.OUT 3.48e-19
C576 Balance_Inverter_0.Inverter_0.OUT Balance_Inverter_4.Inverter_0.OUT 3.46e-19
C577 Balance_Inverter_2.Inverter_0.OUT Balance_Inverter_1.Inverter_0.OUT 0.00442f
C578 Balance_Inverter_1.Inverter_0.OUT Balance_Inverter_0.Inverter_0.OUT 0.00437f
C579 Balance_Inverter_3.Inverter_0.OUT Balance_Inverter_2.Inverter_0.OUT 0.00437f
C580 VDD Gc_2 28.2f
C581 b6b SDc_1 0.00827f
C582 TG_0.IN b1 0.119f
C583 b6 b5 0.0112f
C584 IT OUT6 0.783f
C585 C32_U C32_D 5.52f
C586 TG_0.IN b4 1.31f
C587 TG_1.IN b3 0.794f
C588 SEL_L SD3_1 0.0232f
C589 IT OUT2 0.093f
C590 SEL_L OUT+ 1.34f
C591 TG_0.IN b6b 2.58f
C592 TG_1.IN G1_2 8.68e-23
C593 VDD IT 2.54f
C594 SD3_1 SDn_1 0.297f
C595 b1b OUT1 0.0235f
C596 b3 b3b 0.982f
C597 b1 OUT5 0.0759f
C598 OUT6 b2 0.323f
C599 IT B6 0.485f
C600 IT B4 0.096f
C601 IT B2 0.079f
C602 TG_1.IN b5b 1.25f
C603 TG_1.IN SDn_2 0.00121f
C604 OUT1 G1_1 5.82e-19
C605 b3b G1_2 0.0816f
C606 b2b OUT3 0.00957f
C607 b1b SD1_1 0.223f
C608 b2 OUT2 0.0421f
C609 OUT5 b4 4.5e-19
C610 b1 ITAIL 0.0202f
C611 b1 Balance_Inverter_3.Inverter_0.OUT 0.221f
C612 m1_n558_n5402# VSS 0.0572f $ **FLOATING
C613 C32_D VSS 13f
C614 SDc_2 VSS 0.515f
C615 C32_U VSS 20.1f
C616 Gc_2 VSS 4.39f
C617 Gc_1 VSS 9.04f
C618 SDc_1 VSS 3.4f
C619 Balance_Inverter_5.Inverter_0.OUT VSS 0.553f
C620 B6 VSS 2.85f
C621 Balance_Inverter_4.Inverter_0.OUT VSS 0.553f
C622 B5 VSS 2.26f
C623 Balance_Inverter_0.Inverter_0.OUT VSS 0.562f
C624 B4 VSS 2.65f
C625 Balance_Inverter_1.Inverter_0.OUT VSS 0.55f
C626 B3 VSS 2.52f
C627 Balance_Inverter_2.Inverter_0.OUT VSS 0.549f
C628 B2 VSS 2.61f
C629 Balance_Inverter_3.Inverter_0.OUT VSS 0.552f
C630 B1 VSS 2.26f
C631 b5 VSS 6.56f
C632 b5b VSS 7.46f
C633 b6 VSS 13.7f
C634 b6b VSS 14.4f
C635 SD2_2 VSS 0.0529f
C636 SD2_3 VSS 1.08f
C637 SD2_4 VSS 0.57f
C638 SD2_5 VSS 1.01f
C639 SD2_1 VSS 2.59f
C640 G2 VSS 7.65f
C641 ITAIL VSS 9.62f
C642 SD1_1 VSS 0.746f
C643 OUT4 VSS 3.18f
C644 G1_2 VSS 5.28f
C645 G1_1 VSS 1.57f
C646 b4 VSS 6.35f
C647 b4b VSS 8.37f
C648 OUT2 VSS 1.58f
C649 OUT3 VSS 1.84f
C650 b2b VSS 5.85f
C651 b2 VSS 3.52f
C652 SDn_1 VSS 2.33f
C653 OUT5 VSS 4.71f
C654 OUT1 VSS 1.3f
C655 b3b VSS 5.3f
C656 b3 VSS 7.89f
C657 b1b VSS 4.01f
C658 b1 VSS 4.51f
C659 SD3_1 VSS 3.75f
C660 OUT6 VSS 11.1f
C661 SDn_2 VSS 29.3f
C662 IT VSS 44.9f
C663 OUT+ VSS 14.9f
C664 TG_0.IN VSS 21.8f
C665 OUT- VSS 13.2f
C666 TG_1.IN VSS 24.3f
C667 SEL_L VSS 17.9f
C668 VDD VSS 0.158p
C669 b1.n0 VSS 0.00429f
C670 b1.t2 VSS 0.0263f
C671 b1.n1 VSS 0.0245f
C672 b1.t4 VSS 0.0025f
C673 b1.n2 VSS 0.00755f
C674 b1.n3 VSS 0.38f
C675 b1.t3 VSS 0.0221f
C676 b1.n4 VSS 0.112f
C677 b1.t1 VSS 0.00677f
C678 b1.t0 VSS 0.00536f
C679 b1.n5 VSS 0.116f
C680 b3b.n0 VSS 0.00469f
C681 b3b.n1 VSS 0.0325f
C682 b3b.n2 VSS 0.00523f
C683 b3b.n3 VSS 0.0274f
C684 b3b.t2 VSS 0.00861f
C685 b3b.t4 VSS 0.0172f
C686 b3b.t9 VSS 0.0312f
C687 b3b.t8 VSS 0.0269f
C688 b3b.t5 VSS 0.0376f
C689 b3b.n4 VSS 0.0308f
C690 b3b.t10 VSS 0.0269f
C691 b3b.t7 VSS 0.0375f
C692 b3b.n5 VSS 0.031f
C693 b3b.t6 VSS 0.0311f
C694 b3b.t3 VSS 1.01f
C695 b3b.n6 VSS 2.26f
C696 C32_D.t55 VSS 0.00728f
C697 C32_D.n0 VSS 0.00728f
C698 C32_D.n1 VSS 0.0153f
C699 C32_D.t66 VSS 0.00728f
C700 C32_D.n2 VSS 0.00728f
C701 C32_D.n3 VSS 0.0153f
C702 C32_D.t35 VSS 0.00728f
C703 C32_D.n4 VSS 0.00728f
C704 C32_D.n5 VSS 0.0152f
C705 C32_D.t69 VSS 0.00728f
C706 C32_D.n6 VSS 0.00728f
C707 C32_D.n7 VSS 0.0153f
C708 C32_D.t45 VSS 0.00728f
C709 C32_D.n8 VSS 0.00728f
C710 C32_D.n9 VSS 0.0153f
C711 C32_D.t93 VSS 0.00728f
C712 C32_D.n10 VSS 0.00728f
C713 C32_D.n11 VSS 0.0153f
C714 C32_D.t23 VSS 0.00728f
C715 C32_D.n12 VSS 0.00728f
C716 C32_D.n13 VSS 0.0153f
C717 C32_D.t95 VSS 0.00728f
C718 C32_D.n14 VSS 0.00728f
C719 C32_D.n15 VSS 0.0153f
C720 C32_D.t25 VSS 0.00728f
C721 C32_D.n16 VSS 0.00728f
C722 C32_D.n17 VSS 0.0153f
C723 C32_D.t74 VSS 0.00728f
C724 C32_D.n18 VSS 0.00728f
C725 C32_D.n19 VSS 0.0153f
C726 C32_D.t47 VSS 0.00728f
C727 C32_D.n20 VSS 0.00728f
C728 C32_D.n21 VSS 0.0153f
C729 C32_D.t89 VSS 0.00728f
C730 C32_D.n22 VSS 0.00728f
C731 C32_D.n23 VSS 0.0153f
C732 C32_D.t21 VSS 0.00728f
C733 C32_D.n24 VSS 0.00728f
C734 C32_D.n25 VSS 0.0153f
C735 C32_D.t87 VSS 0.00728f
C736 C32_D.n26 VSS 0.00728f
C737 C32_D.n27 VSS 0.0153f
C738 C32_D.t12 VSS 0.0209f
C739 C32_D.n28 VSS 0.0323f
C740 C32_D.t13 VSS 0.00728f
C741 C32_D.n29 VSS 0.00728f
C742 C32_D.n30 VSS 0.016f
C743 C32_D.n31 VSS 0.0623f
C744 C32_D.t67 VSS 0.00728f
C745 C32_D.n32 VSS 0.00728f
C746 C32_D.n33 VSS 0.016f
C747 C32_D.n34 VSS 0.0331f
C748 C32_D.n35 VSS 0.0179f
C749 C32_D.t42 VSS 0.023f
C750 C32_D.n36 VSS 0.023f
C751 C32_D.n37 VSS 0.0239f
C752 C32_D.n38 VSS 0.0167f
C753 C32_D.t38 VSS 0.023f
C754 C32_D.n39 VSS 0.023f
C755 C32_D.n40 VSS 0.0239f
C756 C32_D.t39 VSS 0.00728f
C757 C32_D.n41 VSS 0.00728f
C758 C32_D.n42 VSS 0.0155f
C759 C32_D.n43 VSS 0.0317f
C760 C32_D.n44 VSS 0.0365f
C761 C32_D.t40 VSS 0.0209f
C762 C32_D.n45 VSS 0.0167f
C763 C32_D.n46 VSS 0.0209f
C764 C32_D.n47 VSS 0.0359f
C765 C32_D.t20 VSS 0.0209f
C766 C32_D.n48 VSS 0.0167f
C767 C32_D.n49 VSS 0.0209f
C768 C32_D.n50 VSS 0.0359f
C769 C32_D.n51 VSS 0.0365f
C770 C32_D.t70 VSS 0.00728f
C771 C32_D.n52 VSS 0.00728f
C772 C32_D.n53 VSS 0.0155f
C773 C32_D.n54 VSS 0.0317f
C774 C32_D.n55 VSS 0.0167f
C775 C32_D.t10 VSS 0.023f
C776 C32_D.n56 VSS 0.023f
C777 C32_D.n57 VSS 0.0239f
C778 C32_D.n58 VSS 0.0167f
C779 C32_D.t48 VSS 0.023f
C780 C32_D.n59 VSS 0.023f
C781 C32_D.n60 VSS 0.0239f
C782 C32_D.t49 VSS 0.00728f
C783 C32_D.n61 VSS 0.00728f
C784 C32_D.n62 VSS 0.0155f
C785 C32_D.n63 VSS 0.0317f
C786 C32_D.n64 VSS 0.0365f
C787 C32_D.t50 VSS 0.0209f
C788 C32_D.n65 VSS 0.0167f
C789 C32_D.n66 VSS 0.0209f
C790 C32_D.n67 VSS 0.0359f
C791 C32_D.t46 VSS 0.0209f
C792 C32_D.n68 VSS 0.0167f
C793 C32_D.n69 VSS 0.0209f
C794 C32_D.n70 VSS 0.0359f
C795 C32_D.n71 VSS 0.0365f
C796 C32_D.t84 VSS 0.00728f
C797 C32_D.n72 VSS 0.00728f
C798 C32_D.n73 VSS 0.0155f
C799 C32_D.n74 VSS 0.0317f
C800 C32_D.n75 VSS 0.0167f
C801 C32_D.t18 VSS 0.023f
C802 C32_D.n76 VSS 0.023f
C803 C32_D.n77 VSS 0.0239f
C804 C32_D.n78 VSS 0.0167f
C805 C32_D.t16 VSS 0.023f
C806 C32_D.n79 VSS 0.023f
C807 C32_D.n80 VSS 0.0239f
C808 C32_D.t17 VSS 0.00728f
C809 C32_D.n81 VSS 0.00728f
C810 C32_D.n82 VSS 0.0155f
C811 C32_D.n83 VSS 0.0317f
C812 C32_D.n84 VSS 0.0365f
C813 C32_D.t30 VSS 0.0209f
C814 C32_D.n85 VSS 0.0167f
C815 C32_D.n86 VSS 0.0209f
C816 C32_D.n87 VSS 0.0359f
C817 C32_D.t24 VSS 0.0209f
C818 C32_D.n88 VSS 0.0167f
C819 C32_D.n89 VSS 0.0209f
C820 C32_D.n90 VSS 0.0359f
C821 C32_D.n91 VSS 0.0365f
C822 C32_D.t76 VSS 0.00728f
C823 C32_D.n92 VSS 0.00728f
C824 C32_D.n93 VSS 0.0155f
C825 C32_D.n94 VSS 0.0317f
C826 C32_D.n95 VSS 0.0167f
C827 C32_D.t52 VSS 0.023f
C828 C32_D.n96 VSS 0.023f
C829 C32_D.n97 VSS 0.0239f
C830 C32_D.n98 VSS 0.0167f
C831 C32_D.t60 VSS 0.023f
C832 C32_D.n99 VSS 0.023f
C833 C32_D.n100 VSS 0.0239f
C834 C32_D.t61 VSS 0.00728f
C835 C32_D.n101 VSS 0.00728f
C836 C32_D.n102 VSS 0.0155f
C837 C32_D.n103 VSS 0.0317f
C838 C32_D.n104 VSS 0.0365f
C839 C32_D.t62 VSS 0.0209f
C840 C32_D.n105 VSS 0.0167f
C841 C32_D.n106 VSS 0.0209f
C842 C32_D.n107 VSS 0.0359f
C843 C32_D.t22 VSS 0.0209f
C844 C32_D.n108 VSS 0.0167f
C845 C32_D.n109 VSS 0.0209f
C846 C32_D.n110 VSS 0.0359f
C847 C32_D.n111 VSS 0.0365f
C848 C32_D.t71 VSS 0.00728f
C849 C32_D.n112 VSS 0.00728f
C850 C32_D.n113 VSS 0.0155f
C851 C32_D.n114 VSS 0.0317f
C852 C32_D.n115 VSS 0.0167f
C853 C32_D.t14 VSS 0.023f
C854 C32_D.n116 VSS 0.023f
C855 C32_D.n117 VSS 0.0239f
C856 C32_D.n118 VSS 0.0167f
C857 C32_D.t58 VSS 0.023f
C858 C32_D.n119 VSS 0.023f
C859 C32_D.n120 VSS 0.0239f
C860 C32_D.t59 VSS 0.00728f
C861 C32_D.n121 VSS 0.00728f
C862 C32_D.n122 VSS 0.0155f
C863 C32_D.n123 VSS 0.0317f
C864 C32_D.n124 VSS 0.0365f
C865 C32_D.t36 VSS 0.0209f
C866 C32_D.n125 VSS 0.0167f
C867 C32_D.n126 VSS 0.0209f
C868 C32_D.n127 VSS 0.0359f
C869 C32_D.t44 VSS 0.0209f
C870 C32_D.n128 VSS 0.0167f
C871 C32_D.n129 VSS 0.0209f
C872 C32_D.n130 VSS 0.0359f
C873 C32_D.n131 VSS 0.0365f
C874 C32_D.t83 VSS 0.00728f
C875 C32_D.n132 VSS 0.00728f
C876 C32_D.n133 VSS 0.0155f
C877 C32_D.n134 VSS 0.0317f
C878 C32_D.n135 VSS 0.0167f
C879 C32_D.t4 VSS 0.023f
C880 C32_D.n136 VSS 0.023f
C881 C32_D.n137 VSS 0.0239f
C882 C32_D.n138 VSS 0.0167f
C883 C32_D.t6 VSS 0.023f
C884 C32_D.n139 VSS 0.023f
C885 C32_D.n140 VSS 0.0239f
C886 C32_D.t7 VSS 0.00728f
C887 C32_D.n141 VSS 0.00728f
C888 C32_D.n142 VSS 0.0155f
C889 C32_D.n143 VSS 0.0317f
C890 C32_D.n144 VSS 0.0365f
C891 C32_D.t56 VSS 0.0209f
C892 C32_D.n145 VSS 0.0167f
C893 C32_D.n146 VSS 0.0209f
C894 C32_D.n147 VSS 0.0359f
C895 C32_D.t34 VSS 0.0205f
C896 C32_D.n148 VSS 0.017f
C897 C32_D.n149 VSS 0.0209f
C898 C32_D.n150 VSS 0.0366f
C899 C32_D.n151 VSS 0.037f
C900 C32_D.t79 VSS 0.00728f
C901 C32_D.n152 VSS 0.00728f
C902 C32_D.n153 VSS 0.0155f
C903 C32_D.n154 VSS 0.0314f
C904 C32_D.n155 VSS 0.0185f
C905 C32_D.t32 VSS 0.0211f
C906 C32_D.n156 VSS 0.023f
C907 C32_D.n157 VSS 0.0239f
C908 C32_D.n158 VSS 0.0175f
C909 C32_D.t0 VSS 0.0222f
C910 C32_D.n159 VSS 0.023f
C911 C32_D.n160 VSS 0.0239f
C912 C32_D.t1 VSS 0.00728f
C913 C32_D.n161 VSS 0.00728f
C914 C32_D.n162 VSS 0.0155f
C915 C32_D.n163 VSS 0.0315f
C916 C32_D.n164 VSS 0.0366f
C917 C32_D.t8 VSS 0.0209f
C918 C32_D.n165 VSS 0.0167f
C919 C32_D.n166 VSS 0.0209f
C920 C32_D.n167 VSS 0.0359f
C921 C32_D.t54 VSS 0.0209f
C922 C32_D.n168 VSS 0.0167f
C923 C32_D.n169 VSS 0.0209f
C924 C32_D.n170 VSS 0.0359f
C925 C32_D.n171 VSS 0.0365f
C926 C32_D.t91 VSS 0.00728f
C927 C32_D.n172 VSS 0.00728f
C928 C32_D.n173 VSS 0.0155f
C929 C32_D.n174 VSS 0.0282f
C930 C32_D.n175 VSS 0.0083f
C931 C32_D.n176 VSS 0.0166f
C932 C32_D.n177 VSS 2.58e-19
C933 C32_D.n178 VSS 0.00361f
C934 C32_D.n179 VSS 0.187f
C935 C32_D.t26 VSS 0.019f
C936 C32_D.n180 VSS 0.0191f
C937 C32_D.n181 VSS 0.00756f
C938 C32_D.n182 VSS 0.0124f
C939 C32_D.t2 VSS 0.0428f
C940 C32_D.n183 VSS 0.0279f
C941 C32_D.t28 VSS 0.023f
C942 C32_D.n184 VSS 0.023f
C943 C32_D.n185 VSS 0.0152f
C944 C32_D.t82 VSS 0.00728f
C945 C32_D.n186 VSS 0.00728f
C946 C32_D.n187 VSS 0.016f
C947 C32_D.t29 VSS 0.00728f
C948 C32_D.n188 VSS 0.00728f
C949 C32_D.n189 VSS 0.0154f
C950 C32_D.n190 VSS 0.0563f
C951 G1_1.t12 VSS 0.109f
C952 G1_1.n0 VSS 0.108f
C953 G1_1.t21 VSS 0.0392f
C954 G1_1.n1 VSS 0.0392f
C955 G1_1.n2 VSS 0.0826f
C956 G1_1.t15 VSS 0.0392f
C957 G1_1.n3 VSS 0.0392f
C958 G1_1.n4 VSS 0.0837f
C959 G1_1.t16 VSS 0.0392f
C960 G1_1.n5 VSS 0.0392f
C961 G1_1.n6 VSS 0.0837f
C962 G1_1.t9 VSS 0.0392f
C963 G1_1.n7 VSS 0.0392f
C964 G1_1.n8 VSS 0.0837f
C965 G1_1.t22 VSS 0.0392f
C966 G1_1.n9 VSS 0.0392f
C967 G1_1.n10 VSS 0.0837f
C968 G1_1.t3 VSS 0.0392f
C969 G1_1.n11 VSS 0.0392f
C970 G1_1.n12 VSS 0.0837f
C971 G1_1.t18 VSS 0.0392f
C972 G1_1.n13 VSS 0.0392f
C973 G1_1.n14 VSS 0.0837f
C974 G1_1.t7 VSS 0.0392f
C975 G1_1.n15 VSS 0.0392f
C976 G1_1.n16 VSS 0.0826f
C977 G1_1.t28 VSS 0.352f
C978 G1_1.t29 VSS 0.128f
C979 G1_1.n17 VSS 0.303f
C980 G1_1.t34 VSS 0.128f
C981 G1_1.n18 VSS 0.275f
C982 G1_1.t32 VSS 0.128f
C983 G1_1.n19 VSS 0.33f
C984 G1_1.n20 VSS 0.242f
C985 G1_1.t14 VSS 0.128f
C986 G1_1.n21 VSS 0.275f
C987 G1_1.t4 VSS 0.128f
C988 G1_1.n22 VSS 0.275f
C989 G1_1.t8 VSS 0.128f
C990 G1_1.n23 VSS 0.275f
C991 G1_1.t0 VSS 0.128f
C992 G1_1.n24 VSS 0.275f
C993 G1_1.t2 VSS 0.128f
C994 G1_1.n25 VSS 0.275f
C995 G1_1.t10 VSS 0.128f
C996 G1_1.n26 VSS 0.275f
C997 G1_1.t24 VSS 0.353f
C998 G1_1.t30 VSS 0.128f
C999 G1_1.n27 VSS 0.303f
C1000 G1_1.t35 VSS 0.128f
C1001 G1_1.n28 VSS 0.275f
C1002 G1_1.t25 VSS 0.128f
C1003 G1_1.n29 VSS 0.325f
C1004 G1_1.n30 VSS 0.236f
C1005 G1_1.t6 VSS 0.109f
C1006 G1_1.n31 VSS 0.111f
C1007 G1_1.n32 VSS 0.353f
C1008 G1_1.n33 VSS 0.328f
C1009 G1_1.n34 VSS 0.33f
C1010 G1_1.n35 VSS 0.33f
C1011 G1_1.n36 VSS 0.33f
C1012 G1_1.n37 VSS 0.33f
C1013 G1_1.n38 VSS 0.304f
C1014 G1_1.n39 VSS 0.148f
C1015 SD1_1.t3 VSS 0.0112f
C1016 SD1_1.n0 VSS 0.0112f
C1017 SD1_1.n1 VSS 0.0224f
C1018 SD1_1.n2 VSS 0.00497f
C1019 SD1_1.n3 VSS 0.022f
C1020 SD1_1.t5 VSS 0.0112f
C1021 SD1_1.n4 VSS 0.0112f
C1022 SD1_1.n5 VSS 0.0297f
C1023 SD1_1.t6 VSS 0.0112f
C1024 SD1_1.n6 VSS 0.0112f
C1025 SD1_1.n7 VSS 0.0308f
C1026 SD1_1.n8 VSS 0.0121f
C1027 SD1_1.t2 VSS 0.0103f
C1028 SD1_1.n9 VSS 0.0453f
C1029 SD1_1.n10 VSS 0.143f
C1030 SD1_1.n11 VSS 0.094f
C1031 SD1_1.t7 VSS 0.0112f
C1032 SD1_1.n12 VSS 0.0112f
C1033 SD1_1.n13 VSS 0.0337f
C1034 SD1_1.n14 VSS 0.559f
C1035 SD1_1.n15 VSS 0.506f
C1036 SD1_1.t8 VSS 0.0104f
C1037 SD1_1.n16 VSS 0.012f
C1038 SD1_1.n17 VSS 0.0519f
C1039 SD1_1.t14 VSS 0.0112f
C1040 SD1_1.n18 VSS 0.0112f
C1041 SD1_1.n19 VSS 0.0347f
C1042 SD1_1.n20 VSS 0.153f
C1043 SD1_1.t13 VSS 0.0112f
C1044 SD1_1.n21 VSS 0.0112f
C1045 SD1_1.n22 VSS 0.0347f
C1046 SD1_1.n23 VSS 0.0988f
C1047 SD1_1.n24 VSS 0.0438f
C1048 G1_2.t31 VSS 0.143f
C1049 G1_2.t26 VSS 0.0827f
C1050 G1_2.n0 VSS 0.212f
C1051 G1_2.t24 VSS 0.0827f
C1052 G1_2.n1 VSS 0.174f
C1053 G1_2.t28 VSS 0.0827f
C1054 G1_2.n2 VSS 0.208f
C1055 G1_2.t12 VSS 0.0827f
C1056 G1_2.t8 VSS 0.0827f
C1057 G1_2.t10 VSS 0.0827f
C1058 G1_2.n3 VSS 0.174f
C1059 G1_2.n4 VSS 0.174f
C1060 G1_2.n5 VSS 0.174f
C1061 G1_2.n6 VSS 0.149f
C1062 G1_2.n7 VSS 0.00736f
C1063 G1_2.n8 VSS 0.012f
C1064 G1_2.t16 VSS 0.0572f
C1065 G1_2.n9 VSS 0.0564f
C1066 G1_2.n10 VSS 0.0239f
C1067 G1_2.t22 VSS 0.0827f
C1068 G1_2.n11 VSS 0.174f
C1069 G1_2.t14 VSS 0.0827f
C1070 G1_2.n12 VSS 0.174f
C1071 G1_2.t18 VSS 0.0827f
C1072 G1_2.n13 VSS 0.174f
C1073 G1_2.t29 VSS 0.143f
C1074 G1_2.t34 VSS 0.0827f
C1075 G1_2.n14 VSS 0.212f
C1076 G1_2.t30 VSS 0.0827f
C1077 G1_2.n15 VSS 0.174f
C1078 G1_2.t32 VSS 0.0827f
C1079 G1_2.n16 VSS 0.204f
C1080 G1_2.n17 VSS 0.146f
C1081 G1_2.n18 VSS 0.00327f
C1082 G1_2.t17 VSS 0.0244f
C1083 G1_2.n19 VSS 0.0244f
C1084 G1_2.n20 VSS 0.0517f
C1085 G1_2.t15 VSS 0.0244f
C1086 G1_2.n21 VSS 0.0244f
C1087 G1_2.n22 VSS 0.0525f
C1088 G1_2.t11 VSS 0.0244f
C1089 G1_2.n23 VSS 0.0244f
C1090 G1_2.n24 VSS 0.0525f
C1091 G1_2.t13 VSS 0.0244f
C1092 G1_2.n25 VSS 0.0244f
C1093 G1_2.n26 VSS 0.0517f
C1094 G1_2.n27 VSS 0.0312f
C1095 G1_2.n28 VSS 0.209f
C1096 G1_2.n29 VSS 0.354f
C1097 G1_2.n30 VSS 0.354f
C1098 G1_2.n31 VSS 0.225f
C1099 G1_2.n32 VSS 0.0327f
C1100 G1_2.n33 VSS 0.0123f
C1101 G1_2.n34 VSS 0.0413f
C1102 G1_2.n35 VSS 0.0557f
C1103 G1_2.n36 VSS 0.0557f
C1104 G1_2.t7 VSS 0.0661f
C1105 G1_2.t0 VSS 0.0557f
C1106 G1_2.n37 VSS 0.376f
C1107 G1_2.n38 VSS 0.279f
C1108 G1_2.n39 VSS 0.434f
C1109 G1_2.n40 VSS 1.28f
C1110 G1_2.t1 VSS 0.0557f
C1111 G1_2.t2 VSS 0.0557f
C1112 G1_2.n41 VSS 0.0661f
C1113 G1_2.n42 VSS 0.0557f
C1114 G1_2.n43 VSS 0.381f
C1115 G1_2.n44 VSS 0.285f
C1116 G1_2.n45 VSS 0.463f
C1117 G1_2.n46 VSS 1.32f
C1118 G1_2.t20 VSS 0.0564f
C1119 G1_2.n47 VSS 0.0548f
C1120 G1_2.n48 VSS 0.0228f
C1121 G1_2.n49 VSS 0.0395f
C1122 b4.n0 VSS 0.00816f
C1123 b4.t11 VSS 0.00241f
C1124 b4.t3 VSS 0.0268f
C1125 b4.t10 VSS 0.098f
C1126 b4.n1 VSS 0.0545f
C1127 b4.n2 VSS 0.0155f
C1128 b4.n3 VSS 0.0276f
C1129 b4.t4 VSS 0.0233f
C1130 b4.n4 VSS 0.11f
C1131 b4.t14 VSS 0.0271f
C1132 b4.t6 VSS 0.031f
C1133 b4.t18 VSS 0.0453f
C1134 b4.t2 VSS 0.0435f
C1135 b4.t8 VSS 0.114f
C1136 b4.t9 VSS 0.0607f
C1137 b4.t17 VSS 0.0754f
C1138 b4.n5 VSS 0.0752f
C1139 b4.t15 VSS 0.0612f
C1140 b4.t13 VSS 0.125f
C1141 b4.t16 VSS 0.107f
C1142 b4.t5 VSS 0.0655f
C1143 b4.n6 VSS 0.102f
C1144 b4.n7 VSS 0.124f
C1145 b4.t7 VSS 0.0762f
C1146 b4.n8 VSS 0.0623f
C1147 b4.n9 VSS 1.11f
C1148 b4.t12 VSS 0.0309f
C1149 b4.n10 VSS 0.0606f
C1150 b4.t1 VSS 0.00966f
C1151 b4.t0 VSS 0.00765f
C1152 b4.n11 VSS 0.165f
C1153 SDn_1.t18 VSS 0.00812f
C1154 SDn_1.n0 VSS 0.00812f
C1155 SDn_1.n1 VSS 0.0163f
C1156 SDn_1.n2 VSS 0.0188f
C1157 SDn_1.t1 VSS 0.00812f
C1158 SDn_1.n3 VSS 0.00812f
C1159 SDn_1.n4 VSS 0.0223f
C1160 SDn_1.t9 VSS 0.00812f
C1161 SDn_1.n5 VSS 0.00812f
C1162 SDn_1.n6 VSS 0.0284f
C1163 SDn_1.t26 VSS 0.00812f
C1164 SDn_1.n7 VSS 0.00812f
C1165 SDn_1.n8 VSS 0.0296f
C1166 SDn_1.t11 VSS 0.00812f
C1167 SDn_1.n9 VSS 0.00812f
C1168 SDn_1.n10 VSS 0.0297f
C1169 SDn_1.t27 VSS 0.00812f
C1170 SDn_1.n11 VSS 0.00812f
C1171 SDn_1.n12 VSS 0.0296f
C1172 SDn_1.t16 VSS 0.00812f
C1173 SDn_1.n13 VSS 0.00812f
C1174 SDn_1.n14 VSS 0.0223f
C1175 SDn_1.t6 VSS 0.00812f
C1176 SDn_1.n15 VSS 0.00812f
C1177 SDn_1.n16 VSS 0.0298f
C1178 SDn_1.n17 VSS 0.109f
C1179 SDn_1.n18 VSS 0.0306f
C1180 SDn_1.n19 VSS 0.0658f
C1181 SDn_1.t3 VSS 0.00812f
C1182 SDn_1.n20 VSS 0.00812f
C1183 SDn_1.n21 VSS 0.0163f
C1184 SDn_1.n22 VSS 0.0137f
C1185 SDn_1.n23 VSS 0.0292f
C1186 SDn_1.n24 VSS 0.03f
C1187 SDn_1.n25 VSS 0.066f
C1188 SDn_1.t28 VSS 0.00812f
C1189 SDn_1.n26 VSS 0.00812f
C1190 SDn_1.n27 VSS 0.0163f
C1191 SDn_1.n28 VSS 0.0137f
C1192 SDn_1.n29 VSS 0.0293f
C1193 SDn_1.t0 VSS 0.00812f
C1194 SDn_1.n30 VSS 0.00812f
C1195 SDn_1.n31 VSS 0.0223f
C1196 SDn_1.t31 VSS 0.00812f
C1197 SDn_1.n32 VSS 0.00812f
C1198 SDn_1.n33 VSS 0.0305f
C1199 SDn_1.n34 VSS 0.078f
C1200 SDn_1.n35 VSS 0.249f
C1201 SDn_1.t29 VSS 0.00812f
C1202 SDn_1.n36 VSS 0.00812f
C1203 SDn_1.n37 VSS 0.0223f
C1204 SDn_1.n38 VSS 0.232f
C1205 SDn_1.n39 VSS 0.00883f
C1206 SDn_1.t8 VSS 0.00751f
C1207 SDn_1.n40 VSS 0.0324f
C1208 SDn_1.n41 VSS 0.0943f
C1209 SDn_1.n42 VSS 0.0294f
C1210 SDn_1.n43 VSS 0.0654f
C1211 SDn_1.t7 VSS 0.00812f
C1212 SDn_1.n44 VSS 0.00812f
C1213 SDn_1.n45 VSS 0.0163f
C1214 SDn_1.n46 VSS 0.0137f
C1215 SDn_1.n47 VSS 0.0324f
C1216 SDn_1.t17 VSS 0.00812f
C1217 SDn_1.n48 VSS 0.00812f
C1218 SDn_1.n49 VSS 0.0163f
C1219 SDn_1.n50 VSS 0.0137f
C1220 SDn_1.n51 VSS 0.0317f
C1221 SDn_1.n52 VSS 0.065f
C1222 SDn_1.n53 VSS 0.0308f
C1223 SDn_1.n54 VSS 0.0689f
C1224 SDn_1.n55 VSS 0.0319f
C1225 b1b.n0 VSS 0.0068f
C1226 b1b.n1 VSS 0.00755f
C1227 b1b.n2 VSS 0.00752f
C1228 b1b.t2 VSS 0.0405f
C1229 b1b.n3 VSS 0.0317f
C1230 b1b.t4 VSS 0.00448f
C1231 b1b.n4 VSS 0.00585f
C1232 b1b.n5 VSS 0.5f
C1233 b1b.n6 VSS 0.0854f
C1234 b1b.n7 VSS 0.0389f
C1235 b1b.t3 VSS 0.0157f
C1236 SDc_1.n0 VSS 0.0101f
C1237 SDc_1.t9 VSS 0.00857f
C1238 SDc_1.n1 VSS 0.0352f
C1239 SDc_1.n2 VSS 0.0101f
C1240 SDc_1.t39 VSS 0.00857f
C1241 SDc_1.n3 VSS 0.0354f
C1242 SDc_1.t7 VSS 0.00927f
C1243 SDc_1.n4 VSS 0.00927f
C1244 SDc_1.n5 VSS 0.0334f
C1245 SDc_1.n6 VSS 0.0101f
C1246 SDc_1.t38 VSS 0.00857f
C1247 SDc_1.n7 VSS 0.0351f
C1248 SDc_1.n8 VSS 0.00998f
C1249 SDc_1.t30 VSS 0.00864f
C1250 SDc_1.n9 VSS 0.0353f
C1251 SDc_1.n10 VSS 0.0101f
C1252 SDc_1.t18 VSS 0.00857f
C1253 SDc_1.n11 VSS 0.0277f
C1254 SDc_1.t45 VSS 0.00927f
C1255 SDc_1.n12 VSS 0.00927f
C1256 SDc_1.n13 VSS 0.0333f
C1257 SDc_1.n14 VSS 0.00998f
C1258 SDc_1.t15 VSS 0.00864f
C1259 SDc_1.n15 VSS 0.0354f
C1260 SDc_1.n16 VSS 0.0101f
C1261 SDc_1.t50 VSS 0.00857f
C1262 SDc_1.n17 VSS 0.0353f
C1263 SDc_1.n18 VSS 0.0101f
C1264 SDc_1.t10 VSS 0.00857f
C1265 SDc_1.n19 VSS 0.0353f
C1266 SDc_1.n20 VSS 0.00998f
C1267 SDc_1.t44 VSS 0.00864f
C1268 SDc_1.n21 VSS 0.0393f
C1269 SDc_1.t41 VSS 0.00927f
C1270 SDc_1.n22 VSS 0.00927f
C1271 SDc_1.n23 VSS 0.0186f
C1272 SDc_1.n24 VSS 0.0155f
C1273 SDc_1.n25 VSS 0.0101f
C1274 SDc_1.t5 VSS 0.00857f
C1275 SDc_1.n26 VSS 0.0353f
C1276 SDc_1.n27 VSS 0.00998f
C1277 SDc_1.t36 VSS 0.00864f
C1278 SDc_1.n28 VSS 0.0355f
C1279 SDc_1.t48 VSS 0.00927f
C1280 SDc_1.n29 VSS 0.00927f
C1281 SDc_1.n30 VSS 0.0265f
C1282 SDc_1.n31 VSS 0.0101f
C1283 SDc_1.t11 VSS 0.00857f
C1284 SDc_1.n32 VSS 0.0353f
C1285 SDc_1.n33 VSS 0.0101f
C1286 SDc_1.t16 VSS 0.00857f
C1287 SDc_1.n34 VSS 0.0315f
C1288 SDc_1.n35 VSS 0.0101f
C1289 SDc_1.t42 VSS 0.00857f
C1290 SDc_1.n36 VSS 0.0358f
C1291 SDc_1.n37 VSS 0.12f
C1292 SDc_1.n38 VSS 0.103f
C1293 SDc_1.n39 VSS 0.0434f
C1294 SDc_1.n40 VSS 0.0369f
C1295 SDc_1.n41 VSS 0.0681f
C1296 SDc_1.n42 VSS 0.00998f
C1297 SDc_1.t12 VSS 0.00864f
C1298 SDc_1.n43 VSS 0.0185f
C1299 SDc_1.n44 VSS 0.0218f
C1300 SDc_1.n45 VSS 0.0333f
C1301 SDc_1.n46 VSS 0.0345f
C1302 SDc_1.n47 VSS 0.0702f
C1303 SDc_1.n48 VSS 0.0342f
C1304 SDc_1.n49 VSS 0.035f
C1305 SDc_1.n50 VSS 0.0713f
C1306 SDc_1.t17 VSS 0.00927f
C1307 SDc_1.n51 VSS 0.00927f
C1308 SDc_1.n52 VSS 0.0186f
C1309 SDc_1.n53 VSS 0.0155f
C1310 SDc_1.n54 VSS 0.035f
C1311 SDc_1.t47 VSS 0.00927f
C1312 SDc_1.n55 VSS 0.00927f
C1313 SDc_1.n56 VSS 0.0186f
C1314 SDc_1.n57 VSS 0.0155f
C1315 SDc_1.n58 VSS 0.0367f
C1316 SDc_1.n59 VSS 0.0674f
C1317 SDc_1.n60 VSS 0.0344f
C1318 SDc_1.n61 VSS 0.0337f
C1319 SDc_1.n62 VSS 0.0704f
C1320 SDc_1.t22 VSS 0.00927f
C1321 SDc_1.n63 VSS 0.00927f
C1322 SDc_1.n64 VSS 0.0186f
C1323 SDc_1.n65 VSS 0.0155f
C1324 SDc_1.n66 VSS 0.0349f
C1325 SDc_1.n67 VSS 0.0101f
C1326 SDc_1.t49 VSS 0.00857f
C1327 SDc_1.n68 VSS 0.0185f
C1328 SDc_1.n69 VSS 0.0155f
C1329 SDc_1.n70 VSS 0.0368f
C1330 SDc_1.n71 VSS 0.0675f
C1331 SDc_1.n72 VSS 0.0349f
C1332 SDc_1.n73 VSS 0.104f
C1333 SDc_1.n74 VSS 0.0427f
C1334 SDc_1.n75 VSS 0.0101f
C1335 SDc_1.t33 VSS 0.00857f
C1336 SDc_1.n76 VSS 0.0185f
C1337 SDc_1.n77 VSS 0.0155f
C1338 SDc_1.n78 VSS 0.037f
C1339 SDc_1.n79 VSS 0.0674f
C1340 SDc_1.n80 VSS 0.0353f
C1341 SDc_1.n81 VSS 0.0101f
C1342 SDc_1.t13 VSS 0.00857f
C1343 SDc_1.n82 VSS 0.0185f
C1344 SDc_1.n83 VSS 0.0155f
C1345 SDc_1.n84 VSS 0.0358f
C1346 SDc_1.n85 VSS 0.0668f
C1347 SDc_1.n86 VSS 0.0354f
C1348 SDc_1.n87 VSS 0.0358f
C1349 SDc_1.n88 VSS 0.0698f
C1350 SDc_1.n89 VSS 0.00998f
C1351 SDc_1.t43 VSS 0.00864f
C1352 SDc_1.n90 VSS 0.0185f
C1353 SDc_1.n91 VSS 0.0155f
C1354 SDc_1.n92 VSS 0.035f
C1355 SDc_1.n93 VSS 0.0364f
C1356 SDc_1.n94 VSS 0.0676f
C1357 SDc_1.n95 VSS 0.00998f
C1358 SDc_1.t14 VSS 0.00864f
C1359 SDc_1.n96 VSS 0.0185f
C1360 SDc_1.n97 VSS 0.0155f
C1361 SDc_1.n98 VSS 0.0349f
C1362 SDc_1.n99 VSS 0.0365f
C1363 SDc_1.n100 VSS 0.0647f
C1364 SDc_1.n101 VSS 0.00998f
C1365 SDc_1.t46 VSS 0.00864f
C1366 SDc_1.n102 VSS 0.0185f
C1367 SDc_1.n103 VSS 0.0155f
C1368 SDc_1.n104 VSS 2.49e-19
C1369 SDc_1.n105 VSS 0.00998f
C1370 SDc_1.t34 VSS 0.00864f
C1371 SDc_1.n106 VSS 0.0393f
C1372 SDc_1.n107 VSS 0.0101f
C1373 SDc_1.t40 VSS 0.00857f
C1374 SDc_1.n108 VSS 0.0278f
C1375 SDc_1.n109 VSS 0.00909f
C1376 SDc_1.n110 VSS 0.00927f
C1377 SDc_1.n111 VSS 0.00412f
C1378 SDc_1.n112 VSS 0.00359f
C1379 SDc_1.t4 VSS 0.00767f
C1380 SDc_1.n113 VSS 0.00694f
C1381 SDc_1.n114 VSS 0.0224f
C1382 SDc_1.n115 VSS 0.108f
C1383 SDc_1.n116 VSS 0.0101f
C1384 SDc_1.t8 VSS 0.00857f
C1385 SDc_1.n117 VSS 0.0185f
C1386 SDc_1.n118 VSS 0.0155f
C1387 SDc_1.n119 VSS 0.0353f
C1388 SDc_1.n120 VSS 0.0686f
C1389 SDc_1.n121 VSS 0.0354f
C1390 SDc_1.n122 VSS 0.0351f
C1391 b2b.t4 VSS 0.0158f
C1392 b2b.t6 VSS 0.0295f
C1393 b2b.n0 VSS 0.0536f
C1394 b2b.t3 VSS 0.0156f
C1395 b2b.n1 VSS 0.0317f
C1396 b2b.t2 VSS 0.0292f
C1397 b2b.n2 VSS 1.55f
C1398 b2b.n3 VSS 0.00819f
C1399 b2b.n4 VSS 0.00916f
C1400 b2b.n5 VSS 0.0899f
C1401 b2b.n6 VSS 0.0691f
C1402 b2b.t5 VSS 0.0194f
C1403 C32_U.t45 VSS 0.0122f
C1404 C32_U.n0 VSS 0.0122f
C1405 C32_U.n1 VSS 0.0273f
C1406 C32_U.t44 VSS 0.0404f
C1407 C32_U.t51 VSS 0.0122f
C1408 C32_U.n2 VSS 0.0122f
C1409 C32_U.n3 VSS 0.0664f
C1410 C32_U.t2 VSS 0.0341f
C1411 C32_U.n4 VSS 0.0682f
C1412 C32_U.t50 VSS 0.0404f
C1413 C32_U.t35 VSS 0.0122f
C1414 C32_U.n5 VSS 0.0122f
C1415 C32_U.n6 VSS 0.0268f
C1416 C32_U.n7 VSS 0.05f
C1417 C32_U.n8 VSS 0.0133f
C1418 C32_U.t55 VSS 0.0122f
C1419 C32_U.n9 VSS 0.0122f
C1420 C32_U.n10 VSS 0.0503f
C1421 C32_U.t54 VSS 0.0341f
C1422 C32_U.n11 VSS 0.0728f
C1423 C32_U.t26 VSS 0.0404f
C1424 C32_U.n12 VSS 0.0867f
C1425 C32_U.t36 VSS 0.0404f
C1426 C32_U.n13 VSS 0.0846f
C1427 C32_U.t37 VSS 0.0122f
C1428 C32_U.n14 VSS 0.0122f
C1429 C32_U.n15 VSS 0.0653f
C1430 C32_U.t0 VSS 0.0341f
C1431 C32_U.n16 VSS 0.0673f
C1432 C32_U.n17 VSS 0.0568f
C1433 C32_U.t40 VSS 0.0404f
C1434 C32_U.n18 VSS 0.0846f
C1435 C32_U.t41 VSS 0.0122f
C1436 C32_U.n19 VSS 0.0122f
C1437 C32_U.n20 VSS 0.0484f
C1438 C32_U.t14 VSS 0.0341f
C1439 C32_U.n21 VSS 0.0526f
C1440 C32_U.n22 VSS 0.0568f
C1441 C32_U.t56 VSS 0.0404f
C1442 C32_U.n23 VSS 0.0846f
C1443 C32_U.t57 VSS 0.0122f
C1444 C32_U.n24 VSS 0.0122f
C1445 C32_U.n25 VSS 0.0652f
C1446 C32_U.t28 VSS 0.0341f
C1447 C32_U.n26 VSS 0.0672f
C1448 C32_U.n27 VSS 0.0568f
C1449 C32_U.t38 VSS 0.0404f
C1450 C32_U.n28 VSS 0.0846f
C1451 C32_U.n29 VSS 0.0562f
C1452 C32_U.n30 VSS 0.00307f
C1453 C32_U.t39 VSS 0.0122f
C1454 C32_U.n31 VSS 0.0122f
C1455 C32_U.n32 VSS 0.0266f
C1456 C32_U.n33 VSS 0.0452f
C1457 C32_U.n34 VSS 0.00271f
C1458 C32_U.n35 VSS 0.00923f
C1459 C32_U.t12 VSS 0.0274f
C1460 C32_U.n36 VSS 0.0269f
C1461 C32_U.n37 VSS 0.0115f
C1462 C32_U.n38 VSS 0.0148f
C1463 C32_U.n39 VSS 0.217f
C1464 C32_U.t46 VSS 0.0441f
C1465 C32_U.t10 VSS 0.0351f
C1466 C32_U.t61 VSS 0.0122f
C1467 C32_U.n40 VSS 0.0122f
C1468 C32_U.n41 VSS 0.0658f
C1469 C32_U.n42 VSS 0.0714f
C1470 C32_U.t60 VSS 0.0441f
C1471 C32_U.t16 VSS 0.0351f
C1472 C32_U.t43 VSS 0.0122f
C1473 C32_U.n43 VSS 0.0122f
C1474 C32_U.n44 VSS 0.0658f
C1475 C32_U.n45 VSS 0.0714f
C1476 C32_U.t42 VSS 0.0441f
C1477 C32_U.t24 VSS 0.0351f
C1478 C32_U.t53 VSS 0.0122f
C1479 C32_U.n46 VSS 0.0122f
C1480 C32_U.n47 VSS 0.0658f
C1481 C32_U.n48 VSS 0.0714f
C1482 C32_U.t52 VSS 0.0441f
C1483 C32_U.n49 VSS 0.0884f
C1484 C32_U.n50 VSS 0.0596f
C1485 C32_U.n51 VSS 0.0884f
C1486 C32_U.n52 VSS 0.0596f
C1487 C32_U.n53 VSS 0.0884f
C1488 C32_U.n54 VSS 0.0596f
C1489 C32_U.n55 VSS 0.0884f
C1490 C32_U.n56 VSS 0.0578f
C1491 C32_U.n57 VSS 0.00735f
C1492 C32_U.t47 VSS 0.0122f
C1493 C32_U.n58 VSS 0.0122f
C1494 C32_U.n59 VSS 0.0273f
C1495 C32_U.n60 VSS 0.0462f
C1496 C32_U.n61 VSS 0.0186f
C1497 C32_U.t22 VSS 0.0282f
C1498 C32_U.n62 VSS 0.0276f
C1499 C32_U.n63 VSS 0.0116f
C1500 C32_U.n64 VSS 0.0071f
C1501 C32_U.n65 VSS 0.169f
C1502 C32_U.t30 VSS 0.0351f
C1503 C32_U.t31 VSS 0.0285f
C1504 C32_U.t66 VSS 0.0122f
C1505 C32_U.n66 VSS 0.0122f
C1506 C32_U.n67 VSS 0.0285f
C1507 C32_U.t81 VSS 0.0122f
C1508 C32_U.n68 VSS 0.0122f
C1509 C32_U.n69 VSS 0.0283f
C1510 C32_U.t68 VSS 0.0122f
C1511 C32_U.n70 VSS 0.0122f
C1512 C32_U.n71 VSS 0.0285f
C1513 C32_U.t93 VSS 0.0122f
C1514 C32_U.n72 VSS 0.0122f
C1515 C32_U.n73 VSS 0.0283f
C1516 C32_U.t95 VSS 0.0122f
C1517 C32_U.n74 VSS 0.0122f
C1518 C32_U.n75 VSS 0.0285f
C1519 C32_U.t69 VSS 0.0122f
C1520 C32_U.n76 VSS 0.0122f
C1521 C32_U.n77 VSS 0.0283f
C1522 C32_U.t92 VSS 0.0122f
C1523 C32_U.n78 VSS 0.0122f
C1524 C32_U.n79 VSS 0.0285f
C1525 C32_U.t64 VSS 0.0122f
C1526 C32_U.n80 VSS 0.0122f
C1527 C32_U.n81 VSS 0.0283f
C1528 C32_U.t73 VSS 0.0122f
C1529 C32_U.n82 VSS 0.0122f
C1530 C32_U.n83 VSS 0.0285f
C1531 C32_U.t75 VSS 0.0122f
C1532 C32_U.n84 VSS 0.0122f
C1533 C32_U.n85 VSS 0.0283f
C1534 C32_U.t91 VSS 0.0122f
C1535 C32_U.n86 VSS 0.0122f
C1536 C32_U.n87 VSS 0.0285f
C1537 C32_U.t71 VSS 0.0122f
C1538 C32_U.n88 VSS 0.0122f
C1539 C32_U.n89 VSS 0.0283f
C1540 C32_U.t87 VSS 0.0122f
C1541 C32_U.n90 VSS 0.0122f
C1542 C32_U.n91 VSS 0.0285f
C1543 C32_U.t72 VSS 0.0122f
C1544 C32_U.n92 VSS 0.0122f
C1545 C32_U.n93 VSS 0.0283f
C1546 C32_U.t83 VSS 0.0122f
C1547 C32_U.n94 VSS 0.0122f
C1548 C32_U.n95 VSS 0.0285f
C1549 C32_U.n96 VSS 0.0292f
C1550 C32_U.n97 VSS 0.0286f
C1551 C32_U.t4 VSS 0.0351f
C1552 C32_U.t8 VSS 0.0351f
C1553 C32_U.t49 VSS 0.0122f
C1554 C32_U.n98 VSS 0.0122f
C1555 C32_U.n99 VSS 0.0659f
C1556 C32_U.n100 VSS 0.0715f
C1557 C32_U.n101 VSS 0.0596f
C1558 C32_U.t48 VSS 0.0441f
C1559 C32_U.n102 VSS 0.09f
C1560 C32_U.n103 VSS 0.0891f
C1561 C32_U.n104 VSS 0.591f
C1562 C32_U.n105 VSS 0.669f
C1563 C32_U.n106 VSS 0.203f
C1564 C32_U.n107 VSS 0.221f
C1565 C32_U.n108 VSS 0.222f
C1566 C32_U.n109 VSS 0.221f
C1567 C32_U.n110 VSS 0.222f
C1568 C32_U.n111 VSS 0.221f
C1569 C32_U.n112 VSS 0.222f
C1570 C32_U.n113 VSS 0.221f
C1571 C32_U.n114 VSS 0.222f
C1572 C32_U.n115 VSS 0.221f
C1573 C32_U.n116 VSS 0.222f
C1574 C32_U.n117 VSS 0.221f
C1575 C32_U.n118 VSS 0.222f
C1576 C32_U.n119 VSS 0.221f
C1577 C32_U.n120 VSS 0.203f
C1578 C32_U.t77 VSS 0.0292f
C1579 C32_U.n121 VSS 0.667f
C1580 C32_U.n122 VSS 0.589f
C1581 C32_U.n123 VSS 0.0892f
C1582 C32_U.t62 VSS 0.0351f
C1583 C32_U.t33 VSS 0.0122f
C1584 C32_U.n124 VSS 0.0122f
C1585 C32_U.n125 VSS 0.0494f
C1586 C32_U.n126 VSS 0.0569f
C1587 C32_U.n127 VSS 0.0612f
C1588 C32_U.t32 VSS 0.0441f
C1589 C32_U.n128 VSS 0.0884f
C1590 C32_U.t58 VSS 0.0441f
C1591 C32_U.n129 VSS 0.0884f
C1592 C32_U.n130 VSS 0.06f
C1593 C32_U.t18 VSS 0.0342f
C1594 C32_U.n131 VSS 0.0383f
C1595 C32_U.t59 VSS 0.0122f
C1596 C32_U.n132 VSS 0.0122f
C1597 C32_U.n133 VSS 0.0282f
C1598 C32_U.n134 VSS 0.0711f
C1599 C32_U.n135 VSS 0.755f
C1600 C32_U.n136 VSS 0.15f
C1601 C32_U.n137 VSS 0.169f
C1602 C32_U.n138 VSS 0.00838f
C1603 C32_U.t6 VSS 0.0312f
C1604 C32_U.n139 VSS 0.0261f
C1605 C32_U.n140 VSS 0.0115f
C1606 C32_U.t34 VSS 0.0404f
C1607 C32_U.n142 VSS 0.0846f
C1608 C32_U.n143 VSS 0.0562f
C1609 C32_U.n144 VSS 0.0846f
C1610 C32_U.n145 VSS 0.0568f
C1611 C32_U.n146 VSS 0.0867f
C1612 C32_U.t20 VSS 0.0341f
C1613 C32_U.n147 VSS 0.0527f
C1614 C32_U.n148 VSS 0.0567f
C1615 b5.t11 VSS 0.0191f
C1616 b5.t5 VSS 0.0149f
C1617 b5.t8 VSS 0.0149f
C1618 b5.t22 VSS 0.0151f
C1619 b5.n0 VSS 0.0315f
C1620 b5.t17 VSS 0.0149f
C1621 b5.n1 VSS 0.0317f
C1622 b5.t7 VSS 0.0953f
C1623 b5.t19 VSS 0.0951f
C1624 b5.n2 VSS 0.0315f
C1625 b5.t15 VSS 0.0149f
C1626 b5.n3 VSS 0.0317f
C1627 b5.t4 VSS 0.0607f
C1628 b5.t25 VSS 0.0185f
C1629 b5.t14 VSS 0.0142f
C1630 b5.t9 VSS 0.0282f
C1631 b5.t6 VSS 0.0571f
C1632 b5.t18 VSS 0.0282f
C1633 b5.t16 VSS 0.0546f
C1634 b5.t13 VSS 0.0198f
C1635 b5.n4 VSS 0.05f
C1636 b5.t21 VSS 0.0198f
C1637 b5.n5 VSS 0.0346f
C1638 b5.n6 VSS 0.034f
C1639 b5.t26 VSS 0.0308f
C1640 b5.t3 VSS 0.0139f
C1641 b5.n7 VSS 0.0329f
C1642 b5.t24 VSS 0.0139f
C1643 b5.n8 VSS 0.0329f
C1644 b5.t20 VSS 0.0308f
C1645 b5.n9 VSS 0.034f
C1646 b5.t12 VSS 0.0198f
C1647 b5.n10 VSS 0.0369f
C1648 b5.t2 VSS 0.00794f
C1649 b5.n11 VSS 0.133f
C1650 b5.n12 VSS 0.0778f
C1651 b5.t23 VSS 0.0195f
C1652 b5.n13 VSS 0.0673f
C1653 b5.t10 VSS 0.0195f
C1654 b5.n14 VSS 0.0654f
C1655 b5.n15 VSS 0.0344f
C1656 b5.n16 VSS 0.365f
C1657 b5.t0 VSS 0.00597f
C1658 b5.t1 VSS 0.00472f
C1659 b5.n17 VSS 0.0923f
C1660 b5.n18 VSS 0.168f
C1661 OUT4.n0 VSS 0.0146f
C1662 OUT4.n1 VSS 0.0124f
C1663 OUT4.n2 VSS 0.0464f
C1664 OUT4.n3 VSS 0.0124f
C1665 OUT4.n4 VSS 0.0124f
C1666 OUT4.t15 VSS 0.0147f
C1667 OUT4.t14 VSS 0.0124f
C1668 OUT4.n5 VSS 0.0986f
C1669 OUT4.n6 VSS 0.0701f
C1670 OUT4.n7 VSS 0.0384f
C1671 OUT4.t7 VSS 0.00542f
C1672 OUT4.n8 VSS 0.00542f
C1673 OUT4.n9 VSS 0.0108f
C1674 OUT4.t23 VSS 0.00542f
C1675 OUT4.n10 VSS 0.00542f
C1676 OUT4.n11 VSS 0.0108f
C1677 OUT4.t17 VSS 0.00542f
C1678 OUT4.n12 VSS 0.00542f
C1679 OUT4.n13 VSS 0.0108f
C1680 OUT4.t4 VSS 0.00542f
C1681 OUT4.n14 VSS 0.00542f
C1682 OUT4.n15 VSS 0.0147f
C1683 OUT4.n16 VSS 0.0475f
C1684 OUT4.n17 VSS 0.0297f
C1685 OUT4.n18 VSS 0.0433f
C1686 OUT4.t22 VSS 0.00542f
C1687 OUT4.n19 VSS 0.00542f
C1688 OUT4.n20 VSS 0.0108f
C1689 OUT4.t3 VSS 0.00542f
C1690 OUT4.n21 VSS 0.00542f
C1691 OUT4.n22 VSS 0.0108f
C1692 OUT4.t0 VSS 0.00542f
C1693 OUT4.n23 VSS 0.00542f
C1694 OUT4.n24 VSS 0.0108f
C1695 OUT4.t19 VSS 0.00542f
C1696 OUT4.n25 VSS 0.00542f
C1697 OUT4.n26 VSS 0.0145f
C1698 OUT4.n27 VSS 0.0454f
C1699 OUT4.n28 VSS 0.0289f
C1700 OUT4.n29 VSS 0.0203f
C1701 OUT4.n30 VSS 0.366f
C1702 OUT4.n31 VSS 0.678f
C1703 OUT4.t12 VSS 0.0124f
C1704 OUT4.n32 VSS 0.188f
C1705 OUT4.t9 VSS 0.0124f
C1706 OUT4.n33 VSS 0.0613f
C1707 b4b.t5 VSS 0.0217f
C1708 b4b.t15 VSS 0.0237f
C1709 b4b.n0 VSS 0.0437f
C1710 b4b.t17 VSS 0.0237f
C1711 b4b.n1 VSS 0.0437f
C1712 b4b.t13 VSS 0.0821f
C1713 b4b.t10 VSS 0.161f
C1714 b4b.t2 VSS 0.0386f
C1715 b4b.n2 VSS 0.151f
C1716 b4b.t8 VSS 0.112f
C1717 b4b.n3 VSS 0.16f
C1718 b4b.t3 VSS 0.0986f
C1719 b4b.t7 VSS 0.0817f
C1720 b4b.t18 VSS 0.0132f
C1721 b4b.n4 VSS 0.0407f
C1722 b4b.t14 VSS 0.0124f
C1723 b4b.n5 VSS 0.0367f
C1724 b4b.t4 VSS 0.0738f
C1725 b4b.t12 VSS 0.184f
C1726 b4b.t6 VSS 0.0298f
C1727 b4b.n6 VSS 0.222f
C1728 b4b.t16 VSS 0.0976f
C1729 b4b.t11 VSS 0.0369f
C1730 b4b.n7 VSS 0.0917f
C1731 b4b.n8 VSS 0.74f
C1732 b4b.n9 VSS 1.15f
C1733 b4b.n11 VSS 0.00307f
C1734 b4b.n12 VSS 0.0118f
C1735 b4b.n13 VSS 0.00771f
C1736 b4b.n14 VSS 0.00293f
C1737 b4b.n15 VSS 0.0103f
C1738 b4b.n16 VSS 0.00858f
C1739 b4b.n17 VSS 0.0672f
C1740 b4b.n18 VSS 0.0436f
C1741 b4b.n19 VSS 0.00866f
C1742 b4b.t9 VSS 0.0178f
C1743 SDc_2.t11 VSS 0.0142f
C1744 SDc_2.n0 VSS 0.0142f
C1745 SDc_2.n1 VSS 0.0593f
C1746 SDc_2.t48 VSS 0.0142f
C1747 SDc_2.n2 VSS 0.0142f
C1748 SDc_2.n3 VSS 0.0287f
C1749 SDc_2.n4 VSS 0.0328f
C1750 SDc_2.t50 VSS 0.0142f
C1751 SDc_2.n5 VSS 0.0142f
C1752 SDc_2.n6 VSS 0.0578f
C1753 SDc_2.t51 VSS 0.0142f
C1754 SDc_2.n7 VSS 0.0142f
C1755 SDc_2.n8 VSS 0.0288f
C1756 SDc_2.n9 VSS 0.0353f
C1757 SDc_2.t3 VSS 0.0142f
C1758 SDc_2.n10 VSS 0.0142f
C1759 SDc_2.n11 VSS 0.0587f
C1760 SDc_2.t15 VSS 0.0142f
C1761 SDc_2.n12 VSS 0.0142f
C1762 SDc_2.n13 VSS 0.0288f
C1763 SDc_2.n14 VSS 0.0348f
C1764 SDc_2.t62 VSS 0.0142f
C1765 SDc_2.n15 VSS 0.0142f
C1766 SDc_2.n16 VSS 0.0586f
C1767 SDc_2.t53 VSS 0.0142f
C1768 SDc_2.n17 VSS 0.0142f
C1769 SDc_2.n18 VSS 0.0474f
C1770 SDc_2.t30 VSS 0.0142f
C1771 SDc_2.n19 VSS 0.0142f
C1772 SDc_2.n20 VSS 0.0588f
C1773 SDc_2.t6 VSS 0.0142f
C1774 SDc_2.n21 VSS 0.0142f
C1775 SDc_2.n22 VSS 0.047f
C1776 SDc_2.t52 VSS 0.0142f
C1777 SDc_2.n23 VSS 0.0142f
C1778 SDc_2.n24 VSS 0.0588f
C1779 SDc_2.t13 VSS 0.0142f
C1780 SDc_2.n25 VSS 0.0142f
C1781 SDc_2.n26 VSS 0.0589f
C1782 SDc_2.t12 VSS 0.0142f
C1783 SDc_2.n27 VSS 0.0142f
C1784 SDc_2.n28 VSS 0.0287f
C1785 SDc_2.n29 VSS 0.034f
C1786 SDc_2.t54 VSS 0.0142f
C1787 SDc_2.n30 VSS 0.0142f
C1788 SDc_2.n31 VSS 0.0587f
C1789 SDc_2.t56 VSS 0.0142f
C1790 SDc_2.n32 VSS 0.0142f
C1791 SDc_2.n33 VSS 0.0287f
C1792 SDc_2.n34 VSS 0.0336f
C1793 SDc_2.t29 VSS 0.0142f
C1794 SDc_2.n35 VSS 0.0142f
C1795 SDc_2.n36 VSS 0.0588f
C1796 SDc_2.t61 VSS 0.0142f
C1797 SDc_2.n37 VSS 0.0142f
C1798 SDc_2.n38 VSS 0.058f
C1799 SDc_2.t10 VSS 0.0142f
C1800 SDc_2.n39 VSS 0.0142f
C1801 SDc_2.n40 VSS 0.0592f
C1802 SDc_2.t23 VSS 0.0142f
C1803 SDc_2.n41 VSS 0.0142f
C1804 SDc_2.n42 VSS 0.0287f
C1805 SDc_2.n43 VSS 0.0324f
C1806 SDc_2.t58 VSS 0.0142f
C1807 SDc_2.n44 VSS 0.0142f
C1808 SDc_2.n45 VSS 0.059f
C1809 SDc_2.t55 VSS 0.0142f
C1810 SDc_2.n46 VSS 0.0142f
C1811 SDc_2.n47 VSS 0.0288f
C1812 SDc_2.n48 VSS 0.0344f
C1813 SDc_2.t21 VSS 0.0142f
C1814 SDc_2.n49 VSS 0.0142f
C1815 SDc_2.n50 VSS 0.0587f
C1816 SDc_2.t19 VSS 0.0142f
C1817 SDc_2.n51 VSS 0.0142f
C1818 SDc_2.n52 VSS 0.0474f
C1819 SDc_2.t63 VSS 0.0142f
C1820 SDc_2.n53 VSS 0.0142f
C1821 SDc_2.n54 VSS 0.0588f
C1822 SDc_2.t59 VSS 0.0142f
C1823 SDc_2.n55 VSS 0.0142f
C1824 SDc_2.n56 VSS 0.0446f
C1825 SDc_2.t18 VSS 0.0142f
C1826 SDc_2.n57 VSS 0.0142f
C1827 SDc_2.n58 VSS 0.0586f
C1828 SDc_2.n59 VSS 0.216f
C1829 SDc_2.n60 VSS 0.186f
C1830 SDc_2.n61 VSS 0.0673f
C1831 SDc_2.n62 VSS 0.0523f
C1832 SDc_2.n63 VSS 0.134f
C1833 SDc_2.n64 VSS 0.0523f
C1834 SDc_2.n65 VSS 0.0529f
C1835 SDc_2.n66 VSS 0.136f
C1836 SDc_2.n67 VSS 0.0525f
C1837 SDc_2.n68 VSS 0.0527f
C1838 SDc_2.n69 VSS 0.137f
C1839 SDc_2.t57 VSS 0.0142f
C1840 SDc_2.n70 VSS 0.0142f
C1841 SDc_2.n71 VSS 0.0287f
C1842 SDc_2.n72 VSS 0.0328f
C1843 SDc_2.n73 VSS 0.0514f
C1844 SDc_2.n74 VSS 0.0516f
C1845 SDc_2.n75 VSS 0.137f
C1846 SDc_2.t17 VSS 0.0142f
C1847 SDc_2.n76 VSS 0.0142f
C1848 SDc_2.n77 VSS 0.0287f
C1849 SDc_2.n78 VSS 0.0328f
C1850 SDc_2.n79 VSS 0.0508f
C1851 SDc_2.n80 VSS 0.052f
C1852 SDc_2.n81 VSS 0.135f
C1853 SDc_2.n82 VSS 0.0522f
C1854 SDc_2.n83 VSS 0.0526f
C1855 SDc_2.n84 VSS 0.134f
C1856 SDc_2.n85 VSS 0.0517f
C1857 SDc_2.n86 VSS 0.0527f
C1858 SDc_2.n87 VSS 0.135f
C1859 SDc_2.t60 VSS 0.0142f
C1860 SDc_2.n88 VSS 0.0142f
C1861 SDc_2.n89 VSS 0.0287f
C1862 SDc_2.n90 VSS 0.0328f
C1863 SDc_2.n91 VSS 0.0538f
C1864 SDc_2.n92 VSS 0.186f
C1865 SDc_2.n93 VSS 0.0691f
C1866 SDc_2.n94 VSS 0.186f
C1867 SDc_2.n95 VSS 0.067f
C1868 SDc_2.n96 VSS 0.0528f
C1869 SDc_2.n97 VSS 0.134f
C1870 SDc_2.n98 VSS 0.0512f
C1871 SDc_2.n99 VSS 0.0526f
C1872 SDc_2.n100 VSS 0.134f
C1873 SDc_2.n101 VSS 0.0542f
C1874 SDc_2.n102 VSS 0.0554f
C1875 SDc_2.n103 VSS 0.132f
C1876 SDc_2.t26 VSS 0.0142f
C1877 SDc_2.n104 VSS 0.0142f
C1878 SDc_2.n105 VSS 0.0287f
C1879 SDc_2.n106 VSS 0.034f
C1880 SDc_2.n107 VSS 0.0522f
C1881 SDc_2.n108 VSS 0.0521f
C1882 SDc_2.t49 VSS 0.0142f
C1883 SDc_2.n109 VSS 0.0142f
C1884 SDc_2.n110 VSS 0.0598f
C1885 SDc_2.t2 VSS 0.0142f
C1886 SDc_2.n111 VSS 0.0142f
C1887 SDc_2.n112 VSS 0.0285f
C1888 SDc_2.n113 VSS 0.0244f
C1889 SDc_2.n114 VSS 0.197f
C1890 SDc_2.n115 VSS 0.053f
C1891 Gc_2.t71 VSS 0.0328f
C1892 Gc_2.n0 VSS 0.0328f
C1893 Gc_2.n1 VSS 0.0656f
C1894 Gc_2.n2 VSS 0.121f
C1895 Gc_2.t76 VSS 0.0328f
C1896 Gc_2.n3 VSS 0.0328f
C1897 Gc_2.n4 VSS 0.0656f
C1898 Gc_2.t15 VSS 0.0328f
C1899 Gc_2.n5 VSS 0.0328f
C1900 Gc_2.n6 VSS 0.0706f
C1901 Gc_2.t49 VSS 0.0328f
C1902 Gc_2.n7 VSS 0.0328f
C1903 Gc_2.n8 VSS 0.084f
C1904 Gc_2.t79 VSS 0.0328f
C1905 Gc_2.n9 VSS 0.0328f
C1906 Gc_2.n10 VSS 0.0656f
C1907 Gc_2.t60 VSS 0.0862f
C1908 Gc_2.t14 VSS 0.0967f
C1909 Gc_2.n11 VSS 0.225f
C1910 Gc_2.n12 VSS 0.0616f
C1911 Gc_2.n13 VSS 0.0933f
C1912 Gc_2.n14 VSS 0.00566f
C1913 Gc_2.n15 VSS 0.105f
C1914 Gc_2.n16 VSS 0.0285f
C1915 Gc_2.n17 VSS 0.0117f
C1916 Gc_2.n18 VSS 0.133f
C1917 Gc_2.t35 VSS 0.0328f
C1918 Gc_2.n19 VSS 0.0328f
C1919 Gc_2.n20 VSS 0.0706f
C1920 Gc_2.t48 VSS 0.107f
C1921 Gc_2.n21 VSS 0.234f
C1922 Gc_2.n22 VSS 0.189f
C1923 Gc_2.t0 VSS 0.0925f
C1924 Gc_2.n23 VSS 0.0931f
C1925 Gc_2.t84 VSS 0.0328f
C1926 Gc_2.n24 VSS 0.0328f
C1927 Gc_2.n25 VSS 0.0656f
C1928 Gc_2.n26 VSS 0.176f
C1929 Gc_2.t29 VSS 0.0328f
C1930 Gc_2.n27 VSS 0.0328f
C1931 Gc_2.n28 VSS 0.084f
C1932 Gc_2.t69 VSS 0.0328f
C1933 Gc_2.n29 VSS 0.0328f
C1934 Gc_2.n30 VSS 0.0656f
C1935 Gc_2.t6 VSS 0.0867f
C1936 Gc_2.t34 VSS 0.0967f
C1937 Gc_2.n31 VSS 0.221f
C1938 Gc_2.n32 VSS 0.0613f
C1939 Gc_2.n33 VSS 0.0929f
C1940 Gc_2.n34 VSS 0.00577f
C1941 Gc_2.n35 VSS 0.104f
C1942 Gc_2.n36 VSS 0.0295f
C1943 Gc_2.n37 VSS 0.0122f
C1944 Gc_2.n38 VSS 0.14f
C1945 Gc_2.t51 VSS 0.0328f
C1946 Gc_2.n39 VSS 0.0328f
C1947 Gc_2.n40 VSS 0.0706f
C1948 Gc_2.t28 VSS 0.107f
C1949 Gc_2.n41 VSS 0.233f
C1950 Gc_2.n42 VSS 0.196f
C1951 Gc_2.t18 VSS 0.0919f
C1952 Gc_2.n43 VSS 0.0855f
C1953 Gc_2.t92 VSS 0.0328f
C1954 Gc_2.n44 VSS 0.0328f
C1955 Gc_2.n45 VSS 0.0656f
C1956 Gc_2.n46 VSS 0.162f
C1957 Gc_2.t41 VSS 0.0328f
C1958 Gc_2.n47 VSS 0.0328f
C1959 Gc_2.n48 VSS 0.084f
C1960 Gc_2.t77 VSS 0.0328f
C1961 Gc_2.n49 VSS 0.0328f
C1962 Gc_2.n50 VSS 0.0656f
C1963 Gc_2.t2 VSS 0.0862f
C1964 Gc_2.t50 VSS 0.0967f
C1965 Gc_2.n51 VSS 0.221f
C1966 Gc_2.n52 VSS 0.0615f
C1967 Gc_2.n53 VSS 0.0942f
C1968 Gc_2.n54 VSS 0.00602f
C1969 Gc_2.n55 VSS 0.104f
C1970 Gc_2.n56 VSS 0.0295f
C1971 Gc_2.n57 VSS 0.0121f
C1972 Gc_2.n58 VSS 0.166f
C1973 Gc_2.t43 VSS 0.0328f
C1974 Gc_2.n59 VSS 0.0328f
C1975 Gc_2.n60 VSS 0.0706f
C1976 Gc_2.t40 VSS 0.107f
C1977 Gc_2.n61 VSS 0.232f
C1978 Gc_2.n62 VSS 0.194f
C1979 Gc_2.t20 VSS 0.0919f
C1980 Gc_2.n63 VSS 0.0865f
C1981 Gc_2.t89 VSS 0.0328f
C1982 Gc_2.n64 VSS 0.0328f
C1983 Gc_2.n65 VSS 0.0656f
C1984 Gc_2.n66 VSS 0.163f
C1985 Gc_2.t55 VSS 0.0328f
C1986 Gc_2.n67 VSS 0.0328f
C1987 Gc_2.n68 VSS 0.084f
C1988 Gc_2.t82 VSS 0.0328f
C1989 Gc_2.n69 VSS 0.0328f
C1990 Gc_2.n70 VSS 0.0656f
C1991 Gc_2.t24 VSS 0.0862f
C1992 Gc_2.t42 VSS 0.0967f
C1993 Gc_2.n71 VSS 0.221f
C1994 Gc_2.n72 VSS 0.0616f
C1995 Gc_2.n73 VSS 0.0927f
C1996 Gc_2.n74 VSS 0.00543f
C1997 Gc_2.n75 VSS 0.105f
C1998 Gc_2.n76 VSS 0.0279f
C1999 Gc_2.n77 VSS 0.00871f
C2000 Gc_2.n78 VSS 0.103f
C2001 Gc_2.t45 VSS 0.0328f
C2002 Gc_2.n79 VSS 0.0328f
C2003 Gc_2.n80 VSS 0.0706f
C2004 Gc_2.t54 VSS 0.107f
C2005 Gc_2.n81 VSS 0.233f
C2006 Gc_2.n82 VSS 0.197f
C2007 Gc_2.t16 VSS 0.0909f
C2008 Gc_2.n83 VSS 0.0862f
C2009 Gc_2.t90 VSS 0.0328f
C2010 Gc_2.n84 VSS 0.0328f
C2011 Gc_2.n85 VSS 0.0656f
C2012 Gc_2.n86 VSS 0.163f
C2013 Gc_2.t63 VSS 0.0328f
C2014 Gc_2.n87 VSS 0.0328f
C2015 Gc_2.n88 VSS 0.084f
C2016 Gc_2.t88 VSS 0.0328f
C2017 Gc_2.n89 VSS 0.0328f
C2018 Gc_2.n90 VSS 0.0656f
C2019 Gc_2.t10 VSS 0.0862f
C2020 Gc_2.t44 VSS 0.0967f
C2021 Gc_2.n91 VSS 0.222f
C2022 Gc_2.n92 VSS 0.0615f
C2023 Gc_2.n93 VSS 0.0948f
C2024 Gc_2.n94 VSS 0.00625f
C2025 Gc_2.n95 VSS 0.104f
C2026 Gc_2.n96 VSS 0.0301f
C2027 Gc_2.n97 VSS 0.0139f
C2028 Gc_2.n98 VSS 0.164f
C2029 Gc_2.t37 VSS 0.0328f
C2030 Gc_2.n99 VSS 0.0328f
C2031 Gc_2.n100 VSS 0.0706f
C2032 Gc_2.t32 VSS 0.187f
C2033 Gc_2.t56 VSS 0.107f
C2034 Gc_2.n101 VSS 0.278f
C2035 Gc_2.t62 VSS 0.107f
C2036 Gc_2.n102 VSS 0.233f
C2037 Gc_2.n103 VSS 0.199f
C2038 Gc_2.t26 VSS 0.0909f
C2039 Gc_2.n104 VSS 0.0843f
C2040 Gc_2.t86 VSS 0.0328f
C2041 Gc_2.n105 VSS 0.0328f
C2042 Gc_2.n106 VSS 0.0656f
C2043 Gc_2.n107 VSS 0.163f
C2044 Gc_2.t57 VSS 0.0328f
C2045 Gc_2.n108 VSS 0.0328f
C2046 Gc_2.n109 VSS 0.084f
C2047 Gc_2.t83 VSS 0.0328f
C2048 Gc_2.n110 VSS 0.0328f
C2049 Gc_2.n111 VSS 0.0656f
C2050 Gc_2.t46 VSS 0.287f
C2051 Gc_2.n112 VSS 0.138f
C2052 Gc_2.n113 VSS 0.0138f
C2053 Gc_2.t12 VSS 0.0872f
C2054 Gc_2.t36 VSS 0.0967f
C2055 Gc_2.n114 VSS 0.22f
C2056 Gc_2.n115 VSS 0.0591f
C2057 Gc_2.n116 VSS 0.0216f
C2058 Gc_2.n117 VSS 0.0709f
C2059 Gc_2.n118 VSS 0.0356f
C2060 Gc_2.t127 VSS 0.097f
C2061 Gc_2.t121 VSS 0.107f
C2062 Gc_2.n119 VSS 0.233f
C2063 Gc_2.t140 VSS 0.107f
C2064 Gc_2.n120 VSS 0.233f
C2065 Gc_2.t113 VSS 0.107f
C2066 Gc_2.n121 VSS 0.233f
C2067 Gc_2.t96 VSS 0.107f
C2068 Gc_2.n122 VSS 0.233f
C2069 Gc_2.t106 VSS 0.107f
C2070 Gc_2.n123 VSS 0.233f
C2071 Gc_2.t134 VSS 0.107f
C2072 Gc_2.n124 VSS 0.233f
C2073 Gc_2.t111 VSS 0.107f
C2074 Gc_2.n125 VSS 0.236f
C2075 Gc_2.n126 VSS 0.364f
C2076 Gc_2.n127 VSS 0.568f
C2077 Gc_2.n128 VSS 0.0835f
C2078 Gc_2.t91 VSS 0.0328f
C2079 Gc_2.n129 VSS 0.0328f
C2080 Gc_2.n130 VSS 0.084f
C2081 Gc_2.t47 VSS 0.0328f
C2082 Gc_2.n131 VSS 0.0328f
C2083 Gc_2.n132 VSS 0.0706f
C2084 Gc_2.n133 VSS 0.436f
C2085 Gc_2.n134 VSS 0.54f
C2086 Gc_2.n135 VSS 0.512f
C2087 Gc_2.n136 VSS 0.54f
C2088 Gc_2.n137 VSS 0.512f
C2089 Gc_2.n138 VSS 0.54f
C2090 Gc_2.n139 VSS 0.512f
C2091 Gc_2.n140 VSS 0.54f
C2092 Gc_2.n141 VSS 0.512f
C2093 Gc_2.n142 VSS 0.54f
C2094 Gc_2.n143 VSS 0.512f
C2095 Gc_2.n144 VSS 0.54f
C2096 Gc_2.t9 VSS 0.0328f
C2097 Gc_2.n145 VSS 0.0328f
C2098 Gc_2.n146 VSS 0.084f
C2099 Gc_2.t94 VSS 0.0328f
C2100 Gc_2.n147 VSS 0.0328f
C2101 Gc_2.n148 VSS 0.0656f
C2102 Gc_2.n149 VSS 0.0599f
C2103 Gc_2.t38 VSS 0.0877f
C2104 Gc_2.n150 VSS 0.0934f
C2105 Gc_2.n151 VSS 0.122f
C2106 Gc_2.n152 VSS 0.0156f
C2107 Gc_2.t108 VSS 0.107f
C2108 Gc_2.t101 VSS 0.107f
C2109 Gc_2.t115 VSS 0.107f
C2110 Gc_2.t116 VSS 0.107f
C2111 Gc_2.t104 VSS 0.107f
C2112 Gc_2.t132 VSS 0.107f
C2113 Gc_2.t143 VSS 0.107f
C2114 Gc_2.n153 VSS 0.233f
C2115 Gc_2.n154 VSS 0.233f
C2116 Gc_2.n155 VSS 0.233f
C2117 Gc_2.n156 VSS 0.233f
C2118 Gc_2.n157 VSS 0.233f
C2119 Gc_2.n158 VSS 0.233f
C2120 Gc_2.n159 VSS 0.235f
C2121 Gc_2.t139 VSS 0.101f
C2122 Gc_2.n160 VSS 0.215f
C2123 Gc_2.t112 VSS 0.295f
C2124 Gc_2.t124 VSS 0.107f
C2125 Gc_2.n161 VSS 0.257f
C2126 Gc_2.t109 VSS 0.107f
C2127 Gc_2.n162 VSS 0.233f
C2128 Gc_2.t100 VSS 0.107f
C2129 Gc_2.n163 VSS 0.233f
C2130 Gc_2.t123 VSS 0.107f
C2131 Gc_2.n164 VSS 0.233f
C2132 Gc_2.t110 VSS 0.107f
C2133 Gc_2.n165 VSS 0.233f
C2134 Gc_2.t98 VSS 0.107f
C2135 Gc_2.n166 VSS 0.233f
C2136 Gc_2.t117 VSS 0.107f
C2137 Gc_2.n167 VSS 0.233f
C2138 Gc_2.t119 VSS 0.107f
C2139 Gc_2.n168 VSS 0.233f
C2140 Gc_2.t99 VSS 0.107f
C2141 Gc_2.n169 VSS 0.233f
C2142 Gc_2.t97 VSS 0.107f
C2143 Gc_2.n170 VSS 0.233f
C2144 Gc_2.t126 VSS 0.107f
C2145 Gc_2.n171 VSS 0.233f
C2146 Gc_2.t138 VSS 0.107f
C2147 Gc_2.n172 VSS 0.233f
C2148 Gc_2.t105 VSS 0.107f
C2149 Gc_2.n173 VSS 0.233f
C2150 Gc_2.t122 VSS 0.107f
C2151 Gc_2.n174 VSS 0.227f
C2152 Gc_2.t137 VSS 0.106f
C2153 Gc_2.n175 VSS 0.404f
C2154 Gc_2.n176 VSS 1.04f
C2155 Gc_2.n177 VSS 0.33f
C2156 Gc_2.n178 VSS 0.0445f
C2157 Gc_2.n179 VSS 0.0303f
C2158 Gc_2.n180 VSS 0.0246f
C2159 Gc_2.n181 VSS 0.0477f
C2160 Gc_2.n182 VSS 0.0804f
C2161 Gc_2.t5 VSS 0.0328f
C2162 Gc_2.n183 VSS 0.0328f
C2163 Gc_2.n184 VSS 0.0706f
C2164 Gc_2.t23 VSS 0.0328f
C2165 Gc_2.n185 VSS 0.0328f
C2166 Gc_2.n186 VSS 0.084f
C2167 Gc_2.t66 VSS 0.0328f
C2168 Gc_2.n187 VSS 0.0328f
C2169 Gc_2.n188 VSS 0.0656f
C2170 Gc_2.t4 VSS 0.0967f
C2171 Gc_2.n189 VSS 0.23f
C2172 Gc_2.t30 VSS 0.103f
C2173 Gc_2.n190 VSS 0.254f
C2174 Gc_2.n191 VSS 0.176f
C2175 Gc_2.n192 VSS 0.382f
C2176 Gc_2.n193 VSS 0.417f
C2177 Gc_2.n194 VSS 0.457f
C2178 Gc_2.n195 VSS 0.512f
C2179 Gc_2.n196 VSS 0.177f
C2180 Gc_2.t52 VSS 0.0935f
C2181 Gc_2.n197 VSS 0.0887f
C2182 Gc_2.n198 VSS 0.186f
C2183 Gc_2.t8 VSS 0.107f
C2184 Gc_2.n199 VSS 0.233f
C2185 Gc_2.t22 VSS 0.192f
C2186 Gc_2.n200 VSS 0.238f
C2187 Gc_2.t58 VSS 0.0935f
C2188 Gc_2.n201 VSS 0.0772f
C2189 Gc_2.n202 VSS 0.0394f
C2190 Gc_1.n0 VSS 0.031f
C2191 Gc_1.t87 VSS 0.0229f
C2192 Gc_1.n1 VSS 0.0547f
C2193 Gc_1.t29 VSS 0.0551f
C2194 Gc_1.t24 VSS 0.0229f
C2195 Gc_1.n2 VSS 0.0229f
C2196 Gc_1.n3 VSS 0.0496f
C2197 Gc_1.t25 VSS 0.0229f
C2198 Gc_1.n4 VSS 0.0229f
C2199 Gc_1.n5 VSS 0.0491f
C2200 Gc_1.t20 VSS 0.0229f
C2201 Gc_1.n6 VSS 0.0229f
C2202 Gc_1.n7 VSS 0.0496f
C2203 Gc_1.t23 VSS 0.0229f
C2204 Gc_1.n8 VSS 0.0229f
C2205 Gc_1.n9 VSS 0.0491f
C2206 Gc_1.t27 VSS 0.0229f
C2207 Gc_1.n10 VSS 0.0229f
C2208 Gc_1.n11 VSS 0.0496f
C2209 Gc_1.t30 VSS 0.0229f
C2210 Gc_1.n12 VSS 0.0229f
C2211 Gc_1.n13 VSS 0.0491f
C2212 Gc_1.t15 VSS 0.0229f
C2213 Gc_1.n14 VSS 0.0229f
C2214 Gc_1.n15 VSS 0.0496f
C2215 Gc_1.t19 VSS 0.0229f
C2216 Gc_1.n16 VSS 0.0229f
C2217 Gc_1.n17 VSS 0.0491f
C2218 Gc_1.t17 VSS 0.0229f
C2219 Gc_1.n18 VSS 0.0229f
C2220 Gc_1.n19 VSS 0.0496f
C2221 Gc_1.t18 VSS 0.0229f
C2222 Gc_1.n20 VSS 0.0229f
C2223 Gc_1.n21 VSS 0.0491f
C2224 Gc_1.t21 VSS 0.0229f
C2225 Gc_1.n22 VSS 0.0229f
C2226 Gc_1.n23 VSS 0.0496f
C2227 Gc_1.t28 VSS 0.0229f
C2228 Gc_1.n24 VSS 0.0229f
C2229 Gc_1.n25 VSS 0.0491f
C2230 Gc_1.t26 VSS 0.0229f
C2231 Gc_1.n26 VSS 0.0229f
C2232 Gc_1.n27 VSS 0.0496f
C2233 Gc_1.t16 VSS 0.0229f
C2234 Gc_1.n28 VSS 0.0229f
C2235 Gc_1.n29 VSS 0.0491f
C2236 Gc_1.t22 VSS 0.0229f
C2237 Gc_1.n30 VSS 0.0229f
C2238 Gc_1.n31 VSS 0.0496f
C2239 Gc_1.n32 VSS 0.0551f
C2240 Gc_1.t143 VSS 0.0807f
C2241 Gc_1.n33 VSS 0.149f
C2242 Gc_1.t123 VSS 0.135f
C2243 Gc_1.n34 VSS 0.203f
C2244 Gc_1.t133 VSS 0.135f
C2245 Gc_1.n35 VSS 0.203f
C2246 Gc_1.t119 VSS 0.0807f
C2247 Gc_1.n36 VSS 0.149f
C2248 Gc_1.t129 VSS 0.0807f
C2249 Gc_1.n37 VSS 0.149f
C2250 Gc_1.t109 VSS 0.135f
C2251 Gc_1.n38 VSS 0.203f
C2252 Gc_1.t107 VSS 0.135f
C2253 Gc_1.n39 VSS 0.203f
C2254 Gc_1.t116 VSS 0.0807f
C2255 Gc_1.n40 VSS 0.149f
C2256 Gc_1.t135 VSS 0.0807f
C2257 Gc_1.n41 VSS 0.149f
C2258 Gc_1.t114 VSS 0.135f
C2259 Gc_1.n42 VSS 0.203f
C2260 Gc_1.t112 VSS 0.135f
C2261 Gc_1.n43 VSS 0.203f
C2262 Gc_1.t121 VSS 0.0807f
C2263 Gc_1.n44 VSS 0.149f
C2264 Gc_1.t134 VSS 0.0807f
C2265 Gc_1.n45 VSS 0.149f
C2266 Gc_1.t97 VSS 0.135f
C2267 Gc_1.n46 VSS 0.203f
C2268 Gc_1.t118 VSS 0.135f
C2269 Gc_1.n47 VSS 0.203f
C2270 Gc_1.t113 VSS 0.0807f
C2271 Gc_1.n48 VSS 0.23f
C2272 Gc_1.n49 VSS 0.0389f
C2273 Gc_1.t75 VSS 0.0229f
C2274 Gc_1.n50 VSS 0.0229f
C2275 Gc_1.n51 VSS 0.087f
C2276 Gc_1.t71 VSS 0.0229f
C2277 Gc_1.n52 VSS 0.0229f
C2278 Gc_1.n53 VSS 0.0861f
C2279 Gc_1.t79 VSS 0.0229f
C2280 Gc_1.n54 VSS 0.0229f
C2281 Gc_1.n55 VSS 0.0511f
C2282 Gc_1.t34 VSS 0.128f
C2283 Gc_1.n56 VSS 0.202f
C2284 Gc_1.t78 VSS 0.0814f
C2285 Gc_1.n57 VSS 0.144f
C2286 Gc_1.t38 VSS 0.0814f
C2287 Gc_1.t94 VSS 0.128f
C2288 Gc_1.n58 VSS 0.202f
C2289 Gc_1.n59 VSS 0.139f
C2290 Gc_1.n60 VSS 0.029f
C2291 Gc_1.n61 VSS 0.0507f
C2292 Gc_1.n62 VSS 0.0853f
C2293 Gc_1.t95 VSS 0.0229f
C2294 Gc_1.n63 VSS 0.0229f
C2295 Gc_1.n64 VSS 0.0866f
C2296 Gc_1.t83 VSS 0.0229f
C2297 Gc_1.n65 VSS 0.0229f
C2298 Gc_1.n66 VSS 0.0511f
C2299 Gc_1.t58 VSS 0.128f
C2300 Gc_1.n67 VSS 0.202f
C2301 Gc_1.t82 VSS 0.0814f
C2302 Gc_1.n68 VSS 0.141f
C2303 Gc_1.t36 VSS 0.0814f
C2304 Gc_1.t66 VSS 0.128f
C2305 Gc_1.n69 VSS 0.202f
C2306 Gc_1.n70 VSS 0.142f
C2307 Gc_1.n71 VSS 0.029f
C2308 Gc_1.n72 VSS 0.0522f
C2309 Gc_1.n73 VSS 0.0844f
C2310 Gc_1.t67 VSS 0.0229f
C2311 Gc_1.n74 VSS 0.0229f
C2312 Gc_1.n75 VSS 0.0852f
C2313 Gc_1.t73 VSS 0.0229f
C2314 Gc_1.n76 VSS 0.0229f
C2315 Gc_1.n77 VSS 0.051f
C2316 Gc_1.t54 VSS 0.128f
C2317 Gc_1.n78 VSS 0.202f
C2318 Gc_1.t72 VSS 0.0814f
C2319 Gc_1.n79 VSS 0.142f
C2320 Gc_1.t42 VSS 0.0814f
C2321 Gc_1.t64 VSS 0.128f
C2322 Gc_1.n80 VSS 0.202f
C2323 Gc_1.n81 VSS 0.14f
C2324 Gc_1.n82 VSS 0.029f
C2325 Gc_1.n83 VSS 0.0492f
C2326 Gc_1.n84 VSS 0.0861f
C2327 Gc_1.t65 VSS 0.0229f
C2328 Gc_1.n85 VSS 0.0229f
C2329 Gc_1.n86 VSS 0.0875f
C2330 Gc_1.t77 VSS 0.0229f
C2331 Gc_1.n87 VSS 0.0229f
C2332 Gc_1.n88 VSS 0.0511f
C2333 Gc_1.t48 VSS 0.128f
C2334 Gc_1.n89 VSS 0.202f
C2335 Gc_1.t76 VSS 0.0814f
C2336 Gc_1.n90 VSS 0.142f
C2337 Gc_1.t62 VSS 0.0814f
C2338 Gc_1.t92 VSS 0.128f
C2339 Gc_1.n91 VSS 0.202f
C2340 Gc_1.n92 VSS 0.141f
C2341 Gc_1.n93 VSS 0.029f
C2342 Gc_1.n94 VSS 0.0507f
C2343 Gc_1.n95 VSS 0.0853f
C2344 Gc_1.t93 VSS 0.0229f
C2345 Gc_1.n96 VSS 0.0229f
C2346 Gc_1.n97 VSS 0.0856f
C2347 Gc_1.t85 VSS 0.0229f
C2348 Gc_1.n98 VSS 0.0229f
C2349 Gc_1.n99 VSS 0.0889f
C2350 Gc_1.t91 VSS 0.0229f
C2351 Gc_1.n100 VSS 0.0229f
C2352 Gc_1.n101 VSS 0.051f
C2353 Gc_1.t44 VSS 0.128f
C2354 Gc_1.n102 VSS 0.202f
C2355 Gc_1.t90 VSS 0.0814f
C2356 Gc_1.n103 VSS 0.141f
C2357 Gc_1.t86 VSS 0.134f
C2358 Gc_1.t46 VSS 0.128f
C2359 Gc_1.n104 VSS 0.276f
C2360 Gc_1.t88 VSS 0.128f
C2361 Gc_1.n105 VSS 0.202f
C2362 Gc_1.t50 VSS 0.0814f
C2363 Gc_1.n106 VSS 0.142f
C2364 Gc_1.n107 VSS 0.029f
C2365 Gc_1.n108 VSS 0.0485f
C2366 Gc_1.n109 VSS 0.0865f
C2367 Gc_1.t89 VSS 0.0229f
C2368 Gc_1.n110 VSS 0.0229f
C2369 Gc_1.n111 VSS 0.0861f
C2370 Gc_1.n112 VSS 0.141f
C2371 Gc_1.n113 VSS 0.395f
C2372 Gc_1.n114 VSS 0.123f
C2373 Gc_1.n115 VSS 0.0219f
C2374 Gc_1.n116 VSS 0.118f
C2375 Gc_1.n117 VSS 0.368f
C2376 Gc_1.t69 VSS 0.0229f
C2377 Gc_1.n118 VSS 0.0229f
C2378 Gc_1.n119 VSS 0.0501f
C2379 Gc_1.n120 VSS 0.101f
C2380 Gc_1.t56 VSS 0.128f
C2381 Gc_1.n121 VSS 0.202f
C2382 Gc_1.t68 VSS 0.0814f
C2383 Gc_1.n122 VSS 0.144f
C2384 Gc_1.t52 VSS 0.0814f
C2385 Gc_1.t84 VSS 0.128f
C2386 Gc_1.n123 VSS 0.202f
C2387 Gc_1.n124 VSS 0.139f
C2388 Gc_1.n125 VSS 0.029f
C2389 Gc_1.n126 VSS 0.0398f
C2390 Gc_1.n127 VSS 0.133f
C2391 Gc_1.n128 VSS 0.0817f
C2392 Gc_1.n129 VSS 0.41f
C2393 Gc_1.n130 VSS 0.12f
C2394 Gc_1.n131 VSS 0.0219f
C2395 Gc_1.n132 VSS 0.118f
C2396 Gc_1.n133 VSS 0.363f
C2397 Gc_1.n134 VSS 0.121f
C2398 Gc_1.n135 VSS 0.0219f
C2399 Gc_1.n136 VSS 0.121f
C2400 Gc_1.n137 VSS 0.362f
C2401 Gc_1.n138 VSS 0.122f
C2402 Gc_1.n139 VSS 0.0219f
C2403 Gc_1.n140 VSS 0.119f
C2404 Gc_1.n141 VSS 0.359f
C2405 Gc_1.n142 VSS 0.119f
C2406 Gc_1.n143 VSS 0.0219f
C2407 Gc_1.n144 VSS 0.121f
C2408 Gc_1.n145 VSS 0.365f
C2409 Gc_1.t81 VSS 0.0229f
C2410 Gc_1.n146 VSS 0.0229f
C2411 Gc_1.n147 VSS 0.0499f
C2412 Gc_1.n148 VSS 0.0952f
C2413 Gc_1.t40 VSS 0.134f
C2414 Gc_1.t74 VSS 0.128f
C2415 Gc_1.n149 VSS 0.276f
C2416 Gc_1.t60 VSS 0.128f
C2417 Gc_1.n150 VSS 0.202f
C2418 Gc_1.t80 VSS 0.0814f
C2419 Gc_1.n151 VSS 0.146f
C2420 Gc_1.t32 VSS 0.0814f
C2421 Gc_1.t70 VSS 0.128f
C2422 Gc_1.n152 VSS 0.202f
C2423 Gc_1.n153 VSS 0.136f
C2424 Gc_1.n154 VSS 0.029f
C2425 Gc_1.n155 VSS 0.0403f
C2426 Gc_1.n156 VSS 0.132f
C2427 Gc_1.n157 VSS 0.0873f
C2428 Gc_1.n158 VSS 0.575f
C2429 Gc_1.n159 VSS 0.199f
C2430 Gc_1.n160 VSS 1.23f
C2431 Gc_1.n161 VSS 0.523f
C2432 Gc_1.n162 VSS 0.276f
C2433 Gc_1.n163 VSS 0.272f
C2434 Gc_1.n164 VSS 0.276f
C2435 Gc_1.n165 VSS 0.272f
C2436 Gc_1.n166 VSS 0.276f
C2437 Gc_1.n167 VSS 0.272f
C2438 Gc_1.n168 VSS 0.276f
C2439 Gc_1.n169 VSS 0.272f
C2440 Gc_1.n170 VSS 0.276f
C2441 Gc_1.n171 VSS 0.272f
C2442 Gc_1.n172 VSS 0.276f
C2443 Gc_1.n173 VSS 0.272f
C2444 Gc_1.n174 VSS 0.276f
C2445 Gc_1.n175 VSS 0.272f
C2446 Gc_1.n176 VSS 0.276f
C2447 Gc_1.n177 VSS 0.547f
C2448 Gc_1.t125 VSS 0.0807f
C2449 Gc_1.t139 VSS 0.135f
C2450 Gc_1.t141 VSS 0.135f
C2451 Gc_1.t142 VSS 0.0807f
C2452 Gc_1.t120 VSS 0.0807f
C2453 Gc_1.t136 VSS 0.135f
C2454 Gc_1.t138 VSS 0.135f
C2455 Gc_1.t132 VSS 0.0807f
C2456 Gc_1.t99 VSS 0.0807f
C2457 Gc_1.t108 VSS 0.135f
C2458 Gc_1.t96 VSS 0.135f
C2459 Gc_1.t124 VSS 0.0807f
C2460 Gc_1.t137 VSS 0.0807f
C2461 Gc_1.t127 VSS 0.135f
C2462 Gc_1.t104 VSS 0.135f
C2463 Gc_1.t110 VSS 0.0807f
C2464 Gc_1.n178 VSS 0.149f
C2465 Gc_1.n179 VSS 0.203f
C2466 Gc_1.n180 VSS 0.203f
C2467 Gc_1.n181 VSS 0.149f
C2468 Gc_1.n182 VSS 0.149f
C2469 Gc_1.n183 VSS 0.203f
C2470 Gc_1.n184 VSS 0.203f
C2471 Gc_1.n185 VSS 0.149f
C2472 Gc_1.n186 VSS 0.149f
C2473 Gc_1.n187 VSS 0.203f
C2474 Gc_1.n188 VSS 0.203f
C2475 Gc_1.n189 VSS 0.149f
C2476 Gc_1.n190 VSS 0.149f
C2477 Gc_1.n191 VSS 0.203f
C2478 Gc_1.n192 VSS 0.203f
C2479 Gc_1.n193 VSS 0.224f
C2480 Gc_1.n194 VSS 1.21f
C2481 Gc_1.n195 VSS 0.0562f
C2482 Gc_1.n196 VSS 0.021f
C2483 Gc_1.n197 VSS 0.00195f
C2484 Gc_1.n198 VSS 0.00225f
C2485 Gc_1.n199 VSS 0.0149f
C2486 OUT5.t34 VSS 0.00776f
C2487 OUT5.n0 VSS 0.00776f
C2488 OUT5.n1 VSS 0.0155f
C2489 OUT5.t19 VSS 0.00776f
C2490 OUT5.n2 VSS 0.00776f
C2491 OUT5.n3 VSS 0.0155f
C2492 OUT5.t20 VSS 0.00776f
C2493 OUT5.n4 VSS 0.00776f
C2494 OUT5.n5 VSS 0.0155f
C2495 OUT5.t42 VSS 0.00776f
C2496 OUT5.n6 VSS 0.00776f
C2497 OUT5.n7 VSS 0.0212f
C2498 OUT5.n8 VSS 0.0641f
C2499 OUT5.n9 VSS 0.0398f
C2500 OUT5.n10 VSS 0.0603f
C2501 OUT5.t26 VSS 0.00776f
C2502 OUT5.n11 VSS 0.00776f
C2503 OUT5.n12 VSS 0.0155f
C2504 OUT5.t38 VSS 0.00776f
C2505 OUT5.n13 VSS 0.00776f
C2506 OUT5.n14 VSS 0.0155f
C2507 OUT5.t36 VSS 0.00776f
C2508 OUT5.n15 VSS 0.00776f
C2509 OUT5.n16 VSS 0.0155f
C2510 OUT5.t28 VSS 0.00776f
C2511 OUT5.n17 VSS 0.00776f
C2512 OUT5.n18 VSS 0.0212f
C2513 OUT5.n19 VSS 0.0639f
C2514 OUT5.n20 VSS 0.0398f
C2515 OUT5.n21 VSS 0.0354f
C2516 OUT5.n22 VSS 0.0695f
C2517 OUT5.t47 VSS 0.00776f
C2518 OUT5.n23 VSS 0.00776f
C2519 OUT5.n24 VSS 0.0155f
C2520 OUT5.t25 VSS 0.00776f
C2521 OUT5.n25 VSS 0.00776f
C2522 OUT5.n26 VSS 0.0155f
C2523 OUT5.t31 VSS 0.00776f
C2524 OUT5.n27 VSS 0.00776f
C2525 OUT5.n28 VSS 0.0155f
C2526 OUT5.t39 VSS 0.00776f
C2527 OUT5.n29 VSS 0.00776f
C2528 OUT5.n30 VSS 0.0214f
C2529 OUT5.n31 VSS 0.0726f
C2530 OUT5.n32 VSS 0.0399f
C2531 OUT5.n33 VSS 0.0376f
C2532 OUT5.t22 VSS 0.00776f
C2533 OUT5.n34 VSS 0.00776f
C2534 OUT5.n35 VSS 0.0155f
C2535 OUT5.t35 VSS 0.00776f
C2536 OUT5.n36 VSS 0.00776f
C2537 OUT5.n37 VSS 0.0155f
C2538 OUT5.t32 VSS 0.00776f
C2539 OUT5.n38 VSS 0.00776f
C2540 OUT5.n39 VSS 0.0155f
C2541 OUT5.t2 VSS 0.00776f
C2542 OUT5.n40 VSS 0.00776f
C2543 OUT5.n41 VSS 0.0212f
C2544 OUT5.n42 VSS 0.0639f
C2545 OUT5.n43 VSS 0.0491f
C2546 OUT5.n44 VSS 0.0609f
C2547 OUT5.n45 VSS 0.0593f
C2548 OUT5.n46 VSS 0.856f
C2549 OUT5.n47 VSS 0.0185f
C2550 OUT5.t6 VSS 0.00776f
C2551 OUT5.n48 VSS 0.00776f
C2552 OUT5.n49 VSS 0.0169f
C2553 OUT5.t10 VSS 0.00776f
C2554 OUT5.n50 VSS 0.00776f
C2555 OUT5.n51 VSS 0.0164f
C2556 OUT5.t11 VSS 0.00776f
C2557 OUT5.n52 VSS 0.00776f
C2558 OUT5.n53 VSS 0.0169f
C2559 OUT5.t9 VSS 0.00776f
C2560 OUT5.n54 VSS 0.00776f
C2561 OUT5.n55 VSS 0.0175f
C2562 OUT5.n56 VSS 0.0247f
C2563 OUT5.n57 VSS 0.103f
C2564 OUT5.t12 VSS 0.00776f
C2565 OUT5.n58 VSS 0.00776f
C2566 OUT5.n59 VSS 0.0164f
C2567 OUT5.t8 VSS 0.00776f
C2568 OUT5.n60 VSS 0.00776f
C2569 OUT5.n61 VSS 0.0169f
C2570 OUT5.t7 VSS 0.0237f
C2571 OUT5.n62 VSS 0.205f
C2572 OUT5.n63 VSS 0.118f
C2573 OUT5.n64 VSS 0.272f
C2574 OUT5.t5 VSS 0.0186f
C2575 OUT5.n65 VSS 0.265f
C2576 OUT5.n66 VSS 0.121f
C2577 OUT5.n67 VSS 0.118f
C2578 OUT5.n68 VSS 0.122f
C2579 OUT5.n69 VSS 0.0949f
C2580 a_n2265_3941.t0 VSS 0.0419f
C2581 a_n2265_3941.t4 VSS 0.0419f
C2582 a_n2265_3941.n0 VSS 0.0419f
C2583 a_n2265_3941.n1 VSS 0.0935f
C2584 a_n2265_3941.t10 VSS 0.0419f
C2585 a_n2265_3941.n2 VSS 0.0419f
C2586 a_n2265_3941.n3 VSS 0.0948f
C2587 a_n2265_3941.t3 VSS 0.0419f
C2588 a_n2265_3941.n4 VSS 0.0419f
C2589 a_n2265_3941.n5 VSS 0.0935f
C2590 a_n2265_3941.t9 VSS 0.0419f
C2591 a_n2265_3941.n6 VSS 0.0419f
C2592 a_n2265_3941.n7 VSS 0.0948f
C2593 a_n2265_3941.t6 VSS 0.0419f
C2594 a_n2265_3941.n8 VSS 0.0419f
C2595 a_n2265_3941.n9 VSS 0.112f
C2596 a_n2265_3941.n10 VSS 0.309f
C2597 a_n2265_3941.n11 VSS 0.216f
C2598 a_n2265_3941.t45 VSS 0.0577f
C2599 a_n2265_3941.t16 VSS 0.0577f
C2600 a_n2265_3941.t27 VSS 0.0577f
C2601 a_n2265_3941.t29 VSS 0.0577f
C2602 a_n2265_3941.t41 VSS 0.0577f
C2603 a_n2265_3941.t43 VSS 0.0577f
C2604 a_n2265_3941.t39 VSS 0.0577f
C2605 a_n2265_3941.t51 VSS 0.0577f
C2606 a_n2265_3941.t12 VSS 0.0577f
C2607 a_n2265_3941.t24 VSS 0.0577f
C2608 a_n2265_3941.t25 VSS 0.0577f
C2609 a_n2265_3941.t38 VSS 0.0577f
C2610 a_n2265_3941.t33 VSS 0.0577f
C2611 a_n2265_3941.t36 VSS 0.0577f
C2612 a_n2265_3941.t47 VSS 0.0577f
C2613 a_n2265_3941.t50 VSS 0.0577f
C2614 a_n2265_3941.t21 VSS 0.0577f
C2615 a_n2265_3941.t31 VSS 0.0577f
C2616 a_n2265_3941.t35 VSS 0.0577f
C2617 a_n2265_3941.t46 VSS 0.0577f
C2618 a_n2265_3941.t49 VSS 0.0577f
C2619 a_n2265_3941.t20 VSS 0.0577f
C2620 a_n2265_3941.t30 VSS 0.0577f
C2621 a_n2265_3941.t32 VSS 0.0577f
C2622 a_n2265_3941.t14 VSS 0.0577f
C2623 a_n2265_3941.t19 VSS 0.0577f
C2624 a_n2265_3941.t48 VSS 0.0577f
C2625 a_n2265_3941.t37 VSS 0.0577f
C2626 a_n2265_3941.t34 VSS 0.0577f
C2627 a_n2265_3941.t23 VSS 0.0577f
C2628 a_n2265_3941.t22 VSS 0.0577f
C2629 a_n2265_3941.t13 VSS 0.0577f
C2630 a_n2265_3941.t42 VSS 0.0577f
C2631 a_n2265_3941.t40 VSS 0.0577f
C2632 a_n2265_3941.t28 VSS 0.0577f
C2633 a_n2265_3941.t26 VSS 0.0577f
C2634 a_n2265_3941.t15 VSS 0.0577f
C2635 a_n2265_3941.t18 VSS 0.0577f
C2636 a_n2265_3941.t17 VSS 0.0797f
C2637 a_n2265_3941.n12 VSS 0.0911f
C2638 a_n2265_3941.n13 VSS 0.0621f
C2639 a_n2265_3941.n14 VSS 0.0621f
C2640 a_n2265_3941.n15 VSS 0.0621f
C2641 a_n2265_3941.n16 VSS 0.0621f
C2642 a_n2265_3941.n17 VSS 0.0621f
C2643 a_n2265_3941.n18 VSS 0.0621f
C2644 a_n2265_3941.n19 VSS 0.0621f
C2645 a_n2265_3941.n20 VSS 0.0621f
C2646 a_n2265_3941.n21 VSS 0.0621f
C2647 a_n2265_3941.n22 VSS 0.0621f
C2648 a_n2265_3941.n23 VSS 0.0621f
C2649 a_n2265_3941.n24 VSS 0.0621f
C2650 a_n2265_3941.n25 VSS 0.0621f
C2651 a_n2265_3941.n26 VSS 0.0621f
C2652 a_n2265_3941.n27 VSS 0.0621f
C2653 a_n2265_3941.n28 VSS 0.0621f
C2654 a_n2265_3941.n29 VSS 0.0621f
C2655 a_n2265_3941.n30 VSS 0.0621f
C2656 a_n2265_3941.n31 VSS 0.0621f
C2657 a_n2265_3941.n32 VSS 0.0621f
C2658 a_n2265_3941.n33 VSS 0.0621f
C2659 a_n2265_3941.n34 VSS 0.0621f
C2660 a_n2265_3941.n35 VSS 0.0621f
C2661 a_n2265_3941.n36 VSS 0.0621f
C2662 a_n2265_3941.n37 VSS 0.0621f
C2663 a_n2265_3941.n38 VSS 0.0621f
C2664 a_n2265_3941.n39 VSS 0.0621f
C2665 a_n2265_3941.n40 VSS 0.0621f
C2666 a_n2265_3941.n41 VSS 0.0621f
C2667 a_n2265_3941.n42 VSS 0.0621f
C2668 a_n2265_3941.n43 VSS 0.0621f
C2669 a_n2265_3941.n44 VSS 0.0621f
C2670 a_n2265_3941.n45 VSS 0.0621f
C2671 a_n2265_3941.n46 VSS 0.0621f
C2672 a_n2265_3941.n47 VSS 0.0621f
C2673 a_n2265_3941.n48 VSS 0.0621f
C2674 a_n2265_3941.n49 VSS 0.0911f
C2675 a_n2265_3941.t44 VSS 0.143f
C2676 a_n2265_3941.n50 VSS 0.255f
C2677 a_n2265_3941.n51 VSS 0.0944f
C2678 a_n2265_3941.n52 VSS 0.0419f
C2679 b2.t3 VSS 0.0437f
C2680 b2.n0 VSS 0.0996f
C2681 b2.n1 VSS 0.00542f
C2682 b2.n2 VSS 0.0111f
C2683 b2.n3 VSS 0.00733f
C2684 b2.t6 VSS 0.0659f
C2685 b2.t4 VSS 0.0147f
C2686 b2.n4 VSS 0.0232f
C2687 b2.n5 VSS 0.00477f
C2688 b2.n6 VSS 0.0497f
C2689 b2.n7 VSS 0.0115f
C2690 b2.n8 VSS 0.115f
C2691 b2.t5 VSS 4.33e-19
C2692 b2.t2 VSS 0.0732f
C2693 b2.n9 VSS 0.143f
C2694 b2.n10 VSS 4.25f
C2695 b2.t1 VSS 0.015f
C2696 b2.t0 VSS 0.0119f
C2697 b2.n11 VSS 0.202f
C2698 b2.n12 VSS 3.18f
C2699 b6b.t49 VSS 0.18f
C2700 b6b.t29 VSS 0.0418f
C2701 b6b.n0 VSS 0.209f
C2702 b6b.t46 VSS 0.0418f
C2703 b6b.n1 VSS 0.181f
C2704 b6b.t28 VSS 0.0418f
C2705 b6b.n2 VSS 0.221f
C2706 b6b.n3 VSS 0.333f
C2707 b6b.n4 VSS 0.0159f
C2708 b6b.t20 VSS 0.0239f
C2709 b6b.t21 VSS 0.123f
C2710 b6b.t15 VSS 0.0319f
C2711 b6b.t45 VSS 0.0342f
C2712 b6b.n5 VSS 0.0687f
C2713 b6b.t30 VSS 0.0319f
C2714 b6b.n6 VSS 0.0687f
C2715 b6b.t11 VSS 0.0641f
C2716 b6b.n7 VSS 0.163f
C2717 b6b.t2 VSS 0.0419f
C2718 b6b.n8 VSS 0.0996f
C2719 b6b.n9 VSS 0.102f
C2720 b6b.t44 VSS 0.0319f
C2721 b6b.t27 VSS 0.0342f
C2722 b6b.n10 VSS 0.0693f
C2723 b6b.t26 VSS 0.0319f
C2724 b6b.n11 VSS 0.0693f
C2725 b6b.t9 VSS 0.0641f
C2726 b6b.n12 VSS 0.143f
C2727 b6b.t50 VSS 0.0407f
C2728 b6b.n13 VSS 0.124f
C2729 b6b.n14 VSS 0.0214f
C2730 b6b.n15 VSS 0.0155f
C2731 b6b.n16 VSS 0.0961f
C2732 b6b.t4 VSS 0.125f
C2733 b6b.t39 VSS 0.04f
C2734 b6b.n17 VSS 0.134f
C2735 b6b.t10 VSS 0.04f
C2736 b6b.n18 VSS 0.116f
C2737 b6b.t19 VSS 0.04f
C2738 b6b.n19 VSS 0.131f
C2739 b6b.n20 VSS 0.299f
C2740 b6b.t24 VSS 0.0671f
C2741 b6b.t25 VSS 0.16f
C2742 b6b.t23 VSS 0.0338f
C2743 b6b.t42 VSS 0.0332f
C2744 b6b.n21 VSS 0.0714f
C2745 b6b.t48 VSS 0.0338f
C2746 b6b.n22 VSS 0.0714f
C2747 b6b.t17 VSS 0.062f
C2748 b6b.n23 VSS 0.127f
C2749 b6b.t14 VSS 0.0658f
C2750 b6b.n24 VSS 0.0763f
C2751 b6b.t12 VSS 0.0385f
C2752 b6b.n25 VSS 0.0791f
C2753 b6b.t31 VSS 0.0385f
C2754 b6b.n26 VSS 0.0791f
C2755 b6b.t33 VSS 0.0658f
C2756 b6b.n27 VSS 0.0763f
C2757 b6b.t37 VSS 0.0334f
C2758 b6b.t7 VSS 0.0336f
C2759 b6b.n28 VSS 0.0706f
C2760 b6b.t18 VSS 0.0334f
C2761 b6b.n29 VSS 0.0706f
C2762 b6b.t36 VSS 0.0624f
C2763 b6b.n30 VSS 0.0998f
C2764 b6b.t38 VSS 0.0668f
C2765 b6b.t40 VSS 0.098f
C2766 b6b.n31 VSS 0.131f
C2767 b6b.n32 VSS 0.398f
C2768 b6b.n33 VSS 0.178f
C2769 b6b.n34 VSS 0.0109f
C2770 b6b.n35 VSS 0.0121f
C2771 b6b.n36 VSS 0.125f
C2772 b6b.t43 VSS 0.0249f
C2773 b6b.n37 VSS 0.156f
C2774 b6b.t47 VSS 0.103f
C2775 b6b.t41 VSS 0.0342f
C2776 b6b.t8 VSS 0.0329f
C2777 b6b.n38 VSS 0.0708f
C2778 b6b.t16 VSS 0.0342f
C2779 b6b.n39 VSS 0.0708f
C2780 b6b.t32 VSS 0.0609f
C2781 b6b.n40 VSS 0.111f
C2782 b6b.t34 VSS 0.0439f
C2783 b6b.n41 VSS 0.0709f
C2784 b6b.t5 VSS 0.0439f
C2785 b6b.n42 VSS 0.0709f
C2786 b6b.t6 VSS 0.0314f
C2787 b6b.t22 VSS 0.0357f
C2788 b6b.n43 VSS 0.0695f
C2789 b6b.t35 VSS 0.0314f
C2790 b6b.n44 VSS 0.0695f
C2791 b6b.t3 VSS 0.0637f
C2792 b6b.n45 VSS 0.0883f
C2793 b6b.t13 VSS 0.0439f
C2794 b6b.n46 VSS 0.114f
C2795 b6b.n47 VSS 0.0618f
C2796 b6b.n48 VSS 0.0113f
C2797 b6b.n49 VSS 0.148f
C2798 OUT6.t2 VSS 0.0157f
C2799 OUT6.n0 VSS 0.0157f
C2800 OUT6.n1 VSS 0.0484f
C2801 OUT6.t68 VSS 0.0157f
C2802 OUT6.n2 VSS 0.0157f
C2803 OUT6.n3 VSS 0.0314f
C2804 OUT6.t1 VSS 0.0157f
C2805 OUT6.n4 VSS 0.0157f
C2806 OUT6.n5 VSS 0.0314f
C2807 OUT6.t93 VSS 0.0157f
C2808 OUT6.n6 VSS 0.0157f
C2809 OUT6.n7 VSS 0.0314f
C2810 OUT6.t52 VSS 0.0157f
C2811 OUT6.n8 VSS 0.0157f
C2812 OUT6.n9 VSS 0.0314f
C2813 OUT6.t53 VSS 0.0157f
C2814 OUT6.n10 VSS 0.0157f
C2815 OUT6.n11 VSS 0.0314f
C2816 OUT6.t77 VSS 0.0157f
C2817 OUT6.n12 VSS 0.0157f
C2818 OUT6.n13 VSS 0.0401f
C2819 OUT6.t76 VSS 0.0157f
C2820 OUT6.n14 VSS 0.0157f
C2821 OUT6.n15 VSS 0.0314f
C2822 OUT6.n16 VSS 0.184f
C2823 OUT6.n17 VSS 0.131f
C2824 OUT6.n18 VSS 0.0731f
C2825 OUT6.t48 VSS 0.0157f
C2826 OUT6.n19 VSS 0.0157f
C2827 OUT6.n20 VSS 0.0391f
C2828 OUT6.t66 VSS 0.0157f
C2829 OUT6.n21 VSS 0.0157f
C2830 OUT6.n22 VSS 0.0314f
C2831 OUT6.n23 VSS 0.159f
C2832 OUT6.n24 VSS 0.119f
C2833 OUT6.n25 VSS 0.0526f
C2834 OUT6.n26 VSS 0.0888f
C2835 OUT6.n27 VSS 0.0668f
C2836 OUT6.n28 VSS 0.163f
C2837 OUT6.t7 VSS 0.0157f
C2838 OUT6.n29 VSS 0.0157f
C2839 OUT6.n30 VSS 0.0314f
C2840 OUT6.t44 VSS 0.0157f
C2841 OUT6.n31 VSS 0.0157f
C2842 OUT6.n32 VSS 0.0314f
C2843 OUT6.t63 VSS 0.0157f
C2844 OUT6.n33 VSS 0.0157f
C2845 OUT6.n34 VSS 0.0314f
C2846 OUT6.t84 VSS 0.0157f
C2847 OUT6.n35 VSS 0.0157f
C2848 OUT6.n36 VSS 0.0389f
C2849 OUT6.t5 VSS 0.0157f
C2850 OUT6.n37 VSS 0.0157f
C2851 OUT6.n38 VSS 0.0314f
C2852 OUT6.n39 VSS 0.155f
C2853 OUT6.t80 VSS 0.0157f
C2854 OUT6.n40 VSS 0.0157f
C2855 OUT6.n41 VSS 0.0314f
C2856 OUT6.t92 VSS 0.0157f
C2857 OUT6.n42 VSS 0.0157f
C2858 OUT6.n43 VSS 0.0342f
C2859 OUT6.t79 VSS 0.0157f
C2860 OUT6.n44 VSS 0.0157f
C2861 OUT6.n45 VSS 0.0314f
C2862 OUT6.t72 VSS 0.0157f
C2863 OUT6.n46 VSS 0.0157f
C2864 OUT6.n47 VSS 0.0314f
C2865 OUT6.t0 VSS 0.0157f
C2866 OUT6.n48 VSS 0.0157f
C2867 OUT6.n49 VSS 0.0575f
C2868 OUT6.n50 VSS 0.199f
C2869 OUT6.t67 VSS 0.0157f
C2870 OUT6.n51 VSS 0.0157f
C2871 OUT6.n52 VSS 0.0393f
C2872 OUT6.t57 VSS 0.0157f
C2873 OUT6.n53 VSS 0.0157f
C2874 OUT6.n54 VSS 0.0314f
C2875 OUT6.n55 VSS 0.163f
C2876 OUT6.n56 VSS 0.121f
C2877 OUT6.n57 VSS 0.0315f
C2878 OUT6.n58 VSS 0.101f
C2879 OUT6.t64 VSS 0.0157f
C2880 OUT6.n59 VSS 0.0157f
C2881 OUT6.n60 VSS 0.0341f
C2882 OUT6.t51 VSS 0.0157f
C2883 OUT6.n61 VSS 0.0157f
C2884 OUT6.n62 VSS 0.0314f
C2885 OUT6.t4 VSS 0.0157f
C2886 OUT6.n63 VSS 0.0157f
C2887 OUT6.n64 VSS 0.0392f
C2888 OUT6.t74 VSS 0.0157f
C2889 OUT6.n65 VSS 0.0157f
C2890 OUT6.n66 VSS 0.0314f
C2891 OUT6.n67 VSS 0.159f
C2892 OUT6.t3 VSS 0.0157f
C2893 OUT6.n68 VSS 0.0157f
C2894 OUT6.n69 VSS 0.0314f
C2895 OUT6.t47 VSS 0.0157f
C2896 OUT6.n70 VSS 0.0157f
C2897 OUT6.n71 VSS 0.0579f
C2898 OUT6.n72 VSS 0.197f
C2899 OUT6.n73 VSS 0.117f
C2900 OUT6.n74 VSS 0.0367f
C2901 OUT6.n75 VSS 0.0837f
C2902 OUT6.n76 VSS 0.306f
C2903 OUT6.t78 VSS 0.0157f
C2904 OUT6.n77 VSS 0.0157f
C2905 OUT6.n78 VSS 0.0314f
C2906 OUT6.t61 VSS 0.0157f
C2907 OUT6.n79 VSS 0.0157f
C2908 OUT6.n80 VSS 0.0402f
C2909 OUT6.t62 VSS 0.0157f
C2910 OUT6.n81 VSS 0.0157f
C2911 OUT6.n82 VSS 0.0314f
C2912 OUT6.n83 VSS 0.18f
C2913 OUT6.n84 VSS 0.11f
C2914 OUT6.n85 VSS 0.0919f
C2915 OUT6.n86 VSS 0.0543f
C2916 OUT6.n87 VSS 0.117f
C2917 OUT6.n88 VSS 0.0578f
C2918 OUT6.n89 VSS 0.0899f
C2919 OUT6.n90 VSS 0.0625f
C2920 OUT6.t43 VSS 0.0157f
C2921 OUT6.n91 VSS 0.0157f
C2922 OUT6.n92 VSS 0.0503f
C2923 OUT6.n93 VSS 0.186f
C2924 OUT6.n94 VSS 2.24f
C2925 OUT6.n95 VSS 0.0374f
C2926 OUT6.t10 VSS 0.0157f
C2927 OUT6.n96 VSS 0.0157f
C2928 OUT6.n97 VSS 0.0351f
C2929 OUT6.t22 VSS 0.0157f
C2930 OUT6.n98 VSS 0.0157f
C2931 OUT6.n99 VSS 0.0332f
C2932 OUT6.t24 VSS 0.0157f
C2933 OUT6.n100 VSS 0.0157f
C2934 OUT6.n101 VSS 0.0351f
C2935 OUT6.t38 VSS 0.0157f
C2936 OUT6.n102 VSS 0.0157f
C2937 OUT6.n103 VSS 0.0332f
C2938 OUT6.t36 VSS 0.0157f
C2939 OUT6.n104 VSS 0.0157f
C2940 OUT6.n105 VSS 0.0351f
C2941 OUT6.t35 VSS 0.0157f
C2942 OUT6.n106 VSS 0.0157f
C2943 OUT6.n107 VSS 0.0332f
C2944 OUT6.t20 VSS 0.0157f
C2945 OUT6.n108 VSS 0.0157f
C2946 OUT6.n109 VSS 0.0351f
C2947 OUT6.t19 VSS 0.0157f
C2948 OUT6.n110 VSS 0.0157f
C2949 OUT6.n111 VSS 0.0332f
C2950 OUT6.t34 VSS 0.0157f
C2951 OUT6.n112 VSS 0.0157f
C2952 OUT6.n113 VSS 0.0351f
C2953 OUT6.t30 VSS 0.0157f
C2954 OUT6.n114 VSS 0.0157f
C2955 OUT6.n115 VSS 0.0332f
C2956 OUT6.t18 VSS 0.0157f
C2957 OUT6.n116 VSS 0.0157f
C2958 OUT6.n117 VSS 0.0351f
C2959 OUT6.t40 VSS 0.0157f
C2960 OUT6.n118 VSS 0.0157f
C2961 OUT6.n119 VSS 0.0332f
C2962 OUT6.t27 VSS 0.0157f
C2963 OUT6.n120 VSS 0.0157f
C2964 OUT6.n121 VSS 0.0351f
C2965 OUT6.t26 VSS 0.0157f
C2966 OUT6.n122 VSS 0.0157f
C2967 OUT6.n123 VSS 0.0332f
C2968 OUT6.t16 VSS 0.0157f
C2969 OUT6.n124 VSS 0.0157f
C2970 OUT6.n125 VSS 0.0351f
C2971 OUT6.t15 VSS 0.0474f
C2972 OUT6.n126 VSS 0.381f
C2973 OUT6.n127 VSS 0.219f
C2974 OUT6.n128 VSS 0.234f
C2975 OUT6.n129 VSS 0.219f
C2976 OUT6.n130 VSS 0.234f
C2977 OUT6.n131 VSS 0.219f
C2978 OUT6.n132 VSS 0.234f
C2979 OUT6.n133 VSS 0.219f
C2980 OUT6.n134 VSS 0.234f
C2981 OUT6.n135 VSS 0.219f
C2982 OUT6.n136 VSS 0.234f
C2983 OUT6.n137 VSS 0.219f
C2984 OUT6.n138 VSS 0.234f
C2985 OUT6.n139 VSS 0.219f
C2986 OUT6.n140 VSS 0.234f
C2987 OUT6.n141 VSS 0.175f
C2988 IT.t36 VSS 0.0204f
C2989 IT.t74 VSS 0.0641f
C2990 IT.t106 VSS 0.0245f
C2991 IT.n0 VSS 0.0545f
C2992 IT.t82 VSS 0.0245f
C2993 IT.n1 VSS 0.0491f
C2994 IT.t37 VSS 0.0245f
C2995 IT.n2 VSS 0.0491f
C2996 IT.t65 VSS 0.0245f
C2997 IT.n3 VSS 0.0491f
C2998 IT.t97 VSS 0.0245f
C2999 IT.n4 VSS 0.0491f
C3000 IT.t53 VSS 0.0245f
C3001 IT.n5 VSS 0.0491f
C3002 IT.t94 VSS 0.0245f
C3003 IT.n6 VSS 0.0491f
C3004 IT.t64 VSS 0.0245f
C3005 IT.n7 VSS 0.0491f
C3006 IT.t28 VSS 0.0245f
C3007 IT.n8 VSS 0.0491f
C3008 IT.t80 VSS 0.0245f
C3009 IT.n9 VSS 0.0491f
C3010 IT.t52 VSS 0.0245f
C3011 IT.n10 VSS 0.0491f
C3012 IT.t77 VSS 0.0245f
C3013 IT.n11 VSS 0.0491f
C3014 IT.t48 VSS 0.0245f
C3015 IT.n12 VSS 0.0491f
C3016 IT.t86 VSS 0.0245f
C3017 IT.n13 VSS 0.0496f
C3018 IT.n14 VSS 0.0834f
C3019 IT.t96 VSS 0.017f
C3020 IT.n15 VSS 0.0136f
C3021 IT.t55 VSS 0.0392f
C3022 IT.t83 VSS 0.0224f
C3023 IT.n16 VSS 0.0571f
C3024 IT.t46 VSS 0.0224f
C3025 IT.n17 VSS 0.047f
C3026 IT.t95 VSS 0.0224f
C3027 IT.n18 VSS 0.047f
C3028 IT.t56 VSS 0.0224f
C3029 IT.n19 VSS 0.047f
C3030 IT.t84 VSS 0.0224f
C3031 IT.n20 VSS 0.047f
C3032 IT.t104 VSS 0.0224f
C3033 IT.n21 VSS 0.047f
C3034 IT.t75 VSS 0.0224f
C3035 IT.n22 VSS 0.047f
C3036 IT.t107 VSS 0.0224f
C3037 IT.n23 VSS 0.047f
C3038 IT.t32 VSS 0.0224f
C3039 IT.n24 VSS 0.047f
C3040 IT.t39 VSS 0.0224f
C3041 IT.n25 VSS 0.047f
C3042 IT.t87 VSS 0.0224f
C3043 IT.n26 VSS 0.047f
C3044 IT.t57 VSS 0.0224f
C3045 IT.n27 VSS 0.047f
C3046 IT.t85 VSS 0.0224f
C3047 IT.n28 VSS 0.047f
C3048 IT.t49 VSS 0.0224f
C3049 IT.n29 VSS 0.0476f
C3050 IT.n30 VSS 0.0115f
C3051 IT.n31 VSS 0.00919f
C3052 IT.n32 VSS 0.00676f
C3053 IT.n33 VSS 0.00823f
C3054 IT.n34 VSS 0.109f
C3055 IT.n35 VSS 1.56f
C3056 IT.t44 VSS 0.0639f
C3057 IT.t68 VSS 0.0244f
C3058 IT.n36 VSS 0.0543f
C3059 IT.t26 VSS 0.0244f
C3060 IT.n37 VSS 0.049f
C3061 IT.t27 VSS 0.0244f
C3062 IT.n38 VSS 0.049f
C3063 IT.t40 VSS 0.0244f
C3064 IT.n39 VSS 0.049f
C3065 IT.t33 VSS 0.0244f
C3066 IT.n40 VSS 0.049f
C3067 IT.t93 VSS 0.0244f
C3068 IT.n41 VSS 0.049f
C3069 IT.t78 VSS 0.0244f
C3070 IT.n42 VSS 0.049f
C3071 IT.t38 VSS 0.0244f
C3072 IT.n43 VSS 0.049f
C3073 IT.t41 VSS 0.0244f
C3074 IT.n44 VSS 0.049f
C3075 IT.t100 VSS 0.0244f
C3076 IT.n45 VSS 0.049f
C3077 IT.t25 VSS 0.0244f
C3078 IT.n46 VSS 0.049f
C3079 IT.t67 VSS 0.0244f
C3080 IT.n47 VSS 0.049f
C3081 IT.t50 VSS 0.0244f
C3082 IT.n48 VSS 0.049f
C3083 IT.t30 VSS 0.0244f
C3084 IT.n49 VSS 0.0493f
C3085 IT.n50 VSS 0.0271f
C3086 IT.n51 VSS 0.00889f
C3087 IT.t90 VSS 0.0174f
C3088 IT.n52 VSS 0.0174f
C3089 IT.n53 VSS 0.00701f
C3090 IT.n54 VSS 0.0399f
C3091 IT.n55 VSS 0.00925f
C3092 IT.t69 VSS 0.0192f
C3093 IT.n56 VSS 0.0164f
C3094 IT.t88 VSS 0.0244f
C3095 IT.t81 VSS 0.0244f
C3096 IT.t45 VSS 0.0244f
C3097 IT.t59 VSS 0.0244f
C3098 IT.t79 VSS 0.0244f
C3099 IT.t98 VSS 0.0244f
C3100 IT.t34 VSS 0.0244f
C3101 IT.t35 VSS 0.0244f
C3102 IT.t76 VSS 0.0244f
C3103 IT.t91 VSS 0.0244f
C3104 IT.t31 VSS 0.0244f
C3105 IT.n57 VSS 0.049f
C3106 IT.n58 VSS 0.049f
C3107 IT.n59 VSS 0.049f
C3108 IT.n60 VSS 0.049f
C3109 IT.n61 VSS 0.049f
C3110 IT.n62 VSS 0.049f
C3111 IT.n63 VSS 0.049f
C3112 IT.n64 VSS 0.049f
C3113 IT.n65 VSS 0.049f
C3114 IT.n66 VSS 0.049f
C3115 IT.n67 VSS 0.049f
C3116 IT.n68 VSS 0.0111f
C3117 IT.n69 VSS 0.00656f
C3118 IT.n70 VSS 0.0084f
C3119 IT.n71 VSS 0.221f
C3120 IT.n72 VSS 1.97f
C3121 IT.t58 VSS 0.0238f
C3122 IT.t54 VSS 0.0238f
C3123 IT.n73 VSS 0.0484f
C3124 IT.n74 VSS 0.0487f
C3125 IT.t63 VSS 0.0231f
C3126 IT.n75 VSS 0.0386f
C3127 IT.t6 VSS 0.015f
C3128 IT.t24 VSS 0.0244f
C3129 IT.n76 VSS 0.049f
C3130 IT.t66 VSS 0.0244f
C3131 IT.n77 VSS 0.049f
C3132 IT.t42 VSS 0.0244f
C3133 IT.n78 VSS 0.0495f
C3134 IT.n79 VSS 0.0107f
C3135 IT.t102 VSS 0.0192f
C3136 IT.n80 VSS 0.0163f
C3137 IT.n81 VSS 0.00903f
C3138 IT.n82 VSS 0.00655f
C3139 IT.n83 VSS 0.12f
C3140 IT.t103 VSS 0.02f
C3141 IT.n84 VSS 0.146f
C3142 IT.t47 VSS 0.024f
C3143 IT.n85 VSS 0.049f
C3144 IT.t62 VSS 0.024f
C3145 IT.n86 VSS 0.0485f
C3146 IT.t101 VSS 0.024f
C3147 IT.n87 VSS 0.0514f
C3148 IT.n88 VSS 0.0326f
C3149 IT.n89 VSS 0.0498f
C3150 IT.n90 VSS 0.0514f
C3151 IT.t12 VSS 0.0222f
C3152 IT.n91 VSS 0.0526f
C3153 IT.t13 VSS 0.00679f
C3154 IT.n92 VSS 0.00679f
C3155 IT.n93 VSS 0.037f
C3156 IT.n94 VSS 0.0294f
C3157 IT.t4 VSS 0.0222f
C3158 IT.n95 VSS 0.0513f
C3159 IT.t2 VSS 0.0217f
C3160 IT.n96 VSS 0.0479f
C3161 IT.n97 VSS 0.00307f
C3162 IT.n98 VSS 0.00287f
C3163 IT.t105 VSS 0.024f
C3164 IT.n99 VSS 0.0517f
C3165 IT.n100 VSS 0.0133f
C3166 IT.t3 VSS 0.0171f
C3167 IT.n101 VSS 0.0296f
C3168 IT.n102 VSS 0.0228f
C3169 IT.n103 VSS 5.75e-19
C3170 IT.n104 VSS 0.00673f
C3171 IT.n105 VSS 0.199f
C3172 IT.t11 VSS 0.00679f
C3173 IT.n106 VSS 0.00679f
C3174 IT.n107 VSS 0.0145f
C3175 IT.t10 VSS 0.0219f
C3176 IT.t73 VSS 0.0411f
C3177 IT.t60 VSS 0.0238f
C3178 IT.n108 VSS 0.0596f
C3179 IT.t43 VSS 0.0238f
C3180 IT.n109 VSS 0.0484f
C3181 IT.t61 VSS 0.0238f
C3182 IT.n110 VSS 0.0538f
C3183 IT.n111 VSS 0.0569f
C3184 IT.t8 VSS 0.0219f
C3185 IT.n112 VSS 0.0515f
C3186 IT.n113 VSS 0.0107f
C3187 IT.n114 VSS 0.101f
C3188 IT.n115 VSS 0.513f
C3189 IT.t51 VSS 0.0238f
C3190 IT.n116 VSS 0.054f
C3191 IT.t0 VSS 0.0223f
C3192 IT.n117 VSS 0.056f
C3193 IT.t14 VSS 0.0223f
C3194 IT.n118 VSS 0.0506f
C3195 IT.n119 VSS 0.00937f
C3196 IT.n120 VSS 0.0142f
C3197 IT.t15 VSS 0.00679f
C3198 IT.n121 VSS 0.00679f
C3199 IT.n122 VSS 0.0147f
C3200 IT.n123 VSS 0.025f
C3201 IT.n124 VSS 0.00866f
C3202 IT.n125 VSS 0.133f
C3203 IT.n126 VSS 0.507f
C3204 IT.n127 VSS 0.312f
C3205 IT.t17 VSS 0.00679f
C3206 IT.n128 VSS 0.00679f
C3207 IT.n129 VSS 0.0145f
C3208 IT.t18 VSS 0.00679f
C3209 IT.n130 VSS 0.00679f
C3210 IT.n131 VSS 0.0145f
C3211 IT.t19 VSS 0.00679f
C3212 IT.n132 VSS 0.00679f
C3213 IT.n133 VSS 0.0365f
C3214 IT.t20 VSS 0.00679f
C3215 IT.n134 VSS 0.00679f
C3216 IT.n135 VSS 0.0145f
C3217 IT.n136 VSS 0.403f
C3218 IT.n137 VSS 0.58f
C3219 IT.n138 VSS 0.662f
C3220 IT.n139 VSS 1.37f
C3221 IT.n140 VSS 0.161f
C3222 IT.n141 VSS 0.0173f
C3223 IT.n142 VSS 0.0101f
C3224 IT.t89 VSS 0.024f
C3225 IT.t29 VSS 0.024f
C3226 IT.n143 VSS 0.0485f
C3227 IT.n144 VSS 0.0486f
C3228 IT.t70 VSS 0.0233f
C3229 IT.n145 VSS 0.0486f
C3230 IT.n146 VSS 0.00294f
C3231 IT.n147 VSS 3.57e-19
C3232 b6.t38 VSS 0.0391f
C3233 b6.t18 VSS 0.0583f
C3234 b6.t37 VSS 0.136f
C3235 b6.t28 VSS 0.04f
C3236 b6.n0 VSS 0.113f
C3237 b6.t41 VSS 0.04f
C3238 b6.n1 VSS 0.0863f
C3239 b6.t45 VSS 0.0583f
C3240 b6.t16 VSS 0.0878f
C3241 b6.n2 VSS 0.0874f
C3242 b6.t17 VSS 0.0583f
C3243 b6.t36 VSS 0.0878f
C3244 b6.n3 VSS 0.088f
C3245 b6.n4 VSS 0.081f
C3246 b6.t9 VSS 0.0391f
C3247 b6.t43 VSS 0.0583f
C3248 b6.t14 VSS 0.137f
C3249 b6.n5 VSS 0.11f
C3250 b6.n6 VSS 0.0655f
C3251 b6.t2 VSS 0.0668f
C3252 b6.t15 VSS 0.0413f
C3253 b6.n7 VSS 0.23f
C3254 b6.t12 VSS 0.0413f
C3255 b6.n8 VSS 0.181f
C3256 b6.t32 VSS 0.0546f
C3257 b6.n9 VSS 0.0701f
C3258 b6.n10 VSS 0.566f
C3259 b6.t25 VSS 0.0592f
C3260 b6.t6 VSS 0.116f
C3261 b6.t49 VSS 0.0404f
C3262 b6.n11 VSS 0.112f
C3263 b6.t27 VSS 0.0404f
C3264 b6.n12 VSS 0.0751f
C3265 b6.t48 VSS 0.0625f
C3266 b6.n13 VSS 0.0767f
C3267 b6.t20 VSS 0.0326f
C3268 b6.n14 VSS 0.0694f
C3269 b6.t47 VSS 0.0326f
C3270 b6.n15 VSS 0.0694f
C3271 b6.t30 VSS 0.0625f
C3272 b6.n16 VSS 0.0767f
C3273 b6.t8 VSS 0.0404f
C3274 b6.n17 VSS 0.0751f
C3275 b6.t35 VSS 0.0404f
C3276 b6.n18 VSS 0.0751f
C3277 b6.t11 VSS 0.0592f
C3278 b6.t40 VSS 0.0892f
C3279 b6.n19 VSS 0.107f
C3280 b6.n20 VSS 0.53f
C3281 b6.n21 VSS 0.175f
C3282 b6.t42 VSS 0.0676f
C3283 b6.t23 VSS 0.0415f
C3284 b6.n22 VSS 0.17f
C3285 b6.t4 VSS 0.0415f
C3286 b6.n23 VSS 0.133f
C3287 b6.t29 VSS 0.0415f
C3288 b6.n24 VSS 0.136f
C3289 b6.t44 VSS 0.0383f
C3290 b6.n25 VSS 0.0935f
C3291 b6.n26 VSS 0.00126f
C3292 b6.t1 VSS 0.0125f
C3293 b6.t0 VSS 0.00523f
C3294 b6.n27 VSS 0.203f
C3295 b6.n28 VSS 0.201f
C3296 b6.n29 VSS 0.0122f
C3297 b6.n30 VSS 0.532f
C3298 b6.n31 VSS 0.673f
C3299 b6.n32 VSS 0.0166f
C3300 b6.t39 VSS 0.059f
C3301 b6.t24 VSS 0.149f
C3302 b6.t22 VSS 0.036f
C3303 b6.t21 VSS 0.0348f
C3304 b6.n33 VSS 0.0778f
C3305 b6.t3 VSS 0.036f
C3306 b6.n34 VSS 0.0778f
C3307 b6.t50 VSS 0.063f
C3308 b6.n35 VSS 0.124f
C3309 b6.t19 VSS 0.0639f
C3310 b6.n36 VSS 0.0743f
C3311 b6.t34 VSS 0.0317f
C3312 b6.n37 VSS 0.0671f
C3313 b6.t13 VSS 0.0317f
C3314 b6.n38 VSS 0.0671f
C3315 b6.t46 VSS 0.0639f
C3316 b6.n39 VSS 0.0743f
C3317 b6.t7 VSS 0.0351f
C3318 b6.t5 VSS 0.0357f
C3319 b6.n40 VSS 0.076f
C3320 b6.t33 VSS 0.0351f
C3321 b6.n41 VSS 0.076f
C3322 b6.t31 VSS 0.0639f
C3323 b6.n42 VSS 0.0971f
C3324 b6.t26 VSS 0.0592f
C3325 b6.t10 VSS 0.0898f
C3326 b6.n43 VSS 0.125f
C3327 b6.n44 VSS 0.0708f
C3328 b6.n46 VSS 0.139f
C3329 SD3_1.t31 VSS 0.00898f
C3330 SD3_1.n0 VSS 0.00898f
C3331 SD3_1.n1 VSS 0.0372f
C3332 SD3_1.t8 VSS 0.00898f
C3333 SD3_1.n2 VSS 0.00898f
C3334 SD3_1.n3 VSS 0.0342f
C3335 SD3_1.t17 VSS 0.00898f
C3336 SD3_1.n4 VSS 0.00898f
C3337 SD3_1.n5 VSS 0.0371f
C3338 SD3_1.t54 VSS 0.00898f
C3339 SD3_1.n6 VSS 0.00898f
C3340 SD3_1.n7 VSS 0.0343f
C3341 SD3_1.t36 VSS 0.00898f
C3342 SD3_1.n8 VSS 0.00898f
C3343 SD3_1.n9 VSS 0.018f
C3344 SD3_1.n10 VSS 0.0222f
C3345 SD3_1.n11 VSS 0.00975f
C3346 SD3_1.t37 VSS 0.0083f
C3347 SD3_1.n12 VSS 0.0363f
C3348 SD3_1.t48 VSS 0.00898f
C3349 SD3_1.n13 VSS 0.00898f
C3350 SD3_1.n14 VSS 0.018f
C3351 SD3_1.n15 VSS 0.0161f
C3352 SD3_1.t63 VSS 0.00898f
C3353 SD3_1.n16 VSS 0.00898f
C3354 SD3_1.n17 VSS 0.0372f
C3355 SD3_1.t18 VSS 0.00898f
C3356 SD3_1.n18 VSS 0.00898f
C3357 SD3_1.n19 VSS 0.018f
C3358 SD3_1.n20 VSS 0.0161f
C3359 SD3_1.t28 VSS 0.00898f
C3360 SD3_1.n21 VSS 0.00898f
C3361 SD3_1.n22 VSS 0.0342f
C3362 SD3_1.t60 VSS 0.00898f
C3363 SD3_1.n23 VSS 0.00898f
C3364 SD3_1.n24 VSS 0.018f
C3365 SD3_1.n25 VSS 0.0222f
C3366 SD3_1.t59 VSS 0.00898f
C3367 SD3_1.n26 VSS 0.00898f
C3368 SD3_1.n27 VSS 0.0342f
C3369 SD3_1.t10 VSS 0.00898f
C3370 SD3_1.n28 VSS 0.00898f
C3371 SD3_1.n29 VSS 0.018f
C3372 SD3_1.n30 VSS 0.0222f
C3373 SD3_1.t38 VSS 0.00898f
C3374 SD3_1.n31 VSS 0.00898f
C3375 SD3_1.n32 VSS 0.034f
C3376 SD3_1.t62 VSS 0.00898f
C3377 SD3_1.n33 VSS 0.00898f
C3378 SD3_1.n34 VSS 0.018f
C3379 SD3_1.n35 VSS 0.0161f
C3380 SD3_1.t61 VSS 0.00898f
C3381 SD3_1.n36 VSS 0.00898f
C3382 SD3_1.n37 VSS 0.0377f
C3383 SD3_1.t19 VSS 0.00898f
C3384 SD3_1.n38 VSS 0.00898f
C3385 SD3_1.n39 VSS 0.0181f
C3386 SD3_1.n40 VSS 0.0229f
C3387 SD3_1.t26 VSS 0.00898f
C3388 SD3_1.n41 VSS 0.00898f
C3389 SD3_1.n42 VSS 0.0375f
C3390 SD3_1.t44 VSS 0.00898f
C3391 SD3_1.n43 VSS 0.00898f
C3392 SD3_1.n44 VSS 0.0373f
C3393 SD3_1.t14 VSS 0.00898f
C3394 SD3_1.n45 VSS 0.00898f
C3395 SD3_1.n46 VSS 0.018f
C3396 SD3_1.n47 VSS 0.0222f
C3397 SD3_1.t34 VSS 0.00898f
C3398 SD3_1.n48 VSS 0.00898f
C3399 SD3_1.n49 VSS 0.034f
C3400 SD3_1.t2 VSS 0.00898f
C3401 SD3_1.n50 VSS 0.00898f
C3402 SD3_1.n51 VSS 0.0374f
C3403 SD3_1.t3 VSS 0.00898f
C3404 SD3_1.n52 VSS 0.00898f
C3405 SD3_1.n53 VSS 0.0251f
C3406 SD3_1.t23 VSS 0.00898f
C3407 SD3_1.n54 VSS 0.00898f
C3408 SD3_1.n55 VSS 0.0343f
C3409 SD3_1.n56 VSS 0.125f
C3410 SD3_1.n57 VSS 0.0341f
C3411 SD3_1.n58 VSS 0.0788f
C3412 SD3_1.t9 VSS 0.00898f
C3413 SD3_1.n59 VSS 0.00898f
C3414 SD3_1.n60 VSS 0.018f
C3415 SD3_1.n61 VSS 0.0161f
C3416 SD3_1.n62 VSS 0.0333f
C3417 SD3_1.n63 VSS 0.0332f
C3418 SD3_1.n64 VSS 0.0762f
C3419 SD3_1.t46 VSS 0.00898f
C3420 SD3_1.n65 VSS 0.00898f
C3421 SD3_1.n66 VSS 0.018f
C3422 SD3_1.n67 VSS 0.0161f
C3423 SD3_1.n68 VSS 0.0338f
C3424 SD3_1.n69 VSS 0.0336f
C3425 SD3_1.n70 VSS 0.0792f
C3426 SD3_1.n71 VSS 0.0337f
C3427 SD3_1.t0 VSS 0.00898f
C3428 SD3_1.n72 VSS 0.00898f
C3429 SD3_1.n73 VSS 0.0181f
C3430 SD3_1.n74 VSS 0.0229f
C3431 SD3_1.n75 VSS 0.0339f
C3432 SD3_1.n76 VSS 0.0792f
C3433 SD3_1.n77 VSS 0.0333f
C3434 SD3_1.n78 VSS 0.0335f
C3435 SD3_1.n79 VSS 0.0793f
C3436 SD3_1.n80 VSS 0.0337f
C3437 SD3_1.n81 VSS 0.034f
C3438 SD3_1.n82 VSS 0.0758f
C3439 SD3_1.n83 VSS 0.0332f
C3440 SD3_1.n84 VSS 0.0338f
C3441 SD3_1.n85 VSS 0.0765f
C3442 SD3_1.n86 VSS 0.0333f
C3443 SD3_1.n87 VSS 0.0343f
C3444 SD3_1.n88 VSS 0.0762f
C3445 SD3_1.n89 VSS 0.033f
C3446 SD3_1.n90 VSS 0.033f
C3447 SD3_1.n91 VSS 0.079f
C3448 SD3_1.n92 VSS 0.034f
C3449 SD3_1.n93 VSS 0.0337f
C3450 SD3_1.n94 VSS 0.0733f
C3451 SD3_1.n95 VSS 0.0335f
C3452 SD3_1.n96 VSS 0.0332f
C3453 SD3_1.n97 VSS 0.0764f
C3454 SD3_1.n98 VSS 0.0342f
C3455 SD3_1.n99 VSS 0.0346f
C3456 SD3_1.n100 VSS 0.0761f
C3457 SD3_1.n101 VSS 0.00975f
C3458 SD3_1.t51 VSS 0.0083f
C3459 SD3_1.n102 VSS 0.0179f
C3460 SD3_1.n103 VSS 0.0161f
C3461 SD3_1.n104 VSS 0.0341f
C3462 SD3_1.t21 VSS 0.00898f
C3463 SD3_1.n105 VSS 0.00898f
C3464 SD3_1.n106 VSS 0.018f
C3465 SD3_1.n107 VSS 0.0161f
C3466 SD3_1.n108 VSS 0.0354f
C3467 SD3_1.n109 VSS 0.0739f
C3468 SD3_1.n110 VSS 0.0336f
C3469 SD3_1.t55 VSS 0.00898f
C3470 SD3_1.n111 VSS 0.00898f
C3471 SD3_1.n112 VSS 0.018f
C3472 SD3_1.n113 VSS 0.00381f
C3473 SD3_1.n114 VSS 0.0166f
C3474 SD3_1.n115 VSS 0.0329f
C3475 SD3_1.t53 VSS 0.00898f
C3476 SD3_1.n116 VSS 0.00898f
C3477 SD3_1.n117 VSS 0.0375f
C3478 SD3_1.t30 VSS 0.00898f
C3479 SD3_1.n118 VSS 0.00898f
C3480 SD3_1.n119 VSS 0.0251f
C3481 SD3_1.n120 VSS 0.126f
C3482 SD3_1.n121 VSS 0.034f
C3483 SDn_2.t16 VSS 0.00619f
C3484 SDn_2.n0 VSS 0.00619f
C3485 SDn_2.n1 VSS 0.0182f
C3486 SDn_2.n2 VSS 0.00607f
C3487 SDn_2.t66 VSS 0.038f
C3488 SDn_2.t89 VSS 0.0232f
C3489 SDn_2.n3 VSS 0.0416f
C3490 SDn_2.t106 VSS 0.0232f
C3491 SDn_2.n4 VSS 0.031f
C3492 SDn_2.t92 VSS 0.0222f
C3493 SDn_2.n5 VSS 0.03f
C3494 SDn_2.t46 VSS 0.0222f
C3495 SDn_2.n6 VSS 0.03f
C3496 SDn_2.t49 VSS 0.0232f
C3497 SDn_2.n7 VSS 0.031f
C3498 SDn_2.t95 VSS 0.0232f
C3499 SDn_2.n8 VSS 0.031f
C3500 SDn_2.t47 VSS 0.0222f
C3501 SDn_2.n9 VSS 0.03f
C3502 SDn_2.t62 VSS 0.0222f
C3503 SDn_2.n10 VSS 0.03f
C3504 SDn_2.t97 VSS 0.0232f
C3505 SDn_2.n11 VSS 0.031f
C3506 SDn_2.t76 VSS 0.0232f
C3507 SDn_2.n12 VSS 0.031f
C3508 SDn_2.t55 VSS 0.0222f
C3509 SDn_2.n13 VSS 0.03f
C3510 SDn_2.t29 VSS 0.0222f
C3511 SDn_2.n14 VSS 0.03f
C3512 SDn_2.t61 VSS 0.0232f
C3513 SDn_2.n15 VSS 0.031f
C3514 SDn_2.t104 VSS 0.0232f
C3515 SDn_2.n16 VSS 0.031f
C3516 SDn_2.t98 VSS 0.0222f
C3517 SDn_2.n17 VSS 0.03f
C3518 SDn_2.t57 VSS 0.0222f
C3519 SDn_2.n18 VSS 0.03f
C3520 SDn_2.t103 VSS 0.0232f
C3521 SDn_2.n19 VSS 0.031f
C3522 SDn_2.t85 VSS 0.0232f
C3523 SDn_2.n20 VSS 0.031f
C3524 SDn_2.t64 VSS 0.0222f
C3525 SDn_2.n21 VSS 0.03f
C3526 SDn_2.t34 VSS 0.0222f
C3527 SDn_2.n22 VSS 0.03f
C3528 SDn_2.t65 VSS 0.0232f
C3529 SDn_2.n23 VSS 0.031f
C3530 SDn_2.t36 VSS 0.0232f
C3531 SDn_2.n24 VSS 0.031f
C3532 SDn_2.t42 VSS 0.0222f
C3533 SDn_2.n25 VSS 0.03f
C3534 SDn_2.t86 VSS 0.0222f
C3535 SDn_2.n26 VSS 0.03f
C3536 SDn_2.t24 VSS 0.0232f
C3537 SDn_2.n27 VSS 0.031f
C3538 SDn_2.t71 VSS 0.0232f
C3539 SDn_2.n28 VSS 0.031f
C3540 SDn_2.t67 VSS 0.0222f
C3541 SDn_2.n29 VSS 0.03f
C3542 SDn_2.t52 VSS 0.0222f
C3543 SDn_2.n30 VSS 0.03f
C3544 SDn_2.t74 VSS 0.0232f
C3545 SDn_2.n31 VSS 0.031f
C3546 SDn_2.t54 VSS 0.0232f
C3547 SDn_2.n32 VSS 0.031f
C3548 SDn_2.t25 VSS 0.0222f
C3549 SDn_2.n33 VSS 0.0402f
C3550 SDn_2.t87 VSS 0.0356f
C3551 SDn_2.t40 VSS 0.0213f
C3552 SDn_2.n34 VSS 0.0383f
C3553 SDn_2.t77 VSS 0.0213f
C3554 SDn_2.n35 VSS 0.0292f
C3555 SDn_2.t31 VSS 0.0203f
C3556 SDn_2.n36 VSS 0.0282f
C3557 SDn_2.t100 VSS 0.0203f
C3558 SDn_2.n37 VSS 0.0282f
C3559 SDn_2.t30 VSS 0.0213f
C3560 SDn_2.n38 VSS 0.0292f
C3561 SDn_2.t90 VSS 0.0213f
C3562 SDn_2.n39 VSS 0.0292f
C3563 SDn_2.t44 VSS 0.0203f
C3564 SDn_2.n40 VSS 0.0282f
C3565 SDn_2.t81 VSS 0.0203f
C3566 SDn_2.n41 VSS 0.0282f
C3567 SDn_2.t43 VSS 0.0213f
C3568 SDn_2.n42 VSS 0.0292f
C3569 SDn_2.t78 VSS 0.0213f
C3570 SDn_2.n43 VSS 0.0292f
C3571 SDn_2.t26 VSS 0.0203f
C3572 SDn_2.n44 VSS 0.0282f
C3573 SDn_2.t63 VSS 0.0203f
C3574 SDn_2.n45 VSS 0.0282f
C3575 SDn_2.t99 VSS 0.0213f
C3576 SDn_2.n46 VSS 0.0292f
C3577 SDn_2.t70 VSS 0.0213f
C3578 SDn_2.n47 VSS 0.0292f
C3579 SDn_2.t107 VSS 0.0203f
C3580 SDn_2.n48 VSS 0.0282f
C3581 SDn_2.t80 VSS 0.0203f
C3582 SDn_2.n49 VSS 0.0282f
C3583 SDn_2.t101 VSS 0.0213f
C3584 SDn_2.n50 VSS 0.0292f
C3585 SDn_2.t105 VSS 0.0213f
C3586 SDn_2.n51 VSS 0.0292f
C3587 SDn_2.t35 VSS 0.0203f
C3588 SDn_2.n52 VSS 0.0282f
C3589 SDn_2.t96 VSS 0.0203f
C3590 SDn_2.n53 VSS 0.0282f
C3591 SDn_2.t27 VSS 0.0213f
C3592 SDn_2.n54 VSS 0.0292f
C3593 SDn_2.t82 VSS 0.0213f
C3594 SDn_2.n55 VSS 0.0292f
C3595 SDn_2.t60 VSS 0.0203f
C3596 SDn_2.n56 VSS 0.0282f
C3597 SDn_2.t93 VSS 0.0203f
C3598 SDn_2.n57 VSS 0.0282f
C3599 SDn_2.t45 VSS 0.0213f
C3600 SDn_2.n58 VSS 0.0292f
C3601 SDn_2.t79 VSS 0.0213f
C3602 SDn_2.n59 VSS 0.0292f
C3603 SDn_2.t59 VSS 0.0203f
C3604 SDn_2.n60 VSS 0.0282f
C3605 SDn_2.t102 VSS 0.0203f
C3606 SDn_2.n61 VSS 0.0282f
C3607 SDn_2.t32 VSS 0.0213f
C3608 SDn_2.n62 VSS 0.0292f
C3609 SDn_2.t91 VSS 0.0213f
C3610 SDn_2.n63 VSS 0.0292f
C3611 SDn_2.t41 VSS 0.0203f
C3612 SDn_2.n64 VSS 0.036f
C3613 SDn_2.n65 VSS 1.68f
C3614 SDn_2.t75 VSS 0.0207f
C3615 SDn_2.n66 VSS 0.0409f
C3616 SDn_2.t94 VSS 0.0227f
C3617 SDn_2.n67 VSS 0.0305f
C3618 SDn_2.t51 VSS 0.0227f
C3619 SDn_2.n68 VSS 0.0305f
C3620 SDn_2.t48 VSS 0.0207f
C3621 SDn_2.n69 VSS 0.0286f
C3622 SDn_2.t37 VSS 0.0207f
C3623 SDn_2.n70 VSS 0.0286f
C3624 SDn_2.t39 VSS 0.0227f
C3625 SDn_2.n71 VSS 0.0305f
C3626 SDn_2.t68 VSS 0.0227f
C3627 SDn_2.n72 VSS 0.0305f
C3628 SDn_2.t33 VSS 0.0207f
C3629 SDn_2.n73 VSS 0.0334f
C3630 SDn_2.t14 VSS 0.0207f
C3631 SDn_2.n74 VSS 0.0334f
C3632 SDn_2.t0 VSS 0.0208f
C3633 SDn_2.n75 VSS 0.0284f
C3634 SDn_2.t10 VSS 0.0227f
C3635 SDn_2.n76 VSS 0.0305f
C3636 SDn_2.n77 VSS 0.0139f
C3637 SDn_2.t8 VSS 0.018f
C3638 SDn_2.n79 VSS 0.0153f
C3639 SDn_2.n80 VSS 0.0084f
C3640 SDn_2.n81 VSS 0.00836f
C3641 SDn_2.n82 VSS 0.063f
C3642 SDn_2.t1 VSS 0.00588f
C3643 SDn_2.n83 VSS 0.00655f
C3644 SDn_2.n84 VSS 0.0258f
C3645 SDn_2.t3 VSS 0.00572f
C3646 SDn_2.n85 VSS 0.00673f
C3647 SDn_2.n86 VSS 0.0205f
C3648 SDn_2.n87 VSS 0.00667f
C3649 SDn_2.t7 VSS 0.00577f
C3650 SDn_2.n88 VSS 0.0236f
C3651 SDn_2.n89 VSS 0.00667f
C3652 SDn_2.t19 VSS 0.00577f
C3653 SDn_2.n90 VSS 0.0178f
C3654 SDn_2.n91 VSS 0.0738f
C3655 SDn_2.n92 VSS 0.00667f
C3656 SDn_2.t20 VSS 0.00577f
C3657 SDn_2.n93 VSS 0.0197f
C3658 SDn_2.t84 VSS 0.0361f
C3659 SDn_2.t69 VSS 0.0227f
C3660 SDn_2.n94 VSS 0.04f
C3661 SDn_2.t88 VSS 0.0227f
C3662 SDn_2.n95 VSS 0.0305f
C3663 SDn_2.t58 VSS 0.0207f
C3664 SDn_2.n96 VSS 0.0286f
C3665 SDn_2.t50 VSS 0.0207f
C3666 SDn_2.n97 VSS 0.0286f
C3667 SDn_2.t72 VSS 0.0227f
C3668 SDn_2.n98 VSS 0.0305f
C3669 SDn_2.t38 VSS 0.0227f
C3670 SDn_2.n99 VSS 0.0305f
C3671 SDn_2.t73 VSS 0.0207f
C3672 SDn_2.n100 VSS 0.0332f
C3673 SDn_2.t6 VSS 0.0208f
C3674 SDn_2.n101 VSS 0.033f
C3675 SDn_2.t12 VSS 0.0227f
C3676 SDn_2.n102 VSS 0.0305f
C3677 SDn_2.t4 VSS 0.0208f
C3678 SDn_2.n103 VSS 0.0284f
C3679 SDn_2.n104 VSS 0.014f
C3680 SDn_2.t2 VSS 0.018f
C3681 SDn_2.n106 VSS 0.0153f
C3682 SDn_2.n107 VSS 0.00823f
C3683 SDn_2.n108 VSS 0.00607f
C3684 SDn_2.n109 VSS 0.00857f
C3685 SDn_2.n110 VSS 0.0624f
C3686 SDn_2.n111 VSS 0.029f
C3687 SDn_2.n112 VSS 0.0291f
C3688 SDn_2.n113 VSS 0.00673f
C3689 SDn_2.t18 VSS 0.00572f
C3690 SDn_2.n114 VSS 0.0123f
C3691 SDn_2.n115 VSS 0.00915f
C3692 SDn_2.n116 VSS 0.0248f
C3693 SDn_2.n117 VSS 0.0461f
C3694 SDn_2.n118 VSS 0.0219f
C3695 SDn_2.n119 VSS 0.022f
C3696 SDn_2.n120 VSS 0.00621f
C3697 SDn_2.t9 VSS 0.00619f
C3698 SDn_2.n121 VSS 0.00619f
C3699 SDn_2.n122 VSS 0.0124f
C3700 SDn_2.n123 VSS 0.00553f
C3701 SDn_2.n124 VSS 0.00998f
C3702 SDn_2.n125 VSS 4.98e-19
C3703 TG_1.IN.n0 VSS 0.296f
C3704 TG_1.IN.t38 VSS 0.0263f
C3705 TG_1.IN.t97 VSS 0.0263f
C3706 TG_1.IN.n1 VSS 0.0217f
C3707 TG_1.IN.t100 VSS 0.0267f
C3708 TG_1.IN.n2 VSS 0.0214f
C3709 TG_1.IN.t2 VSS 0.0157f
C3710 TG_1.IN.n3 VSS 0.0157f
C3711 TG_1.IN.n4 VSS 0.0315f
C3712 TG_1.IN.t262 VSS 0.0157f
C3713 TG_1.IN.n5 VSS 0.0157f
C3714 TG_1.IN.n6 VSS 0.0316f
C3715 TG_1.IN.t260 VSS 0.03f
C3716 TG_1.IN.t118 VSS 0.0337f
C3717 TG_1.IN.n7 VSS 0.133f
C3718 TG_1.IN.t261 VSS 0.0268f
C3719 TG_1.IN.t257 VSS 0.0273f
C3720 TG_1.IN.n8 VSS 0.0207f
C3721 TG_1.IN.n9 VSS 0.118f
C3722 TG_1.IN.n10 VSS 0.132f
C3723 TG_1.IN.t77 VSS 0.0194f
C3724 TG_1.IN.t31 VSS 0.0295f
C3725 TG_1.IN.n11 VSS 0.063f
C3726 TG_1.IN.n12 VSS 0.0302f
C3727 TG_1.IN.t78 VSS 0.0267f
C3728 TG_1.IN.t258 VSS 0.0269f
C3729 TG_1.IN.n13 VSS 0.0216f
C3730 TG_1.IN.n14 VSS 0.0446f
C3731 TG_1.IN.n15 VSS 0.0434f
C3732 TG_1.IN.t32 VSS 0.0271f
C3733 TG_1.IN.t117 VSS 0.027f
C3734 TG_1.IN.n16 VSS 0.0207f
C3735 TG_1.IN.n17 VSS 0.127f
C3736 TG_1.IN.t255 VSS 0.0157f
C3737 TG_1.IN.n18 VSS 0.0157f
C3738 TG_1.IN.n19 VSS 0.0385f
C3739 TG_1.IN.t106 VSS 0.0157f
C3740 TG_1.IN.n20 VSS 0.0157f
C3741 TG_1.IN.n21 VSS 0.0315f
C3742 TG_1.IN.n22 VSS 0.14f
C3743 TG_1.IN.t41 VSS 0.0711f
C3744 TG_1.IN.n23 VSS 0.203f
C3745 TG_1.IN.t42 VSS 0.0558f
C3746 TG_1.IN.n24 VSS 0.0157f
C3747 TG_1.IN.n25 VSS 0.0315f
C3748 TG_1.IN.n26 VSS 0.163f
C3749 TG_1.IN.n27 VSS 0.377f
C3750 TG_1.IN.t12 VSS 0.053f
C3751 TG_1.IN.n28 VSS 0.0157f
C3752 TG_1.IN.n29 VSS 0.0315f
C3753 TG_1.IN.n30 VSS 0.0699f
C3754 TG_1.IN.t11 VSS 0.0874f
C3755 TG_1.IN.n31 VSS 0.168f
C3756 TG_1.IN.n32 VSS 0.0594f
C3757 TG_1.IN.t59 VSS 0.0738f
C3758 TG_1.IN.n33 VSS 0.19f
C3759 TG_1.IN.t45 VSS 0.0633f
C3760 TG_1.IN.n34 VSS 0.186f
C3761 TG_1.IN.t245 VSS 0.0157f
C3762 TG_1.IN.t46 VSS 0.055f
C3763 TG_1.IN.n35 VSS 0.0315f
C3764 TG_1.IN.n36 VSS 0.224f
C3765 TG_1.IN.t107 VSS 0.0157f
C3766 TG_1.IN.t60 VSS 0.0551f
C3767 TG_1.IN.n37 VSS 0.0315f
C3768 TG_1.IN.n38 VSS 0.256f
C3769 TG_1.IN.n39 VSS 0.0524f
C3770 TG_1.IN.n40 VSS 0.155f
C3771 TG_1.IN.n41 VSS 0.159f
C3772 TG_1.IN.t102 VSS 0.0531f
C3773 TG_1.IN.t109 VSS 0.0531f
C3774 TG_1.IN.n42 VSS 0.0336f
C3775 TG_1.IN.t123 VSS 0.0531f
C3776 TG_1.IN.t133 VSS 0.0531f
C3777 TG_1.IN.n43 VSS 0.0315f
C3778 TG_1.IN.t66 VSS 0.0542f
C3779 TG_1.IN.n44 VSS 0.0157f
C3780 TG_1.IN.n45 VSS 0.034f
C3781 TG_1.IN.t36 VSS 0.0536f
C3782 TG_1.IN.t88 VSS 0.0555f
C3783 TG_1.IN.n46 VSS 0.0339f
C3784 TG_1.IN.t87 VSS 0.0668f
C3785 TG_1.IN.n47 VSS 0.17f
C3786 TG_1.IN.n48 VSS 0.0832f
C3787 TG_1.IN.t35 VSS 0.0668f
C3788 TG_1.IN.n49 VSS 0.0821f
C3789 TG_1.IN.n50 VSS 0.1f
C3790 TG_1.IN.n51 VSS 0.112f
C3791 TG_1.IN.t65 VSS 0.0679f
C3792 TG_1.IN.n52 VSS 0.0794f
C3793 TG_1.IN.n53 VSS 0.0847f
C3794 TG_1.IN.t253 VSS 0.0157f
C3795 TG_1.IN.n54 VSS 0.0157f
C3796 TG_1.IN.n55 VSS 0.0315f
C3797 TG_1.IN.t252 VSS 0.0157f
C3798 TG_1.IN.n56 VSS 0.0157f
C3799 TG_1.IN.n57 VSS 0.0315f
C3800 TG_1.IN.t249 VSS 0.0157f
C3801 TG_1.IN.n58 VSS 0.0157f
C3802 TG_1.IN.n59 VSS 0.0315f
C3803 TG_1.IN.t24 VSS 0.0532f
C3804 TG_1.IN.n60 VSS 0.0157f
C3805 TG_1.IN.n61 VSS 0.0315f
C3806 TG_1.IN.t248 VSS 0.0157f
C3807 TG_1.IN.t44 VSS 0.0556f
C3808 TG_1.IN.n62 VSS 0.0338f
C3809 TG_1.IN.t43 VSS 0.0696f
C3810 TG_1.IN.n63 VSS 0.178f
C3811 TG_1.IN.n64 VSS 0.301f
C3812 TG_1.IN.t76 VSS 0.0532f
C3813 TG_1.IN.t50 VSS 0.0552f
C3814 TG_1.IN.n65 VSS 0.0334f
C3815 TG_1.IN.t49 VSS 0.0629f
C3816 TG_1.IN.n66 VSS 0.171f
C3817 TG_1.IN.n67 VSS 0.079f
C3818 TG_1.IN.t75 VSS 0.0627f
C3819 TG_1.IN.n68 VSS 0.0825f
C3820 TG_1.IN.n69 VSS 0.101f
C3821 TG_1.IN.n70 VSS 0.101f
C3822 TG_1.IN.t23 VSS 0.0627f
C3823 TG_1.IN.n71 VSS 0.0819f
C3824 TG_1.IN.n72 VSS 0.267f
C3825 TG_1.IN.n73 VSS 0.0883f
C3826 TG_1.IN.t95 VSS 0.0157f
C3827 TG_1.IN.n74 VSS 0.0157f
C3828 TG_1.IN.n75 VSS 0.078f
C3829 TG_1.IN.n76 VSS 0.344f
C3830 TG_1.IN.n77 VSS 0.0891f
C3831 TG_1.IN.n78 VSS 0.0933f
C3832 TG_1.IN.t98 VSS 0.0157f
C3833 TG_1.IN.n79 VSS 0.0157f
C3834 TG_1.IN.n80 VSS 0.0322f
C3835 TG_1.IN.t251 VSS 0.0157f
C3836 TG_1.IN.n81 VSS 0.0157f
C3837 TG_1.IN.n82 VSS 0.0338f
C3838 TG_1.IN.n83 VSS 0.145f
C3839 TG_1.IN.n84 VSS 0.304f
C3840 TG_1.IN.n85 VSS 0.135f
C3841 TG_1.IN.t250 VSS 0.0157f
C3842 TG_1.IN.t80 VSS 0.0562f
C3843 TG_1.IN.n86 VSS 0.0345f
C3844 TG_1.IN.t79 VSS 0.072f
C3845 TG_1.IN.n87 VSS 0.182f
C3846 TG_1.IN.n88 VSS 0.149f
C3847 TG_1.IN.t104 VSS 0.053f
C3848 TG_1.IN.t137 VSS 0.053f
C3849 TG_1.IN.n89 VSS 0.0331f
C3850 TG_1.IN.n90 VSS 0.166f
C3851 TG_1.IN.n91 VSS 0.17f
C3852 TG_1.IN.n92 VSS 0.119f
C3853 TG_1.IN.t136 VSS 0.0531f
C3854 TG_1.IN.t247 VSS 0.0532f
C3855 TG_1.IN.n93 VSS 0.0315f
C3856 TG_1.IN.n94 VSS 0.0479f
C3857 TG_1.IN.n95 VSS 0.145f
C3858 TG_1.IN.n96 VSS 0.168f
C3859 TG_1.IN.n97 VSS 0.13f
C3860 TG_1.IN.n98 VSS 0.0434f
C3861 TG_1.IN.n99 VSS 0.605f
C3862 TG_1.IN.n100 VSS 0.602f
C3863 TG_1.IN.n101 VSS 0.242f
C3864 TG_1.IN.t142 VSS 0.0516f
C3865 TG_1.IN.n102 VSS 0.0324f
C3866 TG_1.IN.t140 VSS 0.0516f
C3867 TG_1.IN.t131 VSS 0.0516f
C3868 TG_1.IN.t231 VSS 0.0157f
C3869 TG_1.IN.n103 VSS 0.0157f
C3870 TG_1.IN.n104 VSS 0.0359f
C3871 TG_1.IN.t40 VSS 0.053f
C3872 TG_1.IN.n105 VSS 0.0157f
C3873 TG_1.IN.n106 VSS 0.0331f
C3874 TG_1.IN.t90 VSS 0.0601f
C3875 TG_1.IN.t64 VSS 0.0575f
C3876 TG_1.IN.n107 VSS 0.0404f
C3877 TG_1.IN.t63 VSS 0.088f
C3878 TG_1.IN.t89 VSS 0.0436f
C3879 TG_1.IN.n108 VSS 0.105f
C3880 TG_1.IN.n109 VSS 0.206f
C3881 TG_1.IN.n110 VSS 0.0982f
C3882 TG_1.IN.n111 VSS 0.0972f
C3883 TG_1.IN.t39 VSS 0.0599f
C3884 TG_1.IN.n112 VSS 0.0758f
C3885 TG_1.IN.n113 VSS 0.112f
C3886 TG_1.IN.t120 VSS 0.0157f
C3887 TG_1.IN.n114 VSS 0.0157f
C3888 TG_1.IN.n115 VSS 0.0339f
C3889 TG_1.IN.t234 VSS 0.0157f
C3890 TG_1.IN.n116 VSS 0.0157f
C3891 TG_1.IN.n117 VSS 0.0346f
C3892 TG_1.IN.n118 VSS 0.109f
C3893 TG_1.IN.t54 VSS 0.0539f
C3894 TG_1.IN.n119 VSS 0.154f
C3895 TG_1.IN.t19 VSS 0.0466f
C3896 TG_1.IN.t29 VSS 0.0519f
C3897 TG_1.IN.n120 VSS 0.0825f
C3898 TG_1.IN.n121 VSS 0.0285f
C3899 TG_1.IN.t20 VSS 0.0533f
C3900 TG_1.IN.n122 VSS 0.0342f
C3901 TG_1.IN.n123 VSS 0.0664f
C3902 TG_1.IN.t30 VSS 0.0535f
C3903 TG_1.IN.n124 VSS 0.0345f
C3904 TG_1.IN.n125 VSS 0.0697f
C3905 TG_1.IN.t53 VSS 0.0477f
C3906 TG_1.IN.t57 VSS 0.0509f
C3907 TG_1.IN.n126 VSS 0.0825f
C3908 TG_1.IN.n127 VSS 0.0264f
C3909 TG_1.IN.t58 VSS 0.0541f
C3910 TG_1.IN.n128 VSS 0.0871f
C3911 TG_1.IN.n129 VSS 0.0899f
C3912 TG_1.IN.n130 VSS 0.164f
C3913 TG_1.IN.t81 VSS 0.0472f
C3914 TG_1.IN.t85 VSS 0.0514f
C3915 TG_1.IN.n131 VSS 0.0825f
C3916 TG_1.IN.n132 VSS 0.0288f
C3917 TG_1.IN.t82 VSS 0.0532f
C3918 TG_1.IN.n133 VSS 0.0157f
C3919 TG_1.IN.n134 VSS 0.0341f
C3920 TG_1.IN.n135 VSS 0.0682f
C3921 TG_1.IN.t86 VSS 0.0535f
C3922 TG_1.IN.n136 VSS 0.0157f
C3923 TG_1.IN.n137 VSS 0.0315f
C3924 TG_1.IN.t240 VSS 0.0157f
C3925 TG_1.IN.n138 VSS 0.0157f
C3926 TG_1.IN.n139 VSS 0.0404f
C3927 TG_1.IN.t10 VSS 0.0157f
C3928 TG_1.IN.n140 VSS 0.0157f
C3929 TG_1.IN.n141 VSS 0.0315f
C3930 TG_1.IN.n142 VSS 0.12f
C3931 TG_1.IN.t232 VSS 0.0157f
C3932 TG_1.IN.t62 VSS 0.0533f
C3933 TG_1.IN.n143 VSS 0.0334f
C3934 TG_1.IN.t61 VSS 0.0482f
C3935 TG_1.IN.t67 VSS 0.0505f
C3936 TG_1.IN.n144 VSS 0.0817f
C3937 TG_1.IN.n145 VSS 0.157f
C3938 TG_1.IN.n146 VSS 0.0377f
C3939 TG_1.IN.n147 VSS 0.0912f
C3940 TG_1.IN.t230 VSS 0.0157f
C3941 TG_1.IN.t68 VSS 0.0534f
C3942 TG_1.IN.n148 VSS 0.0315f
C3943 TG_1.IN.n149 VSS 0.0993f
C3944 TG_1.IN.t227 VSS 0.0157f
C3945 TG_1.IN.n150 VSS 0.0157f
C3946 TG_1.IN.n151 VSS 0.0315f
C3947 TG_1.IN.t93 VSS 0.0157f
C3948 TG_1.IN.n152 VSS 0.0157f
C3949 TG_1.IN.n153 VSS 0.0391f
C3950 TG_1.IN.n154 VSS 0.108f
C3951 TG_1.IN.n155 VSS 0.157f
C3952 TG_1.IN.n156 VSS 0.128f
C3953 TG_1.IN.t233 VSS 0.0157f
C3954 TG_1.IN.n157 VSS 0.0157f
C3955 TG_1.IN.n158 VSS 0.0315f
C3956 TG_1.IN.t48 VSS 0.0535f
C3957 TG_1.IN.n159 VSS 0.0157f
C3958 TG_1.IN.n160 VSS 0.036f
C3959 TG_1.IN.t15 VSS 0.0877f
C3960 TG_1.IN.t69 VSS 0.0424f
C3961 TG_1.IN.n161 VSS 0.0986f
C3962 TG_1.IN.n162 VSS 0.119f
C3963 TG_1.IN.t47 VSS 0.0793f
C3964 TG_1.IN.n163 VSS 0.151f
C3965 TG_1.IN.n164 VSS 0.113f
C3966 TG_1.IN.n165 VSS 0.0681f
C3967 TG_1.IN.t70 VSS 0.0546f
C3968 TG_1.IN.t16 VSS 0.0529f
C3969 TG_1.IN.n166 VSS 0.0315f
C3970 TG_1.IN.n167 VSS 0.134f
C3971 TG_1.IN.n168 VSS 0.247f
C3972 TG_1.IN.t226 VSS 0.0157f
C3973 TG_1.IN.n169 VSS 0.0157f
C3974 TG_1.IN.n170 VSS 0.0359f
C3975 TG_1.IN.t239 VSS 0.0157f
C3976 TG_1.IN.t26 VSS 0.0546f
C3977 TG_1.IN.n171 VSS 0.0329f
C3978 TG_1.IN.t25 VSS 0.0598f
C3979 TG_1.IN.n172 VSS 0.166f
C3980 TG_1.IN.n173 VSS 0.184f
C3981 TG_1.IN.n174 VSS 0.225f
C3982 TG_1.IN.n175 VSS 0.307f
C3983 TG_1.IN.t8 VSS 0.0157f
C3984 TG_1.IN.n176 VSS 0.0157f
C3985 TG_1.IN.n177 VSS 0.0337f
C3986 TG_1.IN.n178 VSS 0.248f
C3987 TG_1.IN.n179 VSS 0.0384f
C3988 TG_1.IN.n180 VSS 0.158f
C3989 TG_1.IN.n181 VSS 0.104f
C3990 TG_1.IN.n182 VSS 0.0764f
C3991 TG_1.IN.t243 VSS 0.0157f
C3992 TG_1.IN.n183 VSS 0.0157f
C3993 TG_1.IN.n184 VSS 0.0341f
C3994 TG_1.IN.t228 VSS 0.0157f
C3995 TG_1.IN.n185 VSS 0.0157f
C3996 TG_1.IN.n186 VSS 0.0334f
C3997 TG_1.IN.n187 VSS 0.18f
C3998 TG_1.IN.n188 VSS 0.48f
C3999 TG_1.IN.n189 VSS 0.262f
C4000 TG_1.IN.n190 VSS 0.176f
C4001 TG_1.IN.n191 VSS 0.194f
C4002 TG_1.IN.t244 VSS 0.0157f
C4003 TG_1.IN.t14 VSS 0.0523f
C4004 TG_1.IN.n192 VSS 0.0315f
C4005 TG_1.IN.t13 VSS 0.0782f
C4006 TG_1.IN.n193 VSS 0.183f
C4007 TG_1.IN.n194 VSS 0.106f
C4008 TG_1.IN.n195 VSS 0.213f
C4009 TG_1.IN.n196 VSS 0.155f
C4010 TG_1.IN.t139 VSS 0.0516f
C4011 TG_1.IN.n197 VSS 0.0328f
C4012 TG_1.IN.n198 VSS 0.0954f
C4013 TG_1.IN.t126 VSS 0.0525f
C4014 TG_1.IN.n199 VSS 0.12f
C4015 TG_1.IN.n200 VSS 0.0824f
C4016 TG_1.IN.t130 VSS 0.0516f
C4017 TG_1.IN.n201 VSS 0.0337f
C4018 TG_1.IN.t238 VSS 0.0516f
C4019 TG_1.IN.n202 VSS 0.0331f
C4020 TG_1.IN.t129 VSS 0.0532f
C4021 TG_1.IN.n203 VSS 0.0325f
C4022 TG_1.IN.t141 VSS 0.0534f
C4023 TG_1.IN.t72 VSS 0.0528f
C4024 TG_1.IN.n204 VSS 0.0328f
C4025 TG_1.IN.t18 VSS 0.0533f
C4026 TG_1.IN.n205 VSS 0.0335f
C4027 TG_1.IN.n206 VSS 0.143f
C4028 TG_1.IN.t71 VSS 0.0393f
C4029 TG_1.IN.t17 VSS 0.0499f
C4030 TG_1.IN.n207 VSS 0.0731f
C4031 TG_1.IN.n208 VSS 0.0388f
C4032 TG_1.IN.n209 VSS 0.121f
C4033 TG_1.IN.t132 VSS 0.0535f
C4034 TG_1.IN.n210 VSS 0.224f
C4035 TG_1.IN.n211 VSS 0.09f
C4036 TG_1.IN.t236 VSS 0.0516f
C4037 TG_1.IN.n212 VSS 0.123f
C4038 TG_1.IN.n213 VSS 0.0969f
C4039 TG_1.IN.t235 VSS 0.0766f
C4040 TG_1.IN.t128 VSS 0.0583f
C4041 TG_1.IN.n214 VSS 0.156f
C4042 TG_1.IN.n215 VSS 0.242f
C4043 TG_1.IN.n216 VSS 0.061f
C4044 TG_1.IN.n217 VSS 0.135f
C4045 TG_1.IN.n218 VSS 0.0613f
C4046 TG_1.IN.n219 VSS 0.0968f
C4047 TG_1.IN.n220 VSS 0.12f
C4048 TG_1.IN.n221 VSS 0.0922f
C4049 TG_1.IN.t125 VSS 0.0525f
C4050 TG_1.IN.n222 VSS 0.092f
C4051 TG_1.IN.t127 VSS 0.053f
C4052 TG_1.IN.t237 VSS 0.053f
C4053 TG_1.IN.n223 VSS 0.131f
C4054 TG_1.IN.t22 VSS 0.0531f
C4055 TG_1.IN.n224 VSS 0.0332f
C4056 TG_1.IN.t56 VSS 0.0532f
C4057 TG_1.IN.n225 VSS 0.0333f
C4058 TG_1.IN.t21 VSS 0.0444f
C4059 TG_1.IN.t55 VSS 0.0449f
C4060 TG_1.IN.n226 VSS 0.0731f
C4061 TG_1.IN.n227 VSS 0.142f
C4062 TG_1.IN.n228 VSS 0.0346f
C4063 TG_1.IN.n229 VSS 0.12f
C4064 TG_1.IN.n230 VSS 0.0826f
C4065 TG_1.IN.n231 VSS 0.39f
C4066 TG_1.IN.n232 VSS 0.374f
C4067 TG_1.IN.t256 VSS 0.0432f
C4068 TG_1.IN.t259 VSS 0.0383f
C4069 TG_1.IN.n233 VSS 0.221f
C4070 TG_1.IN.n234 VSS 0.131f
C4071 TG_1.IN.n235 VSS 0.152f
C4072 TG_1.IN.n236 VSS 0.0792f
C4073 TG_1.IN.n237 VSS 0.0272f
C4074 TG_1.IN.n238 VSS 0.104f
C4075 TG_1.IN.n239 VSS 0.508f
C4076 TG_1.IN.n240 VSS 0.175f
C4077 TG_1.IN.n241 VSS 0.118f
C4078 TG_1.IN.n242 VSS 0.115f
C4079 TG_1.IN.n243 VSS 0.0948f
C4080 TG_1.IN.t99 VSS 0.0359f
C4081 TG_1.IN.t101 VSS 0.0363f
C4082 TG_1.IN.n244 VSS 0.119f
C4083 TG_1.IN.n245 VSS 0.124f
C4084 TG_1.IN.n246 VSS 0.189f
C4085 TG_1.IN.n247 VSS 0.188f
C4086 TG_1.IN.n248 VSS 0.0573f
C4087 TG_1.IN.n249 VSS 0.057f
C4088 TG_1.IN.t37 VSS 0.0197f
C4089 TG_1.IN.t83 VSS 0.0272f
C4090 TG_1.IN.n250 VSS 0.061f
C4091 TG_1.IN.n251 VSS 0.0293f
C4092 TG_1.IN.t84 VSS 0.0263f
C4093 TG_1.IN.t74 VSS 0.0536f
C4094 TG_1.IN.t52 VSS 0.0315f
C4095 TG_1.IN.n252 VSS 0.0334f
C4096 TG_1.IN.n253 VSS 0.0157f
C4097 TG_1.IN.n254 VSS 0.0324f
C4098 TG_1.IN.t27 VSS 0.0473f
C4099 TG_1.IN.t28 VSS 0.0379f
C4100 TG_1.IN.n255 VSS 0.275f
C4101 TG_1.IN.t124 VSS 0.0351f
C4102 TG_1.IN.n256 VSS 0.238f
C4103 TG_1.IN.n257 VSS 0.177f
C4104 TG_1.IN.t34 VSS 0.0315f
C4105 TG_1.IN.n258 VSS 0.0329f
C4106 TG_1.IN.n259 VSS 0.0715f
C4107 TG_1.IN.t51 VSS 0.0232f
C4108 TG_1.IN.t73 VSS 0.0889f
C4109 TG_1.IN.n260 VSS 0.11f
C4110 TG_1.IN.t33 VSS 0.0644f
C4111 TG_1.IN.n261 VSS 0.0765f
C4112 TG_1.IN.n262 VSS 0.0452f
C4113 TG_1.IN.n263 VSS 0.087f
C4114 TG_1.IN.n264 VSS 0.127f
C4115 TG_1.IN.t135 VSS 0.0157f
C4116 TG_1.IN.n265 VSS 0.0157f
C4117 TG_1.IN.n266 VSS 0.0786f
C4118 TG_1.IN.t115 VSS 0.0365f
C4119 TG_1.IN.t91 VSS 0.0428f
C4120 TG_1.IN.t92 VSS 0.0366f
C4121 TG_1.IN.n267 VSS 0.217f
C4122 TG_1.IN.n268 VSS 0.174f
C4123 TG_1.IN.n269 VSS 0.433f
C4124 TG_1.IN.t116 VSS 0.0356f
C4125 TG_1.IN.n270 VSS 0.26f
C4126 TG_1.IN.n271 VSS 0.155f
C4127 TG_1.IN.n272 VSS 0.0536f
C4128 TG_1.IN.n273 VSS 0.0516f
C4129 TG_1.IN.n274 VSS 1.51f
C4130 TG_1.IN.t197 VSS 0.0524f
C4131 TG_1.IN.n275 VSS 0.0524f
C4132 TG_1.IN.n276 VSS 0.105f
C4133 TG_1.IN.t179 VSS 0.0524f
C4134 TG_1.IN.n277 VSS 0.0524f
C4135 TG_1.IN.n278 VSS 0.138f
C4136 TG_1.IN.n279 VSS 0.186f
C4137 TG_1.IN.t215 VSS 0.0524f
C4138 TG_1.IN.n280 VSS 0.0524f
C4139 TG_1.IN.n281 VSS 0.105f
C4140 TG_1.IN.t157 VSS 0.0524f
C4141 TG_1.IN.n282 VSS 0.0524f
C4142 TG_1.IN.n283 VSS 0.138f
C4143 TG_1.IN.n284 VSS 0.186f
C4144 TG_1.IN.t201 VSS 0.0524f
C4145 TG_1.IN.n285 VSS 0.0524f
C4146 TG_1.IN.n286 VSS 0.105f
C4147 TG_1.IN.t143 VSS 0.0524f
C4148 TG_1.IN.n287 VSS 0.0524f
C4149 TG_1.IN.n288 VSS 0.138f
C4150 TG_1.IN.n289 VSS 0.186f
C4151 TG_1.IN.t202 VSS 0.0524f
C4152 TG_1.IN.n290 VSS 0.0524f
C4153 TG_1.IN.n291 VSS 0.105f
C4154 TG_1.IN.t144 VSS 0.0524f
C4155 TG_1.IN.n292 VSS 0.0524f
C4156 TG_1.IN.n293 VSS 0.138f
C4157 TG_1.IN.n294 VSS 0.186f
C4158 TG_1.IN.t186 VSS 0.0524f
C4159 TG_1.IN.n295 VSS 0.0524f
C4160 TG_1.IN.n296 VSS 0.105f
C4161 TG_1.IN.t168 VSS 0.0524f
C4162 TG_1.IN.n297 VSS 0.0524f
C4163 TG_1.IN.n298 VSS 0.138f
C4164 TG_1.IN.n299 VSS 0.186f
C4165 TG_1.IN.t216 VSS 0.0524f
C4166 TG_1.IN.n300 VSS 0.0524f
C4167 TG_1.IN.n301 VSS 0.105f
C4168 TG_1.IN.t158 VSS 0.0524f
C4169 TG_1.IN.n302 VSS 0.0524f
C4170 TG_1.IN.n303 VSS 0.138f
C4171 TG_1.IN.n304 VSS 0.186f
C4172 TG_1.IN.t206 VSS 0.0524f
C4173 TG_1.IN.n305 VSS 0.0524f
C4174 TG_1.IN.n306 VSS 0.105f
C4175 TG_1.IN.t148 VSS 0.0524f
C4176 TG_1.IN.n307 VSS 0.0524f
C4177 TG_1.IN.n308 VSS 0.138f
C4178 TG_1.IN.n309 VSS 0.186f
C4179 TG_1.IN.t193 VSS 0.0524f
C4180 TG_1.IN.n310 VSS 0.0524f
C4181 TG_1.IN.n311 VSS 0.105f
C4182 TG_1.IN.t175 VSS 0.0524f
C4183 TG_1.IN.n312 VSS 0.0524f
C4184 TG_1.IN.n313 VSS 0.138f
C4185 TG_1.IN.n314 VSS 0.186f
C4186 TG_1.IN.t219 VSS 0.0524f
C4187 TG_1.IN.n315 VSS 0.0524f
C4188 TG_1.IN.n316 VSS 0.105f
C4189 TG_1.IN.t161 VSS 0.0524f
C4190 TG_1.IN.n317 VSS 0.0524f
C4191 TG_1.IN.n318 VSS 0.138f
C4192 TG_1.IN.n319 VSS 0.186f
C4193 TG_1.IN.t205 VSS 0.0524f
C4194 TG_1.IN.n320 VSS 0.0524f
C4195 TG_1.IN.n321 VSS 0.105f
C4196 TG_1.IN.t147 VSS 0.0524f
C4197 TG_1.IN.n322 VSS 0.0524f
C4198 TG_1.IN.n323 VSS 0.138f
C4199 TG_1.IN.n324 VSS 0.186f
C4200 TG_1.IN.t192 VSS 0.0524f
C4201 TG_1.IN.n325 VSS 0.0524f
C4202 TG_1.IN.n326 VSS 0.105f
C4203 TG_1.IN.t174 VSS 0.0524f
C4204 TG_1.IN.n327 VSS 0.0524f
C4205 TG_1.IN.n328 VSS 0.138f
C4206 TG_1.IN.n329 VSS 0.186f
C4207 TG_1.IN.t211 VSS 0.0524f
C4208 TG_1.IN.n330 VSS 0.0524f
C4209 TG_1.IN.n331 VSS 0.105f
C4210 TG_1.IN.t153 VSS 0.0524f
C4211 TG_1.IN.n332 VSS 0.0524f
C4212 TG_1.IN.n333 VSS 0.138f
C4213 TG_1.IN.n334 VSS 0.186f
C4214 TG_1.IN.t194 VSS 0.0524f
C4215 TG_1.IN.n335 VSS 0.0524f
C4216 TG_1.IN.n336 VSS 0.105f
C4217 TG_1.IN.t176 VSS 0.0524f
C4218 TG_1.IN.n337 VSS 0.0524f
C4219 TG_1.IN.n338 VSS 0.138f
C4220 TG_1.IN.n339 VSS 0.186f
C4221 TG_1.IN.t199 VSS 0.0524f
C4222 TG_1.IN.n340 VSS 0.0524f
C4223 TG_1.IN.n341 VSS 0.105f
C4224 TG_1.IN.t181 VSS 0.0524f
C4225 TG_1.IN.n342 VSS 0.0524f
C4226 TG_1.IN.n343 VSS 0.138f
C4227 TG_1.IN.n344 VSS 0.186f
C4228 TG_1.IN.t183 VSS 0.0524f
C4229 TG_1.IN.n345 VSS 0.0524f
C4230 TG_1.IN.n346 VSS 0.105f
C4231 TG_1.IN.t165 VSS 0.0524f
C4232 TG_1.IN.n347 VSS 0.0524f
C4233 TG_1.IN.n348 VSS 0.138f
C4234 TG_1.IN.n349 VSS 0.186f
C4235 TG_1.IN.t207 VSS 0.0524f
C4236 TG_1.IN.n350 VSS 0.0524f
C4237 TG_1.IN.n351 VSS 0.105f
C4238 TG_1.IN.t149 VSS 0.0524f
C4239 TG_1.IN.n352 VSS 0.0524f
C4240 TG_1.IN.n353 VSS 0.138f
C4241 TG_1.IN.n354 VSS 0.186f
C4242 TG_1.IN.t218 VSS 0.0524f
C4243 TG_1.IN.n355 VSS 0.0524f
C4244 TG_1.IN.n356 VSS 0.105f
C4245 TG_1.IN.t160 VSS 0.0524f
C4246 TG_1.IN.n357 VSS 0.0524f
C4247 TG_1.IN.n358 VSS 0.138f
C4248 TG_1.IN.n359 VSS 0.186f
C4249 TG_1.IN.t191 VSS 0.0524f
C4250 TG_1.IN.n360 VSS 0.0524f
C4251 TG_1.IN.n361 VSS 0.105f
C4252 TG_1.IN.t173 VSS 0.0524f
C4253 TG_1.IN.n362 VSS 0.0524f
C4254 TG_1.IN.n363 VSS 0.138f
C4255 TG_1.IN.n364 VSS 0.186f
C4256 TG_1.IN.t190 VSS 0.145f
C4257 TG_1.IN.t172 VSS 0.186f
C4258 TG_1.IN.n365 VSS 0.291f
C4259 TG_1.IN.n366 VSS 0.362f
C4260 TG_1.IN.n367 VSS 0.253f
C4261 TG_1.IN.n368 VSS 0.253f
C4262 TG_1.IN.n369 VSS 0.253f
C4263 TG_1.IN.t155 VSS 0.0524f
C4264 TG_1.IN.n370 VSS 0.0524f
C4265 TG_1.IN.n371 VSS 0.138f
C4266 TG_1.IN.t213 VSS 0.0524f
C4267 TG_1.IN.n372 VSS 0.0524f
C4268 TG_1.IN.n373 VSS 0.105f
C4269 TG_1.IN.n374 VSS 0.186f
C4270 TG_1.IN.n375 VSS 0.253f
C4271 TG_1.IN.n376 VSS 0.253f
C4272 TG_1.IN.n377 VSS 0.253f
C4273 TG_1.IN.n378 VSS 0.253f
C4274 TG_1.IN.n379 VSS 0.253f
C4275 TG_1.IN.n380 VSS 0.253f
C4276 TG_1.IN.n381 VSS 0.253f
C4277 TG_1.IN.n382 VSS 0.253f
C4278 TG_1.IN.n383 VSS 0.253f
C4279 TG_1.IN.n384 VSS 0.253f
C4280 TG_1.IN.n385 VSS 0.253f
C4281 TG_1.IN.n386 VSS 0.253f
C4282 TG_1.IN.n387 VSS 0.253f
C4283 TG_1.IN.n388 VSS 0.253f
C4284 TG_1.IN.n389 VSS 0.371f
C4285 TG_1.IN.n390 VSS 0.145f
C4286 TG_1.IN.n391 VSS 0.349f
C4287 TG_1.IN.n392 VSS 0.154f
C4288 TG_1.IN.n393 VSS 0.527f
C4289 TG_1.IN.n394 VSS 2.4f
C4290 OUT-.t43 VSS 0.0489f
C4291 OUT-.n0 VSS 0.0489f
C4292 OUT-.n1 VSS 0.133f
C4293 OUT-.t14 VSS 0.0489f
C4294 OUT-.n2 VSS 0.0489f
C4295 OUT-.n3 VSS 0.0977f
C4296 OUT-.n4 VSS 0.17f
C4297 OUT-.t57 VSS 0.0489f
C4298 OUT-.n5 VSS 0.0489f
C4299 OUT-.n6 VSS 0.133f
C4300 OUT-.t8 VSS 0.0489f
C4301 OUT-.n7 VSS 0.0489f
C4302 OUT-.n8 VSS 0.0977f
C4303 OUT-.n9 VSS 0.17f
C4304 OUT-.t51 VSS 0.0489f
C4305 OUT-.n10 VSS 0.0489f
C4306 OUT-.n11 VSS 0.133f
C4307 OUT-.t2 VSS 0.0489f
C4308 OUT-.n12 VSS 0.0489f
C4309 OUT-.n13 VSS 0.0977f
C4310 OUT-.n14 VSS 0.17f
C4311 OUT-.t46 VSS 0.0489f
C4312 OUT-.n15 VSS 0.0489f
C4313 OUT-.n16 VSS 0.133f
C4314 OUT-.t17 VSS 0.0489f
C4315 OUT-.n17 VSS 0.0489f
C4316 OUT-.n18 VSS 0.0977f
C4317 OUT-.n19 VSS 0.17f
C4318 OUT-.t59 VSS 0.0489f
C4319 OUT-.n20 VSS 0.0489f
C4320 OUT-.n21 VSS 0.133f
C4321 OUT-.t10 VSS 0.0489f
C4322 OUT-.n22 VSS 0.0489f
C4323 OUT-.n23 VSS 0.0977f
C4324 OUT-.n24 VSS 0.17f
C4325 OUT-.t54 VSS 0.0489f
C4326 OUT-.n25 VSS 0.0489f
C4327 OUT-.n26 VSS 0.133f
C4328 OUT-.t5 VSS 0.0489f
C4329 OUT-.n27 VSS 0.0489f
C4330 OUT-.n28 VSS 0.0977f
C4331 OUT-.n29 VSS 0.17f
C4332 OUT-.t41 VSS 0.0489f
C4333 OUT-.n30 VSS 0.0489f
C4334 OUT-.n31 VSS 0.133f
C4335 OUT-.t12 VSS 0.0489f
C4336 OUT-.n32 VSS 0.0489f
C4337 OUT-.n33 VSS 0.0977f
C4338 OUT-.n34 VSS 0.17f
C4339 OUT-.t52 VSS 0.0489f
C4340 OUT-.n35 VSS 0.0489f
C4341 OUT-.n36 VSS 0.133f
C4342 OUT-.t3 VSS 0.0489f
C4343 OUT-.n37 VSS 0.0489f
C4344 OUT-.n38 VSS 0.0977f
C4345 OUT-.n39 VSS 0.17f
C4346 OUT-.t58 VSS 0.0489f
C4347 OUT-.n40 VSS 0.0489f
C4348 OUT-.n41 VSS 0.133f
C4349 OUT-.t9 VSS 0.0489f
C4350 OUT-.n42 VSS 0.0489f
C4351 OUT-.n43 VSS 0.0977f
C4352 OUT-.n44 VSS 0.17f
C4353 OUT-.t45 VSS 0.0489f
C4354 OUT-.n45 VSS 0.0489f
C4355 OUT-.n46 VSS 0.133f
C4356 OUT-.t16 VSS 0.0489f
C4357 OUT-.n47 VSS 0.0489f
C4358 OUT-.n48 VSS 0.0977f
C4359 OUT-.n49 VSS 0.17f
C4360 OUT-.t53 VSS 0.0489f
C4361 OUT-.n50 VSS 0.0489f
C4362 OUT-.n51 VSS 0.133f
C4363 OUT-.t4 VSS 0.0489f
C4364 OUT-.n52 VSS 0.0489f
C4365 OUT-.n53 VSS 0.0977f
C4366 OUT-.n54 VSS 0.17f
C4367 OUT-.t44 VSS 0.0489f
C4368 OUT-.n55 VSS 0.0489f
C4369 OUT-.n56 VSS 0.133f
C4370 OUT-.t15 VSS 0.0489f
C4371 OUT-.n57 VSS 0.0489f
C4372 OUT-.n58 VSS 0.0977f
C4373 OUT-.n59 VSS 0.17f
C4374 OUT-.t50 VSS 0.0489f
C4375 OUT-.n60 VSS 0.0489f
C4376 OUT-.n61 VSS 0.133f
C4377 OUT-.t1 VSS 0.0489f
C4378 OUT-.n62 VSS 0.0489f
C4379 OUT-.n63 VSS 0.0977f
C4380 OUT-.n64 VSS 0.17f
C4381 OUT-.t49 VSS 0.0489f
C4382 OUT-.n65 VSS 0.0489f
C4383 OUT-.n66 VSS 0.133f
C4384 OUT-.t0 VSS 0.0489f
C4385 OUT-.n67 VSS 0.0489f
C4386 OUT-.n68 VSS 0.0977f
C4387 OUT-.n69 VSS 0.17f
C4388 OUT-.t56 VSS 0.0489f
C4389 OUT-.n70 VSS 0.0489f
C4390 OUT-.n71 VSS 0.133f
C4391 OUT-.t7 VSS 0.0489f
C4392 OUT-.n72 VSS 0.0489f
C4393 OUT-.n73 VSS 0.0977f
C4394 OUT-.n74 VSS 0.17f
C4395 OUT-.t42 VSS 0.0489f
C4396 OUT-.n75 VSS 0.0489f
C4397 OUT-.n76 VSS 0.133f
C4398 OUT-.t13 VSS 0.0489f
C4399 OUT-.n77 VSS 0.0489f
C4400 OUT-.n78 VSS 0.0977f
C4401 OUT-.n79 VSS 0.17f
C4402 OUT-.t48 VSS 0.0489f
C4403 OUT-.n80 VSS 0.0489f
C4404 OUT-.n81 VSS 0.133f
C4405 OUT-.t19 VSS 0.0489f
C4406 OUT-.n82 VSS 0.0489f
C4407 OUT-.n83 VSS 0.0977f
C4408 OUT-.n84 VSS 0.17f
C4409 OUT-.t55 VSS 0.0489f
C4410 OUT-.n85 VSS 0.0489f
C4411 OUT-.n86 VSS 0.133f
C4412 OUT-.t6 VSS 0.0489f
C4413 OUT-.n87 VSS 0.0489f
C4414 OUT-.n88 VSS 0.0977f
C4415 OUT-.n89 VSS 0.17f
C4416 OUT-.t40 VSS 0.0489f
C4417 OUT-.n90 VSS 0.0489f
C4418 OUT-.n91 VSS 0.133f
C4419 OUT-.t11 VSS 0.0489f
C4420 OUT-.n92 VSS 0.0489f
C4421 OUT-.n93 VSS 0.0977f
C4422 OUT-.n94 VSS 0.17f
C4423 OUT-.t47 VSS 0.0489f
C4424 OUT-.n95 VSS 0.0489f
C4425 OUT-.n96 VSS 0.133f
C4426 OUT-.t18 VSS 0.0489f
C4427 OUT-.n97 VSS 0.0489f
C4428 OUT-.n98 VSS 0.0977f
C4429 OUT-.n99 VSS 0.213f
C4430 OUT-.n100 VSS 0.313f
C4431 OUT-.n101 VSS 0.219f
C4432 OUT-.n102 VSS 0.219f
C4433 OUT-.n103 VSS 0.219f
C4434 OUT-.n104 VSS 0.219f
C4435 OUT-.n105 VSS 0.219f
C4436 OUT-.n106 VSS 0.219f
C4437 OUT-.n107 VSS 0.219f
C4438 OUT-.n108 VSS 0.219f
C4439 OUT-.n109 VSS 0.219f
C4440 OUT-.n110 VSS 0.219f
C4441 OUT-.n111 VSS 0.219f
C4442 OUT-.n112 VSS 0.219f
C4443 OUT-.n113 VSS 0.219f
C4444 OUT-.n114 VSS 0.219f
C4445 OUT-.n115 VSS 0.219f
C4446 OUT-.n116 VSS 0.219f
C4447 OUT-.n117 VSS 0.219f
C4448 OUT-.n118 VSS 0.236f
C4449 a_n2280_5855.t4 VSS 0.0419f
C4450 a_n2280_5855.n0 VSS 0.0419f
C4451 a_n2280_5855.n1 VSS 0.0935f
C4452 a_n2280_5855.t9 VSS 0.0419f
C4453 a_n2280_5855.n2 VSS 0.0419f
C4454 a_n2280_5855.n3 VSS 0.0948f
C4455 a_n2280_5855.t5 VSS 0.0419f
C4456 a_n2280_5855.n4 VSS 0.0419f
C4457 a_n2280_5855.n5 VSS 0.0935f
C4458 a_n2280_5855.t10 VSS 0.0419f
C4459 a_n2280_5855.n6 VSS 0.0419f
C4460 a_n2280_5855.n7 VSS 0.0948f
C4461 a_n2280_5855.t1 VSS 0.0419f
C4462 a_n2280_5855.n8 VSS 0.0419f
C4463 a_n2280_5855.n9 VSS 0.0944f
C4464 a_n2280_5855.t37 VSS 0.0577f
C4465 a_n2280_5855.t50 VSS 0.0577f
C4466 a_n2280_5855.t19 VSS 0.0577f
C4467 a_n2280_5855.t20 VSS 0.0577f
C4468 a_n2280_5855.t33 VSS 0.0577f
C4469 a_n2280_5855.t34 VSS 0.0577f
C4470 a_n2280_5855.t32 VSS 0.0577f
C4471 a_n2280_5855.t47 VSS 0.0577f
C4472 a_n2280_5855.t48 VSS 0.0577f
C4473 a_n2280_5855.t17 VSS 0.0577f
C4474 a_n2280_5855.t18 VSS 0.0577f
C4475 a_n2280_5855.t31 VSS 0.0577f
C4476 a_n2280_5855.t28 VSS 0.0577f
C4477 a_n2280_5855.t30 VSS 0.0577f
C4478 a_n2280_5855.t41 VSS 0.0577f
C4479 a_n2280_5855.t45 VSS 0.0577f
C4480 a_n2280_5855.t15 VSS 0.0577f
C4481 a_n2280_5855.t24 VSS 0.0577f
C4482 a_n2280_5855.t29 VSS 0.0577f
C4483 a_n2280_5855.t39 VSS 0.0577f
C4484 a_n2280_5855.t42 VSS 0.0577f
C4485 a_n2280_5855.t13 VSS 0.0577f
C4486 a_n2280_5855.t23 VSS 0.0577f
C4487 a_n2280_5855.t25 VSS 0.0577f
C4488 a_n2280_5855.t40 VSS 0.0577f
C4489 a_n2280_5855.t49 VSS 0.0577f
C4490 a_n2280_5855.t35 VSS 0.0577f
C4491 a_n2280_5855.t22 VSS 0.0577f
C4492 a_n2280_5855.t21 VSS 0.0577f
C4493 a_n2280_5855.t12 VSS 0.0577f
C4494 a_n2280_5855.t51 VSS 0.0577f
C4495 a_n2280_5855.t38 VSS 0.0577f
C4496 a_n2280_5855.t27 VSS 0.0577f
C4497 a_n2280_5855.t26 VSS 0.0577f
C4498 a_n2280_5855.t16 VSS 0.0577f
C4499 a_n2280_5855.t14 VSS 0.0577f
C4500 a_n2280_5855.t43 VSS 0.0577f
C4501 a_n2280_5855.t46 VSS 0.0577f
C4502 a_n2280_5855.t44 VSS 0.0797f
C4503 a_n2280_5855.n10 VSS 0.0911f
C4504 a_n2280_5855.n11 VSS 0.0621f
C4505 a_n2280_5855.n12 VSS 0.0621f
C4506 a_n2280_5855.n13 VSS 0.0621f
C4507 a_n2280_5855.n14 VSS 0.0621f
C4508 a_n2280_5855.n15 VSS 0.0621f
C4509 a_n2280_5855.n16 VSS 0.0621f
C4510 a_n2280_5855.n17 VSS 0.0621f
C4511 a_n2280_5855.n18 VSS 0.0621f
C4512 a_n2280_5855.n19 VSS 0.0621f
C4513 a_n2280_5855.n20 VSS 0.0621f
C4514 a_n2280_5855.n21 VSS 0.0621f
C4515 a_n2280_5855.n22 VSS 0.0621f
C4516 a_n2280_5855.n23 VSS 0.0621f
C4517 a_n2280_5855.n24 VSS 0.0621f
C4518 a_n2280_5855.n25 VSS 0.0621f
C4519 a_n2280_5855.n26 VSS 0.0621f
C4520 a_n2280_5855.n27 VSS 0.0621f
C4521 a_n2280_5855.n28 VSS 0.0621f
C4522 a_n2280_5855.n29 VSS 0.0621f
C4523 a_n2280_5855.n30 VSS 0.0621f
C4524 a_n2280_5855.n31 VSS 0.0621f
C4525 a_n2280_5855.n32 VSS 0.0621f
C4526 a_n2280_5855.n33 VSS 0.0621f
C4527 a_n2280_5855.n34 VSS 0.0621f
C4528 a_n2280_5855.n35 VSS 0.0621f
C4529 a_n2280_5855.n36 VSS 0.0621f
C4530 a_n2280_5855.n37 VSS 0.0621f
C4531 a_n2280_5855.n38 VSS 0.0621f
C4532 a_n2280_5855.n39 VSS 0.0621f
C4533 a_n2280_5855.n40 VSS 0.0621f
C4534 a_n2280_5855.n41 VSS 0.0621f
C4535 a_n2280_5855.n42 VSS 0.0621f
C4536 a_n2280_5855.n43 VSS 0.0621f
C4537 a_n2280_5855.n44 VSS 0.0621f
C4538 a_n2280_5855.n45 VSS 0.0621f
C4539 a_n2280_5855.n46 VSS 0.0621f
C4540 a_n2280_5855.n47 VSS 0.0911f
C4541 a_n2280_5855.t36 VSS 0.143f
C4542 a_n2280_5855.n48 VSS 0.255f
C4543 a_n2280_5855.n49 VSS 0.216f
C4544 a_n2280_5855.n50 VSS 0.309f
C4545 a_n2280_5855.n51 VSS 0.0419f
C4546 a_n2280_5855.n52 VSS 0.112f
C4547 a_n2280_5855.t7 VSS 0.0419f
C4548 VDD.t116 VSS 0.0119f
C4549 VDD.t274 VSS 0.00497f
C4550 VDD.n0 VSS 0.00497f
C4551 VDD.n1 VSS 0.0119f
C4552 VDD.n2 VSS 0.0121f
C4553 VDD.t218 VSS 0.107f
C4554 VDD.n3 VSS 0.282f
C4555 VDD.t216 VSS 0.0987f
C4556 VDD.n4 VSS 0.107f
C4557 VDD.n5 VSS 0.0664f
C4558 VDD.t238 VSS 0.0987f
C4559 VDD.n6 VSS 0.107f
C4560 VDD.n7 VSS 0.0664f
C4561 VDD.t273 VSS 0.0987f
C4562 VDD.n8 VSS 0.107f
C4563 VDD.n9 VSS 0.0598f
C4564 VDD.n10 VSS 0.0471f
C4565 VDD.t233 VSS 0.0987f
C4566 VDD.n11 VSS 0.107f
C4567 VDD.n12 VSS 0.0455f
C4568 VDD.t217 VSS 0.0987f
C4569 VDD.n13 VSS 0.107f
C4570 VDD.n14 VSS 0.0664f
C4571 VDD.t237 VSS 0.0987f
C4572 VDD.n15 VSS 0.107f
C4573 VDD.n16 VSS 0.0664f
C4574 VDD.t115 VSS 0.0987f
C4575 VDD.n17 VSS 0.107f
C4576 VDD.n18 VSS 0.0567f
C4577 VDD.n19 VSS 0.0539f
C4578 VDD.n20 VSS 0.207f
C4579 VDD.n21 VSS 0.0383f
C4580 VDD.n22 VSS 0.0289f
C4581 VDD.n23 VSS 0.0738f
C4582 VDD.t41 VSS 0.129f
C4583 VDD.n24 VSS 0.107f
C4584 VDD.n25 VSS 0.0576f
C4585 VDD.t224 VSS 0.0987f
C4586 VDD.n26 VSS 0.107f
C4587 VDD.n27 VSS 0.0664f
C4588 VDD.t225 VSS 0.0987f
C4589 VDD.n28 VSS 0.107f
C4590 VDD.n29 VSS 0.0648f
C4591 VDD.n30 VSS 0.0274f
C4592 VDD.n31 VSS 0.00755f
C4593 VDD.n32 VSS 0.0715f
C4594 VDD.t145 VSS 0.0931f
C4595 VDD.n33 VSS 0.0245f
C4596 VDD.n34 VSS 0.00599f
C4597 VDD.n35 VSS 0.0216f
C4598 VDD.n36 VSS 0.00748f
C4599 VDD.n37 VSS 0.00671f
C4600 VDD.n38 VSS 0.00714f
C4601 VDD.n39 VSS 0.00536f
C4602 VDD.t146 VSS 0.00458f
C4603 VDD.n40 VSS 0.033f
C4604 VDD.n41 VSS 0.049f
C4605 VDD.t119 VSS 0.0837f
C4606 VDD.n42 VSS 0.107f
C4607 VDD.n43 VSS 0.0606f
C4608 VDD.t240 VSS 0.0987f
C4609 VDD.n44 VSS 0.107f
C4610 VDD.n45 VSS 0.0664f
C4611 VDD.t227 VSS 0.0987f
C4612 VDD.n46 VSS 0.107f
C4613 VDD.n47 VSS 0.064f
C4614 VDD.n48 VSS 0.0274f
C4615 VDD.n49 VSS 0.00587f
C4616 VDD.n50 VSS 0.0602f
C4617 VDD.t211 VSS 0.0903f
C4618 VDD.n51 VSS 0.0357f
C4619 VDD.n52 VSS 0.00525f
C4620 VDD.n53 VSS 0.0216f
C4621 VDD.n54 VSS 0.0101f
C4622 VDD.n55 VSS 0.00663f
C4623 VDD.n56 VSS 0.00625f
C4624 VDD.n57 VSS 0.00541f
C4625 VDD.t212 VSS 0.00454f
C4626 VDD.n58 VSS 0.0335f
C4627 VDD.n59 VSS 0.0504f
C4628 VDD.t112 VSS 0.0865f
C4629 VDD.n60 VSS 0.107f
C4630 VDD.n61 VSS 0.0617f
C4631 VDD.t210 VSS 0.0987f
C4632 VDD.n62 VSS 0.107f
C4633 VDD.n63 VSS 0.0664f
C4634 VDD.t209 VSS 0.0987f
C4635 VDD.n64 VSS 0.107f
C4636 VDD.n65 VSS 0.0619f
C4637 VDD.n66 VSS 0.0274f
C4638 VDD.n67 VSS 0.0258f
C4639 VDD.n68 VSS 0.00792f
C4640 VDD.n69 VSS 0.00576f
C4641 VDD.n70 VSS 0.00532f
C4642 VDD.t40 VSS 0.00462f
C4643 VDD.n71 VSS 0.0399f
C4644 VDD.n72 VSS 0.0282f
C4645 VDD.t39 VSS 0.0828f
C4646 VDD.n73 VSS 0.047f
C4647 VDD.n74 VSS 0.00746f
C4648 VDD.t142 VSS 0.0835f
C4649 VDD.n75 VSS 0.0553f
C4650 VDD.n76 VSS 0.0057f
C4651 VDD.n77 VSS 0.0242f
C4652 VDD.t239 VSS 0.0987f
C4653 VDD.n78 VSS 0.107f
C4654 VDD.n79 VSS 0.0644f
C4655 VDD.t226 VSS 0.0987f
C4656 VDD.n80 VSS 0.107f
C4657 VDD.n81 VSS 0.0664f
C4658 VDD.t147 VSS 0.086f
C4659 VDD.n82 VSS 0.107f
C4660 VDD.n83 VSS 0.0616f
C4661 VDD.t148 VSS 0.0262f
C4662 VDD.n84 VSS 0.0663f
C4663 VDD.n85 VSS 0.00628f
C4664 VDD.n86 VSS 0.104f
C4665 VDD.n87 VSS 0.00718f
C4666 VDD.n88 VSS 0.0583f
C4667 VDD.n89 VSS 0.00552f
C4668 VDD.n90 VSS 0.0216f
C4669 VDD.n91 VSS 0.00841f
C4670 VDD.n92 VSS 0.00667f
C4671 VDD.n93 VSS 0.00523f
C4672 VDD.n94 VSS 0.0119f
C4673 VDD.t228 VSS 0.0987f
C4674 VDD.n95 VSS 0.152f
C4675 VDD.t215 VSS 0.0987f
C4676 VDD.n96 VSS 0.107f
C4677 VDD.t213 VSS 0.0987f
C4678 VDD.n97 VSS 0.107f
C4679 VDD.t231 VSS 0.0969f
C4680 VDD.n98 VSS 0.107f
C4681 VDD.t232 VSS 0.00497f
C4682 VDD.n99 VSS 0.00497f
C4683 VDD.n100 VSS 0.0119f
C4684 VDD.n101 VSS 0.0625f
C4685 VDD.t270 VSS 0.0799f
C4686 VDD.n102 VSS 0.0334f
C4687 VDD.n103 VSS 0.0143f
C4688 VDD.n104 VSS 0.0217f
C4689 VDD.n105 VSS 0.00661f
C4690 VDD.n106 VSS 0.021f
C4691 VDD.n107 VSS 0.0209f
C4692 VDD.n108 VSS 0.0249f
C4693 VDD.n109 VSS 0.00535f
C4694 VDD.n110 VSS 0.0645f
C4695 VDD.n111 VSS 0.0426f
C4696 VDD.n112 VSS 0.00834f
C4697 VDD.n113 VSS 0.147f
C4698 VDD.t167 VSS 0.0166f
C4699 VDD.n114 VSS 0.0166f
C4700 VDD.n115 VSS 0.0368f
C4701 VDD.t177 VSS 0.0166f
C4702 VDD.n116 VSS 0.0166f
C4703 VDD.n117 VSS 0.0368f
C4704 VDD.t192 VSS 0.0166f
C4705 VDD.n118 VSS 0.0166f
C4706 VDD.n119 VSS 0.0368f
C4707 VDD.n120 VSS 0.0499f
C4708 VDD.n121 VSS 0.189f
C4709 VDD.n122 VSS 0.0856f
C4710 VDD.t193 VSS 0.118f
C4711 VDD.t191 VSS 0.114f
C4712 VDD.n123 VSS 0.0912f
C4713 VDD.n124 VSS 0.0281f
C4714 VDD.n125 VSS 0.036f
C4715 VDD.n126 VSS 0.0512f
C4716 VDD.n127 VSS 0.0165f
C4717 VDD.t178 VSS 0.105f
C4718 VDD.n128 VSS 0.0912f
C4719 VDD.n129 VSS 0.0281f
C4720 VDD.t176 VSS 0.0997f
C4721 VDD.n130 VSS 0.0912f
C4722 VDD.n131 VSS 0.0281f
C4723 VDD.n132 VSS 0.0194f
C4724 VDD.n133 VSS 0.0512f
C4725 VDD.t181 VSS 0.114f
C4726 VDD.n134 VSS 0.0912f
C4727 VDD.n135 VSS 0.0281f
C4728 VDD.n136 VSS 0.036f
C4729 VDD.n137 VSS 0.0512f
C4730 VDD.t166 VSS 0.114f
C4731 VDD.t163 VSS 0.114f
C4732 VDD.n138 VSS 0.0912f
C4733 VDD.n139 VSS 0.0281f
C4734 VDD.n140 VSS 0.0242f
C4735 VDD.t156 VSS 0.101f
C4736 VDD.n141 VSS 0.0912f
C4737 VDD.n142 VSS 0.0269f
C4738 VDD.n143 VSS 0.0315f
C4739 VDD.t157 VSS 0.0501f
C4740 VDD.n144 VSS 0.076f
C4741 VDD.n145 VSS 0.257f
C4742 VDD.n146 VSS 0.022f
C4743 VDD.n147 VSS 0.0466f
C4744 VDD.t201 VSS 0.148f
C4745 VDD.n148 VSS 0.192f
C4746 VDD.n149 VSS 0.0281f
C4747 VDD.n150 VSS 0.0449f
C4748 VDD.t202 VSS 0.133f
C4749 VDD.n151 VSS 0.118f
C4750 VDD.n152 VSS 0.0281f
C4751 VDD.n153 VSS 0.0449f
C4752 VDD.t155 VSS 0.133f
C4753 VDD.n154 VSS 0.118f
C4754 VDD.n155 VSS 0.0281f
C4755 VDD.n156 VSS 0.0449f
C4756 VDD.t317 VSS 0.148f
C4757 VDD.n157 VSS 0.118f
C4758 VDD.n158 VSS 0.0281f
C4759 VDD.n159 VSS 0.0449f
C4760 VDD.t308 VSS 0.148f
C4761 VDD.t205 VSS 0.148f
C4762 VDD.n160 VSS 0.118f
C4763 VDD.n161 VSS 0.0281f
C4764 VDD.n162 VSS 0.0449f
C4765 VDD.t206 VSS 0.133f
C4766 VDD.n163 VSS 0.118f
C4767 VDD.n164 VSS 0.0269f
C4768 VDD.n165 VSS 0.0478f
C4769 VDD.t204 VSS 0.151f
C4770 VDD.n166 VSS 0.118f
C4771 VDD.n167 VSS 0.022f
C4772 VDD.n168 VSS 0.0478f
C4773 VDD.t152 VSS 0.148f
C4774 VDD.t153 VSS 0.148f
C4775 VDD.n169 VSS 0.118f
C4776 VDD.n170 VSS 0.0281f
C4777 VDD.n171 VSS 0.0449f
C4778 VDD.t315 VSS 0.144f
C4779 VDD.n172 VSS 0.118f
C4780 VDD.n173 VSS 0.0281f
C4781 VDD.n174 VSS 0.0449f
C4782 VDD.t316 VSS 0.122f
C4783 VDD.n175 VSS 0.118f
C4784 VDD.n176 VSS 0.0281f
C4785 VDD.n177 VSS 0.0449f
C4786 VDD.t97 VSS 0.148f
C4787 VDD.n178 VSS 0.118f
C4788 VDD.n179 VSS 0.0281f
C4789 VDD.n180 VSS 0.0449f
C4790 VDD.t320 VSS 0.148f
C4791 VDD.t96 VSS 0.148f
C4792 VDD.n181 VSS 0.118f
C4793 VDD.n182 VSS 0.0281f
C4794 VDD.n183 VSS 0.0449f
C4795 VDD.t277 VSS 0.144f
C4796 VDD.n184 VSS 0.118f
C4797 VDD.n185 VSS 0.0269f
C4798 VDD.n186 VSS 0.0478f
C4799 VDD.t198 VSS 0.14f
C4800 VDD.n187 VSS 0.118f
C4801 VDD.n188 VSS 0.022f
C4802 VDD.n189 VSS 0.0478f
C4803 VDD.t282 VSS 0.148f
C4804 VDD.t150 VSS 0.148f
C4805 VDD.n190 VSS 0.118f
C4806 VDD.n191 VSS 0.0281f
C4807 VDD.n192 VSS 0.0449f
C4808 VDD.t95 VSS 0.148f
C4809 VDD.n193 VSS 0.118f
C4810 VDD.n194 VSS 0.0281f
C4811 VDD.n195 VSS 0.0449f
C4812 VDD.t275 VSS 0.125f
C4813 VDD.n196 VSS 0.118f
C4814 VDD.n197 VSS 0.0281f
C4815 VDD.n198 VSS 0.0449f
C4816 VDD.t278 VSS 0.14f
C4817 VDD.n199 VSS 0.118f
C4818 VDD.n200 VSS 0.0281f
C4819 VDD.n201 VSS 0.0449f
C4820 VDD.t280 VSS 0.148f
C4821 VDD.t149 VSS 0.148f
C4822 VDD.n202 VSS 0.118f
C4823 VDD.n203 VSS 0.0281f
C4824 VDD.n204 VSS 0.0449f
C4825 VDD.t151 VSS 0.155f
C4826 VDD.n205 VSS 0.118f
C4827 VDD.n206 VSS 0.0269f
C4828 VDD.n207 VSS 0.0478f
C4829 VDD.t276 VSS 0.129f
C4830 VDD.n208 VSS 0.118f
C4831 VDD.n209 VSS 0.022f
C4832 VDD.n210 VSS 0.0478f
C4833 VDD.t154 VSS 0.148f
C4834 VDD.n211 VSS 0.118f
C4835 VDD.n212 VSS 0.0281f
C4836 VDD.n213 VSS 0.0449f
C4837 VDD.t200 VSS 0.148f
C4838 VDD.t310 VSS 0.148f
C4839 VDD.n214 VSS 0.118f
C4840 VDD.n215 VSS 0.0281f
C4841 VDD.n216 VSS 0.0449f
C4842 VDD.t309 VSS 0.137f
C4843 VDD.n217 VSS 0.118f
C4844 VDD.n218 VSS 0.0281f
C4845 VDD.n219 VSS 0.0449f
C4846 VDD.t279 VSS 0.129f
C4847 VDD.n220 VSS 0.118f
C4848 VDD.n221 VSS 0.0281f
C4849 VDD.n222 VSS 0.0449f
C4850 VDD.t311 VSS 0.148f
C4851 VDD.n223 VSS 0.118f
C4852 VDD.n224 VSS 0.0281f
C4853 VDD.n225 VSS 0.0449f
C4854 VDD.t203 VSS 0.148f
C4855 VDD.t319 VSS 0.166f
C4856 VDD.n226 VSS 0.118f
C4857 VDD.n227 VSS 0.0269f
C4858 VDD.n228 VSS 0.0478f
C4859 VDD.t318 VSS 0.236f
C4860 VDD.n229 VSS 0.022f
C4861 VDD.n230 VSS 0.0478f
C4862 VDD.t314 VSS 0.148f
C4863 VDD.n231 VSS 0.118f
C4864 VDD.n232 VSS 0.0281f
C4865 VDD.n233 VSS 0.0354f
C4866 VDD.n234 VSS 0.0303f
C4867 VDD.t281 VSS 0.148f
C4868 VDD.t196 VSS 0.148f
C4869 VDD.n235 VSS 0.118f
C4870 VDD.n236 VSS 0.0281f
C4871 VDD.n237 VSS 0.0365f
C4872 VDD.n238 VSS 0.0276f
C4873 VDD.n239 VSS 0.00834f
C4874 VDD.t199 VSS 0.136f
C4875 VDD.n240 VSS 0.118f
C4876 VDD.n241 VSS 0.0269f
C4877 VDD.n242 VSS 0.0082f
C4878 VDD.n243 VSS 0.0274f
C4879 VDD.n244 VSS 0.118f
C4880 VDD.n245 VSS 0.014f
C4881 VDD.n246 VSS 0.0238f
C4882 VDD.n247 VSS 0.00477f
C4883 VDD.n248 VSS 0.00224f
C4884 VDD.t197 VSS 0.0828f
C4885 VDD.n249 VSS 0.205f
C4886 VDD.n250 VSS 0.0961f
C4887 VDD.n251 VSS 0.0082f
C4888 VDD.n252 VSS 0.0384f
C4889 VDD.n253 VSS 0.0761f
C4890 VDD.n254 VSS 0.454f
C4891 VDD.n255 VSS 0.118f
C4892 VDD.n256 VSS 0.0337f
C4893 VDD.n257 VSS 0.0291f
C4894 VDD.n258 VSS 0.0271f
C4895 VDD.n259 VSS 0.00759f
C4896 VDD.n260 VSS 0.00759f
C4897 VDD.n261 VSS 0.0204f
C4898 VDD.n262 VSS 0.0219f
C4899 VDD.t162 VSS 0.0166f
C4900 VDD.n263 VSS 0.0166f
C4901 VDD.n264 VSS 0.0368f
C4902 VDD.t169 VSS 0.0166f
C4903 VDD.n265 VSS 0.0166f
C4904 VDD.n266 VSS 0.0368f
C4905 VDD.t185 VSS 0.0166f
C4906 VDD.n267 VSS 0.0166f
C4907 VDD.n268 VSS 0.0368f
C4908 VDD.n269 VSS 0.0499f
C4909 VDD.n270 VSS 0.189f
C4910 VDD.n271 VSS 0.0856f
C4911 VDD.t186 VSS 0.118f
C4912 VDD.t184 VSS 0.114f
C4913 VDD.n272 VSS 0.0912f
C4914 VDD.n273 VSS 0.0281f
C4915 VDD.n274 VSS 0.036f
C4916 VDD.n275 VSS 0.0512f
C4917 VDD.n276 VSS 0.0165f
C4918 VDD.t170 VSS 0.105f
C4919 VDD.n277 VSS 0.0912f
C4920 VDD.n278 VSS 0.0281f
C4921 VDD.t168 VSS 0.0997f
C4922 VDD.n279 VSS 0.0912f
C4923 VDD.n280 VSS 0.0281f
C4924 VDD.n281 VSS 0.0194f
C4925 VDD.n282 VSS 0.0512f
C4926 VDD.t173 VSS 0.114f
C4927 VDD.n283 VSS 0.0912f
C4928 VDD.n284 VSS 0.0281f
C4929 VDD.n285 VSS 0.036f
C4930 VDD.n286 VSS 0.0512f
C4931 VDD.t161 VSS 0.114f
C4932 VDD.t158 VSS 0.114f
C4933 VDD.n287 VSS 0.0912f
C4934 VDD.n288 VSS 0.0281f
C4935 VDD.n289 VSS 0.0242f
C4936 VDD.t189 VSS 0.101f
C4937 VDD.n290 VSS 0.0912f
C4938 VDD.n291 VSS 0.0269f
C4939 VDD.n292 VSS 0.0315f
C4940 VDD.t190 VSS 0.0501f
C4941 VDD.n293 VSS 0.076f
C4942 VDD.n294 VSS 0.257f
C4943 VDD.n295 VSS 0.022f
C4944 VDD.n296 VSS 0.0466f
C4945 VDD.t290 VSS 0.148f
C4946 VDD.n297 VSS 0.192f
C4947 VDD.n298 VSS 0.0281f
C4948 VDD.n299 VSS 0.0449f
C4949 VDD.t291 VSS 0.133f
C4950 VDD.n300 VSS 0.118f
C4951 VDD.n301 VSS 0.0281f
C4952 VDD.n302 VSS 0.0449f
C4953 VDD.t305 VSS 0.133f
C4954 VDD.n303 VSS 0.118f
C4955 VDD.n304 VSS 0.0281f
C4956 VDD.n305 VSS 0.0449f
C4957 VDD.t297 VSS 0.148f
C4958 VDD.n306 VSS 0.118f
C4959 VDD.n307 VSS 0.0281f
C4960 VDD.n308 VSS 0.0449f
C4961 VDD.t299 VSS 0.148f
C4962 VDD.t339 VSS 0.148f
C4963 VDD.n309 VSS 0.118f
C4964 VDD.n310 VSS 0.0281f
C4965 VDD.n311 VSS 0.0449f
C4966 VDD.t289 VSS 0.133f
C4967 VDD.n312 VSS 0.118f
C4968 VDD.n313 VSS 0.0269f
C4969 VDD.n314 VSS 0.0478f
C4970 VDD.t337 VSS 0.151f
C4971 VDD.n315 VSS 0.118f
C4972 VDD.n316 VSS 0.022f
C4973 VDD.n317 VSS 0.0478f
C4974 VDD.t139 VSS 0.148f
C4975 VDD.t301 VSS 0.148f
C4976 VDD.n318 VSS 0.118f
C4977 VDD.n319 VSS 0.0281f
C4978 VDD.n320 VSS 0.0449f
C4979 VDD.t288 VSS 0.144f
C4980 VDD.n321 VSS 0.118f
C4981 VDD.n322 VSS 0.0281f
C4982 VDD.n323 VSS 0.0449f
C4983 VDD.t295 VSS 0.122f
C4984 VDD.n324 VSS 0.118f
C4985 VDD.n325 VSS 0.0281f
C4986 VDD.n326 VSS 0.0449f
C4987 VDD.t336 VSS 0.148f
C4988 VDD.n327 VSS 0.118f
C4989 VDD.n328 VSS 0.0281f
C4990 VDD.n329 VSS 0.0449f
C4991 VDD.t108 VSS 0.148f
C4992 VDD.t111 VSS 0.148f
C4993 VDD.n330 VSS 0.118f
C4994 VDD.n331 VSS 0.0281f
C4995 VDD.n332 VSS 0.0449f
C4996 VDD.t293 VSS 0.144f
C4997 VDD.n333 VSS 0.118f
C4998 VDD.n334 VSS 0.0269f
C4999 VDD.n335 VSS 0.0478f
C5000 VDD.t138 VSS 0.14f
C5001 VDD.n336 VSS 0.118f
C5002 VDD.n337 VSS 0.022f
C5003 VDD.n338 VSS 0.0478f
C5004 VDD.t285 VSS 0.148f
C5005 VDD.t106 VSS 0.148f
C5006 VDD.n339 VSS 0.118f
C5007 VDD.n340 VSS 0.0281f
C5008 VDD.n341 VSS 0.0449f
C5009 VDD.t110 VSS 0.148f
C5010 VDD.n342 VSS 0.118f
C5011 VDD.n343 VSS 0.0281f
C5012 VDD.n344 VSS 0.0449f
C5013 VDD.t292 VSS 0.125f
C5014 VDD.n345 VSS 0.118f
C5015 VDD.n346 VSS 0.0281f
C5016 VDD.n347 VSS 0.0449f
C5017 VDD.t137 VSS 0.14f
C5018 VDD.n348 VSS 0.118f
C5019 VDD.n349 VSS 0.0281f
C5020 VDD.n350 VSS 0.0449f
C5021 VDD.t284 VSS 0.148f
C5022 VDD.t300 VSS 0.148f
C5023 VDD.n351 VSS 0.118f
C5024 VDD.n352 VSS 0.0281f
C5025 VDD.n353 VSS 0.0449f
C5026 VDD.t107 VSS 0.155f
C5027 VDD.n354 VSS 0.118f
C5028 VDD.n355 VSS 0.0269f
C5029 VDD.n356 VSS 0.0478f
C5030 VDD.t303 VSS 0.129f
C5031 VDD.n357 VSS 0.118f
C5032 VDD.n358 VSS 0.022f
C5033 VDD.n359 VSS 0.0478f
C5034 VDD.t283 VSS 0.148f
C5035 VDD.n360 VSS 0.118f
C5036 VDD.n361 VSS 0.0281f
C5037 VDD.n362 VSS 0.0449f
C5038 VDD.t294 VSS 0.148f
C5039 VDD.t335 VSS 0.148f
C5040 VDD.n363 VSS 0.118f
C5041 VDD.n364 VSS 0.0281f
C5042 VDD.n365 VSS 0.0449f
C5043 VDD.t109 VSS 0.137f
C5044 VDD.n366 VSS 0.118f
C5045 VDD.n367 VSS 0.0281f
C5046 VDD.n368 VSS 0.0449f
C5047 VDD.t287 VSS 0.129f
C5048 VDD.n369 VSS 0.118f
C5049 VDD.n370 VSS 0.0281f
C5050 VDD.n371 VSS 0.0449f
C5051 VDD.t286 VSS 0.148f
C5052 VDD.n372 VSS 0.118f
C5053 VDD.n373 VSS 0.0281f
C5054 VDD.n374 VSS 0.0449f
C5055 VDD.t302 VSS 0.148f
C5056 VDD.t340 VSS 0.166f
C5057 VDD.n375 VSS 0.118f
C5058 VDD.n376 VSS 0.0269f
C5059 VDD.n377 VSS 0.0478f
C5060 VDD.t338 VSS 0.236f
C5061 VDD.n378 VSS 0.022f
C5062 VDD.n379 VSS 0.0478f
C5063 VDD.t298 VSS 0.148f
C5064 VDD.n380 VSS 0.118f
C5065 VDD.n381 VSS 0.0265f
C5066 VDD.n382 VSS 0.0371f
C5067 VDD.n383 VSS 0.0237f
C5068 VDD.n384 VSS 0.0236f
C5069 VDD.n385 VSS 0.00224f
C5070 VDD.t296 VSS 0.131f
C5071 VDD.n386 VSS 0.059f
C5072 VDD.n387 VSS 0.014f
C5073 VDD.n388 VSS 0.0108f
C5074 VDD.n389 VSS 0.00428f
C5075 VDD.t304 VSS 0.14f
C5076 VDD.n390 VSS 0.059f
C5077 VDD.n391 VSS 0.014f
C5078 VDD.n392 VSS 0.0191f
C5079 VDD.n393 VSS 0.023f
C5080 VDD.n394 VSS 0.00763f
C5081 VDD.t307 VSS 0.148f
C5082 VDD.n395 VSS 0.118f
C5083 VDD.n396 VSS 0.0274f
C5084 VDD.n397 VSS 0.00763f
C5085 VDD.n398 VSS 0.0205f
C5086 VDD.n399 VSS 0.0216f
C5087 VDD.t306 VSS 0.416f
C5088 VDD.n400 VSS 0.0324f
C5089 VDD.n401 VSS 0.0534f
C5090 VDD.n402 VSS 0.0268f
C5091 VDD.n403 VSS 0.25f
C5092 VDD.n404 VSS 1.08f
C5093 VDD.t126 VSS 0.00875f
C5094 VDD.n405 VSS 0.00459f
C5095 VDD.t141 VSS 0.00548f
C5096 VDD.t140 VSS 0.208f
C5097 VDD.t34 VSS 0.208f
C5098 VDD.n406 VSS 0.184f
C5099 VDD.n407 VSS 0.145f
C5100 VDD.n408 VSS 0.0922f
C5101 VDD.t125 VSS 0.167f
C5102 VDD.n409 VSS 0.0645f
C5103 VDD.t128 VSS 0.00875f
C5104 VDD.n410 VSS 0.00459f
C5105 VDD.t79 VSS 0.00548f
C5106 VDD.t78 VSS 0.208f
C5107 VDD.t245 VSS 0.208f
C5108 VDD.n411 VSS 0.184f
C5109 VDD.n412 VSS 0.145f
C5110 VDD.n413 VSS 0.0922f
C5111 VDD.t127 VSS 0.167f
C5112 VDD.n414 VSS 0.0923f
C5113 VDD.t313 VSS 0.00875f
C5114 VDD.n415 VSS 0.00459f
C5115 VDD.t38 VSS 0.00548f
C5116 VDD.t37 VSS 0.208f
C5117 VDD.t343 VSS 0.208f
C5118 VDD.n416 VSS 0.184f
C5119 VDD.n417 VSS 0.145f
C5120 VDD.n418 VSS 0.0922f
C5121 VDD.t312 VSS 0.167f
C5122 VDD.n419 VSS 0.0948f
C5123 VDD.t123 VSS 0.00875f
C5124 VDD.n420 VSS 0.00459f
C5125 VDD.t342 VSS 0.00459f
C5126 VDD.t45 VSS 0.00875f
C5127 VDD.n421 VSS 0.00459f
C5128 VDD.t244 VSS 0.00459f
C5129 VDD.t208 VSS 0.00875f
C5130 VDD.n422 VSS 0.00459f
C5131 VDD.t242 VSS 0.00548f
C5132 VDD.t241 VSS 0.208f
C5133 VDD.t221 VSS 0.208f
C5134 VDD.n423 VSS 0.184f
C5135 VDD.n424 VSS 0.145f
C5136 VDD.n425 VSS 0.0922f
C5137 VDD.t207 VSS 0.167f
C5138 VDD.n426 VSS 0.0723f
C5139 VDD.n427 VSS 0.0897f
C5140 VDD.t243 VSS 0.208f
C5141 VDD.t75 VSS 0.208f
C5142 VDD.n428 VSS 0.184f
C5143 VDD.n429 VSS 0.0574f
C5144 VDD.n430 VSS 0.0922f
C5145 VDD.t44 VSS 0.167f
C5146 VDD.n431 VSS 0.0726f
C5147 VDD.n432 VSS 0.0902f
C5148 VDD.t341 VSS 0.208f
C5149 VDD.t248 VSS 0.208f
C5150 VDD.n433 VSS 0.184f
C5151 VDD.n434 VSS 0.0574f
C5152 VDD.n435 VSS 0.0922f
C5153 VDD.t122 VSS 0.167f
C5154 VDD.n436 VSS 0.0654f
C5155 VDD.n437 VSS 0.123f
C5156 VDD.n438 VSS 0.0286f
C5157 VDD.n439 VSS 0.0257f
C5158 VDD.n440 VSS 0.0295f
C5159 VDD.n441 VSS 0.00945f
C5160 VDD.n442 VSS 0.0286f
C5161 VDD.n443 VSS 0.0333f
C5162 VDD.n444 VSS 0.00945f
C5163 VDD.n445 VSS 0.0175f
C5164 VDD.t102 VSS 0.00497f
C5165 VDD.n446 VSS 0.00497f
C5166 VDD.n447 VSS 0.0118f
C5167 VDD.n448 VSS 0.0126f
C5168 VDD.n449 VSS 0.00925f
C5169 VDD.n450 VSS 0.0197f
C5170 VDD.n451 VSS 0.143f
C5171 VDD.n452 VSS 0.0118f
C5172 VDD.t31 VSS 0.407f
C5173 VDD.n453 VSS 0.101f
C5174 VDD.n454 VSS 0.0462f
C5175 VDD.n455 VSS 0.0966f
C5176 VDD.n456 VSS 0.21f
C5177 VDD.n457 VSS 0.00925f
C5178 VDD.n458 VSS 0.0209f
C5179 VDD.t253 VSS 0.00497f
C5180 VDD.n459 VSS 0.00497f
C5181 VDD.n460 VSS 0.0125f
C5182 VDD.t327 VSS 0.00497f
C5183 VDD.n461 VSS 0.00497f
C5184 VDD.n462 VSS 0.012f
C5185 VDD.t47 VSS 0.00497f
C5186 VDD.n463 VSS 0.00497f
C5187 VDD.n464 VSS 0.0125f
C5188 VDD.t103 VSS 0.00497f
C5189 VDD.n465 VSS 0.00497f
C5190 VDD.n466 VSS 0.012f
C5191 VDD.t16 VSS 0.00497f
C5192 VDD.n467 VSS 0.00497f
C5193 VDD.n468 VSS 0.0125f
C5194 VDD.t25 VSS 0.00497f
C5195 VDD.n469 VSS 0.00497f
C5196 VDD.n470 VSS 0.012f
C5197 VDD.t33 VSS 0.00497f
C5198 VDD.n471 VSS 0.00497f
C5199 VDD.n472 VSS 0.0125f
C5200 VDD.t21 VSS 0.00497f
C5201 VDD.n473 VSS 0.00497f
C5202 VDD.n474 VSS 0.012f
C5203 VDD.t94 VSS 0.00497f
C5204 VDD.n475 VSS 0.00497f
C5205 VDD.n476 VSS 0.0125f
C5206 VDD.t69 VSS 0.00497f
C5207 VDD.n477 VSS 0.00497f
C5208 VDD.n478 VSS 0.012f
C5209 VDD.t1 VSS 0.00497f
C5210 VDD.n479 VSS 0.00497f
C5211 VDD.n480 VSS 0.0125f
C5212 VDD.t265 VSS 0.00497f
C5213 VDD.n481 VSS 0.00497f
C5214 VDD.n482 VSS 0.012f
C5215 VDD.t86 VSS 0.00497f
C5216 VDD.n483 VSS 0.00497f
C5217 VDD.n484 VSS 0.0125f
C5218 VDD.t266 VSS 0.00497f
C5219 VDD.n485 VSS 0.00497f
C5220 VDD.n486 VSS 0.012f
C5221 VDD.t83 VSS 0.00497f
C5222 VDD.n487 VSS 0.00497f
C5223 VDD.n488 VSS 0.0125f
C5224 VDD.n489 VSS 0.0122f
C5225 VDD.t322 VSS 0.00497f
C5226 VDD.n490 VSS 0.00497f
C5227 VDD.n491 VSS 0.0118f
C5228 VDD.t71 VSS 0.00497f
C5229 VDD.n492 VSS 0.00497f
C5230 VDD.n493 VSS 0.0118f
C5231 VDD.t269 VSS 0.00497f
C5232 VDD.n494 VSS 0.00497f
C5233 VDD.n495 VSS 0.0118f
C5234 VDD.t65 VSS 0.00497f
C5235 VDD.n496 VSS 0.00497f
C5236 VDD.n497 VSS 0.0118f
C5237 VDD.t63 VSS 0.00497f
C5238 VDD.n498 VSS 0.00497f
C5239 VDD.n499 VSS 0.0118f
C5240 VDD.t19 VSS 0.00497f
C5241 VDD.n500 VSS 0.00497f
C5242 VDD.n501 VSS 0.0118f
C5243 VDD.t80 VSS 0.483f
C5244 VDD.t89 VSS 0.483f
C5245 VDD.n502 VSS 0.495f
C5246 VDD.t46 VSS 0.441f
C5247 VDD.n503 VSS 0.495f
C5248 VDD.t332 VSS 0.00497f
C5249 VDD.n504 VSS 0.00497f
C5250 VDD.n505 VSS 0.0118f
C5251 VDD.n506 VSS 0.022f
C5252 VDD.t22 VSS 0.393f
C5253 VDD.n507 VSS 0.0252f
C5254 VDD.n508 VSS 0.177f
C5255 VDD.n509 VSS 0.00838f
C5256 VDD.n510 VSS 0.382f
C5257 VDD.n511 VSS 0.0144f
C5258 VDD.n512 VSS 0.0192f
C5259 VDD.n513 VSS 0.0105f
C5260 VDD.n514 VSS 0.0202f
C5261 VDD.n515 VSS 0.0233f
C5262 VDD.n516 VSS 0.0112f
C5263 VDD.n517 VSS 0.428f
C5264 VDD.n518 VSS 0.017f
C5265 VDD.n519 VSS 0.0148f
C5266 VDD.n520 VSS 0.395f
C5267 VDD.n521 VSS 0.0193f
C5268 VDD.t17 VSS 0.0882f
C5269 VDD.n522 VSS 0.118f
C5270 VDD.n523 VSS 0.00838f
C5271 VDD.n524 VSS 0.0105f
C5272 VDD.n525 VSS 0.02f
C5273 VDD.n526 VSS 0.0252f
C5274 VDD.n527 VSS 0.00599f
C5275 VDD.t12 VSS 0.0882f
C5276 VDD.n528 VSS 0.355f
C5277 VDD.n529 VSS 0.017f
C5278 VDD.n530 VSS 0.0151f
C5279 VDD.n531 VSS 0.344f
C5280 VDD.n532 VSS 0.0194f
C5281 VDD.n533 VSS 0.171f
C5282 VDD.n534 VSS 0.00825f
C5283 VDD.n535 VSS 0.0103f
C5284 VDD.n536 VSS 0.0103f
C5285 VDD.n537 VSS 0.0543f
C5286 VDD.n538 VSS 0.0887f
C5287 VDD.n539 VSS 0.0637f
C5288 VDD.n540 VSS 0.089f
C5289 VDD.n541 VSS 0.0577f
C5290 VDD.n542 VSS 0.0677f
C5291 VDD.n543 VSS 0.099f
C5292 VDD.n544 VSS 0.099f
C5293 VDD.n545 VSS 0.0747f
C5294 VDD.n546 VSS 0.0577f
C5295 VDD.n547 VSS 0.085f
C5296 VDD.n548 VSS 0.099f
C5297 VDD.n549 VSS 0.0956f
C5298 VDD.n550 VSS 0.0577f
C5299 VDD.n551 VSS 0.064f
C5300 VDD.n552 VSS 0.099f
C5301 VDD.n553 VSS 0.099f
C5302 VDD.n554 VSS 0.0783f
C5303 VDD.n555 VSS 0.0577f
C5304 VDD.n556 VSS 0.0813f
C5305 VDD.n557 VSS 0.099f
C5306 VDD.n558 VSS 0.099f
C5307 VDD.n559 VSS 0.061f
C5308 VDD.n560 VSS 0.0577f
C5309 VDD.n561 VSS 0.0986f
C5310 VDD.n562 VSS 0.099f
C5311 VDD.n563 VSS 0.082f
C5312 VDD.n564 VSS 0.0577f
C5313 VDD.n565 VSS 0.0705f
C5314 VDD.n566 VSS 0.0383f
C5315 VDD.n567 VSS 0.00766f
C5316 VDD.n568 VSS 0.107f
C5317 VDD.n569 VSS 0.00513f
C5318 VDD.n570 VSS 0.00165f
C5319 VDD.n571 VSS 0.00206f
C5320 VDD.n572 VSS 0.0668f
C5321 VDD.n573 VSS 0.187f
C5322 VDD.n574 VSS 0.0828f
C5323 VDD.n575 VSS 0.0357f
C5324 VDD.t29 VSS 0.0567f
C5325 VDD.n576 VSS 0.0135f
C5326 VDD.n577 VSS 0.0714f
C5327 VDD.n578 VSS 0.468f
C5328 VDD.n579 VSS 0.00955f
C5329 VDD.n580 VSS 0.0735f
C5330 VDD.n581 VSS 0.227f
C5331 VDD.n582 VSS 0.00612f
C5332 VDD.n583 VSS 0.426f
C5333 VDD.n584 VSS 0.0169f
C5334 VDD.n585 VSS 0.00612f
C5335 VDD.n586 VSS 0.0641f
C5336 VDD.n587 VSS 0.0183f
C5337 VDD.n588 VSS 0.0114f
C5338 VDD.n589 VSS 0.0356f
C5339 VDD.t82 VSS 0.888f
C5340 VDD.n590 VSS 0.0697f
C5341 VDD.n591 VSS 0.0579f
C5342 VDD.t98 VSS 0.483f
C5343 VDD.n592 VSS 0.495f
C5344 VDD.n593 VSS 0.0777f
C5345 VDD.t61 VSS 0.483f
C5346 VDD.n594 VSS 0.495f
C5347 VDD.n595 VSS 0.0657f
C5348 VDD.n596 VSS 0.0558f
C5349 VDD.t26 VSS 0.483f
C5350 VDD.n597 VSS 0.495f
C5351 VDD.n598 VSS 0.0854f
C5352 VDD.n599 VSS 0.0579f
C5353 VDD.t70 VSS 0.483f
C5354 VDD.t27 VSS 0.483f
C5355 VDD.n600 VSS 0.495f
C5356 VDD.n601 VSS 0.0582f
C5357 VDD.t10 VSS 0.483f
C5358 VDD.n602 VSS 0.495f
C5359 VDD.n603 VSS 0.0851f
C5360 VDD.n604 VSS 0.0558f
C5361 VDD.t28 VSS 0.483f
C5362 VDD.n605 VSS 0.495f
C5363 VDD.n606 VSS 0.0663f
C5364 VDD.t0 VSS 0.475f
C5365 VDD.n607 VSS 0.495f
C5366 VDD.n608 VSS 0.0771f
C5367 VDD.n609 VSS 0.0579f
C5368 VDD.t124 VSS 0.437f
C5369 VDD.n610 VSS 0.495f
C5370 VDD.n611 VSS 0.0743f
C5371 VDD.t68 VSS 0.483f
C5372 VDD.n612 VSS 0.495f
C5373 VDD.n613 VSS 0.0691f
C5374 VDD.n614 VSS 0.0558f
C5375 VDD.t5 VSS 0.483f
C5376 VDD.n615 VSS 0.495f
C5377 VDD.n616 VSS 0.0823f
C5378 VDD.t64 VSS 0.483f
C5379 VDD.n617 VSS 0.495f
C5380 VDD.n618 VSS 0.061f
C5381 VDD.n619 VSS 0.0579f
C5382 VDD.t54 VSS 0.483f
C5383 VDD.t20 VSS 0.483f
C5384 VDD.n620 VSS 0.495f
C5385 VDD.n621 VSS 0.0854f
C5386 VDD.n622 VSS 0.0558f
C5387 VDD.t30 VSS 0.483f
C5388 VDD.n623 VSS 0.495f
C5389 VDD.n624 VSS 0.0629f
C5390 VDD.t32 VSS 0.483f
C5391 VDD.n625 VSS 0.495f
C5392 VDD.n626 VSS 0.0805f
C5393 VDD.n627 VSS 0.0579f
C5394 VDD.t72 VSS 0.466f
C5395 VDD.n628 VSS 0.495f
C5396 VDD.n629 VSS 0.0709f
C5397 VDD.t8 VSS 0.445f
C5398 VDD.n630 VSS 0.495f
C5399 VDD.n631 VSS 0.0725f
C5400 VDD.n632 VSS 0.0558f
C5401 VDD.t2 VSS 0.483f
C5402 VDD.n633 VSS 0.495f
C5403 VDD.n634 VSS 0.0789f
C5404 VDD.t15 VSS 0.483f
C5405 VDD.n635 VSS 0.495f
C5406 VDD.n636 VSS 0.0644f
C5407 VDD.n637 VSS 0.0579f
C5408 VDD.t48 VSS 0.483f
C5409 VDD.n638 VSS 0.495f
C5410 VDD.n639 VSS 0.0854f
C5411 VDD.n640 VSS 0.0558f
C5412 VDD.n641 VSS 0.0595f
C5413 VDD.n642 VSS 0.0839f
C5414 VDD.n643 VSS 0.0579f
C5415 VDD.n644 VSS 0.0675f
C5416 VDD.n645 VSS 0.0759f
C5417 VDD.n646 VSS 0.0558f
C5418 VDD.n647 VSS 0.0755f
C5419 VDD.n648 VSS 0.0678f
C5420 VDD.n649 VSS 0.0545f
C5421 VDD.n650 VSS 0.0257f
C5422 VDD.n651 VSS 0.0112f
C5423 VDD.n652 VSS 0.00681f
C5424 VDD.t321 VSS 0.0121f
C5425 VDD.n653 VSS 0.116f
C5426 VDD.n654 VSS 0.0293f
C5427 VDD.n655 VSS 0.00353f
C5428 VDD.t18 VSS 0.00497f
C5429 VDD.n656 VSS 0.00497f
C5430 VDD.n657 VSS 0.012f
C5431 VDD.t81 VSS 0.00497f
C5432 VDD.n658 VSS 0.00497f
C5433 VDD.n659 VSS 0.012f
C5434 VDD.t9 VSS 0.00497f
C5435 VDD.n660 VSS 0.00497f
C5436 VDD.n661 VSS 0.012f
C5437 VDD.t51 VSS 0.00497f
C5438 VDD.n662 VSS 0.00497f
C5439 VDD.n663 VSS 0.012f
C5440 VDD.t256 VSS 0.00497f
C5441 VDD.n664 VSS 0.00497f
C5442 VDD.n665 VSS 0.012f
C5443 VDD.t11 VSS 0.00497f
C5444 VDD.n666 VSS 0.00497f
C5445 VDD.n667 VSS 0.012f
C5446 VDD.t62 VSS 0.00497f
C5447 VDD.n668 VSS 0.00497f
C5448 VDD.n669 VSS 0.012f
C5449 VDD.n670 VSS 0.0121f
C5450 VDD.n671 VSS 0.073f
C5451 VDD.n672 VSS 0.00433f
C5452 VDD.n673 VSS 0.00557f
C5453 VDD.n674 VSS 0.0122f
C5454 VDD.n675 VSS 0.00923f
C5455 VDD.n676 VSS 0.0202f
C5456 VDD.n677 VSS 0.0111f
C5457 VDD.n678 VSS 0.0356f
C5458 VDD.n679 VSS 0.0893f
C5459 VDD.n680 VSS 0.0935f
C5460 VDD.n681 VSS 0.0657f
C5461 VDD.n682 VSS 0.0558f
C5462 VDD.n683 VSS 0.0858f
C5463 VDD.n684 VSS 0.0935f
C5464 VDD.n685 VSS 0.0851f
C5465 VDD.n686 VSS 0.0558f
C5466 VDD.n687 VSS 0.0663f
C5467 VDD.n688 VSS 0.0935f
C5468 VDD.n689 VSS 0.0935f
C5469 VDD.n690 VSS 0.0691f
C5470 VDD.n691 VSS 0.0558f
C5471 VDD.n692 VSS 0.0823f
C5472 VDD.n693 VSS 0.0935f
C5473 VDD.n694 VSS 0.0885f
C5474 VDD.n695 VSS 0.0558f
C5475 VDD.n696 VSS 0.0629f
C5476 VDD.n697 VSS 0.0935f
C5477 VDD.n698 VSS 0.0935f
C5478 VDD.n699 VSS 0.0725f
C5479 VDD.n700 VSS 0.0558f
C5480 VDD.n701 VSS 0.0789f
C5481 VDD.n702 VSS 0.0935f
C5482 VDD.n703 VSS 0.0919f
C5483 VDD.n704 VSS 0.0558f
C5484 VDD.n705 VSS 0.0595f
C5485 VDD.n706 VSS 0.0935f
C5486 VDD.n707 VSS 0.0935f
C5487 VDD.n708 VSS 0.0759f
C5488 VDD.n709 VSS 0.0558f
C5489 VDD.n710 VSS 0.0755f
C5490 VDD.n711 VSS 0.0935f
C5491 VDD.n712 VSS 0.0839f
C5492 VDD.n713 VSS 0.0305f
C5493 VDD.t88 VSS 0.012f
C5494 VDD.n714 VSS 0.11f
C5495 VDD.n715 VSS 0.00696f
C5496 VDD.n716 VSS 0.0508f
C5497 VDD.n717 VSS 0.113f
C5498 VDD.n718 VSS 0.116f
C5499 VDD.t87 VSS 0.256f
C5500 VDD.n719 VSS 0.12f
C5501 VDD.n720 VSS 0.00945f
C5502 VDD.n721 VSS 0.13f
C5503 VDD.n722 VSS 0.00825f
C5504 VDD.n723 VSS 0.00825f
C5505 VDD.n724 VSS 0.295f
C5506 VDD.n725 VSS 0.359f
C5507 VDD.n726 VSS 0.18f
C5508 VDD.n727 VSS 0.0112f
C5509 VDD.n728 VSS 0.0117f
C5510 VDD.n729 VSS 0.0277f
C5511 VDD.n730 VSS 0.0527f
C5512 VDD.n731 VSS 0.0107f
C5513 VDD.n732 VSS 0.349f
C5514 VDD.n733 VSS 0.0208f
C5515 VDD.n734 VSS 0.154f
C5516 VDD.n735 VSS 0.00825f
C5517 VDD.n736 VSS 0.0103f
C5518 VDD.t101 VSS 0.101f
C5519 VDD.n737 VSS 0.273f
C5520 VDD.n738 VSS 0.0157f
C5521 VDD.n739 VSS 0.017f
C5522 VDD.n740 VSS 0.00478f
C5523 VDD.n741 VSS 0.0351f
C5524 VDD.n742 VSS 0.621f
C5525 VDD.n743 VSS 0.86f
C5526 VDD.n744 VSS 0.175f
C5527 VDD.n745 VSS 0.169f
C5528 VDD.n746 VSS 0.244f
C5529 VDD.n747 VSS 0.817f
C5530 VDD.n748 VSS 1.05f
C5531 VDD.n749 VSS 0.0174f
C5532 VDD.t236 VSS 0.0987f
C5533 VDD.n750 VSS 0.107f
C5534 VDD.t117 VSS 0.236f
C5535 VDD.n751 VSS 0.107f
C5536 VDD.t118 VSS 0.013f
C5537 VDD.n752 VSS 0.137f
C5538 VDD.n753 VSS 0.0648f
C5539 VDD.n754 VSS 0.0233f
C5540 VDD.t214 VSS 0.0987f
C5541 VDD.n755 VSS 0.107f
C5542 VDD.n756 VSS 0.0231f
C5543 VDD.n757 VSS 0.0222f
C5544 VDD.n758 VSS 0.0216f
C5545 VDD.n759 VSS 0.00677f
C5546 VDD.n760 VSS 0.00196f
C5547 VDD.n761 VSS 0.00353f
C5548 VDD.n762 VSS 0.0248f
C5549 VDD.n763 VSS 0.0235f
C5550 VDD.n764 VSS 0.0592f
C5551 VDD.n765 VSS 0.0664f
C5552 VDD.n766 VSS 0.0664f
C5553 VDD.n767 VSS 0.0398f
C5554 VDD.n768 VSS 0.0501f
C5555 OUT+.t73 VSS 0.0455f
C5556 OUT+.n0 VSS 0.0455f
C5557 OUT+.n1 VSS 0.124f
C5558 OUT+.t24 VSS 0.0455f
C5559 OUT+.n2 VSS 0.0455f
C5560 OUT+.n3 VSS 0.0909f
C5561 OUT+.n4 VSS 0.158f
C5562 OUT+.t62 VSS 0.0455f
C5563 OUT+.n5 VSS 0.0455f
C5564 OUT+.n6 VSS 0.124f
C5565 OUT+.t16 VSS 0.0455f
C5566 OUT+.n7 VSS 0.0455f
C5567 OUT+.n8 VSS 0.0909f
C5568 OUT+.n9 VSS 0.158f
C5569 OUT+.t77 VSS 0.0455f
C5570 OUT+.n10 VSS 0.0455f
C5571 OUT+.n11 VSS 0.124f
C5572 OUT+.t42 VSS 0.0455f
C5573 OUT+.n12 VSS 0.0455f
C5574 OUT+.n13 VSS 0.0909f
C5575 OUT+.n14 VSS 0.158f
C5576 OUT+.t68 VSS 0.0455f
C5577 OUT+.n15 VSS 0.0455f
C5578 OUT+.n16 VSS 0.124f
C5579 OUT+.t29 VSS 0.0455f
C5580 OUT+.n17 VSS 0.0455f
C5581 OUT+.n18 VSS 0.0909f
C5582 OUT+.n19 VSS 0.158f
C5583 OUT+.t53 VSS 0.0455f
C5584 OUT+.n20 VSS 0.0455f
C5585 OUT+.n21 VSS 0.124f
C5586 OUT+.t19 VSS 0.0455f
C5587 OUT+.n22 VSS 0.0455f
C5588 OUT+.n23 VSS 0.0909f
C5589 OUT+.n24 VSS 0.158f
C5590 OUT+.t74 VSS 0.0455f
C5591 OUT+.n25 VSS 0.0455f
C5592 OUT+.n26 VSS 0.124f
C5593 OUT+.t45 VSS 0.0455f
C5594 OUT+.n27 VSS 0.0455f
C5595 OUT+.n28 VSS 0.0909f
C5596 OUT+.n29 VSS 0.158f
C5597 OUT+.t49 VSS 0.0455f
C5598 OUT+.n30 VSS 0.0455f
C5599 OUT+.n31 VSS 0.124f
C5600 OUT+.t23 VSS 0.0455f
C5601 OUT+.n32 VSS 0.0455f
C5602 OUT+.n33 VSS 0.0909f
C5603 OUT+.n34 VSS 0.158f
C5604 OUT+.t1 VSS 0.0455f
C5605 OUT+.n35 VSS 0.0455f
C5606 OUT+.n36 VSS 0.124f
C5607 OUT+.t10 VSS 0.0455f
C5608 OUT+.n37 VSS 0.0455f
C5609 OUT+.n38 VSS 0.0909f
C5610 OUT+.n39 VSS 0.158f
C5611 OUT+.t50 VSS 0.0455f
C5612 OUT+.n40 VSS 0.0455f
C5613 OUT+.n41 VSS 0.124f
C5614 OUT+.t22 VSS 0.0455f
C5615 OUT+.n42 VSS 0.0455f
C5616 OUT+.n43 VSS 0.0909f
C5617 OUT+.n44 VSS 0.158f
C5618 OUT+.t58 VSS 0.0455f
C5619 OUT+.n45 VSS 0.0455f
C5620 OUT+.n46 VSS 0.124f
C5621 OUT+.t36 VSS 0.0455f
C5622 OUT+.n47 VSS 0.0455f
C5623 OUT+.n48 VSS 0.0909f
C5624 OUT+.n49 VSS 0.158f
C5625 OUT+.t0 VSS 0.0455f
C5626 OUT+.n50 VSS 0.0455f
C5627 OUT+.n51 VSS 0.124f
C5628 OUT+.t11 VSS 0.0455f
C5629 OUT+.n52 VSS 0.0455f
C5630 OUT+.n53 VSS 0.0909f
C5631 OUT+.n54 VSS 0.158f
C5632 OUT+.t7 VSS 0.0455f
C5633 OUT+.n55 VSS 0.0455f
C5634 OUT+.n56 VSS 0.124f
C5635 OUT+.t32 VSS 0.0455f
C5636 OUT+.n57 VSS 0.0455f
C5637 OUT+.n58 VSS 0.0909f
C5638 OUT+.n59 VSS 0.158f
C5639 OUT+.t5 VSS 0.0455f
C5640 OUT+.n60 VSS 0.0455f
C5641 OUT+.n61 VSS 0.124f
C5642 OUT+.t46 VSS 0.0455f
C5643 OUT+.n62 VSS 0.0455f
C5644 OUT+.n63 VSS 0.0909f
C5645 OUT+.n64 VSS 0.158f
C5646 OUT+.t75 VSS 0.0455f
C5647 OUT+.n65 VSS 0.0455f
C5648 OUT+.n66 VSS 0.124f
C5649 OUT+.t44 VSS 0.0455f
C5650 OUT+.n67 VSS 0.0455f
C5651 OUT+.n68 VSS 0.0909f
C5652 OUT+.n69 VSS 0.158f
C5653 OUT+.t54 VSS 0.0455f
C5654 OUT+.n70 VSS 0.0455f
C5655 OUT+.n71 VSS 0.124f
C5656 OUT+.t18 VSS 0.0455f
C5657 OUT+.n72 VSS 0.0455f
C5658 OUT+.n73 VSS 0.0909f
C5659 OUT+.n74 VSS 0.158f
C5660 OUT+.t8 VSS 0.0455f
C5661 OUT+.n75 VSS 0.0455f
C5662 OUT+.n76 VSS 0.124f
C5663 OUT+.t31 VSS 0.0455f
C5664 OUT+.n77 VSS 0.0455f
C5665 OUT+.n78 VSS 0.0909f
C5666 OUT+.n79 VSS 0.158f
C5667 OUT+.t55 VSS 0.0455f
C5668 OUT+.n80 VSS 0.0455f
C5669 OUT+.n81 VSS 0.124f
C5670 OUT+.t39 VSS 0.0455f
C5671 OUT+.n82 VSS 0.0455f
C5672 OUT+.n83 VSS 0.0909f
C5673 OUT+.n84 VSS 0.158f
C5674 OUT+.t65 VSS 0.0455f
C5675 OUT+.n85 VSS 0.0455f
C5676 OUT+.n86 VSS 0.124f
C5677 OUT+.t13 VSS 0.0455f
C5678 OUT+.n87 VSS 0.0455f
C5679 OUT+.n88 VSS 0.0909f
C5680 OUT+.n89 VSS 0.158f
C5681 OUT+.t71 VSS 0.0455f
C5682 OUT+.n90 VSS 0.0455f
C5683 OUT+.n91 VSS 0.124f
C5684 OUT+.t26 VSS 0.0455f
C5685 OUT+.n92 VSS 0.0455f
C5686 OUT+.n93 VSS 0.0909f
C5687 OUT+.n94 VSS 0.158f
C5688 OUT+.t56 VSS 0.0455f
C5689 OUT+.n95 VSS 0.0455f
C5690 OUT+.n96 VSS 0.124f
C5691 OUT+.t38 VSS 0.0455f
C5692 OUT+.n97 VSS 0.0455f
C5693 OUT+.n98 VSS 0.0909f
C5694 OUT+.n99 VSS 0.198f
C5695 OUT+.n100 VSS 0.291f
C5696 OUT+.n101 VSS 0.204f
C5697 OUT+.n102 VSS 0.204f
C5698 OUT+.n103 VSS 0.204f
C5699 OUT+.n104 VSS 0.204f
C5700 OUT+.n105 VSS 0.204f
C5701 OUT+.n106 VSS 0.204f
C5702 OUT+.n107 VSS 0.204f
C5703 OUT+.n108 VSS 0.204f
C5704 OUT+.n109 VSS 0.204f
C5705 OUT+.n110 VSS 0.204f
C5706 OUT+.n111 VSS 0.204f
C5707 OUT+.n112 VSS 0.204f
C5708 OUT+.n113 VSS 0.204f
C5709 OUT+.n114 VSS 0.204f
C5710 OUT+.n115 VSS 0.204f
C5711 OUT+.n116 VSS 0.204f
C5712 OUT+.n117 VSS 0.204f
C5713 OUT+.n118 VSS 0.219f
C5714 SEL_L.t3 VSS 0.0118f
C5715 SEL_L.t10 VSS 0.0118f
C5716 SEL_L.t40 VSS 0.0118f
C5717 SEL_L.t78 VSS 0.0139f
C5718 SEL_L.t45 VSS 0.0118f
C5719 SEL_L.t84 VSS 0.0139f
C5720 SEL_L.t39 VSS 0.0118f
C5721 SEL_L.t76 VSS 0.0139f
C5722 SEL_L.t65 VSS 0.0118f
C5723 SEL_L.t9 VSS 0.0139f
C5724 SEL_L.t68 VSS 0.0118f
C5725 SEL_L.t100 VSS 0.0158f
C5726 SEL_L.n0 VSS 0.0178f
C5727 SEL_L.n1 VSS 0.0192f
C5728 SEL_L.n2 VSS 0.0192f
C5729 SEL_L.n3 VSS 0.0192f
C5730 SEL_L.n4 VSS 0.0192f
C5731 SEL_L.n5 VSS 0.012f
C5732 SEL_L.n6 VSS 0.0155f
C5733 SEL_L.t6 VSS 0.0118f
C5734 SEL_L.t29 VSS 0.015f
C5735 SEL_L.t31 VSS 0.0124f
C5736 SEL_L.n7 VSS 0.0177f
C5737 SEL_L.t27 VSS 0.0124f
C5738 SEL_L.n8 VSS 0.0113f
C5739 SEL_L.t53 VSS 0.0124f
C5740 SEL_L.n9 VSS 0.0113f
C5741 SEL_L.t59 VSS 0.0124f
C5742 SEL_L.n10 VSS 0.0113f
C5743 SEL_L.t86 VSS 0.0124f
C5744 SEL_L.n11 VSS 0.0113f
C5745 SEL_L.t89 VSS 0.0124f
C5746 SEL_L.n12 VSS 0.0113f
C5747 SEL_L.t16 VSS 0.0124f
C5748 SEL_L.n13 VSS 0.0113f
C5749 SEL_L.t43 VSS 0.0124f
C5750 SEL_L.n14 VSS 0.0113f
C5751 SEL_L.t46 VSS 0.0124f
C5752 SEL_L.n15 VSS 0.0113f
C5753 SEL_L.t71 VSS 0.0124f
C5754 SEL_L.n16 VSS 0.0113f
C5755 SEL_L.t74 VSS 0.0124f
C5756 SEL_L.n17 VSS 0.0113f
C5757 SEL_L.t5 VSS 0.0124f
C5758 SEL_L.n18 VSS 0.0113f
C5759 SEL_L.t36 VSS 0.0124f
C5760 SEL_L.n19 VSS 0.0113f
C5761 SEL_L.t23 VSS 0.0124f
C5762 SEL_L.n20 VSS 0.0113f
C5763 SEL_L.t85 VSS 0.0124f
C5764 SEL_L.n21 VSS 0.0113f
C5765 SEL_L.t79 VSS 0.0124f
C5766 SEL_L.n22 VSS 0.0113f
C5767 SEL_L.t51 VSS 0.0124f
C5768 SEL_L.n23 VSS 0.0113f
C5769 SEL_L.t25 VSS 0.0124f
C5770 SEL_L.n24 VSS 0.0113f
C5771 SEL_L.t19 VSS 0.0124f
C5772 SEL_L.n25 VSS 0.0113f
C5773 SEL_L.t91 VSS 0.0124f
C5774 SEL_L.n26 VSS 0.0113f
C5775 SEL_L.t83 VSS 0.0124f
C5776 SEL_L.n27 VSS 0.0113f
C5777 SEL_L.t57 VSS 0.0124f
C5778 SEL_L.n28 VSS 0.0113f
C5779 SEL_L.t30 VSS 0.0124f
C5780 SEL_L.n29 VSS 0.0113f
C5781 SEL_L.t24 VSS 0.0124f
C5782 SEL_L.n30 VSS 0.0113f
C5783 SEL_L.t93 VSS 0.0124f
C5784 SEL_L.n31 VSS 0.0113f
C5785 SEL_L.t90 VSS 0.0124f
C5786 SEL_L.n32 VSS 0.0113f
C5787 SEL_L.t96 VSS 0.0124f
C5788 SEL_L.n33 VSS 0.0113f
C5789 SEL_L.t63 VSS 0.0124f
C5790 SEL_L.n34 VSS 0.0113f
C5791 SEL_L.t61 VSS 0.0124f
C5792 SEL_L.n35 VSS 0.0113f
C5793 SEL_L.t34 VSS 0.0124f
C5794 SEL_L.n36 VSS 0.0113f
C5795 SEL_L.t32 VSS 0.0124f
C5796 SEL_L.n37 VSS 0.0113f
C5797 SEL_L.t101 VSS 0.0124f
C5798 SEL_L.n38 VSS 0.0113f
C5799 SEL_L.t2 VSS 0.0124f
C5800 SEL_L.n39 VSS 0.0113f
C5801 SEL_L.t102 VSS 0.0124f
C5802 SEL_L.n40 VSS 0.0113f
C5803 SEL_L.t70 VSS 0.0124f
C5804 SEL_L.n41 VSS 0.0113f
C5805 SEL_L.t67 VSS 0.0124f
C5806 SEL_L.n42 VSS 0.0113f
C5807 SEL_L.t42 VSS 0.0124f
C5808 SEL_L.n43 VSS 0.0113f
C5809 SEL_L.t11 VSS 0.0124f
C5810 SEL_L.n44 VSS 0.0118f
C5811 SEL_L.n45 VSS 0.0276f
C5812 SEL_L.n46 VSS 0.107f
C5813 SEL_L.n47 VSS 0.155f
C5814 SEL_L.t20 VSS 0.0118f
C5815 SEL_L.t26 VSS 0.0118f
C5816 SEL_L.t52 VSS 0.0118f
C5817 SEL_L.t94 VSS 0.0139f
C5818 SEL_L.t58 VSS 0.0118f
C5819 SEL_L.t98 VSS 0.0139f
C5820 SEL_L.t50 VSS 0.0118f
C5821 SEL_L.t92 VSS 0.0139f
C5822 SEL_L.t77 VSS 0.0118f
C5823 SEL_L.t22 VSS 0.0139f
C5824 SEL_L.t82 VSS 0.0118f
C5825 SEL_L.t12 VSS 0.0158f
C5826 SEL_L.n48 VSS 0.0178f
C5827 SEL_L.n49 VSS 0.0192f
C5828 SEL_L.n50 VSS 0.0192f
C5829 SEL_L.n51 VSS 0.0192f
C5830 SEL_L.n52 VSS 0.0192f
C5831 SEL_L.n53 VSS 0.012f
C5832 SEL_L.n54 VSS 0.0155f
C5833 SEL_L.t21 VSS 0.0118f
C5834 SEL_L.t56 VSS 0.015f
C5835 SEL_L.t60 VSS 0.0124f
C5836 SEL_L.n55 VSS 0.0177f
C5837 SEL_L.t54 VSS 0.0124f
C5838 SEL_L.n56 VSS 0.0113f
C5839 SEL_L.t80 VSS 0.0124f
C5840 SEL_L.n57 VSS 0.0113f
C5841 SEL_L.t87 VSS 0.0124f
C5842 SEL_L.n58 VSS 0.0113f
C5843 SEL_L.t14 VSS 0.0124f
C5844 SEL_L.n59 VSS 0.0113f
C5845 SEL_L.t17 VSS 0.0124f
C5846 SEL_L.n60 VSS 0.0113f
C5847 SEL_L.t48 VSS 0.0124f
C5848 SEL_L.n61 VSS 0.0113f
C5849 SEL_L.t69 VSS 0.0124f
C5850 SEL_L.n62 VSS 0.0113f
C5851 SEL_L.t72 VSS 0.0124f
C5852 SEL_L.n63 VSS 0.0113f
C5853 SEL_L.t0 VSS 0.0124f
C5854 SEL_L.n64 VSS 0.0113f
C5855 SEL_L.t7 VSS 0.0124f
C5856 SEL_L.n65 VSS 0.0113f
C5857 SEL_L.t37 VSS 0.0124f
C5858 SEL_L.n66 VSS 0.0113f
C5859 SEL_L.t62 VSS 0.0124f
C5860 SEL_L.n67 VSS 0.0113f
C5861 SEL_L.t49 VSS 0.0124f
C5862 SEL_L.n68 VSS 0.0113f
C5863 SEL_L.t99 VSS 0.0124f
C5864 SEL_L.n69 VSS 0.0113f
C5865 SEL_L.t95 VSS 0.0124f
C5866 SEL_L.n70 VSS 0.0113f
C5867 SEL_L.t64 VSS 0.0124f
C5868 SEL_L.n71 VSS 0.0113f
C5869 SEL_L.t38 VSS 0.0124f
C5870 SEL_L.n72 VSS 0.0113f
C5871 SEL_L.t33 VSS 0.0124f
C5872 SEL_L.n73 VSS 0.0113f
C5873 SEL_L.t1 VSS 0.0124f
C5874 SEL_L.n74 VSS 0.0113f
C5875 SEL_L.t97 VSS 0.0124f
C5876 SEL_L.n75 VSS 0.0113f
C5877 SEL_L.t66 VSS 0.0124f
C5878 SEL_L.n76 VSS 0.0113f
C5879 SEL_L.t41 VSS 0.0124f
C5880 SEL_L.n77 VSS 0.0113f
C5881 SEL_L.t35 VSS 0.0124f
C5882 SEL_L.n78 VSS 0.0113f
C5883 SEL_L.t4 VSS 0.0124f
C5884 SEL_L.n79 VSS 0.0113f
C5885 SEL_L.t103 VSS 0.0124f
C5886 SEL_L.n80 VSS 0.0113f
C5887 SEL_L.t8 VSS 0.0124f
C5888 SEL_L.n81 VSS 0.0113f
C5889 SEL_L.t75 VSS 0.0124f
C5890 SEL_L.n82 VSS 0.0113f
C5891 SEL_L.t73 VSS 0.0124f
C5892 SEL_L.n83 VSS 0.0113f
C5893 SEL_L.t47 VSS 0.0124f
C5894 SEL_L.n84 VSS 0.0113f
C5895 SEL_L.t44 VSS 0.0124f
C5896 SEL_L.n85 VSS 0.0113f
C5897 SEL_L.t13 VSS 0.0124f
C5898 SEL_L.n86 VSS 0.0113f
C5899 SEL_L.t18 VSS 0.0124f
C5900 SEL_L.n87 VSS 0.0113f
C5901 SEL_L.t15 VSS 0.0124f
C5902 SEL_L.n88 VSS 0.0113f
C5903 SEL_L.t88 VSS 0.0124f
C5904 SEL_L.n89 VSS 0.0113f
C5905 SEL_L.t81 VSS 0.0124f
C5906 SEL_L.n90 VSS 0.0113f
C5907 SEL_L.t55 VSS 0.0124f
C5908 SEL_L.n91 VSS 0.0113f
C5909 SEL_L.t28 VSS 0.0124f
C5910 SEL_L.n92 VSS 0.0118f
C5911 SEL_L.n93 VSS 0.0255f
C5912 SEL_L.n94 VSS 0.109f
.ends

