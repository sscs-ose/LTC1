magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1149 1019 1149
<< metal1 >>
rect -19 143 19 149
rect -19 -143 -13 143
rect 13 -143 19 143
rect -19 -149 19 -143
<< via1 >>
rect -13 -143 13 143
<< metal2 >>
rect -19 143 19 149
rect -19 -143 -13 143
rect 13 -143 19 143
rect -19 -149 19 -143
<< end >>
