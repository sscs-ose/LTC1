magic
tech gf180mcuC
magscale 1 10
timestamp 1692617267
<< nwell >>
rect -986 -1586 986 1586
<< pmos >>
rect -812 830 -700 1456
rect -596 830 -484 1456
rect -380 830 -268 1456
rect -164 830 -52 1456
rect 52 830 164 1456
rect 268 830 380 1456
rect 484 830 596 1456
rect 700 830 812 1456
rect -812 68 -700 694
rect -596 68 -484 694
rect -380 68 -268 694
rect -164 68 -52 694
rect 52 68 164 694
rect 268 68 380 694
rect 484 68 596 694
rect 700 68 812 694
rect -812 -694 -700 -68
rect -596 -694 -484 -68
rect -380 -694 -268 -68
rect -164 -694 -52 -68
rect 52 -694 164 -68
rect 268 -694 380 -68
rect 484 -694 596 -68
rect 700 -694 812 -68
rect -812 -1456 -700 -830
rect -596 -1456 -484 -830
rect -380 -1456 -268 -830
rect -164 -1456 -52 -830
rect 52 -1456 164 -830
rect 268 -1456 380 -830
rect 484 -1456 596 -830
rect 700 -1456 812 -830
<< pdiff >>
rect -900 1443 -812 1456
rect -900 843 -887 1443
rect -841 843 -812 1443
rect -900 830 -812 843
rect -700 1443 -596 1456
rect -700 843 -671 1443
rect -625 843 -596 1443
rect -700 830 -596 843
rect -484 1443 -380 1456
rect -484 843 -455 1443
rect -409 843 -380 1443
rect -484 830 -380 843
rect -268 1443 -164 1456
rect -268 843 -239 1443
rect -193 843 -164 1443
rect -268 830 -164 843
rect -52 1443 52 1456
rect -52 843 -23 1443
rect 23 843 52 1443
rect -52 830 52 843
rect 164 1443 268 1456
rect 164 843 193 1443
rect 239 843 268 1443
rect 164 830 268 843
rect 380 1443 484 1456
rect 380 843 409 1443
rect 455 843 484 1443
rect 380 830 484 843
rect 596 1443 700 1456
rect 596 843 625 1443
rect 671 843 700 1443
rect 596 830 700 843
rect 812 1443 900 1456
rect 812 843 841 1443
rect 887 843 900 1443
rect 812 830 900 843
rect -900 681 -812 694
rect -900 81 -887 681
rect -841 81 -812 681
rect -900 68 -812 81
rect -700 681 -596 694
rect -700 81 -671 681
rect -625 81 -596 681
rect -700 68 -596 81
rect -484 681 -380 694
rect -484 81 -455 681
rect -409 81 -380 681
rect -484 68 -380 81
rect -268 681 -164 694
rect -268 81 -239 681
rect -193 81 -164 681
rect -268 68 -164 81
rect -52 681 52 694
rect -52 81 -23 681
rect 23 81 52 681
rect -52 68 52 81
rect 164 681 268 694
rect 164 81 193 681
rect 239 81 268 681
rect 164 68 268 81
rect 380 681 484 694
rect 380 81 409 681
rect 455 81 484 681
rect 380 68 484 81
rect 596 681 700 694
rect 596 81 625 681
rect 671 81 700 681
rect 596 68 700 81
rect 812 681 900 694
rect 812 81 841 681
rect 887 81 900 681
rect 812 68 900 81
rect -900 -81 -812 -68
rect -900 -681 -887 -81
rect -841 -681 -812 -81
rect -900 -694 -812 -681
rect -700 -81 -596 -68
rect -700 -681 -671 -81
rect -625 -681 -596 -81
rect -700 -694 -596 -681
rect -484 -81 -380 -68
rect -484 -681 -455 -81
rect -409 -681 -380 -81
rect -484 -694 -380 -681
rect -268 -81 -164 -68
rect -268 -681 -239 -81
rect -193 -681 -164 -81
rect -268 -694 -164 -681
rect -52 -81 52 -68
rect -52 -681 -23 -81
rect 23 -681 52 -81
rect -52 -694 52 -681
rect 164 -81 268 -68
rect 164 -681 193 -81
rect 239 -681 268 -81
rect 164 -694 268 -681
rect 380 -81 484 -68
rect 380 -681 409 -81
rect 455 -681 484 -81
rect 380 -694 484 -681
rect 596 -81 700 -68
rect 596 -681 625 -81
rect 671 -681 700 -81
rect 596 -694 700 -681
rect 812 -81 900 -68
rect 812 -681 841 -81
rect 887 -681 900 -81
rect 812 -694 900 -681
rect -900 -843 -812 -830
rect -900 -1443 -887 -843
rect -841 -1443 -812 -843
rect -900 -1456 -812 -1443
rect -700 -843 -596 -830
rect -700 -1443 -671 -843
rect -625 -1443 -596 -843
rect -700 -1456 -596 -1443
rect -484 -843 -380 -830
rect -484 -1443 -455 -843
rect -409 -1443 -380 -843
rect -484 -1456 -380 -1443
rect -268 -843 -164 -830
rect -268 -1443 -239 -843
rect -193 -1443 -164 -843
rect -268 -1456 -164 -1443
rect -52 -843 52 -830
rect -52 -1443 -23 -843
rect 23 -1443 52 -843
rect -52 -1456 52 -1443
rect 164 -843 268 -830
rect 164 -1443 193 -843
rect 239 -1443 268 -843
rect 164 -1456 268 -1443
rect 380 -843 484 -830
rect 380 -1443 409 -843
rect 455 -1443 484 -843
rect 380 -1456 484 -1443
rect 596 -843 700 -830
rect 596 -1443 625 -843
rect 671 -1443 700 -843
rect 596 -1456 700 -1443
rect 812 -843 900 -830
rect 812 -1443 841 -843
rect 887 -1443 900 -843
rect 812 -1456 900 -1443
<< pdiffc >>
rect -887 843 -841 1443
rect -671 843 -625 1443
rect -455 843 -409 1443
rect -239 843 -193 1443
rect -23 843 23 1443
rect 193 843 239 1443
rect 409 843 455 1443
rect 625 843 671 1443
rect 841 843 887 1443
rect -887 81 -841 681
rect -671 81 -625 681
rect -455 81 -409 681
rect -239 81 -193 681
rect -23 81 23 681
rect 193 81 239 681
rect 409 81 455 681
rect 625 81 671 681
rect 841 81 887 681
rect -887 -681 -841 -81
rect -671 -681 -625 -81
rect -455 -681 -409 -81
rect -239 -681 -193 -81
rect -23 -681 23 -81
rect 193 -681 239 -81
rect 409 -681 455 -81
rect 625 -681 671 -81
rect 841 -681 887 -81
rect -887 -1443 -841 -843
rect -671 -1443 -625 -843
rect -455 -1443 -409 -843
rect -239 -1443 -193 -843
rect -23 -1443 23 -843
rect 193 -1443 239 -843
rect 409 -1443 455 -843
rect 625 -1443 671 -843
rect 841 -1443 887 -843
<< polysilicon >>
rect -812 1456 -700 1500
rect -596 1456 -484 1500
rect -380 1456 -268 1500
rect -164 1456 -52 1500
rect 52 1456 164 1500
rect 268 1456 380 1500
rect 484 1456 596 1500
rect 700 1456 812 1500
rect -812 786 -700 830
rect -596 786 -484 830
rect -380 786 -268 830
rect -164 786 -52 830
rect 52 786 164 830
rect 268 786 380 830
rect 484 786 596 830
rect 700 786 812 830
rect -812 694 -700 738
rect -596 694 -484 738
rect -380 694 -268 738
rect -164 694 -52 738
rect 52 694 164 738
rect 268 694 380 738
rect 484 694 596 738
rect 700 694 812 738
rect -812 24 -700 68
rect -596 24 -484 68
rect -380 24 -268 68
rect -164 24 -52 68
rect 52 24 164 68
rect 268 24 380 68
rect 484 24 596 68
rect 700 24 812 68
rect -812 -68 -700 -24
rect -596 -68 -484 -24
rect -380 -68 -268 -24
rect -164 -68 -52 -24
rect 52 -68 164 -24
rect 268 -68 380 -24
rect 484 -68 596 -24
rect 700 -68 812 -24
rect -812 -738 -700 -694
rect -596 -738 -484 -694
rect -380 -738 -268 -694
rect -164 -738 -52 -694
rect 52 -738 164 -694
rect 268 -738 380 -694
rect 484 -738 596 -694
rect 700 -738 812 -694
rect -812 -830 -700 -786
rect -596 -830 -484 -786
rect -380 -830 -268 -786
rect -164 -830 -52 -786
rect 52 -830 164 -786
rect 268 -830 380 -786
rect 484 -830 596 -786
rect 700 -830 812 -786
rect -812 -1500 -700 -1456
rect -596 -1500 -484 -1456
rect -380 -1500 -268 -1456
rect -164 -1500 -52 -1456
rect 52 -1500 164 -1456
rect 268 -1500 380 -1456
rect 484 -1500 596 -1456
rect 700 -1500 812 -1456
<< metal1 >>
rect -887 1443 -841 1454
rect -887 832 -841 843
rect -671 1443 -625 1454
rect -671 832 -625 843
rect -455 1443 -409 1454
rect -455 832 -409 843
rect -239 1443 -193 1454
rect -239 832 -193 843
rect -23 1443 23 1454
rect -23 832 23 843
rect 193 1443 239 1454
rect 193 832 239 843
rect 409 1443 455 1454
rect 409 832 455 843
rect 625 1443 671 1454
rect 625 832 671 843
rect 841 1443 887 1454
rect 841 832 887 843
rect -887 681 -841 692
rect -887 70 -841 81
rect -671 681 -625 692
rect -671 70 -625 81
rect -455 681 -409 692
rect -455 70 -409 81
rect -239 681 -193 692
rect -239 70 -193 81
rect -23 681 23 692
rect -23 70 23 81
rect 193 681 239 692
rect 193 70 239 81
rect 409 681 455 692
rect 409 70 455 81
rect 625 681 671 692
rect 625 70 671 81
rect 841 681 887 692
rect 841 70 887 81
rect -887 -81 -841 -70
rect -887 -692 -841 -681
rect -671 -81 -625 -70
rect -671 -692 -625 -681
rect -455 -81 -409 -70
rect -455 -692 -409 -681
rect -239 -81 -193 -70
rect -239 -692 -193 -681
rect -23 -81 23 -70
rect -23 -692 23 -681
rect 193 -81 239 -70
rect 193 -692 239 -681
rect 409 -81 455 -70
rect 409 -692 455 -681
rect 625 -81 671 -70
rect 625 -692 671 -681
rect 841 -81 887 -70
rect 841 -692 887 -681
rect -887 -843 -841 -832
rect -887 -1454 -841 -1443
rect -671 -843 -625 -832
rect -671 -1454 -625 -1443
rect -455 -843 -409 -832
rect -455 -1454 -409 -1443
rect -239 -843 -193 -832
rect -239 -1454 -193 -1443
rect -23 -843 23 -832
rect -23 -1454 23 -1443
rect 193 -843 239 -832
rect 193 -1454 239 -1443
rect 409 -843 455 -832
rect 409 -1454 455 -1443
rect 625 -843 671 -832
rect 625 -1454 671 -1443
rect 841 -843 887 -832
rect 841 -1454 887 -1443
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 3.125 l 0.56 m 4 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
