magic
tech gf180mcuC
magscale 1 10
timestamp 1700416336
<< pwell >>
rect 114165 1654 114402 1661
<< psubdiff >>
rect 113240 2838 116409 2856
rect 113240 2777 113387 2838
rect 113450 2777 113517 2838
rect 113580 2777 113647 2838
rect 113710 2777 113777 2838
rect 113840 2777 113907 2838
rect 113970 2777 114037 2838
rect 114100 2777 114167 2838
rect 114230 2777 114297 2838
rect 114360 2777 114427 2838
rect 114490 2777 114557 2838
rect 114620 2777 114687 2838
rect 114750 2777 114817 2838
rect 114880 2777 114947 2838
rect 115010 2777 115077 2838
rect 115140 2777 115207 2838
rect 115270 2777 115337 2838
rect 115400 2777 115467 2838
rect 115530 2777 115597 2838
rect 115660 2777 115727 2838
rect 115790 2777 115857 2838
rect 115920 2777 115987 2838
rect 116050 2777 116117 2838
rect 116180 2793 116409 2838
rect 116180 2777 116329 2793
rect 113240 2775 116329 2777
rect 113240 2714 113258 2775
rect 113321 2758 116329 2775
rect 113321 2714 113338 2758
rect 113240 2645 113338 2714
rect 113240 2584 113258 2645
rect 113321 2584 113338 2645
rect 113240 2515 113338 2584
rect 113240 2454 113258 2515
rect 113321 2454 113338 2515
rect 113240 2385 113338 2454
rect 113240 2324 113258 2385
rect 113321 2324 113338 2385
rect 113240 2255 113338 2324
rect 113240 2194 113258 2255
rect 113321 2194 113338 2255
rect 113240 2125 113338 2194
rect 113240 2064 113258 2125
rect 113321 2064 113338 2125
rect 113240 1995 113338 2064
rect 113240 1934 113258 1995
rect 113321 1934 113338 1995
rect 113240 1865 113338 1934
rect 113240 1804 113258 1865
rect 113321 1804 113338 1865
rect 116311 2732 116329 2758
rect 116392 2732 116409 2793
rect 116311 2663 116409 2732
rect 116311 2602 116329 2663
rect 116392 2602 116409 2663
rect 116311 2533 116409 2602
rect 116311 2472 116329 2533
rect 116392 2472 116409 2533
rect 116311 2403 116409 2472
rect 116311 2342 116329 2403
rect 116392 2342 116409 2403
rect 116311 2273 116409 2342
rect 116311 2212 116329 2273
rect 116392 2212 116409 2273
rect 116311 2143 116409 2212
rect 116311 2082 116329 2143
rect 116392 2082 116409 2143
rect 116311 2013 116409 2082
rect 116311 1952 116329 2013
rect 116392 1952 116409 2013
rect 116311 1883 116409 1952
rect 113240 1735 113338 1804
rect 113240 1674 113258 1735
rect 113321 1674 113338 1735
rect 113240 1605 113338 1674
rect 113240 1544 113258 1605
rect 113321 1544 113338 1605
rect 116311 1822 116329 1883
rect 116392 1822 116409 1883
rect 116311 1753 116409 1822
rect 116311 1692 116329 1753
rect 116392 1692 116409 1753
rect 116311 1623 116409 1692
rect 116311 1562 116329 1623
rect 116392 1562 116409 1623
rect 113240 1475 113338 1544
rect 113240 1414 113258 1475
rect 113321 1414 113338 1475
rect 113240 1345 113338 1414
rect 113240 1284 113258 1345
rect 113321 1284 113338 1345
rect 113240 1215 113338 1284
rect 113240 1154 113258 1215
rect 113321 1154 113338 1215
rect 113240 1085 113338 1154
rect 113240 1024 113258 1085
rect 113321 1024 113338 1085
rect 113240 955 113338 1024
rect 113240 894 113258 955
rect 113321 894 113338 955
rect 113240 879 113338 894
rect 116311 1493 116409 1562
rect 116311 1432 116329 1493
rect 116392 1432 116409 1493
rect 116311 1363 116409 1432
rect 116311 1302 116329 1363
rect 116392 1302 116409 1363
rect 116311 1233 116409 1302
rect 116311 1172 116329 1233
rect 116392 1172 116409 1233
rect 116311 1103 116409 1172
rect 116311 1042 116329 1103
rect 116392 1042 116409 1103
rect 116311 973 116409 1042
rect 116311 912 116329 973
rect 116392 912 116409 973
rect 116311 879 116409 912
rect 113240 859 116409 879
rect 113240 798 113371 859
rect 113434 798 113501 859
rect 113564 798 113631 859
rect 113694 798 113761 859
rect 113824 798 113891 859
rect 113954 798 114021 859
rect 114084 798 114151 859
rect 114214 798 114281 859
rect 114344 798 114411 859
rect 114474 798 114541 859
rect 114604 798 114671 859
rect 114734 798 114801 859
rect 114864 798 114931 859
rect 114994 798 115061 859
rect 115124 798 115191 859
rect 115254 798 115321 859
rect 115384 798 115451 859
rect 115514 798 115581 859
rect 115644 798 115711 859
rect 115774 798 115841 859
rect 115904 798 115971 859
rect 116034 798 116101 859
rect 116164 798 116231 859
rect 116294 798 116409 859
rect 113240 778 116409 798
<< psubdiffcont >>
rect 113387 2777 113450 2838
rect 113517 2777 113580 2838
rect 113647 2777 113710 2838
rect 113777 2777 113840 2838
rect 113907 2777 113970 2838
rect 114037 2777 114100 2838
rect 114167 2777 114230 2838
rect 114297 2777 114360 2838
rect 114427 2777 114490 2838
rect 114557 2777 114620 2838
rect 114687 2777 114750 2838
rect 114817 2777 114880 2838
rect 114947 2777 115010 2838
rect 115077 2777 115140 2838
rect 115207 2777 115270 2838
rect 115337 2777 115400 2838
rect 115467 2777 115530 2838
rect 115597 2777 115660 2838
rect 115727 2777 115790 2838
rect 115857 2777 115920 2838
rect 115987 2777 116050 2838
rect 116117 2777 116180 2838
rect 113258 2714 113321 2775
rect 113258 2584 113321 2645
rect 113258 2454 113321 2515
rect 113258 2324 113321 2385
rect 113258 2194 113321 2255
rect 113258 2064 113321 2125
rect 113258 1934 113321 1995
rect 113258 1804 113321 1865
rect 116329 2732 116392 2793
rect 116329 2602 116392 2663
rect 116329 2472 116392 2533
rect 116329 2342 116392 2403
rect 116329 2212 116392 2273
rect 116329 2082 116392 2143
rect 116329 1952 116392 2013
rect 113258 1674 113321 1735
rect 113258 1544 113321 1605
rect 116329 1822 116392 1883
rect 116329 1692 116392 1753
rect 116329 1562 116392 1623
rect 113258 1414 113321 1475
rect 113258 1284 113321 1345
rect 113258 1154 113321 1215
rect 113258 1024 113321 1085
rect 113258 894 113321 955
rect 116329 1432 116392 1493
rect 116329 1302 116392 1363
rect 116329 1172 116392 1233
rect 116329 1042 116392 1103
rect 116329 912 116392 973
rect 113371 798 113434 859
rect 113501 798 113564 859
rect 113631 798 113694 859
rect 113761 798 113824 859
rect 113891 798 113954 859
rect 114021 798 114084 859
rect 114151 798 114214 859
rect 114281 798 114344 859
rect 114411 798 114474 859
rect 114541 798 114604 859
rect 114671 798 114734 859
rect 114801 798 114864 859
rect 114931 798 114994 859
rect 115061 798 115124 859
rect 115191 798 115254 859
rect 115321 798 115384 859
rect 115451 798 115514 859
rect 115581 798 115644 859
rect 115711 798 115774 859
rect 115841 798 115904 859
rect 115971 798 116034 859
rect 116101 798 116164 859
rect 116231 798 116294 859
<< polysilicon >>
rect 113528 1729 113628 1842
rect 113528 1671 113547 1729
rect 113606 1671 113628 1729
rect 113859 1810 115782 1842
rect 113859 1747 115006 1810
rect 115069 1808 115782 1810
rect 115069 1747 115144 1808
rect 113859 1745 115144 1747
rect 115207 1745 115782 1808
rect 113859 1726 115782 1745
rect 113528 1550 113628 1671
rect 116015 1722 116115 1842
rect 113860 1646 115783 1666
rect 113860 1583 114184 1646
rect 114247 1644 115783 1646
rect 114247 1583 114322 1644
rect 113860 1581 114322 1583
rect 114385 1581 115783 1644
rect 113860 1550 115783 1581
rect 116015 1664 116034 1722
rect 116093 1664 116115 1722
rect 116015 1550 116115 1664
<< polycontact >>
rect 113547 1671 113606 1729
rect 115006 1747 115069 1810
rect 115144 1745 115207 1808
rect 114184 1583 114247 1646
rect 114322 1581 114385 1644
rect 116034 1664 116093 1722
<< metal1 >>
rect 56587 16439 92016 17147
rect 56587 16113 57295 16439
rect 59737 16113 60445 16439
rect 62978 16113 63686 16439
rect 68397 16113 69105 16439
rect 72016 16113 72724 16439
rect 75401 16113 76109 16439
rect 78264 16113 78972 16439
rect 81847 16113 82555 16439
rect 85772 16113 86480 16439
rect 88922 16113 89630 16439
rect 91308 16113 92016 16439
rect 127187 16313 158887 17021
rect 127187 16113 127895 16313
rect 131718 16113 132426 16313
rect 134509 16113 135217 16313
rect 137771 16113 138479 16313
rect 140744 16113 141452 16313
rect 143317 16113 144025 16313
rect 145637 16113 146345 16313
rect 147921 16113 148629 16313
rect 151292 16113 152000 16313
rect 154627 16113 155335 16313
rect 158179 16113 158887 16313
rect 12617 15405 189263 16113
rect 12617 13631 13325 15405
rect 15224 15081 15932 15405
rect 18778 15081 19486 15405
rect 21309 15081 22017 15405
rect 23500 15081 24208 15405
rect 27065 15081 27773 15405
rect 29769 15081 30477 15405
rect 32838 15081 33546 15405
rect 40835 15081 41543 15405
rect 45268 15081 45976 15405
rect 50677 15081 51385 15405
rect 56905 15081 57613 15405
rect 59353 15081 60061 15405
rect 13804 14373 60061 15081
rect 88646 14698 89354 15405
rect 91864 14698 92572 15405
rect 94959 14698 95667 15405
rect 98938 14698 99646 15405
rect 102899 14698 103607 15405
rect 107638 14698 108346 15405
rect 112112 14698 112820 15405
rect 117400 14698 118108 15405
rect 119700 14698 120408 15405
rect 121800 14698 122508 15405
rect 123104 14698 123812 15405
rect 124469 14698 125177 15405
rect 127390 14698 128098 15405
rect 128672 14698 129380 15405
rect 13804 13631 14512 14373
rect 17117 13631 17825 14373
rect 558 13370 884 13480
rect 558 13318 599 13370
rect 651 13318 703 13370
rect 755 13318 807 13370
rect 859 13318 884 13370
rect 558 13266 884 13318
rect 558 13214 599 13266
rect 651 13214 703 13266
rect 755 13214 807 13266
rect 859 13214 884 13266
rect 558 13162 884 13214
rect 558 13110 599 13162
rect 651 13110 703 13162
rect 755 13110 807 13162
rect 859 13110 884 13162
rect 558 -3337 884 13110
rect 12617 12923 17825 13631
rect 12617 11465 13325 12923
rect 13804 11328 14512 12923
rect 17117 12546 17825 12923
rect 18778 12546 19486 14373
rect 21309 12992 22017 14373
rect 23500 12744 24208 14373
rect 27065 12777 27773 14373
rect 29769 12702 30477 14373
rect 32838 12801 33546 14373
rect 40835 13008 41543 14373
rect 45268 12901 45976 14373
rect 50677 13000 51385 14373
rect 56905 13629 57613 14373
rect 59353 13182 60061 14373
rect 61675 13660 84753 14376
rect 61675 13135 62391 13660
rect 65909 13111 66625 13660
rect 69460 13120 70176 13660
rect 73269 13034 73985 13660
rect 76858 13073 77574 13660
rect 79913 12987 80629 13660
rect 17117 11838 19486 12546
rect 15882 10624 15981 10640
rect 15882 10558 15899 10624
rect 15966 10558 15981 10624
rect 15882 10542 15981 10558
rect 17117 9676 17825 11838
rect 18778 11458 19486 11838
rect 18778 10750 20842 11458
rect 18778 9676 19486 10750
rect 17117 8968 19486 9676
rect 15870 8288 15969 8304
rect 15870 8222 15887 8288
rect 15954 8222 15969 8288
rect 15870 8206 15969 8222
rect 17117 7364 17825 8968
rect 18778 7894 19486 8968
rect 50610 10606 51318 12969
rect 84037 12939 84753 13660
rect 88646 13990 129380 14698
rect 157382 14737 158090 15405
rect 162130 14737 162838 15405
rect 167096 14737 167804 15405
rect 169996 14737 170704 15405
rect 173476 14737 174184 15405
rect 178297 14737 179005 15405
rect 182465 14737 183173 15405
rect 188555 14737 189263 15405
rect 88646 12616 89354 13990
rect 91864 12581 92572 13990
rect 94959 12528 95667 13990
rect 98938 12599 99646 13990
rect 102899 12563 103607 13990
rect 107638 12599 108346 13990
rect 112112 12616 112820 13990
rect 117400 12563 118108 13990
rect 119700 12565 120408 13990
rect 121800 13468 122508 13990
rect 123104 13604 123812 13990
rect 124469 13604 125177 13990
rect 123104 13468 125177 13604
rect 127390 13570 128098 13990
rect 128672 13570 129380 13990
rect 130357 14443 154005 14577
rect 130357 14442 139232 14443
rect 130357 14440 138898 14442
rect 130357 14439 134010 14440
rect 130357 14437 133676 14439
rect 130357 14349 133349 14437
rect 133436 14349 133529 14437
rect 133616 14351 133676 14437
rect 133763 14351 133856 14439
rect 133943 14352 134010 14439
rect 134097 14424 138571 14440
rect 134097 14423 136516 14424
rect 134097 14421 136182 14423
rect 134097 14352 135855 14421
rect 133943 14351 135855 14352
rect 133616 14349 135855 14351
rect 130357 14333 135855 14349
rect 135942 14333 136035 14421
rect 136122 14335 136182 14421
rect 136269 14335 136362 14423
rect 136449 14336 136516 14423
rect 136603 14352 138571 14424
rect 138658 14352 138751 14440
rect 138838 14354 138898 14440
rect 138985 14354 139078 14442
rect 139165 14355 139232 14442
rect 139319 14355 154005 14443
rect 139165 14354 154005 14355
rect 138838 14352 154005 14354
rect 136603 14336 154005 14352
rect 136449 14335 154005 14336
rect 136122 14333 154005 14335
rect 130357 14263 154005 14333
rect 130357 14262 139232 14263
rect 130357 14260 138898 14262
rect 130357 14259 134010 14260
rect 130357 14257 133676 14259
rect 130357 13868 130677 14257
rect 131815 13890 132135 14257
rect 133251 14169 133349 14257
rect 133436 14169 133529 14257
rect 133616 14171 133676 14257
rect 133763 14171 133856 14259
rect 133943 14172 134010 14259
rect 134097 14257 138571 14260
rect 134097 14172 134136 14257
rect 133943 14171 134136 14172
rect 133616 14169 134136 14171
rect 133251 14047 134136 14169
rect 133251 14046 133992 14047
rect 133251 14044 133658 14046
rect 133251 13956 133331 14044
rect 133418 13956 133511 14044
rect 133598 13958 133658 14044
rect 133745 13958 133838 14046
rect 133925 13959 133992 14046
rect 134079 13959 134136 14047
rect 133925 13958 134136 13959
rect 133598 13956 134136 13958
rect 133251 13867 134136 13956
rect 133251 13866 133992 13867
rect 133251 13864 133658 13866
rect 133251 13776 133331 13864
rect 133418 13776 133511 13864
rect 133598 13778 133658 13864
rect 133745 13778 133838 13866
rect 133925 13779 133992 13866
rect 134079 13779 134136 13867
rect 133925 13778 134136 13779
rect 133598 13776 134136 13778
rect 133251 13698 134136 13776
rect 133251 13685 133571 13698
rect 134893 13628 135213 14257
rect 135785 14244 136642 14257
rect 135785 14243 136516 14244
rect 135785 14241 136182 14243
rect 135785 14153 135855 14241
rect 135942 14153 136035 14241
rect 136122 14155 136182 14241
rect 136269 14155 136362 14243
rect 136449 14156 136516 14243
rect 136603 14156 136642 14244
rect 136449 14155 136642 14156
rect 136122 14153 136642 14155
rect 135785 14031 136642 14153
rect 135785 14030 136498 14031
rect 135785 14028 136164 14030
rect 135785 13940 135837 14028
rect 135924 13940 136017 14028
rect 136104 13942 136164 14028
rect 136251 13942 136344 14030
rect 136431 13943 136498 14030
rect 136585 13943 136642 14031
rect 136431 13942 136642 13943
rect 136104 13940 136642 13942
rect 135785 13851 136642 13940
rect 135785 13850 136498 13851
rect 135785 13848 136164 13850
rect 135785 13768 135837 13848
rect 135784 13760 135837 13768
rect 135924 13760 136017 13848
rect 136104 13762 136164 13848
rect 136251 13762 136344 13850
rect 136431 13763 136498 13850
rect 136585 13763 136642 13851
rect 137874 13847 138194 14257
rect 138501 14172 138571 14257
rect 138658 14172 138751 14260
rect 138838 14174 138898 14260
rect 138985 14174 139078 14262
rect 139165 14175 139232 14262
rect 139319 14257 154005 14263
rect 139319 14175 139358 14257
rect 139165 14174 139358 14175
rect 138838 14172 139358 14174
rect 138501 14050 139358 14172
rect 138501 14049 139214 14050
rect 138501 14047 138880 14049
rect 138501 13959 138553 14047
rect 138640 13959 138733 14047
rect 138820 13961 138880 14047
rect 138967 13961 139060 14049
rect 139147 13962 139214 14049
rect 139301 13962 139358 14050
rect 139147 13961 139358 13962
rect 138820 13959 139358 13961
rect 138501 13870 139358 13959
rect 138501 13869 139214 13870
rect 138501 13867 138880 13869
rect 138501 13787 138553 13867
rect 136431 13762 136642 13763
rect 136104 13760 136642 13762
rect 135784 13682 136642 13760
rect 138500 13779 138553 13787
rect 138640 13779 138733 13867
rect 138820 13781 138880 13867
rect 138967 13781 139060 13869
rect 139147 13782 139214 13869
rect 139301 13782 139358 13870
rect 139147 13781 139358 13782
rect 138820 13779 139358 13781
rect 138500 13701 139358 13779
rect 139915 13760 140235 14257
rect 141589 13814 141909 14257
rect 143900 13804 144220 14257
rect 146417 13771 146737 14257
rect 148479 13793 148799 14257
rect 151179 13836 151499 14257
rect 153685 13814 154005 14257
rect 157382 14029 189263 14737
rect 121800 12896 125177 13468
rect 157382 13377 158090 14029
rect 162130 13304 162838 14029
rect 167096 13268 167804 14029
rect 169996 13377 170704 14029
rect 173476 13449 174184 14029
rect 178297 13341 179005 14029
rect 182465 13341 183173 14029
rect 188555 13377 189263 14029
rect 121800 12760 123812 12896
rect 50610 9898 56230 10606
rect 18778 7364 20867 7894
rect 15873 7207 15972 7223
rect 15873 7141 15890 7207
rect 15957 7141 15972 7207
rect 15873 7125 15972 7141
rect 17117 7186 20867 7364
rect 50610 7754 51318 9898
rect 121800 9665 122508 12760
rect 123104 11863 123812 12760
rect 124469 11863 125177 12896
rect 123104 11155 125177 11863
rect 123104 9678 123812 11155
rect 124469 10121 125177 11155
rect 123104 9665 124465 9678
rect 121800 9622 124465 9665
rect 120448 8970 124465 9622
rect 120448 8957 123812 8970
rect 120448 8914 122508 8957
rect 17117 6656 19486 7186
rect 11871 5470 12579 5919
rect 14552 5470 15260 5899
rect 17117 5470 17825 6656
rect 11745 5216 17825 5470
rect 18778 6107 19486 6656
rect 50610 7046 55201 7754
rect 18778 5399 20859 6107
rect 18778 5216 19486 5399
rect 11745 4762 19486 5216
rect 17117 4508 19486 4762
rect 17117 2437 17825 4508
rect 18778 2437 19486 4508
rect 50610 3535 51318 7046
rect 121800 7040 122508 8914
rect 123104 8294 123812 8957
rect 123104 7586 124465 8294
rect 120484 6332 122508 7040
rect 150298 6671 151141 6731
rect 150298 6670 151003 6671
rect 150298 6668 150669 6670
rect 150298 6580 150342 6668
rect 150429 6580 150522 6668
rect 150609 6582 150669 6668
rect 150756 6582 150849 6670
rect 150936 6583 151003 6670
rect 151090 6583 151141 6671
rect 150936 6582 151141 6583
rect 150609 6580 151141 6582
rect 150298 6491 151141 6580
rect 150298 6490 151003 6491
rect 150298 6488 150669 6490
rect 150298 6400 150342 6488
rect 150429 6400 150522 6488
rect 150609 6402 150669 6488
rect 150756 6402 150849 6490
rect 150936 6403 151003 6490
rect 151090 6403 151141 6491
rect 150936 6402 151141 6403
rect 150609 6400 151141 6402
rect 150298 6356 151141 6400
rect 80879 6043 81977 6073
rect 75608 5997 76748 6038
rect 75608 5996 76309 5997
rect 75608 5994 75975 5996
rect 75608 5906 75648 5994
rect 75735 5906 75828 5994
rect 75915 5908 75975 5994
rect 76062 5908 76155 5996
rect 76242 5909 76309 5996
rect 76396 5996 76748 5997
rect 76396 5909 76449 5996
rect 76242 5908 76449 5909
rect 76536 5994 76748 5996
rect 76536 5908 76590 5994
rect 75915 5906 76590 5908
rect 76677 5906 76748 5994
rect 75608 5817 76748 5906
rect 75608 5816 76309 5817
rect 75608 5814 75975 5816
rect 75608 5726 75648 5814
rect 75735 5726 75828 5814
rect 75915 5728 75975 5814
rect 76062 5728 76155 5816
rect 76242 5729 76309 5816
rect 76396 5816 76748 5817
rect 76396 5729 76449 5816
rect 76242 5728 76449 5729
rect 76536 5814 76748 5816
rect 76536 5728 76590 5814
rect 75915 5726 76590 5728
rect 76677 5726 76748 5814
rect 75608 5683 76748 5726
rect 80879 6033 81982 6043
rect 80879 6032 81734 6033
rect 80879 6031 81580 6032
rect 80879 6029 81246 6031
rect 80879 5941 80919 6029
rect 81006 5941 81099 6029
rect 81186 5943 81246 6029
rect 81333 5943 81426 6031
rect 81513 5944 81580 6031
rect 81667 5945 81734 6032
rect 81821 6031 81982 6033
rect 81821 5945 81882 6031
rect 81667 5944 81882 5945
rect 81513 5943 81882 5944
rect 81969 5943 81982 6031
rect 81186 5941 81982 5943
rect 80879 5853 81982 5941
rect 80879 5852 81734 5853
rect 80879 5851 81580 5852
rect 80879 5849 81246 5851
rect 80879 5761 80919 5849
rect 81006 5761 81099 5849
rect 81186 5763 81246 5849
rect 81333 5763 81426 5851
rect 81513 5764 81580 5851
rect 81667 5765 81734 5852
rect 81821 5851 81982 5853
rect 81821 5765 81882 5851
rect 81667 5764 81882 5765
rect 81513 5763 81882 5764
rect 81969 5763 81982 5851
rect 81186 5761 81982 5763
rect 80879 5746 81982 5761
rect 80879 5718 81977 5746
rect 56833 4217 57127 4231
rect 56833 4129 56847 4217
rect 56934 4129 57027 4217
rect 57114 4129 57127 4217
rect 56833 4037 57127 4129
rect 56833 3949 56847 4037
rect 56934 3949 57027 4037
rect 57114 3949 57127 4037
rect 56833 3935 57127 3949
rect 115054 3958 115376 3977
rect 114442 3912 114764 3930
rect 113812 3862 114134 3879
rect 113812 3774 113837 3862
rect 113924 3774 114017 3862
rect 114104 3774 114134 3862
rect 113812 3682 114134 3774
rect 113812 3594 113837 3682
rect 113924 3594 114017 3682
rect 114104 3594 114134 3682
rect 17117 1729 19486 2437
rect 1983 -640 2422 -15
rect 3921 -640 4360 -15
rect 6028 -640 6467 38
rect 8536 -640 8975 -57
rect 10011 -640 10450 -67
rect 12392 -640 12831 -4
rect 14589 -640 15028 17
rect 1983 -1079 15028 -640
rect 17117 -31 17825 1729
rect 18778 -31 19486 1729
rect 44263 2827 55277 3535
rect 113812 3521 114134 3594
rect 113812 3433 113839 3521
rect 113926 3433 114019 3521
rect 114106 3433 114134 3521
rect 113812 3341 114134 3433
rect 113812 3253 113839 3341
rect 113926 3253 114019 3341
rect 114106 3253 114134 3341
rect 114442 3824 114475 3912
rect 114562 3824 114655 3912
rect 114742 3824 114764 3912
rect 114442 3732 114764 3824
rect 114442 3644 114475 3732
rect 114562 3644 114655 3732
rect 114742 3644 114764 3732
rect 114442 3569 114764 3644
rect 114442 3481 114473 3569
rect 114560 3481 114653 3569
rect 114740 3481 114764 3569
rect 114442 3389 114764 3481
rect 114442 3301 114473 3389
rect 114560 3301 114653 3389
rect 114740 3301 114764 3389
rect 115054 3870 115082 3958
rect 115169 3870 115262 3958
rect 115349 3870 115376 3958
rect 115054 3778 115376 3870
rect 115054 3690 115082 3778
rect 115169 3690 115262 3778
rect 115349 3690 115376 3778
rect 115054 3618 115376 3690
rect 115054 3530 115082 3618
rect 115169 3530 115262 3618
rect 115349 3530 115376 3618
rect 115054 3438 115376 3530
rect 115054 3350 115082 3438
rect 115169 3350 115262 3438
rect 115349 3350 115376 3438
rect 115054 3329 115376 3350
rect 115708 3940 116010 3955
rect 115708 3852 115729 3940
rect 115816 3852 115909 3940
rect 115996 3852 116010 3940
rect 115708 3760 116010 3852
rect 115708 3672 115729 3760
rect 115816 3672 115909 3760
rect 115996 3672 116010 3760
rect 115708 3623 116010 3672
rect 119380 3704 120088 5063
rect 121800 4040 122508 6332
rect 126212 4902 126506 4916
rect 126212 4814 126226 4902
rect 126313 4814 126406 4902
rect 126493 4814 126506 4902
rect 126212 4722 126506 4814
rect 126212 4634 126226 4722
rect 126313 4634 126406 4722
rect 126493 4634 126506 4722
rect 126212 4620 126506 4634
rect 121800 3704 124015 4040
rect 115708 3609 116012 3623
rect 115708 3521 115732 3609
rect 115819 3521 115912 3609
rect 115999 3521 116012 3609
rect 115708 3429 116012 3521
rect 115708 3341 115732 3429
rect 115819 3341 115912 3429
rect 115999 3341 116012 3429
rect 115708 3327 116012 3341
rect 119380 3332 124015 3704
rect 115708 3317 116010 3327
rect 114442 3282 114764 3301
rect 113812 3231 114134 3253
rect 119380 2996 122508 3332
rect 113211 2838 116439 2888
rect 44263 2280 44971 2827
rect 50610 2280 51318 2827
rect 52315 2280 53023 2827
rect 113211 2777 113387 2838
rect 113450 2777 113517 2838
rect 113580 2777 113647 2838
rect 113710 2777 113777 2838
rect 113840 2777 113907 2838
rect 113970 2777 114037 2838
rect 114100 2777 114167 2838
rect 114230 2777 114297 2838
rect 114360 2777 114427 2838
rect 114490 2777 114557 2838
rect 114620 2777 114687 2838
rect 114750 2777 114817 2838
rect 114880 2777 114947 2838
rect 115010 2777 115077 2838
rect 115140 2777 115207 2838
rect 115270 2777 115337 2838
rect 115400 2777 115467 2838
rect 115530 2777 115597 2838
rect 115660 2777 115727 2838
rect 115790 2777 115857 2838
rect 115920 2777 115987 2838
rect 116050 2777 116117 2838
rect 116180 2793 116439 2838
rect 116180 2777 116329 2793
rect 113211 2775 116329 2777
rect 113211 2714 113258 2775
rect 113321 2732 116329 2775
rect 116392 2732 116439 2793
rect 113321 2730 116439 2732
rect 113321 2714 113369 2730
rect 113211 2645 113369 2714
rect 113211 2584 113258 2645
rect 113321 2584 113369 2645
rect 113211 2515 113369 2584
rect 113211 2454 113258 2515
rect 113321 2454 113369 2515
rect 113211 2385 113369 2454
rect 113211 2324 113258 2385
rect 113321 2324 113369 2385
rect 44263 1572 55294 2280
rect 113211 2255 113369 2324
rect 113211 2194 113258 2255
rect 113321 2194 113369 2255
rect 113211 2125 113369 2194
rect 113211 2064 113258 2125
rect 113321 2064 113369 2125
rect 113211 1995 113369 2064
rect 113211 1934 113258 1995
rect 113321 1934 113369 1995
rect 113211 1865 113369 1934
rect 113211 1804 113258 1865
rect 113321 1804 113369 1865
rect 113211 1735 113369 1804
rect 113211 1674 113258 1735
rect 113321 1674 113369 1735
rect 113211 1605 113369 1674
rect 17117 -739 19486 -31
rect 28005 680 28862 753
rect 28005 679 28736 680
rect 28005 677 28402 679
rect 28005 589 28075 677
rect 28162 589 28255 677
rect 28342 591 28402 677
rect 28489 591 28582 679
rect 28669 592 28736 679
rect 28823 592 28862 680
rect 28669 591 28862 592
rect 28342 589 28862 591
rect 28005 500 28862 589
rect 28005 499 28736 500
rect 28005 497 28402 499
rect 28005 409 28075 497
rect 28162 409 28255 497
rect 28342 411 28402 497
rect 28489 411 28582 499
rect 28669 412 28736 499
rect 28823 412 28862 500
rect 28669 411 28862 412
rect 28342 409 28862 411
rect 28005 287 28862 409
rect 28005 286 28718 287
rect 28005 284 28384 286
rect 28005 196 28057 284
rect 28144 196 28237 284
rect 28324 198 28384 284
rect 28471 198 28564 286
rect 28651 199 28718 286
rect 28805 199 28862 287
rect 28651 198 28862 199
rect 28324 196 28862 198
rect 28005 107 28862 196
rect 28005 106 28718 107
rect 28005 104 28384 106
rect 28005 16 28057 104
rect 28144 16 28237 104
rect 28324 18 28384 104
rect 28471 18 28564 106
rect 28651 19 28718 106
rect 28805 19 28862 107
rect 28651 18 28862 19
rect 28324 16 28862 18
rect 28005 -63 28862 16
rect 29817 727 30674 793
rect 29817 726 30542 727
rect 29817 724 30208 726
rect 29817 636 29881 724
rect 29968 636 30061 724
rect 30148 638 30208 724
rect 30295 638 30388 726
rect 30475 639 30542 726
rect 30629 639 30674 727
rect 30475 638 30674 639
rect 30148 636 30674 638
rect 29817 547 30674 636
rect 29817 546 30542 547
rect 29817 544 30208 546
rect 29817 456 29881 544
rect 29968 456 30061 544
rect 30148 458 30208 544
rect 30295 458 30388 546
rect 30475 459 30542 546
rect 30629 459 30674 547
rect 30475 458 30674 459
rect 30148 456 30674 458
rect 29817 339 30674 456
rect 29817 338 30548 339
rect 29817 336 30214 338
rect 29817 248 29887 336
rect 29974 248 30067 336
rect 30154 250 30214 336
rect 30301 250 30394 338
rect 30481 251 30548 338
rect 30635 251 30674 339
rect 30481 250 30674 251
rect 30154 248 30674 250
rect 29817 159 30674 248
rect 29817 158 30548 159
rect 29817 156 30214 158
rect 29817 68 29887 156
rect 29974 68 30067 156
rect 30154 70 30214 156
rect 30301 70 30394 158
rect 30481 71 30548 158
rect 30635 71 30674 159
rect 30481 70 30674 71
rect 30154 68 30674 70
rect 29817 -23 30674 68
rect 31572 727 32429 770
rect 31572 726 32279 727
rect 31572 724 31945 726
rect 31572 636 31618 724
rect 31705 636 31798 724
rect 31885 638 31945 724
rect 32032 638 32125 726
rect 32212 639 32279 726
rect 32366 639 32429 727
rect 32212 638 32429 639
rect 31885 636 32429 638
rect 31572 547 32429 636
rect 31572 546 32279 547
rect 31572 544 31945 546
rect 31572 456 31618 544
rect 31705 456 31798 544
rect 31885 458 31945 544
rect 32032 458 32125 546
rect 32212 459 32279 546
rect 32366 459 32429 547
rect 32212 458 32429 459
rect 31885 456 32429 458
rect 31572 339 32429 456
rect 31572 338 32291 339
rect 31572 336 31957 338
rect 31572 248 31630 336
rect 31717 248 31810 336
rect 31897 250 31957 336
rect 32044 250 32137 338
rect 32224 251 32291 338
rect 32378 251 32429 339
rect 32224 250 32429 251
rect 31897 248 32429 250
rect 31572 159 32429 248
rect 31572 158 32291 159
rect 31572 156 31957 158
rect 31572 68 31630 156
rect 31717 68 31810 156
rect 31897 70 31957 156
rect 32044 70 32137 158
rect 32224 71 32291 158
rect 32378 71 32429 159
rect 32224 70 32429 71
rect 31897 68 32429 70
rect 31572 -46 32429 68
rect 1983 -2026 2422 -1079
rect 3921 -2026 4360 -1079
rect 6028 -2026 6467 -1079
rect 8536 -2026 8975 -1079
rect 10011 -2026 10450 -1079
rect 17117 -2624 17825 -739
rect 18778 -798 19486 -739
rect 44263 -798 44971 1572
rect 47306 923 47412 1103
rect 47550 476 47726 948
rect 47817 862 48021 969
rect 47817 810 47846 862
rect 47898 810 47950 862
rect 48002 810 48021 862
rect 47817 758 48021 810
rect 47817 706 47846 758
rect 47898 706 47950 758
rect 48002 706 48021 758
rect 47817 674 48021 706
rect 48111 476 48287 947
rect 48383 825 48568 953
rect 48665 825 48850 951
rect 48986 927 49092 1107
rect 48383 764 48850 825
rect 48383 699 48410 764
rect 48475 699 48535 764
rect 48600 699 48660 764
rect 48725 699 48850 764
rect 48383 640 48850 699
rect 47550 300 48287 476
rect 47830 -477 48573 -297
rect 18778 -1506 46711 -798
rect 47299 -1067 47405 -887
rect 47581 -1069 47690 -885
rect 47830 -911 48010 -477
rect 48100 -624 48295 -601
rect 48100 -676 48120 -624
rect 48172 -676 48224 -624
rect 48276 -676 48295 -624
rect 48100 -728 48295 -676
rect 48100 -780 48120 -728
rect 48172 -780 48224 -728
rect 48276 -780 48295 -728
rect 48100 -903 48295 -780
rect 48393 -914 48573 -477
rect 48661 -631 48856 -602
rect 48661 -683 48678 -631
rect 48730 -683 48782 -631
rect 48834 -683 48856 -631
rect 48661 -735 48856 -683
rect 48661 -787 48678 -735
rect 48730 -787 48782 -735
rect 48834 -787 48856 -735
rect 48661 -904 48856 -787
rect 18778 -2624 19486 -1506
rect 20705 -2176 21413 -1506
rect 22947 -2142 23655 -1506
rect 27130 -2176 27838 -1506
rect 29171 -2209 29879 -1506
rect 31112 -2326 31820 -1506
rect 33069 -2192 33777 -1506
rect 34977 -2259 35685 -1506
rect 38172 -2042 38880 -1506
rect 40598 -2042 41306 -1506
rect 42874 -1874 43582 -1506
rect 46003 -1975 46711 -1506
rect 47944 -1835 48339 -1049
rect 48982 -1060 49088 -880
rect 50610 -2186 51318 1572
rect 11741 -3332 20561 -2624
rect 558 -3349 934 -3337
rect 558 -3401 662 -3349
rect 714 -3401 766 -3349
rect 818 -3401 870 -3349
rect 922 -3401 934 -3349
rect 558 -3453 934 -3401
rect 558 -3505 662 -3453
rect 714 -3505 766 -3453
rect 818 -3505 870 -3453
rect 922 -3505 934 -3453
rect 558 -3557 934 -3505
rect 558 -3609 662 -3557
rect 714 -3609 766 -3557
rect 818 -3609 870 -3557
rect 922 -3609 934 -3557
rect 558 -3621 934 -3609
rect 558 -18230 884 -3621
rect 11741 -3827 12449 -3332
rect 14802 -3827 15510 -3332
rect 17117 -3827 17825 -3332
rect 11741 -4535 17825 -3827
rect 11741 -5353 12449 -4535
rect 14802 -5392 15510 -4535
rect 52315 -6069 53023 1572
rect 113211 1544 113258 1605
rect 113321 1544 113369 1605
rect 113211 1475 113369 1544
rect 113211 1414 113258 1475
rect 113321 1414 113369 1475
rect 113211 1345 113369 1414
rect 113211 1284 113258 1345
rect 113321 1284 113369 1345
rect 113211 1215 113369 1284
rect 113211 1154 113258 1215
rect 113321 1154 113369 1215
rect 113211 1085 113369 1154
rect 113211 1024 113258 1085
rect 113321 1024 113369 1085
rect 113211 955 113369 1024
rect 113211 894 113258 955
rect 113321 910 113369 955
rect 113453 1755 113499 2730
rect 113657 1755 113703 2730
rect 113897 2660 114113 2675
rect 113897 2595 113912 2660
rect 113974 2595 114037 2660
rect 114099 2595 114113 2660
rect 113897 2535 114113 2595
rect 113897 2470 113912 2535
rect 113974 2470 114037 2535
rect 114099 2470 114113 2535
rect 113897 2456 114113 2470
rect 114443 2660 114659 2675
rect 114443 2595 114458 2660
rect 114520 2595 114583 2660
rect 114645 2595 114659 2660
rect 114443 2535 114659 2595
rect 114443 2470 114458 2535
rect 114520 2470 114583 2535
rect 114645 2470 114659 2535
rect 114443 2456 114659 2470
rect 114971 2651 115187 2666
rect 114971 2586 114986 2651
rect 115048 2586 115111 2651
rect 115173 2586 115187 2651
rect 114971 2526 115187 2586
rect 114971 2461 114986 2526
rect 115048 2461 115111 2526
rect 115173 2461 115187 2526
rect 113975 1888 114052 2456
rect 113453 1729 113703 1755
rect 113453 1671 113547 1729
rect 113606 1671 113703 1729
rect 113785 1819 113831 1888
rect 114193 1819 114239 1888
rect 113785 1713 114239 1819
rect 114325 1825 114371 1888
rect 114515 1886 114592 2456
rect 114971 2447 115187 2461
rect 115520 2653 115736 2668
rect 115520 2588 115535 2653
rect 115597 2588 115660 2653
rect 115722 2588 115736 2653
rect 115520 2528 115736 2588
rect 115520 2463 115535 2528
rect 115597 2463 115660 2528
rect 115722 2463 115736 2528
rect 115520 2449 115736 2463
rect 114733 1825 114779 1888
rect 114325 1719 114779 1825
rect 113453 1642 113703 1671
rect 113453 910 113499 1642
rect 113657 910 113703 1642
rect 113767 910 113844 1513
rect 113974 1020 114051 1713
rect 114165 1646 114402 1661
rect 114165 1583 114184 1646
rect 114247 1644 114402 1646
rect 114247 1583 114322 1644
rect 114165 1581 114322 1583
rect 114385 1581 114402 1644
rect 114165 1569 114402 1581
rect 114176 910 114253 1517
rect 114307 910 114384 1513
rect 114514 1020 114591 1719
rect 114865 1672 114911 1888
rect 115055 1874 115132 2447
rect 114987 1810 115224 1825
rect 114987 1747 115006 1810
rect 115069 1808 115224 1810
rect 115069 1747 115144 1808
rect 114987 1745 115144 1747
rect 115207 1745 115224 1808
rect 114987 1733 115224 1745
rect 115273 1672 115319 1888
rect 114865 1566 115319 1672
rect 115404 1756 115450 1888
rect 115594 1874 115671 2449
rect 115812 1756 115858 1888
rect 115404 1650 115858 1756
rect 115940 1748 115986 2730
rect 116144 1748 116190 2730
rect 115940 1722 116190 1748
rect 115940 1664 116034 1722
rect 116093 1664 116190 1722
rect 114716 910 114793 1517
rect 114847 910 114924 1506
rect 115054 1020 115131 1566
rect 115256 910 115333 1507
rect 115386 910 115463 1513
rect 115593 1020 115670 1650
rect 115940 1635 116190 1664
rect 115795 910 115872 1517
rect 115940 910 115986 1635
rect 116144 910 116190 1635
rect 116281 2663 116439 2730
rect 116281 2602 116329 2663
rect 116392 2602 116439 2663
rect 116281 2533 116439 2602
rect 116281 2472 116329 2533
rect 116392 2472 116439 2533
rect 116281 2403 116439 2472
rect 116281 2342 116329 2403
rect 116392 2342 116439 2403
rect 116281 2273 116439 2342
rect 116281 2212 116329 2273
rect 116392 2212 116439 2273
rect 116281 2143 116439 2212
rect 116281 2082 116329 2143
rect 116392 2082 116439 2143
rect 116281 2013 116439 2082
rect 116281 1952 116329 2013
rect 116392 1952 116439 2013
rect 116281 1883 116439 1952
rect 116281 1822 116329 1883
rect 116392 1822 116439 1883
rect 116281 1753 116439 1822
rect 116281 1692 116329 1753
rect 116392 1692 116439 1753
rect 116281 1623 116439 1692
rect 116281 1562 116329 1623
rect 116392 1562 116439 1623
rect 116281 1493 116439 1562
rect 116281 1432 116329 1493
rect 116392 1432 116439 1493
rect 116281 1363 116439 1432
rect 116281 1302 116329 1363
rect 116392 1302 116439 1363
rect 116281 1233 116439 1302
rect 116281 1172 116329 1233
rect 116392 1172 116439 1233
rect 116281 1103 116439 1172
rect 116281 1042 116329 1103
rect 116392 1042 116439 1103
rect 116281 973 116439 1042
rect 116281 912 116329 973
rect 116392 912 116439 973
rect 116281 910 116439 912
rect 113321 894 116439 910
rect 113211 859 116439 894
rect 113211 798 113371 859
rect 113434 798 113501 859
rect 113564 798 113631 859
rect 113694 798 113761 859
rect 113824 798 113891 859
rect 113954 798 114021 859
rect 114084 798 114151 859
rect 114214 798 114281 859
rect 114344 798 114411 859
rect 114474 798 114541 859
rect 114604 798 114671 859
rect 114734 798 114801 859
rect 114864 798 114931 859
rect 114994 798 115061 859
rect 115124 798 115191 859
rect 115254 798 115321 859
rect 115384 798 115451 859
rect 115514 798 115581 859
rect 115644 798 115711 859
rect 115774 798 115841 859
rect 115904 798 115971 859
rect 116034 798 116101 859
rect 116164 798 116231 859
rect 116294 798 116439 859
rect 113211 752 116439 798
rect 113735 -864 114443 752
rect 115168 58 115876 752
rect 115168 -125 116924 58
rect 115168 -127 116292 -125
rect 115168 -179 115977 -127
rect 116029 -179 116081 -127
rect 116133 -179 116185 -127
rect 116237 -177 116292 -127
rect 116344 -177 116396 -125
rect 116448 -177 116500 -125
rect 116552 -177 116607 -125
rect 116659 -177 116711 -125
rect 116763 -177 116815 -125
rect 116867 -177 116924 -125
rect 116237 -179 116924 -177
rect 115168 -229 116924 -179
rect 115168 -231 116292 -229
rect 115168 -283 115977 -231
rect 116029 -283 116081 -231
rect 116133 -283 116185 -231
rect 116237 -281 116292 -231
rect 116344 -281 116396 -229
rect 116448 -281 116500 -229
rect 116552 -281 116607 -229
rect 116659 -281 116711 -229
rect 116763 -281 116815 -229
rect 116867 -281 116924 -229
rect 116237 -283 116924 -281
rect 115168 -333 116924 -283
rect 115168 -335 116292 -333
rect 115168 -387 115977 -335
rect 116029 -387 116081 -335
rect 116133 -387 116185 -335
rect 116237 -385 116292 -335
rect 116344 -385 116396 -333
rect 116448 -385 116500 -333
rect 116552 -385 116607 -333
rect 116659 -385 116711 -333
rect 116763 -385 116815 -333
rect 116867 -385 116924 -333
rect 116237 -387 116924 -385
rect 115168 -621 116924 -387
rect 115168 -864 115876 -621
rect 113735 -1572 115876 -864
rect 55067 -3335 55775 -1833
rect 55067 -4043 58644 -3335
rect 55067 -6069 55775 -4043
rect 113735 -4392 114443 -1572
rect 115168 -4392 115876 -1572
rect 113735 -5100 115876 -4392
rect 16024 -6142 16123 -6126
rect 16024 -6208 16041 -6142
rect 16108 -6208 16123 -6142
rect 16024 -6224 16123 -6208
rect 52315 -6777 57395 -6069
rect 16028 -8484 16127 -8468
rect 16028 -8550 16045 -8484
rect 16112 -8550 16127 -8484
rect 16028 -8566 16127 -8550
rect 55067 -9090 55775 -6777
rect 113735 -7892 114443 -5100
rect 115168 -7892 115876 -5100
rect 113735 -8600 115876 -7892
rect 16041 -9562 16140 -9546
rect 16041 -9628 16058 -9562
rect 16125 -9628 16140 -9562
rect 16041 -9644 16140 -9628
rect 55067 -9798 57412 -9090
rect 113735 -9858 114443 -8600
rect 115168 -9858 115876 -8600
rect 86265 -10566 115876 -9858
rect 86265 -12576 86973 -10566
rect 90080 -12576 90788 -10566
rect 94470 -12576 95178 -10566
rect 98233 -12576 98941 -10566
rect 102205 -12576 102913 -10566
rect 106856 -12576 107564 -10566
rect 110201 -12576 110909 -10566
rect 113735 -12301 114443 -10566
rect 115168 -12301 115876 -10566
rect 119380 -3576 120088 2996
rect 121800 1587 122508 2996
rect 121800 879 123892 1587
rect 129992 310 130341 530
rect 127066 268 130341 310
rect 127066 266 127460 268
rect 127066 214 127145 266
rect 127197 214 127249 266
rect 127301 214 127353 266
rect 127405 216 127460 266
rect 127512 216 127564 268
rect 127616 216 127668 268
rect 127720 216 127775 268
rect 127827 216 127879 268
rect 127931 216 127983 268
rect 128035 216 130341 268
rect 127405 214 130341 216
rect 127066 164 130341 214
rect 127066 162 127460 164
rect 127066 110 127145 162
rect 127197 110 127249 162
rect 127301 110 127353 162
rect 127405 112 127460 162
rect 127512 112 127564 164
rect 127616 112 127668 164
rect 127720 112 127775 164
rect 127827 112 127879 164
rect 127931 112 127983 164
rect 128035 112 130341 164
rect 127405 110 130341 112
rect 127066 60 130341 110
rect 127066 58 127460 60
rect 127066 6 127145 58
rect 127197 6 127249 58
rect 127301 6 127353 58
rect 127405 8 127460 58
rect 127512 8 127564 60
rect 127616 8 127668 60
rect 127720 8 127775 60
rect 127827 8 127879 60
rect 127931 8 127983 60
rect 128035 8 130341 60
rect 127405 6 130341 8
rect 127066 -39 130341 6
rect 120821 -3185 120962 -3012
rect 121086 -3506 121279 -3167
rect 121365 -3241 121560 -3158
rect 121365 -3293 121385 -3241
rect 121437 -3293 121489 -3241
rect 121541 -3293 121560 -3241
rect 121365 -3345 121560 -3293
rect 121365 -3397 121385 -3345
rect 121437 -3397 121489 -3345
rect 121541 -3397 121560 -3345
rect 121365 -3420 121560 -3397
rect 121645 -3506 121838 -3170
rect 121926 -3234 122121 -3158
rect 121926 -3286 121943 -3234
rect 121995 -3286 122047 -3234
rect 122099 -3286 122121 -3234
rect 121926 -3338 122121 -3286
rect 121926 -3390 121943 -3338
rect 121995 -3390 122047 -3338
rect 122099 -3390 122121 -3338
rect 122203 -3171 122402 -3149
rect 122482 -3171 122681 -3154
rect 122203 -3240 122681 -3171
rect 122784 -3187 122925 -3014
rect 122203 -3307 122342 -3240
rect 122406 -3245 122681 -3240
rect 122406 -3307 122474 -3245
rect 122203 -3312 122474 -3307
rect 122538 -3312 122681 -3245
rect 122203 -3364 122681 -3312
rect 122203 -3365 122472 -3364
rect 122203 -3370 122347 -3365
rect 121926 -3419 122121 -3390
rect 122311 -3432 122347 -3370
rect 122411 -3431 122472 -3365
rect 122536 -3370 122681 -3364
rect 122536 -3431 122558 -3370
rect 122411 -3432 122558 -3431
rect 122311 -3441 122558 -3432
rect 122319 -3466 122556 -3441
rect 119380 -4284 120687 -3576
rect 121086 -3699 121838 -3506
rect 121003 -3877 121260 -3833
rect 121003 -3880 121167 -3877
rect 121003 -3946 121036 -3880
rect 121102 -3943 121167 -3880
rect 121233 -3911 121260 -3877
rect 121233 -3943 121298 -3911
rect 121102 -3946 121298 -3943
rect 121003 -4009 121298 -3946
rect 121003 -4075 121035 -4009
rect 121101 -4075 121169 -4009
rect 121235 -4028 121298 -4009
rect 121235 -4075 121569 -4028
rect 121003 -4137 121569 -4075
rect 121003 -4203 121032 -4137
rect 121098 -4203 121167 -4137
rect 121233 -4203 121569 -4137
rect 121003 -4239 121569 -4203
rect 121003 -4274 121260 -4239
rect 119380 -10248 120088 -4284
rect 120832 -4875 120973 -4709
rect 121111 -4875 121252 -4706
rect 121358 -4752 121569 -4239
rect 121645 -4396 122398 -4203
rect 121645 -4735 121838 -4396
rect 121923 -4485 122118 -4462
rect 121923 -4537 121943 -4485
rect 121995 -4537 122047 -4485
rect 122099 -4537 122118 -4485
rect 121923 -4589 122118 -4537
rect 121923 -4641 121943 -4589
rect 121995 -4641 122047 -4589
rect 122099 -4641 122118 -4589
rect 121923 -4744 122118 -4641
rect 122205 -4734 122398 -4396
rect 122484 -4492 122679 -4463
rect 123072 -4478 123818 -3915
rect 168112 -4239 173993 -3531
rect 122484 -4544 122501 -4492
rect 122553 -4544 122605 -4492
rect 122657 -4544 122679 -4492
rect 122484 -4596 122679 -4544
rect 122484 -4648 122501 -4596
rect 122553 -4648 122605 -4596
rect 122657 -4648 122679 -4596
rect 122484 -4744 122679 -4648
rect 120832 -4879 121252 -4875
rect 120832 -4882 121203 -4879
rect 120876 -5317 121203 -4882
rect 122797 -4885 122938 -4712
rect 120876 -5644 123858 -5317
rect 172133 -7987 172841 -4239
rect 173285 -7987 173993 -4239
rect 172133 -8695 173993 -7987
rect 145837 -8792 146487 -8759
rect 145837 -8844 145860 -8792
rect 145912 -8844 145964 -8792
rect 146016 -8844 146068 -8792
rect 146120 -8844 146201 -8792
rect 146253 -8844 146305 -8792
rect 146357 -8844 146409 -8792
rect 146461 -8844 146487 -8792
rect 145837 -8896 146487 -8844
rect 145837 -8948 145860 -8896
rect 145912 -8948 145964 -8896
rect 146016 -8948 146068 -8896
rect 146120 -8948 146201 -8896
rect 146253 -8948 146305 -8896
rect 146357 -8948 146409 -8896
rect 146461 -8948 146487 -8896
rect 145837 -9000 146487 -8948
rect 145837 -9052 145860 -9000
rect 145912 -9052 145964 -9000
rect 146016 -9052 146068 -9000
rect 146120 -9052 146201 -9000
rect 146253 -9052 146305 -9000
rect 146357 -9052 146409 -9000
rect 146461 -9052 146487 -9000
rect 145837 -9075 146487 -9052
rect 119380 -10956 124421 -10248
rect 113735 -12576 115876 -12301
rect 86265 -13009 115876 -12576
rect 86265 -13284 114443 -13009
rect 20515 -14849 21039 -14033
rect 24264 -14849 24972 -14367
rect 27785 -14849 28493 -14292
rect 31251 -14849 31959 -14236
rect 34301 -14849 35009 -14349
rect 41646 -14849 42354 -14236
rect 45017 -14849 45725 -14405
rect 50742 -14849 51450 -14236
rect 54979 -14849 55687 -14311
rect 59405 -14849 60113 -14349
rect 63529 -14849 64237 -14273
rect 69273 -14849 69981 -14198
rect 73002 -14849 73710 -14254
rect 75550 -14725 76478 -14704
rect 75550 -14813 75573 -14725
rect 75660 -14813 75733 -14725
rect 75820 -14813 75893 -14725
rect 75980 -14813 76053 -14725
rect 76140 -14813 76213 -14725
rect 76300 -14813 76373 -14725
rect 76460 -14813 76478 -14725
rect 75550 -14849 76478 -14813
rect 86265 -14849 86973 -13284
rect 90080 -14849 90788 -13284
rect 94470 -14849 95178 -13284
rect 98233 -14849 98941 -13284
rect 102205 -14849 102913 -13284
rect 106856 -14849 107564 -13284
rect 110201 -14849 110909 -13284
rect 113735 -13501 114443 -13284
rect 115168 -13501 115876 -13009
rect 133308 -13430 134166 -13355
rect 133308 -13431 134040 -13430
rect 133308 -13433 133706 -13431
rect 133308 -13501 133379 -13433
rect 113735 -13521 133379 -13501
rect 133466 -13521 133559 -13433
rect 133646 -13519 133706 -13433
rect 133793 -13519 133886 -13431
rect 133973 -13518 134040 -13431
rect 134127 -13501 134166 -13430
rect 135746 -13435 136604 -13360
rect 135746 -13436 136478 -13435
rect 135746 -13438 136144 -13436
rect 135746 -13501 135817 -13438
rect 134127 -13518 135817 -13501
rect 133973 -13519 135817 -13518
rect 133646 -13521 135817 -13519
rect 113735 -13526 135817 -13521
rect 135904 -13526 135997 -13438
rect 136084 -13524 136144 -13438
rect 136231 -13524 136324 -13436
rect 136411 -13523 136478 -13436
rect 136565 -13501 136604 -13435
rect 138468 -13441 139326 -13366
rect 138468 -13442 139200 -13441
rect 138468 -13444 138866 -13442
rect 138468 -13501 138539 -13444
rect 136565 -13523 138539 -13501
rect 136411 -13524 138539 -13523
rect 136084 -13526 138539 -13524
rect 113735 -13532 138539 -13526
rect 138626 -13532 138719 -13444
rect 138806 -13530 138866 -13444
rect 138953 -13530 139046 -13442
rect 139133 -13529 139200 -13442
rect 139287 -13501 139326 -13441
rect 150251 -13408 151108 -13335
rect 150251 -13409 150982 -13408
rect 150251 -13411 150648 -13409
rect 150251 -13499 150321 -13411
rect 150408 -13499 150501 -13411
rect 150588 -13497 150648 -13411
rect 150735 -13497 150828 -13409
rect 150915 -13496 150982 -13409
rect 151069 -13496 151108 -13408
rect 150915 -13497 151108 -13496
rect 150588 -13499 151108 -13497
rect 150251 -13501 151108 -13499
rect 172133 -13501 172841 -8695
rect 173285 -13501 173993 -8695
rect 139287 -13529 173993 -13501
rect 139133 -13530 173993 -13529
rect 138806 -13532 173993 -13530
rect 113735 -13588 173993 -13532
rect 113735 -13589 150982 -13588
rect 113735 -13591 150648 -13589
rect 113735 -13604 150321 -13591
rect 113735 -13610 145840 -13604
rect 113735 -13611 134040 -13610
rect 113735 -13613 133706 -13611
rect 113735 -13701 133379 -13613
rect 133466 -13701 133559 -13613
rect 133646 -13699 133706 -13613
rect 133793 -13699 133886 -13611
rect 133973 -13698 134040 -13611
rect 134127 -13615 145840 -13610
rect 134127 -13616 136478 -13615
rect 134127 -13618 136144 -13616
rect 134127 -13698 135817 -13618
rect 133973 -13699 135817 -13698
rect 133646 -13701 135817 -13699
rect 113735 -13706 135817 -13701
rect 135904 -13706 135997 -13618
rect 136084 -13704 136144 -13618
rect 136231 -13704 136324 -13616
rect 136411 -13703 136478 -13616
rect 136565 -13621 145840 -13615
rect 136565 -13622 139200 -13621
rect 136565 -13624 138866 -13622
rect 136565 -13703 138539 -13624
rect 136411 -13704 138539 -13703
rect 136084 -13706 138539 -13704
rect 113735 -13712 138539 -13706
rect 138626 -13712 138719 -13624
rect 138806 -13710 138866 -13624
rect 138953 -13710 139046 -13622
rect 139133 -13709 139200 -13622
rect 139287 -13656 145840 -13621
rect 145892 -13656 145944 -13604
rect 145996 -13656 146048 -13604
rect 146100 -13656 146181 -13604
rect 146233 -13656 146285 -13604
rect 146337 -13656 146389 -13604
rect 146441 -13656 150321 -13604
rect 139287 -13679 150321 -13656
rect 150408 -13679 150501 -13591
rect 150588 -13677 150648 -13591
rect 150735 -13677 150828 -13589
rect 150915 -13676 150982 -13589
rect 151069 -13676 173993 -13588
rect 150915 -13677 173993 -13676
rect 150588 -13679 173993 -13677
rect 139287 -13708 173993 -13679
rect 139287 -13709 145840 -13708
rect 139133 -13710 145840 -13709
rect 138806 -13712 145840 -13710
rect 113735 -13760 145840 -13712
rect 145892 -13760 145944 -13708
rect 145996 -13760 146048 -13708
rect 146100 -13760 146181 -13708
rect 146233 -13760 146285 -13708
rect 146337 -13760 146389 -13708
rect 146441 -13760 173993 -13708
rect 113735 -13801 173993 -13760
rect 113735 -13802 150964 -13801
rect 113735 -13804 150630 -13802
rect 113735 -13812 150303 -13804
rect 113735 -13823 145840 -13812
rect 113735 -13824 134022 -13823
rect 113735 -13826 133688 -13824
rect 113735 -13914 133361 -13826
rect 133448 -13914 133541 -13826
rect 133628 -13912 133688 -13826
rect 133775 -13912 133868 -13824
rect 133955 -13911 134022 -13824
rect 134109 -13828 145840 -13823
rect 134109 -13829 136460 -13828
rect 134109 -13831 136126 -13829
rect 134109 -13911 135799 -13831
rect 133955 -13912 135799 -13911
rect 133628 -13914 135799 -13912
rect 113735 -13919 135799 -13914
rect 135886 -13919 135979 -13831
rect 136066 -13917 136126 -13831
rect 136213 -13917 136306 -13829
rect 136393 -13916 136460 -13829
rect 136547 -13834 145840 -13828
rect 136547 -13835 139182 -13834
rect 136547 -13837 138848 -13835
rect 136547 -13916 138521 -13837
rect 136393 -13917 138521 -13916
rect 136066 -13919 138521 -13917
rect 113735 -13925 138521 -13919
rect 138608 -13925 138701 -13837
rect 138788 -13923 138848 -13837
rect 138935 -13923 139028 -13835
rect 139115 -13922 139182 -13835
rect 139269 -13864 145840 -13834
rect 145892 -13864 145944 -13812
rect 145996 -13864 146048 -13812
rect 146100 -13864 146181 -13812
rect 146233 -13864 146285 -13812
rect 146337 -13864 146389 -13812
rect 146441 -13864 150303 -13812
rect 139269 -13892 150303 -13864
rect 150390 -13892 150483 -13804
rect 150570 -13890 150630 -13804
rect 150717 -13890 150810 -13802
rect 150897 -13889 150964 -13802
rect 151051 -13889 173993 -13801
rect 150897 -13890 173993 -13889
rect 150570 -13892 173993 -13890
rect 139269 -13922 173993 -13892
rect 139115 -13923 173993 -13922
rect 138788 -13925 173993 -13923
rect 113735 -13981 173993 -13925
rect 113735 -13982 150964 -13981
rect 113735 -13984 150630 -13982
rect 113735 -14003 150303 -13984
rect 113735 -14004 134022 -14003
rect 113735 -14006 133688 -14004
rect 113735 -14094 133361 -14006
rect 133448 -14094 133541 -14006
rect 133628 -14092 133688 -14006
rect 133775 -14092 133868 -14004
rect 133955 -14091 134022 -14004
rect 134109 -14008 150303 -14003
rect 134109 -14009 136460 -14008
rect 134109 -14011 136126 -14009
rect 134109 -14091 135799 -14011
rect 133955 -14092 135799 -14091
rect 133628 -14094 135799 -14092
rect 113735 -14099 135799 -14094
rect 135886 -14099 135979 -14011
rect 136066 -14097 136126 -14011
rect 136213 -14097 136306 -14009
rect 136393 -14096 136460 -14009
rect 136547 -14014 150303 -14008
rect 136547 -14015 139182 -14014
rect 136547 -14017 138848 -14015
rect 136547 -14096 138521 -14017
rect 136393 -14097 138521 -14096
rect 136066 -14099 138521 -14097
rect 113735 -14105 138521 -14099
rect 138608 -14105 138701 -14017
rect 138788 -14103 138848 -14017
rect 138935 -14103 139028 -14015
rect 139115 -14102 139182 -14015
rect 139269 -14072 150303 -14014
rect 150390 -14072 150483 -13984
rect 150570 -14070 150630 -13984
rect 150717 -14070 150810 -13982
rect 150897 -14069 150964 -13982
rect 151051 -14069 173993 -13981
rect 150897 -14070 173993 -14069
rect 150570 -14072 173993 -14070
rect 139269 -14102 173993 -14072
rect 139115 -14103 173993 -14102
rect 138788 -14105 173993 -14103
rect 113735 -14209 173993 -14105
rect 113735 -14849 114443 -14209
rect 115168 -14849 115876 -14209
rect 120089 -14849 120797 -14209
rect 128589 -14849 129297 -14209
rect 134435 -14849 135143 -14209
rect 140249 -14849 140957 -14209
rect 145147 -14849 145855 -14209
rect 149254 -14849 149962 -14209
rect 152138 -14849 152846 -14209
rect 156331 -14849 157039 -14209
rect 162222 -14849 162930 -14209
rect 167574 -14849 168282 -14209
rect 172133 -14849 172841 -14209
rect 173285 -14849 173993 -14209
rect 17096 -14885 173993 -14849
rect 17096 -14973 75573 -14885
rect 75660 -14973 75733 -14885
rect 75820 -14973 75893 -14885
rect 75980 -14973 76053 -14885
rect 76140 -14973 76213 -14885
rect 76300 -14973 76373 -14885
rect 76460 -14936 173993 -14885
rect 76460 -14937 81435 -14936
rect 76460 -14939 81101 -14937
rect 76460 -14973 80774 -14939
rect 17096 -15027 80774 -14973
rect 80861 -15027 80954 -14939
rect 81041 -15025 81101 -14939
rect 81188 -15025 81281 -14937
rect 81368 -15024 81435 -14937
rect 81522 -14938 173993 -14936
rect 81522 -14939 81759 -14938
rect 81522 -15024 81605 -14939
rect 81368 -15025 81605 -15024
rect 81041 -15027 81605 -15025
rect 81692 -15026 81759 -14939
rect 81846 -15026 173993 -14938
rect 81692 -15027 173993 -15026
rect 17096 -15045 173993 -15027
rect 17096 -15133 75573 -15045
rect 75660 -15133 75733 -15045
rect 75820 -15133 75893 -15045
rect 75980 -15133 76053 -15045
rect 76140 -15133 76213 -15045
rect 76300 -15133 76373 -15045
rect 76460 -15116 173993 -15045
rect 76460 -15117 81435 -15116
rect 76460 -15119 81101 -15117
rect 76460 -15133 80774 -15119
rect 17096 -15205 80774 -15133
rect 17096 -15275 75573 -15205
rect 17096 -15361 31543 -15275
rect 17096 -15449 29831 -15361
rect 29918 -15449 29991 -15361
rect 30078 -15449 30151 -15361
rect 30238 -15449 30311 -15361
rect 30398 -15449 30471 -15361
rect 30558 -15449 30631 -15361
rect 30718 -15363 31543 -15361
rect 31630 -15363 31703 -15275
rect 31790 -15363 31863 -15275
rect 31950 -15363 32023 -15275
rect 32110 -15363 32183 -15275
rect 32270 -15363 32343 -15275
rect 32430 -15293 75573 -15275
rect 75660 -15293 75733 -15205
rect 75820 -15293 75893 -15205
rect 75980 -15293 76053 -15205
rect 76140 -15293 76213 -15205
rect 76300 -15293 76373 -15205
rect 76460 -15207 80774 -15205
rect 80861 -15207 80954 -15119
rect 81041 -15205 81101 -15119
rect 81188 -15205 81281 -15117
rect 81368 -15204 81435 -15117
rect 81522 -15118 173993 -15116
rect 81522 -15119 81759 -15118
rect 81522 -15204 81605 -15119
rect 81368 -15205 81605 -15204
rect 81041 -15207 81605 -15205
rect 81692 -15206 81759 -15119
rect 81846 -15206 173993 -15118
rect 81692 -15207 173993 -15206
rect 76460 -15293 173993 -15207
rect 32430 -15294 81429 -15293
rect 32430 -15296 81095 -15294
rect 32430 -15363 80768 -15296
rect 30718 -15365 80768 -15363
rect 30718 -15435 75573 -15365
rect 30718 -15449 31543 -15435
rect 17096 -15478 31543 -15449
rect 17096 -15557 28009 -15478
rect 17096 -16083 17804 -15557
rect 18872 -16083 19580 -15557
rect 25936 -16083 26644 -15557
rect 27885 -15566 28009 -15557
rect 28096 -15566 28169 -15478
rect 28256 -15566 28329 -15478
rect 28416 -15566 28489 -15478
rect 28576 -15566 28649 -15478
rect 28736 -15566 28809 -15478
rect 28896 -15521 31543 -15478
rect 28896 -15557 29831 -15521
rect 28896 -15566 29050 -15557
rect 27885 -15638 29050 -15566
rect 27885 -15726 28009 -15638
rect 28096 -15726 28169 -15638
rect 28256 -15726 28329 -15638
rect 28416 -15726 28489 -15638
rect 28576 -15726 28649 -15638
rect 28736 -15726 28809 -15638
rect 28896 -15726 29050 -15638
rect 27885 -15798 29050 -15726
rect 27885 -15886 28009 -15798
rect 28096 -15886 28169 -15798
rect 28256 -15886 28329 -15798
rect 28416 -15886 28489 -15798
rect 28576 -15886 28649 -15798
rect 28736 -15886 28809 -15798
rect 28896 -15886 29050 -15798
rect 27885 -15958 29050 -15886
rect 27885 -16046 28009 -15958
rect 28096 -16046 28169 -15958
rect 28256 -16046 28329 -15958
rect 28416 -16046 28489 -15958
rect 28576 -16046 28649 -15958
rect 28736 -16046 28809 -15958
rect 28896 -16046 29050 -15958
rect 27885 -16083 29050 -16046
rect 29808 -15609 29831 -15557
rect 29918 -15609 29991 -15521
rect 30078 -15609 30151 -15521
rect 30238 -15609 30311 -15521
rect 30398 -15609 30471 -15521
rect 30558 -15609 30631 -15521
rect 30718 -15523 31543 -15521
rect 31630 -15523 31703 -15435
rect 31790 -15523 31863 -15435
rect 31950 -15523 32023 -15435
rect 32110 -15523 32183 -15435
rect 32270 -15523 32343 -15435
rect 32430 -15453 75573 -15435
rect 75660 -15453 75733 -15365
rect 75820 -15453 75893 -15365
rect 75980 -15453 76053 -15365
rect 76140 -15453 76213 -15365
rect 76300 -15453 76373 -15365
rect 76460 -15384 80768 -15365
rect 80855 -15384 80948 -15296
rect 81035 -15382 81095 -15296
rect 81182 -15382 81275 -15294
rect 81362 -15381 81429 -15294
rect 81516 -15295 173993 -15293
rect 81516 -15296 81753 -15295
rect 81516 -15381 81599 -15296
rect 81362 -15382 81599 -15381
rect 81035 -15384 81599 -15382
rect 81686 -15383 81753 -15296
rect 81840 -15383 173993 -15295
rect 81686 -15384 173993 -15383
rect 76460 -15453 173993 -15384
rect 32430 -15523 173993 -15453
rect 30718 -15525 173993 -15523
rect 30718 -15557 75573 -15525
rect 30718 -15609 30736 -15557
rect 29808 -15681 30736 -15609
rect 29808 -15769 29831 -15681
rect 29918 -15769 29991 -15681
rect 30078 -15769 30151 -15681
rect 30238 -15769 30311 -15681
rect 30398 -15769 30471 -15681
rect 30558 -15769 30631 -15681
rect 30718 -15769 30736 -15681
rect 29808 -15841 30736 -15769
rect 29808 -15929 29831 -15841
rect 29918 -15929 29991 -15841
rect 30078 -15929 30151 -15841
rect 30238 -15929 30311 -15841
rect 30398 -15929 30471 -15841
rect 30558 -15929 30631 -15841
rect 30718 -15929 30736 -15841
rect 29808 -16001 30736 -15929
rect 29808 -16083 29831 -16001
rect 17096 -16089 29831 -16083
rect 29918 -16089 29991 -16001
rect 30078 -16089 30151 -16001
rect 30238 -16089 30311 -16001
rect 30398 -16089 30471 -16001
rect 30558 -16089 30631 -16001
rect 30718 -16083 30736 -16001
rect 31520 -15595 32448 -15557
rect 31520 -15683 31543 -15595
rect 31630 -15683 31703 -15595
rect 31790 -15683 31863 -15595
rect 31950 -15683 32023 -15595
rect 32110 -15683 32183 -15595
rect 32270 -15683 32343 -15595
rect 32430 -15683 32448 -15595
rect 31520 -15755 32448 -15683
rect 31520 -15843 31543 -15755
rect 31630 -15843 31703 -15755
rect 31790 -15843 31863 -15755
rect 31950 -15843 32023 -15755
rect 32110 -15843 32183 -15755
rect 32270 -15843 32343 -15755
rect 32430 -15843 32448 -15755
rect 31520 -15915 32448 -15843
rect 31520 -16003 31543 -15915
rect 31630 -16003 31703 -15915
rect 31790 -16003 31863 -15915
rect 31950 -16003 32023 -15915
rect 32110 -16003 32183 -15915
rect 32270 -16003 32343 -15915
rect 32430 -16003 32448 -15915
rect 31520 -16075 32448 -16003
rect 31520 -16083 31543 -16075
rect 30718 -16089 31543 -16083
rect 17096 -16118 31543 -16089
rect 17096 -16206 28009 -16118
rect 28096 -16206 28169 -16118
rect 28256 -16206 28329 -16118
rect 28416 -16206 28489 -16118
rect 28576 -16206 28649 -16118
rect 28736 -16206 28809 -16118
rect 28896 -16161 31543 -16118
rect 28896 -16206 29831 -16161
rect 17096 -16249 29831 -16206
rect 29918 -16249 29991 -16161
rect 30078 -16249 30151 -16161
rect 30238 -16249 30311 -16161
rect 30398 -16249 30471 -16161
rect 30558 -16249 30631 -16161
rect 30718 -16163 31543 -16161
rect 31630 -16163 31703 -16075
rect 31790 -16163 31863 -16075
rect 31950 -16163 32023 -16075
rect 32110 -16163 32183 -16075
rect 32270 -16163 32343 -16075
rect 32430 -16083 32448 -16075
rect 32660 -16083 33368 -15557
rect 39937 -16083 40645 -15557
rect 46788 -16083 47496 -15557
rect 51852 -16083 52560 -15557
rect 56704 -16083 57412 -15557
rect 61342 -16083 62050 -15557
rect 66832 -16083 67540 -15557
rect 73003 -16083 73711 -15557
rect 75550 -15613 75573 -15557
rect 75660 -15613 75733 -15525
rect 75820 -15613 75893 -15525
rect 75980 -15613 76053 -15525
rect 76140 -15613 76213 -15525
rect 76300 -15613 76373 -15525
rect 76460 -15557 173993 -15525
rect 76460 -15613 76478 -15557
rect 75550 -15635 76478 -15613
rect 78321 -16083 79029 -15557
rect 80861 -15965 81789 -15944
rect 80861 -16053 80884 -15965
rect 80971 -16053 81044 -15965
rect 81131 -16053 81204 -15965
rect 81291 -16053 81364 -15965
rect 81451 -16053 81524 -15965
rect 81611 -16053 81684 -15965
rect 81771 -16053 81789 -15965
rect 80861 -16083 81789 -16053
rect 83171 -16083 83879 -15557
rect 87856 -16083 88564 -15557
rect 92872 -16083 93580 -15557
rect 97530 -16083 98238 -15557
rect 102077 -16083 102785 -15557
rect 106927 -16083 107635 -15557
rect 111227 -16083 111935 -15557
rect 115168 -16083 115876 -15557
rect 32430 -16125 115876 -16083
rect 32430 -16163 80884 -16125
rect 30718 -16213 80884 -16163
rect 80971 -16213 81044 -16125
rect 81131 -16213 81204 -16125
rect 81291 -16213 81364 -16125
rect 81451 -16213 81524 -16125
rect 81611 -16213 81684 -16125
rect 81771 -16213 115876 -16125
rect 30718 -16249 115876 -16213
rect 17096 -16264 115876 -16249
rect 17096 -16265 76313 -16264
rect 17096 -16267 75979 -16265
rect 17096 -16278 75652 -16267
rect 17096 -16366 28009 -16278
rect 28096 -16366 28169 -16278
rect 28256 -16366 28329 -16278
rect 28416 -16366 28489 -16278
rect 28576 -16366 28649 -16278
rect 28736 -16366 28809 -16278
rect 28896 -16355 75652 -16278
rect 75739 -16355 75832 -16267
rect 75919 -16353 75979 -16267
rect 76066 -16353 76159 -16265
rect 76246 -16352 76313 -16265
rect 76400 -16266 115876 -16264
rect 76400 -16267 76637 -16266
rect 76400 -16352 76483 -16267
rect 76246 -16353 76483 -16352
rect 75919 -16355 76483 -16353
rect 76570 -16354 76637 -16267
rect 76724 -16285 115876 -16266
rect 76724 -16354 80884 -16285
rect 76570 -16355 80884 -16354
rect 28896 -16366 80884 -16355
rect 17096 -16373 80884 -16366
rect 80971 -16373 81044 -16285
rect 81131 -16373 81204 -16285
rect 81291 -16373 81364 -16285
rect 81451 -16373 81524 -16285
rect 81611 -16373 81684 -16285
rect 81771 -16373 115876 -16285
rect 17096 -16444 115876 -16373
rect 17096 -16445 76313 -16444
rect 17096 -16447 75979 -16445
rect 17096 -16535 75652 -16447
rect 75739 -16535 75832 -16447
rect 75919 -16533 75979 -16447
rect 76066 -16533 76159 -16445
rect 76246 -16532 76313 -16445
rect 76400 -16445 115876 -16444
rect 76400 -16446 80884 -16445
rect 76400 -16447 76637 -16446
rect 76400 -16532 76483 -16447
rect 76246 -16533 76483 -16532
rect 75919 -16535 76483 -16533
rect 76570 -16534 76637 -16447
rect 76724 -16533 80884 -16446
rect 80971 -16533 81044 -16445
rect 81131 -16533 81204 -16445
rect 81291 -16533 81364 -16445
rect 81451 -16533 81524 -16445
rect 81611 -16533 81684 -16445
rect 81771 -16533 115876 -16445
rect 76724 -16534 115876 -16533
rect 76570 -16535 115876 -16534
rect 17096 -16605 115876 -16535
rect 17096 -16621 80884 -16605
rect 17096 -16622 76307 -16621
rect 17096 -16624 75973 -16622
rect 1373 -17133 2081 -16731
rect 3955 -17133 4663 -16731
rect 7066 -17133 7774 -16731
rect 11806 -17133 12514 -16710
rect 17096 -16712 75646 -16624
rect 75733 -16712 75826 -16624
rect 75913 -16710 75973 -16624
rect 76060 -16710 76153 -16622
rect 76240 -16709 76307 -16622
rect 76394 -16623 80884 -16621
rect 76394 -16624 76631 -16623
rect 76394 -16709 76477 -16624
rect 76240 -16710 76477 -16709
rect 75913 -16712 76477 -16710
rect 76564 -16711 76631 -16624
rect 76718 -16693 80884 -16623
rect 80971 -16693 81044 -16605
rect 81131 -16693 81204 -16605
rect 81291 -16693 81364 -16605
rect 81451 -16693 81524 -16605
rect 81611 -16693 81684 -16605
rect 81771 -16693 115876 -16605
rect 76718 -16711 115876 -16693
rect 76564 -16712 115876 -16711
rect 17096 -16765 115876 -16712
rect 17096 -16791 80884 -16765
rect 17096 -17133 17804 -16791
rect 18872 -17133 19580 -16791
rect 80861 -16853 80884 -16791
rect 80971 -16853 81044 -16765
rect 81131 -16853 81204 -16765
rect 81291 -16853 81364 -16765
rect 81451 -16853 81524 -16765
rect 81611 -16853 81684 -16765
rect 81771 -16791 115876 -16765
rect 81771 -16853 81789 -16791
rect 80861 -16875 81789 -16853
rect 1373 -17841 19580 -17133
rect 27267 -18163 28195 -18142
rect 454 -18329 967 -18230
rect 27267 -18251 27290 -18163
rect 27377 -18251 27450 -18163
rect 27537 -18251 27610 -18163
rect 27697 -18251 27770 -18163
rect 27857 -18251 27930 -18163
rect 28017 -18251 28090 -18163
rect 28177 -18251 28195 -18163
rect 27267 -18323 28195 -18251
rect 290 -18349 1099 -18329
rect 290 -18432 312 -18349
rect 395 -18432 482 -18349
rect 565 -18432 652 -18349
rect 735 -18432 822 -18349
rect 905 -18432 992 -18349
rect 1075 -18432 1099 -18349
rect 290 -18519 1099 -18432
rect 290 -18602 312 -18519
rect 395 -18602 482 -18519
rect 565 -18602 652 -18519
rect 735 -18602 822 -18519
rect 905 -18602 992 -18519
rect 1075 -18602 1099 -18519
rect 290 -18689 1099 -18602
rect 290 -18772 312 -18689
rect 395 -18772 482 -18689
rect 565 -18772 652 -18689
rect 735 -18772 822 -18689
rect 905 -18772 992 -18689
rect 1075 -18772 1099 -18689
rect 290 -18859 1099 -18772
rect 290 -18942 312 -18859
rect 395 -18942 482 -18859
rect 565 -18942 652 -18859
rect 735 -18942 822 -18859
rect 905 -18942 992 -18859
rect 1075 -18942 1099 -18859
rect 290 -19029 1099 -18942
rect 290 -19112 312 -19029
rect 395 -19112 482 -19029
rect 565 -19112 652 -19029
rect 735 -19112 822 -19029
rect 905 -19112 992 -19029
rect 1075 -19112 1099 -19029
rect 27267 -18411 27290 -18323
rect 27377 -18411 27450 -18323
rect 27537 -18411 27610 -18323
rect 27697 -18411 27770 -18323
rect 27857 -18411 27930 -18323
rect 28017 -18411 28090 -18323
rect 28177 -18411 28195 -18323
rect 27267 -18483 28195 -18411
rect 27267 -18571 27290 -18483
rect 27377 -18571 27450 -18483
rect 27537 -18571 27610 -18483
rect 27697 -18571 27770 -18483
rect 27857 -18571 27930 -18483
rect 28017 -18571 28090 -18483
rect 28177 -18571 28195 -18483
rect 27267 -18643 28195 -18571
rect 27267 -18731 27290 -18643
rect 27377 -18731 27450 -18643
rect 27537 -18731 27610 -18643
rect 27697 -18731 27770 -18643
rect 27857 -18731 27930 -18643
rect 28017 -18731 28090 -18643
rect 28177 -18731 28195 -18643
rect 27267 -18803 28195 -18731
rect 27267 -18891 27290 -18803
rect 27377 -18891 27450 -18803
rect 27537 -18891 27610 -18803
rect 27697 -18891 27770 -18803
rect 27857 -18891 27930 -18803
rect 28017 -18891 28090 -18803
rect 28177 -18891 28195 -18803
rect 27267 -18963 28195 -18891
rect 27267 -19051 27290 -18963
rect 27377 -19051 27450 -18963
rect 27537 -19051 27610 -18963
rect 27697 -19051 27770 -18963
rect 27857 -19051 27930 -18963
rect 28017 -19051 28090 -18963
rect 28177 -19051 28195 -18963
rect 27267 -19073 28195 -19051
rect 290 -19134 1099 -19112
rect 27896 -19446 28694 -19411
rect 27896 -19447 28594 -19446
rect 27896 -19449 28260 -19447
rect 27896 -19537 27933 -19449
rect 28020 -19537 28113 -19449
rect 28200 -19535 28260 -19449
rect 28347 -19535 28440 -19447
rect 28527 -19534 28594 -19447
rect 28681 -19534 28694 -19446
rect 28527 -19535 28694 -19534
rect 28200 -19537 28694 -19535
rect 27896 -19569 28694 -19537
<< via1 >>
rect 599 13318 651 13370
rect 703 13318 755 13370
rect 807 13318 859 13370
rect 599 13214 651 13266
rect 703 13214 755 13266
rect 807 13214 859 13266
rect 599 13110 651 13162
rect 703 13110 755 13162
rect 807 13110 859 13162
rect 15899 10558 15966 10624
rect 15887 8222 15954 8288
rect 133349 14349 133436 14437
rect 133529 14349 133616 14437
rect 133676 14351 133763 14439
rect 133856 14351 133943 14439
rect 134010 14352 134097 14440
rect 135855 14333 135942 14421
rect 136035 14333 136122 14421
rect 136182 14335 136269 14423
rect 136362 14335 136449 14423
rect 136516 14336 136603 14424
rect 138571 14352 138658 14440
rect 138751 14352 138838 14440
rect 138898 14354 138985 14442
rect 139078 14354 139165 14442
rect 139232 14355 139319 14443
rect 133349 14169 133436 14257
rect 133529 14169 133616 14257
rect 133676 14171 133763 14259
rect 133856 14171 133943 14259
rect 134010 14172 134097 14260
rect 133331 13956 133418 14044
rect 133511 13956 133598 14044
rect 133658 13958 133745 14046
rect 133838 13958 133925 14046
rect 133992 13959 134079 14047
rect 133331 13776 133418 13864
rect 133511 13776 133598 13864
rect 133658 13778 133745 13866
rect 133838 13778 133925 13866
rect 133992 13779 134079 13867
rect 135855 14153 135942 14241
rect 136035 14153 136122 14241
rect 136182 14155 136269 14243
rect 136362 14155 136449 14243
rect 136516 14156 136603 14244
rect 135837 13940 135924 14028
rect 136017 13940 136104 14028
rect 136164 13942 136251 14030
rect 136344 13942 136431 14030
rect 136498 13943 136585 14031
rect 135837 13760 135924 13848
rect 136017 13760 136104 13848
rect 136164 13762 136251 13850
rect 136344 13762 136431 13850
rect 136498 13763 136585 13851
rect 138571 14172 138658 14260
rect 138751 14172 138838 14260
rect 138898 14174 138985 14262
rect 139078 14174 139165 14262
rect 139232 14175 139319 14263
rect 138553 13959 138640 14047
rect 138733 13959 138820 14047
rect 138880 13961 138967 14049
rect 139060 13961 139147 14049
rect 139214 13962 139301 14050
rect 138553 13779 138640 13867
rect 138733 13779 138820 13867
rect 138880 13781 138967 13869
rect 139060 13781 139147 13869
rect 139214 13782 139301 13870
rect 15890 7141 15957 7207
rect 150342 6580 150429 6668
rect 150522 6580 150609 6668
rect 150669 6582 150756 6670
rect 150849 6582 150936 6670
rect 151003 6583 151090 6671
rect 150342 6400 150429 6488
rect 150522 6400 150609 6488
rect 150669 6402 150756 6490
rect 150849 6402 150936 6490
rect 151003 6403 151090 6491
rect 75648 5906 75735 5994
rect 75828 5906 75915 5994
rect 75975 5908 76062 5996
rect 76155 5908 76242 5996
rect 76309 5909 76396 5997
rect 76449 5908 76536 5996
rect 76590 5906 76677 5994
rect 75648 5726 75735 5814
rect 75828 5726 75915 5814
rect 75975 5728 76062 5816
rect 76155 5728 76242 5816
rect 76309 5729 76396 5817
rect 76449 5728 76536 5816
rect 76590 5726 76677 5814
rect 80919 5941 81006 6029
rect 81099 5941 81186 6029
rect 81246 5943 81333 6031
rect 81426 5943 81513 6031
rect 81580 5944 81667 6032
rect 81734 5945 81821 6033
rect 81882 5943 81969 6031
rect 80919 5761 81006 5849
rect 81099 5761 81186 5849
rect 81246 5763 81333 5851
rect 81426 5763 81513 5851
rect 81580 5764 81667 5852
rect 81734 5765 81821 5853
rect 81882 5763 81969 5851
rect 56847 4129 56934 4217
rect 57027 4129 57114 4217
rect 56847 3949 56934 4037
rect 57027 3949 57114 4037
rect 113837 3774 113924 3862
rect 114017 3774 114104 3862
rect 113837 3594 113924 3682
rect 114017 3594 114104 3682
rect 113839 3433 113926 3521
rect 114019 3433 114106 3521
rect 113839 3253 113926 3341
rect 114019 3253 114106 3341
rect 114475 3824 114562 3912
rect 114655 3824 114742 3912
rect 114475 3644 114562 3732
rect 114655 3644 114742 3732
rect 114473 3481 114560 3569
rect 114653 3481 114740 3569
rect 114473 3301 114560 3389
rect 114653 3301 114740 3389
rect 115082 3870 115169 3958
rect 115262 3870 115349 3958
rect 115082 3690 115169 3778
rect 115262 3690 115349 3778
rect 115082 3530 115169 3618
rect 115262 3530 115349 3618
rect 115082 3350 115169 3438
rect 115262 3350 115349 3438
rect 115729 3852 115816 3940
rect 115909 3852 115996 3940
rect 115729 3672 115816 3760
rect 115909 3672 115996 3760
rect 126226 4814 126313 4902
rect 126406 4814 126493 4902
rect 126226 4634 126313 4722
rect 126406 4634 126493 4722
rect 115732 3521 115819 3609
rect 115912 3521 115999 3609
rect 115732 3341 115819 3429
rect 115912 3341 115999 3429
rect 28075 589 28162 677
rect 28255 589 28342 677
rect 28402 591 28489 679
rect 28582 591 28669 679
rect 28736 592 28823 680
rect 28075 409 28162 497
rect 28255 409 28342 497
rect 28402 411 28489 499
rect 28582 411 28669 499
rect 28736 412 28823 500
rect 28057 196 28144 284
rect 28237 196 28324 284
rect 28384 198 28471 286
rect 28564 198 28651 286
rect 28718 199 28805 287
rect 28057 16 28144 104
rect 28237 16 28324 104
rect 28384 18 28471 106
rect 28564 18 28651 106
rect 28718 19 28805 107
rect 29881 636 29968 724
rect 30061 636 30148 724
rect 30208 638 30295 726
rect 30388 638 30475 726
rect 30542 639 30629 727
rect 29881 456 29968 544
rect 30061 456 30148 544
rect 30208 458 30295 546
rect 30388 458 30475 546
rect 30542 459 30629 547
rect 29887 248 29974 336
rect 30067 248 30154 336
rect 30214 250 30301 338
rect 30394 250 30481 338
rect 30548 251 30635 339
rect 29887 68 29974 156
rect 30067 68 30154 156
rect 30214 70 30301 158
rect 30394 70 30481 158
rect 30548 71 30635 159
rect 31618 636 31705 724
rect 31798 636 31885 724
rect 31945 638 32032 726
rect 32125 638 32212 726
rect 32279 639 32366 727
rect 31618 456 31705 544
rect 31798 456 31885 544
rect 31945 458 32032 546
rect 32125 458 32212 546
rect 32279 459 32366 547
rect 31630 248 31717 336
rect 31810 248 31897 336
rect 31957 250 32044 338
rect 32137 250 32224 338
rect 32291 251 32378 339
rect 31630 68 31717 156
rect 31810 68 31897 156
rect 31957 70 32044 158
rect 32137 70 32224 158
rect 32291 71 32378 159
rect 47846 810 47898 862
rect 47950 810 48002 862
rect 47846 706 47898 758
rect 47950 706 48002 758
rect 48410 699 48475 764
rect 48535 699 48600 764
rect 48660 699 48725 764
rect 48120 -676 48172 -624
rect 48224 -676 48276 -624
rect 48120 -780 48172 -728
rect 48224 -780 48276 -728
rect 48678 -683 48730 -631
rect 48782 -683 48834 -631
rect 48678 -787 48730 -735
rect 48782 -787 48834 -735
rect 662 -3401 714 -3349
rect 766 -3401 818 -3349
rect 870 -3401 922 -3349
rect 662 -3505 714 -3453
rect 766 -3505 818 -3453
rect 870 -3505 922 -3453
rect 662 -3609 714 -3557
rect 766 -3609 818 -3557
rect 870 -3609 922 -3557
rect 113912 2595 113974 2660
rect 114037 2595 114099 2660
rect 113912 2470 113974 2535
rect 114037 2470 114099 2535
rect 114458 2595 114520 2660
rect 114583 2595 114645 2660
rect 114458 2470 114520 2535
rect 114583 2470 114645 2535
rect 114986 2586 115048 2651
rect 115111 2586 115173 2651
rect 114986 2461 115048 2526
rect 115111 2461 115173 2526
rect 115535 2588 115597 2653
rect 115660 2588 115722 2653
rect 115535 2463 115597 2528
rect 115660 2463 115722 2528
rect 114184 1583 114247 1646
rect 114322 1581 114385 1644
rect 115006 1747 115069 1810
rect 115144 1745 115207 1808
rect 115977 -179 116029 -127
rect 116081 -179 116133 -127
rect 116185 -179 116237 -127
rect 116292 -177 116344 -125
rect 116396 -177 116448 -125
rect 116500 -177 116552 -125
rect 116607 -177 116659 -125
rect 116711 -177 116763 -125
rect 116815 -177 116867 -125
rect 115977 -283 116029 -231
rect 116081 -283 116133 -231
rect 116185 -283 116237 -231
rect 116292 -281 116344 -229
rect 116396 -281 116448 -229
rect 116500 -281 116552 -229
rect 116607 -281 116659 -229
rect 116711 -281 116763 -229
rect 116815 -281 116867 -229
rect 115977 -387 116029 -335
rect 116081 -387 116133 -335
rect 116185 -387 116237 -335
rect 116292 -385 116344 -333
rect 116396 -385 116448 -333
rect 116500 -385 116552 -333
rect 116607 -385 116659 -333
rect 116711 -385 116763 -333
rect 116815 -385 116867 -333
rect 16041 -6208 16108 -6142
rect 16045 -8550 16112 -8484
rect 16058 -9628 16125 -9562
rect 127145 214 127197 266
rect 127249 214 127301 266
rect 127353 214 127405 266
rect 127460 216 127512 268
rect 127564 216 127616 268
rect 127668 216 127720 268
rect 127775 216 127827 268
rect 127879 216 127931 268
rect 127983 216 128035 268
rect 127145 110 127197 162
rect 127249 110 127301 162
rect 127353 110 127405 162
rect 127460 112 127512 164
rect 127564 112 127616 164
rect 127668 112 127720 164
rect 127775 112 127827 164
rect 127879 112 127931 164
rect 127983 112 128035 164
rect 127145 6 127197 58
rect 127249 6 127301 58
rect 127353 6 127405 58
rect 127460 8 127512 60
rect 127564 8 127616 60
rect 127668 8 127720 60
rect 127775 8 127827 60
rect 127879 8 127931 60
rect 127983 8 128035 60
rect 121385 -3293 121437 -3241
rect 121489 -3293 121541 -3241
rect 121385 -3397 121437 -3345
rect 121489 -3397 121541 -3345
rect 121943 -3286 121995 -3234
rect 122047 -3286 122099 -3234
rect 121943 -3390 121995 -3338
rect 122047 -3390 122099 -3338
rect 122342 -3307 122406 -3240
rect 122474 -3312 122538 -3245
rect 122347 -3432 122411 -3365
rect 122472 -3431 122536 -3364
rect 121036 -3946 121102 -3880
rect 121167 -3943 121233 -3877
rect 121035 -4075 121101 -4009
rect 121169 -4075 121235 -4009
rect 121032 -4203 121098 -4137
rect 121167 -4203 121233 -4137
rect 121943 -4537 121995 -4485
rect 122047 -4537 122099 -4485
rect 121943 -4641 121995 -4589
rect 122047 -4641 122099 -4589
rect 122501 -4544 122553 -4492
rect 122605 -4544 122657 -4492
rect 122501 -4648 122553 -4596
rect 122605 -4648 122657 -4596
rect 145860 -8844 145912 -8792
rect 145964 -8844 146016 -8792
rect 146068 -8844 146120 -8792
rect 146201 -8844 146253 -8792
rect 146305 -8844 146357 -8792
rect 146409 -8844 146461 -8792
rect 145860 -8948 145912 -8896
rect 145964 -8948 146016 -8896
rect 146068 -8948 146120 -8896
rect 146201 -8948 146253 -8896
rect 146305 -8948 146357 -8896
rect 146409 -8948 146461 -8896
rect 145860 -9052 145912 -9000
rect 145964 -9052 146016 -9000
rect 146068 -9052 146120 -9000
rect 146201 -9052 146253 -9000
rect 146305 -9052 146357 -9000
rect 146409 -9052 146461 -9000
rect 75573 -14813 75660 -14725
rect 75733 -14813 75820 -14725
rect 75893 -14813 75980 -14725
rect 76053 -14813 76140 -14725
rect 76213 -14813 76300 -14725
rect 76373 -14813 76460 -14725
rect 133379 -13521 133466 -13433
rect 133559 -13521 133646 -13433
rect 133706 -13519 133793 -13431
rect 133886 -13519 133973 -13431
rect 134040 -13518 134127 -13430
rect 135817 -13526 135904 -13438
rect 135997 -13526 136084 -13438
rect 136144 -13524 136231 -13436
rect 136324 -13524 136411 -13436
rect 136478 -13523 136565 -13435
rect 138539 -13532 138626 -13444
rect 138719 -13532 138806 -13444
rect 138866 -13530 138953 -13442
rect 139046 -13530 139133 -13442
rect 139200 -13529 139287 -13441
rect 150321 -13499 150408 -13411
rect 150501 -13499 150588 -13411
rect 150648 -13497 150735 -13409
rect 150828 -13497 150915 -13409
rect 150982 -13496 151069 -13408
rect 133379 -13701 133466 -13613
rect 133559 -13701 133646 -13613
rect 133706 -13699 133793 -13611
rect 133886 -13699 133973 -13611
rect 134040 -13698 134127 -13610
rect 135817 -13706 135904 -13618
rect 135997 -13706 136084 -13618
rect 136144 -13704 136231 -13616
rect 136324 -13704 136411 -13616
rect 136478 -13703 136565 -13615
rect 138539 -13712 138626 -13624
rect 138719 -13712 138806 -13624
rect 138866 -13710 138953 -13622
rect 139046 -13710 139133 -13622
rect 139200 -13709 139287 -13621
rect 145840 -13656 145892 -13604
rect 145944 -13656 145996 -13604
rect 146048 -13656 146100 -13604
rect 146181 -13656 146233 -13604
rect 146285 -13656 146337 -13604
rect 146389 -13656 146441 -13604
rect 150321 -13679 150408 -13591
rect 150501 -13679 150588 -13591
rect 150648 -13677 150735 -13589
rect 150828 -13677 150915 -13589
rect 150982 -13676 151069 -13588
rect 145840 -13760 145892 -13708
rect 145944 -13760 145996 -13708
rect 146048 -13760 146100 -13708
rect 146181 -13760 146233 -13708
rect 146285 -13760 146337 -13708
rect 146389 -13760 146441 -13708
rect 133361 -13914 133448 -13826
rect 133541 -13914 133628 -13826
rect 133688 -13912 133775 -13824
rect 133868 -13912 133955 -13824
rect 134022 -13911 134109 -13823
rect 135799 -13919 135886 -13831
rect 135979 -13919 136066 -13831
rect 136126 -13917 136213 -13829
rect 136306 -13917 136393 -13829
rect 136460 -13916 136547 -13828
rect 138521 -13925 138608 -13837
rect 138701 -13925 138788 -13837
rect 138848 -13923 138935 -13835
rect 139028 -13923 139115 -13835
rect 139182 -13922 139269 -13834
rect 145840 -13864 145892 -13812
rect 145944 -13864 145996 -13812
rect 146048 -13864 146100 -13812
rect 146181 -13864 146233 -13812
rect 146285 -13864 146337 -13812
rect 146389 -13864 146441 -13812
rect 150303 -13892 150390 -13804
rect 150483 -13892 150570 -13804
rect 150630 -13890 150717 -13802
rect 150810 -13890 150897 -13802
rect 150964 -13889 151051 -13801
rect 133361 -14094 133448 -14006
rect 133541 -14094 133628 -14006
rect 133688 -14092 133775 -14004
rect 133868 -14092 133955 -14004
rect 134022 -14091 134109 -14003
rect 135799 -14099 135886 -14011
rect 135979 -14099 136066 -14011
rect 136126 -14097 136213 -14009
rect 136306 -14097 136393 -14009
rect 136460 -14096 136547 -14008
rect 138521 -14105 138608 -14017
rect 138701 -14105 138788 -14017
rect 138848 -14103 138935 -14015
rect 139028 -14103 139115 -14015
rect 139182 -14102 139269 -14014
rect 150303 -14072 150390 -13984
rect 150483 -14072 150570 -13984
rect 150630 -14070 150717 -13982
rect 150810 -14070 150897 -13982
rect 150964 -14069 151051 -13981
rect 75573 -14973 75660 -14885
rect 75733 -14973 75820 -14885
rect 75893 -14973 75980 -14885
rect 76053 -14973 76140 -14885
rect 76213 -14973 76300 -14885
rect 76373 -14973 76460 -14885
rect 80774 -15027 80861 -14939
rect 80954 -15027 81041 -14939
rect 81101 -15025 81188 -14937
rect 81281 -15025 81368 -14937
rect 81435 -15024 81522 -14936
rect 81605 -15027 81692 -14939
rect 81759 -15026 81846 -14938
rect 75573 -15133 75660 -15045
rect 75733 -15133 75820 -15045
rect 75893 -15133 75980 -15045
rect 76053 -15133 76140 -15045
rect 76213 -15133 76300 -15045
rect 76373 -15133 76460 -15045
rect 29831 -15449 29918 -15361
rect 29991 -15449 30078 -15361
rect 30151 -15449 30238 -15361
rect 30311 -15449 30398 -15361
rect 30471 -15449 30558 -15361
rect 30631 -15449 30718 -15361
rect 31543 -15363 31630 -15275
rect 31703 -15363 31790 -15275
rect 31863 -15363 31950 -15275
rect 32023 -15363 32110 -15275
rect 32183 -15363 32270 -15275
rect 32343 -15363 32430 -15275
rect 75573 -15293 75660 -15205
rect 75733 -15293 75820 -15205
rect 75893 -15293 75980 -15205
rect 76053 -15293 76140 -15205
rect 76213 -15293 76300 -15205
rect 76373 -15293 76460 -15205
rect 80774 -15207 80861 -15119
rect 80954 -15207 81041 -15119
rect 81101 -15205 81188 -15117
rect 81281 -15205 81368 -15117
rect 81435 -15204 81522 -15116
rect 81605 -15207 81692 -15119
rect 81759 -15206 81846 -15118
rect 28009 -15566 28096 -15478
rect 28169 -15566 28256 -15478
rect 28329 -15566 28416 -15478
rect 28489 -15566 28576 -15478
rect 28649 -15566 28736 -15478
rect 28809 -15566 28896 -15478
rect 28009 -15726 28096 -15638
rect 28169 -15726 28256 -15638
rect 28329 -15726 28416 -15638
rect 28489 -15726 28576 -15638
rect 28649 -15726 28736 -15638
rect 28809 -15726 28896 -15638
rect 28009 -15886 28096 -15798
rect 28169 -15886 28256 -15798
rect 28329 -15886 28416 -15798
rect 28489 -15886 28576 -15798
rect 28649 -15886 28736 -15798
rect 28809 -15886 28896 -15798
rect 28009 -16046 28096 -15958
rect 28169 -16046 28256 -15958
rect 28329 -16046 28416 -15958
rect 28489 -16046 28576 -15958
rect 28649 -16046 28736 -15958
rect 28809 -16046 28896 -15958
rect 29831 -15609 29918 -15521
rect 29991 -15609 30078 -15521
rect 30151 -15609 30238 -15521
rect 30311 -15609 30398 -15521
rect 30471 -15609 30558 -15521
rect 30631 -15609 30718 -15521
rect 31543 -15523 31630 -15435
rect 31703 -15523 31790 -15435
rect 31863 -15523 31950 -15435
rect 32023 -15523 32110 -15435
rect 32183 -15523 32270 -15435
rect 32343 -15523 32430 -15435
rect 75573 -15453 75660 -15365
rect 75733 -15453 75820 -15365
rect 75893 -15453 75980 -15365
rect 76053 -15453 76140 -15365
rect 76213 -15453 76300 -15365
rect 76373 -15453 76460 -15365
rect 80768 -15384 80855 -15296
rect 80948 -15384 81035 -15296
rect 81095 -15382 81182 -15294
rect 81275 -15382 81362 -15294
rect 81429 -15381 81516 -15293
rect 81599 -15384 81686 -15296
rect 81753 -15383 81840 -15295
rect 29831 -15769 29918 -15681
rect 29991 -15769 30078 -15681
rect 30151 -15769 30238 -15681
rect 30311 -15769 30398 -15681
rect 30471 -15769 30558 -15681
rect 30631 -15769 30718 -15681
rect 29831 -15929 29918 -15841
rect 29991 -15929 30078 -15841
rect 30151 -15929 30238 -15841
rect 30311 -15929 30398 -15841
rect 30471 -15929 30558 -15841
rect 30631 -15929 30718 -15841
rect 29831 -16089 29918 -16001
rect 29991 -16089 30078 -16001
rect 30151 -16089 30238 -16001
rect 30311 -16089 30398 -16001
rect 30471 -16089 30558 -16001
rect 30631 -16089 30718 -16001
rect 31543 -15683 31630 -15595
rect 31703 -15683 31790 -15595
rect 31863 -15683 31950 -15595
rect 32023 -15683 32110 -15595
rect 32183 -15683 32270 -15595
rect 32343 -15683 32430 -15595
rect 31543 -15843 31630 -15755
rect 31703 -15843 31790 -15755
rect 31863 -15843 31950 -15755
rect 32023 -15843 32110 -15755
rect 32183 -15843 32270 -15755
rect 32343 -15843 32430 -15755
rect 31543 -16003 31630 -15915
rect 31703 -16003 31790 -15915
rect 31863 -16003 31950 -15915
rect 32023 -16003 32110 -15915
rect 32183 -16003 32270 -15915
rect 32343 -16003 32430 -15915
rect 28009 -16206 28096 -16118
rect 28169 -16206 28256 -16118
rect 28329 -16206 28416 -16118
rect 28489 -16206 28576 -16118
rect 28649 -16206 28736 -16118
rect 28809 -16206 28896 -16118
rect 29831 -16249 29918 -16161
rect 29991 -16249 30078 -16161
rect 30151 -16249 30238 -16161
rect 30311 -16249 30398 -16161
rect 30471 -16249 30558 -16161
rect 30631 -16249 30718 -16161
rect 31543 -16163 31630 -16075
rect 31703 -16163 31790 -16075
rect 31863 -16163 31950 -16075
rect 32023 -16163 32110 -16075
rect 32183 -16163 32270 -16075
rect 32343 -16163 32430 -16075
rect 75573 -15613 75660 -15525
rect 75733 -15613 75820 -15525
rect 75893 -15613 75980 -15525
rect 76053 -15613 76140 -15525
rect 76213 -15613 76300 -15525
rect 76373 -15613 76460 -15525
rect 80884 -16053 80971 -15965
rect 81044 -16053 81131 -15965
rect 81204 -16053 81291 -15965
rect 81364 -16053 81451 -15965
rect 81524 -16053 81611 -15965
rect 81684 -16053 81771 -15965
rect 80884 -16213 80971 -16125
rect 81044 -16213 81131 -16125
rect 81204 -16213 81291 -16125
rect 81364 -16213 81451 -16125
rect 81524 -16213 81611 -16125
rect 81684 -16213 81771 -16125
rect 28009 -16366 28096 -16278
rect 28169 -16366 28256 -16278
rect 28329 -16366 28416 -16278
rect 28489 -16366 28576 -16278
rect 28649 -16366 28736 -16278
rect 28809 -16366 28896 -16278
rect 75652 -16355 75739 -16267
rect 75832 -16355 75919 -16267
rect 75979 -16353 76066 -16265
rect 76159 -16353 76246 -16265
rect 76313 -16352 76400 -16264
rect 76483 -16355 76570 -16267
rect 76637 -16354 76724 -16266
rect 80884 -16373 80971 -16285
rect 81044 -16373 81131 -16285
rect 81204 -16373 81291 -16285
rect 81364 -16373 81451 -16285
rect 81524 -16373 81611 -16285
rect 81684 -16373 81771 -16285
rect 75652 -16535 75739 -16447
rect 75832 -16535 75919 -16447
rect 75979 -16533 76066 -16445
rect 76159 -16533 76246 -16445
rect 76313 -16532 76400 -16444
rect 76483 -16535 76570 -16447
rect 76637 -16534 76724 -16446
rect 80884 -16533 80971 -16445
rect 81044 -16533 81131 -16445
rect 81204 -16533 81291 -16445
rect 81364 -16533 81451 -16445
rect 81524 -16533 81611 -16445
rect 81684 -16533 81771 -16445
rect 75646 -16712 75733 -16624
rect 75826 -16712 75913 -16624
rect 75973 -16710 76060 -16622
rect 76153 -16710 76240 -16622
rect 76307 -16709 76394 -16621
rect 76477 -16712 76564 -16624
rect 76631 -16711 76718 -16623
rect 80884 -16693 80971 -16605
rect 81044 -16693 81131 -16605
rect 81204 -16693 81291 -16605
rect 81364 -16693 81451 -16605
rect 81524 -16693 81611 -16605
rect 81684 -16693 81771 -16605
rect 80884 -16853 80971 -16765
rect 81044 -16853 81131 -16765
rect 81204 -16853 81291 -16765
rect 81364 -16853 81451 -16765
rect 81524 -16853 81611 -16765
rect 81684 -16853 81771 -16765
rect 27290 -18251 27377 -18163
rect 27450 -18251 27537 -18163
rect 27610 -18251 27697 -18163
rect 27770 -18251 27857 -18163
rect 27930 -18251 28017 -18163
rect 28090 -18251 28177 -18163
rect 312 -18432 395 -18349
rect 482 -18432 565 -18349
rect 652 -18432 735 -18349
rect 822 -18432 905 -18349
rect 992 -18432 1075 -18349
rect 312 -18602 395 -18519
rect 482 -18602 565 -18519
rect 652 -18602 735 -18519
rect 822 -18602 905 -18519
rect 992 -18602 1075 -18519
rect 312 -18772 395 -18689
rect 482 -18772 565 -18689
rect 652 -18772 735 -18689
rect 822 -18772 905 -18689
rect 992 -18772 1075 -18689
rect 312 -18942 395 -18859
rect 482 -18942 565 -18859
rect 652 -18942 735 -18859
rect 822 -18942 905 -18859
rect 992 -18942 1075 -18859
rect 312 -19112 395 -19029
rect 482 -19112 565 -19029
rect 652 -19112 735 -19029
rect 822 -19112 905 -19029
rect 992 -19112 1075 -19029
rect 27290 -18411 27377 -18323
rect 27450 -18411 27537 -18323
rect 27610 -18411 27697 -18323
rect 27770 -18411 27857 -18323
rect 27930 -18411 28017 -18323
rect 28090 -18411 28177 -18323
rect 27290 -18571 27377 -18483
rect 27450 -18571 27537 -18483
rect 27610 -18571 27697 -18483
rect 27770 -18571 27857 -18483
rect 27930 -18571 28017 -18483
rect 28090 -18571 28177 -18483
rect 27290 -18731 27377 -18643
rect 27450 -18731 27537 -18643
rect 27610 -18731 27697 -18643
rect 27770 -18731 27857 -18643
rect 27930 -18731 28017 -18643
rect 28090 -18731 28177 -18643
rect 27290 -18891 27377 -18803
rect 27450 -18891 27537 -18803
rect 27610 -18891 27697 -18803
rect 27770 -18891 27857 -18803
rect 27930 -18891 28017 -18803
rect 28090 -18891 28177 -18803
rect 27290 -19051 27377 -18963
rect 27450 -19051 27537 -18963
rect 27610 -19051 27697 -18963
rect 27770 -19051 27857 -18963
rect 27930 -19051 28017 -18963
rect 28090 -19051 28177 -18963
rect 27933 -19537 28020 -19449
rect 28113 -19537 28200 -19449
rect 28260 -19535 28347 -19447
rect 28440 -19535 28527 -19447
rect 28594 -19534 28681 -19446
<< metal2 >>
rect 1898 17585 2709 17608
rect 1898 17502 1922 17585
rect 2005 17502 2092 17585
rect 2175 17502 2262 17585
rect 2345 17502 2432 17585
rect 2515 17502 2602 17585
rect 2685 17502 2709 17585
rect 1898 17415 2709 17502
rect 1898 17332 1922 17415
rect 2005 17332 2092 17415
rect 2175 17332 2262 17415
rect 2345 17332 2432 17415
rect 2515 17332 2602 17415
rect 2685 17332 2709 17415
rect 1898 17245 2709 17332
rect 1898 17162 1922 17245
rect 2005 17162 2092 17245
rect 2175 17162 2262 17245
rect 2345 17162 2432 17245
rect 2515 17162 2602 17245
rect 2685 17162 2709 17245
rect 1898 17075 2709 17162
rect 1898 16992 1922 17075
rect 2005 16992 2092 17075
rect 2175 16992 2262 17075
rect 2345 16992 2432 17075
rect 2515 16992 2602 17075
rect 2685 16992 2709 17075
rect 1898 16905 2709 16992
rect 1898 16822 1922 16905
rect 2005 16822 2092 16905
rect 2175 16822 2262 16905
rect 2345 16822 2432 16905
rect 2515 16822 2602 16905
rect 2685 16822 2709 16905
rect 1898 16799 2709 16822
rect 4041 17567 4852 17590
rect 4041 17484 4065 17567
rect 4148 17484 4235 17567
rect 4318 17484 4405 17567
rect 4488 17484 4575 17567
rect 4658 17484 4745 17567
rect 4828 17484 4852 17567
rect 4041 17397 4852 17484
rect 4041 17314 4065 17397
rect 4148 17314 4235 17397
rect 4318 17314 4405 17397
rect 4488 17314 4575 17397
rect 4658 17314 4745 17397
rect 4828 17314 4852 17397
rect 4041 17227 4852 17314
rect 85623 17368 86434 17391
rect 4041 17144 4065 17227
rect 4148 17144 4235 17227
rect 4318 17144 4405 17227
rect 4488 17144 4575 17227
rect 4658 17144 4745 17227
rect 4828 17144 4852 17227
rect 4041 17057 4852 17144
rect 4041 16974 4065 17057
rect 4148 16974 4235 17057
rect 4318 16974 4405 17057
rect 4488 16974 4575 17057
rect 4658 16974 4745 17057
rect 4828 16974 4852 17057
rect 4041 16887 4852 16974
rect 4041 16804 4065 16887
rect 4148 16804 4235 16887
rect 4318 16804 4405 16887
rect 4488 16804 4575 16887
rect 4658 16804 4745 16887
rect 4828 16804 4852 16887
rect -608 15781 -319 15799
rect -608 15725 -597 15781
rect -541 15725 -493 15781
rect -437 15725 -389 15781
rect -333 15743 -319 15781
rect 2186 15743 2404 16799
rect 4041 16781 4852 16804
rect 17976 17285 18787 17308
rect 17976 17202 18000 17285
rect 18083 17202 18170 17285
rect 18253 17202 18340 17285
rect 18423 17202 18510 17285
rect 18593 17202 18680 17285
rect 18763 17202 18787 17285
rect 85623 17285 85647 17368
rect 85730 17285 85817 17368
rect 85900 17285 85987 17368
rect 86070 17285 86157 17368
rect 86240 17285 86327 17368
rect 86410 17285 86434 17368
rect 17976 17115 18787 17202
rect 17976 17032 18000 17115
rect 18083 17032 18170 17115
rect 18253 17032 18340 17115
rect 18423 17032 18510 17115
rect 18593 17032 18680 17115
rect 18763 17032 18787 17115
rect 17976 16945 18787 17032
rect 17976 16862 18000 16945
rect 18083 16862 18170 16945
rect 18253 16862 18340 16945
rect 18423 16862 18510 16945
rect 18593 16862 18680 16945
rect 18763 16862 18787 16945
rect -333 15725 2404 15743
rect -4959 15658 -4150 15682
rect -4959 15575 -4936 15658
rect -4853 15575 -4766 15658
rect -4683 15575 -4596 15658
rect -4513 15575 -4426 15658
rect -4343 15575 -4256 15658
rect -4173 15575 -4150 15658
rect -4959 15488 -4150 15575
rect -608 15677 2404 15725
rect -608 15621 -597 15677
rect -541 15621 -493 15677
rect -437 15621 -389 15677
rect -333 15621 2404 15677
rect -608 15573 2404 15621
rect -608 15517 -597 15573
rect -541 15517 -493 15573
rect -437 15517 -389 15573
rect -333 15525 2404 15573
rect -333 15517 -319 15525
rect -608 15505 -319 15517
rect -4959 15405 -4936 15488
rect -4853 15405 -4766 15488
rect -4683 15405 -4596 15488
rect -4513 15405 -4426 15488
rect -4343 15405 -4256 15488
rect -4173 15405 -4150 15488
rect -4959 15318 -4150 15405
rect -172 15352 117 15370
rect -4959 15235 -4936 15318
rect -4853 15235 -4766 15318
rect -4683 15235 -4596 15318
rect -4513 15235 -4426 15318
rect -4343 15235 -4256 15318
rect -4173 15314 -4150 15318
rect -3549 15314 -3260 15322
rect -4173 15304 -3260 15314
rect -4173 15248 -3538 15304
rect -3482 15248 -3434 15304
rect -3378 15248 -3330 15304
rect -3274 15248 -3260 15304
rect -4173 15235 -3260 15248
rect -4959 15200 -3260 15235
rect -4959 15148 -3538 15200
rect -4959 15065 -4936 15148
rect -4853 15065 -4766 15148
rect -4683 15065 -4596 15148
rect -4513 15065 -4426 15148
rect -4343 15065 -4256 15148
rect -4173 15144 -3538 15148
rect -3482 15144 -3434 15200
rect -3378 15144 -3330 15200
rect -3274 15144 -3260 15200
rect -4173 15096 -3260 15144
rect -4173 15065 -3538 15096
rect -4959 15056 -3538 15065
rect -4959 14978 -4150 15056
rect -3549 15040 -3538 15056
rect -3482 15040 -3434 15096
rect -3378 15040 -3330 15096
rect -3274 15040 -3260 15096
rect -172 15296 -161 15352
rect -105 15296 -57 15352
rect -1 15296 47 15352
rect 103 15316 117 15352
rect 4392 15316 4610 16781
rect 17976 16775 18787 16862
rect 17976 16692 18000 16775
rect 18083 16692 18170 16775
rect 18253 16692 18340 16775
rect 18423 16692 18510 16775
rect 18593 16692 18680 16775
rect 18763 16692 18787 16775
rect 17976 16605 18787 16692
rect 17976 16522 18000 16605
rect 18083 16522 18170 16605
rect 18253 16522 18340 16605
rect 18423 16522 18510 16605
rect 18593 16522 18680 16605
rect 18763 16522 18787 16605
rect 17976 16499 18787 16522
rect 21980 17221 22791 17244
rect 21980 17138 22004 17221
rect 22087 17138 22174 17221
rect 22257 17138 22344 17221
rect 22427 17138 22514 17221
rect 22597 17138 22684 17221
rect 22767 17138 22791 17221
rect 21980 17051 22791 17138
rect 21980 16968 22004 17051
rect 22087 16968 22174 17051
rect 22257 16968 22344 17051
rect 22427 16968 22514 17051
rect 22597 16968 22684 17051
rect 22767 16968 22791 17051
rect 21980 16881 22791 16968
rect 21980 16798 22004 16881
rect 22087 16798 22174 16881
rect 22257 16798 22344 16881
rect 22427 16798 22514 16881
rect 22597 16798 22684 16881
rect 22767 16798 22791 16881
rect 21980 16711 22791 16798
rect 21980 16628 22004 16711
rect 22087 16628 22174 16711
rect 22257 16628 22344 16711
rect 22427 16628 22514 16711
rect 22597 16628 22684 16711
rect 22767 16628 22791 16711
rect 21980 16541 22791 16628
rect 85623 17198 86434 17285
rect 85623 17115 85647 17198
rect 85730 17115 85817 17198
rect 85900 17115 85987 17198
rect 86070 17115 86157 17198
rect 86240 17115 86327 17198
rect 86410 17115 86434 17198
rect 85623 17028 86434 17115
rect 85623 16945 85647 17028
rect 85730 16945 85817 17028
rect 85900 16945 85987 17028
rect 86070 16945 86157 17028
rect 86240 16945 86327 17028
rect 86410 16945 86434 17028
rect 85623 16858 86434 16945
rect 85623 16775 85647 16858
rect 85730 16775 85817 16858
rect 85900 16775 85987 16858
rect 86070 16775 86157 16858
rect 86240 16775 86327 16858
rect 86410 16775 86434 16858
rect 85623 16688 86434 16775
rect 85623 16605 85647 16688
rect 85730 16605 85817 16688
rect 85900 16605 85987 16688
rect 86070 16605 86157 16688
rect 86240 16605 86327 16688
rect 86410 16605 86434 16688
rect 85623 16582 86434 16605
rect 89240 17359 90051 17382
rect 89240 17276 89264 17359
rect 89347 17276 89434 17359
rect 89517 17276 89604 17359
rect 89687 17276 89774 17359
rect 89857 17276 89944 17359
rect 90027 17276 90051 17359
rect 89240 17189 90051 17276
rect 89240 17106 89264 17189
rect 89347 17106 89434 17189
rect 89517 17106 89604 17189
rect 89687 17106 89774 17189
rect 89857 17106 89944 17189
rect 90027 17106 90051 17189
rect 89240 17019 90051 17106
rect 89240 16936 89264 17019
rect 89347 16936 89434 17019
rect 89517 16936 89604 17019
rect 89687 16936 89774 17019
rect 89857 16936 89944 17019
rect 90027 16936 90051 17019
rect 89240 16849 90051 16936
rect 89240 16766 89264 16849
rect 89347 16766 89434 16849
rect 89517 16766 89604 16849
rect 89687 16766 89774 16849
rect 89857 16766 89944 16849
rect 90027 16766 90051 16849
rect 89240 16679 90051 16766
rect 89240 16596 89264 16679
rect 89347 16596 89434 16679
rect 89517 16596 89604 16679
rect 89687 16596 89774 16679
rect 89857 16596 89944 16679
rect 90027 16596 90051 16679
rect 103 15296 4610 15316
rect -172 15248 4610 15296
rect -172 15192 -161 15248
rect -105 15192 -57 15248
rect -1 15192 47 15248
rect 103 15192 4610 15248
rect -172 15144 4610 15192
rect -172 15088 -161 15144
rect -105 15088 -57 15144
rect -1 15088 47 15144
rect 103 15098 4610 15144
rect 103 15088 117 15098
rect -172 15076 117 15088
rect -3549 15028 -3260 15040
rect -4959 14895 -4936 14978
rect -4853 14895 -4766 14978
rect -4683 14895 -4596 14978
rect -4513 14895 -4426 14978
rect -4343 14895 -4256 14978
rect -4173 14895 -4150 14978
rect -4959 14871 -4150 14895
rect -2468 14747 852 14766
rect -2486 14729 852 14747
rect -2486 14673 -2475 14729
rect -2419 14673 -2371 14729
rect -2315 14673 -2267 14729
rect -2211 14673 852 14729
rect -2486 14625 852 14673
rect -2486 14569 -2475 14625
rect -2419 14569 -2371 14625
rect -2315 14569 -2267 14625
rect -2211 14569 852 14625
rect -2486 14521 852 14569
rect -2486 14465 -2475 14521
rect -2419 14465 -2371 14521
rect -2315 14465 -2267 14521
rect -2211 14465 852 14521
rect -2486 14453 852 14465
rect -2468 14448 852 14453
rect -3026 14328 -2737 14346
rect -3026 14272 -3015 14328
rect -2959 14272 -2911 14328
rect -2855 14272 -2807 14328
rect -2751 14292 -2737 14328
rect -2751 14272 310 14292
rect -3026 14224 310 14272
rect -3026 14168 -3015 14224
rect -2959 14168 -2911 14224
rect -2855 14168 -2807 14224
rect -2751 14168 310 14224
rect -3026 14120 310 14168
rect 514 14276 852 14448
rect 514 14166 964 14276
rect -3026 14064 -3015 14120
rect -2959 14064 -2911 14120
rect -2855 14064 -2807 14120
rect -2751 14076 310 14120
rect -2751 14067 1013 14076
rect -2751 14064 -2737 14067
rect -3026 14052 -2737 14064
rect 154 13966 1013 14067
rect -1051 13919 -762 13937
rect -1051 13863 -1040 13919
rect -984 13863 -936 13919
rect -880 13863 -832 13919
rect -776 13876 -762 13919
rect -776 13863 964 13876
rect -1051 13815 964 13863
rect -1051 13759 -1040 13815
rect -984 13759 -936 13815
rect -880 13759 -832 13815
rect -776 13766 964 13815
rect -776 13759 -762 13766
rect -1051 13711 -762 13759
rect -1051 13655 -1040 13711
rect -984 13655 -936 13711
rect -880 13655 -832 13711
rect -776 13655 -762 13711
rect -1051 13643 -762 13655
rect 210 13566 1067 13676
rect -1455 13365 -1166 13383
rect -1455 13309 -1444 13365
rect -1388 13309 -1340 13365
rect -1284 13309 -1236 13365
rect -1180 13337 -1166 13365
rect 210 13337 320 13566
rect -1180 13309 320 13337
rect -1455 13261 320 13309
rect -1455 13205 -1444 13261
rect -1388 13205 -1340 13261
rect -1284 13205 -1236 13261
rect -1180 13205 320 13261
rect -1455 13157 320 13205
rect -1455 13101 -1444 13157
rect -1388 13101 -1340 13157
rect -1284 13101 -1236 13157
rect -1180 13146 320 13157
rect 580 13370 1186 13401
rect 580 13318 599 13370
rect 651 13318 703 13370
rect 755 13318 807 13370
rect 859 13318 1186 13370
rect 580 13303 1186 13318
rect 580 13266 871 13303
rect 580 13214 599 13266
rect 651 13214 703 13266
rect 755 13214 807 13266
rect 859 13214 871 13266
rect 580 13162 871 13214
rect -1180 13101 -1166 13146
rect -1455 13089 -1166 13101
rect 580 13110 599 13162
rect 651 13110 703 13162
rect 755 13110 807 13162
rect 859 13110 871 13162
rect 580 13100 871 13110
rect 587 13098 871 13100
rect -4976 12724 -4167 12748
rect -4976 12641 -4953 12724
rect -4870 12641 -4783 12724
rect -4700 12641 -4613 12724
rect -4530 12641 -4443 12724
rect -4360 12641 -4273 12724
rect -4190 12641 -4167 12724
rect -4976 12554 -4167 12641
rect -4976 12471 -4953 12554
rect -4870 12471 -4783 12554
rect -4700 12471 -4613 12554
rect -4530 12471 -4443 12554
rect -4360 12471 -4273 12554
rect -4190 12471 -4167 12554
rect -4976 12400 -4167 12471
rect -3003 12400 -2714 12406
rect -4976 12388 -2714 12400
rect -4976 12384 -2992 12388
rect -4976 12301 -4953 12384
rect -4870 12301 -4783 12384
rect -4700 12301 -4613 12384
rect -4530 12301 -4443 12384
rect -4360 12301 -4273 12384
rect -4190 12332 -2992 12384
rect -2936 12332 -2888 12388
rect -2832 12332 -2784 12388
rect -2728 12332 -2714 12388
rect -4190 12301 -2714 12332
rect -4976 12284 -2714 12301
rect -4976 12228 -2992 12284
rect -2936 12228 -2888 12284
rect -2832 12228 -2784 12284
rect -2728 12228 -2714 12284
rect -4976 12214 -2714 12228
rect -4976 12131 -4953 12214
rect -4870 12131 -4783 12214
rect -4700 12131 -4613 12214
rect -4530 12131 -4443 12214
rect -4360 12131 -4273 12214
rect -4190 12180 -2714 12214
rect -4190 12142 -2992 12180
rect -4190 12131 -4167 12142
rect -4976 12044 -4167 12131
rect -3003 12124 -2992 12142
rect -2936 12124 -2888 12180
rect -2832 12124 -2784 12180
rect -2728 12124 -2714 12180
rect -3003 12112 -2714 12124
rect -4976 11961 -4953 12044
rect -4870 11961 -4783 12044
rect -4700 11961 -4613 12044
rect -4530 11961 -4443 12044
rect -4360 11961 -4273 12044
rect -4190 11961 -4167 12044
rect -4976 11937 -4167 11961
rect -1970 11839 1053 11870
rect -1970 11834 527 11839
rect -1970 11778 -1957 11834
rect -1901 11778 -1853 11834
rect -1797 11778 -1749 11834
rect -1693 11783 527 11834
rect 583 11783 631 11839
rect 687 11783 735 11839
rect 791 11783 1053 11839
rect -1693 11778 1053 11783
rect -1970 11735 1053 11778
rect -1970 11730 527 11735
rect -1970 11674 -1957 11730
rect -1901 11674 -1853 11730
rect -1797 11674 -1749 11730
rect -1693 11679 527 11730
rect 583 11679 631 11735
rect 687 11679 735 11735
rect 791 11679 1053 11735
rect -1693 11674 1053 11679
rect -1970 11631 1053 11674
rect -1970 11626 527 11631
rect -1970 11570 -1957 11626
rect -1901 11570 -1853 11626
rect -1797 11570 -1749 11626
rect -1693 11575 527 11626
rect 583 11575 631 11631
rect 687 11575 735 11631
rect 791 11575 1053 11631
rect -1693 11570 1053 11575
rect -1970 11552 1053 11570
rect 15882 10624 15981 10640
rect 15882 10558 15899 10624
rect 15966 10558 15981 10624
rect 15882 10542 15981 10558
rect 16441 10609 16670 11694
rect 16441 10543 16529 10609
rect 16596 10543 16670 10609
rect -4976 9352 -4167 9376
rect -4976 9269 -4953 9352
rect -4870 9269 -4783 9352
rect -4700 9269 -4613 9352
rect -4530 9269 -4443 9352
rect -4360 9269 -4273 9352
rect -4190 9269 -4167 9352
rect -4976 9182 -4167 9269
rect -4976 9099 -4953 9182
rect -4870 9099 -4783 9182
rect -4700 9099 -4613 9182
rect -4530 9099 -4443 9182
rect -4360 9099 -4273 9182
rect -4190 9099 -4167 9182
rect -4976 9085 -4167 9099
rect -2981 9085 -2692 9101
rect -4976 9083 -2692 9085
rect -4976 9027 -2970 9083
rect -2914 9027 -2866 9083
rect -2810 9027 -2762 9083
rect -2706 9027 -2692 9083
rect -4976 9012 -2692 9027
rect -4976 8929 -4953 9012
rect -4870 8929 -4783 9012
rect -4700 8929 -4613 9012
rect -4530 8929 -4443 9012
rect -4360 8929 -4273 9012
rect -4190 8979 -2692 9012
rect -4190 8929 -2970 8979
rect -4976 8923 -2970 8929
rect -2914 8923 -2866 8979
rect -2810 8923 -2762 8979
rect -2706 8923 -2692 8979
rect -4976 8875 -2692 8923
rect -4976 8842 -2970 8875
rect -4976 8759 -4953 8842
rect -4870 8759 -4783 8842
rect -4700 8759 -4613 8842
rect -4530 8759 -4443 8842
rect -4360 8759 -4273 8842
rect -4190 8827 -2970 8842
rect -4190 8759 -4167 8827
rect -2981 8819 -2970 8827
rect -2914 8819 -2866 8875
rect -2810 8819 -2762 8875
rect -2706 8819 -2692 8875
rect -2981 8807 -2692 8819
rect -4976 8672 -4167 8759
rect -4976 8589 -4953 8672
rect -4870 8589 -4783 8672
rect -4700 8589 -4613 8672
rect -4530 8589 -4443 8672
rect -4360 8589 -4273 8672
rect -4190 8589 -4167 8672
rect -4976 8565 -4167 8589
rect 15870 8288 15969 8304
rect 15870 8222 15887 8288
rect 15954 8222 15969 8288
rect 15870 8206 15969 8222
rect 15873 7207 15972 7223
rect 15873 7141 15890 7207
rect 15957 7141 15972 7207
rect 15873 7125 15972 7141
rect -5044 7042 -4235 7066
rect -5044 6959 -5021 7042
rect -4938 6959 -4851 7042
rect -4768 6959 -4681 7042
rect -4598 6959 -4511 7042
rect -4428 6959 -4341 7042
rect -4258 6959 -4235 7042
rect -5044 6872 -4235 6959
rect -5044 6789 -5021 6872
rect -4938 6789 -4851 6872
rect -4768 6789 -4681 6872
rect -4598 6789 -4511 6872
rect -4428 6789 -4341 6872
rect -4258 6817 -4235 6872
rect -4258 6789 958 6817
rect -5044 6787 958 6789
rect -5044 6731 614 6787
rect 670 6731 718 6787
rect 774 6731 822 6787
rect 878 6731 958 6787
rect -5044 6702 958 6731
rect -5044 6619 -5021 6702
rect -4938 6619 -4851 6702
rect -4768 6619 -4681 6702
rect -4598 6619 -4511 6702
rect -4428 6619 -4341 6702
rect -4258 6683 958 6702
rect -4258 6627 614 6683
rect 670 6627 718 6683
rect 774 6627 822 6683
rect 878 6627 958 6683
rect -4258 6619 958 6627
rect -5044 6579 958 6619
rect -5044 6532 614 6579
rect -5044 6449 -5021 6532
rect -4938 6449 -4851 6532
rect -4768 6449 -4681 6532
rect -4598 6449 -4511 6532
rect -4428 6449 -4341 6532
rect -4258 6523 614 6532
rect 670 6523 718 6579
rect 774 6523 822 6579
rect 878 6523 958 6579
rect -4258 6502 958 6523
rect -4258 6449 -4235 6502
rect -5044 6362 -4235 6449
rect -5044 6279 -5021 6362
rect -4938 6279 -4851 6362
rect -4768 6279 -4681 6362
rect -4598 6279 -4511 6362
rect -4428 6279 -4341 6362
rect -4258 6279 -4235 6362
rect -5044 6255 -4235 6279
rect -5027 5290 -4218 5314
rect -5027 5207 -5004 5290
rect -4921 5207 -4834 5290
rect -4751 5207 -4664 5290
rect -4581 5207 -4494 5290
rect -4411 5207 -4324 5290
rect -4241 5207 -4218 5290
rect -5027 5120 -4218 5207
rect -5027 5037 -5004 5120
rect -4921 5037 -4834 5120
rect -4751 5037 -4664 5120
rect -4581 5037 -4494 5120
rect -4411 5037 -4324 5120
rect -4241 5037 -4218 5120
rect -5027 4981 -4218 5037
rect -5027 4968 -2217 4981
rect -5027 4950 -2192 4968
rect -5027 4867 -5004 4950
rect -4921 4867 -4834 4950
rect -4751 4867 -4664 4950
rect -4581 4867 -4494 4950
rect -4411 4867 -4324 4950
rect -4241 4894 -2470 4950
rect -2414 4894 -2366 4950
rect -2310 4894 -2262 4950
rect -2206 4894 -2192 4950
rect -4241 4867 -2192 4894
rect -5027 4846 -2192 4867
rect -5027 4790 -2470 4846
rect -2414 4790 -2366 4846
rect -2310 4790 -2262 4846
rect -2206 4790 -2192 4846
rect -5027 4780 -2192 4790
rect -5027 4697 -5004 4780
rect -4921 4697 -4834 4780
rect -4751 4697 -4664 4780
rect -4581 4697 -4494 4780
rect -4411 4697 -4324 4780
rect -4241 4742 -2192 4780
rect -4241 4697 -2470 4742
rect -5027 4686 -2470 4697
rect -2414 4686 -2366 4742
rect -2310 4686 -2262 4742
rect -2206 4686 -2192 4742
rect -5027 4674 -2192 4686
rect -5027 4666 -2217 4674
rect -5027 4610 -4218 4666
rect -5027 4527 -5004 4610
rect -4921 4527 -4834 4610
rect -4751 4527 -4664 4610
rect -4581 4527 -4494 4610
rect -4411 4527 -4324 4610
rect -4241 4527 -4218 4610
rect -5027 4503 -4218 4527
rect -5178 2777 -4369 2801
rect -5178 2694 -5155 2777
rect -5072 2694 -4985 2777
rect -4902 2694 -4815 2777
rect -4732 2694 -4645 2777
rect -4562 2694 -4475 2777
rect -4392 2694 -4369 2777
rect -5178 2607 -4369 2694
rect -5178 2524 -5155 2607
rect -5072 2524 -4985 2607
rect -4902 2524 -4815 2607
rect -4732 2524 -4645 2607
rect -4562 2524 -4475 2607
rect -4392 2524 -4369 2607
rect -5178 2486 -4369 2524
rect -5178 2470 108 2486
rect -5178 2452 113 2470
rect -5178 2437 -165 2452
rect -5178 2354 -5155 2437
rect -5072 2354 -4985 2437
rect -4902 2354 -4815 2437
rect -4732 2354 -4645 2437
rect -4562 2354 -4475 2437
rect -4392 2396 -165 2437
rect -109 2396 -61 2452
rect -5 2396 43 2452
rect 99 2396 113 2452
rect -4392 2354 113 2396
rect -5178 2348 113 2354
rect -5178 2292 -165 2348
rect -109 2292 -61 2348
rect -5 2292 43 2348
rect 99 2292 113 2348
rect -5178 2267 113 2292
rect -5178 2184 -5155 2267
rect -5072 2184 -4985 2267
rect -4902 2184 -4815 2267
rect -4732 2184 -4645 2267
rect -4562 2184 -4475 2267
rect -4392 2244 113 2267
rect -4392 2188 -165 2244
rect -109 2188 -61 2244
rect -5 2188 43 2244
rect 99 2188 113 2244
rect -4392 2184 113 2188
rect -5178 2176 113 2184
rect -5178 2171 108 2176
rect -5178 2097 -4369 2171
rect -5178 2014 -5155 2097
rect -5072 2014 -4985 2097
rect -4902 2014 -4815 2097
rect -4732 2014 -4645 2097
rect -4562 2014 -4475 2097
rect -4392 2014 -4369 2097
rect -5178 1990 -4369 2014
rect -2472 1074 922 1082
rect -2481 1057 922 1074
rect -2481 1056 943 1057
rect -2481 1000 -2470 1056
rect -2414 1000 -2366 1056
rect -2310 1000 -2262 1056
rect -2206 1039 943 1056
rect -2206 1000 665 1039
rect -2481 983 665 1000
rect 721 983 769 1039
rect 825 983 873 1039
rect 929 983 943 1039
rect -2481 952 943 983
rect -2481 896 -2470 952
rect -2414 896 -2366 952
rect -2310 896 -2262 952
rect -2206 935 943 952
rect -2206 896 665 935
rect -2481 879 665 896
rect 721 879 769 935
rect 825 879 873 935
rect 929 879 943 935
rect -2481 848 943 879
rect -2481 792 -2470 848
rect -2414 792 -2366 848
rect -2310 792 -2262 848
rect -2206 831 943 848
rect -2206 792 665 831
rect -2481 780 665 792
rect -2472 775 665 780
rect 721 775 769 831
rect 825 775 873 831
rect 929 775 943 831
rect -2472 767 943 775
rect 654 763 943 767
rect -5178 -1641 -4369 -1617
rect -5178 -1724 -5155 -1641
rect -5072 -1724 -4985 -1641
rect -4902 -1724 -4815 -1641
rect -4732 -1724 -4645 -1641
rect -4562 -1724 -4475 -1641
rect -4392 -1724 -4369 -1641
rect -5178 -1811 -4369 -1724
rect -5178 -1894 -5155 -1811
rect -5072 -1894 -4985 -1811
rect -4902 -1894 -4815 -1811
rect -4732 -1894 -4645 -1811
rect -4562 -1894 -4475 -1811
rect -4392 -1876 -4369 -1811
rect -4392 -1894 -1682 -1876
rect -5178 -1897 -1682 -1894
rect -5178 -1953 -1966 -1897
rect -1910 -1953 -1862 -1897
rect -1806 -1953 -1758 -1897
rect -1702 -1953 -1682 -1897
rect -5178 -1981 -1682 -1953
rect -5178 -2064 -5155 -1981
rect -5072 -2064 -4985 -1981
rect -4902 -2064 -4815 -1981
rect -4732 -2064 -4645 -1981
rect -4562 -2064 -4475 -1981
rect -4392 -2001 -1682 -1981
rect -4392 -2057 -1966 -2001
rect -1910 -2057 -1862 -2001
rect -1806 -2057 -1758 -2001
rect -1702 -2057 -1682 -2001
rect -4392 -2064 -1682 -2057
rect -5178 -2105 -1682 -2064
rect -5178 -2151 -1966 -2105
rect -5178 -2234 -5155 -2151
rect -5072 -2234 -4985 -2151
rect -4902 -2234 -4815 -2151
rect -4732 -2234 -4645 -2151
rect -4562 -2234 -4475 -2151
rect -4392 -2161 -1966 -2151
rect -1910 -2161 -1862 -2105
rect -1806 -2161 -1758 -2105
rect -1702 -2161 -1682 -2105
rect -4392 -2191 -1682 -2161
rect -4392 -2234 -4369 -2191
rect -5178 -2321 -4369 -2234
rect -5178 -2404 -5155 -2321
rect -5072 -2404 -4985 -2321
rect -4902 -2404 -4815 -2321
rect -4732 -2404 -4645 -2321
rect -4562 -2404 -4475 -2321
rect -4392 -2404 -4369 -2321
rect -5178 -2428 -4369 -2404
rect -163 -2262 126 -2244
rect -163 -2318 -152 -2262
rect -96 -2318 -48 -2262
rect 8 -2318 56 -2262
rect 112 -2318 126 -2262
rect -163 -2366 126 -2318
rect -163 -2422 -152 -2366
rect -96 -2422 -48 -2366
rect 8 -2422 56 -2366
rect 112 -2422 126 -2366
rect -163 -2470 126 -2422
rect -163 -2526 -152 -2470
rect -96 -2526 -48 -2470
rect 8 -2526 56 -2470
rect 112 -2493 126 -2470
rect 112 -2526 1118 -2493
rect -163 -2538 1118 -2526
rect -3586 -2604 -372 -2578
rect -106 -2603 1118 -2538
rect -3586 -2660 -3569 -2604
rect -3513 -2660 -3465 -2604
rect -3409 -2660 -3361 -2604
rect -3305 -2660 -372 -2604
rect -3586 -2693 -372 -2660
rect -3586 -2708 1200 -2693
rect -3586 -2764 -3569 -2708
rect -3513 -2764 -3465 -2708
rect -3409 -2764 -3361 -2708
rect -3305 -2764 1200 -2708
rect -3586 -2803 1200 -2764
rect -3586 -2812 -372 -2803
rect -3586 -2868 -3569 -2812
rect -3513 -2868 -3465 -2812
rect -3409 -2868 -3361 -2812
rect -3305 -2868 -372 -2812
rect -3586 -2893 -372 -2868
rect 46 -2929 1176 -2893
rect -68 -2947 1176 -2929
rect -68 -3003 -57 -2947
rect -1 -3003 47 -2947
rect 103 -3003 151 -2947
rect 207 -3003 1176 -2947
rect -1914 -3063 -1625 -3045
rect -1914 -3119 -1903 -3063
rect -1847 -3119 -1799 -3063
rect -1743 -3119 -1695 -3063
rect -1639 -3093 -1625 -3063
rect -68 -3051 221 -3003
rect -1639 -3119 -627 -3093
rect -1914 -3167 -627 -3119
rect -1914 -3223 -1903 -3167
rect -1847 -3223 -1799 -3167
rect -1743 -3223 -1695 -3167
rect -1639 -3203 -627 -3167
rect -1639 -3223 -1625 -3203
rect -1914 -3271 -1625 -3223
rect -1914 -3327 -1903 -3271
rect -1847 -3327 -1799 -3271
rect -1743 -3327 -1695 -3271
rect -1639 -3327 -1625 -3271
rect -1914 -3339 -1625 -3327
rect -737 -3456 -627 -3203
rect -68 -3107 -57 -3051
rect -1 -3107 47 -3051
rect 103 -3107 151 -3051
rect 207 -3107 221 -3051
rect -68 -3155 221 -3107
rect -68 -3211 -57 -3155
rect -1 -3211 47 -3155
rect 103 -3211 151 -3155
rect 207 -3211 221 -3155
rect -68 -3223 221 -3211
rect 390 -3203 1252 -3093
rect 390 -3456 500 -3203
rect -737 -3566 500 -3456
rect 650 -3349 934 -3337
rect 650 -3401 662 -3349
rect 714 -3401 766 -3349
rect 818 -3401 870 -3349
rect 922 -3401 934 -3349
rect 650 -3453 934 -3401
rect 650 -3505 662 -3453
rect 714 -3505 766 -3453
rect 818 -3505 870 -3453
rect 922 -3505 934 -3453
rect 650 -3557 934 -3505
rect 650 -3609 662 -3557
rect 714 -3609 766 -3557
rect 818 -3609 870 -3557
rect 922 -3609 934 -3557
rect 650 -3621 934 -3609
rect -5147 -4702 -4338 -4678
rect -5147 -4785 -5124 -4702
rect -5041 -4785 -4954 -4702
rect -4871 -4785 -4784 -4702
rect -4701 -4785 -4614 -4702
rect -4531 -4785 -4444 -4702
rect -4361 -4785 -4338 -4702
rect -5147 -4872 -4338 -4785
rect -5147 -4955 -5124 -4872
rect -5041 -4955 -4954 -4872
rect -4871 -4955 -4784 -4872
rect -4701 -4955 -4614 -4872
rect -4531 -4955 -4444 -4872
rect -4361 -4935 -4338 -4872
rect -4361 -4955 1066 -4935
rect -5147 -4976 1066 -4955
rect -5147 -5032 731 -4976
rect 787 -5032 835 -4976
rect 891 -5032 939 -4976
rect 995 -5032 1066 -4976
rect -5147 -5042 1066 -5032
rect -5147 -5125 -5124 -5042
rect -5041 -5125 -4954 -5042
rect -4871 -5125 -4784 -5042
rect -4701 -5125 -4614 -5042
rect -4531 -5125 -4444 -5042
rect -4361 -5080 1066 -5042
rect -4361 -5125 731 -5080
rect -5147 -5136 731 -5125
rect 787 -5136 835 -5080
rect 891 -5136 939 -5080
rect 995 -5136 1066 -5080
rect -5147 -5184 1066 -5136
rect -5147 -5212 731 -5184
rect -5147 -5295 -5124 -5212
rect -5041 -5295 -4954 -5212
rect -4871 -5295 -4784 -5212
rect -4701 -5295 -4614 -5212
rect -4531 -5295 -4444 -5212
rect -4361 -5240 731 -5212
rect 787 -5240 835 -5184
rect 891 -5240 939 -5184
rect 995 -5240 1066 -5184
rect -4361 -5263 1066 -5240
rect -4361 -5295 -4338 -5263
rect -5147 -5382 -4338 -5295
rect -5147 -5465 -5124 -5382
rect -5041 -5465 -4954 -5382
rect -4871 -5465 -4784 -5382
rect -4701 -5465 -4614 -5382
rect -4531 -5465 -4444 -5382
rect -4361 -5465 -4338 -5382
rect -5147 -5489 -4338 -5465
rect 16024 -6142 16123 -6126
rect 16024 -6208 16041 -6142
rect 16108 -6208 16123 -6142
rect 16024 -6224 16123 -6208
rect 16441 -6142 16670 10543
rect 16441 -6208 16538 -6142
rect 16605 -6208 16670 -6142
rect -5122 -7571 -4313 -7547
rect -5122 -7654 -5099 -7571
rect -5016 -7654 -4929 -7571
rect -4846 -7654 -4759 -7571
rect -4676 -7654 -4589 -7571
rect -4506 -7654 -4419 -7571
rect -4336 -7654 -4313 -7571
rect -5122 -7741 -4313 -7654
rect -5122 -7824 -5099 -7741
rect -5016 -7824 -4929 -7741
rect -4846 -7824 -4759 -7741
rect -4676 -7824 -4589 -7741
rect -4506 -7824 -4419 -7741
rect -4336 -7824 -4313 -7741
rect -5122 -7832 -4313 -7824
rect -5122 -7858 -2240 -7832
rect -5122 -7876 -2215 -7858
rect -5122 -7911 -2493 -7876
rect -5122 -7994 -5099 -7911
rect -5016 -7994 -4929 -7911
rect -4846 -7994 -4759 -7911
rect -4676 -7994 -4589 -7911
rect -4506 -7994 -4419 -7911
rect -4336 -7932 -2493 -7911
rect -2437 -7932 -2389 -7876
rect -2333 -7932 -2285 -7876
rect -2229 -7932 -2215 -7876
rect -4336 -7980 -2215 -7932
rect -4336 -7994 -2493 -7980
rect -5122 -8036 -2493 -7994
rect -2437 -8036 -2389 -7980
rect -2333 -8036 -2285 -7980
rect -2229 -8036 -2215 -7980
rect -5122 -8081 -2215 -8036
rect -5122 -8164 -5099 -8081
rect -5016 -8164 -4929 -8081
rect -4846 -8164 -4759 -8081
rect -4676 -8164 -4589 -8081
rect -4506 -8164 -4419 -8081
rect -4336 -8084 -2215 -8081
rect -4336 -8140 -2493 -8084
rect -2437 -8140 -2389 -8084
rect -2333 -8140 -2285 -8084
rect -2229 -8140 -2215 -8084
rect -4336 -8152 -2215 -8140
rect -4336 -8160 -2240 -8152
rect -4336 -8164 -4313 -8160
rect -5122 -8251 -4313 -8164
rect -5122 -8334 -5099 -8251
rect -5016 -8334 -4929 -8251
rect -4846 -8334 -4759 -8251
rect -4676 -8334 -4589 -8251
rect -4506 -8334 -4419 -8251
rect -4336 -8334 -4313 -8251
rect -5122 -8358 -4313 -8334
rect -622 -8254 -333 -8236
rect -622 -8310 -611 -8254
rect -555 -8310 -507 -8254
rect -451 -8310 -403 -8254
rect -347 -8310 -333 -8254
rect -622 -8325 -333 -8310
rect 702 -8312 991 -8294
rect 702 -8325 713 -8312
rect -622 -8358 713 -8325
rect -622 -8414 -611 -8358
rect -555 -8414 -507 -8358
rect -451 -8414 -403 -8358
rect -347 -8368 713 -8358
rect 769 -8368 817 -8312
rect 873 -8368 921 -8312
rect 977 -8325 991 -8312
rect 977 -8368 1235 -8325
rect -347 -8414 1235 -8368
rect -622 -8416 1235 -8414
rect -622 -8462 713 -8416
rect -622 -8518 -611 -8462
rect -555 -8518 -507 -8462
rect -451 -8518 -403 -8462
rect -347 -8472 713 -8462
rect 769 -8472 817 -8416
rect 873 -8472 921 -8416
rect 977 -8472 1235 -8416
rect -347 -8518 1235 -8472
rect -622 -8520 1235 -8518
rect -622 -8530 713 -8520
rect -612 -8539 713 -8530
rect 702 -8576 713 -8539
rect 769 -8576 817 -8520
rect 873 -8576 921 -8520
rect 977 -8539 1235 -8520
rect 16028 -8484 16127 -8468
rect 977 -8576 991 -8539
rect 16028 -8550 16045 -8484
rect 16112 -8550 16127 -8484
rect 16028 -8566 16127 -8550
rect 702 -8588 991 -8576
rect -2994 -9073 1088 -9024
rect -2994 -9082 789 -9073
rect -2994 -9138 -2983 -9082
rect -2927 -9138 -2879 -9082
rect -2823 -9138 -2775 -9082
rect -2719 -9129 789 -9082
rect 845 -9129 893 -9073
rect 949 -9129 997 -9073
rect 1053 -9129 1088 -9073
rect -2719 -9138 1088 -9129
rect -2994 -9177 1088 -9138
rect -2994 -9186 789 -9177
rect -2994 -9242 -2983 -9186
rect -2927 -9242 -2879 -9186
rect -2823 -9242 -2775 -9186
rect -2719 -9233 789 -9186
rect 845 -9233 893 -9177
rect 949 -9233 997 -9177
rect 1053 -9233 1088 -9177
rect -2719 -9242 1088 -9233
rect -2994 -9281 1088 -9242
rect -2994 -9290 789 -9281
rect -2994 -9346 -2983 -9290
rect -2927 -9346 -2879 -9290
rect -2823 -9346 -2775 -9290
rect -2719 -9337 789 -9290
rect 845 -9337 893 -9281
rect 949 -9337 997 -9281
rect 1053 -9337 1088 -9281
rect -2719 -9346 1088 -9337
rect -2994 -9354 1088 -9346
rect -2994 -9358 -2705 -9354
rect 16041 -9562 16140 -9546
rect 16041 -9628 16058 -9562
rect 16125 -9628 16140 -9562
rect 16041 -9644 16140 -9628
rect -5099 -9675 -4290 -9651
rect -5099 -9758 -5076 -9675
rect -4993 -9758 -4906 -9675
rect -4823 -9758 -4736 -9675
rect -4653 -9758 -4566 -9675
rect -4483 -9758 -4396 -9675
rect -4313 -9758 -4290 -9675
rect -5099 -9845 -4290 -9758
rect -5099 -9928 -5076 -9845
rect -4993 -9928 -4906 -9845
rect -4823 -9928 -4736 -9845
rect -4653 -9928 -4566 -9845
rect -4483 -9928 -4396 -9845
rect -4313 -9928 -4290 -9845
rect -5099 -9936 -4290 -9928
rect -5099 -10015 -2693 -9936
rect -5099 -10098 -5076 -10015
rect -4993 -10098 -4906 -10015
rect -4823 -10098 -4736 -10015
rect -4653 -10098 -4566 -10015
rect -4483 -10098 -4396 -10015
rect -4313 -10098 -2693 -10015
rect -5099 -10185 -2693 -10098
rect -5099 -10268 -5076 -10185
rect -4993 -10268 -4906 -10185
rect -4823 -10268 -4736 -10185
rect -4653 -10268 -4566 -10185
rect -4483 -10268 -4396 -10185
rect -4313 -10264 -2693 -10185
rect -4313 -10268 -4290 -10264
rect -5099 -10355 -4290 -10268
rect -5099 -10438 -5076 -10355
rect -4993 -10438 -4906 -10355
rect -4823 -10438 -4736 -10355
rect -4653 -10438 -4566 -10355
rect -4483 -10438 -4396 -10355
rect -4313 -10438 -4290 -10355
rect -5099 -10462 -4290 -10438
rect -2988 -10720 -2693 -10264
rect 1143 -10720 1432 -10717
rect -2988 -10735 1432 -10720
rect -2988 -10791 1154 -10735
rect 1210 -10791 1258 -10735
rect 1314 -10791 1362 -10735
rect 1418 -10791 1432 -10735
rect -2988 -10839 1432 -10791
rect -2988 -10895 1154 -10839
rect 1210 -10895 1258 -10839
rect 1314 -10895 1362 -10839
rect 1418 -10895 1432 -10839
rect -2988 -10943 1432 -10895
rect -2988 -10999 1154 -10943
rect 1210 -10999 1258 -10943
rect 1314 -10999 1362 -10943
rect 1418 -10999 1432 -10943
rect -2988 -11011 1432 -10999
rect -2988 -11015 1406 -11011
rect -5076 -11849 -4267 -11825
rect -5076 -11932 -5053 -11849
rect -4970 -11932 -4883 -11849
rect -4800 -11932 -4713 -11849
rect -4630 -11932 -4543 -11849
rect -4460 -11932 -4373 -11849
rect -4290 -11932 -4267 -11849
rect -5076 -12019 -4267 -11932
rect -5076 -12102 -5053 -12019
rect -4970 -12102 -4883 -12019
rect -4800 -12102 -4713 -12019
rect -4630 -12102 -4543 -12019
rect -4460 -12102 -4373 -12019
rect -4290 -12102 -4267 -12019
rect -5076 -12110 -4267 -12102
rect -5076 -12126 -1735 -12110
rect -5076 -12144 -1647 -12126
rect -5076 -12189 -1925 -12144
rect -5076 -12272 -5053 -12189
rect -4970 -12272 -4883 -12189
rect -4800 -12272 -4713 -12189
rect -4630 -12272 -4543 -12189
rect -4460 -12272 -4373 -12189
rect -4290 -12200 -1925 -12189
rect -1869 -12200 -1821 -12144
rect -1765 -12200 -1717 -12144
rect -1661 -12200 -1647 -12144
rect -4290 -12248 -1647 -12200
rect -4290 -12272 -1925 -12248
rect -5076 -12304 -1925 -12272
rect -1869 -12304 -1821 -12248
rect -1765 -12304 -1717 -12248
rect -1661 -12304 -1647 -12248
rect -5076 -12352 -1647 -12304
rect -5076 -12359 -1925 -12352
rect -5076 -12442 -5053 -12359
rect -4970 -12442 -4883 -12359
rect -4800 -12442 -4713 -12359
rect -4630 -12442 -4543 -12359
rect -4460 -12442 -4373 -12359
rect -4290 -12408 -1925 -12359
rect -1869 -12408 -1821 -12352
rect -1765 -12408 -1717 -12352
rect -1661 -12408 -1647 -12352
rect -4290 -12420 -1647 -12408
rect -4290 -12438 -1735 -12420
rect -4290 -12442 -4267 -12438
rect -5076 -12529 -4267 -12442
rect -5076 -12612 -5053 -12529
rect -4970 -12612 -4883 -12529
rect -4800 -12612 -4713 -12529
rect -4630 -12612 -4543 -12529
rect -4460 -12612 -4373 -12529
rect -4290 -12612 -4267 -12529
rect -5076 -12636 -4267 -12612
rect -5122 -13653 -4313 -13629
rect -5122 -13736 -5099 -13653
rect -5016 -13736 -4929 -13653
rect -4846 -13736 -4759 -13653
rect -4676 -13736 -4589 -13653
rect -4506 -13736 -4419 -13653
rect -4336 -13736 -4313 -13653
rect -5122 -13823 -4313 -13736
rect -5122 -13906 -5099 -13823
rect -5016 -13906 -4929 -13823
rect -4846 -13906 -4759 -13823
rect -4676 -13906 -4589 -13823
rect -4506 -13906 -4419 -13823
rect -4336 -13906 -4313 -13823
rect -5122 -13920 -4313 -13906
rect -5122 -13931 -1340 -13920
rect -5122 -13949 -1193 -13931
rect -5122 -13993 -1471 -13949
rect -5122 -14076 -5099 -13993
rect -5016 -14076 -4929 -13993
rect -4846 -14076 -4759 -13993
rect -4676 -14076 -4589 -13993
rect -4506 -14076 -4419 -13993
rect -4336 -14005 -1471 -13993
rect -1415 -14005 -1367 -13949
rect -1311 -14005 -1263 -13949
rect -1207 -14005 -1193 -13949
rect -4336 -14053 -1193 -14005
rect -4336 -14076 -1471 -14053
rect -5122 -14109 -1471 -14076
rect -1415 -14109 -1367 -14053
rect -1311 -14109 -1263 -14053
rect -1207 -14109 -1193 -14053
rect -5122 -14157 -1193 -14109
rect -5122 -14163 -1471 -14157
rect -5122 -14246 -5099 -14163
rect -5016 -14246 -4929 -14163
rect -4846 -14246 -4759 -14163
rect -4676 -14246 -4589 -14163
rect -4506 -14246 -4419 -14163
rect -4336 -14213 -1471 -14163
rect -1415 -14213 -1367 -14157
rect -1311 -14213 -1263 -14157
rect -1207 -14213 -1193 -14157
rect -4336 -14225 -1193 -14213
rect -4336 -14238 -1340 -14225
rect -4336 -14246 -4313 -14238
rect -5122 -14333 -4313 -14246
rect -5122 -14416 -5099 -14333
rect -5016 -14416 -4929 -14333
rect -4846 -14416 -4759 -14333
rect -4676 -14416 -4589 -14333
rect -4506 -14416 -4419 -14333
rect -4336 -14416 -4313 -14333
rect -5122 -14440 -4313 -14416
rect -5076 -15425 -4267 -15401
rect -5076 -15508 -5053 -15425
rect -4970 -15508 -4883 -15425
rect -4800 -15508 -4713 -15425
rect -4630 -15508 -4543 -15425
rect -4460 -15508 -4373 -15425
rect -4290 -15508 -4267 -15425
rect -5076 -15595 -4267 -15508
rect -5076 -15678 -5053 -15595
rect -4970 -15678 -4883 -15595
rect -4800 -15678 -4713 -15595
rect -4630 -15678 -4543 -15595
rect -4460 -15678 -4373 -15595
rect -4290 -15678 -4267 -15595
rect -5076 -15686 -4267 -15678
rect -5076 -15718 241 -15686
rect -5076 -15765 -66 -15718
rect -5076 -15848 -5053 -15765
rect -4970 -15848 -4883 -15765
rect -4800 -15848 -4713 -15765
rect -4630 -15848 -4543 -15765
rect -4460 -15848 -4373 -15765
rect -4290 -15774 -66 -15765
rect -10 -15774 38 -15718
rect 94 -15774 142 -15718
rect 198 -15774 241 -15718
rect -4290 -15822 241 -15774
rect -4290 -15848 -66 -15822
rect -5076 -15878 -66 -15848
rect -10 -15878 38 -15822
rect 94 -15878 142 -15822
rect 198 -15878 241 -15822
rect -5076 -15926 241 -15878
rect -5076 -15935 -66 -15926
rect -5076 -16018 -5053 -15935
rect -4970 -16018 -4883 -15935
rect -4800 -16018 -4713 -15935
rect -4630 -16018 -4543 -15935
rect -4460 -16018 -4373 -15935
rect -4290 -15982 -66 -15935
rect -10 -15982 38 -15926
rect 94 -15982 142 -15926
rect 198 -15982 241 -15926
rect -4290 -16014 241 -15982
rect -4290 -16018 -4267 -16014
rect -5076 -16105 -4267 -16018
rect -5076 -16188 -5053 -16105
rect -4970 -16188 -4883 -16105
rect -4800 -16188 -4713 -16105
rect -4630 -16188 -4543 -16105
rect -4460 -16188 -4373 -16105
rect -4290 -16188 -4267 -16105
rect -5076 -16212 -4267 -16188
rect 16441 -16980 16670 -6208
rect 16963 8279 17192 11691
rect 16963 8213 17047 8279
rect 17114 8213 17192 8279
rect 16963 -8484 17192 8213
rect 16963 -8550 17013 -8484
rect 17080 -8550 17192 -8484
rect 16963 -15496 17192 -8550
rect 17492 7207 17721 11693
rect 17492 7141 17599 7207
rect 17666 7141 17721 7207
rect 17492 -9562 17721 7141
rect 18170 -5742 18536 16499
rect 21980 16458 22004 16541
rect 22087 16458 22174 16541
rect 22257 16458 22344 16541
rect 22427 16458 22514 16541
rect 22597 16458 22684 16541
rect 22767 16458 22791 16541
rect 21980 16435 22791 16458
rect 22199 14862 22564 16435
rect 52321 16332 53132 16355
rect 49167 16304 49978 16327
rect 49167 16221 49191 16304
rect 49274 16221 49361 16304
rect 49444 16221 49531 16304
rect 49614 16221 49701 16304
rect 49784 16221 49871 16304
rect 49954 16221 49978 16304
rect 49167 16134 49978 16221
rect 49167 16051 49191 16134
rect 49274 16051 49361 16134
rect 49444 16051 49531 16134
rect 49614 16051 49701 16134
rect 49784 16051 49871 16134
rect 49954 16051 49978 16134
rect 49167 15964 49978 16051
rect 49167 15881 49191 15964
rect 49274 15881 49361 15964
rect 49444 15881 49531 15964
rect 49614 15881 49701 15964
rect 49784 15881 49871 15964
rect 49954 15881 49978 15964
rect 49167 15794 49978 15881
rect 49167 15711 49191 15794
rect 49274 15711 49361 15794
rect 49444 15711 49531 15794
rect 49614 15711 49701 15794
rect 49784 15711 49871 15794
rect 49954 15711 49978 15794
rect 49167 15624 49978 15711
rect 49167 15541 49191 15624
rect 49274 15541 49361 15624
rect 49444 15541 49531 15624
rect 49614 15541 49701 15624
rect 49784 15541 49871 15624
rect 49954 15541 49978 15624
rect 52321 16249 52345 16332
rect 52428 16249 52515 16332
rect 52598 16249 52685 16332
rect 52768 16249 52855 16332
rect 52938 16249 53025 16332
rect 53108 16249 53132 16332
rect 52321 16162 53132 16249
rect 52321 16079 52345 16162
rect 52428 16079 52515 16162
rect 52598 16079 52685 16162
rect 52768 16079 52855 16162
rect 52938 16079 53025 16162
rect 53108 16079 53132 16162
rect 52321 15992 53132 16079
rect 52321 15909 52345 15992
rect 52428 15909 52515 15992
rect 52598 15909 52685 15992
rect 52768 15909 52855 15992
rect 52938 15909 53025 15992
rect 53108 15909 53132 15992
rect 52321 15822 53132 15909
rect 52321 15739 52345 15822
rect 52428 15739 52515 15822
rect 52598 15739 52685 15822
rect 52768 15739 52855 15822
rect 52938 15739 53025 15822
rect 53108 15739 53132 15822
rect 52321 15652 53132 15739
rect 52321 15569 52345 15652
rect 52428 15569 52515 15652
rect 52598 15569 52685 15652
rect 52768 15569 52855 15652
rect 52938 15569 53025 15652
rect 53108 15569 53132 15652
rect 52321 15546 53132 15569
rect 49167 15518 49978 15541
rect 18872 14497 22564 14862
rect 18872 9352 19237 14497
rect 85851 13414 86135 16582
rect 89240 16573 90051 16596
rect 154944 17163 155755 17186
rect 154944 17080 154968 17163
rect 155051 17080 155138 17163
rect 155221 17080 155308 17163
rect 155391 17080 155478 17163
rect 155561 17080 155648 17163
rect 155731 17080 155755 17163
rect 154944 16993 155755 17080
rect 154944 16910 154968 16993
rect 155051 16910 155138 16993
rect 155221 16910 155308 16993
rect 155391 16910 155478 16993
rect 155561 16910 155648 16993
rect 155731 16910 155755 16993
rect 154944 16823 155755 16910
rect 154944 16740 154968 16823
rect 155051 16740 155138 16823
rect 155221 16740 155308 16823
rect 155391 16740 155478 16823
rect 155561 16740 155648 16823
rect 155731 16740 155755 16823
rect 154944 16653 155755 16740
rect 89467 14497 89745 16573
rect 154944 16570 154968 16653
rect 155051 16570 155138 16653
rect 155221 16570 155308 16653
rect 155391 16570 155478 16653
rect 155561 16570 155648 16653
rect 155731 16570 155755 16653
rect 154944 16483 155755 16570
rect 154944 16400 154968 16483
rect 155051 16400 155138 16483
rect 155221 16400 155308 16483
rect 155391 16400 155478 16483
rect 155561 16400 155648 16483
rect 155731 16400 155755 16483
rect 154944 16377 155755 16400
rect 157319 17163 158130 17186
rect 157319 17080 157343 17163
rect 157426 17080 157513 17163
rect 157596 17080 157683 17163
rect 157766 17080 157853 17163
rect 157936 17080 158023 17163
rect 158106 17080 158130 17163
rect 157319 16993 158130 17080
rect 157319 16910 157343 16993
rect 157426 16910 157513 16993
rect 157596 16910 157683 16993
rect 157766 16910 157853 16993
rect 157936 16910 158023 16993
rect 158106 16910 158130 16993
rect 157319 16823 158130 16910
rect 157319 16740 157343 16823
rect 157426 16740 157513 16823
rect 157596 16740 157683 16823
rect 157766 16740 157853 16823
rect 157936 16740 158023 16823
rect 158106 16740 158130 16823
rect 157319 16653 158130 16740
rect 157319 16570 157343 16653
rect 157426 16570 157513 16653
rect 157596 16570 157683 16653
rect 157766 16570 157853 16653
rect 157936 16570 158023 16653
rect 158106 16570 158130 16653
rect 157319 16483 158130 16570
rect 157319 16400 157343 16483
rect 157426 16400 157513 16483
rect 157596 16400 157683 16483
rect 157766 16400 157853 16483
rect 157936 16400 158023 16483
rect 158106 16400 158130 16483
rect 157319 16377 158130 16400
rect 86765 14219 89745 14497
rect 133279 14440 134136 14513
rect 133279 14439 134010 14440
rect 133279 14437 133676 14439
rect 133279 14349 133349 14437
rect 133436 14349 133529 14437
rect 133616 14351 133676 14437
rect 133763 14351 133856 14439
rect 133943 14352 134010 14439
rect 134097 14352 134136 14440
rect 133943 14351 134136 14352
rect 133616 14349 134136 14351
rect 133279 14260 134136 14349
rect 133279 14259 134010 14260
rect 133279 14257 133676 14259
rect 86765 13094 87043 14219
rect 133279 14169 133349 14257
rect 133436 14169 133529 14257
rect 133616 14171 133676 14257
rect 133763 14171 133856 14259
rect 133943 14172 134010 14259
rect 134097 14172 134136 14260
rect 133943 14171 134136 14172
rect 133616 14169 134136 14171
rect 133279 14047 134136 14169
rect 133279 14046 133992 14047
rect 133279 14044 133658 14046
rect 133279 13956 133331 14044
rect 133418 13956 133511 14044
rect 133598 13958 133658 14044
rect 133745 13958 133838 14046
rect 133925 13959 133992 14046
rect 134079 13959 134136 14047
rect 133925 13958 134136 13959
rect 133598 13956 134136 13958
rect 133279 13867 134136 13956
rect 133279 13866 133992 13867
rect 133279 13864 133658 13866
rect 133279 13776 133331 13864
rect 133418 13776 133511 13864
rect 133598 13778 133658 13864
rect 133745 13778 133838 13866
rect 133925 13779 133992 13866
rect 134079 13779 134136 13867
rect 133925 13778 134136 13779
rect 133598 13776 134136 13778
rect 133279 13698 134136 13776
rect 135785 14424 136642 14497
rect 135785 14423 136516 14424
rect 135785 14421 136182 14423
rect 135785 14333 135855 14421
rect 135942 14333 136035 14421
rect 136122 14335 136182 14421
rect 136269 14335 136362 14423
rect 136449 14336 136516 14423
rect 136603 14336 136642 14424
rect 136449 14335 136642 14336
rect 136122 14333 136642 14335
rect 135785 14244 136642 14333
rect 135785 14243 136516 14244
rect 135785 14241 136182 14243
rect 135785 14153 135855 14241
rect 135942 14153 136035 14241
rect 136122 14155 136182 14241
rect 136269 14155 136362 14243
rect 136449 14156 136516 14243
rect 136603 14156 136642 14244
rect 136449 14155 136642 14156
rect 136122 14153 136642 14155
rect 135785 14031 136642 14153
rect 135785 14030 136498 14031
rect 135785 14028 136164 14030
rect 135785 13940 135837 14028
rect 135924 13940 136017 14028
rect 136104 13942 136164 14028
rect 136251 13942 136344 14030
rect 136431 13943 136498 14030
rect 136585 13943 136642 14031
rect 136431 13942 136642 13943
rect 136104 13940 136642 13942
rect 135785 13851 136642 13940
rect 135785 13850 136498 13851
rect 135785 13848 136164 13850
rect 135785 13760 135837 13848
rect 135924 13760 136017 13848
rect 136104 13762 136164 13848
rect 136251 13762 136344 13850
rect 136431 13763 136498 13850
rect 136585 13763 136642 13851
rect 136431 13762 136642 13763
rect 136104 13760 136642 13762
rect 135785 13682 136642 13760
rect 138501 14443 139358 14516
rect 138501 14442 139232 14443
rect 138501 14440 138898 14442
rect 138501 14352 138571 14440
rect 138658 14352 138751 14440
rect 138838 14354 138898 14440
rect 138985 14354 139078 14442
rect 139165 14355 139232 14442
rect 139319 14355 139358 14443
rect 139165 14354 139358 14355
rect 138838 14352 139358 14354
rect 138501 14263 139358 14352
rect 138501 14262 139232 14263
rect 138501 14260 138898 14262
rect 138501 14172 138571 14260
rect 138658 14172 138751 14260
rect 138838 14174 138898 14260
rect 138985 14174 139078 14262
rect 139165 14175 139232 14262
rect 139319 14175 139358 14263
rect 139165 14174 139358 14175
rect 138838 14172 139358 14174
rect 138501 14050 139358 14172
rect 155138 14084 155422 16377
rect 157543 14928 157821 16377
rect 156052 14650 157821 14928
rect 138501 14049 139214 14050
rect 138501 14047 138880 14049
rect 138501 13959 138553 14047
rect 138640 13959 138733 14047
rect 138820 13961 138880 14047
rect 138967 13961 139060 14049
rect 139147 13962 139214 14049
rect 139301 13962 139358 14050
rect 139147 13961 139358 13962
rect 138820 13959 139358 13961
rect 138501 13870 139358 13959
rect 138501 13869 139214 13870
rect 138501 13867 138880 13869
rect 138501 13779 138553 13867
rect 138640 13779 138733 13867
rect 138820 13781 138880 13867
rect 138967 13781 139060 13869
rect 139147 13782 139214 13869
rect 139301 13782 139358 13870
rect 156052 13845 156330 14650
rect 139147 13781 139358 13782
rect 138820 13779 139358 13781
rect 138501 13701 139358 13779
rect 23334 12875 23628 12889
rect 23334 12787 23348 12875
rect 23435 12787 23528 12875
rect 23615 12787 23628 12875
rect 23334 12695 23628 12787
rect 23334 12607 23348 12695
rect 23435 12607 23528 12695
rect 23615 12607 23628 12695
rect 23334 12593 23628 12607
rect 18781 9293 19303 9352
rect 18781 9210 18836 9293
rect 18919 9210 19006 9293
rect 19089 9210 19176 9293
rect 19259 9210 19303 9293
rect 18781 9123 19303 9210
rect 18781 9040 18836 9123
rect 18919 9040 19006 9123
rect 19089 9040 19176 9123
rect 19259 9040 19303 9123
rect 18781 8953 19303 9040
rect 18781 8870 18836 8953
rect 18919 8870 19006 8953
rect 19089 8870 19176 8953
rect 19259 8870 19303 8953
rect 18781 8714 19303 8870
rect 18781 8631 18838 8714
rect 18921 8631 19008 8714
rect 19091 8631 19178 8714
rect 19261 8631 19303 8714
rect 18781 8544 19303 8631
rect 18781 8461 18838 8544
rect 18921 8461 19008 8544
rect 19091 8461 19178 8544
rect 19261 8461 19303 8544
rect 18781 8374 19303 8461
rect 18781 8291 18838 8374
rect 18921 8291 19008 8374
rect 19091 8291 19178 8374
rect 19261 8291 19303 8374
rect 18781 8226 19303 8291
rect 150298 6671 151141 6731
rect 150298 6670 151003 6671
rect 150298 6668 150669 6670
rect 150298 6580 150342 6668
rect 150429 6580 150522 6668
rect 150609 6582 150669 6668
rect 150756 6582 150849 6670
rect 150936 6583 151003 6670
rect 151090 6583 151141 6671
rect 150936 6582 151141 6583
rect 150609 6580 151141 6582
rect 150298 6491 151141 6580
rect 150298 6490 151003 6491
rect 150298 6488 150669 6490
rect 150298 6400 150342 6488
rect 150429 6400 150522 6488
rect 150609 6402 150669 6488
rect 150756 6402 150849 6490
rect 150936 6403 151003 6490
rect 151090 6403 151141 6491
rect 150936 6402 151141 6403
rect 150609 6400 151141 6402
rect 150298 6356 151141 6400
rect 80879 6043 81977 6073
rect 75608 5997 76748 6038
rect 75608 5996 76309 5997
rect 75608 5994 75975 5996
rect 75608 5906 75648 5994
rect 75735 5906 75828 5994
rect 75915 5908 75975 5994
rect 76062 5908 76155 5996
rect 76242 5909 76309 5996
rect 76396 5996 76748 5997
rect 76396 5909 76449 5996
rect 76242 5908 76449 5909
rect 76536 5994 76748 5996
rect 76536 5908 76590 5994
rect 75915 5906 76590 5908
rect 76677 5906 76748 5994
rect 75608 5817 76748 5906
rect 75608 5816 76309 5817
rect 75608 5814 75975 5816
rect 75608 5726 75648 5814
rect 75735 5726 75828 5814
rect 75915 5728 75975 5814
rect 76062 5728 76155 5816
rect 76242 5729 76309 5816
rect 76396 5816 76748 5817
rect 76396 5729 76449 5816
rect 76242 5728 76449 5729
rect 76536 5814 76748 5816
rect 76536 5728 76590 5814
rect 75915 5726 76590 5728
rect 76677 5726 76748 5814
rect 75608 5683 76748 5726
rect 80879 6033 81982 6043
rect 80879 6032 81734 6033
rect 80879 6031 81580 6032
rect 80879 6029 81246 6031
rect 80879 5941 80919 6029
rect 81006 5941 81099 6029
rect 81186 5943 81246 6029
rect 81333 5943 81426 6031
rect 81513 5944 81580 6031
rect 81667 5945 81734 6032
rect 81821 6031 81982 6033
rect 81821 5945 81882 6031
rect 81667 5944 81882 5945
rect 81513 5943 81882 5944
rect 81969 5943 81982 6031
rect 81186 5941 81982 5943
rect 80879 5853 81982 5941
rect 80879 5852 81734 5853
rect 80879 5851 81580 5852
rect 80879 5849 81246 5851
rect 80879 5761 80919 5849
rect 81006 5761 81099 5849
rect 81186 5763 81246 5849
rect 81333 5763 81426 5851
rect 81513 5764 81580 5851
rect 81667 5765 81734 5852
rect 81821 5851 81982 5853
rect 81821 5765 81882 5851
rect 81667 5764 81882 5765
rect 81513 5763 81882 5764
rect 81969 5763 81982 5851
rect 81186 5761 81982 5763
rect 80879 5746 81982 5761
rect 80879 5718 81977 5746
rect 126076 4902 126522 4934
rect 126076 4814 126226 4902
rect 126313 4814 126406 4902
rect 126493 4814 126522 4902
rect 126076 4722 126522 4814
rect 126076 4634 126226 4722
rect 126313 4634 126406 4722
rect 126493 4634 126522 4722
rect 126076 4333 126522 4634
rect 56786 4217 57185 4277
rect 56786 4129 56847 4217
rect 56934 4129 57027 4217
rect 57114 4129 57185 4217
rect 56786 4037 57185 4129
rect 56786 3949 56847 4037
rect 56934 3949 57027 4037
rect 57114 3949 57185 4037
rect 56786 3600 57185 3949
rect 115054 3958 115376 3977
rect 114442 3912 114764 3930
rect 113812 3862 114134 3879
rect 113812 3774 113837 3862
rect 113924 3774 114017 3862
rect 114104 3774 114134 3862
rect 113812 3682 114134 3774
rect 113812 3594 113837 3682
rect 113924 3594 114017 3682
rect 114104 3594 114134 3682
rect 113812 3521 114134 3594
rect 113812 3433 113839 3521
rect 113926 3433 114019 3521
rect 114106 3433 114134 3521
rect 113812 3341 114134 3433
rect 113812 3253 113839 3341
rect 113926 3253 114019 3341
rect 114106 3253 114134 3341
rect 114442 3824 114475 3912
rect 114562 3824 114655 3912
rect 114742 3824 114764 3912
rect 114442 3732 114764 3824
rect 114442 3644 114475 3732
rect 114562 3644 114655 3732
rect 114742 3644 114764 3732
rect 114442 3569 114764 3644
rect 114442 3481 114473 3569
rect 114560 3481 114653 3569
rect 114740 3481 114764 3569
rect 114442 3389 114764 3481
rect 114442 3301 114473 3389
rect 114560 3301 114653 3389
rect 114740 3301 114764 3389
rect 115054 3870 115082 3958
rect 115169 3870 115262 3958
rect 115349 3870 115376 3958
rect 115054 3778 115376 3870
rect 115054 3690 115082 3778
rect 115169 3690 115262 3778
rect 115349 3690 115376 3778
rect 115054 3618 115376 3690
rect 115054 3530 115082 3618
rect 115169 3530 115262 3618
rect 115349 3530 115376 3618
rect 115054 3438 115376 3530
rect 115054 3350 115082 3438
rect 115169 3350 115262 3438
rect 115349 3350 115376 3438
rect 115054 3329 115376 3350
rect 115708 3940 116010 3955
rect 115708 3852 115729 3940
rect 115816 3852 115909 3940
rect 115996 3852 116010 3940
rect 115708 3760 116010 3852
rect 115708 3672 115729 3760
rect 115816 3672 115909 3760
rect 115996 3672 116010 3760
rect 115708 3623 116010 3672
rect 115708 3609 116012 3623
rect 115708 3521 115732 3609
rect 115819 3521 115912 3609
rect 115999 3521 116012 3609
rect 115708 3429 116012 3521
rect 115708 3341 115732 3429
rect 115819 3341 115912 3429
rect 115999 3341 116012 3429
rect 114442 3282 114764 3301
rect 113812 3231 114134 3253
rect 113913 2675 114096 3231
rect 114555 3143 114738 3282
rect 114463 2960 114738 3143
rect 115142 3025 115325 3329
rect 115708 3327 116012 3341
rect 115708 3317 116010 3327
rect 115761 3050 115944 3317
rect 114463 2675 114646 2960
rect 114985 2842 115325 3025
rect 115536 2867 115944 3050
rect 113897 2660 114113 2675
rect 113897 2595 113912 2660
rect 113974 2595 114037 2660
rect 114099 2595 114113 2660
rect 113897 2535 114113 2595
rect 113897 2470 113912 2535
rect 113974 2470 114037 2535
rect 114099 2470 114113 2535
rect 113897 2456 114113 2470
rect 114443 2660 114659 2675
rect 114985 2666 115168 2842
rect 115536 2668 115719 2867
rect 114443 2595 114458 2660
rect 114520 2595 114583 2660
rect 114645 2595 114659 2660
rect 114443 2535 114659 2595
rect 114443 2470 114458 2535
rect 114520 2470 114583 2535
rect 114645 2470 114659 2535
rect 114443 2456 114659 2470
rect 114971 2651 115187 2666
rect 114971 2586 114986 2651
rect 115048 2586 115111 2651
rect 115173 2586 115187 2651
rect 114971 2526 115187 2586
rect 114971 2461 114986 2526
rect 115048 2461 115111 2526
rect 115173 2461 115187 2526
rect 114971 2447 115187 2461
rect 115520 2653 115736 2668
rect 115520 2588 115535 2653
rect 115597 2588 115660 2653
rect 115722 2588 115736 2653
rect 115520 2528 115736 2588
rect 115520 2463 115535 2528
rect 115597 2463 115660 2528
rect 115722 2463 115736 2528
rect 115520 2449 115736 2463
rect 114987 1810 115224 1825
rect 114987 1747 115006 1810
rect 115069 1808 115224 1810
rect 115069 1747 115144 1808
rect 114987 1745 115144 1747
rect 115207 1745 115224 1808
rect 114987 1733 115224 1745
rect 114165 1646 114402 1661
rect 114165 1583 114184 1646
rect 114247 1644 114402 1646
rect 114247 1583 114322 1644
rect 114165 1581 114322 1583
rect 114385 1581 114402 1644
rect 114165 1569 114402 1581
rect 47817 1118 50889 1322
rect 47817 862 48021 1118
rect 47817 810 47846 862
rect 47898 810 47950 862
rect 48002 810 48021 862
rect 28005 680 28862 753
rect 28005 679 28736 680
rect 28005 677 28402 679
rect 28005 589 28075 677
rect 28162 589 28255 677
rect 28342 591 28402 677
rect 28489 591 28582 679
rect 28669 592 28736 679
rect 28823 592 28862 680
rect 28669 591 28862 592
rect 28342 589 28862 591
rect 28005 500 28862 589
rect 28005 499 28736 500
rect 28005 497 28402 499
rect 28005 409 28075 497
rect 28162 409 28255 497
rect 28342 411 28402 497
rect 28489 411 28582 499
rect 28669 412 28736 499
rect 28823 412 28862 500
rect 28669 411 28862 412
rect 28342 409 28862 411
rect 28005 287 28862 409
rect 28005 286 28718 287
rect 28005 284 28384 286
rect 28005 196 28057 284
rect 28144 196 28237 284
rect 28324 198 28384 284
rect 28471 198 28564 286
rect 28651 199 28718 286
rect 28805 199 28862 287
rect 28651 198 28862 199
rect 28324 196 28862 198
rect 28005 107 28862 196
rect 28005 106 28718 107
rect 28005 104 28384 106
rect 28005 16 28057 104
rect 28144 16 28237 104
rect 28324 18 28384 104
rect 28471 18 28564 106
rect 28651 19 28718 106
rect 28805 19 28862 107
rect 28651 18 28862 19
rect 28324 16 28862 18
rect 28005 -63 28862 16
rect 29817 727 30674 793
rect 29817 726 30542 727
rect 29817 724 30208 726
rect 29817 636 29881 724
rect 29968 636 30061 724
rect 30148 638 30208 724
rect 30295 638 30388 726
rect 30475 639 30542 726
rect 30629 639 30674 727
rect 30475 638 30674 639
rect 30148 636 30674 638
rect 29817 547 30674 636
rect 29817 546 30542 547
rect 29817 544 30208 546
rect 29817 456 29881 544
rect 29968 456 30061 544
rect 30148 458 30208 544
rect 30295 458 30388 546
rect 30475 459 30542 546
rect 30629 459 30674 547
rect 30475 458 30674 459
rect 30148 456 30674 458
rect 29817 339 30674 456
rect 29817 338 30548 339
rect 29817 336 30214 338
rect 29817 248 29887 336
rect 29974 248 30067 336
rect 30154 250 30214 336
rect 30301 250 30394 338
rect 30481 251 30548 338
rect 30635 251 30674 339
rect 30481 250 30674 251
rect 30154 248 30674 250
rect 29817 159 30674 248
rect 29817 158 30548 159
rect 29817 156 30214 158
rect 29817 68 29887 156
rect 29974 68 30067 156
rect 30154 70 30214 156
rect 30301 70 30394 158
rect 30481 71 30548 158
rect 30635 71 30674 159
rect 30481 70 30674 71
rect 30154 68 30674 70
rect 29817 -23 30674 68
rect 31572 727 32429 770
rect 31572 726 32279 727
rect 31572 724 31945 726
rect 31572 636 31618 724
rect 31705 636 31798 724
rect 31885 638 31945 724
rect 32032 638 32125 726
rect 32212 639 32279 726
rect 32366 639 32429 727
rect 47817 758 48021 810
rect 47817 706 47846 758
rect 47898 706 47950 758
rect 48002 706 48021 758
rect 47817 674 48021 706
rect 48388 764 48752 791
rect 48388 699 48410 764
rect 48475 699 48535 764
rect 48600 699 48660 764
rect 48725 699 48752 764
rect 48388 675 48752 699
rect 32212 638 32429 639
rect 31885 636 32429 638
rect 31572 547 32429 636
rect 31572 546 32279 547
rect 31572 544 31945 546
rect 31572 456 31618 544
rect 31705 456 31798 544
rect 31885 458 31945 544
rect 32032 458 32125 546
rect 32212 459 32279 546
rect 32366 459 32429 547
rect 32212 458 32429 459
rect 31885 456 32429 458
rect 31572 339 32429 456
rect 31572 338 32291 339
rect 31572 336 31957 338
rect 31572 248 31630 336
rect 31717 248 31810 336
rect 31897 250 31957 336
rect 32044 250 32137 338
rect 32224 251 32291 338
rect 32378 251 32429 339
rect 32224 250 32429 251
rect 31897 248 32429 250
rect 31572 159 32429 248
rect 31572 158 32291 159
rect 31572 156 31957 158
rect 31572 68 31630 156
rect 31717 68 31810 156
rect 31897 70 31957 156
rect 32044 70 32137 158
rect 32224 71 32291 158
rect 32378 71 32429 159
rect 32224 70 32429 71
rect 31897 68 32429 70
rect 31572 -46 32429 68
rect 48101 -624 48851 -611
rect 48101 -676 48120 -624
rect 48172 -676 48224 -624
rect 48276 -631 48851 -624
rect 48276 -676 48678 -631
rect 48101 -683 48678 -676
rect 48730 -683 48782 -631
rect 48834 -683 48851 -631
rect 48101 -728 48851 -683
rect 48101 -780 48120 -728
rect 48172 -780 48224 -728
rect 48276 -735 48851 -728
rect 48276 -780 48678 -735
rect 48101 -787 48678 -780
rect 48730 -787 48782 -735
rect 48834 -787 48851 -735
rect 48101 -799 48851 -787
rect 64649 -1261 64809 1569
rect 64609 -1280 64825 -1261
rect 64609 -1336 64643 -1280
rect 64699 -1336 64747 -1280
rect 64803 -1336 64825 -1280
rect 64609 -1384 64825 -1336
rect 64609 -1440 64643 -1384
rect 64699 -1440 64747 -1384
rect 64803 -1440 64825 -1384
rect 64609 -1514 64825 -1440
rect 64609 -1570 64645 -1514
rect 64701 -1570 64749 -1514
rect 64805 -1570 64825 -1514
rect 64609 -1618 64825 -1570
rect 64609 -1674 64645 -1618
rect 64701 -1674 64749 -1618
rect 64805 -1674 64825 -1618
rect 64609 -1703 64825 -1674
rect 23075 -2069 23369 -2055
rect 23075 -2157 23089 -2069
rect 23176 -2157 23269 -2069
rect 23356 -2157 23369 -2069
rect 23075 -2249 23369 -2157
rect 23075 -2337 23089 -2249
rect 23176 -2337 23269 -2249
rect 23356 -2337 23369 -2249
rect 23075 -2351 23369 -2337
rect 85851 -3243 86135 -432
rect 86759 -2092 87043 -361
rect 86665 -2131 87681 -2092
rect 86665 -2219 86691 -2131
rect 86778 -2219 86871 -2131
rect 86958 -2219 87037 -2131
rect 87124 -2219 87217 -2131
rect 87304 -2134 87681 -2131
rect 87304 -2219 87390 -2134
rect 86665 -2222 87390 -2219
rect 87477 -2222 87570 -2134
rect 87657 -2222 87681 -2134
rect 86665 -2311 87681 -2222
rect 86665 -2399 86691 -2311
rect 86778 -2399 86871 -2311
rect 86958 -2399 87037 -2311
rect 87124 -2399 87217 -2311
rect 87304 -2314 87681 -2311
rect 87304 -2399 87390 -2314
rect 86665 -2402 87390 -2399
rect 87477 -2402 87570 -2314
rect 87657 -2402 87681 -2314
rect 86665 -2431 87681 -2402
rect 86759 -2497 87043 -2431
rect 85723 -3282 86739 -3243
rect 85723 -3370 85749 -3282
rect 85836 -3370 85929 -3282
rect 86016 -3370 86095 -3282
rect 86182 -3370 86275 -3282
rect 86362 -3285 86739 -3282
rect 86362 -3370 86448 -3285
rect 85723 -3373 86448 -3370
rect 86535 -3373 86628 -3285
rect 86715 -3373 86739 -3285
rect 85723 -3462 86739 -3373
rect 85723 -3550 85749 -3462
rect 85836 -3550 85929 -3462
rect 86016 -3550 86095 -3462
rect 86182 -3550 86275 -3462
rect 86362 -3465 86739 -3462
rect 86362 -3550 86448 -3465
rect 85723 -3553 86448 -3550
rect 86535 -3553 86628 -3465
rect 86715 -3553 86739 -3465
rect 85723 -3582 86739 -3553
rect 18093 -5810 18615 -5742
rect 18093 -5893 18142 -5810
rect 18225 -5893 18312 -5810
rect 18395 -5893 18482 -5810
rect 18565 -5893 18615 -5810
rect 18093 -5980 18615 -5893
rect 18093 -6063 18142 -5980
rect 18225 -6063 18312 -5980
rect 18395 -6063 18482 -5980
rect 18565 -6063 18615 -5980
rect 18093 -6150 18615 -6063
rect 18093 -6233 18142 -6150
rect 18225 -6233 18312 -6150
rect 18395 -6233 18482 -6150
rect 18565 -6233 18615 -6150
rect 18093 -6392 18615 -6233
rect 18093 -6475 18151 -6392
rect 18234 -6475 18321 -6392
rect 18404 -6475 18491 -6392
rect 18574 -6475 18615 -6392
rect 18093 -6562 18615 -6475
rect 18093 -6645 18151 -6562
rect 18234 -6645 18321 -6562
rect 18404 -6645 18491 -6562
rect 18574 -6645 18615 -6562
rect 18093 -6732 18615 -6645
rect 18093 -6815 18151 -6732
rect 18234 -6815 18321 -6732
rect 18404 -6815 18491 -6732
rect 18574 -6815 18615 -6732
rect 18093 -6868 18615 -6815
rect 17492 -9628 17557 -9562
rect 17624 -9628 17721 -9562
rect 17492 -14720 17721 -9628
rect 114186 -13748 114380 1569
rect 113311 -13942 114380 -13748
rect 115006 -13734 115200 1733
rect 127066 270 128070 310
rect 127066 268 127458 270
rect 127066 212 127143 268
rect 127199 212 127247 268
rect 127303 212 127351 268
rect 127407 214 127458 268
rect 127514 214 127562 270
rect 127618 214 127666 270
rect 127722 214 127773 270
rect 127829 214 127877 270
rect 127933 214 127981 270
rect 128037 214 128070 270
rect 127407 212 128070 214
rect 127066 166 128070 212
rect 127066 164 127458 166
rect 127066 108 127143 164
rect 127199 108 127247 164
rect 127303 108 127351 164
rect 127407 110 127458 164
rect 127514 110 127562 166
rect 127618 110 127666 166
rect 127722 110 127773 166
rect 127829 110 127877 166
rect 127933 110 127981 166
rect 128037 110 128070 166
rect 127407 108 128070 110
rect 127066 62 128070 108
rect 127066 60 127458 62
rect 127066 4 127143 60
rect 127199 4 127247 60
rect 127303 4 127351 60
rect 127407 6 127458 60
rect 127514 6 127562 62
rect 127618 6 127666 62
rect 127722 6 127773 62
rect 127829 6 127877 62
rect 127933 6 127981 62
rect 128037 6 128070 62
rect 127407 4 128070 6
rect 127066 -39 128070 4
rect 115944 -123 116895 -97
rect 115944 -125 116290 -123
rect 115944 -181 115975 -125
rect 116031 -181 116079 -125
rect 116135 -181 116183 -125
rect 116239 -179 116290 -125
rect 116346 -179 116394 -123
rect 116450 -179 116498 -123
rect 116554 -179 116605 -123
rect 116661 -179 116709 -123
rect 116765 -179 116813 -123
rect 116869 -179 116895 -123
rect 116239 -181 116895 -179
rect 115944 -227 116895 -181
rect 115944 -229 116290 -227
rect 115944 -285 115975 -229
rect 116031 -285 116079 -229
rect 116135 -285 116183 -229
rect 116239 -283 116290 -229
rect 116346 -283 116394 -227
rect 116450 -283 116498 -227
rect 116554 -283 116605 -227
rect 116661 -283 116709 -227
rect 116765 -283 116813 -227
rect 116869 -283 116895 -227
rect 116239 -285 116895 -283
rect 115944 -331 116895 -285
rect 115944 -333 116290 -331
rect 115944 -389 115975 -333
rect 116031 -389 116079 -333
rect 116135 -389 116183 -333
rect 116239 -387 116290 -333
rect 116346 -387 116394 -331
rect 116450 -387 116498 -331
rect 116554 -387 116605 -331
rect 116661 -387 116709 -331
rect 116765 -387 116813 -331
rect 116869 -387 116895 -331
rect 116239 -389 116895 -387
rect 115944 -423 116895 -389
rect 133936 -568 134096 2329
rect 133906 -588 134342 -568
rect 133906 -644 133929 -588
rect 133985 -644 134033 -588
rect 134089 -591 134342 -588
rect 134089 -644 134165 -591
rect 133906 -647 134165 -644
rect 134221 -647 134269 -591
rect 134325 -647 134342 -591
rect 133906 -692 134342 -647
rect 133906 -748 133929 -692
rect 133985 -748 134033 -692
rect 134089 -695 134342 -692
rect 134089 -748 134165 -695
rect 133906 -751 134165 -748
rect 134221 -751 134269 -695
rect 134325 -751 134342 -695
rect 133906 -765 134342 -751
rect 121366 -3234 122116 -3222
rect 121366 -3241 121943 -3234
rect 121366 -3293 121385 -3241
rect 121437 -3293 121489 -3241
rect 121541 -3286 121943 -3241
rect 121995 -3286 122047 -3234
rect 122099 -3286 122116 -3234
rect 121541 -3293 122116 -3286
rect 121366 -3338 122116 -3293
rect 121366 -3345 121943 -3338
rect 121366 -3397 121385 -3345
rect 121437 -3397 121489 -3345
rect 121541 -3390 121943 -3345
rect 121995 -3390 122047 -3338
rect 122099 -3390 122116 -3338
rect 121541 -3397 122116 -3390
rect 121366 -3410 122116 -3397
rect 122319 -3240 122556 -3222
rect 122319 -3307 122342 -3240
rect 122406 -3245 122556 -3240
rect 122406 -3307 122474 -3245
rect 122319 -3312 122474 -3307
rect 122538 -3312 122556 -3245
rect 122319 -3364 122556 -3312
rect 122319 -3365 122472 -3364
rect 122319 -3432 122347 -3365
rect 122411 -3431 122472 -3365
rect 122536 -3431 122556 -3364
rect 122411 -3432 122556 -3431
rect 122319 -3466 122556 -3432
rect 121003 -3877 121260 -3833
rect 121003 -3880 121167 -3877
rect 121003 -3946 121036 -3880
rect 121102 -3943 121167 -3880
rect 121233 -3943 121260 -3877
rect 121102 -3946 121260 -3943
rect 121003 -4009 121260 -3946
rect 121003 -4075 121035 -4009
rect 121101 -4075 121169 -4009
rect 121235 -4075 121260 -4009
rect 121003 -4137 121260 -4075
rect 121003 -4203 121032 -4137
rect 121098 -4203 121167 -4137
rect 121233 -4203 121260 -4137
rect 121003 -4274 121260 -4203
rect 121924 -4485 122674 -4472
rect 121924 -4537 121943 -4485
rect 121995 -4537 122047 -4485
rect 122099 -4492 122674 -4485
rect 122099 -4537 122501 -4492
rect 121924 -4544 122501 -4537
rect 122553 -4544 122605 -4492
rect 122657 -4544 122674 -4492
rect 121924 -4589 122674 -4544
rect 121924 -4641 121943 -4589
rect 121995 -4641 122047 -4589
rect 122099 -4596 122674 -4589
rect 122099 -4641 122501 -4596
rect 121924 -4648 122501 -4641
rect 122553 -4648 122605 -4596
rect 122657 -4648 122674 -4596
rect 121924 -4660 122674 -4648
rect 121601 -7081 122617 -7042
rect 121601 -7169 121627 -7081
rect 121714 -7169 121807 -7081
rect 121894 -7169 121973 -7081
rect 122060 -7169 122153 -7081
rect 122240 -7084 122617 -7081
rect 122240 -7169 122326 -7084
rect 121601 -7172 122326 -7169
rect 122413 -7172 122506 -7084
rect 122593 -7125 122617 -7084
rect 122593 -7172 124635 -7125
rect 121601 -7261 124635 -7172
rect 121601 -7349 121627 -7261
rect 121714 -7349 121807 -7261
rect 121894 -7349 121973 -7261
rect 122060 -7349 122153 -7261
rect 122240 -7264 124635 -7261
rect 122240 -7349 122326 -7264
rect 121601 -7352 122326 -7349
rect 122413 -7352 122506 -7264
rect 122593 -7325 124635 -7264
rect 122593 -7352 122617 -7325
rect 121601 -7381 122617 -7352
rect 145049 -8986 145105 -6615
rect 170266 -7085 171282 -7046
rect 170266 -7173 170292 -7085
rect 170379 -7173 170472 -7085
rect 170559 -7173 170638 -7085
rect 170725 -7173 170818 -7085
rect 170905 -7088 171282 -7085
rect 170905 -7173 170991 -7088
rect 170266 -7176 170991 -7173
rect 171078 -7176 171171 -7088
rect 171258 -7176 171282 -7088
rect 170266 -7265 171282 -7176
rect 170266 -7353 170292 -7265
rect 170379 -7353 170472 -7265
rect 170559 -7353 170638 -7265
rect 170725 -7353 170818 -7265
rect 170905 -7268 171282 -7265
rect 170905 -7353 170991 -7268
rect 170266 -7356 170991 -7353
rect 171078 -7356 171171 -7268
rect 171258 -7356 171282 -7268
rect 170266 -7385 171282 -7356
rect 144607 -9042 145105 -8986
rect 144607 -9351 144663 -9042
rect 144521 -12839 144771 -9351
rect 145185 -9361 145241 -7533
rect 146488 -8737 146600 -8532
rect 145819 -8792 146600 -8737
rect 145819 -8844 145860 -8792
rect 145912 -8844 145964 -8792
rect 146016 -8844 146068 -8792
rect 146120 -8844 146201 -8792
rect 146253 -8844 146305 -8792
rect 146357 -8844 146409 -8792
rect 146461 -8844 146600 -8792
rect 145819 -8896 146600 -8844
rect 145819 -8948 145860 -8896
rect 145912 -8948 145964 -8896
rect 146016 -8948 146068 -8896
rect 146120 -8948 146201 -8896
rect 146253 -8948 146305 -8896
rect 146357 -8948 146409 -8896
rect 146461 -8948 146600 -8896
rect 145819 -9000 146600 -8948
rect 145819 -9019 145860 -9000
rect 145749 -9052 145860 -9019
rect 145912 -9052 145964 -9000
rect 146016 -9052 146068 -9000
rect 146120 -9052 146201 -9000
rect 146253 -9052 146305 -9000
rect 146357 -9052 146409 -9000
rect 146461 -9052 146600 -9000
rect 145749 -9212 146600 -9052
rect 143034 -13089 144771 -12839
rect 133309 -13430 134166 -13357
rect 133309 -13431 134040 -13430
rect 133309 -13433 133706 -13431
rect 133309 -13521 133379 -13433
rect 133466 -13521 133559 -13433
rect 133646 -13519 133706 -13433
rect 133793 -13519 133886 -13431
rect 133973 -13518 134040 -13431
rect 134127 -13518 134166 -13430
rect 133973 -13519 134166 -13518
rect 133646 -13521 134166 -13519
rect 133309 -13610 134166 -13521
rect 133309 -13611 134040 -13610
rect 133309 -13613 133706 -13611
rect 133309 -13701 133379 -13613
rect 133466 -13701 133559 -13613
rect 133646 -13699 133706 -13613
rect 133793 -13699 133886 -13611
rect 133973 -13698 134040 -13611
rect 134127 -13698 134166 -13610
rect 133973 -13699 134166 -13698
rect 133646 -13701 134166 -13699
rect 115006 -13928 117188 -13734
rect 17492 -14949 20417 -14720
rect 16963 -15725 18346 -15496
rect 16080 -17003 16891 -16980
rect 18117 -16988 18346 -15725
rect 20188 -16964 20417 -14949
rect 75550 -14725 76478 -14704
rect 75550 -14813 75573 -14725
rect 75660 -14813 75733 -14725
rect 75820 -14813 75893 -14725
rect 75980 -14813 76053 -14725
rect 76140 -14813 76213 -14725
rect 76300 -14813 76373 -14725
rect 76460 -14813 76478 -14725
rect 75550 -14885 76478 -14813
rect 75550 -14973 75573 -14885
rect 75660 -14973 75733 -14885
rect 75820 -14973 75893 -14885
rect 75980 -14973 76053 -14885
rect 76140 -14973 76213 -14885
rect 76300 -14973 76373 -14885
rect 76460 -14973 76478 -14885
rect 75550 -15045 76478 -14973
rect 75550 -15133 75573 -15045
rect 75660 -15133 75733 -15045
rect 75820 -15133 75893 -15045
rect 75980 -15133 76053 -15045
rect 76140 -15133 76213 -15045
rect 76300 -15133 76373 -15045
rect 76460 -15133 76478 -15045
rect 75550 -15205 76478 -15133
rect 31520 -15275 32448 -15254
rect 29808 -15361 30736 -15340
rect 29808 -15449 29831 -15361
rect 29918 -15449 29991 -15361
rect 30078 -15449 30151 -15361
rect 30238 -15449 30311 -15361
rect 30398 -15449 30471 -15361
rect 30558 -15449 30631 -15361
rect 30718 -15449 30736 -15361
rect 27986 -15478 28914 -15457
rect 27986 -15566 28009 -15478
rect 28096 -15566 28169 -15478
rect 28256 -15566 28329 -15478
rect 28416 -15566 28489 -15478
rect 28576 -15566 28649 -15478
rect 28736 -15566 28809 -15478
rect 28896 -15566 28914 -15478
rect 27986 -15638 28914 -15566
rect 27986 -15726 28009 -15638
rect 28096 -15726 28169 -15638
rect 28256 -15726 28329 -15638
rect 28416 -15726 28489 -15638
rect 28576 -15726 28649 -15638
rect 28736 -15726 28809 -15638
rect 28896 -15726 28914 -15638
rect 27986 -15798 28914 -15726
rect 27986 -15886 28009 -15798
rect 28096 -15886 28169 -15798
rect 28256 -15886 28329 -15798
rect 28416 -15886 28489 -15798
rect 28576 -15886 28649 -15798
rect 28736 -15886 28809 -15798
rect 28896 -15886 28914 -15798
rect 27986 -15958 28914 -15886
rect 27986 -16046 28009 -15958
rect 28096 -16046 28169 -15958
rect 28256 -16046 28329 -15958
rect 28416 -16046 28489 -15958
rect 28576 -16046 28649 -15958
rect 28736 -16046 28809 -15958
rect 28896 -16046 28914 -15958
rect 27986 -16118 28914 -16046
rect 27986 -16206 28009 -16118
rect 28096 -16206 28169 -16118
rect 28256 -16206 28329 -16118
rect 28416 -16206 28489 -16118
rect 28576 -16206 28649 -16118
rect 28736 -16206 28809 -16118
rect 28896 -16206 28914 -16118
rect 27986 -16278 28914 -16206
rect 29808 -15521 30736 -15449
rect 29808 -15609 29831 -15521
rect 29918 -15609 29991 -15521
rect 30078 -15609 30151 -15521
rect 30238 -15609 30311 -15521
rect 30398 -15609 30471 -15521
rect 30558 -15609 30631 -15521
rect 30718 -15609 30736 -15521
rect 29808 -15681 30736 -15609
rect 29808 -15769 29831 -15681
rect 29918 -15769 29991 -15681
rect 30078 -15769 30151 -15681
rect 30238 -15769 30311 -15681
rect 30398 -15769 30471 -15681
rect 30558 -15769 30631 -15681
rect 30718 -15769 30736 -15681
rect 29808 -15841 30736 -15769
rect 29808 -15929 29831 -15841
rect 29918 -15929 29991 -15841
rect 30078 -15929 30151 -15841
rect 30238 -15929 30311 -15841
rect 30398 -15929 30471 -15841
rect 30558 -15929 30631 -15841
rect 30718 -15929 30736 -15841
rect 29808 -16001 30736 -15929
rect 29808 -16089 29831 -16001
rect 29918 -16089 29991 -16001
rect 30078 -16089 30151 -16001
rect 30238 -16089 30311 -16001
rect 30398 -16089 30471 -16001
rect 30558 -16089 30631 -16001
rect 30718 -16089 30736 -16001
rect 29808 -16161 30736 -16089
rect 29808 -16249 29831 -16161
rect 29918 -16249 29991 -16161
rect 30078 -16249 30151 -16161
rect 30238 -16249 30311 -16161
rect 30398 -16249 30471 -16161
rect 30558 -16249 30631 -16161
rect 30718 -16249 30736 -16161
rect 31520 -15363 31543 -15275
rect 31630 -15363 31703 -15275
rect 31790 -15363 31863 -15275
rect 31950 -15363 32023 -15275
rect 32110 -15363 32183 -15275
rect 32270 -15363 32343 -15275
rect 32430 -15363 32448 -15275
rect 31520 -15435 32448 -15363
rect 31520 -15523 31543 -15435
rect 31630 -15523 31703 -15435
rect 31790 -15523 31863 -15435
rect 31950 -15523 32023 -15435
rect 32110 -15523 32183 -15435
rect 32270 -15523 32343 -15435
rect 32430 -15523 32448 -15435
rect 31520 -15595 32448 -15523
rect 31520 -15683 31543 -15595
rect 31630 -15683 31703 -15595
rect 31790 -15683 31863 -15595
rect 31950 -15683 32023 -15595
rect 32110 -15683 32183 -15595
rect 32270 -15683 32343 -15595
rect 32430 -15683 32448 -15595
rect 75550 -15293 75573 -15205
rect 75660 -15293 75733 -15205
rect 75820 -15293 75893 -15205
rect 75980 -15293 76053 -15205
rect 76140 -15293 76213 -15205
rect 76300 -15293 76373 -15205
rect 76460 -15293 76478 -15205
rect 75550 -15365 76478 -15293
rect 75550 -15453 75573 -15365
rect 75660 -15453 75733 -15365
rect 75820 -15453 75893 -15365
rect 75980 -15453 76053 -15365
rect 76140 -15453 76213 -15365
rect 76300 -15453 76373 -15365
rect 76460 -15453 76478 -15365
rect 80725 -14936 81871 -14901
rect 80725 -14937 81435 -14936
rect 80725 -14939 81101 -14937
rect 80725 -15027 80774 -14939
rect 80861 -15027 80954 -14939
rect 81041 -15025 81101 -14939
rect 81188 -15025 81281 -14937
rect 81368 -15024 81435 -14937
rect 81522 -14938 81871 -14936
rect 81522 -14939 81759 -14938
rect 81522 -15024 81605 -14939
rect 81368 -15025 81605 -15024
rect 81041 -15027 81605 -15025
rect 81692 -15026 81759 -14939
rect 81846 -15026 81871 -14938
rect 81692 -15027 81871 -15026
rect 80725 -15116 81871 -15027
rect 80725 -15117 81435 -15116
rect 80725 -15119 81101 -15117
rect 80725 -15207 80774 -15119
rect 80861 -15207 80954 -15119
rect 81041 -15205 81101 -15119
rect 81188 -15205 81281 -15117
rect 81368 -15204 81435 -15117
rect 81522 -15118 81871 -15116
rect 81522 -15119 81759 -15118
rect 81522 -15204 81605 -15119
rect 81368 -15205 81605 -15204
rect 81041 -15207 81605 -15205
rect 81692 -15206 81759 -15119
rect 81846 -15206 81871 -15118
rect 81692 -15207 81871 -15206
rect 80725 -15293 81871 -15207
rect 80725 -15294 81429 -15293
rect 80725 -15296 81095 -15294
rect 80725 -15384 80768 -15296
rect 80855 -15384 80948 -15296
rect 81035 -15382 81095 -15296
rect 81182 -15382 81275 -15294
rect 81362 -15381 81429 -15294
rect 81516 -15295 81871 -15293
rect 81516 -15296 81753 -15295
rect 81516 -15381 81599 -15296
rect 81362 -15382 81599 -15381
rect 81035 -15384 81599 -15382
rect 81686 -15383 81753 -15296
rect 81840 -15383 81871 -15295
rect 81686 -15384 81871 -15383
rect 80725 -15423 81871 -15384
rect 75550 -15525 76478 -15453
rect 75550 -15613 75573 -15525
rect 75660 -15613 75733 -15525
rect 75820 -15613 75893 -15525
rect 75980 -15613 76053 -15525
rect 76140 -15613 76213 -15525
rect 76300 -15613 76373 -15525
rect 76460 -15613 76478 -15525
rect 75550 -15635 76478 -15613
rect 113311 -15672 113505 -13942
rect 31520 -15755 32448 -15683
rect 31520 -15843 31543 -15755
rect 31630 -15843 31703 -15755
rect 31790 -15843 31863 -15755
rect 31950 -15843 32023 -15755
rect 32110 -15843 32183 -15755
rect 32270 -15843 32343 -15755
rect 32430 -15843 32448 -15755
rect 31520 -15915 32448 -15843
rect 31520 -16003 31543 -15915
rect 31630 -16003 31703 -15915
rect 31790 -16003 31863 -15915
rect 31950 -16003 32023 -15915
rect 32110 -16003 32183 -15915
rect 32270 -16003 32343 -15915
rect 32430 -16003 32448 -15915
rect 112965 -15695 113776 -15672
rect 112965 -15778 112989 -15695
rect 113072 -15778 113159 -15695
rect 113242 -15778 113329 -15695
rect 113412 -15778 113499 -15695
rect 113582 -15778 113669 -15695
rect 113752 -15778 113776 -15695
rect 116994 -15707 117188 -13928
rect 133309 -13823 134166 -13701
rect 133309 -13824 134022 -13823
rect 133309 -13826 133688 -13824
rect 133309 -13914 133361 -13826
rect 133448 -13914 133541 -13826
rect 133628 -13912 133688 -13826
rect 133775 -13912 133868 -13824
rect 133955 -13911 134022 -13824
rect 134109 -13911 134166 -13823
rect 133955 -13912 134166 -13911
rect 133628 -13914 134166 -13912
rect 133309 -14003 134166 -13914
rect 133309 -14004 134022 -14003
rect 133309 -14006 133688 -14004
rect 133309 -14094 133361 -14006
rect 133448 -14094 133541 -14006
rect 133628 -14092 133688 -14006
rect 133775 -14092 133868 -14004
rect 133955 -14091 134022 -14004
rect 134109 -14091 134166 -14003
rect 133955 -14092 134166 -14091
rect 133628 -14094 134166 -14092
rect 133309 -14172 134166 -14094
rect 135747 -13435 136604 -13362
rect 135747 -13436 136478 -13435
rect 135747 -13438 136144 -13436
rect 135747 -13526 135817 -13438
rect 135904 -13526 135997 -13438
rect 136084 -13524 136144 -13438
rect 136231 -13524 136324 -13436
rect 136411 -13523 136478 -13436
rect 136565 -13523 136604 -13435
rect 136411 -13524 136604 -13523
rect 136084 -13526 136604 -13524
rect 135747 -13615 136604 -13526
rect 135747 -13616 136478 -13615
rect 135747 -13618 136144 -13616
rect 135747 -13706 135817 -13618
rect 135904 -13706 135997 -13618
rect 136084 -13704 136144 -13618
rect 136231 -13704 136324 -13616
rect 136411 -13703 136478 -13616
rect 136565 -13703 136604 -13615
rect 136411 -13704 136604 -13703
rect 136084 -13706 136604 -13704
rect 135747 -13828 136604 -13706
rect 135747 -13829 136460 -13828
rect 135747 -13831 136126 -13829
rect 135747 -13919 135799 -13831
rect 135886 -13919 135979 -13831
rect 136066 -13917 136126 -13831
rect 136213 -13917 136306 -13829
rect 136393 -13916 136460 -13829
rect 136547 -13916 136604 -13828
rect 136393 -13917 136604 -13916
rect 136066 -13919 136604 -13917
rect 135747 -14008 136604 -13919
rect 135747 -14009 136460 -14008
rect 135747 -14011 136126 -14009
rect 135747 -14099 135799 -14011
rect 135886 -14099 135979 -14011
rect 136066 -14097 136126 -14011
rect 136213 -14097 136306 -14009
rect 136393 -14096 136460 -14009
rect 136547 -14096 136604 -14008
rect 136393 -14097 136604 -14096
rect 136066 -14099 136604 -14097
rect 135747 -14177 136604 -14099
rect 138469 -13441 139326 -13368
rect 138469 -13442 139200 -13441
rect 138469 -13444 138866 -13442
rect 138469 -13532 138539 -13444
rect 138626 -13532 138719 -13444
rect 138806 -13530 138866 -13444
rect 138953 -13530 139046 -13442
rect 139133 -13529 139200 -13442
rect 139287 -13529 139326 -13441
rect 139133 -13530 139326 -13529
rect 138806 -13532 139326 -13530
rect 138469 -13621 139326 -13532
rect 138469 -13622 139200 -13621
rect 138469 -13624 138866 -13622
rect 138469 -13712 138539 -13624
rect 138626 -13712 138719 -13624
rect 138806 -13710 138866 -13624
rect 138953 -13710 139046 -13622
rect 139133 -13709 139200 -13622
rect 139287 -13709 139326 -13621
rect 139133 -13710 139326 -13709
rect 138806 -13712 139326 -13710
rect 138469 -13834 139326 -13712
rect 138469 -13835 139182 -13834
rect 138469 -13837 138848 -13835
rect 138469 -13925 138521 -13837
rect 138608 -13925 138701 -13837
rect 138788 -13923 138848 -13837
rect 138935 -13923 139028 -13835
rect 139115 -13922 139182 -13835
rect 139269 -13922 139326 -13834
rect 139115 -13923 139326 -13922
rect 138788 -13925 139326 -13923
rect 138469 -14014 139326 -13925
rect 138469 -14015 139182 -14014
rect 138469 -14017 138848 -14015
rect 138469 -14105 138521 -14017
rect 138608 -14105 138701 -14017
rect 138788 -14103 138848 -14017
rect 138935 -14103 139028 -14015
rect 139115 -14102 139182 -14015
rect 139269 -14102 139326 -14014
rect 139115 -14103 139326 -14102
rect 138788 -14105 139326 -14103
rect 138469 -14183 139326 -14105
rect 143034 -14930 143284 -13089
rect 145106 -14908 145356 -9361
rect 145749 -13604 146527 -9212
rect 147149 -9319 147205 -7969
rect 145749 -13656 145840 -13604
rect 145892 -13656 145944 -13604
rect 145996 -13656 146048 -13604
rect 146100 -13656 146181 -13604
rect 146233 -13656 146285 -13604
rect 146337 -13656 146389 -13604
rect 146441 -13656 146527 -13604
rect 145749 -13708 146527 -13656
rect 145749 -13760 145840 -13708
rect 145892 -13760 145944 -13708
rect 145996 -13760 146048 -13708
rect 146100 -13760 146181 -13708
rect 146233 -13760 146285 -13708
rect 146337 -13760 146389 -13708
rect 146441 -13760 146527 -13708
rect 145749 -13812 146527 -13760
rect 145749 -13864 145840 -13812
rect 145892 -13864 145944 -13812
rect 145996 -13864 146048 -13812
rect 146100 -13864 146181 -13812
rect 146233 -13864 146285 -13812
rect 146337 -13864 146389 -13812
rect 146441 -13864 146527 -13812
rect 145749 -13890 146527 -13864
rect 147122 -14887 147372 -9319
rect 150251 -13408 151108 -13335
rect 150251 -13409 150982 -13408
rect 150251 -13411 150648 -13409
rect 150251 -13499 150321 -13411
rect 150408 -13499 150501 -13411
rect 150588 -13497 150648 -13411
rect 150735 -13497 150828 -13409
rect 150915 -13496 150982 -13409
rect 151069 -13496 151108 -13408
rect 150915 -13497 151108 -13496
rect 150588 -13499 151108 -13497
rect 150251 -13588 151108 -13499
rect 150251 -13589 150982 -13588
rect 150251 -13591 150648 -13589
rect 150251 -13679 150321 -13591
rect 150408 -13679 150501 -13591
rect 150588 -13677 150648 -13591
rect 150735 -13677 150828 -13589
rect 150915 -13676 150982 -13589
rect 151069 -13676 151108 -13588
rect 150915 -13677 151108 -13676
rect 150588 -13679 151108 -13677
rect 150251 -13801 151108 -13679
rect 150251 -13802 150964 -13801
rect 150251 -13804 150630 -13802
rect 150251 -13892 150303 -13804
rect 150390 -13892 150483 -13804
rect 150570 -13890 150630 -13804
rect 150717 -13890 150810 -13802
rect 150897 -13889 150964 -13802
rect 151051 -13889 151108 -13801
rect 150897 -13890 151108 -13889
rect 150570 -13892 151108 -13890
rect 150251 -13981 151108 -13892
rect 150251 -13982 150964 -13981
rect 150251 -13984 150630 -13982
rect 150251 -14072 150303 -13984
rect 150390 -14072 150483 -13984
rect 150570 -14070 150630 -13984
rect 150717 -14070 150810 -13982
rect 150897 -14069 150964 -13982
rect 151051 -14069 151108 -13981
rect 150897 -14070 151108 -14069
rect 150570 -14072 151108 -14070
rect 150251 -14150 151108 -14072
rect 142756 -14953 143567 -14930
rect 142756 -15036 142780 -14953
rect 142863 -15036 142950 -14953
rect 143033 -15036 143120 -14953
rect 143203 -15036 143290 -14953
rect 143373 -15036 143460 -14953
rect 143543 -15036 143567 -14953
rect 142756 -15123 143567 -15036
rect 142756 -15206 142780 -15123
rect 142863 -15206 142950 -15123
rect 143033 -15206 143120 -15123
rect 143203 -15206 143290 -15123
rect 143373 -15206 143460 -15123
rect 143543 -15206 143567 -15123
rect 142756 -15293 143567 -15206
rect 142756 -15376 142780 -15293
rect 142863 -15376 142950 -15293
rect 143033 -15376 143120 -15293
rect 143203 -15376 143290 -15293
rect 143373 -15376 143460 -15293
rect 143543 -15376 143567 -15293
rect 142756 -15463 143567 -15376
rect 142756 -15546 142780 -15463
rect 142863 -15546 142950 -15463
rect 143033 -15546 143120 -15463
rect 143203 -15546 143290 -15463
rect 143373 -15546 143460 -15463
rect 143543 -15546 143567 -15463
rect 142756 -15633 143567 -15546
rect 112965 -15865 113776 -15778
rect 80861 -15965 81789 -15944
rect 31520 -16075 32448 -16003
rect 31520 -16163 31543 -16075
rect 31630 -16163 31703 -16075
rect 31790 -16163 31863 -16075
rect 31950 -16163 32023 -16075
rect 32110 -16163 32183 -16075
rect 32270 -16163 32343 -16075
rect 32430 -16163 32448 -16075
rect 31520 -16185 32448 -16163
rect 65068 -16002 65879 -15979
rect 65068 -16085 65092 -16002
rect 65175 -16085 65262 -16002
rect 65345 -16085 65432 -16002
rect 65515 -16085 65602 -16002
rect 65685 -16085 65772 -16002
rect 65855 -16085 65879 -16002
rect 65068 -16172 65879 -16085
rect 29808 -16271 30736 -16249
rect 65068 -16255 65092 -16172
rect 65175 -16255 65262 -16172
rect 65345 -16255 65432 -16172
rect 65515 -16255 65602 -16172
rect 65685 -16255 65772 -16172
rect 65855 -16255 65879 -16172
rect 80861 -16053 80884 -15965
rect 80971 -16053 81044 -15965
rect 81131 -16053 81204 -15965
rect 81291 -16053 81364 -15965
rect 81451 -16053 81524 -15965
rect 81611 -16053 81684 -15965
rect 81771 -16053 81789 -15965
rect 80861 -16125 81789 -16053
rect 27986 -16366 28009 -16278
rect 28096 -16366 28169 -16278
rect 28256 -16366 28329 -16278
rect 28416 -16366 28489 -16278
rect 28576 -16366 28649 -16278
rect 28736 -16366 28809 -16278
rect 28896 -16366 28914 -16278
rect 27986 -16388 28914 -16366
rect 65068 -16342 65879 -16255
rect 65068 -16425 65092 -16342
rect 65175 -16425 65262 -16342
rect 65345 -16425 65432 -16342
rect 65515 -16425 65602 -16342
rect 65685 -16425 65772 -16342
rect 65855 -16425 65879 -16342
rect 65068 -16512 65879 -16425
rect 65068 -16595 65092 -16512
rect 65175 -16595 65262 -16512
rect 65345 -16595 65432 -16512
rect 65515 -16595 65602 -16512
rect 65685 -16595 65772 -16512
rect 65855 -16595 65879 -16512
rect 65068 -16682 65879 -16595
rect 65068 -16765 65092 -16682
rect 65175 -16765 65262 -16682
rect 65345 -16765 65432 -16682
rect 65515 -16765 65602 -16682
rect 65685 -16765 65772 -16682
rect 65855 -16765 65879 -16682
rect 65068 -16788 65879 -16765
rect 75576 -16264 76755 -16205
rect 75576 -16265 76313 -16264
rect 75576 -16267 75979 -16265
rect 75576 -16355 75652 -16267
rect 75739 -16355 75832 -16267
rect 75919 -16353 75979 -16267
rect 76066 -16353 76159 -16265
rect 76246 -16352 76313 -16265
rect 76400 -16266 76755 -16264
rect 76400 -16267 76637 -16266
rect 76400 -16352 76483 -16267
rect 76246 -16353 76483 -16352
rect 75919 -16355 76483 -16353
rect 76570 -16354 76637 -16267
rect 76724 -16354 76755 -16266
rect 76570 -16355 76755 -16354
rect 75576 -16444 76755 -16355
rect 75576 -16445 76313 -16444
rect 75576 -16447 75979 -16445
rect 75576 -16535 75652 -16447
rect 75739 -16535 75832 -16447
rect 75919 -16533 75979 -16447
rect 76066 -16533 76159 -16445
rect 76246 -16532 76313 -16445
rect 76400 -16446 76755 -16444
rect 76400 -16447 76637 -16446
rect 76400 -16532 76483 -16447
rect 76246 -16533 76483 -16532
rect 75919 -16535 76483 -16533
rect 76570 -16534 76637 -16447
rect 76724 -16534 76755 -16446
rect 76570 -16535 76755 -16534
rect 75576 -16621 76755 -16535
rect 75576 -16622 76307 -16621
rect 75576 -16624 75973 -16622
rect 75576 -16712 75646 -16624
rect 75733 -16712 75826 -16624
rect 75913 -16710 75973 -16624
rect 76060 -16710 76153 -16622
rect 76240 -16709 76307 -16622
rect 76394 -16623 76755 -16621
rect 76394 -16624 76631 -16623
rect 76394 -16709 76477 -16624
rect 76240 -16710 76477 -16709
rect 75913 -16712 76477 -16710
rect 76564 -16711 76631 -16624
rect 76718 -16711 76755 -16623
rect 76564 -16712 76755 -16711
rect 75576 -16768 76755 -16712
rect 80861 -16213 80884 -16125
rect 80971 -16213 81044 -16125
rect 81131 -16213 81204 -16125
rect 81291 -16213 81364 -16125
rect 81451 -16213 81524 -16125
rect 81611 -16213 81684 -16125
rect 81771 -16213 81789 -16125
rect 80861 -16285 81789 -16213
rect 80861 -16373 80884 -16285
rect 80971 -16373 81044 -16285
rect 81131 -16373 81204 -16285
rect 81291 -16373 81364 -16285
rect 81451 -16373 81524 -16285
rect 81611 -16373 81684 -16285
rect 81771 -16373 81789 -16285
rect 80861 -16445 81789 -16373
rect 80861 -16533 80884 -16445
rect 80971 -16533 81044 -16445
rect 81131 -16533 81204 -16445
rect 81291 -16533 81364 -16445
rect 81451 -16533 81524 -16445
rect 81611 -16533 81684 -16445
rect 81771 -16533 81789 -16445
rect 112965 -15948 112989 -15865
rect 113072 -15948 113159 -15865
rect 113242 -15948 113329 -15865
rect 113412 -15948 113499 -15865
rect 113582 -15948 113669 -15865
rect 113752 -15948 113776 -15865
rect 112965 -16035 113776 -15948
rect 112965 -16118 112989 -16035
rect 113072 -16118 113159 -16035
rect 113242 -16118 113329 -16035
rect 113412 -16118 113499 -16035
rect 113582 -16118 113669 -16035
rect 113752 -16118 113776 -16035
rect 112965 -16205 113776 -16118
rect 112965 -16288 112989 -16205
rect 113072 -16288 113159 -16205
rect 113242 -16288 113329 -16205
rect 113412 -16288 113499 -16205
rect 113582 -16288 113669 -16205
rect 113752 -16288 113776 -16205
rect 112965 -16375 113776 -16288
rect 112965 -16458 112989 -16375
rect 113072 -16458 113159 -16375
rect 113242 -16458 113329 -16375
rect 113412 -16458 113499 -16375
rect 113582 -16458 113669 -16375
rect 113752 -16458 113776 -16375
rect 112965 -16481 113776 -16458
rect 116695 -15730 117506 -15707
rect 116695 -15813 116719 -15730
rect 116802 -15813 116889 -15730
rect 116972 -15813 117059 -15730
rect 117142 -15813 117229 -15730
rect 117312 -15813 117399 -15730
rect 117482 -15813 117506 -15730
rect 142756 -15716 142780 -15633
rect 142863 -15716 142950 -15633
rect 143033 -15716 143120 -15633
rect 143203 -15716 143290 -15633
rect 143373 -15716 143460 -15633
rect 143543 -15716 143567 -15633
rect 142756 -15739 143567 -15716
rect 144802 -14931 145613 -14908
rect 144802 -15014 144826 -14931
rect 144909 -15014 144996 -14931
rect 145079 -15014 145166 -14931
rect 145249 -15014 145336 -14931
rect 145419 -15014 145506 -14931
rect 145589 -15014 145613 -14931
rect 144802 -15101 145613 -15014
rect 144802 -15184 144826 -15101
rect 144909 -15184 144996 -15101
rect 145079 -15184 145166 -15101
rect 145249 -15184 145336 -15101
rect 145419 -15184 145506 -15101
rect 145589 -15184 145613 -15101
rect 144802 -15271 145613 -15184
rect 144802 -15354 144826 -15271
rect 144909 -15354 144996 -15271
rect 145079 -15354 145166 -15271
rect 145249 -15354 145336 -15271
rect 145419 -15354 145506 -15271
rect 145589 -15354 145613 -15271
rect 144802 -15441 145613 -15354
rect 144802 -15524 144826 -15441
rect 144909 -15524 144996 -15441
rect 145079 -15524 145166 -15441
rect 145249 -15524 145336 -15441
rect 145419 -15524 145506 -15441
rect 145589 -15524 145613 -15441
rect 144802 -15611 145613 -15524
rect 144802 -15694 144826 -15611
rect 144909 -15694 144996 -15611
rect 145079 -15694 145166 -15611
rect 145249 -15694 145336 -15611
rect 145419 -15694 145506 -15611
rect 145589 -15694 145613 -15611
rect 144802 -15717 145613 -15694
rect 146936 -14910 147747 -14887
rect 146936 -14993 146960 -14910
rect 147043 -14993 147130 -14910
rect 147213 -14993 147300 -14910
rect 147383 -14993 147470 -14910
rect 147553 -14993 147640 -14910
rect 147723 -14993 147747 -14910
rect 146936 -15080 147747 -14993
rect 146936 -15163 146960 -15080
rect 147043 -15163 147130 -15080
rect 147213 -15163 147300 -15080
rect 147383 -15163 147470 -15080
rect 147553 -15163 147640 -15080
rect 147723 -15163 147747 -15080
rect 146936 -15250 147747 -15163
rect 146936 -15333 146960 -15250
rect 147043 -15333 147130 -15250
rect 147213 -15333 147300 -15250
rect 147383 -15333 147470 -15250
rect 147553 -15333 147640 -15250
rect 147723 -15333 147747 -15250
rect 146936 -15420 147747 -15333
rect 146936 -15503 146960 -15420
rect 147043 -15503 147130 -15420
rect 147213 -15503 147300 -15420
rect 147383 -15503 147470 -15420
rect 147553 -15503 147640 -15420
rect 147723 -15503 147747 -15420
rect 146936 -15590 147747 -15503
rect 146936 -15673 146960 -15590
rect 147043 -15673 147130 -15590
rect 147213 -15673 147300 -15590
rect 147383 -15673 147470 -15590
rect 147553 -15673 147640 -15590
rect 147723 -15673 147747 -15590
rect 146936 -15696 147747 -15673
rect 116695 -15900 117506 -15813
rect 116695 -15983 116719 -15900
rect 116802 -15983 116889 -15900
rect 116972 -15983 117059 -15900
rect 117142 -15983 117229 -15900
rect 117312 -15983 117399 -15900
rect 117482 -15983 117506 -15900
rect 116695 -16070 117506 -15983
rect 116695 -16153 116719 -16070
rect 116802 -16153 116889 -16070
rect 116972 -16153 117059 -16070
rect 117142 -16153 117229 -16070
rect 117312 -16153 117399 -16070
rect 117482 -16153 117506 -16070
rect 116695 -16240 117506 -16153
rect 116695 -16323 116719 -16240
rect 116802 -16323 116889 -16240
rect 116972 -16323 117059 -16240
rect 117142 -16323 117229 -16240
rect 117312 -16323 117399 -16240
rect 117482 -16323 117506 -16240
rect 116695 -16410 117506 -16323
rect 116695 -16493 116719 -16410
rect 116802 -16493 116889 -16410
rect 116972 -16493 117059 -16410
rect 117142 -16493 117229 -16410
rect 117312 -16493 117399 -16410
rect 117482 -16493 117506 -16410
rect 116695 -16516 117506 -16493
rect 80861 -16605 81789 -16533
rect 80861 -16693 80884 -16605
rect 80971 -16693 81044 -16605
rect 81131 -16693 81204 -16605
rect 81291 -16693 81364 -16605
rect 81451 -16693 81524 -16605
rect 81611 -16693 81684 -16605
rect 81771 -16693 81789 -16605
rect 80861 -16765 81789 -16693
rect 80861 -16853 80884 -16765
rect 80971 -16853 81044 -16765
rect 81131 -16853 81204 -16765
rect 81291 -16853 81364 -16765
rect 81451 -16853 81524 -16765
rect 81611 -16853 81684 -16765
rect 81771 -16853 81789 -16765
rect 80861 -16875 81789 -16853
rect 20058 -16987 20869 -16964
rect 16080 -17086 16104 -17003
rect 16187 -17086 16274 -17003
rect 16357 -17086 16444 -17003
rect 16527 -17086 16614 -17003
rect 16697 -17086 16784 -17003
rect 16867 -17086 16891 -17003
rect 16080 -17173 16891 -17086
rect -5122 -17229 -4313 -17205
rect -5122 -17312 -5099 -17229
rect -5016 -17312 -4929 -17229
rect -4846 -17312 -4759 -17229
rect -4676 -17312 -4589 -17229
rect -4506 -17312 -4419 -17229
rect -4336 -17312 -4313 -17229
rect -5122 -17399 -4313 -17312
rect -5122 -17482 -5099 -17399
rect -5016 -17482 -4929 -17399
rect -4846 -17482 -4759 -17399
rect -4676 -17482 -4589 -17399
rect -4506 -17482 -4419 -17399
rect -4336 -17482 -4313 -17399
rect -5122 -17496 -4313 -17482
rect 16080 -17256 16104 -17173
rect 16187 -17256 16274 -17173
rect 16357 -17256 16444 -17173
rect 16527 -17256 16614 -17173
rect 16697 -17256 16784 -17173
rect 16867 -17256 16891 -17173
rect 16080 -17343 16891 -17256
rect 16080 -17426 16104 -17343
rect 16187 -17426 16274 -17343
rect 16357 -17426 16444 -17343
rect 16527 -17426 16614 -17343
rect 16697 -17426 16784 -17343
rect 16867 -17426 16891 -17343
rect -5122 -17524 -817 -17496
rect -5122 -17569 -1129 -17524
rect -5122 -17652 -5099 -17569
rect -5016 -17652 -4929 -17569
rect -4846 -17652 -4759 -17569
rect -4676 -17652 -4589 -17569
rect -4506 -17652 -4419 -17569
rect -4336 -17580 -1129 -17569
rect -1073 -17580 -1025 -17524
rect -969 -17580 -921 -17524
rect -865 -17580 -817 -17524
rect -4336 -17628 -817 -17580
rect -4336 -17652 -1129 -17628
rect -5122 -17684 -1129 -17652
rect -1073 -17684 -1025 -17628
rect -969 -17684 -921 -17628
rect -865 -17684 -817 -17628
rect -5122 -17732 -817 -17684
rect -5122 -17739 -1129 -17732
rect -5122 -17822 -5099 -17739
rect -5016 -17822 -4929 -17739
rect -4846 -17822 -4759 -17739
rect -4676 -17822 -4589 -17739
rect -4506 -17822 -4419 -17739
rect -4336 -17788 -1129 -17739
rect -1073 -17788 -1025 -17732
rect -969 -17788 -921 -17732
rect -865 -17788 -817 -17732
rect -4336 -17814 -817 -17788
rect 16080 -17513 16891 -17426
rect 16080 -17596 16104 -17513
rect 16187 -17596 16274 -17513
rect 16357 -17596 16444 -17513
rect 16527 -17596 16614 -17513
rect 16697 -17596 16784 -17513
rect 16867 -17596 16891 -17513
rect 16080 -17683 16891 -17596
rect 16080 -17766 16104 -17683
rect 16187 -17766 16274 -17683
rect 16357 -17766 16444 -17683
rect 16527 -17766 16614 -17683
rect 16697 -17766 16784 -17683
rect 16867 -17766 16891 -17683
rect 16080 -17789 16891 -17766
rect 17986 -17011 18797 -16988
rect 17986 -17094 18010 -17011
rect 18093 -17094 18180 -17011
rect 18263 -17094 18350 -17011
rect 18433 -17094 18520 -17011
rect 18603 -17094 18690 -17011
rect 18773 -17094 18797 -17011
rect 17986 -17181 18797 -17094
rect 17986 -17264 18010 -17181
rect 18093 -17264 18180 -17181
rect 18263 -17264 18350 -17181
rect 18433 -17264 18520 -17181
rect 18603 -17264 18690 -17181
rect 18773 -17264 18797 -17181
rect 17986 -17351 18797 -17264
rect 17986 -17434 18010 -17351
rect 18093 -17434 18180 -17351
rect 18263 -17434 18350 -17351
rect 18433 -17434 18520 -17351
rect 18603 -17434 18690 -17351
rect 18773 -17434 18797 -17351
rect 17986 -17521 18797 -17434
rect 17986 -17604 18010 -17521
rect 18093 -17604 18180 -17521
rect 18263 -17604 18350 -17521
rect 18433 -17604 18520 -17521
rect 18603 -17604 18690 -17521
rect 18773 -17604 18797 -17521
rect 17986 -17691 18797 -17604
rect 17986 -17774 18010 -17691
rect 18093 -17774 18180 -17691
rect 18263 -17774 18350 -17691
rect 18433 -17774 18520 -17691
rect 18603 -17774 18690 -17691
rect 18773 -17774 18797 -17691
rect 20058 -17070 20082 -16987
rect 20165 -17070 20252 -16987
rect 20335 -17070 20422 -16987
rect 20505 -17070 20592 -16987
rect 20675 -17070 20762 -16987
rect 20845 -17070 20869 -16987
rect 20058 -17157 20869 -17070
rect 20058 -17240 20082 -17157
rect 20165 -17240 20252 -17157
rect 20335 -17240 20422 -17157
rect 20505 -17240 20592 -17157
rect 20675 -17240 20762 -17157
rect 20845 -17240 20869 -17157
rect 20058 -17327 20869 -17240
rect 20058 -17410 20082 -17327
rect 20165 -17410 20252 -17327
rect 20335 -17410 20422 -17327
rect 20505 -17410 20592 -17327
rect 20675 -17410 20762 -17327
rect 20845 -17410 20869 -17327
rect 20058 -17497 20869 -17410
rect 20058 -17580 20082 -17497
rect 20165 -17580 20252 -17497
rect 20335 -17580 20422 -17497
rect 20505 -17580 20592 -17497
rect 20675 -17580 20762 -17497
rect 20845 -17580 20869 -17497
rect 20058 -17667 20869 -17580
rect 20058 -17750 20082 -17667
rect 20165 -17750 20252 -17667
rect 20335 -17750 20422 -17667
rect 20505 -17750 20592 -17667
rect 20675 -17750 20762 -17667
rect 20845 -17750 20869 -17667
rect 20058 -17773 20869 -17750
rect 17986 -17797 18797 -17774
rect -4336 -17822 -4313 -17814
rect -5122 -17909 -4313 -17822
rect -5122 -17992 -5099 -17909
rect -5016 -17992 -4929 -17909
rect -4846 -17992 -4759 -17909
rect -4676 -17992 -4589 -17909
rect -4506 -17992 -4419 -17909
rect -4336 -17992 -4313 -17909
rect -5122 -18016 -4313 -17992
rect 27267 -18163 28195 -18142
rect 27267 -18251 27290 -18163
rect 27377 -18251 27450 -18163
rect 27537 -18251 27610 -18163
rect 27697 -18251 27770 -18163
rect 27857 -18251 27930 -18163
rect 28017 -18251 28090 -18163
rect 28177 -18251 28195 -18163
rect 27267 -18323 28195 -18251
rect 288 -18349 1099 -18326
rect 288 -18432 312 -18349
rect 395 -18432 482 -18349
rect 565 -18432 652 -18349
rect 735 -18432 822 -18349
rect 905 -18432 992 -18349
rect 1075 -18432 1099 -18349
rect 288 -18519 1099 -18432
rect 288 -18602 312 -18519
rect 395 -18602 482 -18519
rect 565 -18602 652 -18519
rect 735 -18602 822 -18519
rect 905 -18602 992 -18519
rect 1075 -18602 1099 -18519
rect 288 -18689 1099 -18602
rect 288 -18772 312 -18689
rect 395 -18772 482 -18689
rect 565 -18772 652 -18689
rect 735 -18772 822 -18689
rect 905 -18772 992 -18689
rect 1075 -18772 1099 -18689
rect 288 -18859 1099 -18772
rect 288 -18942 312 -18859
rect 395 -18942 482 -18859
rect 565 -18942 652 -18859
rect 735 -18942 822 -18859
rect 905 -18942 992 -18859
rect 1075 -18942 1099 -18859
rect 288 -19029 1099 -18942
rect 288 -19112 312 -19029
rect 395 -19112 482 -19029
rect 565 -19112 652 -19029
rect 735 -19112 822 -19029
rect 905 -19112 992 -19029
rect 1075 -19112 1099 -19029
rect 27267 -18411 27290 -18323
rect 27377 -18411 27450 -18323
rect 27537 -18411 27610 -18323
rect 27697 -18411 27770 -18323
rect 27857 -18411 27930 -18323
rect 28017 -18411 28090 -18323
rect 28177 -18411 28195 -18323
rect 27267 -18483 28195 -18411
rect 27267 -18571 27290 -18483
rect 27377 -18571 27450 -18483
rect 27537 -18571 27610 -18483
rect 27697 -18571 27770 -18483
rect 27857 -18571 27930 -18483
rect 28017 -18571 28090 -18483
rect 28177 -18571 28195 -18483
rect 27267 -18643 28195 -18571
rect 27267 -18731 27290 -18643
rect 27377 -18731 27450 -18643
rect 27537 -18731 27610 -18643
rect 27697 -18731 27770 -18643
rect 27857 -18731 27930 -18643
rect 28017 -18731 28090 -18643
rect 28177 -18731 28195 -18643
rect 27267 -18803 28195 -18731
rect 27267 -18891 27290 -18803
rect 27377 -18891 27450 -18803
rect 27537 -18891 27610 -18803
rect 27697 -18891 27770 -18803
rect 27857 -18891 27930 -18803
rect 28017 -18891 28090 -18803
rect 28177 -18891 28195 -18803
rect 27267 -18963 28195 -18891
rect 27267 -19051 27290 -18963
rect 27377 -19051 27450 -18963
rect 27537 -19051 27610 -18963
rect 27697 -19051 27770 -18963
rect 27857 -19051 27930 -18963
rect 28017 -19051 28090 -18963
rect 28177 -19051 28195 -18963
rect 27267 -19073 28195 -19051
rect 288 -19135 1099 -19112
rect 27896 -19446 28694 -19411
rect 27896 -19447 28594 -19446
rect 27896 -19449 28260 -19447
rect 27896 -19537 27933 -19449
rect 28020 -19537 28113 -19449
rect 28200 -19535 28260 -19449
rect 28347 -19535 28440 -19447
rect 28527 -19534 28594 -19447
rect 28681 -19534 28694 -19446
rect 28527 -19535 28694 -19534
rect 28200 -19537 28694 -19535
rect 27896 -19569 28694 -19537
<< via2 >>
rect 1922 17502 2005 17585
rect 2092 17502 2175 17585
rect 2262 17502 2345 17585
rect 2432 17502 2515 17585
rect 2602 17502 2685 17585
rect 1922 17332 2005 17415
rect 2092 17332 2175 17415
rect 2262 17332 2345 17415
rect 2432 17332 2515 17415
rect 2602 17332 2685 17415
rect 1922 17162 2005 17245
rect 2092 17162 2175 17245
rect 2262 17162 2345 17245
rect 2432 17162 2515 17245
rect 2602 17162 2685 17245
rect 1922 16992 2005 17075
rect 2092 16992 2175 17075
rect 2262 16992 2345 17075
rect 2432 16992 2515 17075
rect 2602 16992 2685 17075
rect 1922 16822 2005 16905
rect 2092 16822 2175 16905
rect 2262 16822 2345 16905
rect 2432 16822 2515 16905
rect 2602 16822 2685 16905
rect 4065 17484 4148 17567
rect 4235 17484 4318 17567
rect 4405 17484 4488 17567
rect 4575 17484 4658 17567
rect 4745 17484 4828 17567
rect 4065 17314 4148 17397
rect 4235 17314 4318 17397
rect 4405 17314 4488 17397
rect 4575 17314 4658 17397
rect 4745 17314 4828 17397
rect 4065 17144 4148 17227
rect 4235 17144 4318 17227
rect 4405 17144 4488 17227
rect 4575 17144 4658 17227
rect 4745 17144 4828 17227
rect 4065 16974 4148 17057
rect 4235 16974 4318 17057
rect 4405 16974 4488 17057
rect 4575 16974 4658 17057
rect 4745 16974 4828 17057
rect 4065 16804 4148 16887
rect 4235 16804 4318 16887
rect 4405 16804 4488 16887
rect 4575 16804 4658 16887
rect 4745 16804 4828 16887
rect -597 15725 -541 15781
rect -493 15725 -437 15781
rect -389 15725 -333 15781
rect 18000 17202 18083 17285
rect 18170 17202 18253 17285
rect 18340 17202 18423 17285
rect 18510 17202 18593 17285
rect 18680 17202 18763 17285
rect 85647 17285 85730 17368
rect 85817 17285 85900 17368
rect 85987 17285 86070 17368
rect 86157 17285 86240 17368
rect 86327 17285 86410 17368
rect 18000 17032 18083 17115
rect 18170 17032 18253 17115
rect 18340 17032 18423 17115
rect 18510 17032 18593 17115
rect 18680 17032 18763 17115
rect 18000 16862 18083 16945
rect 18170 16862 18253 16945
rect 18340 16862 18423 16945
rect 18510 16862 18593 16945
rect 18680 16862 18763 16945
rect -4936 15575 -4853 15658
rect -4766 15575 -4683 15658
rect -4596 15575 -4513 15658
rect -4426 15575 -4343 15658
rect -4256 15575 -4173 15658
rect -597 15621 -541 15677
rect -493 15621 -437 15677
rect -389 15621 -333 15677
rect -597 15517 -541 15573
rect -493 15517 -437 15573
rect -389 15517 -333 15573
rect -4936 15405 -4853 15488
rect -4766 15405 -4683 15488
rect -4596 15405 -4513 15488
rect -4426 15405 -4343 15488
rect -4256 15405 -4173 15488
rect -4936 15235 -4853 15318
rect -4766 15235 -4683 15318
rect -4596 15235 -4513 15318
rect -4426 15235 -4343 15318
rect -4256 15235 -4173 15318
rect -3538 15248 -3482 15304
rect -3434 15248 -3378 15304
rect -3330 15248 -3274 15304
rect -4936 15065 -4853 15148
rect -4766 15065 -4683 15148
rect -4596 15065 -4513 15148
rect -4426 15065 -4343 15148
rect -4256 15065 -4173 15148
rect -3538 15144 -3482 15200
rect -3434 15144 -3378 15200
rect -3330 15144 -3274 15200
rect -3538 15040 -3482 15096
rect -3434 15040 -3378 15096
rect -3330 15040 -3274 15096
rect -161 15296 -105 15352
rect -57 15296 -1 15352
rect 47 15296 103 15352
rect 18000 16692 18083 16775
rect 18170 16692 18253 16775
rect 18340 16692 18423 16775
rect 18510 16692 18593 16775
rect 18680 16692 18763 16775
rect 18000 16522 18083 16605
rect 18170 16522 18253 16605
rect 18340 16522 18423 16605
rect 18510 16522 18593 16605
rect 18680 16522 18763 16605
rect 22004 17138 22087 17221
rect 22174 17138 22257 17221
rect 22344 17138 22427 17221
rect 22514 17138 22597 17221
rect 22684 17138 22767 17221
rect 22004 16968 22087 17051
rect 22174 16968 22257 17051
rect 22344 16968 22427 17051
rect 22514 16968 22597 17051
rect 22684 16968 22767 17051
rect 22004 16798 22087 16881
rect 22174 16798 22257 16881
rect 22344 16798 22427 16881
rect 22514 16798 22597 16881
rect 22684 16798 22767 16881
rect 22004 16628 22087 16711
rect 22174 16628 22257 16711
rect 22344 16628 22427 16711
rect 22514 16628 22597 16711
rect 22684 16628 22767 16711
rect 85647 17115 85730 17198
rect 85817 17115 85900 17198
rect 85987 17115 86070 17198
rect 86157 17115 86240 17198
rect 86327 17115 86410 17198
rect 85647 16945 85730 17028
rect 85817 16945 85900 17028
rect 85987 16945 86070 17028
rect 86157 16945 86240 17028
rect 86327 16945 86410 17028
rect 85647 16775 85730 16858
rect 85817 16775 85900 16858
rect 85987 16775 86070 16858
rect 86157 16775 86240 16858
rect 86327 16775 86410 16858
rect 85647 16605 85730 16688
rect 85817 16605 85900 16688
rect 85987 16605 86070 16688
rect 86157 16605 86240 16688
rect 86327 16605 86410 16688
rect 89264 17276 89347 17359
rect 89434 17276 89517 17359
rect 89604 17276 89687 17359
rect 89774 17276 89857 17359
rect 89944 17276 90027 17359
rect 89264 17106 89347 17189
rect 89434 17106 89517 17189
rect 89604 17106 89687 17189
rect 89774 17106 89857 17189
rect 89944 17106 90027 17189
rect 89264 16936 89347 17019
rect 89434 16936 89517 17019
rect 89604 16936 89687 17019
rect 89774 16936 89857 17019
rect 89944 16936 90027 17019
rect 89264 16766 89347 16849
rect 89434 16766 89517 16849
rect 89604 16766 89687 16849
rect 89774 16766 89857 16849
rect 89944 16766 90027 16849
rect 89264 16596 89347 16679
rect 89434 16596 89517 16679
rect 89604 16596 89687 16679
rect 89774 16596 89857 16679
rect 89944 16596 90027 16679
rect -161 15192 -105 15248
rect -57 15192 -1 15248
rect 47 15192 103 15248
rect -161 15088 -105 15144
rect -57 15088 -1 15144
rect 47 15088 103 15144
rect -4936 14895 -4853 14978
rect -4766 14895 -4683 14978
rect -4596 14895 -4513 14978
rect -4426 14895 -4343 14978
rect -4256 14895 -4173 14978
rect -2475 14673 -2419 14729
rect -2371 14673 -2315 14729
rect -2267 14673 -2211 14729
rect -2475 14569 -2419 14625
rect -2371 14569 -2315 14625
rect -2267 14569 -2211 14625
rect -2475 14465 -2419 14521
rect -2371 14465 -2315 14521
rect -2267 14465 -2211 14521
rect -3015 14272 -2959 14328
rect -2911 14272 -2855 14328
rect -2807 14272 -2751 14328
rect -3015 14168 -2959 14224
rect -2911 14168 -2855 14224
rect -2807 14168 -2751 14224
rect -3015 14064 -2959 14120
rect -2911 14064 -2855 14120
rect -2807 14064 -2751 14120
rect -1040 13863 -984 13919
rect -936 13863 -880 13919
rect -832 13863 -776 13919
rect -1040 13759 -984 13815
rect -936 13759 -880 13815
rect -832 13759 -776 13815
rect -1040 13655 -984 13711
rect -936 13655 -880 13711
rect -832 13655 -776 13711
rect -1444 13309 -1388 13365
rect -1340 13309 -1284 13365
rect -1236 13309 -1180 13365
rect -1444 13205 -1388 13261
rect -1340 13205 -1284 13261
rect -1236 13205 -1180 13261
rect -1444 13101 -1388 13157
rect -1340 13101 -1284 13157
rect -1236 13101 -1180 13157
rect -4953 12641 -4870 12724
rect -4783 12641 -4700 12724
rect -4613 12641 -4530 12724
rect -4443 12641 -4360 12724
rect -4273 12641 -4190 12724
rect -4953 12471 -4870 12554
rect -4783 12471 -4700 12554
rect -4613 12471 -4530 12554
rect -4443 12471 -4360 12554
rect -4273 12471 -4190 12554
rect -4953 12301 -4870 12384
rect -4783 12301 -4700 12384
rect -4613 12301 -4530 12384
rect -4443 12301 -4360 12384
rect -4273 12301 -4190 12384
rect -2992 12332 -2936 12388
rect -2888 12332 -2832 12388
rect -2784 12332 -2728 12388
rect -2992 12228 -2936 12284
rect -2888 12228 -2832 12284
rect -2784 12228 -2728 12284
rect -4953 12131 -4870 12214
rect -4783 12131 -4700 12214
rect -4613 12131 -4530 12214
rect -4443 12131 -4360 12214
rect -4273 12131 -4190 12214
rect -2992 12124 -2936 12180
rect -2888 12124 -2832 12180
rect -2784 12124 -2728 12180
rect -4953 11961 -4870 12044
rect -4783 11961 -4700 12044
rect -4613 11961 -4530 12044
rect -4443 11961 -4360 12044
rect -4273 11961 -4190 12044
rect -1957 11778 -1901 11834
rect -1853 11778 -1797 11834
rect -1749 11778 -1693 11834
rect 527 11783 583 11839
rect 631 11783 687 11839
rect 735 11783 791 11839
rect -1957 11674 -1901 11730
rect -1853 11674 -1797 11730
rect -1749 11674 -1693 11730
rect 527 11679 583 11735
rect 631 11679 687 11735
rect 735 11679 791 11735
rect -1957 11570 -1901 11626
rect -1853 11570 -1797 11626
rect -1749 11570 -1693 11626
rect 527 11575 583 11631
rect 631 11575 687 11631
rect 735 11575 791 11631
rect 15899 10558 15966 10624
rect 16529 10543 16596 10609
rect -4953 9269 -4870 9352
rect -4783 9269 -4700 9352
rect -4613 9269 -4530 9352
rect -4443 9269 -4360 9352
rect -4273 9269 -4190 9352
rect -4953 9099 -4870 9182
rect -4783 9099 -4700 9182
rect -4613 9099 -4530 9182
rect -4443 9099 -4360 9182
rect -4273 9099 -4190 9182
rect -2970 9027 -2914 9083
rect -2866 9027 -2810 9083
rect -2762 9027 -2706 9083
rect -4953 8929 -4870 9012
rect -4783 8929 -4700 9012
rect -4613 8929 -4530 9012
rect -4443 8929 -4360 9012
rect -4273 8929 -4190 9012
rect -2970 8923 -2914 8979
rect -2866 8923 -2810 8979
rect -2762 8923 -2706 8979
rect -4953 8759 -4870 8842
rect -4783 8759 -4700 8842
rect -4613 8759 -4530 8842
rect -4443 8759 -4360 8842
rect -4273 8759 -4190 8842
rect -2970 8819 -2914 8875
rect -2866 8819 -2810 8875
rect -2762 8819 -2706 8875
rect -4953 8589 -4870 8672
rect -4783 8589 -4700 8672
rect -4613 8589 -4530 8672
rect -4443 8589 -4360 8672
rect -4273 8589 -4190 8672
rect 15887 8222 15954 8288
rect 15890 7141 15957 7207
rect -5021 6959 -4938 7042
rect -4851 6959 -4768 7042
rect -4681 6959 -4598 7042
rect -4511 6959 -4428 7042
rect -4341 6959 -4258 7042
rect -5021 6789 -4938 6872
rect -4851 6789 -4768 6872
rect -4681 6789 -4598 6872
rect -4511 6789 -4428 6872
rect -4341 6789 -4258 6872
rect 614 6731 670 6787
rect 718 6731 774 6787
rect 822 6731 878 6787
rect -5021 6619 -4938 6702
rect -4851 6619 -4768 6702
rect -4681 6619 -4598 6702
rect -4511 6619 -4428 6702
rect -4341 6619 -4258 6702
rect 614 6627 670 6683
rect 718 6627 774 6683
rect 822 6627 878 6683
rect -5021 6449 -4938 6532
rect -4851 6449 -4768 6532
rect -4681 6449 -4598 6532
rect -4511 6449 -4428 6532
rect -4341 6449 -4258 6532
rect 614 6523 670 6579
rect 718 6523 774 6579
rect 822 6523 878 6579
rect -5021 6279 -4938 6362
rect -4851 6279 -4768 6362
rect -4681 6279 -4598 6362
rect -4511 6279 -4428 6362
rect -4341 6279 -4258 6362
rect -5004 5207 -4921 5290
rect -4834 5207 -4751 5290
rect -4664 5207 -4581 5290
rect -4494 5207 -4411 5290
rect -4324 5207 -4241 5290
rect -5004 5037 -4921 5120
rect -4834 5037 -4751 5120
rect -4664 5037 -4581 5120
rect -4494 5037 -4411 5120
rect -4324 5037 -4241 5120
rect -5004 4867 -4921 4950
rect -4834 4867 -4751 4950
rect -4664 4867 -4581 4950
rect -4494 4867 -4411 4950
rect -4324 4867 -4241 4950
rect -2470 4894 -2414 4950
rect -2366 4894 -2310 4950
rect -2262 4894 -2206 4950
rect -2470 4790 -2414 4846
rect -2366 4790 -2310 4846
rect -2262 4790 -2206 4846
rect -5004 4697 -4921 4780
rect -4834 4697 -4751 4780
rect -4664 4697 -4581 4780
rect -4494 4697 -4411 4780
rect -4324 4697 -4241 4780
rect -2470 4686 -2414 4742
rect -2366 4686 -2310 4742
rect -2262 4686 -2206 4742
rect -5004 4527 -4921 4610
rect -4834 4527 -4751 4610
rect -4664 4527 -4581 4610
rect -4494 4527 -4411 4610
rect -4324 4527 -4241 4610
rect -5155 2694 -5072 2777
rect -4985 2694 -4902 2777
rect -4815 2694 -4732 2777
rect -4645 2694 -4562 2777
rect -4475 2694 -4392 2777
rect -5155 2524 -5072 2607
rect -4985 2524 -4902 2607
rect -4815 2524 -4732 2607
rect -4645 2524 -4562 2607
rect -4475 2524 -4392 2607
rect -5155 2354 -5072 2437
rect -4985 2354 -4902 2437
rect -4815 2354 -4732 2437
rect -4645 2354 -4562 2437
rect -4475 2354 -4392 2437
rect -165 2396 -109 2452
rect -61 2396 -5 2452
rect 43 2396 99 2452
rect -165 2292 -109 2348
rect -61 2292 -5 2348
rect 43 2292 99 2348
rect -5155 2184 -5072 2267
rect -4985 2184 -4902 2267
rect -4815 2184 -4732 2267
rect -4645 2184 -4562 2267
rect -4475 2184 -4392 2267
rect -165 2188 -109 2244
rect -61 2188 -5 2244
rect 43 2188 99 2244
rect -5155 2014 -5072 2097
rect -4985 2014 -4902 2097
rect -4815 2014 -4732 2097
rect -4645 2014 -4562 2097
rect -4475 2014 -4392 2097
rect -2470 1000 -2414 1056
rect -2366 1000 -2310 1056
rect -2262 1000 -2206 1056
rect 665 983 721 1039
rect 769 983 825 1039
rect 873 983 929 1039
rect -2470 896 -2414 952
rect -2366 896 -2310 952
rect -2262 896 -2206 952
rect 665 879 721 935
rect 769 879 825 935
rect 873 879 929 935
rect -2470 792 -2414 848
rect -2366 792 -2310 848
rect -2262 792 -2206 848
rect 665 775 721 831
rect 769 775 825 831
rect 873 775 929 831
rect -5155 -1724 -5072 -1641
rect -4985 -1724 -4902 -1641
rect -4815 -1724 -4732 -1641
rect -4645 -1724 -4562 -1641
rect -4475 -1724 -4392 -1641
rect -5155 -1894 -5072 -1811
rect -4985 -1894 -4902 -1811
rect -4815 -1894 -4732 -1811
rect -4645 -1894 -4562 -1811
rect -4475 -1894 -4392 -1811
rect -1966 -1953 -1910 -1897
rect -1862 -1953 -1806 -1897
rect -1758 -1953 -1702 -1897
rect -5155 -2064 -5072 -1981
rect -4985 -2064 -4902 -1981
rect -4815 -2064 -4732 -1981
rect -4645 -2064 -4562 -1981
rect -4475 -2064 -4392 -1981
rect -1966 -2057 -1910 -2001
rect -1862 -2057 -1806 -2001
rect -1758 -2057 -1702 -2001
rect -5155 -2234 -5072 -2151
rect -4985 -2234 -4902 -2151
rect -4815 -2234 -4732 -2151
rect -4645 -2234 -4562 -2151
rect -4475 -2234 -4392 -2151
rect -1966 -2161 -1910 -2105
rect -1862 -2161 -1806 -2105
rect -1758 -2161 -1702 -2105
rect -5155 -2404 -5072 -2321
rect -4985 -2404 -4902 -2321
rect -4815 -2404 -4732 -2321
rect -4645 -2404 -4562 -2321
rect -4475 -2404 -4392 -2321
rect -152 -2318 -96 -2262
rect -48 -2318 8 -2262
rect 56 -2318 112 -2262
rect -152 -2422 -96 -2366
rect -48 -2422 8 -2366
rect 56 -2422 112 -2366
rect -152 -2526 -96 -2470
rect -48 -2526 8 -2470
rect 56 -2526 112 -2470
rect -3569 -2660 -3513 -2604
rect -3465 -2660 -3409 -2604
rect -3361 -2660 -3305 -2604
rect -3569 -2764 -3513 -2708
rect -3465 -2764 -3409 -2708
rect -3361 -2764 -3305 -2708
rect -3569 -2868 -3513 -2812
rect -3465 -2868 -3409 -2812
rect -3361 -2868 -3305 -2812
rect -57 -3003 -1 -2947
rect 47 -3003 103 -2947
rect 151 -3003 207 -2947
rect -1903 -3119 -1847 -3063
rect -1799 -3119 -1743 -3063
rect -1695 -3119 -1639 -3063
rect -1903 -3223 -1847 -3167
rect -1799 -3223 -1743 -3167
rect -1695 -3223 -1639 -3167
rect -1903 -3327 -1847 -3271
rect -1799 -3327 -1743 -3271
rect -1695 -3327 -1639 -3271
rect -57 -3107 -1 -3051
rect 47 -3107 103 -3051
rect 151 -3107 207 -3051
rect -57 -3211 -1 -3155
rect 47 -3211 103 -3155
rect 151 -3211 207 -3155
rect -5124 -4785 -5041 -4702
rect -4954 -4785 -4871 -4702
rect -4784 -4785 -4701 -4702
rect -4614 -4785 -4531 -4702
rect -4444 -4785 -4361 -4702
rect -5124 -4955 -5041 -4872
rect -4954 -4955 -4871 -4872
rect -4784 -4955 -4701 -4872
rect -4614 -4955 -4531 -4872
rect -4444 -4955 -4361 -4872
rect 731 -5032 787 -4976
rect 835 -5032 891 -4976
rect 939 -5032 995 -4976
rect -5124 -5125 -5041 -5042
rect -4954 -5125 -4871 -5042
rect -4784 -5125 -4701 -5042
rect -4614 -5125 -4531 -5042
rect -4444 -5125 -4361 -5042
rect 731 -5136 787 -5080
rect 835 -5136 891 -5080
rect 939 -5136 995 -5080
rect -5124 -5295 -5041 -5212
rect -4954 -5295 -4871 -5212
rect -4784 -5295 -4701 -5212
rect -4614 -5295 -4531 -5212
rect -4444 -5295 -4361 -5212
rect 731 -5240 787 -5184
rect 835 -5240 891 -5184
rect 939 -5240 995 -5184
rect -5124 -5465 -5041 -5382
rect -4954 -5465 -4871 -5382
rect -4784 -5465 -4701 -5382
rect -4614 -5465 -4531 -5382
rect -4444 -5465 -4361 -5382
rect 16041 -6208 16108 -6142
rect 16538 -6208 16605 -6142
rect -5099 -7654 -5016 -7571
rect -4929 -7654 -4846 -7571
rect -4759 -7654 -4676 -7571
rect -4589 -7654 -4506 -7571
rect -4419 -7654 -4336 -7571
rect -5099 -7824 -5016 -7741
rect -4929 -7824 -4846 -7741
rect -4759 -7824 -4676 -7741
rect -4589 -7824 -4506 -7741
rect -4419 -7824 -4336 -7741
rect -5099 -7994 -5016 -7911
rect -4929 -7994 -4846 -7911
rect -4759 -7994 -4676 -7911
rect -4589 -7994 -4506 -7911
rect -4419 -7994 -4336 -7911
rect -2493 -7932 -2437 -7876
rect -2389 -7932 -2333 -7876
rect -2285 -7932 -2229 -7876
rect -2493 -8036 -2437 -7980
rect -2389 -8036 -2333 -7980
rect -2285 -8036 -2229 -7980
rect -5099 -8164 -5016 -8081
rect -4929 -8164 -4846 -8081
rect -4759 -8164 -4676 -8081
rect -4589 -8164 -4506 -8081
rect -4419 -8164 -4336 -8081
rect -2493 -8140 -2437 -8084
rect -2389 -8140 -2333 -8084
rect -2285 -8140 -2229 -8084
rect -5099 -8334 -5016 -8251
rect -4929 -8334 -4846 -8251
rect -4759 -8334 -4676 -8251
rect -4589 -8334 -4506 -8251
rect -4419 -8334 -4336 -8251
rect -611 -8310 -555 -8254
rect -507 -8310 -451 -8254
rect -403 -8310 -347 -8254
rect -611 -8414 -555 -8358
rect -507 -8414 -451 -8358
rect -403 -8414 -347 -8358
rect 713 -8368 769 -8312
rect 817 -8368 873 -8312
rect 921 -8368 977 -8312
rect -611 -8518 -555 -8462
rect -507 -8518 -451 -8462
rect -403 -8518 -347 -8462
rect 713 -8472 769 -8416
rect 817 -8472 873 -8416
rect 921 -8472 977 -8416
rect 713 -8576 769 -8520
rect 817 -8576 873 -8520
rect 921 -8576 977 -8520
rect 16045 -8550 16112 -8484
rect -2983 -9138 -2927 -9082
rect -2879 -9138 -2823 -9082
rect -2775 -9138 -2719 -9082
rect 789 -9129 845 -9073
rect 893 -9129 949 -9073
rect 997 -9129 1053 -9073
rect -2983 -9242 -2927 -9186
rect -2879 -9242 -2823 -9186
rect -2775 -9242 -2719 -9186
rect 789 -9233 845 -9177
rect 893 -9233 949 -9177
rect 997 -9233 1053 -9177
rect -2983 -9346 -2927 -9290
rect -2879 -9346 -2823 -9290
rect -2775 -9346 -2719 -9290
rect 789 -9337 845 -9281
rect 893 -9337 949 -9281
rect 997 -9337 1053 -9281
rect 16058 -9628 16125 -9562
rect -5076 -9758 -4993 -9675
rect -4906 -9758 -4823 -9675
rect -4736 -9758 -4653 -9675
rect -4566 -9758 -4483 -9675
rect -4396 -9758 -4313 -9675
rect -5076 -9928 -4993 -9845
rect -4906 -9928 -4823 -9845
rect -4736 -9928 -4653 -9845
rect -4566 -9928 -4483 -9845
rect -4396 -9928 -4313 -9845
rect -5076 -10098 -4993 -10015
rect -4906 -10098 -4823 -10015
rect -4736 -10098 -4653 -10015
rect -4566 -10098 -4483 -10015
rect -4396 -10098 -4313 -10015
rect -5076 -10268 -4993 -10185
rect -4906 -10268 -4823 -10185
rect -4736 -10268 -4653 -10185
rect -4566 -10268 -4483 -10185
rect -4396 -10268 -4313 -10185
rect -5076 -10438 -4993 -10355
rect -4906 -10438 -4823 -10355
rect -4736 -10438 -4653 -10355
rect -4566 -10438 -4483 -10355
rect -4396 -10438 -4313 -10355
rect 1154 -10791 1210 -10735
rect 1258 -10791 1314 -10735
rect 1362 -10791 1418 -10735
rect 1154 -10895 1210 -10839
rect 1258 -10895 1314 -10839
rect 1362 -10895 1418 -10839
rect 1154 -10999 1210 -10943
rect 1258 -10999 1314 -10943
rect 1362 -10999 1418 -10943
rect -5053 -11932 -4970 -11849
rect -4883 -11932 -4800 -11849
rect -4713 -11932 -4630 -11849
rect -4543 -11932 -4460 -11849
rect -4373 -11932 -4290 -11849
rect -5053 -12102 -4970 -12019
rect -4883 -12102 -4800 -12019
rect -4713 -12102 -4630 -12019
rect -4543 -12102 -4460 -12019
rect -4373 -12102 -4290 -12019
rect -5053 -12272 -4970 -12189
rect -4883 -12272 -4800 -12189
rect -4713 -12272 -4630 -12189
rect -4543 -12272 -4460 -12189
rect -4373 -12272 -4290 -12189
rect -1925 -12200 -1869 -12144
rect -1821 -12200 -1765 -12144
rect -1717 -12200 -1661 -12144
rect -1925 -12304 -1869 -12248
rect -1821 -12304 -1765 -12248
rect -1717 -12304 -1661 -12248
rect -5053 -12442 -4970 -12359
rect -4883 -12442 -4800 -12359
rect -4713 -12442 -4630 -12359
rect -4543 -12442 -4460 -12359
rect -4373 -12442 -4290 -12359
rect -1925 -12408 -1869 -12352
rect -1821 -12408 -1765 -12352
rect -1717 -12408 -1661 -12352
rect -5053 -12612 -4970 -12529
rect -4883 -12612 -4800 -12529
rect -4713 -12612 -4630 -12529
rect -4543 -12612 -4460 -12529
rect -4373 -12612 -4290 -12529
rect -5099 -13736 -5016 -13653
rect -4929 -13736 -4846 -13653
rect -4759 -13736 -4676 -13653
rect -4589 -13736 -4506 -13653
rect -4419 -13736 -4336 -13653
rect -5099 -13906 -5016 -13823
rect -4929 -13906 -4846 -13823
rect -4759 -13906 -4676 -13823
rect -4589 -13906 -4506 -13823
rect -4419 -13906 -4336 -13823
rect -5099 -14076 -5016 -13993
rect -4929 -14076 -4846 -13993
rect -4759 -14076 -4676 -13993
rect -4589 -14076 -4506 -13993
rect -4419 -14076 -4336 -13993
rect -1471 -14005 -1415 -13949
rect -1367 -14005 -1311 -13949
rect -1263 -14005 -1207 -13949
rect -1471 -14109 -1415 -14053
rect -1367 -14109 -1311 -14053
rect -1263 -14109 -1207 -14053
rect -5099 -14246 -5016 -14163
rect -4929 -14246 -4846 -14163
rect -4759 -14246 -4676 -14163
rect -4589 -14246 -4506 -14163
rect -4419 -14246 -4336 -14163
rect -1471 -14213 -1415 -14157
rect -1367 -14213 -1311 -14157
rect -1263 -14213 -1207 -14157
rect -5099 -14416 -5016 -14333
rect -4929 -14416 -4846 -14333
rect -4759 -14416 -4676 -14333
rect -4589 -14416 -4506 -14333
rect -4419 -14416 -4336 -14333
rect -5053 -15508 -4970 -15425
rect -4883 -15508 -4800 -15425
rect -4713 -15508 -4630 -15425
rect -4543 -15508 -4460 -15425
rect -4373 -15508 -4290 -15425
rect -5053 -15678 -4970 -15595
rect -4883 -15678 -4800 -15595
rect -4713 -15678 -4630 -15595
rect -4543 -15678 -4460 -15595
rect -4373 -15678 -4290 -15595
rect -5053 -15848 -4970 -15765
rect -4883 -15848 -4800 -15765
rect -4713 -15848 -4630 -15765
rect -4543 -15848 -4460 -15765
rect -4373 -15848 -4290 -15765
rect -66 -15774 -10 -15718
rect 38 -15774 94 -15718
rect 142 -15774 198 -15718
rect -66 -15878 -10 -15822
rect 38 -15878 94 -15822
rect 142 -15878 198 -15822
rect -5053 -16018 -4970 -15935
rect -4883 -16018 -4800 -15935
rect -4713 -16018 -4630 -15935
rect -4543 -16018 -4460 -15935
rect -4373 -16018 -4290 -15935
rect -66 -15982 -10 -15926
rect 38 -15982 94 -15926
rect 142 -15982 198 -15926
rect -5053 -16188 -4970 -16105
rect -4883 -16188 -4800 -16105
rect -4713 -16188 -4630 -16105
rect -4543 -16188 -4460 -16105
rect -4373 -16188 -4290 -16105
rect 17047 8213 17114 8279
rect 17013 -8550 17080 -8484
rect 17599 7141 17666 7207
rect 22004 16458 22087 16541
rect 22174 16458 22257 16541
rect 22344 16458 22427 16541
rect 22514 16458 22597 16541
rect 22684 16458 22767 16541
rect 49191 16221 49274 16304
rect 49361 16221 49444 16304
rect 49531 16221 49614 16304
rect 49701 16221 49784 16304
rect 49871 16221 49954 16304
rect 49191 16051 49274 16134
rect 49361 16051 49444 16134
rect 49531 16051 49614 16134
rect 49701 16051 49784 16134
rect 49871 16051 49954 16134
rect 49191 15881 49274 15964
rect 49361 15881 49444 15964
rect 49531 15881 49614 15964
rect 49701 15881 49784 15964
rect 49871 15881 49954 15964
rect 49191 15711 49274 15794
rect 49361 15711 49444 15794
rect 49531 15711 49614 15794
rect 49701 15711 49784 15794
rect 49871 15711 49954 15794
rect 49191 15541 49274 15624
rect 49361 15541 49444 15624
rect 49531 15541 49614 15624
rect 49701 15541 49784 15624
rect 49871 15541 49954 15624
rect 52345 16249 52428 16332
rect 52515 16249 52598 16332
rect 52685 16249 52768 16332
rect 52855 16249 52938 16332
rect 53025 16249 53108 16332
rect 52345 16079 52428 16162
rect 52515 16079 52598 16162
rect 52685 16079 52768 16162
rect 52855 16079 52938 16162
rect 53025 16079 53108 16162
rect 52345 15909 52428 15992
rect 52515 15909 52598 15992
rect 52685 15909 52768 15992
rect 52855 15909 52938 15992
rect 53025 15909 53108 15992
rect 52345 15739 52428 15822
rect 52515 15739 52598 15822
rect 52685 15739 52768 15822
rect 52855 15739 52938 15822
rect 53025 15739 53108 15822
rect 52345 15569 52428 15652
rect 52515 15569 52598 15652
rect 52685 15569 52768 15652
rect 52855 15569 52938 15652
rect 53025 15569 53108 15652
rect 154968 17080 155051 17163
rect 155138 17080 155221 17163
rect 155308 17080 155391 17163
rect 155478 17080 155561 17163
rect 155648 17080 155731 17163
rect 154968 16910 155051 16993
rect 155138 16910 155221 16993
rect 155308 16910 155391 16993
rect 155478 16910 155561 16993
rect 155648 16910 155731 16993
rect 154968 16740 155051 16823
rect 155138 16740 155221 16823
rect 155308 16740 155391 16823
rect 155478 16740 155561 16823
rect 155648 16740 155731 16823
rect 154968 16570 155051 16653
rect 155138 16570 155221 16653
rect 155308 16570 155391 16653
rect 155478 16570 155561 16653
rect 155648 16570 155731 16653
rect 154968 16400 155051 16483
rect 155138 16400 155221 16483
rect 155308 16400 155391 16483
rect 155478 16400 155561 16483
rect 155648 16400 155731 16483
rect 157343 17080 157426 17163
rect 157513 17080 157596 17163
rect 157683 17080 157766 17163
rect 157853 17080 157936 17163
rect 158023 17080 158106 17163
rect 157343 16910 157426 16993
rect 157513 16910 157596 16993
rect 157683 16910 157766 16993
rect 157853 16910 157936 16993
rect 158023 16910 158106 16993
rect 157343 16740 157426 16823
rect 157513 16740 157596 16823
rect 157683 16740 157766 16823
rect 157853 16740 157936 16823
rect 158023 16740 158106 16823
rect 157343 16570 157426 16653
rect 157513 16570 157596 16653
rect 157683 16570 157766 16653
rect 157853 16570 157936 16653
rect 158023 16570 158106 16653
rect 157343 16400 157426 16483
rect 157513 16400 157596 16483
rect 157683 16400 157766 16483
rect 157853 16400 157936 16483
rect 158023 16400 158106 16483
rect 133349 14349 133436 14437
rect 133529 14349 133616 14437
rect 133676 14351 133763 14439
rect 133856 14351 133943 14439
rect 134010 14352 134097 14440
rect 133349 14169 133436 14257
rect 133529 14169 133616 14257
rect 133676 14171 133763 14259
rect 133856 14171 133943 14259
rect 134010 14172 134097 14260
rect 133331 13956 133418 14044
rect 133511 13956 133598 14044
rect 133658 13958 133745 14046
rect 133838 13958 133925 14046
rect 133992 13959 134079 14047
rect 133331 13776 133418 13864
rect 133511 13776 133598 13864
rect 133658 13778 133745 13866
rect 133838 13778 133925 13866
rect 133992 13779 134079 13867
rect 135855 14333 135942 14421
rect 136035 14333 136122 14421
rect 136182 14335 136269 14423
rect 136362 14335 136449 14423
rect 136516 14336 136603 14424
rect 135855 14153 135942 14241
rect 136035 14153 136122 14241
rect 136182 14155 136269 14243
rect 136362 14155 136449 14243
rect 136516 14156 136603 14244
rect 135837 13940 135924 14028
rect 136017 13940 136104 14028
rect 136164 13942 136251 14030
rect 136344 13942 136431 14030
rect 136498 13943 136585 14031
rect 135837 13760 135924 13848
rect 136017 13760 136104 13848
rect 136164 13762 136251 13850
rect 136344 13762 136431 13850
rect 136498 13763 136585 13851
rect 138571 14352 138658 14440
rect 138751 14352 138838 14440
rect 138898 14354 138985 14442
rect 139078 14354 139165 14442
rect 139232 14355 139319 14443
rect 138571 14172 138658 14260
rect 138751 14172 138838 14260
rect 138898 14174 138985 14262
rect 139078 14174 139165 14262
rect 139232 14175 139319 14263
rect 138553 13959 138640 14047
rect 138733 13959 138820 14047
rect 138880 13961 138967 14049
rect 139060 13961 139147 14049
rect 139214 13962 139301 14050
rect 138553 13779 138640 13867
rect 138733 13779 138820 13867
rect 138880 13781 138967 13869
rect 139060 13781 139147 13869
rect 139214 13782 139301 13870
rect 23348 12787 23435 12875
rect 23528 12787 23615 12875
rect 23348 12607 23435 12695
rect 23528 12607 23615 12695
rect 18836 9210 18919 9293
rect 19006 9210 19089 9293
rect 19176 9210 19259 9293
rect 18836 9040 18919 9123
rect 19006 9040 19089 9123
rect 19176 9040 19259 9123
rect 18836 8870 18919 8953
rect 19006 8870 19089 8953
rect 19176 8870 19259 8953
rect 18838 8631 18921 8714
rect 19008 8631 19091 8714
rect 19178 8631 19261 8714
rect 18838 8461 18921 8544
rect 19008 8461 19091 8544
rect 19178 8461 19261 8544
rect 18838 8291 18921 8374
rect 19008 8291 19091 8374
rect 19178 8291 19261 8374
rect 150342 6580 150429 6668
rect 150522 6580 150609 6668
rect 150669 6582 150756 6670
rect 150849 6582 150936 6670
rect 151003 6583 151090 6671
rect 150342 6400 150429 6488
rect 150522 6400 150609 6488
rect 150669 6402 150756 6490
rect 150849 6402 150936 6490
rect 151003 6403 151090 6491
rect 75648 5906 75735 5994
rect 75828 5906 75915 5994
rect 75975 5908 76062 5996
rect 76155 5908 76242 5996
rect 76309 5909 76396 5997
rect 76449 5908 76536 5996
rect 76590 5906 76677 5994
rect 75648 5726 75735 5814
rect 75828 5726 75915 5814
rect 75975 5728 76062 5816
rect 76155 5728 76242 5816
rect 76309 5729 76396 5817
rect 76449 5728 76536 5816
rect 76590 5726 76677 5814
rect 80919 5941 81006 6029
rect 81099 5941 81186 6029
rect 81246 5943 81333 6031
rect 81426 5943 81513 6031
rect 81580 5944 81667 6032
rect 81734 5945 81821 6033
rect 81882 5943 81969 6031
rect 80919 5761 81006 5849
rect 81099 5761 81186 5849
rect 81246 5763 81333 5851
rect 81426 5763 81513 5851
rect 81580 5764 81667 5852
rect 81734 5765 81821 5853
rect 81882 5763 81969 5851
rect 126226 4814 126313 4902
rect 126406 4814 126493 4902
rect 126226 4634 126313 4722
rect 126406 4634 126493 4722
rect 56847 4129 56934 4217
rect 57027 4129 57114 4217
rect 56847 3949 56934 4037
rect 57027 3949 57114 4037
rect 113837 3774 113924 3862
rect 114017 3774 114104 3862
rect 113837 3594 113924 3682
rect 114017 3594 114104 3682
rect 113839 3433 113926 3521
rect 114019 3433 114106 3521
rect 113839 3253 113926 3341
rect 114019 3253 114106 3341
rect 114475 3824 114562 3912
rect 114655 3824 114742 3912
rect 114475 3644 114562 3732
rect 114655 3644 114742 3732
rect 114473 3481 114560 3569
rect 114653 3481 114740 3569
rect 114473 3301 114560 3389
rect 114653 3301 114740 3389
rect 115082 3870 115169 3958
rect 115262 3870 115349 3958
rect 115082 3690 115169 3778
rect 115262 3690 115349 3778
rect 115082 3530 115169 3618
rect 115262 3530 115349 3618
rect 115082 3350 115169 3438
rect 115262 3350 115349 3438
rect 115729 3852 115816 3940
rect 115909 3852 115996 3940
rect 115729 3672 115816 3760
rect 115909 3672 115996 3760
rect 115732 3521 115819 3609
rect 115912 3521 115999 3609
rect 115732 3341 115819 3429
rect 115912 3341 115999 3429
rect 28075 589 28162 677
rect 28255 589 28342 677
rect 28402 591 28489 679
rect 28582 591 28669 679
rect 28736 592 28823 680
rect 28075 409 28162 497
rect 28255 409 28342 497
rect 28402 411 28489 499
rect 28582 411 28669 499
rect 28736 412 28823 500
rect 28057 196 28144 284
rect 28237 196 28324 284
rect 28384 198 28471 286
rect 28564 198 28651 286
rect 28718 199 28805 287
rect 28057 16 28144 104
rect 28237 16 28324 104
rect 28384 18 28471 106
rect 28564 18 28651 106
rect 28718 19 28805 107
rect 29881 636 29968 724
rect 30061 636 30148 724
rect 30208 638 30295 726
rect 30388 638 30475 726
rect 30542 639 30629 727
rect 29881 456 29968 544
rect 30061 456 30148 544
rect 30208 458 30295 546
rect 30388 458 30475 546
rect 30542 459 30629 547
rect 29887 248 29974 336
rect 30067 248 30154 336
rect 30214 250 30301 338
rect 30394 250 30481 338
rect 30548 251 30635 339
rect 29887 68 29974 156
rect 30067 68 30154 156
rect 30214 70 30301 158
rect 30394 70 30481 158
rect 30548 71 30635 159
rect 31618 636 31705 724
rect 31798 636 31885 724
rect 31945 638 32032 726
rect 32125 638 32212 726
rect 32279 639 32366 727
rect 48410 699 48475 764
rect 48535 699 48600 764
rect 48660 699 48725 764
rect 31618 456 31705 544
rect 31798 456 31885 544
rect 31945 458 32032 546
rect 32125 458 32212 546
rect 32279 459 32366 547
rect 31630 248 31717 336
rect 31810 248 31897 336
rect 31957 250 32044 338
rect 32137 250 32224 338
rect 32291 251 32378 339
rect 31630 68 31717 156
rect 31810 68 31897 156
rect 31957 70 32044 158
rect 32137 70 32224 158
rect 32291 71 32378 159
rect 64643 -1336 64699 -1280
rect 64747 -1336 64803 -1280
rect 64643 -1440 64699 -1384
rect 64747 -1440 64803 -1384
rect 64645 -1570 64701 -1514
rect 64749 -1570 64805 -1514
rect 64645 -1674 64701 -1618
rect 64749 -1674 64805 -1618
rect 23089 -2157 23176 -2069
rect 23269 -2157 23356 -2069
rect 23089 -2337 23176 -2249
rect 23269 -2337 23356 -2249
rect 86691 -2219 86778 -2131
rect 86871 -2219 86958 -2131
rect 87037 -2219 87124 -2131
rect 87217 -2219 87304 -2131
rect 87390 -2222 87477 -2134
rect 87570 -2222 87657 -2134
rect 86691 -2399 86778 -2311
rect 86871 -2399 86958 -2311
rect 87037 -2399 87124 -2311
rect 87217 -2399 87304 -2311
rect 87390 -2402 87477 -2314
rect 87570 -2402 87657 -2314
rect 85749 -3370 85836 -3282
rect 85929 -3370 86016 -3282
rect 86095 -3370 86182 -3282
rect 86275 -3370 86362 -3282
rect 86448 -3373 86535 -3285
rect 86628 -3373 86715 -3285
rect 85749 -3550 85836 -3462
rect 85929 -3550 86016 -3462
rect 86095 -3550 86182 -3462
rect 86275 -3550 86362 -3462
rect 86448 -3553 86535 -3465
rect 86628 -3553 86715 -3465
rect 18142 -5893 18225 -5810
rect 18312 -5893 18395 -5810
rect 18482 -5893 18565 -5810
rect 18142 -6063 18225 -5980
rect 18312 -6063 18395 -5980
rect 18482 -6063 18565 -5980
rect 18142 -6233 18225 -6150
rect 18312 -6233 18395 -6150
rect 18482 -6233 18565 -6150
rect 18151 -6475 18234 -6392
rect 18321 -6475 18404 -6392
rect 18491 -6475 18574 -6392
rect 18151 -6645 18234 -6562
rect 18321 -6645 18404 -6562
rect 18491 -6645 18574 -6562
rect 18151 -6815 18234 -6732
rect 18321 -6815 18404 -6732
rect 18491 -6815 18574 -6732
rect 17557 -9628 17624 -9562
rect 127458 268 127514 270
rect 127143 266 127199 268
rect 127143 214 127145 266
rect 127145 214 127197 266
rect 127197 214 127199 266
rect 127143 212 127199 214
rect 127247 266 127303 268
rect 127247 214 127249 266
rect 127249 214 127301 266
rect 127301 214 127303 266
rect 127247 212 127303 214
rect 127351 266 127407 268
rect 127351 214 127353 266
rect 127353 214 127405 266
rect 127405 214 127407 266
rect 127458 216 127460 268
rect 127460 216 127512 268
rect 127512 216 127514 268
rect 127458 214 127514 216
rect 127562 268 127618 270
rect 127562 216 127564 268
rect 127564 216 127616 268
rect 127616 216 127618 268
rect 127562 214 127618 216
rect 127666 268 127722 270
rect 127666 216 127668 268
rect 127668 216 127720 268
rect 127720 216 127722 268
rect 127666 214 127722 216
rect 127773 268 127829 270
rect 127773 216 127775 268
rect 127775 216 127827 268
rect 127827 216 127829 268
rect 127773 214 127829 216
rect 127877 268 127933 270
rect 127877 216 127879 268
rect 127879 216 127931 268
rect 127931 216 127933 268
rect 127877 214 127933 216
rect 127981 268 128037 270
rect 127981 216 127983 268
rect 127983 216 128035 268
rect 128035 216 128037 268
rect 127981 214 128037 216
rect 127351 212 127407 214
rect 127458 164 127514 166
rect 127143 162 127199 164
rect 127143 110 127145 162
rect 127145 110 127197 162
rect 127197 110 127199 162
rect 127143 108 127199 110
rect 127247 162 127303 164
rect 127247 110 127249 162
rect 127249 110 127301 162
rect 127301 110 127303 162
rect 127247 108 127303 110
rect 127351 162 127407 164
rect 127351 110 127353 162
rect 127353 110 127405 162
rect 127405 110 127407 162
rect 127458 112 127460 164
rect 127460 112 127512 164
rect 127512 112 127514 164
rect 127458 110 127514 112
rect 127562 164 127618 166
rect 127562 112 127564 164
rect 127564 112 127616 164
rect 127616 112 127618 164
rect 127562 110 127618 112
rect 127666 164 127722 166
rect 127666 112 127668 164
rect 127668 112 127720 164
rect 127720 112 127722 164
rect 127666 110 127722 112
rect 127773 164 127829 166
rect 127773 112 127775 164
rect 127775 112 127827 164
rect 127827 112 127829 164
rect 127773 110 127829 112
rect 127877 164 127933 166
rect 127877 112 127879 164
rect 127879 112 127931 164
rect 127931 112 127933 164
rect 127877 110 127933 112
rect 127981 164 128037 166
rect 127981 112 127983 164
rect 127983 112 128035 164
rect 128035 112 128037 164
rect 127981 110 128037 112
rect 127351 108 127407 110
rect 127458 60 127514 62
rect 127143 58 127199 60
rect 127143 6 127145 58
rect 127145 6 127197 58
rect 127197 6 127199 58
rect 127143 4 127199 6
rect 127247 58 127303 60
rect 127247 6 127249 58
rect 127249 6 127301 58
rect 127301 6 127303 58
rect 127247 4 127303 6
rect 127351 58 127407 60
rect 127351 6 127353 58
rect 127353 6 127405 58
rect 127405 6 127407 58
rect 127458 8 127460 60
rect 127460 8 127512 60
rect 127512 8 127514 60
rect 127458 6 127514 8
rect 127562 60 127618 62
rect 127562 8 127564 60
rect 127564 8 127616 60
rect 127616 8 127618 60
rect 127562 6 127618 8
rect 127666 60 127722 62
rect 127666 8 127668 60
rect 127668 8 127720 60
rect 127720 8 127722 60
rect 127666 6 127722 8
rect 127773 60 127829 62
rect 127773 8 127775 60
rect 127775 8 127827 60
rect 127827 8 127829 60
rect 127773 6 127829 8
rect 127877 60 127933 62
rect 127877 8 127879 60
rect 127879 8 127931 60
rect 127931 8 127933 60
rect 127877 6 127933 8
rect 127981 60 128037 62
rect 127981 8 127983 60
rect 127983 8 128035 60
rect 128035 8 128037 60
rect 127981 6 128037 8
rect 127351 4 127407 6
rect 116290 -125 116346 -123
rect 115975 -127 116031 -125
rect 115975 -179 115977 -127
rect 115977 -179 116029 -127
rect 116029 -179 116031 -127
rect 115975 -181 116031 -179
rect 116079 -127 116135 -125
rect 116079 -179 116081 -127
rect 116081 -179 116133 -127
rect 116133 -179 116135 -127
rect 116079 -181 116135 -179
rect 116183 -127 116239 -125
rect 116183 -179 116185 -127
rect 116185 -179 116237 -127
rect 116237 -179 116239 -127
rect 116290 -177 116292 -125
rect 116292 -177 116344 -125
rect 116344 -177 116346 -125
rect 116290 -179 116346 -177
rect 116394 -125 116450 -123
rect 116394 -177 116396 -125
rect 116396 -177 116448 -125
rect 116448 -177 116450 -125
rect 116394 -179 116450 -177
rect 116498 -125 116554 -123
rect 116498 -177 116500 -125
rect 116500 -177 116552 -125
rect 116552 -177 116554 -125
rect 116498 -179 116554 -177
rect 116605 -125 116661 -123
rect 116605 -177 116607 -125
rect 116607 -177 116659 -125
rect 116659 -177 116661 -125
rect 116605 -179 116661 -177
rect 116709 -125 116765 -123
rect 116709 -177 116711 -125
rect 116711 -177 116763 -125
rect 116763 -177 116765 -125
rect 116709 -179 116765 -177
rect 116813 -125 116869 -123
rect 116813 -177 116815 -125
rect 116815 -177 116867 -125
rect 116867 -177 116869 -125
rect 116813 -179 116869 -177
rect 116183 -181 116239 -179
rect 116290 -229 116346 -227
rect 115975 -231 116031 -229
rect 115975 -283 115977 -231
rect 115977 -283 116029 -231
rect 116029 -283 116031 -231
rect 115975 -285 116031 -283
rect 116079 -231 116135 -229
rect 116079 -283 116081 -231
rect 116081 -283 116133 -231
rect 116133 -283 116135 -231
rect 116079 -285 116135 -283
rect 116183 -231 116239 -229
rect 116183 -283 116185 -231
rect 116185 -283 116237 -231
rect 116237 -283 116239 -231
rect 116290 -281 116292 -229
rect 116292 -281 116344 -229
rect 116344 -281 116346 -229
rect 116290 -283 116346 -281
rect 116394 -229 116450 -227
rect 116394 -281 116396 -229
rect 116396 -281 116448 -229
rect 116448 -281 116450 -229
rect 116394 -283 116450 -281
rect 116498 -229 116554 -227
rect 116498 -281 116500 -229
rect 116500 -281 116552 -229
rect 116552 -281 116554 -229
rect 116498 -283 116554 -281
rect 116605 -229 116661 -227
rect 116605 -281 116607 -229
rect 116607 -281 116659 -229
rect 116659 -281 116661 -229
rect 116605 -283 116661 -281
rect 116709 -229 116765 -227
rect 116709 -281 116711 -229
rect 116711 -281 116763 -229
rect 116763 -281 116765 -229
rect 116709 -283 116765 -281
rect 116813 -229 116869 -227
rect 116813 -281 116815 -229
rect 116815 -281 116867 -229
rect 116867 -281 116869 -229
rect 116813 -283 116869 -281
rect 116183 -285 116239 -283
rect 116290 -333 116346 -331
rect 115975 -335 116031 -333
rect 115975 -387 115977 -335
rect 115977 -387 116029 -335
rect 116029 -387 116031 -335
rect 115975 -389 116031 -387
rect 116079 -335 116135 -333
rect 116079 -387 116081 -335
rect 116081 -387 116133 -335
rect 116133 -387 116135 -335
rect 116079 -389 116135 -387
rect 116183 -335 116239 -333
rect 116183 -387 116185 -335
rect 116185 -387 116237 -335
rect 116237 -387 116239 -335
rect 116290 -385 116292 -333
rect 116292 -385 116344 -333
rect 116344 -385 116346 -333
rect 116290 -387 116346 -385
rect 116394 -333 116450 -331
rect 116394 -385 116396 -333
rect 116396 -385 116448 -333
rect 116448 -385 116450 -333
rect 116394 -387 116450 -385
rect 116498 -333 116554 -331
rect 116498 -385 116500 -333
rect 116500 -385 116552 -333
rect 116552 -385 116554 -333
rect 116498 -387 116554 -385
rect 116605 -333 116661 -331
rect 116605 -385 116607 -333
rect 116607 -385 116659 -333
rect 116659 -385 116661 -333
rect 116605 -387 116661 -385
rect 116709 -333 116765 -331
rect 116709 -385 116711 -333
rect 116711 -385 116763 -333
rect 116763 -385 116765 -333
rect 116709 -387 116765 -385
rect 116813 -333 116869 -331
rect 116813 -385 116815 -333
rect 116815 -385 116867 -333
rect 116867 -385 116869 -333
rect 116813 -387 116869 -385
rect 116183 -389 116239 -387
rect 133929 -644 133985 -588
rect 134033 -644 134089 -588
rect 134165 -647 134221 -591
rect 134269 -647 134325 -591
rect 133929 -748 133985 -692
rect 134033 -748 134089 -692
rect 134165 -751 134221 -695
rect 134269 -751 134325 -695
rect 122342 -3307 122406 -3240
rect 122474 -3312 122538 -3245
rect 122347 -3432 122411 -3365
rect 122472 -3431 122536 -3364
rect 121036 -3946 121102 -3880
rect 121167 -3943 121233 -3877
rect 121035 -4075 121101 -4009
rect 121169 -4075 121235 -4009
rect 121032 -4203 121098 -4137
rect 121167 -4203 121233 -4137
rect 121627 -7169 121714 -7081
rect 121807 -7169 121894 -7081
rect 121973 -7169 122060 -7081
rect 122153 -7169 122240 -7081
rect 122326 -7172 122413 -7084
rect 122506 -7172 122593 -7084
rect 121627 -7349 121714 -7261
rect 121807 -7349 121894 -7261
rect 121973 -7349 122060 -7261
rect 122153 -7349 122240 -7261
rect 122326 -7352 122413 -7264
rect 122506 -7352 122593 -7264
rect 170292 -7173 170379 -7085
rect 170472 -7173 170559 -7085
rect 170638 -7173 170725 -7085
rect 170818 -7173 170905 -7085
rect 170991 -7176 171078 -7088
rect 171171 -7176 171258 -7088
rect 170292 -7353 170379 -7265
rect 170472 -7353 170559 -7265
rect 170638 -7353 170725 -7265
rect 170818 -7353 170905 -7265
rect 170991 -7356 171078 -7268
rect 171171 -7356 171258 -7268
rect 133379 -13521 133466 -13433
rect 133559 -13521 133646 -13433
rect 133706 -13519 133793 -13431
rect 133886 -13519 133973 -13431
rect 134040 -13518 134127 -13430
rect 133379 -13701 133466 -13613
rect 133559 -13701 133646 -13613
rect 133706 -13699 133793 -13611
rect 133886 -13699 133973 -13611
rect 134040 -13698 134127 -13610
rect 75573 -14813 75660 -14725
rect 75733 -14813 75820 -14725
rect 75893 -14813 75980 -14725
rect 76053 -14813 76140 -14725
rect 76213 -14813 76300 -14725
rect 76373 -14813 76460 -14725
rect 75573 -14973 75660 -14885
rect 75733 -14973 75820 -14885
rect 75893 -14973 75980 -14885
rect 76053 -14973 76140 -14885
rect 76213 -14973 76300 -14885
rect 76373 -14973 76460 -14885
rect 75573 -15133 75660 -15045
rect 75733 -15133 75820 -15045
rect 75893 -15133 75980 -15045
rect 76053 -15133 76140 -15045
rect 76213 -15133 76300 -15045
rect 76373 -15133 76460 -15045
rect 29831 -15449 29918 -15361
rect 29991 -15449 30078 -15361
rect 30151 -15449 30238 -15361
rect 30311 -15449 30398 -15361
rect 30471 -15449 30558 -15361
rect 30631 -15449 30718 -15361
rect 28009 -15566 28096 -15478
rect 28169 -15566 28256 -15478
rect 28329 -15566 28416 -15478
rect 28489 -15566 28576 -15478
rect 28649 -15566 28736 -15478
rect 28809 -15566 28896 -15478
rect 28009 -15726 28096 -15638
rect 28169 -15726 28256 -15638
rect 28329 -15726 28416 -15638
rect 28489 -15726 28576 -15638
rect 28649 -15726 28736 -15638
rect 28809 -15726 28896 -15638
rect 28009 -15886 28096 -15798
rect 28169 -15886 28256 -15798
rect 28329 -15886 28416 -15798
rect 28489 -15886 28576 -15798
rect 28649 -15886 28736 -15798
rect 28809 -15886 28896 -15798
rect 28009 -16046 28096 -15958
rect 28169 -16046 28256 -15958
rect 28329 -16046 28416 -15958
rect 28489 -16046 28576 -15958
rect 28649 -16046 28736 -15958
rect 28809 -16046 28896 -15958
rect 28009 -16206 28096 -16118
rect 28169 -16206 28256 -16118
rect 28329 -16206 28416 -16118
rect 28489 -16206 28576 -16118
rect 28649 -16206 28736 -16118
rect 28809 -16206 28896 -16118
rect 29831 -15609 29918 -15521
rect 29991 -15609 30078 -15521
rect 30151 -15609 30238 -15521
rect 30311 -15609 30398 -15521
rect 30471 -15609 30558 -15521
rect 30631 -15609 30718 -15521
rect 29831 -15769 29918 -15681
rect 29991 -15769 30078 -15681
rect 30151 -15769 30238 -15681
rect 30311 -15769 30398 -15681
rect 30471 -15769 30558 -15681
rect 30631 -15769 30718 -15681
rect 29831 -15929 29918 -15841
rect 29991 -15929 30078 -15841
rect 30151 -15929 30238 -15841
rect 30311 -15929 30398 -15841
rect 30471 -15929 30558 -15841
rect 30631 -15929 30718 -15841
rect 29831 -16089 29918 -16001
rect 29991 -16089 30078 -16001
rect 30151 -16089 30238 -16001
rect 30311 -16089 30398 -16001
rect 30471 -16089 30558 -16001
rect 30631 -16089 30718 -16001
rect 29831 -16249 29918 -16161
rect 29991 -16249 30078 -16161
rect 30151 -16249 30238 -16161
rect 30311 -16249 30398 -16161
rect 30471 -16249 30558 -16161
rect 30631 -16249 30718 -16161
rect 31543 -15363 31630 -15275
rect 31703 -15363 31790 -15275
rect 31863 -15363 31950 -15275
rect 32023 -15363 32110 -15275
rect 32183 -15363 32270 -15275
rect 32343 -15363 32430 -15275
rect 31543 -15523 31630 -15435
rect 31703 -15523 31790 -15435
rect 31863 -15523 31950 -15435
rect 32023 -15523 32110 -15435
rect 32183 -15523 32270 -15435
rect 32343 -15523 32430 -15435
rect 31543 -15683 31630 -15595
rect 31703 -15683 31790 -15595
rect 31863 -15683 31950 -15595
rect 32023 -15683 32110 -15595
rect 32183 -15683 32270 -15595
rect 32343 -15683 32430 -15595
rect 75573 -15293 75660 -15205
rect 75733 -15293 75820 -15205
rect 75893 -15293 75980 -15205
rect 76053 -15293 76140 -15205
rect 76213 -15293 76300 -15205
rect 76373 -15293 76460 -15205
rect 75573 -15453 75660 -15365
rect 75733 -15453 75820 -15365
rect 75893 -15453 75980 -15365
rect 76053 -15453 76140 -15365
rect 76213 -15453 76300 -15365
rect 76373 -15453 76460 -15365
rect 80774 -15027 80861 -14939
rect 80954 -15027 81041 -14939
rect 81101 -15025 81188 -14937
rect 81281 -15025 81368 -14937
rect 81435 -15024 81522 -14936
rect 81605 -15027 81692 -14939
rect 81759 -15026 81846 -14938
rect 80774 -15207 80861 -15119
rect 80954 -15207 81041 -15119
rect 81101 -15205 81188 -15117
rect 81281 -15205 81368 -15117
rect 81435 -15204 81522 -15116
rect 81605 -15207 81692 -15119
rect 81759 -15206 81846 -15118
rect 80768 -15384 80855 -15296
rect 80948 -15384 81035 -15296
rect 81095 -15382 81182 -15294
rect 81275 -15382 81362 -15294
rect 81429 -15381 81516 -15293
rect 81599 -15384 81686 -15296
rect 81753 -15383 81840 -15295
rect 75573 -15613 75660 -15525
rect 75733 -15613 75820 -15525
rect 75893 -15613 75980 -15525
rect 76053 -15613 76140 -15525
rect 76213 -15613 76300 -15525
rect 76373 -15613 76460 -15525
rect 31543 -15843 31630 -15755
rect 31703 -15843 31790 -15755
rect 31863 -15843 31950 -15755
rect 32023 -15843 32110 -15755
rect 32183 -15843 32270 -15755
rect 32343 -15843 32430 -15755
rect 31543 -16003 31630 -15915
rect 31703 -16003 31790 -15915
rect 31863 -16003 31950 -15915
rect 32023 -16003 32110 -15915
rect 32183 -16003 32270 -15915
rect 32343 -16003 32430 -15915
rect 112989 -15778 113072 -15695
rect 113159 -15778 113242 -15695
rect 113329 -15778 113412 -15695
rect 113499 -15778 113582 -15695
rect 113669 -15778 113752 -15695
rect 133361 -13914 133448 -13826
rect 133541 -13914 133628 -13826
rect 133688 -13912 133775 -13824
rect 133868 -13912 133955 -13824
rect 134022 -13911 134109 -13823
rect 133361 -14094 133448 -14006
rect 133541 -14094 133628 -14006
rect 133688 -14092 133775 -14004
rect 133868 -14092 133955 -14004
rect 134022 -14091 134109 -14003
rect 135817 -13526 135904 -13438
rect 135997 -13526 136084 -13438
rect 136144 -13524 136231 -13436
rect 136324 -13524 136411 -13436
rect 136478 -13523 136565 -13435
rect 135817 -13706 135904 -13618
rect 135997 -13706 136084 -13618
rect 136144 -13704 136231 -13616
rect 136324 -13704 136411 -13616
rect 136478 -13703 136565 -13615
rect 135799 -13919 135886 -13831
rect 135979 -13919 136066 -13831
rect 136126 -13917 136213 -13829
rect 136306 -13917 136393 -13829
rect 136460 -13916 136547 -13828
rect 135799 -14099 135886 -14011
rect 135979 -14099 136066 -14011
rect 136126 -14097 136213 -14009
rect 136306 -14097 136393 -14009
rect 136460 -14096 136547 -14008
rect 138539 -13532 138626 -13444
rect 138719 -13532 138806 -13444
rect 138866 -13530 138953 -13442
rect 139046 -13530 139133 -13442
rect 139200 -13529 139287 -13441
rect 138539 -13712 138626 -13624
rect 138719 -13712 138806 -13624
rect 138866 -13710 138953 -13622
rect 139046 -13710 139133 -13622
rect 139200 -13709 139287 -13621
rect 138521 -13925 138608 -13837
rect 138701 -13925 138788 -13837
rect 138848 -13923 138935 -13835
rect 139028 -13923 139115 -13835
rect 139182 -13922 139269 -13834
rect 138521 -14105 138608 -14017
rect 138701 -14105 138788 -14017
rect 138848 -14103 138935 -14015
rect 139028 -14103 139115 -14015
rect 139182 -14102 139269 -14014
rect 150321 -13499 150408 -13411
rect 150501 -13499 150588 -13411
rect 150648 -13497 150735 -13409
rect 150828 -13497 150915 -13409
rect 150982 -13496 151069 -13408
rect 150321 -13679 150408 -13591
rect 150501 -13679 150588 -13591
rect 150648 -13677 150735 -13589
rect 150828 -13677 150915 -13589
rect 150982 -13676 151069 -13588
rect 150303 -13892 150390 -13804
rect 150483 -13892 150570 -13804
rect 150630 -13890 150717 -13802
rect 150810 -13890 150897 -13802
rect 150964 -13889 151051 -13801
rect 150303 -14072 150390 -13984
rect 150483 -14072 150570 -13984
rect 150630 -14070 150717 -13982
rect 150810 -14070 150897 -13982
rect 150964 -14069 151051 -13981
rect 142780 -15036 142863 -14953
rect 142950 -15036 143033 -14953
rect 143120 -15036 143203 -14953
rect 143290 -15036 143373 -14953
rect 143460 -15036 143543 -14953
rect 142780 -15206 142863 -15123
rect 142950 -15206 143033 -15123
rect 143120 -15206 143203 -15123
rect 143290 -15206 143373 -15123
rect 143460 -15206 143543 -15123
rect 142780 -15376 142863 -15293
rect 142950 -15376 143033 -15293
rect 143120 -15376 143203 -15293
rect 143290 -15376 143373 -15293
rect 143460 -15376 143543 -15293
rect 142780 -15546 142863 -15463
rect 142950 -15546 143033 -15463
rect 143120 -15546 143203 -15463
rect 143290 -15546 143373 -15463
rect 143460 -15546 143543 -15463
rect 31543 -16163 31630 -16075
rect 31703 -16163 31790 -16075
rect 31863 -16163 31950 -16075
rect 32023 -16163 32110 -16075
rect 32183 -16163 32270 -16075
rect 32343 -16163 32430 -16075
rect 65092 -16085 65175 -16002
rect 65262 -16085 65345 -16002
rect 65432 -16085 65515 -16002
rect 65602 -16085 65685 -16002
rect 65772 -16085 65855 -16002
rect 65092 -16255 65175 -16172
rect 65262 -16255 65345 -16172
rect 65432 -16255 65515 -16172
rect 65602 -16255 65685 -16172
rect 65772 -16255 65855 -16172
rect 80884 -16053 80971 -15965
rect 81044 -16053 81131 -15965
rect 81204 -16053 81291 -15965
rect 81364 -16053 81451 -15965
rect 81524 -16053 81611 -15965
rect 81684 -16053 81771 -15965
rect 28009 -16366 28096 -16278
rect 28169 -16366 28256 -16278
rect 28329 -16366 28416 -16278
rect 28489 -16366 28576 -16278
rect 28649 -16366 28736 -16278
rect 28809 -16366 28896 -16278
rect 65092 -16425 65175 -16342
rect 65262 -16425 65345 -16342
rect 65432 -16425 65515 -16342
rect 65602 -16425 65685 -16342
rect 65772 -16425 65855 -16342
rect 65092 -16595 65175 -16512
rect 65262 -16595 65345 -16512
rect 65432 -16595 65515 -16512
rect 65602 -16595 65685 -16512
rect 65772 -16595 65855 -16512
rect 65092 -16765 65175 -16682
rect 65262 -16765 65345 -16682
rect 65432 -16765 65515 -16682
rect 65602 -16765 65685 -16682
rect 65772 -16765 65855 -16682
rect 75652 -16355 75739 -16267
rect 75832 -16355 75919 -16267
rect 75979 -16353 76066 -16265
rect 76159 -16353 76246 -16265
rect 76313 -16352 76400 -16264
rect 76483 -16355 76570 -16267
rect 76637 -16354 76724 -16266
rect 75652 -16535 75739 -16447
rect 75832 -16535 75919 -16447
rect 75979 -16533 76066 -16445
rect 76159 -16533 76246 -16445
rect 76313 -16532 76400 -16444
rect 76483 -16535 76570 -16447
rect 76637 -16534 76724 -16446
rect 75646 -16712 75733 -16624
rect 75826 -16712 75913 -16624
rect 75973 -16710 76060 -16622
rect 76153 -16710 76240 -16622
rect 76307 -16709 76394 -16621
rect 76477 -16712 76564 -16624
rect 76631 -16711 76718 -16623
rect 80884 -16213 80971 -16125
rect 81044 -16213 81131 -16125
rect 81204 -16213 81291 -16125
rect 81364 -16213 81451 -16125
rect 81524 -16213 81611 -16125
rect 81684 -16213 81771 -16125
rect 80884 -16373 80971 -16285
rect 81044 -16373 81131 -16285
rect 81204 -16373 81291 -16285
rect 81364 -16373 81451 -16285
rect 81524 -16373 81611 -16285
rect 81684 -16373 81771 -16285
rect 80884 -16533 80971 -16445
rect 81044 -16533 81131 -16445
rect 81204 -16533 81291 -16445
rect 81364 -16533 81451 -16445
rect 81524 -16533 81611 -16445
rect 81684 -16533 81771 -16445
rect 112989 -15948 113072 -15865
rect 113159 -15948 113242 -15865
rect 113329 -15948 113412 -15865
rect 113499 -15948 113582 -15865
rect 113669 -15948 113752 -15865
rect 112989 -16118 113072 -16035
rect 113159 -16118 113242 -16035
rect 113329 -16118 113412 -16035
rect 113499 -16118 113582 -16035
rect 113669 -16118 113752 -16035
rect 112989 -16288 113072 -16205
rect 113159 -16288 113242 -16205
rect 113329 -16288 113412 -16205
rect 113499 -16288 113582 -16205
rect 113669 -16288 113752 -16205
rect 112989 -16458 113072 -16375
rect 113159 -16458 113242 -16375
rect 113329 -16458 113412 -16375
rect 113499 -16458 113582 -16375
rect 113669 -16458 113752 -16375
rect 116719 -15813 116802 -15730
rect 116889 -15813 116972 -15730
rect 117059 -15813 117142 -15730
rect 117229 -15813 117312 -15730
rect 117399 -15813 117482 -15730
rect 142780 -15716 142863 -15633
rect 142950 -15716 143033 -15633
rect 143120 -15716 143203 -15633
rect 143290 -15716 143373 -15633
rect 143460 -15716 143543 -15633
rect 144826 -15014 144909 -14931
rect 144996 -15014 145079 -14931
rect 145166 -15014 145249 -14931
rect 145336 -15014 145419 -14931
rect 145506 -15014 145589 -14931
rect 144826 -15184 144909 -15101
rect 144996 -15184 145079 -15101
rect 145166 -15184 145249 -15101
rect 145336 -15184 145419 -15101
rect 145506 -15184 145589 -15101
rect 144826 -15354 144909 -15271
rect 144996 -15354 145079 -15271
rect 145166 -15354 145249 -15271
rect 145336 -15354 145419 -15271
rect 145506 -15354 145589 -15271
rect 144826 -15524 144909 -15441
rect 144996 -15524 145079 -15441
rect 145166 -15524 145249 -15441
rect 145336 -15524 145419 -15441
rect 145506 -15524 145589 -15441
rect 144826 -15694 144909 -15611
rect 144996 -15694 145079 -15611
rect 145166 -15694 145249 -15611
rect 145336 -15694 145419 -15611
rect 145506 -15694 145589 -15611
rect 146960 -14993 147043 -14910
rect 147130 -14993 147213 -14910
rect 147300 -14993 147383 -14910
rect 147470 -14993 147553 -14910
rect 147640 -14993 147723 -14910
rect 146960 -15163 147043 -15080
rect 147130 -15163 147213 -15080
rect 147300 -15163 147383 -15080
rect 147470 -15163 147553 -15080
rect 147640 -15163 147723 -15080
rect 146960 -15333 147043 -15250
rect 147130 -15333 147213 -15250
rect 147300 -15333 147383 -15250
rect 147470 -15333 147553 -15250
rect 147640 -15333 147723 -15250
rect 146960 -15503 147043 -15420
rect 147130 -15503 147213 -15420
rect 147300 -15503 147383 -15420
rect 147470 -15503 147553 -15420
rect 147640 -15503 147723 -15420
rect 146960 -15673 147043 -15590
rect 147130 -15673 147213 -15590
rect 147300 -15673 147383 -15590
rect 147470 -15673 147553 -15590
rect 147640 -15673 147723 -15590
rect 116719 -15983 116802 -15900
rect 116889 -15983 116972 -15900
rect 117059 -15983 117142 -15900
rect 117229 -15983 117312 -15900
rect 117399 -15983 117482 -15900
rect 116719 -16153 116802 -16070
rect 116889 -16153 116972 -16070
rect 117059 -16153 117142 -16070
rect 117229 -16153 117312 -16070
rect 117399 -16153 117482 -16070
rect 116719 -16323 116802 -16240
rect 116889 -16323 116972 -16240
rect 117059 -16323 117142 -16240
rect 117229 -16323 117312 -16240
rect 117399 -16323 117482 -16240
rect 116719 -16493 116802 -16410
rect 116889 -16493 116972 -16410
rect 117059 -16493 117142 -16410
rect 117229 -16493 117312 -16410
rect 117399 -16493 117482 -16410
rect 80884 -16693 80971 -16605
rect 81044 -16693 81131 -16605
rect 81204 -16693 81291 -16605
rect 81364 -16693 81451 -16605
rect 81524 -16693 81611 -16605
rect 81684 -16693 81771 -16605
rect 80884 -16853 80971 -16765
rect 81044 -16853 81131 -16765
rect 81204 -16853 81291 -16765
rect 81364 -16853 81451 -16765
rect 81524 -16853 81611 -16765
rect 81684 -16853 81771 -16765
rect 16104 -17086 16187 -17003
rect 16274 -17086 16357 -17003
rect 16444 -17086 16527 -17003
rect 16614 -17086 16697 -17003
rect 16784 -17086 16867 -17003
rect -5099 -17312 -5016 -17229
rect -4929 -17312 -4846 -17229
rect -4759 -17312 -4676 -17229
rect -4589 -17312 -4506 -17229
rect -4419 -17312 -4336 -17229
rect -5099 -17482 -5016 -17399
rect -4929 -17482 -4846 -17399
rect -4759 -17482 -4676 -17399
rect -4589 -17482 -4506 -17399
rect -4419 -17482 -4336 -17399
rect 16104 -17256 16187 -17173
rect 16274 -17256 16357 -17173
rect 16444 -17256 16527 -17173
rect 16614 -17256 16697 -17173
rect 16784 -17256 16867 -17173
rect 16104 -17426 16187 -17343
rect 16274 -17426 16357 -17343
rect 16444 -17426 16527 -17343
rect 16614 -17426 16697 -17343
rect 16784 -17426 16867 -17343
rect -5099 -17652 -5016 -17569
rect -4929 -17652 -4846 -17569
rect -4759 -17652 -4676 -17569
rect -4589 -17652 -4506 -17569
rect -4419 -17652 -4336 -17569
rect -1129 -17580 -1073 -17524
rect -1025 -17580 -969 -17524
rect -921 -17580 -865 -17524
rect -1129 -17684 -1073 -17628
rect -1025 -17684 -969 -17628
rect -921 -17684 -865 -17628
rect -5099 -17822 -5016 -17739
rect -4929 -17822 -4846 -17739
rect -4759 -17822 -4676 -17739
rect -4589 -17822 -4506 -17739
rect -4419 -17822 -4336 -17739
rect -1129 -17788 -1073 -17732
rect -1025 -17788 -969 -17732
rect -921 -17788 -865 -17732
rect 16104 -17596 16187 -17513
rect 16274 -17596 16357 -17513
rect 16444 -17596 16527 -17513
rect 16614 -17596 16697 -17513
rect 16784 -17596 16867 -17513
rect 16104 -17766 16187 -17683
rect 16274 -17766 16357 -17683
rect 16444 -17766 16527 -17683
rect 16614 -17766 16697 -17683
rect 16784 -17766 16867 -17683
rect 18010 -17094 18093 -17011
rect 18180 -17094 18263 -17011
rect 18350 -17094 18433 -17011
rect 18520 -17094 18603 -17011
rect 18690 -17094 18773 -17011
rect 18010 -17264 18093 -17181
rect 18180 -17264 18263 -17181
rect 18350 -17264 18433 -17181
rect 18520 -17264 18603 -17181
rect 18690 -17264 18773 -17181
rect 18010 -17434 18093 -17351
rect 18180 -17434 18263 -17351
rect 18350 -17434 18433 -17351
rect 18520 -17434 18603 -17351
rect 18690 -17434 18773 -17351
rect 18010 -17604 18093 -17521
rect 18180 -17604 18263 -17521
rect 18350 -17604 18433 -17521
rect 18520 -17604 18603 -17521
rect 18690 -17604 18773 -17521
rect 18010 -17774 18093 -17691
rect 18180 -17774 18263 -17691
rect 18350 -17774 18433 -17691
rect 18520 -17774 18603 -17691
rect 18690 -17774 18773 -17691
rect 20082 -17070 20165 -16987
rect 20252 -17070 20335 -16987
rect 20422 -17070 20505 -16987
rect 20592 -17070 20675 -16987
rect 20762 -17070 20845 -16987
rect 20082 -17240 20165 -17157
rect 20252 -17240 20335 -17157
rect 20422 -17240 20505 -17157
rect 20592 -17240 20675 -17157
rect 20762 -17240 20845 -17157
rect 20082 -17410 20165 -17327
rect 20252 -17410 20335 -17327
rect 20422 -17410 20505 -17327
rect 20592 -17410 20675 -17327
rect 20762 -17410 20845 -17327
rect 20082 -17580 20165 -17497
rect 20252 -17580 20335 -17497
rect 20422 -17580 20505 -17497
rect 20592 -17580 20675 -17497
rect 20762 -17580 20845 -17497
rect 20082 -17750 20165 -17667
rect 20252 -17750 20335 -17667
rect 20422 -17750 20505 -17667
rect 20592 -17750 20675 -17667
rect 20762 -17750 20845 -17667
rect -5099 -17992 -5016 -17909
rect -4929 -17992 -4846 -17909
rect -4759 -17992 -4676 -17909
rect -4589 -17992 -4506 -17909
rect -4419 -17992 -4336 -17909
rect 27290 -18251 27377 -18163
rect 27450 -18251 27537 -18163
rect 27610 -18251 27697 -18163
rect 27770 -18251 27857 -18163
rect 27930 -18251 28017 -18163
rect 28090 -18251 28177 -18163
rect 312 -18432 395 -18349
rect 482 -18432 565 -18349
rect 652 -18432 735 -18349
rect 822 -18432 905 -18349
rect 992 -18432 1075 -18349
rect 312 -18602 395 -18519
rect 482 -18602 565 -18519
rect 652 -18602 735 -18519
rect 822 -18602 905 -18519
rect 992 -18602 1075 -18519
rect 312 -18772 395 -18689
rect 482 -18772 565 -18689
rect 652 -18772 735 -18689
rect 822 -18772 905 -18689
rect 992 -18772 1075 -18689
rect 312 -18942 395 -18859
rect 482 -18942 565 -18859
rect 652 -18942 735 -18859
rect 822 -18942 905 -18859
rect 992 -18942 1075 -18859
rect 312 -19112 395 -19029
rect 482 -19112 565 -19029
rect 652 -19112 735 -19029
rect 822 -19112 905 -19029
rect 992 -19112 1075 -19029
rect 27290 -18411 27377 -18323
rect 27450 -18411 27537 -18323
rect 27610 -18411 27697 -18323
rect 27770 -18411 27857 -18323
rect 27930 -18411 28017 -18323
rect 28090 -18411 28177 -18323
rect 27290 -18571 27377 -18483
rect 27450 -18571 27537 -18483
rect 27610 -18571 27697 -18483
rect 27770 -18571 27857 -18483
rect 27930 -18571 28017 -18483
rect 28090 -18571 28177 -18483
rect 27290 -18731 27377 -18643
rect 27450 -18731 27537 -18643
rect 27610 -18731 27697 -18643
rect 27770 -18731 27857 -18643
rect 27930 -18731 28017 -18643
rect 28090 -18731 28177 -18643
rect 27290 -18891 27377 -18803
rect 27450 -18891 27537 -18803
rect 27610 -18891 27697 -18803
rect 27770 -18891 27857 -18803
rect 27930 -18891 28017 -18803
rect 28090 -18891 28177 -18803
rect 27290 -19051 27377 -18963
rect 27450 -19051 27537 -18963
rect 27610 -19051 27697 -18963
rect 27770 -19051 27857 -18963
rect 27930 -19051 28017 -18963
rect 28090 -19051 28177 -18963
rect 27933 -19537 28020 -19449
rect 28113 -19537 28200 -19449
rect 28260 -19535 28347 -19447
rect 28440 -19535 28527 -19447
rect 28594 -19534 28681 -19446
<< metal3 >>
rect 1963 17608 2630 18311
rect 1898 17585 2709 17608
rect 4106 17590 4773 18293
rect 1898 17502 1922 17585
rect 2005 17502 2092 17585
rect 2175 17502 2262 17585
rect 2345 17502 2432 17585
rect 2515 17502 2602 17585
rect 2685 17502 2709 17585
rect 1898 17415 2709 17502
rect 1898 17332 1922 17415
rect 2005 17332 2092 17415
rect 2175 17332 2262 17415
rect 2345 17332 2432 17415
rect 2515 17332 2602 17415
rect 2685 17332 2709 17415
rect 1898 17245 2709 17332
rect 1898 17162 1922 17245
rect 2005 17162 2092 17245
rect 2175 17162 2262 17245
rect 2345 17162 2432 17245
rect 2515 17162 2602 17245
rect 2685 17162 2709 17245
rect 1898 17075 2709 17162
rect 1898 16992 1922 17075
rect 2005 16992 2092 17075
rect 2175 16992 2262 17075
rect 2345 16992 2432 17075
rect 2515 16992 2602 17075
rect 2685 16992 2709 17075
rect 1898 16905 2709 16992
rect 1898 16822 1922 16905
rect 2005 16822 2092 16905
rect 2175 16822 2262 16905
rect 2345 16822 2432 16905
rect 2515 16822 2602 16905
rect 2685 16822 2709 16905
rect 1898 16799 2709 16822
rect 4041 17567 4852 17590
rect 4041 17484 4065 17567
rect 4148 17484 4235 17567
rect 4318 17484 4405 17567
rect 4488 17484 4575 17567
rect 4658 17484 4745 17567
rect 4828 17484 4852 17567
rect 4041 17397 4852 17484
rect 4041 17314 4065 17397
rect 4148 17314 4235 17397
rect 4318 17314 4405 17397
rect 4488 17314 4575 17397
rect 4658 17314 4745 17397
rect 4828 17314 4852 17397
rect 4041 17227 4852 17314
rect 18041 17308 18708 18011
rect 4041 17144 4065 17227
rect 4148 17144 4235 17227
rect 4318 17144 4405 17227
rect 4488 17144 4575 17227
rect 4658 17144 4745 17227
rect 4828 17144 4852 17227
rect 4041 17057 4852 17144
rect 4041 16974 4065 17057
rect 4148 16974 4235 17057
rect 4318 16974 4405 17057
rect 4488 16974 4575 17057
rect 4658 16974 4745 17057
rect 4828 16974 4852 17057
rect 4041 16887 4852 16974
rect 4041 16804 4065 16887
rect 4148 16804 4235 16887
rect 4318 16804 4405 16887
rect 4488 16804 4575 16887
rect 4658 16804 4745 16887
rect 4828 16804 4852 16887
rect 4041 16781 4852 16804
rect 17976 17285 18787 17308
rect 17976 17202 18000 17285
rect 18083 17202 18170 17285
rect 18253 17202 18340 17285
rect 18423 17202 18510 17285
rect 18593 17202 18680 17285
rect 18763 17202 18787 17285
rect 22045 17244 22712 17947
rect 85688 17391 86355 18094
rect 85623 17368 86434 17391
rect 89305 17382 89972 18085
rect 85623 17285 85647 17368
rect 85730 17285 85817 17368
rect 85900 17285 85987 17368
rect 86070 17285 86157 17368
rect 86240 17285 86327 17368
rect 86410 17285 86434 17368
rect 17976 17115 18787 17202
rect 17976 17032 18000 17115
rect 18083 17032 18170 17115
rect 18253 17032 18340 17115
rect 18423 17032 18510 17115
rect 18593 17032 18680 17115
rect 18763 17032 18787 17115
rect 17976 16945 18787 17032
rect 17976 16862 18000 16945
rect 18083 16862 18170 16945
rect 18253 16862 18340 16945
rect 18423 16862 18510 16945
rect 18593 16862 18680 16945
rect 18763 16862 18787 16945
rect 17976 16775 18787 16862
rect 17976 16692 18000 16775
rect 18083 16692 18170 16775
rect 18253 16692 18340 16775
rect 18423 16692 18510 16775
rect 18593 16692 18680 16775
rect 18763 16692 18787 16775
rect 17976 16605 18787 16692
rect 17976 16522 18000 16605
rect 18083 16522 18170 16605
rect 18253 16522 18340 16605
rect 18423 16522 18510 16605
rect 18593 16522 18680 16605
rect 18763 16522 18787 16605
rect 17976 16499 18787 16522
rect 21980 17221 22791 17244
rect 21980 17138 22004 17221
rect 22087 17138 22174 17221
rect 22257 17138 22344 17221
rect 22427 17138 22514 17221
rect 22597 17138 22684 17221
rect 22767 17138 22791 17221
rect 21980 17051 22791 17138
rect 85623 17198 86434 17285
rect 85623 17115 85647 17198
rect 85730 17115 85817 17198
rect 85900 17115 85987 17198
rect 86070 17115 86157 17198
rect 86240 17115 86327 17198
rect 86410 17115 86434 17198
rect 21980 16968 22004 17051
rect 22087 16968 22174 17051
rect 22257 16968 22344 17051
rect 22427 16968 22514 17051
rect 22597 16968 22684 17051
rect 22767 16968 22791 17051
rect 21980 16881 22791 16968
rect 21980 16798 22004 16881
rect 22087 16798 22174 16881
rect 22257 16798 22344 16881
rect 22427 16798 22514 16881
rect 22597 16798 22684 16881
rect 22767 16798 22791 16881
rect 21980 16711 22791 16798
rect 21980 16628 22004 16711
rect 22087 16628 22174 16711
rect 22257 16628 22344 16711
rect 22427 16628 22514 16711
rect 22597 16628 22684 16711
rect 22767 16628 22791 16711
rect 21980 16541 22791 16628
rect 21980 16458 22004 16541
rect 22087 16458 22174 16541
rect 22257 16458 22344 16541
rect 22427 16458 22514 16541
rect 22597 16458 22684 16541
rect 22767 16458 22791 16541
rect 21980 16435 22791 16458
rect 49232 16327 49899 17030
rect 52386 16355 53053 17058
rect 85623 17028 86434 17115
rect 85623 16945 85647 17028
rect 85730 16945 85817 17028
rect 85900 16945 85987 17028
rect 86070 16945 86157 17028
rect 86240 16945 86327 17028
rect 86410 16945 86434 17028
rect 85623 16858 86434 16945
rect 85623 16775 85647 16858
rect 85730 16775 85817 16858
rect 85900 16775 85987 16858
rect 86070 16775 86157 16858
rect 86240 16775 86327 16858
rect 86410 16775 86434 16858
rect 85623 16688 86434 16775
rect 85623 16605 85647 16688
rect 85730 16605 85817 16688
rect 85900 16605 85987 16688
rect 86070 16605 86157 16688
rect 86240 16605 86327 16688
rect 86410 16605 86434 16688
rect 85623 16582 86434 16605
rect 89240 17359 90051 17382
rect 89240 17276 89264 17359
rect 89347 17276 89434 17359
rect 89517 17276 89604 17359
rect 89687 17276 89774 17359
rect 89857 17276 89944 17359
rect 90027 17276 90051 17359
rect 89240 17189 90051 17276
rect 89240 17106 89264 17189
rect 89347 17106 89434 17189
rect 89517 17106 89604 17189
rect 89687 17106 89774 17189
rect 89857 17106 89944 17189
rect 90027 17106 90051 17189
rect 155009 17186 155676 17889
rect 157384 17186 158051 17889
rect 89240 17019 90051 17106
rect 89240 16936 89264 17019
rect 89347 16936 89434 17019
rect 89517 16936 89604 17019
rect 89687 16936 89774 17019
rect 89857 16936 89944 17019
rect 90027 16936 90051 17019
rect 89240 16849 90051 16936
rect 89240 16766 89264 16849
rect 89347 16766 89434 16849
rect 89517 16766 89604 16849
rect 89687 16766 89774 16849
rect 89857 16766 89944 16849
rect 90027 16766 90051 16849
rect 89240 16679 90051 16766
rect 89240 16596 89264 16679
rect 89347 16596 89434 16679
rect 89517 16596 89604 16679
rect 89687 16596 89774 16679
rect 89857 16596 89944 16679
rect 90027 16596 90051 16679
rect 89240 16573 90051 16596
rect 154944 17163 155755 17186
rect 154944 17080 154968 17163
rect 155051 17080 155138 17163
rect 155221 17080 155308 17163
rect 155391 17080 155478 17163
rect 155561 17080 155648 17163
rect 155731 17080 155755 17163
rect 154944 16993 155755 17080
rect 154944 16910 154968 16993
rect 155051 16910 155138 16993
rect 155221 16910 155308 16993
rect 155391 16910 155478 16993
rect 155561 16910 155648 16993
rect 155731 16910 155755 16993
rect 154944 16823 155755 16910
rect 154944 16740 154968 16823
rect 155051 16740 155138 16823
rect 155221 16740 155308 16823
rect 155391 16740 155478 16823
rect 155561 16740 155648 16823
rect 155731 16740 155755 16823
rect 154944 16653 155755 16740
rect 154944 16570 154968 16653
rect 155051 16570 155138 16653
rect 155221 16570 155308 16653
rect 155391 16570 155478 16653
rect 155561 16570 155648 16653
rect 155731 16570 155755 16653
rect 154944 16483 155755 16570
rect 154944 16400 154968 16483
rect 155051 16400 155138 16483
rect 155221 16400 155308 16483
rect 155391 16400 155478 16483
rect 155561 16400 155648 16483
rect 155731 16400 155755 16483
rect 154944 16377 155755 16400
rect 157319 17163 158130 17186
rect 157319 17080 157343 17163
rect 157426 17080 157513 17163
rect 157596 17080 157683 17163
rect 157766 17080 157853 17163
rect 157936 17080 158023 17163
rect 158106 17080 158130 17163
rect 157319 16993 158130 17080
rect 157319 16910 157343 16993
rect 157426 16910 157513 16993
rect 157596 16910 157683 16993
rect 157766 16910 157853 16993
rect 157936 16910 158023 16993
rect 158106 16910 158130 16993
rect 157319 16823 158130 16910
rect 157319 16740 157343 16823
rect 157426 16740 157513 16823
rect 157596 16740 157683 16823
rect 157766 16740 157853 16823
rect 157936 16740 158023 16823
rect 158106 16740 158130 16823
rect 157319 16653 158130 16740
rect 157319 16570 157343 16653
rect 157426 16570 157513 16653
rect 157596 16570 157683 16653
rect 157766 16570 157853 16653
rect 157936 16570 158023 16653
rect 158106 16570 158130 16653
rect 157319 16483 158130 16570
rect 157319 16400 157343 16483
rect 157426 16400 157513 16483
rect 157596 16400 157683 16483
rect 157766 16400 157853 16483
rect 157936 16400 158023 16483
rect 158106 16400 158130 16483
rect 157319 16377 158130 16400
rect 52321 16332 53132 16355
rect 49167 16304 49978 16327
rect 49167 16221 49191 16304
rect 49274 16221 49361 16304
rect 49444 16221 49531 16304
rect 49614 16221 49701 16304
rect 49784 16221 49871 16304
rect 49954 16221 49978 16304
rect 49167 16134 49978 16221
rect 49167 16051 49191 16134
rect 49274 16051 49361 16134
rect 49444 16051 49531 16134
rect 49614 16051 49701 16134
rect 49784 16051 49871 16134
rect 49954 16051 49978 16134
rect 49167 15964 49978 16051
rect 49167 15881 49191 15964
rect 49274 15881 49361 15964
rect 49444 15881 49531 15964
rect 49614 15881 49701 15964
rect 49784 15881 49871 15964
rect 49954 15881 49978 15964
rect -608 15781 -319 15799
rect -608 15725 -597 15781
rect -541 15725 -493 15781
rect -437 15725 -389 15781
rect -333 15725 -319 15781
rect -4959 15658 -4150 15682
rect -4959 15603 -4936 15658
rect -5662 15575 -4936 15603
rect -4853 15575 -4766 15658
rect -4683 15575 -4596 15658
rect -4513 15575 -4426 15658
rect -4343 15575 -4256 15658
rect -4173 15575 -4150 15658
rect -5662 15488 -4150 15575
rect -608 15677 -319 15725
rect -608 15621 -597 15677
rect -541 15621 -493 15677
rect -437 15621 -389 15677
rect -333 15621 -319 15677
rect -608 15573 -319 15621
rect -608 15517 -597 15573
rect -541 15517 -493 15573
rect -437 15517 -389 15573
rect -333 15517 -319 15573
rect 49167 15794 49978 15881
rect 49167 15711 49191 15794
rect 49274 15711 49361 15794
rect 49444 15711 49531 15794
rect 49614 15711 49701 15794
rect 49784 15711 49871 15794
rect 49954 15711 49978 15794
rect 49167 15624 49978 15711
rect 49167 15541 49191 15624
rect 49274 15541 49361 15624
rect 49444 15541 49531 15624
rect 49614 15541 49701 15624
rect 49784 15541 49871 15624
rect 49954 15541 49978 15624
rect 52321 16249 52345 16332
rect 52428 16249 52515 16332
rect 52598 16249 52685 16332
rect 52768 16249 52855 16332
rect 52938 16249 53025 16332
rect 53108 16249 53132 16332
rect 52321 16162 53132 16249
rect 52321 16079 52345 16162
rect 52428 16079 52515 16162
rect 52598 16079 52685 16162
rect 52768 16079 52855 16162
rect 52938 16079 53025 16162
rect 53108 16079 53132 16162
rect 52321 15992 53132 16079
rect 52321 15909 52345 15992
rect 52428 15909 52515 15992
rect 52598 15909 52685 15992
rect 52768 15909 52855 15992
rect 52938 15909 53025 15992
rect 53108 15909 53132 15992
rect 52321 15822 53132 15909
rect 52321 15739 52345 15822
rect 52428 15739 52515 15822
rect 52598 15739 52685 15822
rect 52768 15739 52855 15822
rect 52938 15739 53025 15822
rect 53108 15739 53132 15822
rect 52321 15652 53132 15739
rect 52321 15569 52345 15652
rect 52428 15569 52515 15652
rect 52598 15569 52685 15652
rect 52768 15569 52855 15652
rect 52938 15569 53025 15652
rect 53108 15569 53132 15652
rect 52321 15546 53132 15569
rect 49167 15518 49978 15541
rect -608 15505 -319 15517
rect -5662 15405 -4936 15488
rect -4853 15405 -4766 15488
rect -4683 15405 -4596 15488
rect -4513 15405 -4426 15488
rect -4343 15405 -4256 15488
rect -4173 15405 -4150 15488
rect -5662 15318 -4150 15405
rect -5662 15235 -4936 15318
rect -4853 15235 -4766 15318
rect -4683 15235 -4596 15318
rect -4513 15235 -4426 15318
rect -4343 15235 -4256 15318
rect -4173 15235 -4150 15318
rect -5662 15148 -4150 15235
rect -5662 15065 -4936 15148
rect -4853 15065 -4766 15148
rect -4683 15065 -4596 15148
rect -4513 15065 -4426 15148
rect -4343 15065 -4256 15148
rect -4173 15065 -4150 15148
rect -5662 14978 -4150 15065
rect -3549 15304 -3260 15322
rect -3549 15248 -3538 15304
rect -3482 15248 -3434 15304
rect -3378 15248 -3330 15304
rect -3274 15248 -3260 15304
rect -3549 15200 -3260 15248
rect -3549 15144 -3538 15200
rect -3482 15144 -3434 15200
rect -3378 15144 -3330 15200
rect -3274 15144 -3260 15200
rect -3549 15096 -3260 15144
rect -3549 15040 -3538 15096
rect -3482 15040 -3434 15096
rect -3378 15040 -3330 15096
rect -3274 15040 -3260 15096
rect -3549 15028 -3260 15040
rect -5662 14936 -4936 14978
rect -4959 14895 -4936 14936
rect -4853 14895 -4766 14978
rect -4683 14895 -4596 14978
rect -4513 14895 -4426 14978
rect -4343 14895 -4256 14978
rect -4173 14895 -4150 14978
rect -4959 14871 -4150 14895
rect -4976 12724 -4167 12748
rect -4976 12669 -4953 12724
rect -5679 12641 -4953 12669
rect -4870 12641 -4783 12724
rect -4700 12641 -4613 12724
rect -4530 12641 -4443 12724
rect -4360 12641 -4273 12724
rect -4190 12641 -4167 12724
rect -5679 12554 -4167 12641
rect -5679 12471 -4953 12554
rect -4870 12471 -4783 12554
rect -4700 12471 -4613 12554
rect -4530 12471 -4443 12554
rect -4360 12471 -4273 12554
rect -4190 12471 -4167 12554
rect -5679 12384 -4167 12471
rect -5679 12301 -4953 12384
rect -4870 12301 -4783 12384
rect -4700 12301 -4613 12384
rect -4530 12301 -4443 12384
rect -4360 12301 -4273 12384
rect -4190 12301 -4167 12384
rect -5679 12214 -4167 12301
rect -5679 12131 -4953 12214
rect -4870 12131 -4783 12214
rect -4700 12131 -4613 12214
rect -4530 12131 -4443 12214
rect -4360 12131 -4273 12214
rect -4190 12131 -4167 12214
rect -5679 12044 -4167 12131
rect -5679 12002 -4953 12044
rect -4976 11961 -4953 12002
rect -4870 11961 -4783 12044
rect -4700 11961 -4613 12044
rect -4530 11961 -4443 12044
rect -4360 11961 -4273 12044
rect -4190 11961 -4167 12044
rect -4976 11937 -4167 11961
rect -4976 9352 -4167 9376
rect -4976 9297 -4953 9352
rect -5679 9269 -4953 9297
rect -4870 9269 -4783 9352
rect -4700 9269 -4613 9352
rect -4530 9269 -4443 9352
rect -4360 9269 -4273 9352
rect -4190 9269 -4167 9352
rect -5679 9182 -4167 9269
rect -5679 9099 -4953 9182
rect -4870 9099 -4783 9182
rect -4700 9099 -4613 9182
rect -4530 9099 -4443 9182
rect -4360 9099 -4273 9182
rect -4190 9099 -4167 9182
rect -5679 9012 -4167 9099
rect -5679 8929 -4953 9012
rect -4870 8929 -4783 9012
rect -4700 8929 -4613 9012
rect -4530 8929 -4443 9012
rect -4360 8929 -4273 9012
rect -4190 8929 -4167 9012
rect -5679 8842 -4167 8929
rect -5679 8759 -4953 8842
rect -4870 8759 -4783 8842
rect -4700 8759 -4613 8842
rect -4530 8759 -4443 8842
rect -4360 8759 -4273 8842
rect -4190 8759 -4167 8842
rect -5679 8672 -4167 8759
rect -5679 8630 -4953 8672
rect -4976 8589 -4953 8630
rect -4870 8589 -4783 8672
rect -4700 8589 -4613 8672
rect -4530 8589 -4443 8672
rect -4360 8589 -4273 8672
rect -4190 8589 -4167 8672
rect -4976 8565 -4167 8589
rect -5044 7042 -4235 7066
rect -5044 6987 -5021 7042
rect -5747 6959 -5021 6987
rect -4938 6959 -4851 7042
rect -4768 6959 -4681 7042
rect -4598 6959 -4511 7042
rect -4428 6959 -4341 7042
rect -4258 6959 -4235 7042
rect -5747 6872 -4235 6959
rect -5747 6789 -5021 6872
rect -4938 6789 -4851 6872
rect -4768 6789 -4681 6872
rect -4598 6789 -4511 6872
rect -4428 6789 -4341 6872
rect -4258 6789 -4235 6872
rect -5747 6702 -4235 6789
rect -5747 6619 -5021 6702
rect -4938 6619 -4851 6702
rect -4768 6619 -4681 6702
rect -4598 6619 -4511 6702
rect -4428 6619 -4341 6702
rect -4258 6619 -4235 6702
rect -5747 6532 -4235 6619
rect -5747 6449 -5021 6532
rect -4938 6449 -4851 6532
rect -4768 6449 -4681 6532
rect -4598 6449 -4511 6532
rect -4428 6449 -4341 6532
rect -4258 6449 -4235 6532
rect -5747 6362 -4235 6449
rect -5747 6320 -5021 6362
rect -5044 6279 -5021 6320
rect -4938 6279 -4851 6362
rect -4768 6279 -4681 6362
rect -4598 6279 -4511 6362
rect -4428 6279 -4341 6362
rect -4258 6279 -4235 6362
rect -5044 6255 -4235 6279
rect -5027 5290 -4218 5314
rect -5027 5235 -5004 5290
rect -5730 5207 -5004 5235
rect -4921 5207 -4834 5290
rect -4751 5207 -4664 5290
rect -4581 5207 -4494 5290
rect -4411 5207 -4324 5290
rect -4241 5207 -4218 5290
rect -5730 5120 -4218 5207
rect -5730 5037 -5004 5120
rect -4921 5037 -4834 5120
rect -4751 5037 -4664 5120
rect -4581 5037 -4494 5120
rect -4411 5037 -4324 5120
rect -4241 5037 -4218 5120
rect -5730 4950 -4218 5037
rect -5730 4867 -5004 4950
rect -4921 4867 -4834 4950
rect -4751 4867 -4664 4950
rect -4581 4867 -4494 4950
rect -4411 4867 -4324 4950
rect -4241 4867 -4218 4950
rect -5730 4780 -4218 4867
rect -5730 4697 -5004 4780
rect -4921 4697 -4834 4780
rect -4751 4697 -4664 4780
rect -4581 4697 -4494 4780
rect -4411 4697 -4324 4780
rect -4241 4697 -4218 4780
rect -5730 4610 -4218 4697
rect -5730 4568 -5004 4610
rect -5027 4527 -5004 4568
rect -4921 4527 -4834 4610
rect -4751 4527 -4664 4610
rect -4581 4527 -4494 4610
rect -4411 4527 -4324 4610
rect -4241 4527 -4218 4610
rect -5027 4503 -4218 4527
rect -5178 2777 -4369 2801
rect -5178 2722 -5155 2777
rect -5881 2694 -5155 2722
rect -5072 2694 -4985 2777
rect -4902 2694 -4815 2777
rect -4732 2694 -4645 2777
rect -4562 2694 -4475 2777
rect -4392 2694 -4369 2777
rect -5881 2607 -4369 2694
rect -5881 2524 -5155 2607
rect -5072 2524 -4985 2607
rect -4902 2524 -4815 2607
rect -4732 2524 -4645 2607
rect -4562 2524 -4475 2607
rect -4392 2524 -4369 2607
rect -5881 2437 -4369 2524
rect -5881 2354 -5155 2437
rect -5072 2354 -4985 2437
rect -4902 2354 -4815 2437
rect -4732 2354 -4645 2437
rect -4562 2354 -4475 2437
rect -4392 2354 -4369 2437
rect -5881 2267 -4369 2354
rect -5881 2184 -5155 2267
rect -5072 2184 -4985 2267
rect -4902 2184 -4815 2267
rect -4732 2184 -4645 2267
rect -4562 2184 -4475 2267
rect -4392 2184 -4369 2267
rect -5881 2097 -4369 2184
rect -5881 2055 -5155 2097
rect -5178 2014 -5155 2055
rect -5072 2014 -4985 2097
rect -4902 2014 -4815 2097
rect -4732 2014 -4645 2097
rect -4562 2014 -4475 2097
rect -4392 2014 -4369 2097
rect -5178 1990 -4369 2014
rect -5178 -1641 -4369 -1617
rect -5178 -1696 -5155 -1641
rect -5881 -1724 -5155 -1696
rect -5072 -1724 -4985 -1641
rect -4902 -1724 -4815 -1641
rect -4732 -1724 -4645 -1641
rect -4562 -1724 -4475 -1641
rect -4392 -1724 -4369 -1641
rect -5881 -1811 -4369 -1724
rect -5881 -1894 -5155 -1811
rect -5072 -1894 -4985 -1811
rect -4902 -1894 -4815 -1811
rect -4732 -1894 -4645 -1811
rect -4562 -1894 -4475 -1811
rect -4392 -1894 -4369 -1811
rect -5881 -1981 -4369 -1894
rect -5881 -2064 -5155 -1981
rect -5072 -2064 -4985 -1981
rect -4902 -2064 -4815 -1981
rect -4732 -2064 -4645 -1981
rect -4562 -2064 -4475 -1981
rect -4392 -2064 -4369 -1981
rect -5881 -2151 -4369 -2064
rect -5881 -2234 -5155 -2151
rect -5072 -2234 -4985 -2151
rect -4902 -2234 -4815 -2151
rect -4732 -2234 -4645 -2151
rect -4562 -2234 -4475 -2151
rect -4392 -2234 -4369 -2151
rect -5881 -2321 -4369 -2234
rect -5881 -2363 -5155 -2321
rect -5178 -2404 -5155 -2363
rect -5072 -2404 -4985 -2321
rect -4902 -2404 -4815 -2321
rect -4732 -2404 -4645 -2321
rect -4562 -2404 -4475 -2321
rect -4392 -2404 -4369 -2321
rect -5178 -2428 -4369 -2404
rect -3527 -2586 -3269 15028
rect -2486 14729 -2197 14747
rect -2486 14673 -2475 14729
rect -2419 14673 -2371 14729
rect -2315 14673 -2267 14729
rect -2211 14673 -2197 14729
rect -2486 14625 -2197 14673
rect -2486 14569 -2475 14625
rect -2419 14569 -2371 14625
rect -2315 14569 -2267 14625
rect -2211 14569 -2197 14625
rect -2486 14521 -2197 14569
rect -2486 14465 -2475 14521
rect -2419 14465 -2371 14521
rect -2315 14465 -2267 14521
rect -2211 14465 -2197 14521
rect -2486 14453 -2197 14465
rect -3026 14328 -2737 14346
rect -3026 14272 -3015 14328
rect -2959 14272 -2911 14328
rect -2855 14272 -2807 14328
rect -2751 14272 -2737 14328
rect -3026 14224 -2737 14272
rect -3026 14168 -3015 14224
rect -2959 14168 -2911 14224
rect -2855 14168 -2807 14224
rect -2751 14168 -2737 14224
rect -3026 14120 -2737 14168
rect -3026 14064 -3015 14120
rect -2959 14064 -2911 14120
rect -2855 14064 -2807 14120
rect -2751 14064 -2737 14120
rect -3026 14052 -2737 14064
rect -3012 12406 -2747 14052
rect -3012 12388 -2714 12406
rect -3012 12332 -2992 12388
rect -2936 12332 -2888 12388
rect -2832 12332 -2784 12388
rect -2728 12332 -2714 12388
rect -3012 12284 -2714 12332
rect -3012 12228 -2992 12284
rect -2936 12228 -2888 12284
rect -2832 12228 -2784 12284
rect -2728 12228 -2714 12284
rect -3012 12180 -2714 12228
rect -3012 12124 -2992 12180
rect -2936 12124 -2888 12180
rect -2832 12124 -2784 12180
rect -2728 12124 -2714 12180
rect -3012 12112 -2714 12124
rect -3012 12094 -2747 12112
rect -2981 9083 -2692 9101
rect -2981 9027 -2970 9083
rect -2914 9027 -2866 9083
rect -2810 9027 -2762 9083
rect -2706 9027 -2692 9083
rect -2981 8979 -2692 9027
rect -2981 8923 -2970 8979
rect -2914 8923 -2866 8979
rect -2810 8923 -2762 8979
rect -2706 8923 -2692 8979
rect -2981 8875 -2692 8923
rect -2981 8819 -2970 8875
rect -2914 8819 -2866 8875
rect -2810 8819 -2762 8875
rect -2706 8819 -2692 8875
rect -2981 8807 -2692 8819
rect -3580 -2604 -3269 -2586
rect -3580 -2660 -3569 -2604
rect -3513 -2660 -3465 -2604
rect -3409 -2660 -3361 -2604
rect -3305 -2660 -3269 -2604
rect -3580 -2708 -3269 -2660
rect -3580 -2764 -3569 -2708
rect -3513 -2764 -3465 -2708
rect -3409 -2764 -3361 -2708
rect -3305 -2764 -3269 -2708
rect -3580 -2812 -3269 -2764
rect -3580 -2868 -3569 -2812
rect -3513 -2868 -3465 -2812
rect -3409 -2868 -3361 -2812
rect -3305 -2868 -3269 -2812
rect -3580 -2880 -3269 -2868
rect -3527 -2908 -3269 -2880
rect -5147 -4702 -4338 -4678
rect -5147 -4757 -5124 -4702
rect -5850 -4785 -5124 -4757
rect -5041 -4785 -4954 -4702
rect -4871 -4785 -4784 -4702
rect -4701 -4785 -4614 -4702
rect -4531 -4785 -4444 -4702
rect -4361 -4785 -4338 -4702
rect -5850 -4872 -4338 -4785
rect -5850 -4955 -5124 -4872
rect -5041 -4955 -4954 -4872
rect -4871 -4955 -4784 -4872
rect -4701 -4955 -4614 -4872
rect -4531 -4955 -4444 -4872
rect -4361 -4955 -4338 -4872
rect -5850 -5042 -4338 -4955
rect -5850 -5125 -5124 -5042
rect -5041 -5125 -4954 -5042
rect -4871 -5125 -4784 -5042
rect -4701 -5125 -4614 -5042
rect -4531 -5125 -4444 -5042
rect -4361 -5125 -4338 -5042
rect -5850 -5212 -4338 -5125
rect -5850 -5295 -5124 -5212
rect -5041 -5295 -4954 -5212
rect -4871 -5295 -4784 -5212
rect -4701 -5295 -4614 -5212
rect -4531 -5295 -4444 -5212
rect -4361 -5295 -4338 -5212
rect -5850 -5382 -4338 -5295
rect -5850 -5424 -5124 -5382
rect -5147 -5465 -5124 -5424
rect -5041 -5465 -4954 -5382
rect -4871 -5465 -4784 -5382
rect -4701 -5465 -4614 -5382
rect -4531 -5465 -4444 -5382
rect -4361 -5465 -4338 -5382
rect -5147 -5489 -4338 -5465
rect -5122 -7571 -4313 -7547
rect -5122 -7626 -5099 -7571
rect -5825 -7654 -5099 -7626
rect -5016 -7654 -4929 -7571
rect -4846 -7654 -4759 -7571
rect -4676 -7654 -4589 -7571
rect -4506 -7654 -4419 -7571
rect -4336 -7654 -4313 -7571
rect -5825 -7741 -4313 -7654
rect -5825 -7824 -5099 -7741
rect -5016 -7824 -4929 -7741
rect -4846 -7824 -4759 -7741
rect -4676 -7824 -4589 -7741
rect -4506 -7824 -4419 -7741
rect -4336 -7824 -4313 -7741
rect -5825 -7911 -4313 -7824
rect -5825 -7994 -5099 -7911
rect -5016 -7994 -4929 -7911
rect -4846 -7994 -4759 -7911
rect -4676 -7994 -4589 -7911
rect -4506 -7994 -4419 -7911
rect -4336 -7994 -4313 -7911
rect -5825 -8081 -4313 -7994
rect -5825 -8164 -5099 -8081
rect -5016 -8164 -4929 -8081
rect -4846 -8164 -4759 -8081
rect -4676 -8164 -4589 -8081
rect -4506 -8164 -4419 -8081
rect -4336 -8164 -4313 -8081
rect -5825 -8251 -4313 -8164
rect -5825 -8293 -5099 -8251
rect -5122 -8334 -5099 -8293
rect -5016 -8334 -4929 -8251
rect -4846 -8334 -4759 -8251
rect -4676 -8334 -4589 -8251
rect -4506 -8334 -4419 -8251
rect -4336 -8334 -4313 -8251
rect -5122 -8358 -4313 -8334
rect -2976 -9064 -2718 8807
rect -2459 4968 -2201 14453
rect -1051 13919 -762 13937
rect -1051 13863 -1040 13919
rect -984 13863 -936 13919
rect -880 13863 -832 13919
rect -776 13863 -762 13919
rect -1051 13815 -762 13863
rect -1051 13759 -1040 13815
rect -984 13759 -936 13815
rect -880 13759 -832 13815
rect -776 13759 -762 13815
rect -1051 13711 -762 13759
rect -1051 13655 -1040 13711
rect -984 13655 -936 13711
rect -880 13655 -832 13711
rect -776 13655 -762 13711
rect -1051 13643 -762 13655
rect -1430 13383 -1211 13399
rect -1455 13365 -1166 13383
rect -1455 13309 -1444 13365
rect -1388 13309 -1340 13365
rect -1284 13309 -1236 13365
rect -1180 13309 -1166 13365
rect -1455 13261 -1166 13309
rect -1455 13205 -1444 13261
rect -1388 13205 -1340 13261
rect -1284 13205 -1236 13261
rect -1180 13205 -1166 13261
rect -1455 13157 -1166 13205
rect -1455 13101 -1444 13157
rect -1388 13101 -1340 13157
rect -1284 13101 -1236 13157
rect -1180 13101 -1166 13157
rect -1455 13089 -1166 13101
rect -1953 11852 -1695 11853
rect -1968 11834 -1679 11852
rect -1968 11778 -1957 11834
rect -1901 11778 -1853 11834
rect -1797 11778 -1749 11834
rect -1693 11778 -1679 11834
rect -1968 11730 -1679 11778
rect -1968 11674 -1957 11730
rect -1901 11674 -1853 11730
rect -1797 11674 -1749 11730
rect -1693 11674 -1679 11730
rect -1968 11626 -1679 11674
rect -1968 11570 -1957 11626
rect -1901 11570 -1853 11626
rect -1797 11570 -1749 11626
rect -1693 11570 -1679 11626
rect -1968 11558 -1679 11570
rect -2481 4950 -2192 4968
rect -2481 4894 -2470 4950
rect -2414 4894 -2366 4950
rect -2310 4894 -2262 4950
rect -2206 4894 -2192 4950
rect -2481 4846 -2192 4894
rect -2481 4790 -2470 4846
rect -2414 4790 -2366 4846
rect -2310 4790 -2262 4846
rect -2206 4790 -2192 4846
rect -2481 4742 -2192 4790
rect -2481 4686 -2470 4742
rect -2414 4686 -2366 4742
rect -2310 4686 -2262 4742
rect -2206 4686 -2192 4742
rect -2481 4674 -2192 4686
rect -2459 4622 -2201 4674
rect -2466 1074 -2208 1102
rect -2481 1056 -2192 1074
rect -2481 1000 -2470 1056
rect -2414 1000 -2366 1056
rect -2310 1000 -2262 1056
rect -2206 1000 -2192 1056
rect -2481 952 -2192 1000
rect -2481 896 -2470 952
rect -2414 896 -2366 952
rect -2310 896 -2262 952
rect -2206 896 -2192 952
rect -2481 848 -2192 896
rect -2481 792 -2470 848
rect -2414 792 -2366 848
rect -2310 792 -2262 848
rect -2206 792 -2192 848
rect -2481 780 -2192 792
rect -2466 -7858 -2208 780
rect -1953 -1879 -1695 11558
rect -1977 -1897 -1688 -1879
rect -1977 -1953 -1966 -1897
rect -1910 -1953 -1862 -1897
rect -1806 -1953 -1758 -1897
rect -1702 -1953 -1688 -1897
rect -1977 -2001 -1688 -1953
rect -1977 -2057 -1966 -2001
rect -1910 -2057 -1862 -2001
rect -1806 -2057 -1758 -2001
rect -1702 -2057 -1688 -2001
rect -1977 -2105 -1688 -2057
rect -1977 -2161 -1966 -2105
rect -1910 -2161 -1862 -2105
rect -1806 -2161 -1758 -2105
rect -1702 -2161 -1688 -2105
rect -1977 -2173 -1688 -2161
rect -1914 -3063 -1625 -3045
rect -1914 -3119 -1903 -3063
rect -1847 -3119 -1799 -3063
rect -1743 -3119 -1695 -3063
rect -1639 -3119 -1625 -3063
rect -1914 -3167 -1625 -3119
rect -1914 -3223 -1903 -3167
rect -1847 -3223 -1799 -3167
rect -1743 -3223 -1695 -3167
rect -1639 -3223 -1625 -3167
rect -1914 -3271 -1625 -3223
rect -1914 -3327 -1903 -3271
rect -1847 -3327 -1799 -3271
rect -1743 -3327 -1695 -3271
rect -1639 -3327 -1625 -3271
rect -1914 -3339 -1625 -3327
rect -2504 -7876 -2208 -7858
rect -2504 -7932 -2493 -7876
rect -2437 -7932 -2389 -7876
rect -2333 -7932 -2285 -7876
rect -2229 -7932 -2208 -7876
rect -2504 -7980 -2208 -7932
rect -2504 -8036 -2493 -7980
rect -2437 -8036 -2389 -7980
rect -2333 -8036 -2285 -7980
rect -2229 -8036 -2208 -7980
rect -2504 -8084 -2208 -8036
rect -2504 -8140 -2493 -8084
rect -2437 -8140 -2389 -8084
rect -2333 -8140 -2285 -8084
rect -2229 -8140 -2208 -8084
rect -2504 -8152 -2208 -8140
rect -2466 -8187 -2208 -8152
rect -2994 -9082 -2705 -9064
rect -2994 -9138 -2983 -9082
rect -2927 -9138 -2879 -9082
rect -2823 -9138 -2775 -9082
rect -2719 -9138 -2705 -9082
rect -2994 -9186 -2705 -9138
rect -2994 -9242 -2983 -9186
rect -2927 -9242 -2879 -9186
rect -2823 -9242 -2775 -9186
rect -2719 -9242 -2705 -9186
rect -2994 -9290 -2705 -9242
rect -2994 -9346 -2983 -9290
rect -2927 -9346 -2879 -9290
rect -2823 -9346 -2775 -9290
rect -2719 -9346 -2705 -9290
rect -2994 -9358 -2705 -9346
rect -2976 -9369 -2718 -9358
rect -5099 -9675 -4290 -9651
rect -5099 -9730 -5076 -9675
rect -5802 -9758 -5076 -9730
rect -4993 -9758 -4906 -9675
rect -4823 -9758 -4736 -9675
rect -4653 -9758 -4566 -9675
rect -4483 -9758 -4396 -9675
rect -4313 -9758 -4290 -9675
rect -5802 -9845 -4290 -9758
rect -5802 -9928 -5076 -9845
rect -4993 -9928 -4906 -9845
rect -4823 -9928 -4736 -9845
rect -4653 -9928 -4566 -9845
rect -4483 -9928 -4396 -9845
rect -4313 -9928 -4290 -9845
rect -5802 -10015 -4290 -9928
rect -5802 -10098 -5076 -10015
rect -4993 -10098 -4906 -10015
rect -4823 -10098 -4736 -10015
rect -4653 -10098 -4566 -10015
rect -4483 -10098 -4396 -10015
rect -4313 -10098 -4290 -10015
rect -5802 -10185 -4290 -10098
rect -5802 -10268 -5076 -10185
rect -4993 -10268 -4906 -10185
rect -4823 -10268 -4736 -10185
rect -4653 -10268 -4566 -10185
rect -4483 -10268 -4396 -10185
rect -4313 -10268 -4290 -10185
rect -5802 -10355 -4290 -10268
rect -5802 -10397 -5076 -10355
rect -5099 -10438 -5076 -10397
rect -4993 -10438 -4906 -10355
rect -4823 -10438 -4736 -10355
rect -4653 -10438 -4566 -10355
rect -4483 -10438 -4396 -10355
rect -4313 -10438 -4290 -10355
rect -5099 -10462 -4290 -10438
rect -5076 -11849 -4267 -11825
rect -5076 -11904 -5053 -11849
rect -5779 -11932 -5053 -11904
rect -4970 -11932 -4883 -11849
rect -4800 -11932 -4713 -11849
rect -4630 -11932 -4543 -11849
rect -4460 -11932 -4373 -11849
rect -4290 -11932 -4267 -11849
rect -5779 -12019 -4267 -11932
rect -5779 -12102 -5053 -12019
rect -4970 -12102 -4883 -12019
rect -4800 -12102 -4713 -12019
rect -4630 -12102 -4543 -12019
rect -4460 -12102 -4373 -12019
rect -4290 -12102 -4267 -12019
rect -5779 -12189 -4267 -12102
rect -1878 -12126 -1659 -3339
rect -5779 -12272 -5053 -12189
rect -4970 -12272 -4883 -12189
rect -4800 -12272 -4713 -12189
rect -4630 -12272 -4543 -12189
rect -4460 -12272 -4373 -12189
rect -4290 -12272 -4267 -12189
rect -5779 -12359 -4267 -12272
rect -5779 -12442 -5053 -12359
rect -4970 -12442 -4883 -12359
rect -4800 -12442 -4713 -12359
rect -4630 -12442 -4543 -12359
rect -4460 -12442 -4373 -12359
rect -4290 -12442 -4267 -12359
rect -1936 -12144 -1647 -12126
rect -1936 -12200 -1925 -12144
rect -1869 -12200 -1821 -12144
rect -1765 -12200 -1717 -12144
rect -1661 -12200 -1647 -12144
rect -1936 -12248 -1647 -12200
rect -1936 -12304 -1925 -12248
rect -1869 -12304 -1821 -12248
rect -1765 -12304 -1717 -12248
rect -1661 -12304 -1647 -12248
rect -1936 -12352 -1647 -12304
rect -1936 -12408 -1925 -12352
rect -1869 -12408 -1821 -12352
rect -1765 -12408 -1717 -12352
rect -1661 -12408 -1647 -12352
rect -1936 -12420 -1647 -12408
rect -5779 -12529 -4267 -12442
rect -5779 -12571 -5053 -12529
rect -5076 -12612 -5053 -12571
rect -4970 -12612 -4883 -12529
rect -4800 -12612 -4713 -12529
rect -4630 -12612 -4543 -12529
rect -4460 -12612 -4373 -12529
rect -4290 -12612 -4267 -12529
rect -5076 -12636 -4267 -12612
rect -5122 -13653 -4313 -13629
rect -5122 -13708 -5099 -13653
rect -5825 -13736 -5099 -13708
rect -5016 -13736 -4929 -13653
rect -4846 -13736 -4759 -13653
rect -4676 -13736 -4589 -13653
rect -4506 -13736 -4419 -13653
rect -4336 -13736 -4313 -13653
rect -5825 -13823 -4313 -13736
rect -5825 -13906 -5099 -13823
rect -5016 -13906 -4929 -13823
rect -4846 -13906 -4759 -13823
rect -4676 -13906 -4589 -13823
rect -4506 -13906 -4419 -13823
rect -4336 -13906 -4313 -13823
rect -5825 -13993 -4313 -13906
rect -1430 -13931 -1211 13089
rect -5825 -14076 -5099 -13993
rect -5016 -14076 -4929 -13993
rect -4846 -14076 -4759 -13993
rect -4676 -14076 -4589 -13993
rect -4506 -14076 -4419 -13993
rect -4336 -14076 -4313 -13993
rect -5825 -14163 -4313 -14076
rect -5825 -14246 -5099 -14163
rect -5016 -14246 -4929 -14163
rect -4846 -14246 -4759 -14163
rect -4676 -14246 -4589 -14163
rect -4506 -14246 -4419 -14163
rect -4336 -14246 -4313 -14163
rect -1482 -13949 -1193 -13931
rect -1482 -14005 -1471 -13949
rect -1415 -14005 -1367 -13949
rect -1311 -14005 -1263 -13949
rect -1207 -14005 -1193 -13949
rect -1482 -14053 -1193 -14005
rect -1482 -14109 -1471 -14053
rect -1415 -14109 -1367 -14053
rect -1311 -14109 -1263 -14053
rect -1207 -14109 -1193 -14053
rect -1482 -14157 -1193 -14109
rect -1482 -14213 -1471 -14157
rect -1415 -14213 -1367 -14157
rect -1311 -14213 -1263 -14157
rect -1207 -14213 -1193 -14157
rect -1482 -14225 -1193 -14213
rect -5825 -14333 -4313 -14246
rect -5825 -14375 -5099 -14333
rect -5122 -14416 -5099 -14375
rect -5016 -14416 -4929 -14333
rect -4846 -14416 -4759 -14333
rect -4676 -14416 -4589 -14333
rect -4506 -14416 -4419 -14333
rect -4336 -14416 -4313 -14333
rect -5122 -14440 -4313 -14416
rect -5076 -15425 -4267 -15401
rect -5076 -15480 -5053 -15425
rect -5779 -15508 -5053 -15480
rect -4970 -15508 -4883 -15425
rect -4800 -15508 -4713 -15425
rect -4630 -15508 -4543 -15425
rect -4460 -15508 -4373 -15425
rect -4290 -15508 -4267 -15425
rect -5779 -15595 -4267 -15508
rect -5779 -15678 -5053 -15595
rect -4970 -15678 -4883 -15595
rect -4800 -15678 -4713 -15595
rect -4630 -15678 -4543 -15595
rect -4460 -15678 -4373 -15595
rect -4290 -15678 -4267 -15595
rect -5779 -15765 -4267 -15678
rect -5779 -15848 -5053 -15765
rect -4970 -15848 -4883 -15765
rect -4800 -15848 -4713 -15765
rect -4630 -15848 -4543 -15765
rect -4460 -15848 -4373 -15765
rect -4290 -15848 -4267 -15765
rect -5779 -15935 -4267 -15848
rect -5779 -16018 -5053 -15935
rect -4970 -16018 -4883 -15935
rect -4800 -16018 -4713 -15935
rect -4630 -16018 -4543 -15935
rect -4460 -16018 -4373 -15935
rect -4290 -16018 -4267 -15935
rect -5779 -16105 -4267 -16018
rect -5779 -16147 -5053 -16105
rect -5076 -16188 -5053 -16147
rect -4970 -16188 -4883 -16105
rect -4800 -16188 -4713 -16105
rect -4630 -16188 -4543 -16105
rect -4460 -16188 -4373 -16105
rect -4290 -16188 -4267 -16105
rect -5076 -16212 -4267 -16188
rect -5122 -17229 -4313 -17205
rect -5122 -17284 -5099 -17229
rect -5825 -17312 -5099 -17284
rect -5016 -17312 -4929 -17229
rect -4846 -17312 -4759 -17229
rect -4676 -17312 -4589 -17229
rect -4506 -17312 -4419 -17229
rect -4336 -17312 -4313 -17229
rect -5825 -17399 -4313 -17312
rect -5825 -17482 -5099 -17399
rect -5016 -17482 -4929 -17399
rect -4846 -17482 -4759 -17399
rect -4676 -17482 -4589 -17399
rect -4506 -17482 -4419 -17399
rect -4336 -17482 -4313 -17399
rect -5825 -17569 -4313 -17482
rect -1020 -17506 -802 13643
rect -583 -8236 -365 15505
rect -172 15352 117 15370
rect -172 15296 -161 15352
rect -105 15296 -57 15352
rect -1 15296 47 15352
rect 103 15296 117 15352
rect -172 15248 117 15296
rect -172 15192 -161 15248
rect -105 15192 -57 15248
rect -1 15192 47 15248
rect 103 15192 117 15248
rect -172 15144 117 15192
rect -172 15088 -161 15144
rect -105 15088 -57 15144
rect -1 15088 47 15144
rect 103 15088 117 15144
rect -172 15076 117 15088
rect -157 8398 61 15076
rect 23334 12875 23628 12889
rect 23334 12787 23348 12875
rect 23435 12787 23528 12875
rect 23615 12787 23628 12875
rect 23334 12695 23628 12787
rect 23334 12607 23348 12695
rect 23435 12607 23528 12695
rect 23615 12607 23628 12695
rect 23334 12593 23628 12607
rect 516 11839 805 11857
rect 516 11783 527 11839
rect 583 11783 631 11839
rect 687 11783 735 11839
rect 791 11783 805 11839
rect 516 11735 805 11783
rect 516 11679 527 11735
rect 583 11679 631 11735
rect 687 11679 735 11735
rect 791 11679 805 11735
rect 516 11631 805 11679
rect 516 11575 527 11631
rect 583 11575 631 11631
rect 687 11575 735 11631
rect 791 11575 805 11631
rect 516 11563 805 11575
rect 15882 10631 15981 10640
rect 15882 10624 16625 10631
rect 15882 10558 15899 10624
rect 15966 10609 16625 10624
rect 15966 10558 16529 10609
rect 15882 10552 16529 10558
rect 15882 10542 15981 10552
rect 16512 10543 16529 10552
rect 16596 10552 16625 10609
rect 16596 10543 16611 10552
rect 16512 10527 16611 10543
rect 18781 9293 19303 9352
rect 18781 9210 18836 9293
rect 18919 9210 19006 9293
rect 19089 9210 19176 9293
rect 19259 9210 19303 9293
rect 18781 9123 19303 9210
rect 18781 9040 18836 9123
rect 18919 9040 19006 9123
rect 19089 9040 19176 9123
rect 19259 9040 19303 9123
rect 18781 8953 19303 9040
rect 18781 8870 18836 8953
rect 18919 8870 19006 8953
rect 19089 8870 19176 8953
rect 19259 8870 19303 8953
rect 18781 8714 19303 8870
rect 18781 8631 18838 8714
rect 18921 8631 19008 8714
rect 19091 8631 19178 8714
rect 19261 8631 19303 8714
rect 18781 8544 19303 8631
rect 18781 8461 18838 8544
rect 18921 8461 19008 8544
rect 19091 8461 19178 8544
rect 19261 8461 19303 8544
rect -157 8289 1070 8398
rect 18781 8374 19303 8461
rect 15870 8293 15969 8304
rect 17030 8293 17129 8295
rect -157 8196 61 8289
rect 15870 8288 17129 8293
rect 15870 8222 15887 8288
rect 15954 8279 17129 8288
rect 15954 8222 17047 8279
rect 15870 8214 17047 8222
rect 15870 8206 15969 8214
rect 17030 8213 17047 8214
rect 17114 8213 17129 8279
rect 18781 8291 18838 8374
rect 18921 8291 19008 8374
rect 19091 8291 19178 8374
rect 19261 8291 19303 8374
rect 18781 8226 19303 8291
rect 17030 8197 17129 8213
rect 15873 7213 15972 7223
rect 17582 7213 17681 7223
rect 15873 7207 17681 7213
rect 15873 7141 15890 7207
rect 15957 7141 17599 7207
rect 17666 7141 17681 7207
rect 15873 7132 17681 7141
rect 15873 7125 15972 7132
rect 17582 7125 17681 7132
rect 603 6787 892 6805
rect 603 6731 614 6787
rect 670 6731 718 6787
rect 774 6731 822 6787
rect 878 6731 892 6787
rect 603 6683 892 6731
rect 603 6627 614 6683
rect 670 6627 718 6683
rect 774 6627 822 6683
rect 878 6627 892 6683
rect 603 6579 892 6627
rect 603 6523 614 6579
rect 670 6523 718 6579
rect 774 6523 822 6579
rect 878 6523 892 6579
rect 603 6511 892 6523
rect 19542 3771 19877 9769
rect 49563 7915 49888 15518
rect 52475 14621 52800 15546
rect 45166 7590 49888 7915
rect 50946 14296 52800 14621
rect 133279 14440 134136 14513
rect 133279 14439 134010 14440
rect 133279 14437 133676 14439
rect 133279 14349 133349 14437
rect 133436 14349 133529 14437
rect 133616 14351 133676 14437
rect 133763 14351 133856 14439
rect 133943 14352 134010 14439
rect 134097 14352 134136 14440
rect 133943 14351 134136 14352
rect 133616 14349 134136 14351
rect 50946 6616 51271 14296
rect 133279 14260 134136 14349
rect 133279 14259 134010 14260
rect 133279 14257 133676 14259
rect 133279 14169 133349 14257
rect 133436 14169 133529 14257
rect 133616 14171 133676 14257
rect 133763 14171 133856 14259
rect 133943 14172 134010 14259
rect 134097 14172 134136 14260
rect 133943 14171 134136 14172
rect 133616 14169 134136 14171
rect 133279 14047 134136 14169
rect 133279 14046 133992 14047
rect 133279 14044 133658 14046
rect 133279 13956 133331 14044
rect 133418 13956 133511 14044
rect 133598 13958 133658 14044
rect 133745 13958 133838 14046
rect 133925 13959 133992 14046
rect 134079 13959 134136 14047
rect 133925 13958 134136 13959
rect 133598 13956 134136 13958
rect 133279 13867 134136 13956
rect 133279 13866 133992 13867
rect 133279 13864 133658 13866
rect 133279 13776 133331 13864
rect 133418 13776 133511 13864
rect 133598 13778 133658 13864
rect 133745 13778 133838 13866
rect 133925 13779 133992 13866
rect 134079 13779 134136 13867
rect 133925 13778 134136 13779
rect 133598 13776 134136 13778
rect 133279 13698 134136 13776
rect 135785 14424 136642 14497
rect 135785 14423 136516 14424
rect 135785 14421 136182 14423
rect 135785 14333 135855 14421
rect 135942 14333 136035 14421
rect 136122 14335 136182 14421
rect 136269 14335 136362 14423
rect 136449 14336 136516 14423
rect 136603 14336 136642 14424
rect 136449 14335 136642 14336
rect 136122 14333 136642 14335
rect 135785 14244 136642 14333
rect 135785 14243 136516 14244
rect 135785 14241 136182 14243
rect 135785 14153 135855 14241
rect 135942 14153 136035 14241
rect 136122 14155 136182 14241
rect 136269 14155 136362 14243
rect 136449 14156 136516 14243
rect 136603 14156 136642 14244
rect 136449 14155 136642 14156
rect 136122 14153 136642 14155
rect 135785 14031 136642 14153
rect 135785 14030 136498 14031
rect 135785 14028 136164 14030
rect 135785 13940 135837 14028
rect 135924 13940 136017 14028
rect 136104 13942 136164 14028
rect 136251 13942 136344 14030
rect 136431 13943 136498 14030
rect 136585 13943 136642 14031
rect 136431 13942 136642 13943
rect 136104 13940 136642 13942
rect 135785 13851 136642 13940
rect 135785 13850 136498 13851
rect 135785 13848 136164 13850
rect 135785 13760 135837 13848
rect 135924 13760 136017 13848
rect 136104 13762 136164 13848
rect 136251 13762 136344 13850
rect 136431 13763 136498 13850
rect 136585 13763 136642 13851
rect 136431 13762 136642 13763
rect 136104 13760 136642 13762
rect 135785 13682 136642 13760
rect 138501 14443 139358 14516
rect 138501 14442 139232 14443
rect 138501 14440 138898 14442
rect 138501 14352 138571 14440
rect 138658 14352 138751 14440
rect 138838 14354 138898 14440
rect 138985 14354 139078 14442
rect 139165 14355 139232 14442
rect 139319 14355 139358 14443
rect 139165 14354 139358 14355
rect 138838 14352 139358 14354
rect 138501 14263 139358 14352
rect 138501 14262 139232 14263
rect 138501 14260 138898 14262
rect 138501 14172 138571 14260
rect 138658 14172 138751 14260
rect 138838 14174 138898 14260
rect 138985 14174 139078 14262
rect 139165 14175 139232 14262
rect 139319 14175 139358 14263
rect 139165 14174 139358 14175
rect 138838 14172 139358 14174
rect 138501 14050 139358 14172
rect 138501 14049 139214 14050
rect 138501 14047 138880 14049
rect 138501 13959 138553 14047
rect 138640 13959 138733 14047
rect 138820 13961 138880 14047
rect 138967 13961 139060 14049
rect 139147 13962 139214 14049
rect 139301 13962 139358 14050
rect 139147 13961 139358 13962
rect 138820 13959 139358 13961
rect 138501 13870 139358 13959
rect 138501 13869 139214 13870
rect 138501 13867 138880 13869
rect 138501 13779 138553 13867
rect 138640 13779 138733 13867
rect 138820 13781 138880 13867
rect 138967 13781 139060 13869
rect 139147 13782 139214 13869
rect 139301 13782 139358 13870
rect 139147 13781 139358 13782
rect 138820 13779 139358 13781
rect 138501 13701 139358 13779
rect 15138 3436 19877 3771
rect 46665 6291 51271 6616
rect 150298 6671 151141 6731
rect 150298 6670 151003 6671
rect 150298 6668 150669 6670
rect 150298 6580 150342 6668
rect 150429 6580 150522 6668
rect 150609 6582 150669 6668
rect 150756 6582 150849 6670
rect 150936 6583 151003 6670
rect 151090 6583 151141 6671
rect 150936 6582 151141 6583
rect 150609 6580 151141 6582
rect 150298 6491 151141 6580
rect 150298 6490 151003 6491
rect 150298 6488 150669 6490
rect 150298 6400 150342 6488
rect 150429 6400 150522 6488
rect 150609 6402 150669 6488
rect 150756 6402 150849 6490
rect 150936 6403 151003 6490
rect 151090 6403 151141 6491
rect 150936 6402 151141 6403
rect 150609 6400 151141 6402
rect 150298 6356 151141 6400
rect -163 2470 95 2479
rect -176 2452 113 2470
rect -176 2396 -165 2452
rect -109 2396 -61 2452
rect -5 2396 43 2452
rect 99 2396 113 2452
rect -176 2348 113 2396
rect -176 2292 -165 2348
rect -109 2292 -61 2348
rect -5 2292 43 2348
rect 99 2292 113 2348
rect -176 2244 113 2292
rect -176 2188 -165 2244
rect -109 2188 -61 2244
rect -5 2188 43 2244
rect 99 2188 113 2244
rect -176 2176 113 2188
rect -163 -2244 95 2176
rect 654 1039 943 1057
rect 654 983 665 1039
rect 721 983 769 1039
rect 825 983 873 1039
rect 929 983 943 1039
rect 654 935 943 983
rect 654 879 665 935
rect 721 879 769 935
rect 825 879 873 935
rect 929 879 943 935
rect 654 831 943 879
rect 654 775 665 831
rect 721 775 769 831
rect 825 775 873 831
rect 929 775 943 831
rect 654 763 943 775
rect 28005 680 28862 753
rect 28005 679 28736 680
rect 28005 677 28402 679
rect 28005 589 28075 677
rect 28162 589 28255 677
rect 28342 591 28402 677
rect 28489 591 28582 679
rect 28669 592 28736 679
rect 28823 592 28862 680
rect 28669 591 28862 592
rect 28342 589 28862 591
rect 28005 500 28862 589
rect 28005 499 28736 500
rect 28005 497 28402 499
rect 28005 409 28075 497
rect 28162 409 28255 497
rect 28342 411 28402 497
rect 28489 411 28582 499
rect 28669 412 28736 499
rect 28823 412 28862 500
rect 28669 411 28862 412
rect 28342 409 28862 411
rect 28005 287 28862 409
rect 28005 286 28718 287
rect 28005 284 28384 286
rect 28005 196 28057 284
rect 28144 196 28237 284
rect 28324 198 28384 284
rect 28471 198 28564 286
rect 28651 199 28718 286
rect 28805 199 28862 287
rect 28651 198 28862 199
rect 28324 196 28862 198
rect 28005 107 28862 196
rect 28005 106 28718 107
rect 28005 104 28384 106
rect 28005 16 28057 104
rect 28144 16 28237 104
rect 28324 18 28384 104
rect 28471 18 28564 106
rect 28651 19 28718 106
rect 28805 19 28862 107
rect 28651 18 28862 19
rect 28324 16 28862 18
rect 28005 -63 28862 16
rect 29817 727 30674 793
rect 29817 726 30542 727
rect 29817 724 30208 726
rect 29817 636 29881 724
rect 29968 636 30061 724
rect 30148 638 30208 724
rect 30295 638 30388 726
rect 30475 639 30542 726
rect 30629 639 30674 727
rect 30475 638 30674 639
rect 30148 636 30674 638
rect 29817 547 30674 636
rect 29817 546 30542 547
rect 29817 544 30208 546
rect 29817 456 29881 544
rect 29968 456 30061 544
rect 30148 458 30208 544
rect 30295 458 30388 546
rect 30475 459 30542 546
rect 30629 459 30674 547
rect 30475 458 30674 459
rect 30148 456 30674 458
rect 29817 339 30674 456
rect 29817 338 30548 339
rect 29817 336 30214 338
rect 29817 248 29887 336
rect 29974 248 30067 336
rect 30154 250 30214 336
rect 30301 250 30394 338
rect 30481 251 30548 338
rect 30635 251 30674 339
rect 30481 250 30674 251
rect 30154 248 30674 250
rect 29817 159 30674 248
rect 29817 158 30548 159
rect 29817 156 30214 158
rect 29817 68 29887 156
rect 29974 68 30067 156
rect 30154 70 30214 156
rect 30301 70 30394 158
rect 30481 71 30548 158
rect 30635 71 30674 159
rect 30481 70 30674 71
rect 30154 68 30674 70
rect 29817 -23 30674 68
rect 31572 727 32429 770
rect 31572 726 32279 727
rect 31572 724 31945 726
rect 31572 636 31618 724
rect 31705 636 31798 724
rect 31885 638 31945 724
rect 32032 638 32125 726
rect 32212 639 32279 726
rect 32366 639 32429 727
rect 32212 638 32429 639
rect 31885 636 32429 638
rect 31572 547 32429 636
rect 31572 546 32279 547
rect 31572 544 31945 546
rect 31572 456 31618 544
rect 31705 456 31798 544
rect 31885 458 31945 544
rect 32032 458 32125 546
rect 32212 459 32279 546
rect 32366 459 32429 547
rect 32212 458 32429 459
rect 31885 456 32429 458
rect 31572 339 32429 456
rect 31572 338 32291 339
rect 31572 336 31957 338
rect 31572 248 31630 336
rect 31717 248 31810 336
rect 31897 250 31957 336
rect 32044 250 32137 338
rect 32224 251 32291 338
rect 32378 251 32429 339
rect 32224 250 32429 251
rect 31897 248 32429 250
rect 31572 159 32429 248
rect 31572 158 32291 159
rect 31572 156 31957 158
rect 31572 68 31630 156
rect 31717 68 31810 156
rect 31897 70 31957 156
rect 32044 70 32137 158
rect 32224 71 32291 158
rect 32378 71 32429 159
rect 32224 70 32429 71
rect 31897 68 32429 70
rect 31572 -46 32429 68
rect 23075 -2069 23369 -2055
rect 23075 -2157 23089 -2069
rect 23176 -2157 23269 -2069
rect 23356 -2157 23369 -2069
rect -163 -2262 126 -2244
rect -163 -2318 -152 -2262
rect -96 -2318 -48 -2262
rect 8 -2318 56 -2262
rect 112 -2318 126 -2262
rect -163 -2366 126 -2318
rect 23075 -2249 23369 -2157
rect 23075 -2337 23089 -2249
rect 23176 -2337 23269 -2249
rect 23356 -2337 23369 -2249
rect 23075 -2351 23369 -2337
rect -163 -2422 -152 -2366
rect -96 -2422 -48 -2366
rect 8 -2422 56 -2366
rect 112 -2422 126 -2366
rect -163 -2470 126 -2422
rect -163 -2526 -152 -2470
rect -96 -2526 -48 -2470
rect 8 -2526 56 -2470
rect 112 -2526 126 -2470
rect -163 -2538 126 -2526
rect 17 -2929 236 -2893
rect -68 -2947 236 -2929
rect -68 -3003 -57 -2947
rect -1 -3003 47 -2947
rect 103 -3003 151 -2947
rect 207 -3003 236 -2947
rect -68 -3051 236 -3003
rect -68 -3107 -57 -3051
rect -1 -3107 47 -3051
rect 103 -3107 151 -3051
rect 207 -3107 236 -3051
rect -68 -3155 236 -3107
rect -68 -3211 -57 -3155
rect -1 -3211 47 -3155
rect 103 -3211 151 -3155
rect 207 -3211 236 -3155
rect -68 -3223 236 -3211
rect -622 -8254 -333 -8236
rect -622 -8310 -611 -8254
rect -555 -8310 -507 -8254
rect -451 -8310 -403 -8254
rect -347 -8310 -333 -8254
rect -622 -8358 -333 -8310
rect -622 -8414 -611 -8358
rect -555 -8414 -507 -8358
rect -451 -8414 -403 -8358
rect -347 -8414 -333 -8358
rect -622 -8462 -333 -8414
rect -622 -8518 -611 -8462
rect -555 -8518 -507 -8462
rect -451 -8518 -403 -8462
rect -347 -8518 -333 -8462
rect -622 -8530 -333 -8518
rect 17 -15700 236 -3223
rect 720 -4976 1009 -4958
rect 720 -5032 731 -4976
rect 787 -5032 835 -4976
rect 891 -5032 939 -4976
rect 995 -5032 1009 -4976
rect 720 -5080 1009 -5032
rect 720 -5136 731 -5080
rect 787 -5136 835 -5080
rect 891 -5136 939 -5080
rect 995 -5136 1009 -5080
rect 720 -5184 1009 -5136
rect 720 -5240 731 -5184
rect 787 -5240 835 -5184
rect 891 -5240 939 -5184
rect 995 -5240 1009 -5184
rect 720 -5252 1009 -5240
rect 18093 -5810 18615 -5742
rect 18093 -5893 18142 -5810
rect 18225 -5893 18312 -5810
rect 18395 -5893 18482 -5810
rect 18565 -5893 18615 -5810
rect 18093 -5980 18615 -5893
rect 18093 -6063 18142 -5980
rect 18225 -6063 18312 -5980
rect 18395 -6063 18482 -5980
rect 18565 -6063 18615 -5980
rect 16024 -6136 16123 -6126
rect 16521 -6136 16620 -6126
rect 16024 -6142 16620 -6136
rect 16024 -6208 16041 -6142
rect 16108 -6208 16538 -6142
rect 16605 -6208 16620 -6142
rect 16024 -6215 16620 -6208
rect 16024 -6224 16123 -6215
rect 16521 -6224 16620 -6215
rect 18093 -6150 18615 -6063
rect 18093 -6233 18142 -6150
rect 18225 -6233 18312 -6150
rect 18395 -6233 18482 -6150
rect 18565 -6233 18615 -6150
rect 18093 -6392 18615 -6233
rect 18093 -6475 18151 -6392
rect 18234 -6475 18321 -6392
rect 18404 -6475 18491 -6392
rect 18574 -6475 18615 -6392
rect 18093 -6562 18615 -6475
rect 18093 -6645 18151 -6562
rect 18234 -6645 18321 -6562
rect 18404 -6645 18491 -6562
rect 18574 -6645 18615 -6562
rect 18093 -6732 18615 -6645
rect 18093 -6815 18151 -6732
rect 18234 -6815 18321 -6732
rect 18404 -6815 18491 -6732
rect 18574 -6815 18615 -6732
rect 18093 -6868 18615 -6815
rect 702 -8312 991 -8294
rect 702 -8368 713 -8312
rect 769 -8368 817 -8312
rect 873 -8368 921 -8312
rect 977 -8368 991 -8312
rect 702 -8416 991 -8368
rect 702 -8472 713 -8416
rect 769 -8472 817 -8416
rect 873 -8472 921 -8416
rect 977 -8472 991 -8416
rect 702 -8520 991 -8472
rect 702 -8576 713 -8520
rect 769 -8576 817 -8520
rect 873 -8576 921 -8520
rect 977 -8576 991 -8520
rect 16028 -8478 16127 -8468
rect 16996 -8478 17095 -8468
rect 16028 -8484 17095 -8478
rect 16028 -8550 16045 -8484
rect 16112 -8550 17013 -8484
rect 17080 -8550 17095 -8484
rect 16028 -8555 17095 -8550
rect 16028 -8566 16127 -8555
rect 16996 -8566 17095 -8555
rect 702 -8588 991 -8576
rect 778 -9073 1067 -9055
rect 778 -9129 789 -9073
rect 845 -9129 893 -9073
rect 949 -9129 997 -9073
rect 1053 -9085 1067 -9073
rect 1053 -9129 1100 -9085
rect 778 -9177 1100 -9129
rect 778 -9233 789 -9177
rect 845 -9233 893 -9177
rect 949 -9233 997 -9177
rect 1053 -9233 1100 -9177
rect 778 -9281 1100 -9233
rect 778 -9337 789 -9281
rect 845 -9337 893 -9281
rect 949 -9337 997 -9281
rect 1053 -9337 1100 -9281
rect 778 -9349 1100 -9337
rect 795 -10233 1100 -9349
rect 16041 -9555 16140 -9546
rect 17540 -9555 17639 -9546
rect 16041 -9562 17639 -9555
rect 16041 -9628 16058 -9562
rect 16125 -9628 17557 -9562
rect 17624 -9628 17639 -9562
rect 16041 -9635 17639 -9628
rect 16041 -9644 16140 -9635
rect 17540 -9644 17639 -9635
rect 1143 -10735 1432 -10717
rect 1143 -10791 1154 -10735
rect 1210 -10791 1258 -10735
rect 1314 -10791 1362 -10735
rect 1418 -10791 1432 -10735
rect 1143 -10839 1432 -10791
rect 1143 -10895 1154 -10839
rect 1210 -10895 1258 -10839
rect 1314 -10895 1362 -10839
rect 1418 -10895 1432 -10839
rect 1143 -10943 1432 -10895
rect 1143 -10999 1154 -10943
rect 1210 -10999 1258 -10943
rect 1314 -10999 1362 -10943
rect 1418 -10999 1432 -10943
rect 1143 -11011 1432 -10999
rect -77 -15718 236 -15700
rect -77 -15774 -66 -15718
rect -10 -15774 38 -15718
rect 94 -15774 142 -15718
rect 198 -15774 236 -15718
rect -77 -15822 236 -15774
rect -77 -15878 -66 -15822
rect -10 -15878 38 -15822
rect 94 -15878 142 -15822
rect 198 -15878 236 -15822
rect -77 -15926 236 -15878
rect -77 -15982 -66 -15926
rect -10 -15982 38 -15926
rect 94 -15982 142 -15926
rect 198 -15982 236 -15926
rect 1182 -15975 1403 -11011
rect 19264 -12999 19599 -5417
rect 46665 -5426 46990 6291
rect 80879 6043 81977 6073
rect 75608 5997 76748 6038
rect 75608 5996 76309 5997
rect 75608 5994 75975 5996
rect 75608 5906 75648 5994
rect 75735 5906 75828 5994
rect 75915 5908 75975 5994
rect 76062 5908 76155 5996
rect 76242 5909 76309 5996
rect 76396 5996 76748 5997
rect 76396 5909 76449 5996
rect 76242 5908 76449 5909
rect 76536 5994 76748 5996
rect 76536 5908 76590 5994
rect 75915 5906 76590 5908
rect 76677 5906 76748 5994
rect 75608 5817 76748 5906
rect 75608 5816 76309 5817
rect 75608 5814 75975 5816
rect 75608 5726 75648 5814
rect 75735 5726 75828 5814
rect 75915 5728 75975 5814
rect 76062 5728 76155 5816
rect 76242 5729 76309 5816
rect 76396 5816 76748 5817
rect 76396 5729 76449 5816
rect 76242 5728 76449 5729
rect 76536 5814 76748 5816
rect 76536 5728 76590 5814
rect 75915 5726 76590 5728
rect 76677 5726 76748 5814
rect 75608 5683 76748 5726
rect 80879 6033 81982 6043
rect 80879 6032 81734 6033
rect 80879 6031 81580 6032
rect 80879 6029 81246 6031
rect 80879 5941 80919 6029
rect 81006 5941 81099 6029
rect 81186 5943 81246 6029
rect 81333 5943 81426 6031
rect 81513 5944 81580 6031
rect 81667 5945 81734 6032
rect 81821 6031 81982 6033
rect 81821 5945 81882 6031
rect 81667 5944 81882 5945
rect 81513 5943 81882 5944
rect 81969 5943 81982 6031
rect 81186 5941 81982 5943
rect 80879 5853 81982 5941
rect 80879 5852 81734 5853
rect 80879 5851 81580 5852
rect 80879 5849 81246 5851
rect 80879 5761 80919 5849
rect 81006 5761 81099 5849
rect 81186 5763 81246 5849
rect 81333 5763 81426 5851
rect 81513 5764 81580 5851
rect 81667 5765 81734 5852
rect 81821 5851 81982 5853
rect 81821 5765 81882 5851
rect 81667 5764 81882 5765
rect 81513 5763 81882 5764
rect 81969 5763 81982 5851
rect 81186 5761 81982 5763
rect 80879 5746 81982 5761
rect 80879 5718 81977 5746
rect 126212 4902 126506 4916
rect 126212 4901 126226 4902
rect 115729 4814 126226 4901
rect 126313 4814 126406 4902
rect 126493 4814 126506 4902
rect 115729 4722 126506 4814
rect 115729 4634 126226 4722
rect 126313 4634 126406 4722
rect 126493 4634 126506 4722
rect 56833 4217 57127 4231
rect 56833 4129 56847 4217
rect 56934 4129 57027 4217
rect 57114 4129 57127 4217
rect 56833 4037 57127 4129
rect 56833 3949 56847 4037
rect 56934 3949 57027 4037
rect 57114 3949 57127 4037
rect 56833 3935 57127 3949
rect 115054 3958 115376 3977
rect 114442 3912 114764 3930
rect 113812 3862 114134 3879
rect 113812 3774 113837 3862
rect 113924 3774 114017 3862
rect 114104 3774 114134 3862
rect 113812 3682 114134 3774
rect 113812 3594 113837 3682
rect 113924 3594 114017 3682
rect 114104 3594 114134 3682
rect 113812 3521 114134 3594
rect 113812 3433 113839 3521
rect 113926 3433 114019 3521
rect 114106 3433 114134 3521
rect 113812 3341 114134 3433
rect 113812 3253 113839 3341
rect 113926 3253 114019 3341
rect 114106 3253 114134 3341
rect 114442 3824 114475 3912
rect 114562 3824 114655 3912
rect 114742 3824 114764 3912
rect 114442 3732 114764 3824
rect 114442 3644 114475 3732
rect 114562 3644 114655 3732
rect 114742 3644 114764 3732
rect 114442 3569 114764 3644
rect 114442 3481 114473 3569
rect 114560 3481 114653 3569
rect 114740 3481 114764 3569
rect 114442 3389 114764 3481
rect 114442 3301 114473 3389
rect 114560 3301 114653 3389
rect 114740 3301 114764 3389
rect 115054 3870 115082 3958
rect 115169 3870 115262 3958
rect 115349 3870 115376 3958
rect 115729 3955 115996 4634
rect 126212 4620 126506 4634
rect 115054 3778 115376 3870
rect 115054 3690 115082 3778
rect 115169 3690 115262 3778
rect 115349 3690 115376 3778
rect 115054 3618 115376 3690
rect 115054 3530 115082 3618
rect 115169 3530 115262 3618
rect 115349 3530 115376 3618
rect 115054 3438 115376 3530
rect 115054 3350 115082 3438
rect 115169 3350 115262 3438
rect 115349 3350 115376 3438
rect 115054 3329 115376 3350
rect 115708 3940 116010 3955
rect 115708 3852 115729 3940
rect 115816 3852 115909 3940
rect 115996 3852 116010 3940
rect 115708 3760 116010 3852
rect 115708 3672 115729 3760
rect 115816 3672 115909 3760
rect 115996 3672 116010 3760
rect 115708 3623 116010 3672
rect 115708 3609 116012 3623
rect 115708 3521 115732 3609
rect 115819 3521 115912 3609
rect 115999 3521 116012 3609
rect 115708 3429 116012 3521
rect 115708 3341 115732 3429
rect 115819 3341 115912 3429
rect 115999 3341 116012 3429
rect 115708 3327 116012 3341
rect 115708 3317 116010 3327
rect 114442 3282 114764 3301
rect 113812 3231 114134 3253
rect 48377 764 50129 828
rect 48377 699 48410 764
rect 48475 699 48535 764
rect 48600 699 48660 764
rect 48725 699 50129 764
rect 48377 602 50129 699
rect 49903 -1391 50129 602
rect 120761 270 128097 447
rect 120761 268 127458 270
rect 120761 212 127143 268
rect 127199 212 127247 268
rect 127303 212 127351 268
rect 127407 214 127458 268
rect 127514 214 127562 270
rect 127618 214 127666 270
rect 127722 214 127773 270
rect 127829 214 127877 270
rect 127933 214 127981 270
rect 128037 214 128097 270
rect 127407 212 128097 214
rect 120761 166 128097 212
rect 120761 164 127458 166
rect 120761 108 127143 164
rect 127199 108 127247 164
rect 127303 108 127351 164
rect 127407 110 127458 164
rect 127514 110 127562 166
rect 127618 110 127666 166
rect 127722 110 127773 166
rect 127829 110 127877 166
rect 127933 110 127981 166
rect 128037 110 128097 166
rect 127407 108 128097 110
rect 120761 62 128097 108
rect 120761 60 127458 62
rect 120761 55 127143 60
rect 115912 4 127143 55
rect 127199 4 127247 60
rect 127303 4 127351 60
rect 127407 6 127458 60
rect 127514 6 127562 62
rect 127618 6 127666 62
rect 127722 6 127773 62
rect 127829 6 127877 62
rect 127933 6 127981 62
rect 128037 6 128097 62
rect 127407 4 128097 6
rect 115912 -123 128097 4
rect 115912 -125 116290 -123
rect 115912 -181 115975 -125
rect 116031 -181 116079 -125
rect 116135 -181 116183 -125
rect 116239 -179 116290 -125
rect 116346 -179 116394 -123
rect 116450 -179 116498 -123
rect 116554 -179 116605 -123
rect 116661 -179 116709 -123
rect 116765 -179 116813 -123
rect 116869 -179 128097 -123
rect 116239 -181 128097 -179
rect 115912 -227 128097 -181
rect 115912 -229 116290 -227
rect 115912 -285 115975 -229
rect 116031 -285 116079 -229
rect 116135 -285 116183 -229
rect 116239 -283 116290 -229
rect 116346 -283 116394 -227
rect 116450 -283 116498 -227
rect 116554 -283 116605 -227
rect 116661 -283 116709 -227
rect 116765 -283 116813 -227
rect 116869 -229 128097 -227
rect 116869 -283 121437 -229
rect 116239 -285 121437 -283
rect 115912 -331 121437 -285
rect 115912 -333 116290 -331
rect 115912 -389 115975 -333
rect 116031 -389 116079 -333
rect 116135 -389 116183 -333
rect 116239 -387 116290 -333
rect 116346 -387 116394 -331
rect 116450 -387 116498 -331
rect 116554 -387 116605 -331
rect 116661 -387 116709 -331
rect 116765 -387 116813 -331
rect 116869 -387 121437 -331
rect 116239 -389 121437 -387
rect 115912 -621 121437 -389
rect 123050 -588 134370 -551
rect 64609 -1280 64825 -1261
rect 64609 -1336 64643 -1280
rect 64699 -1336 64747 -1280
rect 64803 -1336 64825 -1280
rect 64609 -1384 64825 -1336
rect 64609 -1391 64643 -1384
rect 49903 -1440 64643 -1391
rect 64699 -1440 64747 -1384
rect 64803 -1440 64825 -1384
rect 49903 -1514 64825 -1440
rect 49903 -1570 64645 -1514
rect 64701 -1570 64749 -1514
rect 64805 -1570 64825 -1514
rect 49903 -1617 64825 -1570
rect 64609 -1618 64825 -1617
rect 64609 -1674 64645 -1618
rect 64701 -1674 64749 -1618
rect 64805 -1674 64825 -1618
rect 64609 -1703 64825 -1674
rect 68749 -1972 69427 -1550
rect 68749 -5239 69171 -1972
rect 86665 -2131 87681 -2092
rect 86665 -2219 86691 -2131
rect 86778 -2219 86871 -2131
rect 86958 -2219 87037 -2131
rect 87124 -2219 87217 -2131
rect 87304 -2134 87681 -2131
rect 87304 -2219 87390 -2134
rect 86665 -2222 87390 -2219
rect 87477 -2222 87570 -2134
rect 87657 -2222 87681 -2134
rect 86665 -2311 87681 -2222
rect 86665 -2399 86691 -2311
rect 86778 -2399 86871 -2311
rect 86958 -2399 87037 -2311
rect 87124 -2399 87217 -2311
rect 87304 -2314 87681 -2311
rect 87304 -2399 87390 -2314
rect 86665 -2402 87390 -2399
rect 87477 -2402 87570 -2314
rect 87657 -2402 87681 -2314
rect 86665 -2431 87681 -2402
rect 85602 -3282 117978 -3116
rect 85602 -3370 85749 -3282
rect 85836 -3370 85929 -3282
rect 86016 -3370 86095 -3282
rect 86182 -3370 86275 -3282
rect 86362 -3285 117978 -3282
rect 86362 -3370 86448 -3285
rect 85602 -3373 86448 -3370
rect 86535 -3373 86628 -3285
rect 86715 -3373 117978 -3285
rect 85602 -3462 117978 -3373
rect 85602 -3550 85749 -3462
rect 85836 -3550 85929 -3462
rect 86016 -3550 86095 -3462
rect 86182 -3550 86275 -3462
rect 86362 -3465 117978 -3462
rect 86362 -3550 86448 -3465
rect 85602 -3553 86448 -3550
rect 86535 -3553 86628 -3465
rect 86715 -3553 117978 -3465
rect 85602 -3718 117978 -3553
rect 68749 -5661 69427 -5239
rect 117376 -11604 117978 -3718
rect 120991 -3877 121340 -621
rect 123050 -644 133929 -588
rect 133985 -644 134033 -588
rect 134089 -591 134370 -588
rect 134089 -644 134165 -591
rect 123050 -647 134165 -644
rect 134221 -647 134269 -591
rect 134325 -647 134370 -591
rect 123050 -692 134370 -647
rect 123050 -748 133929 -692
rect 133985 -748 134033 -692
rect 134089 -695 134370 -692
rect 134089 -748 134165 -695
rect 123050 -751 134165 -748
rect 134221 -751 134269 -695
rect 134325 -751 134370 -695
rect 123050 -794 134370 -751
rect 123050 -3203 123293 -794
rect 122319 -3240 123293 -3203
rect 122319 -3307 122342 -3240
rect 122406 -3245 123293 -3240
rect 122406 -3307 122474 -3245
rect 122319 -3312 122474 -3307
rect 122538 -3312 123293 -3245
rect 122319 -3364 123293 -3312
rect 122319 -3365 122472 -3364
rect 122319 -3432 122347 -3365
rect 122411 -3431 122472 -3365
rect 122536 -3431 123293 -3364
rect 122411 -3432 123293 -3431
rect 122319 -3446 123293 -3432
rect 122319 -3466 122556 -3446
rect 120991 -3880 121167 -3877
rect 120991 -3946 121036 -3880
rect 121102 -3943 121167 -3880
rect 121233 -3943 121340 -3877
rect 121102 -3946 121340 -3943
rect 120991 -4009 121340 -3946
rect 120991 -4075 121035 -4009
rect 121101 -4075 121169 -4009
rect 121235 -4075 121340 -4009
rect 120991 -4137 121340 -4075
rect 120991 -4203 121032 -4137
rect 121098 -4203 121167 -4137
rect 121233 -4203 121340 -4137
rect 120991 -4290 121340 -4203
rect 121601 -7081 122617 -7042
rect 121601 -7169 121627 -7081
rect 121714 -7169 121807 -7081
rect 121894 -7169 121973 -7081
rect 122060 -7169 122153 -7081
rect 122240 -7084 122617 -7081
rect 122240 -7169 122326 -7084
rect 121601 -7172 122326 -7169
rect 122413 -7172 122506 -7084
rect 122593 -7172 122617 -7084
rect 121601 -7261 122617 -7172
rect 121601 -7349 121627 -7261
rect 121714 -7349 121807 -7261
rect 121894 -7349 121973 -7261
rect 122060 -7349 122153 -7261
rect 122240 -7264 122617 -7261
rect 122240 -7349 122326 -7264
rect 121601 -7352 122326 -7349
rect 122413 -7352 122506 -7264
rect 122593 -7352 122617 -7264
rect 121601 -7381 122617 -7352
rect 170266 -7085 171282 -7046
rect 170266 -7173 170292 -7085
rect 170379 -7173 170472 -7085
rect 170559 -7173 170638 -7085
rect 170725 -7173 170818 -7085
rect 170905 -7088 171282 -7085
rect 170905 -7173 170991 -7088
rect 170266 -7176 170991 -7173
rect 171078 -7176 171171 -7088
rect 171258 -7176 171282 -7088
rect 170266 -7265 171282 -7176
rect 170266 -7353 170292 -7265
rect 170379 -7353 170472 -7265
rect 170559 -7353 170638 -7265
rect 170725 -7353 170818 -7265
rect 170905 -7268 171282 -7265
rect 170905 -7353 170991 -7268
rect 170266 -7356 170991 -7353
rect 171078 -7356 171171 -7268
rect 171258 -7356 171282 -7268
rect 170266 -7385 171282 -7356
rect 170589 -11604 171132 -7385
rect 117376 -12175 171132 -11604
rect 15308 -13334 19599 -12999
rect 133309 -13430 134166 -13357
rect 133309 -13431 134040 -13430
rect 133309 -13433 133706 -13431
rect 133309 -13521 133379 -13433
rect 133466 -13521 133559 -13433
rect 133646 -13519 133706 -13433
rect 133793 -13519 133886 -13431
rect 133973 -13518 134040 -13431
rect 134127 -13518 134166 -13430
rect 133973 -13519 134166 -13518
rect 133646 -13521 134166 -13519
rect 133309 -13610 134166 -13521
rect 133309 -13611 134040 -13610
rect 133309 -13613 133706 -13611
rect 133309 -13701 133379 -13613
rect 133466 -13701 133559 -13613
rect 133646 -13699 133706 -13613
rect 133793 -13699 133886 -13611
rect 133973 -13698 134040 -13611
rect 134127 -13698 134166 -13610
rect 133973 -13699 134166 -13698
rect 133646 -13701 134166 -13699
rect 133309 -13823 134166 -13701
rect 133309 -13824 134022 -13823
rect 133309 -13826 133688 -13824
rect 133309 -13914 133361 -13826
rect 133448 -13914 133541 -13826
rect 133628 -13912 133688 -13826
rect 133775 -13912 133868 -13824
rect 133955 -13911 134022 -13824
rect 134109 -13911 134166 -13823
rect 133955 -13912 134166 -13911
rect 133628 -13914 134166 -13912
rect 133309 -14003 134166 -13914
rect 133309 -14004 134022 -14003
rect 133309 -14006 133688 -14004
rect 133309 -14094 133361 -14006
rect 133448 -14094 133541 -14006
rect 133628 -14092 133688 -14006
rect 133775 -14092 133868 -14004
rect 133955 -14091 134022 -14004
rect 134109 -14091 134166 -14003
rect 133955 -14092 134166 -14091
rect 133628 -14094 134166 -14092
rect 133309 -14172 134166 -14094
rect 135747 -13435 136604 -13362
rect 135747 -13436 136478 -13435
rect 135747 -13438 136144 -13436
rect 135747 -13526 135817 -13438
rect 135904 -13526 135997 -13438
rect 136084 -13524 136144 -13438
rect 136231 -13524 136324 -13436
rect 136411 -13523 136478 -13436
rect 136565 -13523 136604 -13435
rect 136411 -13524 136604 -13523
rect 136084 -13526 136604 -13524
rect 135747 -13615 136604 -13526
rect 135747 -13616 136478 -13615
rect 135747 -13618 136144 -13616
rect 135747 -13706 135817 -13618
rect 135904 -13706 135997 -13618
rect 136084 -13704 136144 -13618
rect 136231 -13704 136324 -13616
rect 136411 -13703 136478 -13616
rect 136565 -13703 136604 -13615
rect 136411 -13704 136604 -13703
rect 136084 -13706 136604 -13704
rect 135747 -13828 136604 -13706
rect 135747 -13829 136460 -13828
rect 135747 -13831 136126 -13829
rect 135747 -13919 135799 -13831
rect 135886 -13919 135979 -13831
rect 136066 -13917 136126 -13831
rect 136213 -13917 136306 -13829
rect 136393 -13916 136460 -13829
rect 136547 -13916 136604 -13828
rect 136393 -13917 136604 -13916
rect 136066 -13919 136604 -13917
rect 135747 -14008 136604 -13919
rect 135747 -14009 136460 -14008
rect 135747 -14011 136126 -14009
rect 135747 -14099 135799 -14011
rect 135886 -14099 135979 -14011
rect 136066 -14097 136126 -14011
rect 136213 -14097 136306 -14009
rect 136393 -14096 136460 -14009
rect 136547 -14096 136604 -14008
rect 136393 -14097 136604 -14096
rect 136066 -14099 136604 -14097
rect 135747 -14177 136604 -14099
rect 138469 -13441 139326 -13368
rect 138469 -13442 139200 -13441
rect 138469 -13444 138866 -13442
rect 138469 -13532 138539 -13444
rect 138626 -13532 138719 -13444
rect 138806 -13530 138866 -13444
rect 138953 -13530 139046 -13442
rect 139133 -13529 139200 -13442
rect 139287 -13529 139326 -13441
rect 139133 -13530 139326 -13529
rect 138806 -13532 139326 -13530
rect 138469 -13621 139326 -13532
rect 138469 -13622 139200 -13621
rect 138469 -13624 138866 -13622
rect 138469 -13712 138539 -13624
rect 138626 -13712 138719 -13624
rect 138806 -13710 138866 -13624
rect 138953 -13710 139046 -13622
rect 139133 -13709 139200 -13622
rect 139287 -13709 139326 -13621
rect 139133 -13710 139326 -13709
rect 138806 -13712 139326 -13710
rect 138469 -13834 139326 -13712
rect 138469 -13835 139182 -13834
rect 138469 -13837 138848 -13835
rect 138469 -13925 138521 -13837
rect 138608 -13925 138701 -13837
rect 138788 -13923 138848 -13837
rect 138935 -13923 139028 -13835
rect 139115 -13922 139182 -13835
rect 139269 -13922 139326 -13834
rect 139115 -13923 139326 -13922
rect 138788 -13925 139326 -13923
rect 138469 -14014 139326 -13925
rect 138469 -14015 139182 -14014
rect 138469 -14017 138848 -14015
rect 138469 -14105 138521 -14017
rect 138608 -14105 138701 -14017
rect 138788 -14103 138848 -14017
rect 138935 -14103 139028 -14015
rect 139115 -14102 139182 -14015
rect 139269 -14102 139326 -14014
rect 139115 -14103 139326 -14102
rect 138788 -14105 139326 -14103
rect 138469 -14183 139326 -14105
rect 150251 -13408 151108 -13335
rect 150251 -13409 150982 -13408
rect 150251 -13411 150648 -13409
rect 150251 -13499 150321 -13411
rect 150408 -13499 150501 -13411
rect 150588 -13497 150648 -13411
rect 150735 -13497 150828 -13409
rect 150915 -13496 150982 -13409
rect 151069 -13496 151108 -13408
rect 150915 -13497 151108 -13496
rect 150588 -13499 151108 -13497
rect 150251 -13588 151108 -13499
rect 150251 -13589 150982 -13588
rect 150251 -13591 150648 -13589
rect 150251 -13679 150321 -13591
rect 150408 -13679 150501 -13591
rect 150588 -13677 150648 -13591
rect 150735 -13677 150828 -13589
rect 150915 -13676 150982 -13589
rect 151069 -13676 151108 -13588
rect 150915 -13677 151108 -13676
rect 150588 -13679 151108 -13677
rect 150251 -13801 151108 -13679
rect 150251 -13802 150964 -13801
rect 150251 -13804 150630 -13802
rect 150251 -13892 150303 -13804
rect 150390 -13892 150483 -13804
rect 150570 -13890 150630 -13804
rect 150717 -13890 150810 -13802
rect 150897 -13889 150964 -13802
rect 151051 -13889 151108 -13801
rect 150897 -13890 151108 -13889
rect 150570 -13892 151108 -13890
rect 150251 -13981 151108 -13892
rect 150251 -13982 150964 -13981
rect 150251 -13984 150630 -13982
rect 150251 -14072 150303 -13984
rect 150390 -14072 150483 -13984
rect 150570 -14070 150630 -13984
rect 150717 -14070 150810 -13982
rect 150897 -14069 150964 -13982
rect 151051 -14069 151108 -13981
rect 150897 -14070 151108 -14069
rect 150570 -14072 151108 -14070
rect 150251 -14150 151108 -14072
rect 31520 -15275 32448 -15254
rect 29808 -15361 30736 -15340
rect 29808 -15449 29831 -15361
rect 29918 -15449 29991 -15361
rect 30078 -15449 30151 -15361
rect 30238 -15449 30311 -15361
rect 30398 -15449 30471 -15361
rect 30558 -15449 30631 -15361
rect 30718 -15449 30736 -15361
rect 27986 -15478 28914 -15457
rect 27986 -15566 28009 -15478
rect 28096 -15566 28169 -15478
rect 28256 -15566 28329 -15478
rect 28416 -15566 28489 -15478
rect 28576 -15566 28649 -15478
rect 28736 -15566 28809 -15478
rect 28896 -15566 28914 -15478
rect 27986 -15638 28914 -15566
rect 27986 -15726 28009 -15638
rect 28096 -15726 28169 -15638
rect 28256 -15726 28329 -15638
rect 28416 -15726 28489 -15638
rect 28576 -15726 28649 -15638
rect 28736 -15726 28809 -15638
rect 28896 -15726 28914 -15638
rect 27986 -15798 28914 -15726
rect 27986 -15886 28009 -15798
rect 28096 -15886 28169 -15798
rect 28256 -15886 28329 -15798
rect 28416 -15886 28489 -15798
rect 28576 -15886 28649 -15798
rect 28736 -15886 28809 -15798
rect 28896 -15886 28914 -15798
rect 27986 -15958 28914 -15886
rect -77 -15994 236 -15982
rect 17 -16046 236 -15994
rect 27986 -16046 28009 -15958
rect 28096 -16046 28169 -15958
rect 28256 -16046 28329 -15958
rect 28416 -16046 28489 -15958
rect 28576 -16046 28649 -15958
rect 28736 -16046 28809 -15958
rect 28896 -16046 28914 -15958
rect 27986 -16118 28914 -16046
rect 27986 -16206 28009 -16118
rect 28096 -16206 28169 -16118
rect 28256 -16206 28329 -16118
rect 28416 -16206 28489 -16118
rect 28576 -16206 28649 -16118
rect 28736 -16206 28809 -16118
rect 28896 -16206 28914 -16118
rect 27986 -16278 28914 -16206
rect 29808 -15521 30736 -15449
rect 29808 -15609 29831 -15521
rect 29918 -15609 29991 -15521
rect 30078 -15609 30151 -15521
rect 30238 -15609 30311 -15521
rect 30398 -15609 30471 -15521
rect 30558 -15609 30631 -15521
rect 30718 -15609 30736 -15521
rect 29808 -15681 30736 -15609
rect 29808 -15769 29831 -15681
rect 29918 -15769 29991 -15681
rect 30078 -15769 30151 -15681
rect 30238 -15769 30311 -15681
rect 30398 -15769 30471 -15681
rect 30558 -15769 30631 -15681
rect 30718 -15769 30736 -15681
rect 29808 -15841 30736 -15769
rect 29808 -15929 29831 -15841
rect 29918 -15929 29991 -15841
rect 30078 -15929 30151 -15841
rect 30238 -15929 30311 -15841
rect 30398 -15929 30471 -15841
rect 30558 -15929 30631 -15841
rect 30718 -15929 30736 -15841
rect 29808 -16001 30736 -15929
rect 29808 -16089 29831 -16001
rect 29918 -16089 29991 -16001
rect 30078 -16089 30151 -16001
rect 30238 -16089 30311 -16001
rect 30398 -16089 30471 -16001
rect 30558 -16089 30631 -16001
rect 30718 -16089 30736 -16001
rect 29808 -16161 30736 -16089
rect 29808 -16249 29831 -16161
rect 29918 -16249 29991 -16161
rect 30078 -16249 30151 -16161
rect 30238 -16249 30311 -16161
rect 30398 -16249 30471 -16161
rect 30558 -16249 30631 -16161
rect 30718 -16249 30736 -16161
rect 31520 -15363 31543 -15275
rect 31630 -15363 31703 -15275
rect 31790 -15363 31863 -15275
rect 31950 -15363 32023 -15275
rect 32110 -15363 32183 -15275
rect 32270 -15363 32343 -15275
rect 32430 -15363 32448 -15275
rect 31520 -15435 32448 -15363
rect 31520 -15523 31543 -15435
rect 31630 -15523 31703 -15435
rect 31790 -15523 31863 -15435
rect 31950 -15523 32023 -15435
rect 32110 -15523 32183 -15435
rect 32270 -15523 32343 -15435
rect 32430 -15523 32448 -15435
rect 31520 -15595 32448 -15523
rect 31520 -15683 31543 -15595
rect 31630 -15683 31703 -15595
rect 31790 -15683 31863 -15595
rect 31950 -15683 32023 -15595
rect 32110 -15683 32183 -15595
rect 32270 -15683 32343 -15595
rect 32430 -15683 32448 -15595
rect 31520 -15755 32448 -15683
rect 31520 -15843 31543 -15755
rect 31630 -15843 31703 -15755
rect 31790 -15843 31863 -15755
rect 31950 -15843 32023 -15755
rect 32110 -15843 32183 -15755
rect 32270 -15843 32343 -15755
rect 32430 -15843 32448 -15755
rect 31520 -15915 32448 -15843
rect 31520 -16003 31543 -15915
rect 31630 -16003 31703 -15915
rect 31790 -16003 31863 -15915
rect 31950 -16003 32023 -15915
rect 32110 -16003 32183 -15915
rect 32270 -16003 32343 -15915
rect 32430 -16003 32448 -15915
rect 65364 -15979 65646 -14536
rect 75550 -14725 76478 -14704
rect 75550 -14813 75573 -14725
rect 75660 -14813 75733 -14725
rect 75820 -14813 75893 -14725
rect 75980 -14813 76053 -14725
rect 76140 -14813 76213 -14725
rect 76300 -14813 76373 -14725
rect 76460 -14813 76478 -14725
rect 75550 -14885 76478 -14813
rect 75550 -14973 75573 -14885
rect 75660 -14973 75733 -14885
rect 75820 -14973 75893 -14885
rect 75980 -14973 76053 -14885
rect 76140 -14973 76213 -14885
rect 76300 -14973 76373 -14885
rect 76460 -14973 76478 -14885
rect 75550 -15045 76478 -14973
rect 75550 -15133 75573 -15045
rect 75660 -15133 75733 -15045
rect 75820 -15133 75893 -15045
rect 75980 -15133 76053 -15045
rect 76140 -15133 76213 -15045
rect 76300 -15133 76373 -15045
rect 76460 -15133 76478 -15045
rect 75550 -15205 76478 -15133
rect 75550 -15293 75573 -15205
rect 75660 -15293 75733 -15205
rect 75820 -15293 75893 -15205
rect 75980 -15293 76053 -15205
rect 76140 -15293 76213 -15205
rect 76300 -15293 76373 -15205
rect 76460 -15293 76478 -15205
rect 75550 -15365 76478 -15293
rect 75550 -15453 75573 -15365
rect 75660 -15453 75733 -15365
rect 75820 -15453 75893 -15365
rect 75980 -15453 76053 -15365
rect 76140 -15453 76213 -15365
rect 76300 -15453 76373 -15365
rect 76460 -15453 76478 -15365
rect 80725 -14936 81871 -14901
rect 80725 -14937 81435 -14936
rect 80725 -14939 81101 -14937
rect 80725 -15027 80774 -14939
rect 80861 -15027 80954 -14939
rect 81041 -15025 81101 -14939
rect 81188 -15025 81281 -14937
rect 81368 -15024 81435 -14937
rect 81522 -14938 81871 -14936
rect 81522 -14939 81759 -14938
rect 81522 -15024 81605 -14939
rect 81368 -15025 81605 -15024
rect 81041 -15027 81605 -15025
rect 81692 -15026 81759 -14939
rect 81846 -15026 81871 -14938
rect 81692 -15027 81871 -15026
rect 80725 -15116 81871 -15027
rect 80725 -15117 81435 -15116
rect 80725 -15119 81101 -15117
rect 80725 -15207 80774 -15119
rect 80861 -15207 80954 -15119
rect 81041 -15205 81101 -15119
rect 81188 -15205 81281 -15117
rect 81368 -15204 81435 -15117
rect 81522 -15118 81871 -15116
rect 81522 -15119 81759 -15118
rect 81522 -15204 81605 -15119
rect 81368 -15205 81605 -15204
rect 81041 -15207 81605 -15205
rect 81692 -15206 81759 -15119
rect 81846 -15206 81871 -15118
rect 81692 -15207 81871 -15206
rect 80725 -15293 81871 -15207
rect 80725 -15294 81429 -15293
rect 80725 -15296 81095 -15294
rect 80725 -15384 80768 -15296
rect 80855 -15384 80948 -15296
rect 81035 -15382 81095 -15296
rect 81182 -15382 81275 -15294
rect 81362 -15381 81429 -15294
rect 81516 -15295 81871 -15293
rect 81516 -15296 81753 -15295
rect 81516 -15381 81599 -15296
rect 81362 -15382 81599 -15381
rect 81035 -15384 81599 -15382
rect 81686 -15383 81753 -15296
rect 81840 -15383 81871 -15295
rect 81686 -15384 81871 -15383
rect 80725 -15423 81871 -15384
rect 142756 -14953 143567 -14930
rect 142756 -15036 142780 -14953
rect 142863 -15036 142950 -14953
rect 143033 -15036 143120 -14953
rect 143203 -15036 143290 -14953
rect 143373 -15036 143460 -14953
rect 143543 -15036 143567 -14953
rect 142756 -15123 143567 -15036
rect 142756 -15206 142780 -15123
rect 142863 -15206 142950 -15123
rect 143033 -15206 143120 -15123
rect 143203 -15206 143290 -15123
rect 143373 -15206 143460 -15123
rect 143543 -15206 143567 -15123
rect 142756 -15293 143567 -15206
rect 142756 -15376 142780 -15293
rect 142863 -15376 142950 -15293
rect 143033 -15376 143120 -15293
rect 143203 -15376 143290 -15293
rect 143373 -15376 143460 -15293
rect 143543 -15376 143567 -15293
rect 75550 -15525 76478 -15453
rect 75550 -15613 75573 -15525
rect 75660 -15613 75733 -15525
rect 75820 -15613 75893 -15525
rect 75980 -15613 76053 -15525
rect 76140 -15613 76213 -15525
rect 76300 -15613 76373 -15525
rect 76460 -15613 76478 -15525
rect 75550 -15635 76478 -15613
rect 142756 -15463 143567 -15376
rect 142756 -15546 142780 -15463
rect 142863 -15546 142950 -15463
rect 143033 -15546 143120 -15463
rect 143203 -15546 143290 -15463
rect 143373 -15546 143460 -15463
rect 143543 -15546 143567 -15463
rect 142756 -15633 143567 -15546
rect 112965 -15695 113776 -15672
rect 112965 -15778 112989 -15695
rect 113072 -15778 113159 -15695
rect 113242 -15778 113329 -15695
rect 113412 -15778 113499 -15695
rect 113582 -15778 113669 -15695
rect 113752 -15778 113776 -15695
rect 112965 -15865 113776 -15778
rect 80861 -15965 81789 -15944
rect 31520 -16075 32448 -16003
rect 31520 -16163 31543 -16075
rect 31630 -16163 31703 -16075
rect 31790 -16163 31863 -16075
rect 31950 -16163 32023 -16075
rect 32110 -16163 32183 -16075
rect 32270 -16163 32343 -16075
rect 32430 -16163 32448 -16075
rect 31520 -16185 32448 -16163
rect 65068 -16002 65879 -15979
rect 65068 -16085 65092 -16002
rect 65175 -16085 65262 -16002
rect 65345 -16085 65432 -16002
rect 65515 -16085 65602 -16002
rect 65685 -16085 65772 -16002
rect 65855 -16085 65879 -16002
rect 65068 -16172 65879 -16085
rect 29808 -16271 30736 -16249
rect 65068 -16255 65092 -16172
rect 65175 -16255 65262 -16172
rect 65345 -16255 65432 -16172
rect 65515 -16255 65602 -16172
rect 65685 -16255 65772 -16172
rect 65855 -16255 65879 -16172
rect 80861 -16053 80884 -15965
rect 80971 -16053 81044 -15965
rect 81131 -16053 81204 -15965
rect 81291 -16053 81364 -15965
rect 81451 -16053 81524 -15965
rect 81611 -16053 81684 -15965
rect 81771 -16053 81789 -15965
rect 80861 -16125 81789 -16053
rect 27986 -16366 28009 -16278
rect 28096 -16366 28169 -16278
rect 28256 -16366 28329 -16278
rect 28416 -16366 28489 -16278
rect 28576 -16366 28649 -16278
rect 28736 -16366 28809 -16278
rect 28896 -16366 28914 -16278
rect 27986 -16388 28914 -16366
rect 65068 -16342 65879 -16255
rect 65068 -16425 65092 -16342
rect 65175 -16425 65262 -16342
rect 65345 -16425 65432 -16342
rect 65515 -16425 65602 -16342
rect 65685 -16425 65772 -16342
rect 65855 -16425 65879 -16342
rect 65068 -16512 65879 -16425
rect 65068 -16595 65092 -16512
rect 65175 -16595 65262 -16512
rect 65345 -16595 65432 -16512
rect 65515 -16595 65602 -16512
rect 65685 -16595 65772 -16512
rect 65855 -16595 65879 -16512
rect 65068 -16682 65879 -16595
rect 65068 -16765 65092 -16682
rect 65175 -16765 65262 -16682
rect 65345 -16765 65432 -16682
rect 65515 -16765 65602 -16682
rect 65685 -16765 65772 -16682
rect 65855 -16765 65879 -16682
rect 65068 -16788 65879 -16765
rect 75576 -16264 76755 -16205
rect 75576 -16265 76313 -16264
rect 75576 -16267 75979 -16265
rect 75576 -16355 75652 -16267
rect 75739 -16355 75832 -16267
rect 75919 -16353 75979 -16267
rect 76066 -16353 76159 -16265
rect 76246 -16352 76313 -16265
rect 76400 -16266 76755 -16264
rect 76400 -16267 76637 -16266
rect 76400 -16352 76483 -16267
rect 76246 -16353 76483 -16352
rect 75919 -16355 76483 -16353
rect 76570 -16354 76637 -16267
rect 76724 -16354 76755 -16266
rect 76570 -16355 76755 -16354
rect 75576 -16444 76755 -16355
rect 75576 -16445 76313 -16444
rect 75576 -16447 75979 -16445
rect 75576 -16535 75652 -16447
rect 75739 -16535 75832 -16447
rect 75919 -16533 75979 -16447
rect 76066 -16533 76159 -16445
rect 76246 -16532 76313 -16445
rect 76400 -16446 76755 -16444
rect 76400 -16447 76637 -16446
rect 76400 -16532 76483 -16447
rect 76246 -16533 76483 -16532
rect 75919 -16535 76483 -16533
rect 76570 -16534 76637 -16447
rect 76724 -16534 76755 -16446
rect 76570 -16535 76755 -16534
rect 75576 -16621 76755 -16535
rect 75576 -16622 76307 -16621
rect 75576 -16624 75973 -16622
rect 75576 -16712 75646 -16624
rect 75733 -16712 75826 -16624
rect 75913 -16710 75973 -16624
rect 76060 -16710 76153 -16622
rect 76240 -16709 76307 -16622
rect 76394 -16623 76755 -16621
rect 76394 -16624 76631 -16623
rect 76394 -16709 76477 -16624
rect 76240 -16710 76477 -16709
rect 75913 -16712 76477 -16710
rect 76564 -16711 76631 -16624
rect 76718 -16711 76755 -16623
rect 76564 -16712 76755 -16711
rect 75576 -16768 76755 -16712
rect 80861 -16213 80884 -16125
rect 80971 -16213 81044 -16125
rect 81131 -16213 81204 -16125
rect 81291 -16213 81364 -16125
rect 81451 -16213 81524 -16125
rect 81611 -16213 81684 -16125
rect 81771 -16213 81789 -16125
rect 80861 -16285 81789 -16213
rect 80861 -16373 80884 -16285
rect 80971 -16373 81044 -16285
rect 81131 -16373 81204 -16285
rect 81291 -16373 81364 -16285
rect 81451 -16373 81524 -16285
rect 81611 -16373 81684 -16285
rect 81771 -16373 81789 -16285
rect 80861 -16445 81789 -16373
rect 80861 -16533 80884 -16445
rect 80971 -16533 81044 -16445
rect 81131 -16533 81204 -16445
rect 81291 -16533 81364 -16445
rect 81451 -16533 81524 -16445
rect 81611 -16533 81684 -16445
rect 81771 -16533 81789 -16445
rect 112965 -15948 112989 -15865
rect 113072 -15948 113159 -15865
rect 113242 -15948 113329 -15865
rect 113412 -15948 113499 -15865
rect 113582 -15948 113669 -15865
rect 113752 -15948 113776 -15865
rect 112965 -16035 113776 -15948
rect 112965 -16118 112989 -16035
rect 113072 -16118 113159 -16035
rect 113242 -16118 113329 -16035
rect 113412 -16118 113499 -16035
rect 113582 -16118 113669 -16035
rect 113752 -16118 113776 -16035
rect 112965 -16205 113776 -16118
rect 112965 -16288 112989 -16205
rect 113072 -16288 113159 -16205
rect 113242 -16288 113329 -16205
rect 113412 -16288 113499 -16205
rect 113582 -16288 113669 -16205
rect 113752 -16288 113776 -16205
rect 112965 -16375 113776 -16288
rect 112965 -16458 112989 -16375
rect 113072 -16458 113159 -16375
rect 113242 -16458 113329 -16375
rect 113412 -16458 113499 -16375
rect 113582 -16458 113669 -16375
rect 113752 -16458 113776 -16375
rect 112965 -16481 113776 -16458
rect 116695 -15730 117506 -15707
rect 116695 -15813 116719 -15730
rect 116802 -15813 116889 -15730
rect 116972 -15813 117059 -15730
rect 117142 -15813 117229 -15730
rect 117312 -15813 117399 -15730
rect 117482 -15813 117506 -15730
rect 142756 -15716 142780 -15633
rect 142863 -15716 142950 -15633
rect 143033 -15716 143120 -15633
rect 143203 -15716 143290 -15633
rect 143373 -15716 143460 -15633
rect 143543 -15716 143567 -15633
rect 142756 -15739 143567 -15716
rect 144802 -14931 145613 -14908
rect 144802 -15014 144826 -14931
rect 144909 -15014 144996 -14931
rect 145079 -15014 145166 -14931
rect 145249 -15014 145336 -14931
rect 145419 -15014 145506 -14931
rect 145589 -15014 145613 -14931
rect 144802 -15101 145613 -15014
rect 144802 -15184 144826 -15101
rect 144909 -15184 144996 -15101
rect 145079 -15184 145166 -15101
rect 145249 -15184 145336 -15101
rect 145419 -15184 145506 -15101
rect 145589 -15184 145613 -15101
rect 144802 -15271 145613 -15184
rect 144802 -15354 144826 -15271
rect 144909 -15354 144996 -15271
rect 145079 -15354 145166 -15271
rect 145249 -15354 145336 -15271
rect 145419 -15354 145506 -15271
rect 145589 -15354 145613 -15271
rect 144802 -15441 145613 -15354
rect 144802 -15524 144826 -15441
rect 144909 -15524 144996 -15441
rect 145079 -15524 145166 -15441
rect 145249 -15524 145336 -15441
rect 145419 -15524 145506 -15441
rect 145589 -15524 145613 -15441
rect 144802 -15611 145613 -15524
rect 144802 -15694 144826 -15611
rect 144909 -15694 144996 -15611
rect 145079 -15694 145166 -15611
rect 145249 -15694 145336 -15611
rect 145419 -15694 145506 -15611
rect 145589 -15694 145613 -15611
rect 144802 -15717 145613 -15694
rect 146936 -14910 147747 -14887
rect 146936 -14993 146960 -14910
rect 147043 -14993 147130 -14910
rect 147213 -14993 147300 -14910
rect 147383 -14993 147470 -14910
rect 147553 -14993 147640 -14910
rect 147723 -14993 147747 -14910
rect 146936 -15080 147747 -14993
rect 146936 -15163 146960 -15080
rect 147043 -15163 147130 -15080
rect 147213 -15163 147300 -15080
rect 147383 -15163 147470 -15080
rect 147553 -15163 147640 -15080
rect 147723 -15163 147747 -15080
rect 146936 -15250 147747 -15163
rect 146936 -15333 146960 -15250
rect 147043 -15333 147130 -15250
rect 147213 -15333 147300 -15250
rect 147383 -15333 147470 -15250
rect 147553 -15333 147640 -15250
rect 147723 -15333 147747 -15250
rect 146936 -15420 147747 -15333
rect 146936 -15503 146960 -15420
rect 147043 -15503 147130 -15420
rect 147213 -15503 147300 -15420
rect 147383 -15503 147470 -15420
rect 147553 -15503 147640 -15420
rect 147723 -15503 147747 -15420
rect 146936 -15590 147747 -15503
rect 146936 -15673 146960 -15590
rect 147043 -15673 147130 -15590
rect 147213 -15673 147300 -15590
rect 147383 -15673 147470 -15590
rect 147553 -15673 147640 -15590
rect 147723 -15673 147747 -15590
rect 146936 -15696 147747 -15673
rect 116695 -15900 117506 -15813
rect 116695 -15983 116719 -15900
rect 116802 -15983 116889 -15900
rect 116972 -15983 117059 -15900
rect 117142 -15983 117229 -15900
rect 117312 -15983 117399 -15900
rect 117482 -15983 117506 -15900
rect 116695 -16070 117506 -15983
rect 116695 -16153 116719 -16070
rect 116802 -16153 116889 -16070
rect 116972 -16153 117059 -16070
rect 117142 -16153 117229 -16070
rect 117312 -16153 117399 -16070
rect 117482 -16153 117506 -16070
rect 116695 -16240 117506 -16153
rect 116695 -16323 116719 -16240
rect 116802 -16323 116889 -16240
rect 116972 -16323 117059 -16240
rect 117142 -16323 117229 -16240
rect 117312 -16323 117399 -16240
rect 117482 -16323 117506 -16240
rect 116695 -16410 117506 -16323
rect 80861 -16605 81789 -16533
rect 80861 -16693 80884 -16605
rect 80971 -16693 81044 -16605
rect 81131 -16693 81204 -16605
rect 81291 -16693 81364 -16605
rect 81451 -16693 81524 -16605
rect 81611 -16693 81684 -16605
rect 81771 -16693 81789 -16605
rect 80861 -16765 81789 -16693
rect -5825 -17652 -5099 -17569
rect -5016 -17652 -4929 -17569
rect -4846 -17652 -4759 -17569
rect -4676 -17652 -4589 -17569
rect -4506 -17652 -4419 -17569
rect -4336 -17652 -4313 -17569
rect -5825 -17739 -4313 -17652
rect -5825 -17822 -5099 -17739
rect -5016 -17822 -4929 -17739
rect -4846 -17822 -4759 -17739
rect -4676 -17822 -4589 -17739
rect -4506 -17822 -4419 -17739
rect -4336 -17822 -4313 -17739
rect -1140 -17524 -802 -17506
rect -1140 -17580 -1129 -17524
rect -1073 -17580 -1025 -17524
rect -969 -17580 -921 -17524
rect -865 -17580 -802 -17524
rect -1140 -17628 -802 -17580
rect -1140 -17684 -1129 -17628
rect -1073 -17684 -1025 -17628
rect -969 -17684 -921 -17628
rect -865 -17684 -802 -17628
rect -1140 -17732 -802 -17684
rect -1140 -17788 -1129 -17732
rect -1073 -17788 -1025 -17732
rect -969 -17788 -921 -17732
rect -865 -17788 -802 -17732
rect -1140 -17800 -802 -17788
rect 16080 -17003 16891 -16980
rect 20058 -16987 20869 -16964
rect 16080 -17086 16104 -17003
rect 16187 -17086 16274 -17003
rect 16357 -17086 16444 -17003
rect 16527 -17086 16614 -17003
rect 16697 -17086 16784 -17003
rect 16867 -17086 16891 -17003
rect 16080 -17173 16891 -17086
rect 16080 -17256 16104 -17173
rect 16187 -17256 16274 -17173
rect 16357 -17256 16444 -17173
rect 16527 -17256 16614 -17173
rect 16697 -17256 16784 -17173
rect 16867 -17256 16891 -17173
rect 16080 -17343 16891 -17256
rect 16080 -17426 16104 -17343
rect 16187 -17426 16274 -17343
rect 16357 -17426 16444 -17343
rect 16527 -17426 16614 -17343
rect 16697 -17426 16784 -17343
rect 16867 -17426 16891 -17343
rect 16080 -17513 16891 -17426
rect 16080 -17596 16104 -17513
rect 16187 -17596 16274 -17513
rect 16357 -17596 16444 -17513
rect 16527 -17596 16614 -17513
rect 16697 -17596 16784 -17513
rect 16867 -17596 16891 -17513
rect 16080 -17683 16891 -17596
rect 16080 -17766 16104 -17683
rect 16187 -17766 16274 -17683
rect 16357 -17766 16444 -17683
rect 16527 -17766 16614 -17683
rect 16697 -17766 16784 -17683
rect 16867 -17766 16891 -17683
rect 16080 -17789 16891 -17766
rect 17986 -17011 18797 -16988
rect 17986 -17094 18010 -17011
rect 18093 -17094 18180 -17011
rect 18263 -17094 18350 -17011
rect 18433 -17094 18520 -17011
rect 18603 -17094 18690 -17011
rect 18773 -17094 18797 -17011
rect 17986 -17181 18797 -17094
rect 17986 -17264 18010 -17181
rect 18093 -17264 18180 -17181
rect 18263 -17264 18350 -17181
rect 18433 -17264 18520 -17181
rect 18603 -17264 18690 -17181
rect 18773 -17264 18797 -17181
rect 17986 -17351 18797 -17264
rect 17986 -17434 18010 -17351
rect 18093 -17434 18180 -17351
rect 18263 -17434 18350 -17351
rect 18433 -17434 18520 -17351
rect 18603 -17434 18690 -17351
rect 18773 -17434 18797 -17351
rect 17986 -17521 18797 -17434
rect 17986 -17604 18010 -17521
rect 18093 -17604 18180 -17521
rect 18263 -17604 18350 -17521
rect 18433 -17604 18520 -17521
rect 18603 -17604 18690 -17521
rect 18773 -17604 18797 -17521
rect 17986 -17691 18797 -17604
rect 17986 -17774 18010 -17691
rect 18093 -17774 18180 -17691
rect 18263 -17774 18350 -17691
rect 18433 -17774 18520 -17691
rect 18603 -17774 18690 -17691
rect 18773 -17774 18797 -17691
rect 20058 -17070 20082 -16987
rect 20165 -17070 20252 -16987
rect 20335 -17070 20422 -16987
rect 20505 -17070 20592 -16987
rect 20675 -17070 20762 -16987
rect 20845 -17070 20869 -16987
rect 20058 -17157 20869 -17070
rect 20058 -17240 20082 -17157
rect 20165 -17240 20252 -17157
rect 20335 -17240 20422 -17157
rect 20505 -17240 20592 -17157
rect 20675 -17240 20762 -17157
rect 20845 -17240 20869 -17157
rect 20058 -17327 20869 -17240
rect 20058 -17410 20082 -17327
rect 20165 -17410 20252 -17327
rect 20335 -17410 20422 -17327
rect 20505 -17410 20592 -17327
rect 20675 -17410 20762 -17327
rect 20845 -17410 20869 -17327
rect 20058 -17497 20869 -17410
rect 65147 -17491 65814 -16788
rect 80861 -16853 80884 -16765
rect 80971 -16853 81044 -16765
rect 81131 -16853 81204 -16765
rect 81291 -16853 81364 -16765
rect 81451 -16853 81524 -16765
rect 81611 -16853 81684 -16765
rect 81771 -16853 81789 -16765
rect 80861 -16875 81789 -16853
rect 113044 -17184 113711 -16481
rect 116695 -16493 116719 -16410
rect 116802 -16493 116889 -16410
rect 116972 -16493 117059 -16410
rect 117142 -16493 117229 -16410
rect 117312 -16493 117399 -16410
rect 117482 -16493 117506 -16410
rect 142835 -16442 143502 -15739
rect 144881 -16420 145548 -15717
rect 147015 -16399 147682 -15696
rect 116695 -16516 117506 -16493
rect 116774 -17219 117441 -16516
rect 20058 -17580 20082 -17497
rect 20165 -17580 20252 -17497
rect 20335 -17580 20422 -17497
rect 20505 -17580 20592 -17497
rect 20675 -17580 20762 -17497
rect 20845 -17580 20869 -17497
rect 20058 -17667 20869 -17580
rect 20058 -17750 20082 -17667
rect 20165 -17750 20252 -17667
rect 20335 -17750 20422 -17667
rect 20505 -17750 20592 -17667
rect 20675 -17750 20762 -17667
rect 20845 -17750 20869 -17667
rect 20058 -17773 20869 -17750
rect -1020 -17804 -802 -17800
rect -5825 -17909 -4313 -17822
rect -5825 -17951 -5099 -17909
rect -5122 -17992 -5099 -17951
rect -5016 -17992 -4929 -17909
rect -4846 -17992 -4759 -17909
rect -4676 -17992 -4589 -17909
rect -4506 -17992 -4419 -17909
rect -4336 -17992 -4313 -17909
rect -5122 -18016 -4313 -17992
rect 288 -18349 1099 -18326
rect 288 -18432 312 -18349
rect 395 -18432 482 -18349
rect 565 -18432 652 -18349
rect 735 -18432 822 -18349
rect 905 -18432 992 -18349
rect 1075 -18432 1099 -18349
rect 288 -18519 1099 -18432
rect 16159 -18492 16826 -17789
rect 17986 -17797 18797 -17774
rect 18065 -18500 18732 -17797
rect 20137 -18476 20804 -17773
rect 27267 -18163 28195 -18142
rect 27267 -18251 27290 -18163
rect 27377 -18251 27450 -18163
rect 27537 -18251 27610 -18163
rect 27697 -18251 27770 -18163
rect 27857 -18251 27930 -18163
rect 28017 -18251 28090 -18163
rect 28177 -18251 28195 -18163
rect 27267 -18323 28195 -18251
rect 27267 -18411 27290 -18323
rect 27377 -18411 27450 -18323
rect 27537 -18411 27610 -18323
rect 27697 -18411 27770 -18323
rect 27857 -18411 27930 -18323
rect 28017 -18411 28090 -18323
rect 28177 -18411 28195 -18323
rect 27267 -18483 28195 -18411
rect 288 -18602 312 -18519
rect 395 -18602 482 -18519
rect 565 -18602 652 -18519
rect 735 -18602 822 -18519
rect 905 -18602 992 -18519
rect 1075 -18602 1099 -18519
rect 288 -18689 1099 -18602
rect 288 -18772 312 -18689
rect 395 -18772 482 -18689
rect 565 -18772 652 -18689
rect 735 -18772 822 -18689
rect 905 -18772 992 -18689
rect 1075 -18772 1099 -18689
rect 288 -18859 1099 -18772
rect 288 -18942 312 -18859
rect 395 -18942 482 -18859
rect 565 -18942 652 -18859
rect 735 -18942 822 -18859
rect 905 -18942 992 -18859
rect 1075 -18942 1099 -18859
rect 288 -19029 1099 -18942
rect 288 -19112 312 -19029
rect 395 -19112 482 -19029
rect 565 -19112 652 -19029
rect 735 -19112 822 -19029
rect 905 -19112 992 -19029
rect 1075 -19112 1099 -19029
rect 27267 -18571 27290 -18483
rect 27377 -18571 27450 -18483
rect 27537 -18571 27610 -18483
rect 27697 -18571 27770 -18483
rect 27857 -18571 27930 -18483
rect 28017 -18571 28090 -18483
rect 28177 -18571 28195 -18483
rect 27267 -18643 28195 -18571
rect 27267 -18731 27290 -18643
rect 27377 -18731 27450 -18643
rect 27537 -18731 27610 -18643
rect 27697 -18731 27770 -18643
rect 27857 -18731 27930 -18643
rect 28017 -18731 28090 -18643
rect 28177 -18731 28195 -18643
rect 27267 -18803 28195 -18731
rect 27267 -18891 27290 -18803
rect 27377 -18891 27450 -18803
rect 27537 -18891 27610 -18803
rect 27697 -18891 27770 -18803
rect 27857 -18891 27930 -18803
rect 28017 -18891 28090 -18803
rect 28177 -18891 28195 -18803
rect 27267 -18963 28195 -18891
rect 27267 -19051 27290 -18963
rect 27377 -19051 27450 -18963
rect 27537 -19051 27610 -18963
rect 27697 -19051 27770 -18963
rect 27857 -19051 27930 -18963
rect 28017 -19051 28090 -18963
rect 28177 -19051 28195 -18963
rect 27267 -19073 28195 -19051
rect 288 -19135 1099 -19112
rect 367 -19838 1034 -19135
rect 27896 -19446 28694 -19411
rect 27896 -19447 28594 -19446
rect 27896 -19449 28260 -19447
rect 27896 -19537 27933 -19449
rect 28020 -19537 28113 -19449
rect 28200 -19535 28260 -19449
rect 28347 -19535 28440 -19447
rect 28527 -19534 28594 -19447
rect 28681 -19534 28694 -19446
rect 28527 -19535 28694 -19534
rect 28200 -19537 28694 -19535
rect 27896 -19569 28694 -19537
<< via3 >>
rect 23348 12787 23435 12875
rect 23528 12787 23615 12875
rect 23348 12607 23435 12695
rect 23528 12607 23615 12695
rect 133349 14349 133436 14437
rect 133529 14349 133616 14437
rect 133676 14351 133763 14439
rect 133856 14351 133943 14439
rect 134010 14352 134097 14440
rect 133349 14169 133436 14257
rect 133529 14169 133616 14257
rect 133676 14171 133763 14259
rect 133856 14171 133943 14259
rect 134010 14172 134097 14260
rect 133331 13956 133418 14044
rect 133511 13956 133598 14044
rect 133658 13958 133745 14046
rect 133838 13958 133925 14046
rect 133992 13959 134079 14047
rect 133331 13776 133418 13864
rect 133511 13776 133598 13864
rect 133658 13778 133745 13866
rect 133838 13778 133925 13866
rect 133992 13779 134079 13867
rect 135855 14333 135942 14421
rect 136035 14333 136122 14421
rect 136182 14335 136269 14423
rect 136362 14335 136449 14423
rect 136516 14336 136603 14424
rect 135855 14153 135942 14241
rect 136035 14153 136122 14241
rect 136182 14155 136269 14243
rect 136362 14155 136449 14243
rect 136516 14156 136603 14244
rect 135837 13940 135924 14028
rect 136017 13940 136104 14028
rect 136164 13942 136251 14030
rect 136344 13942 136431 14030
rect 136498 13943 136585 14031
rect 135837 13760 135924 13848
rect 136017 13760 136104 13848
rect 136164 13762 136251 13850
rect 136344 13762 136431 13850
rect 136498 13763 136585 13851
rect 138571 14352 138658 14440
rect 138751 14352 138838 14440
rect 138898 14354 138985 14442
rect 139078 14354 139165 14442
rect 139232 14355 139319 14443
rect 138571 14172 138658 14260
rect 138751 14172 138838 14260
rect 138898 14174 138985 14262
rect 139078 14174 139165 14262
rect 139232 14175 139319 14263
rect 138553 13959 138640 14047
rect 138733 13959 138820 14047
rect 138880 13961 138967 14049
rect 139060 13961 139147 14049
rect 139214 13962 139301 14050
rect 138553 13779 138640 13867
rect 138733 13779 138820 13867
rect 138880 13781 138967 13869
rect 139060 13781 139147 13869
rect 139214 13782 139301 13870
rect 150342 6580 150429 6668
rect 150522 6580 150609 6668
rect 150669 6582 150756 6670
rect 150849 6582 150936 6670
rect 151003 6583 151090 6671
rect 150342 6400 150429 6488
rect 150522 6400 150609 6488
rect 150669 6402 150756 6490
rect 150849 6402 150936 6490
rect 151003 6403 151090 6491
rect 28075 589 28162 677
rect 28255 589 28342 677
rect 28402 591 28489 679
rect 28582 591 28669 679
rect 28736 592 28823 680
rect 28075 409 28162 497
rect 28255 409 28342 497
rect 28402 411 28489 499
rect 28582 411 28669 499
rect 28736 412 28823 500
rect 28057 196 28144 284
rect 28237 196 28324 284
rect 28384 198 28471 286
rect 28564 198 28651 286
rect 28718 199 28805 287
rect 28057 16 28144 104
rect 28237 16 28324 104
rect 28384 18 28471 106
rect 28564 18 28651 106
rect 28718 19 28805 107
rect 29881 636 29968 724
rect 30061 636 30148 724
rect 30208 638 30295 726
rect 30388 638 30475 726
rect 30542 639 30629 727
rect 29881 456 29968 544
rect 30061 456 30148 544
rect 30208 458 30295 546
rect 30388 458 30475 546
rect 30542 459 30629 547
rect 29887 248 29974 336
rect 30067 248 30154 336
rect 30214 250 30301 338
rect 30394 250 30481 338
rect 30548 251 30635 339
rect 29887 68 29974 156
rect 30067 68 30154 156
rect 30214 70 30301 158
rect 30394 70 30481 158
rect 30548 71 30635 159
rect 31618 636 31705 724
rect 31798 636 31885 724
rect 31945 638 32032 726
rect 32125 638 32212 726
rect 32279 639 32366 727
rect 31618 456 31705 544
rect 31798 456 31885 544
rect 31945 458 32032 546
rect 32125 458 32212 546
rect 32279 459 32366 547
rect 31630 248 31717 336
rect 31810 248 31897 336
rect 31957 250 32044 338
rect 32137 250 32224 338
rect 32291 251 32378 339
rect 31630 68 31717 156
rect 31810 68 31897 156
rect 31957 70 32044 158
rect 32137 70 32224 158
rect 32291 71 32378 159
rect 23089 -2157 23176 -2069
rect 23269 -2157 23356 -2069
rect 23089 -2337 23176 -2249
rect 23269 -2337 23356 -2249
rect 75648 5906 75735 5994
rect 75828 5906 75915 5994
rect 75975 5908 76062 5996
rect 76155 5908 76242 5996
rect 76309 5909 76396 5997
rect 76449 5908 76536 5996
rect 76590 5906 76677 5994
rect 75648 5726 75735 5814
rect 75828 5726 75915 5814
rect 75975 5728 76062 5816
rect 76155 5728 76242 5816
rect 76309 5729 76396 5817
rect 76449 5728 76536 5816
rect 76590 5726 76677 5814
rect 80919 5941 81006 6029
rect 81099 5941 81186 6029
rect 81246 5943 81333 6031
rect 81426 5943 81513 6031
rect 81580 5944 81667 6032
rect 81734 5945 81821 6033
rect 81882 5943 81969 6031
rect 80919 5761 81006 5849
rect 81099 5761 81186 5849
rect 81246 5763 81333 5851
rect 81426 5763 81513 5851
rect 81580 5764 81667 5852
rect 81734 5765 81821 5853
rect 81882 5763 81969 5851
rect 56847 4129 56934 4217
rect 57027 4129 57114 4217
rect 56847 3949 56934 4037
rect 57027 3949 57114 4037
rect 113837 3774 113924 3862
rect 114017 3774 114104 3862
rect 113837 3594 113924 3682
rect 114017 3594 114104 3682
rect 113839 3433 113926 3521
rect 114019 3433 114106 3521
rect 113839 3253 113926 3341
rect 114019 3253 114106 3341
rect 114475 3824 114562 3912
rect 114655 3824 114742 3912
rect 114475 3644 114562 3732
rect 114655 3644 114742 3732
rect 114473 3481 114560 3569
rect 114653 3481 114740 3569
rect 114473 3301 114560 3389
rect 114653 3301 114740 3389
rect 115082 3870 115169 3958
rect 115262 3870 115349 3958
rect 115082 3690 115169 3778
rect 115262 3690 115349 3778
rect 115082 3530 115169 3618
rect 115262 3530 115349 3618
rect 115082 3350 115169 3438
rect 115262 3350 115349 3438
rect 86691 -2219 86778 -2131
rect 86871 -2219 86958 -2131
rect 87037 -2219 87124 -2131
rect 87217 -2219 87304 -2131
rect 87390 -2222 87477 -2134
rect 87570 -2222 87657 -2134
rect 86691 -2399 86778 -2311
rect 86871 -2399 86958 -2311
rect 87037 -2399 87124 -2311
rect 87217 -2399 87304 -2311
rect 87390 -2402 87477 -2314
rect 87570 -2402 87657 -2314
rect 121627 -7169 121714 -7081
rect 121807 -7169 121894 -7081
rect 121973 -7169 122060 -7081
rect 122153 -7169 122240 -7081
rect 122326 -7172 122413 -7084
rect 122506 -7172 122593 -7084
rect 121627 -7349 121714 -7261
rect 121807 -7349 121894 -7261
rect 121973 -7349 122060 -7261
rect 122153 -7349 122240 -7261
rect 122326 -7352 122413 -7264
rect 122506 -7352 122593 -7264
rect 133379 -13521 133466 -13433
rect 133559 -13521 133646 -13433
rect 133706 -13519 133793 -13431
rect 133886 -13519 133973 -13431
rect 134040 -13518 134127 -13430
rect 133379 -13701 133466 -13613
rect 133559 -13701 133646 -13613
rect 133706 -13699 133793 -13611
rect 133886 -13699 133973 -13611
rect 134040 -13698 134127 -13610
rect 133361 -13914 133448 -13826
rect 133541 -13914 133628 -13826
rect 133688 -13912 133775 -13824
rect 133868 -13912 133955 -13824
rect 134022 -13911 134109 -13823
rect 133361 -14094 133448 -14006
rect 133541 -14094 133628 -14006
rect 133688 -14092 133775 -14004
rect 133868 -14092 133955 -14004
rect 134022 -14091 134109 -14003
rect 135817 -13526 135904 -13438
rect 135997 -13526 136084 -13438
rect 136144 -13524 136231 -13436
rect 136324 -13524 136411 -13436
rect 136478 -13523 136565 -13435
rect 135817 -13706 135904 -13618
rect 135997 -13706 136084 -13618
rect 136144 -13704 136231 -13616
rect 136324 -13704 136411 -13616
rect 136478 -13703 136565 -13615
rect 135799 -13919 135886 -13831
rect 135979 -13919 136066 -13831
rect 136126 -13917 136213 -13829
rect 136306 -13917 136393 -13829
rect 136460 -13916 136547 -13828
rect 135799 -14099 135886 -14011
rect 135979 -14099 136066 -14011
rect 136126 -14097 136213 -14009
rect 136306 -14097 136393 -14009
rect 136460 -14096 136547 -14008
rect 138539 -13532 138626 -13444
rect 138719 -13532 138806 -13444
rect 138866 -13530 138953 -13442
rect 139046 -13530 139133 -13442
rect 139200 -13529 139287 -13441
rect 138539 -13712 138626 -13624
rect 138719 -13712 138806 -13624
rect 138866 -13710 138953 -13622
rect 139046 -13710 139133 -13622
rect 139200 -13709 139287 -13621
rect 138521 -13925 138608 -13837
rect 138701 -13925 138788 -13837
rect 138848 -13923 138935 -13835
rect 139028 -13923 139115 -13835
rect 139182 -13922 139269 -13834
rect 138521 -14105 138608 -14017
rect 138701 -14105 138788 -14017
rect 138848 -14103 138935 -14015
rect 139028 -14103 139115 -14015
rect 139182 -14102 139269 -14014
rect 150321 -13499 150408 -13411
rect 150501 -13499 150588 -13411
rect 150648 -13497 150735 -13409
rect 150828 -13497 150915 -13409
rect 150982 -13496 151069 -13408
rect 150321 -13679 150408 -13591
rect 150501 -13679 150588 -13591
rect 150648 -13677 150735 -13589
rect 150828 -13677 150915 -13589
rect 150982 -13676 151069 -13588
rect 150303 -13892 150390 -13804
rect 150483 -13892 150570 -13804
rect 150630 -13890 150717 -13802
rect 150810 -13890 150897 -13802
rect 150964 -13889 151051 -13801
rect 150303 -14072 150390 -13984
rect 150483 -14072 150570 -13984
rect 150630 -14070 150717 -13982
rect 150810 -14070 150897 -13982
rect 150964 -14069 151051 -13981
rect 29831 -15449 29918 -15361
rect 29991 -15449 30078 -15361
rect 30151 -15449 30238 -15361
rect 30311 -15449 30398 -15361
rect 30471 -15449 30558 -15361
rect 30631 -15449 30718 -15361
rect 28009 -15566 28096 -15478
rect 28169 -15566 28256 -15478
rect 28329 -15566 28416 -15478
rect 28489 -15566 28576 -15478
rect 28649 -15566 28736 -15478
rect 28809 -15566 28896 -15478
rect 28009 -15726 28096 -15638
rect 28169 -15726 28256 -15638
rect 28329 -15726 28416 -15638
rect 28489 -15726 28576 -15638
rect 28649 -15726 28736 -15638
rect 28809 -15726 28896 -15638
rect 28009 -15886 28096 -15798
rect 28169 -15886 28256 -15798
rect 28329 -15886 28416 -15798
rect 28489 -15886 28576 -15798
rect 28649 -15886 28736 -15798
rect 28809 -15886 28896 -15798
rect 28009 -16046 28096 -15958
rect 28169 -16046 28256 -15958
rect 28329 -16046 28416 -15958
rect 28489 -16046 28576 -15958
rect 28649 -16046 28736 -15958
rect 28809 -16046 28896 -15958
rect 28009 -16206 28096 -16118
rect 28169 -16206 28256 -16118
rect 28329 -16206 28416 -16118
rect 28489 -16206 28576 -16118
rect 28649 -16206 28736 -16118
rect 28809 -16206 28896 -16118
rect 29831 -15609 29918 -15521
rect 29991 -15609 30078 -15521
rect 30151 -15609 30238 -15521
rect 30311 -15609 30398 -15521
rect 30471 -15609 30558 -15521
rect 30631 -15609 30718 -15521
rect 29831 -15769 29918 -15681
rect 29991 -15769 30078 -15681
rect 30151 -15769 30238 -15681
rect 30311 -15769 30398 -15681
rect 30471 -15769 30558 -15681
rect 30631 -15769 30718 -15681
rect 29831 -15929 29918 -15841
rect 29991 -15929 30078 -15841
rect 30151 -15929 30238 -15841
rect 30311 -15929 30398 -15841
rect 30471 -15929 30558 -15841
rect 30631 -15929 30718 -15841
rect 29831 -16089 29918 -16001
rect 29991 -16089 30078 -16001
rect 30151 -16089 30238 -16001
rect 30311 -16089 30398 -16001
rect 30471 -16089 30558 -16001
rect 30631 -16089 30718 -16001
rect 29831 -16249 29918 -16161
rect 29991 -16249 30078 -16161
rect 30151 -16249 30238 -16161
rect 30311 -16249 30398 -16161
rect 30471 -16249 30558 -16161
rect 30631 -16249 30718 -16161
rect 31543 -15363 31630 -15275
rect 31703 -15363 31790 -15275
rect 31863 -15363 31950 -15275
rect 32023 -15363 32110 -15275
rect 32183 -15363 32270 -15275
rect 32343 -15363 32430 -15275
rect 31543 -15523 31630 -15435
rect 31703 -15523 31790 -15435
rect 31863 -15523 31950 -15435
rect 32023 -15523 32110 -15435
rect 32183 -15523 32270 -15435
rect 32343 -15523 32430 -15435
rect 31543 -15683 31630 -15595
rect 31703 -15683 31790 -15595
rect 31863 -15683 31950 -15595
rect 32023 -15683 32110 -15595
rect 32183 -15683 32270 -15595
rect 32343 -15683 32430 -15595
rect 31543 -15843 31630 -15755
rect 31703 -15843 31790 -15755
rect 31863 -15843 31950 -15755
rect 32023 -15843 32110 -15755
rect 32183 -15843 32270 -15755
rect 32343 -15843 32430 -15755
rect 31543 -16003 31630 -15915
rect 31703 -16003 31790 -15915
rect 31863 -16003 31950 -15915
rect 32023 -16003 32110 -15915
rect 32183 -16003 32270 -15915
rect 32343 -16003 32430 -15915
rect 75573 -14813 75660 -14725
rect 75733 -14813 75820 -14725
rect 75893 -14813 75980 -14725
rect 76053 -14813 76140 -14725
rect 76213 -14813 76300 -14725
rect 76373 -14813 76460 -14725
rect 75573 -14973 75660 -14885
rect 75733 -14973 75820 -14885
rect 75893 -14973 75980 -14885
rect 76053 -14973 76140 -14885
rect 76213 -14973 76300 -14885
rect 76373 -14973 76460 -14885
rect 75573 -15133 75660 -15045
rect 75733 -15133 75820 -15045
rect 75893 -15133 75980 -15045
rect 76053 -15133 76140 -15045
rect 76213 -15133 76300 -15045
rect 76373 -15133 76460 -15045
rect 75573 -15293 75660 -15205
rect 75733 -15293 75820 -15205
rect 75893 -15293 75980 -15205
rect 76053 -15293 76140 -15205
rect 76213 -15293 76300 -15205
rect 76373 -15293 76460 -15205
rect 75573 -15453 75660 -15365
rect 75733 -15453 75820 -15365
rect 75893 -15453 75980 -15365
rect 76053 -15453 76140 -15365
rect 76213 -15453 76300 -15365
rect 76373 -15453 76460 -15365
rect 80774 -15027 80861 -14939
rect 80954 -15027 81041 -14939
rect 81101 -15025 81188 -14937
rect 81281 -15025 81368 -14937
rect 81435 -15024 81522 -14936
rect 81605 -15027 81692 -14939
rect 81759 -15026 81846 -14938
rect 80774 -15207 80861 -15119
rect 80954 -15207 81041 -15119
rect 81101 -15205 81188 -15117
rect 81281 -15205 81368 -15117
rect 81435 -15204 81522 -15116
rect 81605 -15207 81692 -15119
rect 81759 -15206 81846 -15118
rect 80768 -15384 80855 -15296
rect 80948 -15384 81035 -15296
rect 81095 -15382 81182 -15294
rect 81275 -15382 81362 -15294
rect 81429 -15381 81516 -15293
rect 81599 -15384 81686 -15296
rect 81753 -15383 81840 -15295
rect 75573 -15613 75660 -15525
rect 75733 -15613 75820 -15525
rect 75893 -15613 75980 -15525
rect 76053 -15613 76140 -15525
rect 76213 -15613 76300 -15525
rect 76373 -15613 76460 -15525
rect 31543 -16163 31630 -16075
rect 31703 -16163 31790 -16075
rect 31863 -16163 31950 -16075
rect 32023 -16163 32110 -16075
rect 32183 -16163 32270 -16075
rect 32343 -16163 32430 -16075
rect 80884 -16053 80971 -15965
rect 81044 -16053 81131 -15965
rect 81204 -16053 81291 -15965
rect 81364 -16053 81451 -15965
rect 81524 -16053 81611 -15965
rect 81684 -16053 81771 -15965
rect 28009 -16366 28096 -16278
rect 28169 -16366 28256 -16278
rect 28329 -16366 28416 -16278
rect 28489 -16366 28576 -16278
rect 28649 -16366 28736 -16278
rect 28809 -16366 28896 -16278
rect 75652 -16355 75739 -16267
rect 75832 -16355 75919 -16267
rect 75979 -16353 76066 -16265
rect 76159 -16353 76246 -16265
rect 76313 -16352 76400 -16264
rect 76483 -16355 76570 -16267
rect 76637 -16354 76724 -16266
rect 75652 -16535 75739 -16447
rect 75832 -16535 75919 -16447
rect 75979 -16533 76066 -16445
rect 76159 -16533 76246 -16445
rect 76313 -16532 76400 -16444
rect 76483 -16535 76570 -16447
rect 76637 -16534 76724 -16446
rect 75646 -16712 75733 -16624
rect 75826 -16712 75913 -16624
rect 75973 -16710 76060 -16622
rect 76153 -16710 76240 -16622
rect 76307 -16709 76394 -16621
rect 76477 -16712 76564 -16624
rect 76631 -16711 76718 -16623
rect 80884 -16213 80971 -16125
rect 81044 -16213 81131 -16125
rect 81204 -16213 81291 -16125
rect 81364 -16213 81451 -16125
rect 81524 -16213 81611 -16125
rect 81684 -16213 81771 -16125
rect 80884 -16373 80971 -16285
rect 81044 -16373 81131 -16285
rect 81204 -16373 81291 -16285
rect 81364 -16373 81451 -16285
rect 81524 -16373 81611 -16285
rect 81684 -16373 81771 -16285
rect 80884 -16533 80971 -16445
rect 81044 -16533 81131 -16445
rect 81204 -16533 81291 -16445
rect 81364 -16533 81451 -16445
rect 81524 -16533 81611 -16445
rect 81684 -16533 81771 -16445
rect 80884 -16693 80971 -16605
rect 81044 -16693 81131 -16605
rect 81204 -16693 81291 -16605
rect 81364 -16693 81451 -16605
rect 81524 -16693 81611 -16605
rect 81684 -16693 81771 -16605
rect 80884 -16853 80971 -16765
rect 81044 -16853 81131 -16765
rect 81204 -16853 81291 -16765
rect 81364 -16853 81451 -16765
rect 81524 -16853 81611 -16765
rect 81684 -16853 81771 -16765
rect 27290 -18251 27377 -18163
rect 27450 -18251 27537 -18163
rect 27610 -18251 27697 -18163
rect 27770 -18251 27857 -18163
rect 27930 -18251 28017 -18163
rect 28090 -18251 28177 -18163
rect 27290 -18411 27377 -18323
rect 27450 -18411 27537 -18323
rect 27610 -18411 27697 -18323
rect 27770 -18411 27857 -18323
rect 27930 -18411 28017 -18323
rect 28090 -18411 28177 -18323
rect 27290 -18571 27377 -18483
rect 27450 -18571 27537 -18483
rect 27610 -18571 27697 -18483
rect 27770 -18571 27857 -18483
rect 27930 -18571 28017 -18483
rect 28090 -18571 28177 -18483
rect 27290 -18731 27377 -18643
rect 27450 -18731 27537 -18643
rect 27610 -18731 27697 -18643
rect 27770 -18731 27857 -18643
rect 27930 -18731 28017 -18643
rect 28090 -18731 28177 -18643
rect 27290 -18891 27377 -18803
rect 27450 -18891 27537 -18803
rect 27610 -18891 27697 -18803
rect 27770 -18891 27857 -18803
rect 27930 -18891 28017 -18803
rect 28090 -18891 28177 -18803
rect 27290 -19051 27377 -18963
rect 27450 -19051 27537 -18963
rect 27610 -19051 27697 -18963
rect 27770 -19051 27857 -18963
rect 27930 -19051 28017 -18963
rect 28090 -19051 28177 -18963
rect 27933 -19537 28020 -19449
rect 28113 -19537 28200 -19449
rect 28260 -19535 28347 -19447
rect 28440 -19535 28527 -19447
rect 28594 -19534 28681 -19446
<< metal4 >>
rect 133188 14440 134249 14549
rect 133188 14439 134010 14440
rect 133188 14437 133676 14439
rect 133188 14349 133349 14437
rect 133436 14349 133529 14437
rect 133616 14351 133676 14437
rect 133763 14351 133856 14439
rect 133943 14352 134010 14439
rect 134097 14352 134249 14440
rect 133943 14351 134249 14352
rect 133616 14349 134249 14351
rect 133188 14260 134249 14349
rect 133188 14259 134010 14260
rect 133188 14257 133676 14259
rect 133188 14169 133349 14257
rect 133436 14169 133529 14257
rect 133616 14171 133676 14257
rect 133763 14171 133856 14259
rect 133943 14172 134010 14259
rect 134097 14172 134249 14260
rect 133943 14171 134249 14172
rect 133616 14169 134249 14171
rect 133188 14047 134249 14169
rect 133188 14046 133992 14047
rect 133188 14044 133658 14046
rect 133188 13956 133331 14044
rect 133418 13956 133511 14044
rect 133598 13958 133658 14044
rect 133745 13958 133838 14046
rect 133925 13959 133992 14046
rect 134079 13959 134249 14047
rect 133925 13958 134249 13959
rect 133598 13956 134249 13958
rect 133188 13867 134249 13956
rect 133188 13866 133992 13867
rect 133188 13864 133658 13866
rect 133188 13776 133331 13864
rect 133418 13776 133511 13864
rect 133598 13778 133658 13864
rect 133745 13778 133838 13866
rect 133925 13779 133992 13866
rect 134079 13779 134249 13867
rect 133925 13778 134249 13779
rect 133598 13776 134249 13778
rect 23306 12875 115469 13010
rect 23306 12787 23348 12875
rect 23435 12787 23528 12875
rect 23615 12787 115469 12875
rect 23306 12695 115469 12787
rect 23306 12607 23348 12695
rect 23435 12607 23528 12695
rect 23615 12607 115469 12695
rect 23306 12536 115469 12607
rect 25434 10370 114856 10844
rect 25434 -1934 25908 10370
rect 71760 8163 114171 8546
rect 71760 4283 72143 8163
rect 80879 6043 81977 6073
rect 75608 5997 76748 6038
rect 75608 5996 76309 5997
rect 75608 5994 75975 5996
rect 75608 5988 75648 5994
rect 56785 4217 72143 4283
rect 56785 4129 56847 4217
rect 56934 4129 57027 4217
rect 57114 4129 72143 4217
rect 56785 4037 72143 4129
rect 56785 3949 56847 4037
rect 56934 3949 57027 4037
rect 57114 3949 72143 4037
rect 56785 3900 72143 3949
rect 75575 5906 75648 5988
rect 75735 5906 75828 5994
rect 75915 5908 75975 5994
rect 76062 5908 76155 5996
rect 76242 5909 76309 5996
rect 76396 5996 76748 5997
rect 76396 5909 76449 5996
rect 76242 5908 76449 5909
rect 76536 5994 76748 5996
rect 76536 5908 76590 5994
rect 75915 5906 76590 5908
rect 76677 5906 76748 5994
rect 75575 5817 76748 5906
rect 75575 5816 76309 5817
rect 75575 5814 75975 5816
rect 75575 5726 75648 5814
rect 75735 5726 75828 5814
rect 75915 5728 75975 5814
rect 76062 5728 76155 5816
rect 76242 5729 76309 5816
rect 76396 5816 76748 5817
rect 76396 5729 76449 5816
rect 76242 5728 76449 5729
rect 76536 5814 76748 5816
rect 76536 5728 76590 5814
rect 75915 5726 76590 5728
rect 76677 5726 76748 5814
rect 75575 5683 76748 5726
rect 80849 6033 81982 6043
rect 80849 6032 81734 6033
rect 80849 6031 81580 6032
rect 80849 6029 81246 6031
rect 80849 5941 80919 6029
rect 81006 5941 81099 6029
rect 81186 5943 81246 6029
rect 81333 5943 81426 6031
rect 81513 5944 81580 6031
rect 81667 5945 81734 6032
rect 81821 6031 81982 6033
rect 81821 5945 81882 6031
rect 81667 5944 81882 5945
rect 81513 5943 81882 5944
rect 81969 5943 81982 6031
rect 81186 5941 81982 5943
rect 80849 5853 81982 5941
rect 80849 5852 81734 5853
rect 80849 5851 81580 5852
rect 80849 5849 81246 5851
rect 80849 5761 80919 5849
rect 81006 5761 81099 5849
rect 81186 5763 81246 5849
rect 81333 5763 81426 5851
rect 81513 5764 81580 5851
rect 81667 5765 81734 5852
rect 81821 5851 81982 5853
rect 81821 5765 81882 5851
rect 81667 5764 81882 5765
rect 81513 5763 81882 5764
rect 81969 5763 81982 5851
rect 81186 5761 81982 5763
rect 80849 5746 81982 5761
rect 80849 5718 81977 5746
rect 23047 -2069 25908 -1934
rect 23047 -2157 23089 -2069
rect 23176 -2157 23269 -2069
rect 23356 -2157 25908 -2069
rect 23047 -2249 25908 -2157
rect 23047 -2337 23089 -2249
rect 23176 -2337 23269 -2249
rect 23356 -2337 25908 -2249
rect 23047 -2408 25908 -2337
rect 27974 680 28954 810
rect 27974 679 28736 680
rect 27974 677 28402 679
rect 27974 589 28075 677
rect 28162 589 28255 677
rect 28342 591 28402 677
rect 28489 591 28582 679
rect 28669 592 28736 679
rect 28823 592 28954 680
rect 28669 591 28954 592
rect 28342 589 28954 591
rect 27974 500 28954 589
rect 27974 499 28736 500
rect 27974 497 28402 499
rect 27974 409 28075 497
rect 28162 409 28255 497
rect 28342 411 28402 497
rect 28489 411 28582 499
rect 28669 412 28736 499
rect 28823 412 28954 500
rect 28669 411 28954 412
rect 28342 409 28954 411
rect 27974 287 28954 409
rect 27974 286 28718 287
rect 27974 284 28384 286
rect 27974 196 28057 284
rect 28144 196 28237 284
rect 28324 198 28384 284
rect 28471 198 28564 286
rect 28651 199 28718 286
rect 28805 199 28954 287
rect 28651 198 28954 199
rect 28324 196 28954 198
rect 27974 107 28954 196
rect 27974 106 28718 107
rect 27974 104 28384 106
rect 27974 16 28057 104
rect 28144 16 28237 104
rect 28324 18 28384 104
rect 28471 18 28564 106
rect 28651 19 28718 106
rect 28805 19 28954 107
rect 28651 18 28954 19
rect 28324 16 28954 18
rect 27974 -15478 28954 16
rect 27974 -15566 28009 -15478
rect 28096 -15566 28169 -15478
rect 28256 -15566 28329 -15478
rect 28416 -15566 28489 -15478
rect 28576 -15566 28649 -15478
rect 28736 -15566 28809 -15478
rect 28896 -15566 28954 -15478
rect 27974 -15638 28954 -15566
rect 27974 -15726 28009 -15638
rect 28096 -15726 28169 -15638
rect 28256 -15726 28329 -15638
rect 28416 -15726 28489 -15638
rect 28576 -15726 28649 -15638
rect 28736 -15726 28809 -15638
rect 28896 -15726 28954 -15638
rect 27974 -15798 28954 -15726
rect 27974 -15886 28009 -15798
rect 28096 -15886 28169 -15798
rect 28256 -15886 28329 -15798
rect 28416 -15886 28489 -15798
rect 28576 -15886 28649 -15798
rect 28736 -15886 28809 -15798
rect 28896 -15886 28954 -15798
rect 27974 -15958 28954 -15886
rect 27974 -16046 28009 -15958
rect 28096 -16046 28169 -15958
rect 28256 -16046 28329 -15958
rect 28416 -16046 28489 -15958
rect 28576 -16046 28649 -15958
rect 28736 -16046 28809 -15958
rect 28896 -16046 28954 -15958
rect 27974 -16118 28954 -16046
rect 27974 -16206 28009 -16118
rect 28096 -16206 28169 -16118
rect 28256 -16206 28329 -16118
rect 28416 -16206 28489 -16118
rect 28576 -16206 28649 -16118
rect 28736 -16206 28809 -16118
rect 28896 -16206 28954 -16118
rect 27974 -16278 28954 -16206
rect 27974 -16366 28009 -16278
rect 28096 -16366 28169 -16278
rect 28256 -16366 28329 -16278
rect 28416 -16366 28489 -16278
rect 28576 -16366 28649 -16278
rect 28736 -16366 28809 -16278
rect 28896 -16366 28954 -16278
rect 29757 727 30737 832
rect 29757 726 30542 727
rect 29757 724 30208 726
rect 29757 636 29881 724
rect 29968 636 30061 724
rect 30148 638 30208 724
rect 30295 638 30388 726
rect 30475 639 30542 726
rect 30629 639 30737 727
rect 30475 638 30737 639
rect 30148 636 30737 638
rect 29757 547 30737 636
rect 29757 546 30542 547
rect 29757 544 30208 546
rect 29757 456 29881 544
rect 29968 456 30061 544
rect 30148 458 30208 544
rect 30295 458 30388 546
rect 30475 459 30542 546
rect 30629 459 30737 547
rect 30475 458 30737 459
rect 30148 456 30737 458
rect 29757 339 30737 456
rect 29757 338 30548 339
rect 29757 336 30214 338
rect 29757 248 29887 336
rect 29974 248 30067 336
rect 30154 250 30214 336
rect 30301 250 30394 338
rect 30481 251 30548 338
rect 30635 251 30737 339
rect 30481 250 30737 251
rect 30154 248 30737 250
rect 29757 159 30737 248
rect 29757 158 30548 159
rect 29757 156 30214 158
rect 29757 68 29887 156
rect 29974 68 30067 156
rect 30154 70 30214 156
rect 30301 70 30394 158
rect 30481 71 30548 158
rect 30635 71 30737 159
rect 30481 70 30737 71
rect 30154 68 30737 70
rect 29757 -15361 30737 68
rect 29757 -15449 29831 -15361
rect 29918 -15449 29991 -15361
rect 30078 -15449 30151 -15361
rect 30238 -15449 30311 -15361
rect 30398 -15449 30471 -15361
rect 30558 -15449 30631 -15361
rect 30718 -15449 30737 -15361
rect 29757 -15521 30737 -15449
rect 29757 -15609 29831 -15521
rect 29918 -15609 29991 -15521
rect 30078 -15609 30151 -15521
rect 30238 -15609 30311 -15521
rect 30398 -15609 30471 -15521
rect 30558 -15609 30631 -15521
rect 30718 -15609 30737 -15521
rect 29757 -15681 30737 -15609
rect 29757 -15769 29831 -15681
rect 29918 -15769 29991 -15681
rect 30078 -15769 30151 -15681
rect 30238 -15769 30311 -15681
rect 30398 -15769 30471 -15681
rect 30558 -15769 30631 -15681
rect 30718 -15769 30737 -15681
rect 29757 -15841 30737 -15769
rect 29757 -15929 29831 -15841
rect 29918 -15929 29991 -15841
rect 30078 -15929 30151 -15841
rect 30238 -15929 30311 -15841
rect 30398 -15929 30471 -15841
rect 30558 -15929 30631 -15841
rect 30718 -15929 30737 -15841
rect 29757 -16001 30737 -15929
rect 29757 -16089 29831 -16001
rect 29918 -16089 29991 -16001
rect 30078 -16089 30151 -16001
rect 30238 -16089 30311 -16001
rect 30398 -16089 30471 -16001
rect 30558 -16089 30631 -16001
rect 30718 -16089 30737 -16001
rect 29757 -16161 30737 -16089
rect 29757 -16249 29831 -16161
rect 29918 -16249 29991 -16161
rect 30078 -16249 30151 -16161
rect 30238 -16249 30311 -16161
rect 30398 -16249 30471 -16161
rect 30558 -16249 30631 -16161
rect 30718 -16249 30737 -16161
rect 31495 727 32475 810
rect 31495 726 32279 727
rect 31495 724 31945 726
rect 31495 636 31618 724
rect 31705 636 31798 724
rect 31885 638 31945 724
rect 32032 638 32125 726
rect 32212 639 32279 726
rect 32366 639 32475 727
rect 32212 638 32475 639
rect 31885 636 32475 638
rect 31495 547 32475 636
rect 31495 546 32279 547
rect 31495 544 31945 546
rect 31495 456 31618 544
rect 31705 456 31798 544
rect 31885 458 31945 544
rect 32032 458 32125 546
rect 32212 459 32279 546
rect 32366 459 32475 547
rect 32212 458 32475 459
rect 31885 456 32475 458
rect 31495 339 32475 456
rect 31495 338 32291 339
rect 31495 336 31957 338
rect 31495 248 31630 336
rect 31717 248 31810 336
rect 31897 250 31957 336
rect 32044 250 32137 338
rect 32224 251 32291 338
rect 32378 251 32475 339
rect 32224 250 32475 251
rect 31897 248 32475 250
rect 31495 159 32475 248
rect 31495 158 32291 159
rect 31495 156 31957 158
rect 31495 68 31630 156
rect 31717 68 31810 156
rect 31897 70 31957 156
rect 32044 70 32137 158
rect 32224 71 32291 158
rect 32378 71 32475 159
rect 32224 70 32475 71
rect 31897 68 32475 70
rect 31495 -15275 32475 68
rect 75575 -14704 76466 5683
rect 31495 -15363 31543 -15275
rect 31630 -15363 31703 -15275
rect 31790 -15363 31863 -15275
rect 31950 -15363 32023 -15275
rect 32110 -15363 32183 -15275
rect 32270 -15363 32343 -15275
rect 32430 -15363 32475 -15275
rect 31495 -15435 32475 -15363
rect 31495 -15523 31543 -15435
rect 31630 -15523 31703 -15435
rect 31790 -15523 31863 -15435
rect 31950 -15523 32023 -15435
rect 32110 -15523 32183 -15435
rect 32270 -15523 32343 -15435
rect 32430 -15523 32475 -15435
rect 31495 -15595 32475 -15523
rect 31495 -15683 31543 -15595
rect 31630 -15683 31703 -15595
rect 31790 -15683 31863 -15595
rect 31950 -15683 32023 -15595
rect 32110 -15683 32183 -15595
rect 32270 -15683 32343 -15595
rect 32430 -15683 32475 -15595
rect 75550 -14725 76478 -14704
rect 75550 -14813 75573 -14725
rect 75660 -14813 75733 -14725
rect 75820 -14813 75893 -14725
rect 75980 -14813 76053 -14725
rect 76140 -14813 76213 -14725
rect 76300 -14813 76373 -14725
rect 76460 -14813 76478 -14725
rect 75550 -14885 76478 -14813
rect 75550 -14973 75573 -14885
rect 75660 -14973 75733 -14885
rect 75820 -14973 75893 -14885
rect 75980 -14973 76053 -14885
rect 76140 -14973 76213 -14885
rect 76300 -14973 76373 -14885
rect 76460 -14973 76478 -14885
rect 80849 -14901 81740 5718
rect 113788 3862 114171 8163
rect 113788 3774 113837 3862
rect 113924 3774 114017 3862
rect 114104 3774 114171 3862
rect 113788 3682 114171 3774
rect 113788 3594 113837 3682
rect 113924 3594 114017 3682
rect 114104 3594 114171 3682
rect 113788 3521 114171 3594
rect 113788 3433 113839 3521
rect 113926 3433 114019 3521
rect 114106 3433 114171 3521
rect 113788 3341 114171 3433
rect 113788 3253 113839 3341
rect 113926 3253 114019 3341
rect 114106 3253 114171 3341
rect 113788 3160 114171 3253
rect 114382 3912 114856 10370
rect 114382 3824 114475 3912
rect 114562 3824 114655 3912
rect 114742 3824 114856 3912
rect 114382 3732 114856 3824
rect 114382 3644 114475 3732
rect 114562 3644 114655 3732
rect 114742 3644 114856 3732
rect 114382 3569 114856 3644
rect 114382 3481 114473 3569
rect 114560 3481 114653 3569
rect 114740 3481 114856 3569
rect 114382 3389 114856 3481
rect 114382 3301 114473 3389
rect 114560 3301 114653 3389
rect 114740 3301 114856 3389
rect 114382 3209 114856 3301
rect 114995 3958 115469 12536
rect 114995 3870 115082 3958
rect 115169 3870 115262 3958
rect 115349 3870 115469 3958
rect 114995 3778 115469 3870
rect 114995 3690 115082 3778
rect 115169 3690 115262 3778
rect 115349 3690 115469 3778
rect 114995 3618 115469 3690
rect 114995 3530 115082 3618
rect 115169 3530 115262 3618
rect 115349 3530 115469 3618
rect 114995 3438 115469 3530
rect 114995 3350 115082 3438
rect 115169 3350 115262 3438
rect 115349 3350 115469 3438
rect 114995 3260 115469 3350
rect 86630 -2131 119145 -1980
rect 86630 -2219 86691 -2131
rect 86778 -2219 86871 -2131
rect 86958 -2219 87037 -2131
rect 87124 -2219 87217 -2131
rect 87304 -2134 119145 -2131
rect 87304 -2219 87390 -2134
rect 86630 -2222 87390 -2219
rect 87477 -2222 87570 -2134
rect 87657 -2222 119145 -2134
rect 86630 -2311 119145 -2222
rect 86630 -2399 86691 -2311
rect 86778 -2399 86871 -2311
rect 86958 -2399 87037 -2311
rect 87124 -2399 87217 -2311
rect 87304 -2314 119145 -2311
rect 87304 -2399 87390 -2314
rect 86630 -2402 87390 -2399
rect 87477 -2402 87570 -2314
rect 87657 -2402 119145 -2314
rect 86630 -2610 119145 -2402
rect 118515 -6875 119145 -2610
rect 118515 -7081 122775 -6875
rect 118515 -7169 121627 -7081
rect 121714 -7169 121807 -7081
rect 121894 -7169 121973 -7081
rect 122060 -7169 122153 -7081
rect 122240 -7084 122775 -7081
rect 122240 -7169 122326 -7084
rect 118515 -7172 122326 -7169
rect 122413 -7172 122506 -7084
rect 122593 -7172 122775 -7084
rect 118515 -7261 122775 -7172
rect 118515 -7349 121627 -7261
rect 121714 -7349 121807 -7261
rect 121894 -7349 121973 -7261
rect 122060 -7349 122153 -7261
rect 122240 -7264 122775 -7261
rect 122240 -7349 122326 -7264
rect 118515 -7352 122326 -7349
rect 122413 -7352 122506 -7264
rect 122593 -7352 122775 -7264
rect 118515 -7505 122775 -7352
rect 133188 -13430 134249 13776
rect 133188 -13431 134040 -13430
rect 133188 -13433 133706 -13431
rect 133188 -13521 133379 -13433
rect 133466 -13521 133559 -13433
rect 133646 -13519 133706 -13433
rect 133793 -13519 133886 -13431
rect 133973 -13518 134040 -13431
rect 134127 -13518 134249 -13430
rect 133973 -13519 134249 -13518
rect 133646 -13521 134249 -13519
rect 133188 -13610 134249 -13521
rect 133188 -13611 134040 -13610
rect 133188 -13613 133706 -13611
rect 133188 -13701 133379 -13613
rect 133466 -13701 133559 -13613
rect 133646 -13699 133706 -13613
rect 133793 -13699 133886 -13611
rect 133973 -13698 134040 -13611
rect 134127 -13698 134249 -13610
rect 133973 -13699 134249 -13698
rect 133646 -13701 134249 -13699
rect 133188 -13823 134249 -13701
rect 133188 -13824 134022 -13823
rect 133188 -13826 133688 -13824
rect 133188 -13914 133361 -13826
rect 133448 -13914 133541 -13826
rect 133628 -13912 133688 -13826
rect 133775 -13912 133868 -13824
rect 133955 -13911 134022 -13824
rect 134109 -13911 134249 -13823
rect 133955 -13912 134249 -13911
rect 133628 -13914 134249 -13912
rect 133188 -14003 134249 -13914
rect 133188 -14004 134022 -14003
rect 133188 -14006 133688 -14004
rect 133188 -14094 133361 -14006
rect 133448 -14094 133541 -14006
rect 133628 -14092 133688 -14006
rect 133775 -14092 133868 -14004
rect 133955 -14091 134022 -14004
rect 134109 -14091 134249 -14003
rect 133955 -14092 134249 -14091
rect 133628 -14094 134249 -14092
rect 133188 -14218 134249 -14094
rect 135672 14424 136733 14617
rect 135672 14423 136516 14424
rect 135672 14421 136182 14423
rect 135672 14333 135855 14421
rect 135942 14333 136035 14421
rect 136122 14335 136182 14421
rect 136269 14335 136362 14423
rect 136449 14336 136516 14423
rect 136603 14336 136733 14424
rect 136449 14335 136733 14336
rect 136122 14333 136733 14335
rect 135672 14244 136733 14333
rect 135672 14243 136516 14244
rect 135672 14241 136182 14243
rect 135672 14153 135855 14241
rect 135942 14153 136035 14241
rect 136122 14155 136182 14241
rect 136269 14155 136362 14243
rect 136449 14156 136516 14243
rect 136603 14156 136733 14244
rect 136449 14155 136733 14156
rect 136122 14153 136733 14155
rect 135672 14031 136733 14153
rect 135672 14030 136498 14031
rect 135672 14028 136164 14030
rect 135672 13940 135837 14028
rect 135924 13940 136017 14028
rect 136104 13942 136164 14028
rect 136251 13942 136344 14030
rect 136431 13943 136498 14030
rect 136585 13943 136733 14031
rect 136431 13942 136733 13943
rect 136104 13940 136733 13942
rect 135672 13851 136733 13940
rect 135672 13850 136498 13851
rect 135672 13848 136164 13850
rect 135672 13760 135837 13848
rect 135924 13760 136017 13848
rect 136104 13762 136164 13848
rect 136251 13762 136344 13850
rect 136431 13763 136498 13850
rect 136585 13763 136733 13851
rect 136431 13762 136733 13763
rect 136104 13760 136733 13762
rect 135672 -13435 136733 13760
rect 135672 -13436 136478 -13435
rect 135672 -13438 136144 -13436
rect 135672 -13526 135817 -13438
rect 135904 -13526 135997 -13438
rect 136084 -13524 136144 -13438
rect 136231 -13524 136324 -13436
rect 136411 -13523 136478 -13436
rect 136565 -13523 136733 -13435
rect 136411 -13524 136733 -13523
rect 136084 -13526 136733 -13524
rect 135672 -13615 136733 -13526
rect 135672 -13616 136478 -13615
rect 135672 -13618 136144 -13616
rect 135672 -13706 135817 -13618
rect 135904 -13706 135997 -13618
rect 136084 -13704 136144 -13618
rect 136231 -13704 136324 -13616
rect 136411 -13703 136478 -13616
rect 136565 -13703 136733 -13615
rect 136411 -13704 136733 -13703
rect 136084 -13706 136733 -13704
rect 135672 -13828 136733 -13706
rect 135672 -13829 136460 -13828
rect 135672 -13831 136126 -13829
rect 135672 -13919 135799 -13831
rect 135886 -13919 135979 -13831
rect 136066 -13917 136126 -13831
rect 136213 -13917 136306 -13829
rect 136393 -13916 136460 -13829
rect 136547 -13916 136733 -13828
rect 136393 -13917 136733 -13916
rect 136066 -13919 136733 -13917
rect 135672 -14008 136733 -13919
rect 135672 -14009 136460 -14008
rect 135672 -14011 136126 -14009
rect 135672 -14099 135799 -14011
rect 135886 -14099 135979 -14011
rect 136066 -14097 136126 -14011
rect 136213 -14097 136306 -14009
rect 136393 -14096 136460 -14009
rect 136547 -14096 136733 -14008
rect 136393 -14097 136733 -14096
rect 136066 -14099 136733 -14097
rect 135672 -14218 136733 -14099
rect 138371 14443 139432 14590
rect 138371 14442 139232 14443
rect 138371 14440 138898 14442
rect 138371 14352 138571 14440
rect 138658 14352 138751 14440
rect 138838 14354 138898 14440
rect 138985 14354 139078 14442
rect 139165 14355 139232 14442
rect 139319 14355 139432 14443
rect 139165 14354 139432 14355
rect 138838 14352 139432 14354
rect 138371 14263 139432 14352
rect 138371 14262 139232 14263
rect 138371 14260 138898 14262
rect 138371 14172 138571 14260
rect 138658 14172 138751 14260
rect 138838 14174 138898 14260
rect 138985 14174 139078 14262
rect 139165 14175 139232 14262
rect 139319 14175 139432 14263
rect 139165 14174 139432 14175
rect 138838 14172 139432 14174
rect 138371 14050 139432 14172
rect 138371 14049 139214 14050
rect 138371 14047 138880 14049
rect 138371 13959 138553 14047
rect 138640 13959 138733 14047
rect 138820 13961 138880 14047
rect 138967 13961 139060 14049
rect 139147 13962 139214 14049
rect 139301 13962 139432 14050
rect 139147 13961 139432 13962
rect 138820 13959 139432 13961
rect 138371 13870 139432 13959
rect 138371 13869 139214 13870
rect 138371 13867 138880 13869
rect 138371 13779 138553 13867
rect 138640 13779 138733 13867
rect 138820 13781 138880 13867
rect 138967 13781 139060 13869
rect 139147 13782 139214 13869
rect 139301 13782 139432 13870
rect 139147 13781 139432 13782
rect 138820 13779 139432 13781
rect 138371 -13441 139432 13779
rect 138371 -13442 139200 -13441
rect 138371 -13444 138866 -13442
rect 138371 -13532 138539 -13444
rect 138626 -13532 138719 -13444
rect 138806 -13530 138866 -13444
rect 138953 -13530 139046 -13442
rect 139133 -13529 139200 -13442
rect 139287 -13529 139432 -13441
rect 139133 -13530 139432 -13529
rect 138806 -13532 139432 -13530
rect 138371 -13621 139432 -13532
rect 138371 -13622 139200 -13621
rect 138371 -13624 138866 -13622
rect 138371 -13712 138539 -13624
rect 138626 -13712 138719 -13624
rect 138806 -13710 138866 -13624
rect 138953 -13710 139046 -13622
rect 139133 -13709 139200 -13622
rect 139287 -13709 139432 -13621
rect 139133 -13710 139432 -13709
rect 138806 -13712 139432 -13710
rect 138371 -13834 139432 -13712
rect 138371 -13835 139182 -13834
rect 138371 -13837 138848 -13835
rect 138371 -13925 138521 -13837
rect 138608 -13925 138701 -13837
rect 138788 -13923 138848 -13837
rect 138935 -13923 139028 -13835
rect 139115 -13922 139182 -13835
rect 139269 -13922 139432 -13834
rect 139115 -13923 139432 -13922
rect 138788 -13925 139432 -13923
rect 138371 -14014 139432 -13925
rect 138371 -14015 139182 -14014
rect 138371 -14017 138848 -14015
rect 138371 -14105 138521 -14017
rect 138608 -14105 138701 -14017
rect 138788 -14103 138848 -14017
rect 138935 -14103 139028 -14015
rect 139115 -14102 139182 -14015
rect 139269 -14102 139432 -14014
rect 139115 -14103 139432 -14102
rect 138788 -14105 139432 -14103
rect 138371 -14196 139432 -14105
rect 150164 6671 151228 6773
rect 150164 6670 151003 6671
rect 150164 6668 150669 6670
rect 150164 6580 150342 6668
rect 150429 6580 150522 6668
rect 150609 6582 150669 6668
rect 150756 6582 150849 6670
rect 150936 6583 151003 6670
rect 151090 6583 151228 6671
rect 150936 6582 151228 6583
rect 150609 6580 151228 6582
rect 150164 6491 151228 6580
rect 150164 6490 151003 6491
rect 150164 6488 150669 6490
rect 150164 6400 150342 6488
rect 150429 6400 150522 6488
rect 150609 6402 150669 6488
rect 150756 6402 150849 6490
rect 150936 6403 151003 6490
rect 151090 6403 151228 6491
rect 150936 6402 151228 6403
rect 150609 6400 151228 6402
rect 150164 -13408 151228 6400
rect 150164 -13409 150982 -13408
rect 150164 -13411 150648 -13409
rect 150164 -13499 150321 -13411
rect 150408 -13499 150501 -13411
rect 150588 -13497 150648 -13411
rect 150735 -13497 150828 -13409
rect 150915 -13496 150982 -13409
rect 151069 -13496 151228 -13408
rect 150915 -13497 151228 -13496
rect 150588 -13499 151228 -13497
rect 150164 -13588 151228 -13499
rect 150164 -13589 150982 -13588
rect 150164 -13591 150648 -13589
rect 150164 -13679 150321 -13591
rect 150408 -13679 150501 -13591
rect 150588 -13677 150648 -13591
rect 150735 -13677 150828 -13589
rect 150915 -13676 150982 -13589
rect 151069 -13676 151228 -13588
rect 150915 -13677 151228 -13676
rect 150588 -13679 151228 -13677
rect 150164 -13801 151228 -13679
rect 150164 -13802 150964 -13801
rect 150164 -13804 150630 -13802
rect 150164 -13892 150303 -13804
rect 150390 -13892 150483 -13804
rect 150570 -13890 150630 -13804
rect 150717 -13890 150810 -13802
rect 150897 -13889 150964 -13802
rect 151051 -13889 151228 -13801
rect 150897 -13890 151228 -13889
rect 150570 -13892 151228 -13890
rect 150164 -13981 151228 -13892
rect 150164 -13982 150964 -13981
rect 150164 -13984 150630 -13982
rect 150164 -14072 150303 -13984
rect 150390 -14072 150483 -13984
rect 150570 -14070 150630 -13984
rect 150717 -14070 150810 -13982
rect 150897 -14069 150964 -13982
rect 151051 -14069 151228 -13981
rect 150897 -14070 151228 -14069
rect 150570 -14072 151228 -14070
rect 150164 -14179 151228 -14072
rect 75550 -15045 76478 -14973
rect 75550 -15133 75573 -15045
rect 75660 -15133 75733 -15045
rect 75820 -15133 75893 -15045
rect 75980 -15133 76053 -15045
rect 76140 -15133 76213 -15045
rect 76300 -15133 76373 -15045
rect 76460 -15133 76478 -15045
rect 75550 -15205 76478 -15133
rect 75550 -15293 75573 -15205
rect 75660 -15293 75733 -15205
rect 75820 -15293 75893 -15205
rect 75980 -15293 76053 -15205
rect 76140 -15293 76213 -15205
rect 76300 -15293 76373 -15205
rect 76460 -15293 76478 -15205
rect 75550 -15365 76478 -15293
rect 75550 -15453 75573 -15365
rect 75660 -15453 75733 -15365
rect 75820 -15453 75893 -15365
rect 75980 -15453 76053 -15365
rect 76140 -15453 76213 -15365
rect 76300 -15453 76373 -15365
rect 76460 -15453 76478 -15365
rect 80725 -14936 81871 -14901
rect 80725 -14937 81435 -14936
rect 80725 -14939 81101 -14937
rect 80725 -15027 80774 -14939
rect 80861 -15027 80954 -14939
rect 81041 -15025 81101 -14939
rect 81188 -15025 81281 -14937
rect 81368 -15024 81435 -14937
rect 81522 -14938 81871 -14936
rect 81522 -14939 81759 -14938
rect 81522 -15024 81605 -14939
rect 81368 -15025 81605 -15024
rect 81041 -15027 81605 -15025
rect 81692 -15026 81759 -14939
rect 81846 -15026 81871 -14938
rect 81692 -15027 81871 -15026
rect 80725 -15116 81871 -15027
rect 80725 -15117 81435 -15116
rect 80725 -15119 81101 -15117
rect 80725 -15207 80774 -15119
rect 80861 -15207 80954 -15119
rect 81041 -15205 81101 -15119
rect 81188 -15205 81281 -15117
rect 81368 -15204 81435 -15117
rect 81522 -15118 81871 -15116
rect 81522 -15119 81759 -15118
rect 81522 -15204 81605 -15119
rect 81368 -15205 81605 -15204
rect 81041 -15207 81605 -15205
rect 81692 -15206 81759 -15119
rect 81846 -15206 81871 -15118
rect 81692 -15207 81871 -15206
rect 80725 -15293 81871 -15207
rect 80725 -15294 81429 -15293
rect 80725 -15296 81095 -15294
rect 80725 -15384 80768 -15296
rect 80855 -15384 80948 -15296
rect 81035 -15382 81095 -15296
rect 81182 -15382 81275 -15294
rect 81362 -15381 81429 -15294
rect 81516 -15295 81871 -15293
rect 81516 -15296 81753 -15295
rect 81516 -15381 81599 -15296
rect 81362 -15382 81599 -15381
rect 81035 -15384 81599 -15382
rect 81686 -15383 81753 -15296
rect 81840 -15383 81871 -15295
rect 81686 -15384 81871 -15383
rect 80725 -15423 81871 -15384
rect 75550 -15525 76478 -15453
rect 75550 -15613 75573 -15525
rect 75660 -15613 75733 -15525
rect 75820 -15613 75893 -15525
rect 75980 -15613 76053 -15525
rect 76140 -15613 76213 -15525
rect 76300 -15613 76373 -15525
rect 76460 -15613 76478 -15525
rect 75550 -15635 76478 -15613
rect 31495 -15755 32475 -15683
rect 31495 -15843 31543 -15755
rect 31630 -15843 31703 -15755
rect 31790 -15843 31863 -15755
rect 31950 -15843 32023 -15755
rect 32110 -15843 32183 -15755
rect 32270 -15843 32343 -15755
rect 32430 -15843 32475 -15755
rect 31495 -15915 32475 -15843
rect 31495 -16003 31543 -15915
rect 31630 -16003 31703 -15915
rect 31790 -16003 31863 -15915
rect 31950 -16003 32023 -15915
rect 32110 -16003 32183 -15915
rect 32270 -16003 32343 -15915
rect 32430 -16003 32475 -15915
rect 31495 -16075 32475 -16003
rect 31495 -16163 31543 -16075
rect 31630 -16163 31703 -16075
rect 31790 -16163 31863 -16075
rect 31950 -16163 32023 -16075
rect 32110 -16163 32183 -16075
rect 32270 -16163 32343 -16075
rect 32430 -16163 32475 -16075
rect 31495 -16209 32475 -16163
rect 75575 -16205 76466 -15635
rect 80849 -15944 81740 -15423
rect 80849 -15965 81789 -15944
rect 80849 -16053 80884 -15965
rect 80971 -16053 81044 -15965
rect 81131 -16053 81204 -15965
rect 81291 -16053 81364 -15965
rect 81451 -16053 81524 -15965
rect 81611 -16053 81684 -15965
rect 81771 -16053 81789 -15965
rect 80849 -16125 81789 -16053
rect 29757 -16300 30737 -16249
rect 75575 -16264 76755 -16205
rect 75575 -16265 76313 -16264
rect 75575 -16267 75979 -16265
rect 27974 -16411 28954 -16366
rect 75575 -16355 75652 -16267
rect 75739 -16355 75832 -16267
rect 75919 -16353 75979 -16267
rect 76066 -16353 76159 -16265
rect 76246 -16352 76313 -16265
rect 76400 -16266 76755 -16264
rect 76400 -16267 76637 -16266
rect 76400 -16352 76483 -16267
rect 76246 -16353 76483 -16352
rect 75919 -16355 76483 -16353
rect 76570 -16354 76637 -16267
rect 76724 -16354 76755 -16266
rect 76570 -16355 76755 -16354
rect 75575 -16444 76755 -16355
rect 75575 -16445 76313 -16444
rect 75575 -16447 75979 -16445
rect 75575 -16535 75652 -16447
rect 75739 -16535 75832 -16447
rect 75919 -16533 75979 -16447
rect 76066 -16533 76159 -16445
rect 76246 -16532 76313 -16445
rect 76400 -16446 76755 -16444
rect 76400 -16447 76637 -16446
rect 76400 -16532 76483 -16447
rect 76246 -16533 76483 -16532
rect 75919 -16535 76483 -16533
rect 76570 -16534 76637 -16447
rect 76724 -16534 76755 -16446
rect 76570 -16535 76755 -16534
rect 75575 -16606 76755 -16535
rect 75576 -16621 76755 -16606
rect 75576 -16622 76307 -16621
rect 75576 -16624 75973 -16622
rect 75576 -16712 75646 -16624
rect 75733 -16712 75826 -16624
rect 75913 -16710 75973 -16624
rect 76060 -16710 76153 -16622
rect 76240 -16709 76307 -16622
rect 76394 -16623 76755 -16621
rect 76394 -16624 76631 -16623
rect 76394 -16709 76477 -16624
rect 76240 -16710 76477 -16709
rect 75913 -16712 76477 -16710
rect 76564 -16711 76631 -16624
rect 76718 -16711 76755 -16623
rect 76564 -16712 76755 -16711
rect 75576 -16768 76755 -16712
rect 80849 -16213 80884 -16125
rect 80971 -16213 81044 -16125
rect 81131 -16213 81204 -16125
rect 81291 -16213 81364 -16125
rect 81451 -16213 81524 -16125
rect 81611 -16213 81684 -16125
rect 81771 -16213 81789 -16125
rect 80849 -16285 81789 -16213
rect 80849 -16373 80884 -16285
rect 80971 -16373 81044 -16285
rect 81131 -16373 81204 -16285
rect 81291 -16373 81364 -16285
rect 81451 -16373 81524 -16285
rect 81611 -16373 81684 -16285
rect 81771 -16373 81789 -16285
rect 80849 -16445 81789 -16373
rect 80849 -16533 80884 -16445
rect 80971 -16533 81044 -16445
rect 81131 -16533 81204 -16445
rect 81291 -16533 81364 -16445
rect 81451 -16533 81524 -16445
rect 81611 -16533 81684 -16445
rect 81771 -16533 81789 -16445
rect 80849 -16605 81789 -16533
rect 80849 -16693 80884 -16605
rect 80971 -16693 81044 -16605
rect 81131 -16693 81204 -16605
rect 81291 -16693 81364 -16605
rect 81451 -16693 81524 -16605
rect 81611 -16693 81684 -16605
rect 81771 -16693 81789 -16605
rect 80849 -16765 81789 -16693
rect 80849 -16853 80884 -16765
rect 80971 -16853 81044 -16765
rect 81131 -16853 81204 -16765
rect 81291 -16853 81364 -16765
rect 81451 -16853 81524 -16765
rect 81611 -16853 81684 -16765
rect 81771 -16853 81789 -16765
rect 80849 -16875 81789 -16853
rect 80849 -16919 81740 -16875
rect 27267 -18163 28195 -18142
rect 27267 -18251 27290 -18163
rect 27377 -18251 27450 -18163
rect 27537 -18251 27610 -18163
rect 27697 -18251 27770 -18163
rect 27857 -18251 27930 -18163
rect 28017 -18251 28090 -18163
rect 28177 -18251 28195 -18163
rect 27267 -18323 28195 -18251
rect 27267 -18411 27290 -18323
rect 27377 -18411 27450 -18323
rect 27537 -18411 27610 -18323
rect 27697 -18411 27770 -18323
rect 27857 -18411 27930 -18323
rect 28017 -18411 28090 -18323
rect 28177 -18411 28195 -18323
rect 27267 -18483 28195 -18411
rect 27267 -18571 27290 -18483
rect 27377 -18571 27450 -18483
rect 27537 -18571 27610 -18483
rect 27697 -18571 27770 -18483
rect 27857 -18571 27930 -18483
rect 28017 -18571 28090 -18483
rect 28177 -18571 28195 -18483
rect 27267 -18643 28195 -18571
rect 27267 -18731 27290 -18643
rect 27377 -18731 27450 -18643
rect 27537 -18731 27610 -18643
rect 27697 -18731 27770 -18643
rect 27857 -18731 27930 -18643
rect 28017 -18731 28090 -18643
rect 28177 -18731 28195 -18643
rect 27267 -18803 28195 -18731
rect 27267 -18891 27290 -18803
rect 27377 -18891 27450 -18803
rect 27537 -18891 27610 -18803
rect 27697 -18891 27770 -18803
rect 27857 -18891 27930 -18803
rect 28017 -18891 28090 -18803
rect 28177 -18891 28195 -18803
rect 27267 -18963 28195 -18891
rect 27267 -19051 27290 -18963
rect 27377 -19051 27450 -18963
rect 27537 -19051 27610 -18963
rect 27697 -19051 27770 -18963
rect 27857 -19051 27930 -18963
rect 28017 -19051 28090 -18963
rect 28177 -19051 28195 -18963
rect 27267 -19073 28195 -19051
rect 27896 -19446 28694 -19411
rect 27896 -19447 28594 -19446
rect 27896 -19449 28260 -19447
rect 27896 -19537 27933 -19449
rect 28020 -19537 28113 -19449
rect 28200 -19535 28260 -19449
rect 28347 -19535 28440 -19447
rect 28527 -19534 28594 -19447
rect 28681 -19534 28694 -19446
rect 28527 -19535 28694 -19534
rect 28200 -19537 28694 -19535
rect 27896 -19569 28694 -19537
use MUX_8x1_Layout  MUX_8x1_Layout_0 ~/GF180Projects/Tapeout/Magic/8x1_MUX
timestamp 1699883071
transform -1 0 10959 0 1 -9355
box -5127 -7616 10259 7767
use MUX_8x1_Layout  MUX_8x1_Layout_1
timestamp 1699883071
transform -1 0 10794 0 1 7414
box -5127 -7616 10259 7767
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_0
timestamp 1699877609
transform 1 0 115631 0 1 1266
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_1
timestamp 1699877609
transform 1 0 115631 0 1 2126
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_2
timestamp 1699877609
transform 1 0 114012 0 1 1266
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_3
timestamp 1699877609
transform 1 0 114012 0 1 2126
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_4
timestamp 1699877609
transform 1 0 114552 0 1 2126
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_5
timestamp 1699877609
transform 1 0 114552 0 1 1266
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_6
timestamp 1699877609
transform 1 0 115092 0 1 2126
box -264 -308 264 308
use nfet_03v3_CT75PZ  nfet_03v3_CT75PZ_7
timestamp 1699877609
transform 1 0 115092 0 1 1266
box -264 -308 264 308
use nfet_03v3_CTB5PZ  nfet_03v3_CTB5PZ_0
timestamp 1699882541
transform 1 0 113578 0 1 1266
box -162 -308 162 308
use nfet_03v3_CTB5PZ  nfet_03v3_CTB5PZ_1
timestamp 1699882541
transform 1 0 113578 0 1 2126
box -162 -308 162 308
use nfet_03v3_CTB5PZ  nfet_03v3_CTB5PZ_2
timestamp 1699882541
transform 1 0 116065 0 1 1266
box -162 -308 162 308
use nfet_03v3_CTB5PZ  nfet_03v3_CTB5PZ_3
timestamp 1699882541
transform 1 0 116065 0 1 2126
box -162 -308 162 308
use PGA_block_mag  PGA_block_mag_0 ~/GF180Projects/Tapeout/Magic/PGA_Block
timestamp 1699938486
transform 1 0 123920 0 1 -774
box -2576 -10349 67418 15396
use ppolyf_u_TVCJSY  ppolyf_u_TVCJSY_0
timestamp 1699871744
transform 1 0 121883 0 1 -3950
box -1264 -986 1264 986
use ppolyf_u_WUY3SH  ppolyf_u_WUY3SH_0
timestamp 1699859038
transform 1 0 48199 0 1 19
box -1124 -1136 1124 1136
use trans_block_mag  trans_block_mag_0 ~/GF180Projects/Tapeout/Magic/Transimp_block
timestamp 1699960019
transform 1 0 54633 0 1 -1503
box -36427 -14224 67418 15554
<< labels >>
flabel metal3 155294 17415 155294 17415 0 FreeSans 3200 0 0 0 OUT_P
port 1 nsew
flabel metal3 157743 17706 157743 17706 0 FreeSans 3200 0 0 0 OUT_N
port 2 nsew
flabel metal3 89645 17598 89645 17598 0 FreeSans 3200 0 0 0 TRS_TST1
port 3 nsew
flabel metal3 85975 17581 85975 17581 0 FreeSans 3200 0 0 0 TRS_TST2
port 4 nsew
flabel metal3 49379 16660 49379 16660 0 FreeSans 3200 0 0 0 BUF_TST1
port 5 nsew
flabel metal3 52838 16734 52838 16734 0 FreeSans 3200 0 0 0 BUF_TST2
port 6 nsew
flabel metal3 65447 -17318 65447 -17318 0 FreeSans 3200 0 0 0 TRS
port 7 nsew
flabel metal3 143153 -16247 143153 -16247 0 FreeSans 3200 0 0 0 PGA_2
port 8 nsew
flabel metal3 145244 -16240 145244 -16240 0 FreeSans 3200 0 0 0 PGA_1
port 9 nsew
flabel metal3 147403 -16235 147403 -16235 0 FreeSans 3200 0 0 0 PGA_3
port 10 nsew
flabel metal3 16266 -18321 16266 -18321 0 FreeSans 3200 0 0 0 MUX_1
port 11 nsew
flabel metal3 18533 -18384 18533 -18384 0 FreeSans 3200 0 0 0 MUX_2
port 12 nsew
flabel metal3 20674 -18380 20674 -18380 0 FreeSans 3200 0 0 0 MUX_3
port 13 nsew
flabel metal1 39576 15801 39576 15801 0 FreeSans 4800 0 0 0 VDD
port 14 nsew
flabel metal1 40277 -16553 40277 -16553 0 FreeSans 4800 0 0 0 VSS
port 15 nsew
flabel metal3 113414 -17062 113414 -17062 0 FreeSans 3200 0 0 0 G_sink_dn
port 74 nsew
flabel metal3 117148 -17097 117148 -17097 0 FreeSans 3200 0 0 0 G_sink_up
port 75 nsew
flabel metal3 -5493 -17643 -5493 -17643 0 FreeSans 3200 0 0 0 IN1_1
port 77 nsew
flabel metal3 -5431 -15835 -5431 -15835 0 FreeSans 3200 0 0 0 IN1_2
port 78 nsew
flabel metal3 -5519 -14074 -5519 -14074 0 FreeSans 3200 0 0 0 IN2_1
port 79 nsew
flabel metal3 -5418 -12239 -5418 -12239 0 FreeSans 3200 0 0 0 IN2_2
port 80 nsew
flabel metal3 -5513 -10098 -5513 -10098 0 FreeSans 3200 0 0 0 IN3_2
port 81 nsew
flabel metal3 -5448 -7984 -5448 -7984 0 FreeSans 3200 0 0 0 IN3_1
port 82 nsew
flabel metal3 -5435 -5131 -5435 -5131 0 FreeSans 3200 0 0 0 IN4_2
port 83 nsew
flabel metal3 -5469 -1965 -5469 -1965 0 FreeSans 3200 0 0 0 IN4_1
port 84 nsew
flabel metal3 -5526 2345 -5526 2345 0 FreeSans 3200 0 0 0 IN5_2
port 85 nsew
flabel metal3 -5326 4928 -5326 4928 0 FreeSans 3200 0 0 0 IN5_1
port 86 nsew
flabel metal3 -5438 6610 -5438 6610 0 FreeSans 3200 0 0 0 IN6_1
port 87 nsew
flabel metal3 -5352 8974 -5352 8974 0 FreeSans 3200 0 0 0 IN6_2
port 88 nsew
flabel metal3 -5263 12309 -5263 12309 0 FreeSans 3200 0 0 0 IN7_1
port 89 nsew
flabel metal3 -5366 15229 -5366 15229 0 FreeSans 3200 0 0 0 IN7_2
port 90 nsew
flabel metal3 2259 17910 2259 17910 0 FreeSans 3200 0 0 0 IN8_2
port 91 nsew
flabel metal3 4384 17932 4384 17932 0 FreeSans 3200 0 0 0 IN8_1
port 92 nsew
flabel metal3 22403 17655 22403 17655 0 FreeSans 3200 0 0 0 MUX_TST1
port 93 nsew
flabel metal3 18357 17705 18357 17705 0 FreeSans 3200 0 0 0 MUX_TST2
port 94 nsew
flabel metal3 714 -19559 714 -19559 0 FreeSans 3200 180 0 0 EN
port 76 nsew
<< end >>
