magic
tech gf180mcuC
magscale 1 10
timestamp 1694159936
<< nwell >>
rect -864 -932 864 932
<< nsubdiff >>
rect -840 895 840 908
rect -840 849 -724 895
rect 724 849 840 895
rect -840 836 840 849
rect -840 792 -768 836
rect -840 -792 -827 792
rect -781 -792 -768 792
rect 768 792 840 836
rect -840 -836 -768 -792
rect 768 -792 781 792
rect 827 -792 840 792
rect 768 -836 840 -792
rect -840 -849 840 -836
rect -840 -895 -724 -849
rect 724 -895 840 -849
rect -840 -908 840 -895
<< nsubdiffcont >>
rect -724 849 724 895
rect -827 -792 -781 792
rect 781 -792 827 792
rect -724 -895 724 -849
<< polysilicon >>
rect -680 735 -520 748
rect -680 689 -667 735
rect -533 689 -520 735
rect -680 646 -520 689
rect -680 -689 -520 -646
rect -680 -735 -667 -689
rect -533 -735 -520 -689
rect -680 -748 -520 -735
rect -440 735 -280 748
rect -440 689 -427 735
rect -293 689 -280 735
rect -440 646 -280 689
rect -440 -689 -280 -646
rect -440 -735 -427 -689
rect -293 -735 -280 -689
rect -440 -748 -280 -735
rect -200 735 -40 748
rect -200 689 -187 735
rect -53 689 -40 735
rect -200 646 -40 689
rect -200 -689 -40 -646
rect -200 -735 -187 -689
rect -53 -735 -40 -689
rect -200 -748 -40 -735
rect 40 735 200 748
rect 40 689 53 735
rect 187 689 200 735
rect 40 646 200 689
rect 40 -689 200 -646
rect 40 -735 53 -689
rect 187 -735 200 -689
rect 40 -748 200 -735
rect 280 735 440 748
rect 280 689 293 735
rect 427 689 440 735
rect 280 646 440 689
rect 280 -689 440 -646
rect 280 -735 293 -689
rect 427 -735 440 -689
rect 280 -748 440 -735
rect 520 735 680 748
rect 520 689 533 735
rect 667 689 680 735
rect 520 646 680 689
rect 520 -689 680 -646
rect 520 -735 533 -689
rect 667 -735 680 -689
rect 520 -748 680 -735
<< polycontact >>
rect -667 689 -533 735
rect -667 -735 -533 -689
rect -427 689 -293 735
rect -427 -735 -293 -689
rect -187 689 -53 735
rect -187 -735 -53 -689
rect 53 689 187 735
rect 53 -735 187 -689
rect 293 689 427 735
rect 293 -735 427 -689
rect 533 689 667 735
rect 533 -735 667 -689
<< ppolyres >>
rect -680 -646 -520 646
rect -440 -646 -280 646
rect -200 -646 -40 646
rect 40 -646 200 646
rect 280 -646 440 646
rect 520 -646 680 646
<< metal1 >>
rect -827 849 -724 895
rect 724 849 827 895
rect -827 792 -781 849
rect 781 792 827 849
rect -678 689 -667 735
rect -533 689 -522 735
rect -438 689 -427 735
rect -293 689 -282 735
rect -198 689 -187 735
rect -53 689 -42 735
rect 42 689 53 735
rect 187 689 198 735
rect 282 689 293 735
rect 427 689 438 735
rect 522 689 533 735
rect 667 689 678 735
rect -678 -735 -667 -689
rect -533 -735 -522 -689
rect -438 -735 -427 -689
rect -293 -735 -282 -689
rect -198 -735 -187 -689
rect -53 -735 -42 -689
rect 42 -735 53 -689
rect 187 -735 198 -689
rect 282 -735 293 -689
rect 427 -735 438 -689
rect 522 -735 533 -689
rect 667 -735 678 -689
rect -827 -849 -781 -792
rect 781 -849 827 -792
rect -827 -895 -724 -849
rect 724 -895 827 -849
<< properties >>
string FIXED_BBOX -804 -872 804 872
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 6.459 m 1 nx 6 wmin 0.80 lmin 1.00 rho 315 val 2.787k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1
<< end >>
