* NGSPICE file created from resistor_PGA_new_flat.ext - technology: gf180mcuC

.subckt resistor_PGA_new_flat A B C D E F G H VDD
X0 F.t1 a_12867_13238.t1 VDD.t8 ppolyf_u r_width=1.2u r_length=1u
X1 a_7427_13890.t1 a_6467_13588.t1 VDD.t28 ppolyf_u r_width=1.2u r_length=1u
X2 a_8387_13238.t1 a_8067_14892.t1 VDD.t4 ppolyf_u r_width=1.2u r_length=1u
X3 a_8387_13238.t0 a_8387_12936.t0 VDD.t4 ppolyf_u r_width=1.2u r_length=1u
X4 a_9987_13890.t0 a_9667_13588.t0 VDD.t32 ppolyf_u r_width=1.2u r_length=1u
X5 A.t0 a_6467_13588.t0 VDD.t19 ppolyf_u r_width=1.2u r_length=1u
X6 a_10627_14542.t1 a_9987_13890.t1 VDD.t23 ppolyf_u r_width=1.2u r_length=1u
X7 VDD.t36 VDD.t37 VDD.t5 ppolyf_u r_width=1.2u r_length=1u
X8 VDD.t6 VDD.t7 VDD.t5 ppolyf_u r_width=1.2u r_length=1u
X9 VDD.t30 VDD.t31 VDD.t1 ppolyf_u r_width=1.2u r_length=1u
X10 a_9347_15194.t1 a_10307_14892.t0 VDD.t22 ppolyf_u r_width=1.2u r_length=1u
X11 VDD.t26 VDD.t27 VDD.t1 ppolyf_u r_width=1.2u r_length=1u
X12 a_7107_14892.t1 a_7427_14240.t1 VDD.t28 ppolyf_u r_width=1.2u r_length=1u
X13 a_9987_13238.t1 a_10307_12936.t1 VDD.t22 ppolyf_u r_width=1.2u r_length=1u
X14 a_11907_13890.t1 a_11587_13588.t0 VDD.t12 ppolyf_u r_width=1.2u r_length=1u
X15 a_9667_14542.t0 a_9987_14240.t1 VDD.t32 ppolyf_u r_width=1.2u r_length=1u
X16 a_12547_15194.t1 D.t1 VDD.t14 ppolyf_u r_width=1.2u r_length=1u
X17 a_6787_15194.t0 a_7107_14892.t0 VDD.t17 ppolyf_u r_width=1.2u r_length=1u
X18 a_12867_13238.t0 a_12547_12936.t0 VDD.t14 ppolyf_u r_width=1.2u r_length=1u
X19 G.t3 a_6467_14240.t1 VDD.t19 ppolyf_u r_width=1.2u r_length=1u
X20 a_7107_13238.t0 a_6787_12936.t1 VDD.t17 ppolyf_u r_width=1.2u r_length=1u
X21 a_10947_13890.t0 a_10627_13588.t0 VDD.t15 ppolyf_u r_width=1.2u r_length=1u
X22 a_8067_14240.t0 a_8707_13588.t0 VDD.t20 ppolyf_u r_width=1.2u r_length=1u
X23 a_9667_15194.t0 a_9347_13890.t0 VDD.t18 ppolyf_u r_width=1.2u r_length=1u
X24 A.t1 A.t2 VDD.t11 ppolyf_u r_width=1.2u r_length=1u
X25 a_9347_13238.t1 a_9667_12936.t1 VDD.t18 ppolyf_u r_width=1.2u r_length=1u
X26 G.t0 G.t1 VDD.t11 ppolyf_u r_width=1.2u r_length=1u
X27 a_7107_14240.t1 a_7747_13588.t1 VDD.t25 ppolyf_u r_width=1.2u r_length=1u
X28 a_11587_14542.t0 a_11907_14240.t0 VDD.t12 ppolyf_u r_width=1.2u r_length=1u
X29 a_11267_13890.t1 a_12227_13588.t0 VDD.t24 ppolyf_u r_width=1.2u r_length=1u
X30 B.t0 a_11907_13238.t0 VDD.t8 ppolyf_u r_width=1.2u r_length=1u
X31 H.t2 a_12227_12936.t1 VDD.t8 ppolyf_u r_width=1.2u r_length=1u
X32 E.t5 a_6787_13588.t1 VDD.t0 ppolyf_u r_width=1.2u r_length=1u
X33 a_10627_14542.t0 a_10947_14240.t0 VDD.t15 ppolyf_u r_width=1.2u r_length=1u
X34 a_8707_14542.t0 a_8067_13890.t1 VDD.t20 ppolyf_u r_width=1.2u r_length=1u
X35 a_11267_13890.t0 a_10307_13588.t0 VDD.t29 ppolyf_u r_width=1.2u r_length=1u
X36 a_9027_13890.t1 a_8707_13588.t1 VDD.t33 ppolyf_u r_width=1.2u r_length=1u
X37 a_7747_14542.t0 a_7107_13890.t1 VDD.t25 ppolyf_u r_width=1.2u r_length=1u
X38 a_10627_15194.t1 a_9027_14892.t1 VDD.t23 ppolyf_u r_width=1.2u r_length=1u
X39 a_10307_14240.t1 a_10627_12936.t0 VDD.t23 ppolyf_u r_width=1.2u r_length=1u
X40 a_8067_13890.t0 a_7747_13588.t0 VDD.t21 ppolyf_u r_width=1.2u r_length=1u
X41 a_12227_14542.t0 a_11267_14240.t0 VDD.t24 ppolyf_u r_width=1.2u r_length=1u
X42 a_7427_13238.t1 a_7427_14892.t1 VDD.t28 ppolyf_u r_width=1.2u r_length=1u
X43 a_6787_14542.t0 E.t0 VDD.t0 ppolyf_u r_width=1.2u r_length=1u
X44 a_7427_13238.t0 a_6467_12936.t1 VDD.t28 ppolyf_u r_width=1.2u r_length=1u
X45 a_10947_14892.t1 a_11267_14240.t1 VDD.t29 ppolyf_u r_width=1.2u r_length=1u
X46 a_8707_14542.t1 a_9027_14240.t0 VDD.t33 ppolyf_u r_width=1.2u r_length=1u
X47 a_9667_15194.t1 a_9987_14892.t0 VDD.t32 ppolyf_u r_width=1.2u r_length=1u
X48 C.t1 a_6467_14892.t1 VDD.t19 ppolyf_u r_width=1.2u r_length=1u
X49 a_9987_13238.t0 a_9667_12936.t0 VDD.t32 ppolyf_u r_width=1.2u r_length=1u
X50 G.t2 a_6467_12936.t0 VDD.t19 ppolyf_u r_width=1.2u r_length=1u
X51 a_12867_14240.t0 F.t0 VDD.t13 ppolyf_u r_width=1.2u r_length=1u
X52 a_7747_14542.t1 a_8067_14240.t1 VDD.t21 ppolyf_u r_width=1.2u r_length=1u
X53 a_11907_14240.t1 a_12547_13588.t0 VDD.t16 ppolyf_u r_width=1.2u r_length=1u
X54 a_11587_15194.t1 a_11907_14892.t1 VDD.t12 ppolyf_u r_width=1.2u r_length=1u
X55 a_11907_13238.t1 a_11587_12936.t0 VDD.t12 ppolyf_u r_width=1.2u r_length=1u
X56 a_10947_14240.t1 a_11587_13588.t1 VDD.t9 ppolyf_u r_width=1.2u r_length=1u
X57 a_9347_13890.t1 a_8387_13588.t1 VDD.t10 ppolyf_u r_width=1.2u r_length=1u
X58 D.t0 a_12867_13890.t0 VDD.t13 ppolyf_u r_width=1.2u r_length=1u
X59 a_10627_15194.t0 a_10947_14892.t0 VDD.t15 ppolyf_u r_width=1.2u r_length=1u
X60 a_8707_15194.t0 a_8387_14542.t1 VDD.t20 ppolyf_u r_width=1.2u r_length=1u
X61 a_10947_13238.t1 a_10627_12936.t1 VDD.t15 ppolyf_u r_width=1.2u r_length=1u
X62 a_7107_13238.t1 a_8707_12936.t0 VDD.t20 ppolyf_u r_width=1.2u r_length=1u
X63 a_12547_14542.t0 a_11907_13890.t0 VDD.t16 ppolyf_u r_width=1.2u r_length=1u
X64 a_7427_13890.t0 a_8387_13588.t0 VDD.t4 ppolyf_u r_width=1.2u r_length=1u
X65 a_7747_15194.t1 a_7427_14892.t0 VDD.t25 ppolyf_u r_width=1.2u r_length=1u
X66 a_6467_14892.t0 a_7747_12936.t0 VDD.t25 ppolyf_u r_width=1.2u r_length=1u
X67 a_11587_14542.t1 a_10947_13890.t1 VDD.t9 ppolyf_u r_width=1.2u r_length=1u
X68 a_9347_14542.t1 a_9027_13238.t0 VDD.t10 ppolyf_u r_width=1.2u r_length=1u
X69 a_12227_13238.t1 a_11907_14892.t0 VDD.t24 ppolyf_u r_width=1.2u r_length=1u
X70 a_12227_13238.t0 a_12227_12936.t0 VDD.t24 ppolyf_u r_width=1.2u r_length=1u
X71 a_6787_15194.t1 C.t0 VDD.t0 ppolyf_u r_width=1.2u r_length=1u
X72 VDD.t34 VDD.t35 VDD.t5 ppolyf_u r_width=1.2u r_length=1u
X73 a_6467_14240.t0 a_6787_12936.t0 VDD.t0 ppolyf_u r_width=1.2u r_length=1u
X74 VDD.t2 VDD.t3 VDD.t1 ppolyf_u r_width=1.2u r_length=1u
X75 a_9987_14892.t1 a_10307_13588.t1 VDD.t22 ppolyf_u r_width=1.2u r_length=1u
X76 a_8387_14542.t0 a_7427_14240.t0 VDD.t4 ppolyf_u r_width=1.2u r_length=1u
X77 a_11267_13238.t0 a_11267_14892.t1 VDD.t29 ppolyf_u r_width=1.2u r_length=1u
X78 a_8707_15194.t1 a_9027_14892.t0 VDD.t33 ppolyf_u r_width=1.2u r_length=1u
X79 a_11267_13238.t1 a_10307_12936.t0 VDD.t29 ppolyf_u r_width=1.2u r_length=1u
X80 a_9027_13238.t1 a_8707_12936.t1 VDD.t33 ppolyf_u r_width=1.2u r_length=1u
X81 a_12867_13890.t1 a_12547_13588.t1 VDD.t14 ppolyf_u r_width=1.2u r_length=1u
X82 a_7107_13890.t0 a_6787_13588.t0 VDD.t17 ppolyf_u r_width=1.2u r_length=1u
X83 a_7747_15194.t0 a_8067_14892.t0 VDD.t21 ppolyf_u r_width=1.2u r_length=1u
X84 a_8067_13238.t1 a_7747_12936.t1 VDD.t21 ppolyf_u r_width=1.2u r_length=1u
X85 VDD.t40 VDD.t41 VDD.t5 ppolyf_u r_width=1.2u r_length=1u
X86 a_9027_14240.t1 a_9667_13588.t1 VDD.t18 ppolyf_u r_width=1.2u r_length=1u
X87 VDD.t38 VDD.t39 VDD.t1 ppolyf_u r_width=1.2u r_length=1u
X88 E.t3 E.t4 VDD.t11 ppolyf_u r_width=1.2u r_length=1u
X89 a_9347_14542.t0 a_10307_14240.t0 VDD.t22 ppolyf_u r_width=1.2u r_length=1u
X90 a_12547_14542.t1 a_12867_14240.t1 VDD.t14 ppolyf_u r_width=1.2u r_length=1u
X91 B.t1 B.t2 VDD.t13 ppolyf_u r_width=1.2u r_length=1u
X92 H.t0 H.t1 VDD.t13 ppolyf_u r_width=1.2u r_length=1u
X93 a_6787_14542.t1 a_7107_14240.t0 VDD.t17 ppolyf_u r_width=1.2u r_length=1u
X94 B.t3 a_12227_13588.t1 VDD.t8 ppolyf_u r_width=1.2u r_length=1u
X95 a_9667_14542.t1 a_9027_13890.t0 VDD.t18 ppolyf_u r_width=1.2u r_length=1u
X96 a_12547_15194.t0 a_12227_14542.t1 VDD.t16 ppolyf_u r_width=1.2u r_length=1u
X97 E.t1 E.t2 VDD.t11 ppolyf_u r_width=1.2u r_length=1u
X98 a_10947_13238.t0 a_12547_12936.t1 VDD.t16 ppolyf_u r_width=1.2u r_length=1u
X99 a_9987_14240.t0 a_10627_13588.t1 VDD.t23 ppolyf_u r_width=1.2u r_length=1u
X100 a_11587_15194.t0 a_11267_14892.t0 VDD.t9 ppolyf_u r_width=1.2u r_length=1u
X101 a_9347_15194.t0 a_8067_13238.t0 VDD.t10 ppolyf_u r_width=1.2u r_length=1u
X102 a_10307_14892.t1 a_11587_12936.t1 VDD.t9 ppolyf_u r_width=1.2u r_length=1u
X103 a_9347_13238.t0 a_8387_12936.t1 VDD.t10 ppolyf_u r_width=1.2u r_length=1u
R0 F F.t0 9.63762
R1 F F.t1 6.8369
R2 a_12867_13238.t0 a_12867_13238.t1 10.61
R3 VDD.n276 VDD.t33 14.599
R4 VDD.n330 VDD.t28 14.599
R5 VDD.n225 VDD.t23 13.9643
R6 VDD.n664 VDD.t5 13.9643
R7 VDD.n174 VDD.t24 13.3296
R8 VDD.n122 VDD.t1 12.6949
R9 VDD.n156 VDD.t14 10.7907
R10 VDD.n207 VDD.t29 10.156
R11 VDD.n258 VDD.t18 9.52129
R12 VDD.n348 VDD.t0 9.52129
R13 VDD.n297 VDD.t4 8.88657
R14 VDD.n309 VDD.t21 8.88657
R15 VDD.n246 VDD.t32 8.25185
R16 VDD.n360 VDD.t19 8.25185
R17 VDD.n195 VDD.t9 7.61713
R18 VDD.n144 VDD.t8 6.98241
R19 VDD.n619 VDD.t40 6.7055
R20 VDD.n82 VDD.t31 6.6704
R21 VDD.n37 VDD.t3 6.55272
R22 VDD.n50 VDD.t2 6.54902
R23 VDD.n0 VDD.t38 6.54788
R24 VDD.n17 VDD.t27 6.54322
R25 VDD.n27 VDD.t26 6.53371
R26 VDD.n668 VDD.t37 6.38623
R27 VDD.n125 VDD.t30 6.35318
R28 VDD.n586 VDD.t6 6.16828
R29 VDD.n384 VDD.t7 6.14788
R30 VDD.n382 VDD.t41 6.14246
R31 VDD.n382 VDD.t34 6.12511
R32 VDD.n0 VDD.t39 6.09716
R33 VDD.n590 VDD.t35 6.01571
R34 VDD.n668 VDD.t36 6.008
R35 VDD.n135 VDD.t13 5.07825
R36 VDD.n186 VDD.t12 4.44353
R37 VDD.n237 VDD.t22 3.80882
R38 VDD.n369 VDD.t11 3.80882
R39 VDD.n288 VDD.t20 3.1741
R40 VDD.n318 VDD.t25 3.1741
R41 VDD.n564 VDD.n381 3.1505
R42 VDD.n641 VDD.n640 3.1505
R43 VDD.n639 VDD.n638 3.1505
R44 VDD.n636 VDD.n635 3.1505
R45 VDD.n634 VDD.n633 3.1505
R46 VDD.n631 VDD.n630 3.1505
R47 VDD.n629 VDD.n628 3.1505
R48 VDD.n626 VDD.n625 3.1505
R49 VDD.n624 VDD.n623 3.1505
R50 VDD.n621 VDD.n620 3.1505
R51 VDD.n618 VDD.n617 3.1505
R52 VDD.n615 VDD.n614 3.1505
R53 VDD.n613 VDD.n612 3.1505
R54 VDD.n610 VDD.n609 3.1505
R55 VDD.n608 VDD.n607 3.1505
R56 VDD.n605 VDD.n604 3.1505
R57 VDD.n603 VDD.n602 3.1505
R58 VDD.n600 VDD.n599 3.1505
R59 VDD.n598 VDD.n597 3.1505
R60 VDD.n596 VDD.n595 3.1505
R61 VDD.n594 VDD.n593 3.1505
R62 VDD.n584 VDD.n583 3.1505
R63 VDD.n582 VDD.n581 3.1505
R64 VDD.n580 VDD.n579 3.1505
R65 VDD.n578 VDD.n577 3.1505
R66 VDD.n576 VDD.n575 3.1505
R67 VDD.n574 VDD.n573 3.1505
R68 VDD.n572 VDD.n571 3.1505
R69 VDD.n570 VDD.n569 3.1505
R70 VDD.n568 VDD.n567 3.1505
R71 VDD.n566 VDD.n565 3.1505
R72 VDD.n652 VDD.n651 3.1505
R73 VDD.n8 VDD.n7 3.1505
R74 VDD.n6 VDD.n5 3.1505
R75 VDD.n4 VDD.n3 3.1505
R76 VDD.n2 VDD.n1 3.1505
R77 VDD.n386 VDD.n385 3.1505
R78 VDD.n388 VDD.n387 3.1505
R79 VDD.n390 VDD.n389 3.1505
R80 VDD.n392 VDD.n391 3.1505
R81 VDD.n394 VDD.n393 3.1505
R82 VDD.n396 VDD.n395 3.1505
R83 VDD.n398 VDD.n397 3.1505
R84 VDD.n400 VDD.n399 3.1505
R85 VDD.n402 VDD.n401 3.1505
R86 VDD.n404 VDD.n403 3.1505
R87 VDD.n406 VDD.n405 3.1505
R88 VDD.n408 VDD.n407 3.1505
R89 VDD.n410 VDD.n409 3.1505
R90 VDD.n412 VDD.n411 3.1505
R91 VDD.n414 VDD.n413 3.1505
R92 VDD.n416 VDD.n415 3.1505
R93 VDD.n418 VDD.n417 3.1505
R94 VDD.n420 VDD.n419 3.1505
R95 VDD.n422 VDD.n421 3.1505
R96 VDD.n424 VDD.n423 3.1505
R97 VDD.n426 VDD.n425 3.1505
R98 VDD.n428 VDD.n427 3.1505
R99 VDD.n430 VDD.n429 3.1505
R100 VDD.n432 VDD.n431 3.1505
R101 VDD.n434 VDD.n433 3.1505
R102 VDD.n436 VDD.n435 3.1505
R103 VDD.n438 VDD.n437 3.1505
R104 VDD.n440 VDD.n439 3.1505
R105 VDD.n442 VDD.n441 3.1505
R106 VDD.n444 VDD.n443 3.1505
R107 VDD.n446 VDD.n445 3.1505
R108 VDD.n448 VDD.n447 3.1505
R109 VDD.n450 VDD.n449 3.1505
R110 VDD.n452 VDD.n451 3.1505
R111 VDD.n454 VDD.n453 3.1505
R112 VDD.n456 VDD.n455 3.1505
R113 VDD.n458 VDD.n457 3.1505
R114 VDD.n460 VDD.n459 3.1505
R115 VDD.n462 VDD.n461 3.1505
R116 VDD.n464 VDD.n463 3.1505
R117 VDD.n466 VDD.n465 3.1505
R118 VDD.n468 VDD.n467 3.1505
R119 VDD.n470 VDD.n469 3.1505
R120 VDD.n472 VDD.n471 3.1505
R121 VDD.n474 VDD.n473 3.1505
R122 VDD.n476 VDD.n475 3.1505
R123 VDD.n478 VDD.n477 3.1505
R124 VDD.n480 VDD.n479 3.1505
R125 VDD.n482 VDD.n481 3.1505
R126 VDD.n484 VDD.n483 3.1505
R127 VDD.n486 VDD.n485 3.1505
R128 VDD.n488 VDD.n487 3.1505
R129 VDD.n490 VDD.n489 3.1505
R130 VDD.n492 VDD.n491 3.1505
R131 VDD.n494 VDD.n493 3.1505
R132 VDD.n496 VDD.n495 3.1505
R133 VDD.n498 VDD.n497 3.1505
R134 VDD.n500 VDD.n499 3.1505
R135 VDD.n502 VDD.n501 3.1505
R136 VDD.n504 VDD.n503 3.1505
R137 VDD.n506 VDD.n505 3.1505
R138 VDD.n508 VDD.n507 3.1505
R139 VDD.n510 VDD.n509 3.1505
R140 VDD.n512 VDD.n511 3.1505
R141 VDD.n514 VDD.n513 3.1505
R142 VDD.n516 VDD.n515 3.1505
R143 VDD.n518 VDD.n517 3.1505
R144 VDD.n520 VDD.n519 3.1505
R145 VDD.n522 VDD.n521 3.1505
R146 VDD.n524 VDD.n523 3.1505
R147 VDD.n526 VDD.n525 3.1505
R148 VDD.n528 VDD.n527 3.1505
R149 VDD.n530 VDD.n529 3.1505
R150 VDD.n532 VDD.n531 3.1505
R151 VDD.n534 VDD.n533 3.1505
R152 VDD.n536 VDD.n535 3.1505
R153 VDD.n538 VDD.n537 3.1505
R154 VDD.n540 VDD.n539 3.1505
R155 VDD.n542 VDD.n541 3.1505
R156 VDD.n544 VDD.n543 3.1505
R157 VDD.n546 VDD.n545 3.1505
R158 VDD.n548 VDD.n547 3.1505
R159 VDD.n550 VDD.n549 3.1505
R160 VDD.n552 VDD.n551 3.1505
R161 VDD.n554 VDD.n553 3.1505
R162 VDD.n557 VDD.n556 3.1505
R163 VDD.n559 VDD.n558 3.1505
R164 VDD.n561 VDD.n560 3.1505
R165 VDD.n563 VDD.n562 3.1505
R166 VDD.n10 VDD.n9 3.1505
R167 VDD.n12 VDD.n11 3.1505
R168 VDD.n14 VDD.n13 3.1505
R169 VDD.n16 VDD.n15 3.1505
R170 VDD.n19 VDD.n18 3.1505
R171 VDD.n21 VDD.n20 3.1505
R172 VDD.n23 VDD.n22 3.1505
R173 VDD.n26 VDD.n25 3.1505
R174 VDD.n30 VDD.n29 3.1505
R175 VDD.n33 VDD.n32 3.1505
R176 VDD.n36 VDD.n35 3.1505
R177 VDD.n40 VDD.n39 3.1505
R178 VDD.n43 VDD.n42 3.1505
R179 VDD.n46 VDD.n45 3.1505
R180 VDD.n49 VDD.n48 3.1505
R181 VDD.n53 VDD.n52 3.1505
R182 VDD.n56 VDD.n55 3.1505
R183 VDD.n59 VDD.n58 3.1505
R184 VDD.n63 VDD.n62 3.1505
R185 VDD.n66 VDD.n65 3.1505
R186 VDD.n69 VDD.n68 3.1505
R187 VDD.n72 VDD.n71 3.1505
R188 VDD.n75 VDD.n74 3.1505
R189 VDD.n78 VDD.n77 3.1505
R190 VDD.n81 VDD.n80 3.1505
R191 VDD.n85 VDD.n84 3.1505
R192 VDD.n88 VDD.n87 3.1505
R193 VDD.n91 VDD.n90 3.1505
R194 VDD.n94 VDD.n93 3.1505
R195 VDD.n97 VDD.n96 3.1505
R196 VDD.n100 VDD.n99 3.1505
R197 VDD.n110 VDD.n109 3.1505
R198 VDD.n112 VDD.n111 3.1505
R199 VDD.n115 VDD.n114 3.1505
R200 VDD.n114 VDD.n113 3.1505
R201 VDD.n118 VDD.n117 3.1505
R202 VDD.n117 VDD.n116 3.1505
R203 VDD.n121 VDD.n120 3.1505
R204 VDD.n120 VDD.n119 3.1505
R205 VDD.n124 VDD.n123 3.1505
R206 VDD.n123 VDD.n122 3.1505
R207 VDD.n128 VDD.n127 3.1505
R208 VDD.n127 VDD.n126 3.1505
R209 VDD.n131 VDD.n130 3.1505
R210 VDD.n130 VDD.n129 3.1505
R211 VDD.n134 VDD.n133 3.1505
R212 VDD.n133 VDD.n132 3.1505
R213 VDD.n137 VDD.n136 3.1505
R214 VDD.n136 VDD.n135 3.1505
R215 VDD.n140 VDD.n139 3.1505
R216 VDD.n139 VDD.n138 3.1505
R217 VDD.n143 VDD.n142 3.1505
R218 VDD.n142 VDD.n141 3.1505
R219 VDD.n146 VDD.n145 3.1505
R220 VDD.n145 VDD.n144 3.1505
R221 VDD.n149 VDD.n148 3.1505
R222 VDD.n148 VDD.n147 3.1505
R223 VDD.n152 VDD.n151 3.1505
R224 VDD.n151 VDD.n150 3.1505
R225 VDD.n155 VDD.n154 3.1505
R226 VDD.n154 VDD.n153 3.1505
R227 VDD.n158 VDD.n157 3.1505
R228 VDD.n157 VDD.n156 3.1505
R229 VDD.n161 VDD.n160 3.1505
R230 VDD.n160 VDD.n159 3.1505
R231 VDD.n164 VDD.n163 3.1505
R232 VDD.n163 VDD.n162 3.1505
R233 VDD.n167 VDD.n166 3.1505
R234 VDD.n166 VDD.n165 3.1505
R235 VDD.n170 VDD.n169 3.1505
R236 VDD.n169 VDD.n168 3.1505
R237 VDD.n173 VDD.n172 3.1505
R238 VDD.n172 VDD.n171 3.1505
R239 VDD.n176 VDD.n175 3.1505
R240 VDD.n175 VDD.n174 3.1505
R241 VDD.n179 VDD.n178 3.1505
R242 VDD.n178 VDD.n177 3.1505
R243 VDD.n182 VDD.n181 3.1505
R244 VDD.n181 VDD.n180 3.1505
R245 VDD.n185 VDD.n184 3.1505
R246 VDD.n184 VDD.n183 3.1505
R247 VDD.n188 VDD.n187 3.1505
R248 VDD.n187 VDD.n186 3.1505
R249 VDD.n191 VDD.n190 3.1505
R250 VDD.n190 VDD.n189 3.1505
R251 VDD.n194 VDD.n193 3.1505
R252 VDD.n193 VDD.n192 3.1505
R253 VDD.n197 VDD.n196 3.1505
R254 VDD.n196 VDD.n195 3.1505
R255 VDD.n200 VDD.n199 3.1505
R256 VDD.n199 VDD.n198 3.1505
R257 VDD.n203 VDD.n202 3.1505
R258 VDD.n202 VDD.n201 3.1505
R259 VDD.n206 VDD.n205 3.1505
R260 VDD.n205 VDD.n204 3.1505
R261 VDD.n209 VDD.n208 3.1505
R262 VDD.n208 VDD.n207 3.1505
R263 VDD.n212 VDD.n211 3.1505
R264 VDD.n211 VDD.n210 3.1505
R265 VDD.n215 VDD.n214 3.1505
R266 VDD.n214 VDD.n213 3.1505
R267 VDD.n218 VDD.n217 3.1505
R268 VDD.n217 VDD.n216 3.1505
R269 VDD.n221 VDD.n220 3.1505
R270 VDD.n220 VDD.n219 3.1505
R271 VDD.n224 VDD.n223 3.1505
R272 VDD.n223 VDD.n222 3.1505
R273 VDD.n227 VDD.n226 3.1505
R274 VDD.n226 VDD.n225 3.1505
R275 VDD.n230 VDD.n229 3.1505
R276 VDD.n229 VDD.n228 3.1505
R277 VDD.n233 VDD.n232 3.1505
R278 VDD.n232 VDD.n231 3.1505
R279 VDD.n236 VDD.n235 3.1505
R280 VDD.n235 VDD.n234 3.1505
R281 VDD.n239 VDD.n238 3.1505
R282 VDD.n238 VDD.n237 3.1505
R283 VDD.n242 VDD.n241 3.1505
R284 VDD.n241 VDD.n240 3.1505
R285 VDD.n245 VDD.n244 3.1505
R286 VDD.n244 VDD.n243 3.1505
R287 VDD.n248 VDD.n247 3.1505
R288 VDD.n247 VDD.n246 3.1505
R289 VDD.n251 VDD.n250 3.1505
R290 VDD.n250 VDD.n249 3.1505
R291 VDD.n254 VDD.n253 3.1505
R292 VDD.n253 VDD.n252 3.1505
R293 VDD.n257 VDD.n256 3.1505
R294 VDD.n256 VDD.n255 3.1505
R295 VDD.n260 VDD.n259 3.1505
R296 VDD.n259 VDD.n258 3.1505
R297 VDD.n263 VDD.n262 3.1505
R298 VDD.n262 VDD.n261 3.1505
R299 VDD.n266 VDD.n265 3.1505
R300 VDD.n265 VDD.n264 3.1505
R301 VDD.n269 VDD.n268 3.1505
R302 VDD.n268 VDD.n267 3.1505
R303 VDD.n272 VDD.n271 3.1505
R304 VDD.n271 VDD.n270 3.1505
R305 VDD.n275 VDD.n274 3.1505
R306 VDD.n274 VDD.n273 3.1505
R307 VDD.n278 VDD.n277 3.1505
R308 VDD.n277 VDD.n276 3.1505
R309 VDD.n281 VDD.n280 3.1505
R310 VDD.n280 VDD.n279 3.1505
R311 VDD.n284 VDD.n283 3.1505
R312 VDD.n283 VDD.n282 3.1505
R313 VDD.n287 VDD.n286 3.1505
R314 VDD.n286 VDD.n285 3.1505
R315 VDD.n290 VDD.n289 3.1505
R316 VDD.n289 VDD.n288 3.1505
R317 VDD.n293 VDD.n292 3.1505
R318 VDD.n292 VDD.n291 3.1505
R319 VDD.n296 VDD.n295 3.1505
R320 VDD.n295 VDD.n294 3.1505
R321 VDD.n299 VDD.n298 3.1505
R322 VDD.n298 VDD.n297 3.1505
R323 VDD.n302 VDD.n301 3.1505
R324 VDD.n301 VDD.n300 3.1505
R325 VDD.n305 VDD.n304 3.1505
R326 VDD.n304 VDD.n303 3.1505
R327 VDD.n308 VDD.n307 3.1505
R328 VDD.n307 VDD.n306 3.1505
R329 VDD.n311 VDD.n310 3.1505
R330 VDD.n310 VDD.n309 3.1505
R331 VDD.n314 VDD.n313 3.1505
R332 VDD.n313 VDD.n312 3.1505
R333 VDD.n317 VDD.n316 3.1505
R334 VDD.n316 VDD.n315 3.1505
R335 VDD.n320 VDD.n319 3.1505
R336 VDD.n319 VDD.n318 3.1505
R337 VDD.n323 VDD.n322 3.1505
R338 VDD.n322 VDD.n321 3.1505
R339 VDD.n326 VDD.n325 3.1505
R340 VDD.n325 VDD.n324 3.1505
R341 VDD.n329 VDD.n328 3.1505
R342 VDD.n328 VDD.n327 3.1505
R343 VDD.n332 VDD.n331 3.1505
R344 VDD.n331 VDD.n330 3.1505
R345 VDD.n335 VDD.n334 3.1505
R346 VDD.n334 VDD.n333 3.1505
R347 VDD.n338 VDD.n337 3.1505
R348 VDD.n337 VDD.n336 3.1505
R349 VDD.n341 VDD.n340 3.1505
R350 VDD.n340 VDD.n339 3.1505
R351 VDD.n344 VDD.n343 3.1505
R352 VDD.n343 VDD.n342 3.1505
R353 VDD.n347 VDD.n346 3.1505
R354 VDD.n346 VDD.n345 3.1505
R355 VDD.n350 VDD.n349 3.1505
R356 VDD.n349 VDD.n348 3.1505
R357 VDD.n353 VDD.n352 3.1505
R358 VDD.n352 VDD.n351 3.1505
R359 VDD.n356 VDD.n355 3.1505
R360 VDD.n355 VDD.n354 3.1505
R361 VDD.n359 VDD.n358 3.1505
R362 VDD.n358 VDD.n357 3.1505
R363 VDD.n362 VDD.n361 3.1505
R364 VDD.n361 VDD.n360 3.1505
R365 VDD.n365 VDD.n364 3.1505
R366 VDD.n364 VDD.n363 3.1505
R367 VDD.n368 VDD.n367 3.1505
R368 VDD.n367 VDD.n366 3.1505
R369 VDD.n371 VDD.n370 3.1505
R370 VDD.n370 VDD.n369 3.1505
R371 VDD.n374 VDD.n373 3.1505
R372 VDD.n373 VDD.n372 3.1505
R373 VDD.n377 VDD.n376 3.1505
R374 VDD.n376 VDD.n375 3.1505
R375 VDD.n380 VDD.n379 3.1505
R376 VDD.n379 VDD.n378 3.1505
R377 VDD.n666 VDD.n665 3.1505
R378 VDD.n665 VDD.n664 3.1505
R379 VDD.n663 VDD.n662 3.1505
R380 VDD.n662 VDD.n661 3.1505
R381 VDD.n660 VDD.n659 3.1505
R382 VDD.n659 VDD.n658 3.1505
R383 VDD.n657 VDD.n656 3.1505
R384 VDD.n656 VDD.n655 3.1505
R385 VDD.n654 VDD.n653 3.1505
R386 VDD.n267 VDD.t10 2.53938
R387 VDD.n339 VDD.t17 2.53938
R388 VDD.n99 VDD.n98 2.40832
R389 VDD.n96 VDD.n95 2.40832
R390 VDD.n93 VDD.n92 2.40832
R391 VDD.n90 VDD.n89 2.40832
R392 VDD.n87 VDD.n86 2.40832
R393 VDD.n84 VDD.n83 2.40832
R394 VDD.n80 VDD.n79 2.40832
R395 VDD.n77 VDD.n76 2.40832
R396 VDD.n74 VDD.n73 2.40832
R397 VDD.n71 VDD.n70 2.40832
R398 VDD.n68 VDD.n67 2.40832
R399 VDD.n65 VDD.n64 2.40832
R400 VDD.n62 VDD.n61 2.40832
R401 VDD.n58 VDD.n57 2.40832
R402 VDD.n55 VDD.n54 2.40832
R403 VDD.n52 VDD.n51 2.40832
R404 VDD.n48 VDD.n47 2.40832
R405 VDD.n45 VDD.n44 2.40832
R406 VDD.n42 VDD.n41 2.40832
R407 VDD.n39 VDD.n38 2.40832
R408 VDD.n35 VDD.n34 2.40832
R409 VDD.n32 VDD.n31 2.40832
R410 VDD.n29 VDD.n28 2.40832
R411 VDD.n25 VDD.n24 2.40832
R412 VDD.n107 VDD.n103 1.94734
R413 VDD.n107 VDD.n104 1.94734
R414 VDD.n107 VDD.n105 1.94734
R415 VDD.n107 VDD.n106 1.94734
R416 VDD.n216 VDD.t15 1.90466
R417 VDD.n638 VDD.n637 1.74343
R418 VDD.n633 VDD.n632 1.74343
R419 VDD.n628 VDD.n627 1.74343
R420 VDD.n623 VDD.n622 1.74343
R421 VDD.n617 VDD.n616 1.74343
R422 VDD.n612 VDD.n611 1.74343
R423 VDD.n607 VDD.n606 1.74343
R424 VDD.n602 VDD.n601 1.74343
R425 VDD.n651 VDD.n650 1.7429
R426 VDD.n383 VDD.n382 1.6665
R427 VDD.n384 VDD.n383 1.66598
R428 VDD.n109 VDD.n108 1.42472
R429 VDD.n165 VDD.t16 1.26994
R430 VDD.n108 VDD.n107 1.15215
R431 VDD.n107 VDD.n102 1.15196
R432 VDD.n649 VDD.n648 0.705355
R433 VDD.n649 VDD.n647 0.705355
R434 VDD.n649 VDD.n646 0.705355
R435 VDD.n649 VDD.n645 0.705355
R436 VDD.n649 VDD.n644 0.705355
R437 VDD.n649 VDD.n643 0.705355
R438 VDD.n650 VDD.n649 0.705355
R439 VDD.n592 VDD.n591 0.481929
R440 VDD VDD.n668 0.365057
R441 VDD.n60 VDD.n0 0.361929
R442 VDD.n107 VDD.n101 0.31786
R443 VDD.n649 VDD.n642 0.31786
R444 VDD.n589 VDD.n587 0.173577
R445 VDD.n590 VDD.n589 0.1265
R446 VDD.n652 VDD.n641 0.0868265
R447 VDD.n641 VDD.n639 0.0868265
R448 VDD.n639 VDD.n636 0.0868265
R449 VDD.n636 VDD.n634 0.0868265
R450 VDD.n634 VDD.n631 0.0868265
R451 VDD.n631 VDD.n629 0.0868265
R452 VDD.n629 VDD.n626 0.0868265
R453 VDD.n626 VDD.n624 0.0868265
R454 VDD.n624 VDD.n621 0.0868265
R455 VDD.n618 VDD.n615 0.0868265
R456 VDD.n615 VDD.n613 0.0868265
R457 VDD.n613 VDD.n610 0.0868265
R458 VDD.n610 VDD.n608 0.0868265
R459 VDD.n608 VDD.n605 0.0868265
R460 VDD.n605 VDD.n603 0.0868265
R461 VDD.n603 VDD.n600 0.0868265
R462 VDD.n600 VDD.n598 0.0868265
R463 VDD.n598 VDD.n596 0.0868265
R464 VDD.n596 VDD.n594 0.0868265
R465 VDD.n584 VDD.n582 0.0868265
R466 VDD.n582 VDD.n580 0.0868265
R467 VDD.n580 VDD.n578 0.0868265
R468 VDD.n578 VDD.n576 0.0868265
R469 VDD.n576 VDD.n574 0.0868265
R470 VDD.n574 VDD.n572 0.0868265
R471 VDD.n572 VDD.n570 0.0868265
R472 VDD.n570 VDD.n568 0.0868265
R473 VDD.n568 VDD.n566 0.0868265
R474 VDD.n566 VDD.n564 0.0868265
R475 VDD.n10 VDD.n8 0.0868265
R476 VDD.n8 VDD.n6 0.0868265
R477 VDD.n6 VDD.n4 0.0868265
R478 VDD.n4 VDD.n2 0.0868265
R479 VDD.n388 VDD.n386 0.0868265
R480 VDD.n390 VDD.n388 0.0868265
R481 VDD.n392 VDD.n390 0.0868265
R482 VDD.n394 VDD.n392 0.0868265
R483 VDD.n396 VDD.n394 0.0868265
R484 VDD.n398 VDD.n396 0.0868265
R485 VDD.n400 VDD.n398 0.0868265
R486 VDD.n402 VDD.n400 0.0868265
R487 VDD.n404 VDD.n402 0.0868265
R488 VDD.n406 VDD.n404 0.0868265
R489 VDD.n408 VDD.n406 0.0868265
R490 VDD.n410 VDD.n408 0.0868265
R491 VDD.n412 VDD.n410 0.0868265
R492 VDD.n414 VDD.n412 0.0868265
R493 VDD.n416 VDD.n414 0.0868265
R494 VDD.n418 VDD.n416 0.0868265
R495 VDD.n420 VDD.n418 0.0868265
R496 VDD.n422 VDD.n420 0.0868265
R497 VDD.n424 VDD.n422 0.0868265
R498 VDD.n426 VDD.n424 0.0868265
R499 VDD.n428 VDD.n426 0.0868265
R500 VDD.n430 VDD.n428 0.0868265
R501 VDD.n432 VDD.n430 0.0868265
R502 VDD.n434 VDD.n432 0.0868265
R503 VDD.n436 VDD.n434 0.0868265
R504 VDD.n438 VDD.n436 0.0868265
R505 VDD.n440 VDD.n438 0.0868265
R506 VDD.n442 VDD.n440 0.0868265
R507 VDD.n444 VDD.n442 0.0868265
R508 VDD.n446 VDD.n444 0.0868265
R509 VDD.n448 VDD.n446 0.0868265
R510 VDD.n450 VDD.n448 0.0868265
R511 VDD.n452 VDD.n450 0.0868265
R512 VDD.n454 VDD.n452 0.0868265
R513 VDD.n456 VDD.n454 0.0868265
R514 VDD.n458 VDD.n456 0.0868265
R515 VDD.n460 VDD.n458 0.0868265
R516 VDD.n462 VDD.n460 0.0868265
R517 VDD.n464 VDD.n462 0.0868265
R518 VDD.n466 VDD.n464 0.0868265
R519 VDD.n468 VDD.n466 0.0868265
R520 VDD.n470 VDD.n468 0.0868265
R521 VDD.n472 VDD.n470 0.0868265
R522 VDD.n474 VDD.n472 0.0868265
R523 VDD.n476 VDD.n474 0.0868265
R524 VDD.n478 VDD.n476 0.0868265
R525 VDD.n480 VDD.n478 0.0868265
R526 VDD.n482 VDD.n480 0.0868265
R527 VDD.n484 VDD.n482 0.0868265
R528 VDD.n486 VDD.n484 0.0868265
R529 VDD.n488 VDD.n486 0.0868265
R530 VDD.n490 VDD.n488 0.0868265
R531 VDD.n492 VDD.n490 0.0868265
R532 VDD.n494 VDD.n492 0.0868265
R533 VDD.n496 VDD.n494 0.0868265
R534 VDD.n498 VDD.n496 0.0868265
R535 VDD.n500 VDD.n498 0.0868265
R536 VDD.n502 VDD.n500 0.0868265
R537 VDD.n504 VDD.n502 0.0868265
R538 VDD.n506 VDD.n504 0.0868265
R539 VDD.n508 VDD.n506 0.0868265
R540 VDD.n510 VDD.n508 0.0868265
R541 VDD.n512 VDD.n510 0.0868265
R542 VDD.n514 VDD.n512 0.0868265
R543 VDD.n516 VDD.n514 0.0868265
R544 VDD.n518 VDD.n516 0.0868265
R545 VDD.n520 VDD.n518 0.0868265
R546 VDD.n522 VDD.n520 0.0868265
R547 VDD.n524 VDD.n522 0.0868265
R548 VDD.n526 VDD.n524 0.0868265
R549 VDD.n528 VDD.n526 0.0868265
R550 VDD.n530 VDD.n528 0.0868265
R551 VDD.n532 VDD.n530 0.0868265
R552 VDD.n534 VDD.n532 0.0868265
R553 VDD.n536 VDD.n534 0.0868265
R554 VDD.n538 VDD.n536 0.0868265
R555 VDD.n540 VDD.n538 0.0868265
R556 VDD.n542 VDD.n540 0.0868265
R557 VDD.n544 VDD.n542 0.0868265
R558 VDD.n546 VDD.n544 0.0868265
R559 VDD.n548 VDD.n546 0.0868265
R560 VDD.n550 VDD.n548 0.0868265
R561 VDD.n552 VDD.n550 0.0868265
R562 VDD.n554 VDD.n552 0.0868265
R563 VDD.n559 VDD.n557 0.0868265
R564 VDD.n561 VDD.n559 0.0868265
R565 VDD.n563 VDD.n561 0.0868265
R566 VDD.n110 VDD.n100 0.0868265
R567 VDD.n100 VDD.n97 0.0868265
R568 VDD.n97 VDD.n94 0.0868265
R569 VDD.n94 VDD.n91 0.0868265
R570 VDD.n91 VDD.n88 0.0868265
R571 VDD.n88 VDD.n85 0.0868265
R572 VDD.n81 VDD.n78 0.0868265
R573 VDD.n78 VDD.n75 0.0868265
R574 VDD.n75 VDD.n72 0.0868265
R575 VDD.n72 VDD.n69 0.0868265
R576 VDD.n69 VDD.n66 0.0868265
R577 VDD.n66 VDD.n63 0.0868265
R578 VDD.n59 VDD.n56 0.0868265
R579 VDD.n56 VDD.n53 0.0868265
R580 VDD.n49 VDD.n46 0.0868265
R581 VDD.n46 VDD.n43 0.0868265
R582 VDD.n43 VDD.n40 0.0868265
R583 VDD.n36 VDD.n33 0.0868265
R584 VDD.n33 VDD.n30 0.0868265
R585 VDD.n26 VDD.n23 0.0868265
R586 VDD.n23 VDD.n21 0.0868265
R587 VDD.n21 VDD.n19 0.0868265
R588 VDD.n16 VDD.n14 0.0868265
R589 VDD.n14 VDD.n12 0.0868265
R590 VDD.n115 VDD.n112 0.0868265
R591 VDD.n118 VDD.n115 0.0868265
R592 VDD.n121 VDD.n118 0.0868265
R593 VDD.n124 VDD.n121 0.0868265
R594 VDD.n131 VDD.n128 0.0868265
R595 VDD.n134 VDD.n131 0.0868265
R596 VDD.n137 VDD.n134 0.0868265
R597 VDD.n140 VDD.n137 0.0868265
R598 VDD.n143 VDD.n140 0.0868265
R599 VDD.n146 VDD.n143 0.0868265
R600 VDD.n149 VDD.n146 0.0868265
R601 VDD.n152 VDD.n149 0.0868265
R602 VDD.n155 VDD.n152 0.0868265
R603 VDD.n158 VDD.n155 0.0868265
R604 VDD.n161 VDD.n158 0.0868265
R605 VDD.n164 VDD.n161 0.0868265
R606 VDD.n167 VDD.n164 0.0868265
R607 VDD.n170 VDD.n167 0.0868265
R608 VDD.n173 VDD.n170 0.0868265
R609 VDD.n176 VDD.n173 0.0868265
R610 VDD.n179 VDD.n176 0.0868265
R611 VDD.n182 VDD.n179 0.0868265
R612 VDD.n185 VDD.n182 0.0868265
R613 VDD.n188 VDD.n185 0.0868265
R614 VDD.n191 VDD.n188 0.0868265
R615 VDD.n194 VDD.n191 0.0868265
R616 VDD.n197 VDD.n194 0.0868265
R617 VDD.n200 VDD.n197 0.0868265
R618 VDD.n203 VDD.n200 0.0868265
R619 VDD.n206 VDD.n203 0.0868265
R620 VDD.n209 VDD.n206 0.0868265
R621 VDD.n212 VDD.n209 0.0868265
R622 VDD.n215 VDD.n212 0.0868265
R623 VDD.n218 VDD.n215 0.0868265
R624 VDD.n221 VDD.n218 0.0868265
R625 VDD.n224 VDD.n221 0.0868265
R626 VDD.n227 VDD.n224 0.0868265
R627 VDD.n230 VDD.n227 0.0868265
R628 VDD.n233 VDD.n230 0.0868265
R629 VDD.n236 VDD.n233 0.0868265
R630 VDD.n239 VDD.n236 0.0868265
R631 VDD.n242 VDD.n239 0.0868265
R632 VDD.n245 VDD.n242 0.0868265
R633 VDD.n248 VDD.n245 0.0868265
R634 VDD.n251 VDD.n248 0.0868265
R635 VDD.n254 VDD.n251 0.0868265
R636 VDD.n257 VDD.n254 0.0868265
R637 VDD.n260 VDD.n257 0.0868265
R638 VDD.n263 VDD.n260 0.0868265
R639 VDD.n266 VDD.n263 0.0868265
R640 VDD.n269 VDD.n266 0.0868265
R641 VDD.n272 VDD.n269 0.0868265
R642 VDD.n275 VDD.n272 0.0868265
R643 VDD.n278 VDD.n275 0.0868265
R644 VDD.n281 VDD.n278 0.0868265
R645 VDD.n284 VDD.n281 0.0868265
R646 VDD.n287 VDD.n284 0.0868265
R647 VDD.n290 VDD.n287 0.0868265
R648 VDD.n293 VDD.n290 0.0868265
R649 VDD.n296 VDD.n293 0.0868265
R650 VDD.n299 VDD.n296 0.0868265
R651 VDD.n302 VDD.n299 0.0868265
R652 VDD.n305 VDD.n302 0.0868265
R653 VDD.n308 VDD.n305 0.0868265
R654 VDD.n311 VDD.n308 0.0868265
R655 VDD.n314 VDD.n311 0.0868265
R656 VDD.n317 VDD.n314 0.0868265
R657 VDD.n320 VDD.n317 0.0868265
R658 VDD.n323 VDD.n320 0.0868265
R659 VDD.n326 VDD.n323 0.0868265
R660 VDD.n329 VDD.n326 0.0868265
R661 VDD.n332 VDD.n329 0.0868265
R662 VDD.n335 VDD.n332 0.0868265
R663 VDD.n338 VDD.n335 0.0868265
R664 VDD.n341 VDD.n338 0.0868265
R665 VDD.n344 VDD.n341 0.0868265
R666 VDD.n347 VDD.n344 0.0868265
R667 VDD.n350 VDD.n347 0.0868265
R668 VDD.n353 VDD.n350 0.0868265
R669 VDD.n356 VDD.n353 0.0868265
R670 VDD.n359 VDD.n356 0.0868265
R671 VDD.n362 VDD.n359 0.0868265
R672 VDD.n365 VDD.n362 0.0868265
R673 VDD.n368 VDD.n365 0.0868265
R674 VDD.n371 VDD.n368 0.0868265
R675 VDD.n374 VDD.n371 0.0868265
R676 VDD.n377 VDD.n374 0.0868265
R677 VDD.n380 VDD.n377 0.0868265
R678 VDD.n666 VDD.n663 0.0868265
R679 VDD.n663 VDD.n660 0.0868265
R680 VDD.n660 VDD.n657 0.0868265
R681 VDD.n657 VDD.n654 0.0868265
R682 VDD.n555 VDD.n384 0.0861626
R683 VDD.n621 VDD.n619 0.0813163
R684 VDD.n53 VDD.n50 0.0748878
R685 VDD.n30 VDD.n27 0.0712143
R686 VDD.n589 VDD.n588 0.0699286
R687 VDD.n128 VDD.n125 0.0601939
R688 VDD.n17 VDD.n16 0.0574388
R689 VDD.n592 VDD.n584 0.0537653
R690 VDD.n555 VDD.n554 0.0537653
R691 VDD.n37 VDD.n36 0.0519286
R692 VDD.n667 VDD.n380 0.0500918
R693 VDD.n60 VDD.n59 0.0473367
R694 VDD.n85 VDD.n82 0.0455
R695 VDD.n564 VDD.n563 0.0427449
R696 VDD.n654 VDD.n652 0.0427449
R697 VDD.n12 VDD.n10 0.0427449
R698 VDD.n112 VDD.n110 0.0427449
R699 VDD.n82 VDD.n81 0.0418265
R700 VDD.n63 VDD.n60 0.0399898
R701 VDD.n667 VDD.n666 0.0372347
R702 VDD.n40 VDD.n37 0.035398
R703 VDD.n594 VDD.n592 0.0335612
R704 VDD.n557 VDD.n555 0.0335612
R705 VDD.n19 VDD.n17 0.0298878
R706 VDD.n125 VDD.n124 0.0271327
R707 VDD.n27 VDD.n26 0.0161122
R708 VDD.n50 VDD.n49 0.0124388
R709 VDD.n586 VDD.n585 0.0111513
R710 VDD.n587 VDD.n586 0.00926768
R711 VDD.n591 VDD.n590 0.00764286
R712 VDD VDD.n667 0.00733544
R713 VDD.n619 VDD.n618 0.0060102
R714 a_7427_13890.t0 a_7427_13890.t1 12.9075
R715 a_6467_13588.t0 a_6467_13588.t1 13.0784
R716 a_8387_13238.t0 a_8387_13238.t1 11.4969
R717 a_8067_14892.t0 a_8067_14892.t1 12.3428
R718 a_8387_12936.t0 a_8387_12936.t1 12.8783
R719 a_9987_13890.t0 a_9987_13890.t1 12.6832
R720 a_9667_13588.t0 a_9667_13588.t1 12.3428
R721 A.n5 A.t1 6.008
R722 A.n0 A.t0 5.06153
R723 A.n1 A.t2 2.008
R724 A.n2 A.n1 1.67436
R725 A.n2 A.n0 1.12905
R726 A.n5 A.n4 0.2957
R727 A A.n5 0.0635
R728 A.n4 A.n3 0.0158409
R729 A.n4 A.n2 0.00989489
R730 a_10627_14542.t0 a_10627_14542.t1 12.3428
R731 a_9347_15194.t0 a_9347_15194.t1 13.0919
R732 a_10307_14892.t0 a_10307_14892.t1 12.269
R733 a_7107_14892.t0 a_7107_14892.t1 12.5042
R734 a_7427_14240.t0 a_7427_14240.t1 13.0955
R735 a_9987_13238.t0 a_9987_13238.t1 12.3428
R736 a_10307_12936.t0 a_10307_12936.t1 12.8783
R737 a_11907_13890.t0 a_11907_13890.t1 8.16893
R738 a_11587_13588.t0 a_11587_13588.t1 12.3428
R739 a_9667_14542.t0 a_9667_14542.t1 12.3428
R740 a_9987_14240.t0 a_9987_14240.t1 8.39018
R741 a_12547_15194.t0 a_12547_15194.t1 12.3428
R742 D.n0 D.t0 8.7261
R743 D.n0 D.t1 3.74328
R744 D D.n0 0.1814
R745 a_6787_15194.t0 a_6787_15194.t1 12.3428
R746 a_12547_12936.t0 a_12547_12936.t1 12.3428
R747 G G.t3 6.8171
R748 G.n0 G.t2 6.29266
R749 G.n1 G.t1 6.116
R750 G.n0 G.t0 6.008
R751 G G.n1 4.48949
R752 G.n1 G.n0 0.117026
R753 a_6467_14240.t0 a_6467_14240.t1 10.61
R754 a_7107_13238.t0 a_7107_13238.t1 13.4549
R755 a_6787_12936.t0 a_6787_12936.t1 12.3428
R756 a_10947_13890.t0 a_10947_13890.t1 10.611
R757 a_10627_13588.t0 a_10627_13588.t1 12.3428
R758 a_8067_14240.t0 a_8067_14240.t1 10.6102
R759 a_8707_13588.t0 a_8707_13588.t1 12.3428
R760 a_9667_15194.t0 a_9667_15194.t1 12.3428
R761 a_9347_13890.t0 a_9347_13890.t1 8.7002
R762 a_9347_13238.t0 a_9347_13238.t1 12.3428
R763 a_9667_12936.t0 a_9667_12936.t1 12.3428
R764 a_7107_14240.t0 a_7107_14240.t1 8.16961
R765 a_7747_13588.t0 a_7747_13588.t1 12.3428
R766 a_11587_14542.t0 a_11587_14542.t1 12.3428
R767 a_11907_14240.t0 a_11907_14240.t1 10.6123
R768 a_11267_13890.t0 a_11267_13890.t1 12.9075
R769 a_12227_13588.t0 a_12227_13588.t1 13.0784
R770 B.n6 B.t0 6.16
R771 B.n5 B.t1 6.0089
R772 B.n2 B.t3 4.95996
R773 B.n0 B.t2 2.008
R774 B.n1 B.n0 1.67431
R775 B.n3 B.n2 1.13153
R776 B.n5 B.n4 0.2948
R777 B.n6 B.n5 0.1175
R778 B B.n6 0.0355
R779 B.n4 B.n3 0.0158409
R780 B.n4 B.n1 0.00989506
R781 a_11907_13238.t0 a_11907_13238.t1 12.269
R782 H.n0 H.t2 6.29675
R783 H.n1 H.t1 6.11695
R784 H.n0 H.t0 6.008
R785 H H.n1 0.495974
R786 H.n1 H.n0 0.116079
R787 a_12227_12936.t0 a_12227_12936.t1 12.8783
R788 E.n6 E.t0 6.74076
R789 E.n7 E.t4 6.1187
R790 E.n5 E.t1 6.10756
R791 E.n6 E.t3 6.008
R792 E.n0 E.t5 4.7503
R793 E.n1 E.t2 2.008
R794 E.n2 E.n1 1.67429
R795 E.n2 E.n0 1.1377
R796 E E.n7 1.0166
R797 E E.n5 0.4658
R798 E.n5 E.n4 0.1085
R799 E.n7 E.n6 0.0779
R800 E.n4 E.n3 0.0178864
R801 E.n4 E.n2 0.0087093
R802 a_6787_13588.t0 a_6787_13588.t1 12.3428
R803 a_10947_14240.t0 a_10947_14240.t1 8.16961
R804 a_8707_14542.t0 a_8707_14542.t1 12.3428
R805 a_8067_13890.t0 a_8067_13890.t1 8.16868
R806 a_10307_13588.t0 a_10307_13588.t1 13.0784
R807 a_9027_13890.t0 a_9027_13890.t1 8.38962
R808 a_7747_14542.t0 a_7747_14542.t1 12.3428
R809 a_7107_13890.t0 a_7107_13890.t1 10.611
R810 a_10627_15194.t0 a_10627_15194.t1 12.3428
R811 a_9027_14892.t0 a_9027_14892.t1 9.5196
R812 a_10307_14240.t0 a_10307_14240.t1 10.6105
R813 a_10627_12936.t0 a_10627_12936.t1 12.3428
R814 a_12227_14542.t0 a_12227_14542.t1 12.5042
R815 a_11267_14240.t0 a_11267_14240.t1 13.0955
R816 a_7427_13238.t0 a_7427_13238.t1 11.4973
R817 a_7427_14892.t0 a_7427_14892.t1 12.3428
R818 a_6787_14542.t0 a_6787_14542.t1 12.3428
R819 a_6467_12936.t0 a_6467_12936.t1 12.8783
R820 a_10947_14892.t0 a_10947_14892.t1 12.5042
R821 a_9027_14240.t0 a_9027_14240.t1 12.6832
R822 a_9987_14892.t0 a_9987_14892.t1 8.6992
R823 C.n0 C.t0 6.5003
R824 C.n0 C.t1 6.008
R825 C C.n0 0.0716
R826 a_6467_14892.t0 a_6467_14892.t1 12.268
R827 a_12867_14240.t0 a_12867_14240.t1 12.6832
R828 a_12547_13588.t0 a_12547_13588.t1 12.3428
R829 a_11587_15194.t0 a_11587_15194.t1 12.3428
R830 a_11907_14892.t0 a_11907_14892.t1 12.3428
R831 a_11587_12936.t0 a_11587_12936.t1 12.3428
R832 a_8387_13588.t0 a_8387_13588.t1 13.0784
R833 a_12867_13890.t0 a_12867_13890.t1 8.38962
R834 a_8707_15194.t0 a_8707_15194.t1 12.3428
R835 a_8387_14542.t0 a_8387_14542.t1 12.5042
R836 a_10947_13238.t0 a_10947_13238.t1 13.4549
R837 a_8707_12936.t0 a_8707_12936.t1 12.3428
R838 a_12547_14542.t0 a_12547_14542.t1 12.3428
R839 a_7747_15194.t0 a_7747_15194.t1 12.3428
R840 a_7747_12936.t0 a_7747_12936.t1 12.3428
R841 a_9347_14542.t0 a_9347_14542.t1 13.0703
R842 a_9027_13238.t0 a_9027_13238.t1 10.6105
R843 a_12227_13238.t0 a_12227_13238.t1 11.4969
R844 a_11267_13238.t0 a_11267_13238.t1 11.497
R845 a_11267_14892.t0 a_11267_14892.t1 12.3428
R846 a_8067_13238.t0 a_8067_13238.t1 12.269
C0 VDD E 3.08f
C1 VDD F 1.96f
C2 A G 0.302f
C3 C E 0.00425f
C4 B H 1.57e-20
C5 VDD C 0.444f
C6 D H 3.48e-19
C7 D B 0.395f
C8 E G 0.472f
C9 VDD G 2.72f
C10 A E 0.921f
C11 F H 0.0598f
C12 VDD H 1.22f
C13 C G 5.14e-20
C14 B F 0.278f
C15 VDD A 0.863f
C16 D F 0.355f
C17 VDD B 1.1f
C18 VDD D 0.805f
C19 A C 0.113f
C20 H VSUBS 0.291f
C21 F VSUBS 0.371f
C22 G VSUBS 1.78f
C23 E VSUBS 0.997f
C24 B VSUBS 0.408f
C25 D VSUBS 0.404f
C26 C VSUBS 0.227f
C27 A VSUBS 0.324f
C28 VDD VSUBS 90.1f
C29 E.t1 VSUBS 0.0909f
C30 E.t5 VSUBS 0.202f
C31 E.n0 VSUBS 0.752f
C32 E.t2 VSUBS 0.0375f
C33 E.n1 VSUBS 0.0786f
C34 E.n2 VSUBS 0.0202f
C35 E.n3 VSUBS 0.0196f
C36 E.n4 VSUBS 0.0556f
C37 E.n5 VSUBS 0.269f
C38 E.t0 VSUBS 0.114f
C39 E.t3 VSUBS 0.0898f
C40 E.n6 VSUBS 0.455f
C41 E.t4 VSUBS 0.0907f
C42 E.n7 VSUBS 0.4f
C43 G.t3 VSUBS 0.135f
C44 G.t2 VSUBS 0.108f
C45 G.t0 VSUBS 0.103f
C46 G.n0 VSUBS 0.252f
C47 G.t1 VSUBS 0.104f
C48 G.n1 VSUBS 0.873f
C49 VDD.t30 VSUBS 0.00343f
C50 VDD.t31 VSUBS 0.0035f
C51 VDD.t39 VSUBS 0.00332f
C52 VDD.t38 VSUBS 0.00363f
C53 VDD.n0 VSUBS 0.0101f
C54 VDD.t2 VSUBS 0.00361f
C55 VDD.t3 VSUBS 0.0036f
C56 VDD.t26 VSUBS 0.00346f
C57 VDD.t27 VSUBS 0.00361f
C58 VDD.n1 VSUBS 0.00124f
C59 VDD.n2 VSUBS 0.0016f
C60 VDD.n3 VSUBS 0.00124f
C61 VDD.n4 VSUBS 0.0016f
C62 VDD.n5 VSUBS 0.00124f
C63 VDD.n6 VSUBS 0.0016f
C64 VDD.n7 VSUBS 0.00124f
C65 VDD.n8 VSUBS 0.0016f
C66 VDD.n9 VSUBS 0.00149f
C67 VDD.n10 VSUBS 0.00201f
C68 VDD.n11 VSUBS 0.00101f
C69 VDD.n12 VSUBS 0.00121f
C70 VDD.n13 VSUBS 0.00124f
C71 VDD.n14 VSUBS 0.0016f
C72 VDD.n15 VSUBS 0.00124f
C73 VDD.n16 VSUBS 0.00133f
C74 VDD.n17 VSUBS 0.00637f
C75 VDD.n18 VSUBS 0.00124f
C76 VDD.n19 VSUBS 0.00107f
C77 VDD.n20 VSUBS 0.00124f
C78 VDD.n21 VSUBS 0.0016f
C79 VDD.n22 VSUBS 0.00124f
C80 VDD.n23 VSUBS 0.0016f
C81 VDD.n25 VSUBS 0.00124f
C82 VDD.n26 VSUBS 9.45e-19
C83 VDD.n27 VSUBS 0.0047f
C84 VDD.n29 VSUBS 0.00124f
C85 VDD.n30 VSUBS 0.00146f
C86 VDD.n32 VSUBS 0.00124f
C87 VDD.n33 VSUBS 0.0016f
C88 VDD.n35 VSUBS 0.00124f
C89 VDD.n36 VSUBS 0.00128f
C90 VDD.n37 VSUBS 0.00632f
C91 VDD.n39 VSUBS 0.00124f
C92 VDD.n40 VSUBS 0.00112f
C93 VDD.n42 VSUBS 0.00124f
C94 VDD.n43 VSUBS 0.0016f
C95 VDD.n45 VSUBS 0.00124f
C96 VDD.n46 VSUBS 0.0016f
C97 VDD.n48 VSUBS 0.00124f
C98 VDD.n49 VSUBS 9.11e-19
C99 VDD.n50 VSUBS 0.00634f
C100 VDD.n52 VSUBS 0.00124f
C101 VDD.n53 VSUBS 0.00149f
C102 VDD.n55 VSUBS 0.00124f
C103 VDD.n56 VSUBS 0.0016f
C104 VDD.n58 VSUBS 0.00124f
C105 VDD.n59 VSUBS 0.00123f
C106 VDD.n60 VSUBS 0.00219f
C107 VDD.n62 VSUBS 0.00124f
C108 VDD.n63 VSUBS 0.00117f
C109 VDD.n65 VSUBS 0.00124f
C110 VDD.n66 VSUBS 0.0016f
C111 VDD.n68 VSUBS 0.00124f
C112 VDD.n69 VSUBS 0.0016f
C113 VDD.n71 VSUBS 0.00124f
C114 VDD.n72 VSUBS 0.0016f
C115 VDD.n74 VSUBS 0.00124f
C116 VDD.n75 VSUBS 0.0016f
C117 VDD.n77 VSUBS 0.00124f
C118 VDD.n78 VSUBS 0.0016f
C119 VDD.n80 VSUBS 0.00124f
C120 VDD.n81 VSUBS 0.00118f
C121 VDD.n82 VSUBS 0.00431f
C122 VDD.n84 VSUBS 0.00124f
C123 VDD.n85 VSUBS 0.00122f
C124 VDD.n87 VSUBS 0.00124f
C125 VDD.n88 VSUBS 0.0016f
C126 VDD.n90 VSUBS 0.00124f
C127 VDD.n91 VSUBS 0.0016f
C128 VDD.n93 VSUBS 0.00124f
C129 VDD.n94 VSUBS 0.0016f
C130 VDD.n96 VSUBS 0.00124f
C131 VDD.n97 VSUBS 0.0016f
C132 VDD.n99 VSUBS 0.00124f
C133 VDD.n100 VSUBS 0.0016f
C134 VDD.n101 VSUBS 0.026f
C135 VDD.n107 VSUBS 0.0348f
C136 VDD.n109 VSUBS 0.00101f
C137 VDD.n110 VSUBS 0.00121f
C138 VDD.n111 VSUBS 0.00149f
C139 VDD.n112 VSUBS 0.00201f
C140 VDD.n113 VSUBS 0.0515f
C141 VDD.n114 VSUBS 0.00124f
C142 VDD.n115 VSUBS 0.0016f
C143 VDD.n116 VSUBS 0.0515f
C144 VDD.n117 VSUBS 0.00124f
C145 VDD.n118 VSUBS 0.0016f
C146 VDD.n119 VSUBS 0.0515f
C147 VDD.n120 VSUBS 0.00124f
C148 VDD.n121 VSUBS 0.0016f
C149 VDD.t1 VSUBS 0.0257f
C150 VDD.n122 VSUBS 0.0367f
C151 VDD.n123 VSUBS 0.00124f
C152 VDD.n124 VSUBS 0.00105f
C153 VDD.n125 VSUBS 0.00557f
C154 VDD.n126 VSUBS 0.0405f
C155 VDD.n127 VSUBS 0.00124f
C156 VDD.n128 VSUBS 0.00135f
C157 VDD.n129 VSUBS 0.0515f
C158 VDD.n130 VSUBS 0.00124f
C159 VDD.n131 VSUBS 0.0016f
C160 VDD.n132 VSUBS 0.0471f
C161 VDD.n133 VSUBS 0.00124f
C162 VDD.n134 VSUBS 0.0016f
C163 VDD.t13 VSUBS 0.0257f
C164 VDD.n135 VSUBS 0.0301f
C165 VDD.n136 VSUBS 0.00124f
C166 VDD.n137 VSUBS 0.0016f
C167 VDD.n138 VSUBS 0.0515f
C168 VDD.n139 VSUBS 0.00124f
C169 VDD.n140 VSUBS 0.0016f
C170 VDD.n141 VSUBS 0.0515f
C171 VDD.n142 VSUBS 0.00124f
C172 VDD.n143 VSUBS 0.0016f
C173 VDD.t8 VSUBS 0.0257f
C174 VDD.n144 VSUBS 0.0318f
C175 VDD.n145 VSUBS 0.00124f
C176 VDD.n146 VSUBS 0.0016f
C177 VDD.n147 VSUBS 0.0454f
C178 VDD.n148 VSUBS 0.00124f
C179 VDD.n149 VSUBS 0.0016f
C180 VDD.n150 VSUBS 0.0515f
C181 VDD.n151 VSUBS 0.00124f
C182 VDD.n152 VSUBS 0.0016f
C183 VDD.n153 VSUBS 0.0422f
C184 VDD.n154 VSUBS 0.00124f
C185 VDD.n155 VSUBS 0.0016f
C186 VDD.t14 VSUBS 0.0257f
C187 VDD.n156 VSUBS 0.035f
C188 VDD.n157 VSUBS 0.00124f
C189 VDD.n158 VSUBS 0.0016f
C190 VDD.n159 VSUBS 0.0515f
C191 VDD.n160 VSUBS 0.00124f
C192 VDD.n161 VSUBS 0.0016f
C193 VDD.n162 VSUBS 0.0515f
C194 VDD.n163 VSUBS 0.00124f
C195 VDD.n164 VSUBS 0.0016f
C196 VDD.t16 VSUBS 0.0257f
C197 VDD.n165 VSUBS 0.0268f
C198 VDD.n166 VSUBS 0.00124f
C199 VDD.n167 VSUBS 0.0016f
C200 VDD.n168 VSUBS 0.0504f
C201 VDD.n169 VSUBS 0.00124f
C202 VDD.n170 VSUBS 0.0016f
C203 VDD.n171 VSUBS 0.0515f
C204 VDD.n172 VSUBS 0.00124f
C205 VDD.n173 VSUBS 0.0016f
C206 VDD.t24 VSUBS 0.0257f
C207 VDD.n174 VSUBS 0.0372f
C208 VDD.n175 VSUBS 0.00124f
C209 VDD.n176 VSUBS 0.0016f
C210 VDD.n177 VSUBS 0.04f
C211 VDD.n178 VSUBS 0.00124f
C212 VDD.n179 VSUBS 0.0016f
C213 VDD.n180 VSUBS 0.0515f
C214 VDD.n181 VSUBS 0.00124f
C215 VDD.n182 VSUBS 0.0016f
C216 VDD.n183 VSUBS 0.0476f
C217 VDD.n184 VSUBS 0.00124f
C218 VDD.n185 VSUBS 0.0016f
C219 VDD.t12 VSUBS 0.0257f
C220 VDD.n186 VSUBS 0.0296f
C221 VDD.n187 VSUBS 0.00124f
C222 VDD.n188 VSUBS 0.0016f
C223 VDD.n189 VSUBS 0.0515f
C224 VDD.n190 VSUBS 0.00124f
C225 VDD.n191 VSUBS 0.0016f
C226 VDD.n192 VSUBS 0.0515f
C227 VDD.n193 VSUBS 0.00124f
C228 VDD.n194 VSUBS 0.0016f
C229 VDD.t9 VSUBS 0.0257f
C230 VDD.n195 VSUBS 0.0323f
C231 VDD.n196 VSUBS 0.00124f
C232 VDD.n197 VSUBS 0.0016f
C233 VDD.n198 VSUBS 0.0449f
C234 VDD.n199 VSUBS 0.00124f
C235 VDD.n200 VSUBS 0.0016f
C236 VDD.n201 VSUBS 0.0515f
C237 VDD.n202 VSUBS 0.00124f
C238 VDD.n203 VSUBS 0.0016f
C239 VDD.n204 VSUBS 0.0427f
C240 VDD.n205 VSUBS 0.00124f
C241 VDD.n206 VSUBS 0.0016f
C242 VDD.t29 VSUBS 0.0257f
C243 VDD.n207 VSUBS 0.0345f
C244 VDD.n208 VSUBS 0.00124f
C245 VDD.n209 VSUBS 0.0016f
C246 VDD.n210 VSUBS 0.0515f
C247 VDD.n211 VSUBS 0.00124f
C248 VDD.n212 VSUBS 0.0016f
C249 VDD.n213 VSUBS 0.0515f
C250 VDD.n214 VSUBS 0.00124f
C251 VDD.n215 VSUBS 0.0016f
C252 VDD.t15 VSUBS 0.0257f
C253 VDD.n216 VSUBS 0.0274f
C254 VDD.n217 VSUBS 0.00124f
C255 VDD.n218 VSUBS 0.0016f
C256 VDD.n219 VSUBS 0.0498f
C257 VDD.n220 VSUBS 0.00124f
C258 VDD.n221 VSUBS 0.0016f
C259 VDD.n222 VSUBS 0.0515f
C260 VDD.n223 VSUBS 0.00124f
C261 VDD.n224 VSUBS 0.0016f
C262 VDD.t23 VSUBS 0.0257f
C263 VDD.n225 VSUBS 0.0378f
C264 VDD.n226 VSUBS 0.00124f
C265 VDD.n227 VSUBS 0.0016f
C266 VDD.n228 VSUBS 0.0394f
C267 VDD.n229 VSUBS 0.00124f
C268 VDD.n230 VSUBS 0.0016f
C269 VDD.n231 VSUBS 0.0515f
C270 VDD.n232 VSUBS 0.00124f
C271 VDD.n233 VSUBS 0.0016f
C272 VDD.n234 VSUBS 0.0482f
C273 VDD.n235 VSUBS 0.00124f
C274 VDD.n236 VSUBS 0.0016f
C275 VDD.t22 VSUBS 0.0257f
C276 VDD.n237 VSUBS 0.029f
C277 VDD.n238 VSUBS 0.00124f
C278 VDD.n239 VSUBS 0.0016f
C279 VDD.n240 VSUBS 0.0515f
C280 VDD.n241 VSUBS 0.00124f
C281 VDD.n242 VSUBS 0.0016f
C282 VDD.n243 VSUBS 0.0515f
C283 VDD.n244 VSUBS 0.00124f
C284 VDD.n245 VSUBS 0.0016f
C285 VDD.t32 VSUBS 0.0257f
C286 VDD.n246 VSUBS 0.0329f
C287 VDD.n247 VSUBS 0.00124f
C288 VDD.n248 VSUBS 0.0016f
C289 VDD.n249 VSUBS 0.0444f
C290 VDD.n250 VSUBS 0.00124f
C291 VDD.n251 VSUBS 0.0016f
C292 VDD.n252 VSUBS 0.0515f
C293 VDD.n253 VSUBS 0.00124f
C294 VDD.n254 VSUBS 0.0016f
C295 VDD.n255 VSUBS 0.0433f
C296 VDD.n256 VSUBS 0.00124f
C297 VDD.n257 VSUBS 0.0016f
C298 VDD.t18 VSUBS 0.0257f
C299 VDD.n258 VSUBS 0.034f
C300 VDD.n259 VSUBS 0.00124f
C301 VDD.n260 VSUBS 0.0016f
C302 VDD.n261 VSUBS 0.0515f
C303 VDD.n262 VSUBS 0.00124f
C304 VDD.n263 VSUBS 0.0016f
C305 VDD.n264 VSUBS 0.0515f
C306 VDD.n265 VSUBS 0.00124f
C307 VDD.n266 VSUBS 0.0016f
C308 VDD.t10 VSUBS 0.0257f
C309 VDD.n267 VSUBS 0.0279f
C310 VDD.n268 VSUBS 0.00124f
C311 VDD.n269 VSUBS 0.0016f
C312 VDD.n270 VSUBS 0.0493f
C313 VDD.n271 VSUBS 0.00124f
C314 VDD.n272 VSUBS 0.0016f
C315 VDD.n273 VSUBS 0.0515f
C316 VDD.n274 VSUBS 0.00124f
C317 VDD.n275 VSUBS 0.0016f
C318 VDD.t33 VSUBS 0.0257f
C319 VDD.n276 VSUBS 0.0383f
C320 VDD.n277 VSUBS 0.00124f
C321 VDD.n278 VSUBS 0.0016f
C322 VDD.n279 VSUBS 0.0389f
C323 VDD.n280 VSUBS 0.00124f
C324 VDD.n281 VSUBS 0.0016f
C325 VDD.n282 VSUBS 0.0515f
C326 VDD.n283 VSUBS 0.00124f
C327 VDD.n284 VSUBS 0.0016f
C328 VDD.n285 VSUBS 0.0487f
C329 VDD.n286 VSUBS 0.00124f
C330 VDD.n287 VSUBS 0.0016f
C331 VDD.t20 VSUBS 0.0257f
C332 VDD.n288 VSUBS 0.0285f
C333 VDD.n289 VSUBS 0.00124f
C334 VDD.n290 VSUBS 0.0016f
C335 VDD.n291 VSUBS 0.0515f
C336 VDD.n292 VSUBS 0.00124f
C337 VDD.n293 VSUBS 0.0016f
C338 VDD.n294 VSUBS 0.0515f
C339 VDD.n295 VSUBS 0.00124f
C340 VDD.n296 VSUBS 0.0016f
C341 VDD.t4 VSUBS 0.0257f
C342 VDD.n297 VSUBS 0.0334f
C343 VDD.n298 VSUBS 0.00124f
C344 VDD.n299 VSUBS 0.0016f
C345 VDD.n300 VSUBS 0.0438f
C346 VDD.n301 VSUBS 0.00124f
C347 VDD.n302 VSUBS 0.0016f
C348 VDD.n303 VSUBS 0.0515f
C349 VDD.n304 VSUBS 0.00124f
C350 VDD.n305 VSUBS 0.0016f
C351 VDD.n306 VSUBS 0.0438f
C352 VDD.n307 VSUBS 0.00124f
C353 VDD.n308 VSUBS 0.0016f
C354 VDD.t21 VSUBS 0.0257f
C355 VDD.n309 VSUBS 0.0334f
C356 VDD.n310 VSUBS 0.00124f
C357 VDD.n311 VSUBS 0.0016f
C358 VDD.n312 VSUBS 0.0515f
C359 VDD.n313 VSUBS 0.00124f
C360 VDD.n314 VSUBS 0.0016f
C361 VDD.n315 VSUBS 0.0515f
C362 VDD.n316 VSUBS 0.00124f
C363 VDD.n317 VSUBS 0.0016f
C364 VDD.t25 VSUBS 0.0257f
C365 VDD.n318 VSUBS 0.0285f
C366 VDD.n319 VSUBS 0.00124f
C367 VDD.n320 VSUBS 0.0016f
C368 VDD.n321 VSUBS 0.0487f
C369 VDD.n322 VSUBS 0.00124f
C370 VDD.n323 VSUBS 0.0016f
C371 VDD.n324 VSUBS 0.0515f
C372 VDD.n325 VSUBS 0.00124f
C373 VDD.n326 VSUBS 0.0016f
C374 VDD.n327 VSUBS 0.0389f
C375 VDD.n328 VSUBS 0.00124f
C376 VDD.n329 VSUBS 0.0016f
C377 VDD.t28 VSUBS 0.0257f
C378 VDD.n330 VSUBS 0.0383f
C379 VDD.n331 VSUBS 0.00124f
C380 VDD.n332 VSUBS 0.0016f
C381 VDD.n333 VSUBS 0.0515f
C382 VDD.n334 VSUBS 0.00124f
C383 VDD.n335 VSUBS 0.0016f
C384 VDD.n336 VSUBS 0.0493f
C385 VDD.n337 VSUBS 0.00124f
C386 VDD.n338 VSUBS 0.0016f
C387 VDD.t17 VSUBS 0.0257f
C388 VDD.n339 VSUBS 0.0279f
C389 VDD.n340 VSUBS 0.00124f
C390 VDD.n341 VSUBS 0.0016f
C391 VDD.n342 VSUBS 0.0515f
C392 VDD.n343 VSUBS 0.00124f
C393 VDD.n344 VSUBS 0.0016f
C394 VDD.n345 VSUBS 0.0515f
C395 VDD.n346 VSUBS 0.00124f
C396 VDD.n347 VSUBS 0.0016f
C397 VDD.t0 VSUBS 0.0257f
C398 VDD.n348 VSUBS 0.034f
C399 VDD.n349 VSUBS 0.00124f
C400 VDD.n350 VSUBS 0.0016f
C401 VDD.n351 VSUBS 0.0433f
C402 VDD.n352 VSUBS 0.00124f
C403 VDD.n353 VSUBS 0.0016f
C404 VDD.n354 VSUBS 0.0515f
C405 VDD.n355 VSUBS 0.00124f
C406 VDD.n356 VSUBS 0.0016f
C407 VDD.n357 VSUBS 0.0444f
C408 VDD.n358 VSUBS 0.00124f
C409 VDD.n359 VSUBS 0.0016f
C410 VDD.t19 VSUBS 0.0257f
C411 VDD.n360 VSUBS 0.0329f
C412 VDD.n361 VSUBS 0.00124f
C413 VDD.n362 VSUBS 0.0016f
C414 VDD.n363 VSUBS 0.0515f
C415 VDD.n364 VSUBS 0.00124f
C416 VDD.n365 VSUBS 0.0016f
C417 VDD.n366 VSUBS 0.0515f
C418 VDD.n367 VSUBS 0.00124f
C419 VDD.n368 VSUBS 0.0016f
C420 VDD.t11 VSUBS 0.0257f
C421 VDD.n369 VSUBS 0.029f
C422 VDD.n370 VSUBS 0.00124f
C423 VDD.n371 VSUBS 0.0016f
C424 VDD.n372 VSUBS 0.0482f
C425 VDD.n373 VSUBS 0.00124f
C426 VDD.n374 VSUBS 0.0016f
C427 VDD.n375 VSUBS 0.0515f
C428 VDD.n376 VSUBS 0.00124f
C429 VDD.n377 VSUBS 0.0016f
C430 VDD.n378 VSUBS 0.0394f
C431 VDD.n379 VSUBS 0.00124f
C432 VDD.n380 VSUBS 0.00126f
C433 VDD.t40 VSUBS 0.00349f
C434 VDD.n381 VSUBS 0.00149f
C435 VDD.t7 VSUBS 0.00332f
C436 VDD.t41 VSUBS 0.00331f
C437 VDD.t34 VSUBS 0.00331f
C438 VDD.n382 VSUBS 0.0095f
C439 VDD.n383 VSUBS 0.0277f
C440 VDD.n384 VSUBS 0.00853f
C441 VDD.n385 VSUBS 0.00124f
C442 VDD.n386 VSUBS 0.0016f
C443 VDD.n387 VSUBS 0.00124f
C444 VDD.n388 VSUBS 0.0016f
C445 VDD.n389 VSUBS 0.00124f
C446 VDD.n390 VSUBS 0.0016f
C447 VDD.n391 VSUBS 0.00124f
C448 VDD.n392 VSUBS 0.0016f
C449 VDD.n393 VSUBS 0.00124f
C450 VDD.n394 VSUBS 0.0016f
C451 VDD.n395 VSUBS 0.00124f
C452 VDD.n396 VSUBS 0.0016f
C453 VDD.n397 VSUBS 0.00124f
C454 VDD.n398 VSUBS 0.0016f
C455 VDD.n399 VSUBS 0.00124f
C456 VDD.n400 VSUBS 0.0016f
C457 VDD.n401 VSUBS 0.00124f
C458 VDD.n402 VSUBS 0.0016f
C459 VDD.n403 VSUBS 0.00124f
C460 VDD.n404 VSUBS 0.0016f
C461 VDD.n405 VSUBS 0.00124f
C462 VDD.n406 VSUBS 0.0016f
C463 VDD.n407 VSUBS 0.00124f
C464 VDD.n408 VSUBS 0.0016f
C465 VDD.n409 VSUBS 0.00124f
C466 VDD.n410 VSUBS 0.0016f
C467 VDD.n411 VSUBS 0.00124f
C468 VDD.n412 VSUBS 0.0016f
C469 VDD.n413 VSUBS 0.00124f
C470 VDD.n414 VSUBS 0.0016f
C471 VDD.n415 VSUBS 0.00124f
C472 VDD.n416 VSUBS 0.0016f
C473 VDD.n417 VSUBS 0.00124f
C474 VDD.n418 VSUBS 0.0016f
C475 VDD.n419 VSUBS 0.00124f
C476 VDD.n420 VSUBS 0.0016f
C477 VDD.n421 VSUBS 0.00124f
C478 VDD.n422 VSUBS 0.0016f
C479 VDD.n423 VSUBS 0.00124f
C480 VDD.n424 VSUBS 0.0016f
C481 VDD.n425 VSUBS 0.00124f
C482 VDD.n426 VSUBS 0.0016f
C483 VDD.n427 VSUBS 0.00124f
C484 VDD.n428 VSUBS 0.0016f
C485 VDD.n429 VSUBS 0.00124f
C486 VDD.n430 VSUBS 0.0016f
C487 VDD.n431 VSUBS 0.00124f
C488 VDD.n432 VSUBS 0.0016f
C489 VDD.n433 VSUBS 0.00124f
C490 VDD.n434 VSUBS 0.0016f
C491 VDD.n435 VSUBS 0.00124f
C492 VDD.n436 VSUBS 0.0016f
C493 VDD.n437 VSUBS 0.00124f
C494 VDD.n438 VSUBS 0.0016f
C495 VDD.n439 VSUBS 0.00124f
C496 VDD.n440 VSUBS 0.0016f
C497 VDD.n441 VSUBS 0.00124f
C498 VDD.n442 VSUBS 0.0016f
C499 VDD.n443 VSUBS 0.00124f
C500 VDD.n444 VSUBS 0.0016f
C501 VDD.n445 VSUBS 0.00124f
C502 VDD.n446 VSUBS 0.0016f
C503 VDD.n447 VSUBS 0.00124f
C504 VDD.n448 VSUBS 0.0016f
C505 VDD.n449 VSUBS 0.00124f
C506 VDD.n450 VSUBS 0.0016f
C507 VDD.n451 VSUBS 0.00124f
C508 VDD.n452 VSUBS 0.0016f
C509 VDD.n453 VSUBS 0.00124f
C510 VDD.n454 VSUBS 0.0016f
C511 VDD.n455 VSUBS 0.00124f
C512 VDD.n456 VSUBS 0.0016f
C513 VDD.n457 VSUBS 0.00124f
C514 VDD.n458 VSUBS 0.0016f
C515 VDD.n459 VSUBS 0.00124f
C516 VDD.n460 VSUBS 0.0016f
C517 VDD.n461 VSUBS 0.00124f
C518 VDD.n462 VSUBS 0.0016f
C519 VDD.n463 VSUBS 0.00124f
C520 VDD.n464 VSUBS 0.0016f
C521 VDD.n465 VSUBS 0.00124f
C522 VDD.n466 VSUBS 0.0016f
C523 VDD.n467 VSUBS 0.00124f
C524 VDD.n468 VSUBS 0.0016f
C525 VDD.n469 VSUBS 0.00124f
C526 VDD.n470 VSUBS 0.0016f
C527 VDD.n471 VSUBS 0.00124f
C528 VDD.n472 VSUBS 0.0016f
C529 VDD.n473 VSUBS 0.00124f
C530 VDD.n474 VSUBS 0.0016f
C531 VDD.n475 VSUBS 0.00124f
C532 VDD.n476 VSUBS 0.0016f
C533 VDD.n477 VSUBS 0.00124f
C534 VDD.n478 VSUBS 0.0016f
C535 VDD.n479 VSUBS 0.00124f
C536 VDD.n480 VSUBS 0.0016f
C537 VDD.n481 VSUBS 0.00124f
C538 VDD.n482 VSUBS 0.0016f
C539 VDD.n483 VSUBS 0.00124f
C540 VDD.n484 VSUBS 0.0016f
C541 VDD.n485 VSUBS 0.00124f
C542 VDD.n486 VSUBS 0.0016f
C543 VDD.n487 VSUBS 0.00124f
C544 VDD.n488 VSUBS 0.0016f
C545 VDD.n489 VSUBS 0.00124f
C546 VDD.n490 VSUBS 0.0016f
C547 VDD.n491 VSUBS 0.00124f
C548 VDD.n492 VSUBS 0.0016f
C549 VDD.n493 VSUBS 0.00124f
C550 VDD.n494 VSUBS 0.0016f
C551 VDD.n495 VSUBS 0.00124f
C552 VDD.n496 VSUBS 0.0016f
C553 VDD.n497 VSUBS 0.00124f
C554 VDD.n498 VSUBS 0.0016f
C555 VDD.n499 VSUBS 0.00124f
C556 VDD.n500 VSUBS 0.0016f
C557 VDD.n501 VSUBS 0.00124f
C558 VDD.n502 VSUBS 0.0016f
C559 VDD.n503 VSUBS 0.00124f
C560 VDD.n504 VSUBS 0.0016f
C561 VDD.n505 VSUBS 0.00124f
C562 VDD.n506 VSUBS 0.0016f
C563 VDD.n507 VSUBS 0.00124f
C564 VDD.n508 VSUBS 0.0016f
C565 VDD.n509 VSUBS 0.00124f
C566 VDD.n510 VSUBS 0.0016f
C567 VDD.n511 VSUBS 0.00124f
C568 VDD.n512 VSUBS 0.0016f
C569 VDD.n513 VSUBS 0.00124f
C570 VDD.n514 VSUBS 0.0016f
C571 VDD.n515 VSUBS 0.00124f
C572 VDD.n516 VSUBS 0.0016f
C573 VDD.n517 VSUBS 0.00124f
C574 VDD.n518 VSUBS 0.0016f
C575 VDD.n519 VSUBS 0.00124f
C576 VDD.n520 VSUBS 0.0016f
C577 VDD.n521 VSUBS 0.00124f
C578 VDD.n522 VSUBS 0.0016f
C579 VDD.n523 VSUBS 0.00124f
C580 VDD.n524 VSUBS 0.0016f
C581 VDD.n525 VSUBS 0.00124f
C582 VDD.n526 VSUBS 0.0016f
C583 VDD.n527 VSUBS 0.00124f
C584 VDD.n528 VSUBS 0.0016f
C585 VDD.n529 VSUBS 0.00124f
C586 VDD.n530 VSUBS 0.0016f
C587 VDD.n531 VSUBS 0.00124f
C588 VDD.n532 VSUBS 0.0016f
C589 VDD.n533 VSUBS 0.00124f
C590 VDD.n534 VSUBS 0.0016f
C591 VDD.n535 VSUBS 0.00124f
C592 VDD.n536 VSUBS 0.0016f
C593 VDD.n537 VSUBS 0.00124f
C594 VDD.n538 VSUBS 0.0016f
C595 VDD.n539 VSUBS 0.00124f
C596 VDD.n540 VSUBS 0.0016f
C597 VDD.n541 VSUBS 0.00124f
C598 VDD.n542 VSUBS 0.0016f
C599 VDD.n543 VSUBS 0.00124f
C600 VDD.n544 VSUBS 0.0016f
C601 VDD.n545 VSUBS 0.00124f
C602 VDD.n546 VSUBS 0.0016f
C603 VDD.n547 VSUBS 0.00124f
C604 VDD.n548 VSUBS 0.0016f
C605 VDD.n549 VSUBS 0.00124f
C606 VDD.n550 VSUBS 0.0016f
C607 VDD.n551 VSUBS 0.00124f
C608 VDD.n552 VSUBS 0.0016f
C609 VDD.n553 VSUBS 0.00124f
C610 VDD.n554 VSUBS 0.00129f
C611 VDD.n555 VSUBS 0.00137f
C612 VDD.n556 VSUBS 0.00124f
C613 VDD.n557 VSUBS 0.00111f
C614 VDD.n558 VSUBS 0.00124f
C615 VDD.n559 VSUBS 0.0016f
C616 VDD.n560 VSUBS 0.00124f
C617 VDD.n561 VSUBS 0.0016f
C618 VDD.n562 VSUBS 0.00124f
C619 VDD.n563 VSUBS 0.00119f
C620 VDD.n564 VSUBS 0.00203f
C621 VDD.n565 VSUBS 0.00101f
C622 VDD.n566 VSUBS 0.0016f
C623 VDD.n567 VSUBS 0.00124f
C624 VDD.n568 VSUBS 0.0016f
C625 VDD.n569 VSUBS 0.00124f
C626 VDD.n570 VSUBS 0.0016f
C627 VDD.n571 VSUBS 0.00124f
C628 VDD.n572 VSUBS 0.0016f
C629 VDD.n573 VSUBS 0.00124f
C630 VDD.n574 VSUBS 0.0016f
C631 VDD.n575 VSUBS 0.00124f
C632 VDD.n576 VSUBS 0.0016f
C633 VDD.n577 VSUBS 0.00124f
C634 VDD.n578 VSUBS 0.0016f
C635 VDD.n579 VSUBS 0.00124f
C636 VDD.n580 VSUBS 0.0016f
C637 VDD.n581 VSUBS 0.00124f
C638 VDD.n582 VSUBS 0.0016f
C639 VDD.n583 VSUBS 0.00124f
C640 VDD.n584 VSUBS 0.00129f
C641 VDD.t35 VSUBS 0.00329f
C642 VDD.t6 VSUBS 0.00335f
C643 VDD.n585 VSUBS 0.00152f
C644 VDD.n586 VSUBS 0.00247f
C645 VDD.n587 VSUBS 0.00239f
C646 VDD.n588 VSUBS 4.7e-19
C647 VDD.n589 VSUBS 4.02e-19
C648 VDD.n590 VSUBS 0.00131f
C649 VDD.n591 VSUBS 0.00191f
C650 VDD.n592 VSUBS 0.00265f
C651 VDD.n593 VSUBS 0.00124f
C652 VDD.n594 VSUBS 0.00111f
C653 VDD.n595 VSUBS 0.00124f
C654 VDD.n596 VSUBS 0.0016f
C655 VDD.n597 VSUBS 0.00124f
C656 VDD.n598 VSUBS 0.0016f
C657 VDD.n599 VSUBS 0.00124f
C658 VDD.n600 VSUBS 0.0016f
C659 VDD.n602 VSUBS 0.00124f
C660 VDD.n603 VSUBS 0.0016f
C661 VDD.n604 VSUBS 0.00124f
C662 VDD.n605 VSUBS 0.0016f
C663 VDD.n607 VSUBS 0.00124f
C664 VDD.n608 VSUBS 0.0016f
C665 VDD.n609 VSUBS 0.00124f
C666 VDD.n610 VSUBS 0.0016f
C667 VDD.n612 VSUBS 0.00124f
C668 VDD.n613 VSUBS 0.0016f
C669 VDD.n614 VSUBS 0.00124f
C670 VDD.n615 VSUBS 0.0016f
C671 VDD.n617 VSUBS 0.00124f
C672 VDD.n618 VSUBS 8.52e-19
C673 VDD.n619 VSUBS 0.0041f
C674 VDD.n620 VSUBS 0.00124f
C675 VDD.n621 VSUBS 0.00155f
C676 VDD.n623 VSUBS 0.00124f
C677 VDD.n624 VSUBS 0.0016f
C678 VDD.n625 VSUBS 0.00124f
C679 VDD.n626 VSUBS 0.0016f
C680 VDD.n628 VSUBS 0.00124f
C681 VDD.n629 VSUBS 0.0016f
C682 VDD.n630 VSUBS 0.00124f
C683 VDD.n631 VSUBS 0.0016f
C684 VDD.n633 VSUBS 0.00124f
C685 VDD.n634 VSUBS 0.0016f
C686 VDD.n635 VSUBS 0.00124f
C687 VDD.n636 VSUBS 0.0016f
C688 VDD.n638 VSUBS 0.00124f
C689 VDD.n639 VSUBS 0.0016f
C690 VDD.n640 VSUBS 0.00124f
C691 VDD.n641 VSUBS 0.0016f
C692 VDD.n642 VSUBS 0.026f
C693 VDD.n649 VSUBS 0.0441f
C694 VDD.n651 VSUBS 0.00101f
C695 VDD.n652 VSUBS 0.00121f
C696 VDD.n653 VSUBS 0.00149f
C697 VDD.n654 VSUBS 0.00201f
C698 VDD.n655 VSUBS 0.0515f
C699 VDD.n656 VSUBS 0.00124f
C700 VDD.n657 VSUBS 0.0016f
C701 VDD.n658 VSUBS 0.0515f
C702 VDD.n659 VSUBS 0.00124f
C703 VDD.n660 VSUBS 0.0016f
C704 VDD.n661 VSUBS 0.0515f
C705 VDD.n662 VSUBS 0.00124f
C706 VDD.n663 VSUBS 0.0016f
C707 VDD.t5 VSUBS 0.0257f
C708 VDD.n664 VSUBS 0.0378f
C709 VDD.n665 VSUBS 0.00124f
C710 VDD.n666 VSUBS 0.00114f
C711 VDD.n667 VSUBS 8.42e-19
C712 VDD.t36 VSUBS 0.00329f
C713 VDD.t37 VSUBS 0.00343f
C714 VDD.n668 VSUBS 0.00635f
.ends

