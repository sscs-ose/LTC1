magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2374 -2045 2374 2045
<< psubdiff >>
rect -374 23 374 45
rect -374 -23 -352 23
rect 352 -23 374 23
rect -374 -45 374 -23
<< psubdiffcont >>
rect -352 -23 352 23
<< metal1 >>
rect -363 23 363 34
rect -363 -23 -352 23
rect 352 -23 363 23
rect -363 -34 363 -23
<< end >>
