magic
tech gf180mcuC
magscale 1 10
timestamp 1700063835
<< nwell >>
rect -73266 61805 -58779 62054
rect -73258 58003 -58787 61805
rect -73258 57988 -59591 58003
rect -73258 57977 -72761 57988
rect -70093 57871 -68828 57988
rect -64256 57871 -62991 57988
rect -71203 11821 -71102 11883
rect -71733 11589 -71082 11821
<< nsubdiff >>
rect -73028 61775 -58932 61903
rect -73028 61655 -71678 61775
rect -73028 61098 -72827 61655
rect -73022 61059 -72827 61098
rect -72225 61250 -71678 61655
rect -71087 61250 -70778 61775
rect -70187 61250 -69878 61775
rect -69287 61250 -68978 61775
rect -68387 61250 -68078 61775
rect -67487 61250 -67178 61775
rect -66587 61250 -66278 61775
rect -65687 61250 -65378 61775
rect -64787 61250 -64478 61775
rect -63887 61250 -63578 61775
rect -62987 61250 -62678 61775
rect -62087 61250 -61778 61775
rect -61187 61250 -60878 61775
rect -60287 61250 -59978 61775
rect -59387 61250 -58932 61775
rect -72225 61098 -58932 61250
rect -72225 61059 -72072 61098
rect -73022 60637 -72072 61059
rect -73022 60041 -72854 60637
rect -72252 60041 -72072 60637
rect -73022 59751 -72072 60041
rect -73022 59155 -72860 59751
rect -72258 59155 -72072 59751
rect -73022 58810 -72072 59155
rect -73022 58214 -72860 58810
rect -72258 58214 -72072 58810
rect -73022 58109 -72072 58214
rect -59619 60975 -58932 61098
rect -59619 60450 -59558 60975
rect -58967 60450 -58932 60975
rect -59619 60122 -58932 60450
rect -59619 59597 -59570 60122
rect -58979 59597 -58932 60122
rect -59619 59364 -58932 59597
rect -59619 58839 -59576 59364
rect -58985 58839 -58932 59364
rect -59619 58677 -58932 58839
rect -59619 58152 -59576 58677
rect -58985 58152 -58932 58677
rect -59619 58114 -58932 58152
rect -71528 11733 -71386 11748
rect -71528 11633 -71510 11733
rect -71399 11633 -71386 11733
rect -71528 11617 -71386 11633
rect -71271 11735 -71129 11750
rect -71271 11635 -71253 11735
rect -71142 11635 -71129 11735
rect -71271 11619 -71129 11635
<< nsubdiffcont >>
rect -72827 61059 -72225 61655
rect -71678 61250 -71087 61775
rect -70778 61250 -70187 61775
rect -69878 61250 -69287 61775
rect -68978 61250 -68387 61775
rect -68078 61250 -67487 61775
rect -67178 61250 -66587 61775
rect -66278 61250 -65687 61775
rect -65378 61250 -64787 61775
rect -64478 61250 -63887 61775
rect -63578 61250 -62987 61775
rect -62678 61250 -62087 61775
rect -61778 61250 -61187 61775
rect -60878 61250 -60287 61775
rect -59978 61250 -59387 61775
rect -72854 60041 -72252 60637
rect -72860 59155 -72258 59751
rect -72860 58214 -72258 58810
rect -59558 60450 -58967 60975
rect -59570 59597 -58979 60122
rect -59576 58839 -58985 59364
rect -59576 58152 -58985 58677
rect -71510 11633 -71399 11733
rect -71253 11635 -71142 11735
<< polysilicon >>
rect -56814 21654 -56200 21754
rect -56300 21619 -56200 21654
rect -56300 21547 -56286 21619
rect -56214 21547 -56200 21619
rect -56300 21533 -56200 21547
rect -71355 12314 -71255 12332
rect -71355 12263 -71333 12314
rect -71275 12263 -71255 12314
rect -71559 12224 -71459 12243
rect -71559 12176 -71539 12224
rect -71480 12176 -71459 12224
rect -71559 12110 -71459 12176
rect -71355 12110 -71255 12263
rect -17915 9817 -17815 9831
rect -17915 9770 -17901 9817
rect -17829 9770 -17815 9817
rect -17915 9756 -17815 9770
<< polycontact >>
rect -56286 21547 -56214 21619
rect -71333 12263 -71275 12314
rect -71539 12176 -71480 12224
rect -17901 9770 -17829 9817
<< metal1 >>
rect -59631 61923 -58871 61933
rect -72080 61918 -58871 61923
rect -73185 61775 -58871 61918
rect -73185 61655 -71678 61775
rect -73185 61133 -72827 61655
rect -73186 61059 -72827 61133
rect -72225 61250 -71678 61655
rect -71087 61250 -70778 61775
rect -70187 61250 -69878 61775
rect -69287 61250 -68978 61775
rect -68387 61250 -68078 61775
rect -67487 61250 -67178 61775
rect -66587 61250 -66278 61775
rect -65687 61250 -65378 61775
rect -64787 61250 -64478 61775
rect -63887 61250 -63578 61775
rect -62987 61250 -62678 61775
rect -62087 61250 -61778 61775
rect -61187 61250 -60878 61775
rect -60287 61250 -59978 61775
rect -59387 61250 -58871 61775
rect -72225 61134 -58871 61250
rect -72225 61059 -72081 61134
rect -73186 60637 -72081 61059
rect -67448 60876 -67063 61134
rect -59631 60975 -58871 61134
rect -73186 60041 -72854 60637
rect -72252 60041 -72081 60637
rect -70993 60800 -61181 60876
rect -70993 60795 -66142 60800
rect -70993 60691 -66351 60795
rect -66237 60696 -66142 60795
rect -66028 60696 -61181 60800
rect -66237 60691 -61181 60696
rect -70993 60630 -61181 60691
rect -70993 60526 -66354 60630
rect -66240 60629 -61181 60630
rect -66240 60526 -66141 60629
rect -70993 60525 -66141 60526
rect -66027 60525 -61181 60629
rect -70993 60505 -61181 60525
rect -70992 60491 -61181 60505
rect -70991 60318 -70621 60491
rect -73186 59751 -72081 60041
rect -70542 60122 -70174 60418
rect -70091 60315 -69721 60491
rect -69641 60122 -69271 60419
rect -69193 60314 -68822 60491
rect -68737 60122 -68367 60421
rect -68291 60315 -67925 60491
rect -67839 60122 -67469 60425
rect -67389 60307 -67023 60491
rect -66948 60122 -66578 60425
rect -65154 60318 -64784 60491
rect -64705 60122 -64337 60418
rect -64254 60315 -63884 60491
rect -63804 60122 -63434 60419
rect -63356 60314 -62985 60491
rect -62900 60122 -62530 60421
rect -62454 60315 -62088 60491
rect -62002 60122 -61632 60425
rect -61552 60307 -61186 60491
rect -59631 60450 -59558 60975
rect -58967 60450 -58871 60975
rect -61111 60122 -60741 60425
rect -59631 60122 -58871 60450
rect -70542 60104 -60733 60122
rect -70542 60000 -66351 60104
rect -66237 60000 -66128 60104
rect -66014 60000 -60733 60104
rect -70542 59948 -60733 60000
rect -70542 59947 -66128 59948
rect -70542 59906 -66350 59947
rect -70540 59843 -66350 59906
rect -66236 59844 -66128 59947
rect -66014 59844 -60733 59948
rect -66236 59843 -60733 59844
rect -70540 59814 -60733 59843
rect -73186 59155 -72860 59751
rect -72258 59155 -72081 59751
rect -73186 58810 -72081 59155
rect -59631 59597 -59570 60122
rect -58979 59597 -58871 60122
rect -59631 59364 -58871 59597
rect -73186 58214 -72860 58810
rect -72258 58214 -72081 58810
rect -70990 58794 -61183 58981
rect -73186 58046 -72081 58214
rect -70991 58622 -61183 58794
rect -59631 58839 -59576 59364
rect -58985 58839 -58871 59364
rect -59631 58677 -58871 58839
rect -70991 58508 -61182 58622
rect -70991 57148 -70621 58508
rect -70541 58118 -70170 58316
rect -70090 58222 -69720 58508
rect -69638 58118 -69273 58317
rect -69191 58214 -68819 58508
rect -68743 58118 -68372 58320
rect -68292 58214 -67920 58508
rect -67842 58118 -67471 58320
rect -67391 58212 -67019 58508
rect -66941 58118 -66571 58313
rect -65154 58214 -64784 58508
rect -64704 58118 -64333 58316
rect -64253 58222 -63883 58508
rect -63801 58118 -63436 58317
rect -63354 58214 -62982 58508
rect -62906 58118 -62535 58320
rect -62455 58214 -62083 58508
rect -62005 58118 -61634 58320
rect -61554 58212 -61182 58508
rect -61104 58118 -60734 58313
rect -70545 58011 -60734 58118
rect -59631 58152 -59576 58677
rect -58985 58152 -58871 58677
rect -59631 58036 -58871 58152
rect -70550 57733 -60734 58011
rect -70228 57148 -69832 57733
rect -66381 57176 -65982 57186
rect -66381 57175 -66214 57176
rect -70991 57141 -70510 57148
rect -70991 57140 -70742 57141
rect -70991 57087 -70897 57140
rect -70844 57088 -70742 57140
rect -70689 57088 -70584 57141
rect -70531 57088 -70510 57141
rect -70844 57087 -70510 57088
rect -70991 57034 -70510 57087
rect -70991 56981 -70895 57034
rect -70842 57031 -70510 57034
rect -70842 56981 -70738 57031
rect -70991 56978 -70738 56981
rect -70685 56978 -70585 57031
rect -70532 56978 -70510 57031
rect -70991 56926 -70510 56978
rect -70991 56925 -70738 56926
rect -70991 56872 -70896 56925
rect -70843 56873 -70738 56925
rect -70685 56924 -70510 56926
rect -70685 56873 -70586 56924
rect -70843 56872 -70586 56873
rect -70991 56871 -70586 56872
rect -70533 56871 -70510 56924
rect -70991 56816 -70510 56871
rect -70991 56797 -70893 56816
rect -70909 56763 -70893 56797
rect -70840 56815 -70510 56816
rect -70840 56763 -70737 56815
rect -70909 56762 -70737 56763
rect -70684 56762 -70584 56815
rect -70531 56762 -70510 56815
rect -70909 56749 -70510 56762
rect -70228 57140 -69824 57148
rect -70228 57139 -70055 57140
rect -70228 57086 -70210 57139
rect -70157 57087 -70055 57139
rect -70002 57087 -69897 57140
rect -69844 57087 -69824 57140
rect -70157 57086 -69824 57087
rect -70228 57033 -69824 57086
rect -70228 56980 -70208 57033
rect -70155 57030 -69824 57033
rect -70155 56980 -70051 57030
rect -70228 56977 -70051 56980
rect -69998 56977 -69898 57030
rect -69845 56977 -69824 57030
rect -70228 56925 -69824 56977
rect -70228 56924 -70051 56925
rect -70228 56871 -70209 56924
rect -70156 56872 -70051 56924
rect -69998 56923 -69824 56925
rect -69998 56872 -69899 56923
rect -70156 56871 -69899 56872
rect -70228 56870 -69899 56871
rect -69846 56870 -69824 56923
rect -70228 56815 -69824 56870
rect -70228 56762 -70206 56815
rect -70153 56814 -69824 56815
rect -70153 56762 -70050 56814
rect -70228 56761 -70050 56762
rect -69997 56761 -69897 56814
rect -69844 56761 -69824 56814
rect -66381 57122 -66369 57175
rect -66316 57123 -66214 57175
rect -66161 57123 -66056 57176
rect -66003 57123 -65982 57176
rect -66316 57122 -65982 57123
rect -66381 57069 -65982 57122
rect -66381 57016 -66367 57069
rect -66314 57066 -65982 57069
rect -66314 57016 -66210 57066
rect -66381 57013 -66210 57016
rect -66157 57013 -66057 57066
rect -66004 57013 -65982 57066
rect -66381 56961 -65982 57013
rect -66381 56960 -66210 56961
rect -66381 56907 -66368 56960
rect -66315 56908 -66210 56960
rect -66157 56959 -65982 56961
rect -66157 56908 -66058 56959
rect -66315 56907 -66058 56908
rect -66381 56906 -66058 56907
rect -66005 56906 -65982 56959
rect -66381 56851 -65982 56906
rect -66381 56798 -66365 56851
rect -66312 56850 -65982 56851
rect -66312 56798 -66209 56850
rect -66381 56797 -66209 56798
rect -66156 56797 -66056 56850
rect -66003 56797 -65982 56850
rect -66381 56787 -65982 56797
rect -65695 57172 -65296 57182
rect -65695 57171 -65528 57172
rect -65695 57118 -65683 57171
rect -65630 57119 -65528 57171
rect -65475 57119 -65370 57172
rect -65317 57119 -65296 57172
rect -65630 57118 -65296 57119
rect -65695 57065 -65296 57118
rect -65695 57012 -65681 57065
rect -65628 57062 -65296 57065
rect -65628 57012 -65524 57062
rect -65695 57009 -65524 57012
rect -65471 57009 -65371 57062
rect -65318 57009 -65296 57062
rect -65695 56957 -65296 57009
rect -65695 56956 -65524 56957
rect -65695 56903 -65682 56956
rect -65629 56904 -65524 56956
rect -65471 56955 -65296 56957
rect -65471 56904 -65372 56955
rect -65629 56903 -65372 56904
rect -65695 56902 -65372 56903
rect -65319 56902 -65296 56955
rect -65695 56847 -65296 56902
rect -65695 56794 -65679 56847
rect -65626 56846 -65296 56847
rect -65626 56794 -65523 56846
rect -65695 56793 -65523 56794
rect -65470 56793 -65370 56846
rect -65317 56793 -65296 56846
rect -65695 56783 -65296 56793
rect -70228 56749 -69824 56761
rect -8574 56766 -8343 56775
rect -70228 56736 -69832 56749
rect -8574 56713 -8560 56766
rect -8508 56765 -8343 56766
rect -8508 56713 -8423 56765
rect -8574 56712 -8423 56713
rect -8371 56712 -8343 56765
rect -8574 56620 -8343 56712
rect -8574 56567 -8555 56620
rect -8503 56567 -8409 56620
rect -8357 56567 -8343 56620
rect -8574 56544 -8343 56567
rect -43768 52594 -43665 52615
rect -43768 52520 -43752 52594
rect -43678 52520 -43665 52594
rect -53949 52420 -53842 52442
rect -43768 52420 -43665 52520
rect 16644 52468 17105 52473
rect -4656 52461 -4553 52465
rect 6502 52461 6774 52463
rect 16644 52461 17106 52468
rect -4667 52450 16664 52461
rect -4667 52449 6516 52450
rect -32412 52424 -32065 52431
rect -18447 52424 -18336 52439
rect -32412 52423 -18336 52424
rect -32412 52420 -18434 52423
rect -53949 52416 -18434 52420
rect -53949 52415 -32393 52416
rect -53949 52343 -53932 52415
rect -53860 52343 -43752 52415
rect -53949 52341 -43752 52343
rect -43678 52342 -32393 52415
rect -32319 52342 -32152 52416
rect -32078 52342 -18434 52416
rect -43678 52341 -18434 52342
rect -53949 52339 -18434 52341
rect -53949 52194 -53842 52339
rect -43768 52323 -43665 52339
rect -32412 52336 -18434 52339
rect -18347 52336 -18336 52423
rect -4667 52373 -4639 52449
rect -4563 52373 6516 52449
rect -4667 52372 6516 52373
rect 6594 52372 6681 52450
rect 6759 52372 16664 52450
rect -4667 52362 16664 52372
rect 16763 52460 17106 52461
rect 16763 52363 16857 52460
rect 16954 52363 17106 52460
rect 16763 52362 17106 52363
rect -32412 52335 -18336 52336
rect -32412 52331 -32065 52335
rect -53949 52120 -53933 52194
rect -53859 52120 -53842 52194
rect -18447 52221 -18336 52335
rect -53949 52105 -53842 52120
rect -53685 52166 -53551 52183
rect -43467 52166 -43344 52179
rect -32652 52166 -32293 52180
rect -18790 52166 -18663 52181
rect -53685 52165 -32642 52166
rect -53685 52067 -53671 52165
rect -53573 52067 -43453 52165
rect -43355 52067 -32642 52165
rect -53685 52066 -32642 52067
rect -32542 52066 -32415 52166
rect -32315 52165 -18663 52166
rect -32315 52067 -18775 52165
rect -18677 52067 -18663 52165
rect -18447 52132 -18434 52221
rect -18345 52132 -18336 52221
rect -4656 52251 -4553 52362
rect 6502 52357 6774 52362
rect 16644 52348 17106 52362
rect -4656 52173 -4640 52251
rect -4562 52173 -4553 52251
rect -4656 52165 -4553 52173
rect -4381 52196 -4248 52213
rect 6356 52196 6489 52215
rect 17262 52196 17412 52214
rect -4381 52195 6370 52196
rect -18447 52117 -18336 52132
rect -32315 52066 -18663 52067
rect -53685 51987 -53551 52066
rect -53685 51887 -53672 51987
rect -53572 51887 -53551 51987
rect -53685 51877 -53551 51887
rect -43467 51951 -43344 52066
rect -32652 52052 -32293 52066
rect -43467 51851 -43454 51951
rect -43354 51851 -43344 51951
rect -43467 51842 -43344 51851
rect -18790 51928 -18663 52066
rect -18790 51828 -18776 51928
rect -18676 51828 -18663 51928
rect -4381 52090 -4366 52195
rect -4261 52090 6370 52195
rect -4381 52089 6370 52090
rect 6477 52195 17412 52196
rect 6477 52090 17284 52195
rect 17389 52090 17412 52195
rect 6477 52089 17412 52090
rect -4381 51970 -4248 52089
rect -4381 51863 -4366 51970
rect -4259 51863 -4248 51970
rect 6356 51989 6489 52089
rect 6356 51884 6371 51989
rect 6476 51884 6489 51989
rect 6356 51868 6489 51884
rect 17262 51993 17412 52089
rect 17262 51886 17283 51993
rect 17390 51886 17412 51993
rect 17262 51875 17412 51886
rect -4381 51851 -4248 51863
rect -32166 51817 -32065 51825
rect -32166 51743 -32152 51817
rect -32078 51743 -32065 51817
rect -18790 51814 -18663 51828
rect 6673 51771 6769 51780
rect -32166 51644 -32065 51743
rect 6672 51770 6769 51771
rect 6672 51692 6681 51770
rect 6759 51692 6769 51770
rect 6672 51691 6769 51692
rect -32166 51643 -30936 51644
rect -32166 51571 -32151 51643
rect -32079 51571 -30936 51643
rect 6673 51606 6769 51691
rect -32166 51570 -30936 51571
rect -32166 51556 -32065 51570
rect 6673 51530 6682 51606
rect 6758 51604 6977 51606
rect 6758 51530 7910 51604
rect 6673 51529 6977 51530
rect 6673 51518 6769 51529
rect -46054 51363 -40254 51388
rect -46054 51360 -44929 51363
rect -46130 51314 -44929 51360
rect -46054 51306 -44929 51314
rect -44876 51306 -44814 51363
rect -44761 51362 -40254 51363
rect -44761 51306 -44678 51362
rect -46054 51305 -44678 51306
rect -44625 51317 -40254 51362
rect 3146 51319 5233 51334
rect -44625 51305 -40024 51317
rect -46054 51287 -40024 51305
rect 3146 51316 5158 51319
rect -40355 51216 -40024 51287
rect -35684 51264 -34300 51278
rect -35684 51261 -34395 51264
rect -35684 51258 -34546 51261
rect -35684 51247 -34692 51258
rect -36151 51201 -34692 51247
rect -35684 51187 -34692 51201
rect -34618 51190 -34546 51258
rect -34472 51193 -34395 51261
rect -34321 51193 -34300 51264
rect -34472 51190 -34300 51193
rect -34618 51187 -34300 51190
rect -24775 51273 -15407 51288
rect -24775 51271 -23234 51273
rect -24775 51196 -23385 51271
rect -23314 51198 -23234 51271
rect -23163 51272 -15407 51273
rect -23163 51198 -23089 51272
rect -23314 51197 -23089 51198
rect -23018 51197 -15407 51272
rect -10856 51263 -1331 51277
rect -10856 51261 -6869 51263
rect -10856 51247 -7131 51261
rect -10939 51201 -7131 51247
rect -23314 51196 -15407 51197
rect -35684 51171 -34300 51187
rect -32439 51168 -32291 51188
rect -24775 51179 -15407 51196
rect -10856 51185 -7131 51201
rect -7078 51260 -6869 51261
rect -7078 51185 -7009 51260
rect -10856 51184 -7009 51185
rect -6956 51187 -6869 51260
rect -6816 51187 -1331 51263
rect 3146 51240 4845 51316
rect 4907 51315 5158 51316
rect 4907 51240 4973 51315
rect 3146 51239 4973 51240
rect 5035 51243 5158 51315
rect 5220 51243 5233 51319
rect 5035 51239 5233 51243
rect 3146 51227 5233 51239
rect 14057 51242 20405 51274
rect 24950 51265 26424 51278
rect 24950 51262 26325 51265
rect 24950 51260 26161 51262
rect 24950 51247 26024 51260
rect -6956 51184 -1331 51187
rect -10856 51171 -1331 51184
rect -32439 51057 -32421 51168
rect -32310 51057 -32291 51168
rect -1437 51095 -1331 51171
rect 14057 51153 15334 51242
rect 15395 51241 20405 51242
rect 15395 51153 15482 51241
rect 14057 51152 15482 51153
rect 15543 51152 15644 51241
rect 15705 51152 20405 51241
rect 24862 51201 26024 51247
rect 24950 51178 26024 51201
rect 26083 51180 26161 51260
rect 26220 51183 26325 51262
rect 26384 51183 26424 51265
rect 26220 51180 26424 51183
rect 26083 51178 26424 51180
rect 24950 51170 26424 51178
rect 6351 51129 6497 51144
rect 14057 51137 20405 51152
rect -32439 50943 -32291 51057
rect 6351 51018 6368 51129
rect 6479 51018 6497 51129
rect -32439 50942 -31553 50943
rect -32439 50833 -32421 50942
rect -32312 50833 -31553 50942
rect -32439 50832 -31553 50833
rect 6351 50903 6497 51018
rect 20268 51013 20405 51137
rect 6351 50902 7293 50903
rect -32439 50815 -32291 50832
rect 6351 50793 6369 50902
rect 6478 50793 7293 50902
rect 6351 50792 7293 50793
rect 6351 50772 6497 50792
rect -55956 50421 -52524 50479
rect -55956 50418 -55769 50421
rect -55956 50355 -55901 50418
rect -55841 50358 -55769 50418
rect -55709 50418 -52524 50421
rect -55709 50358 -55635 50418
rect -55841 50355 -55635 50358
rect -55575 50355 -52524 50418
rect -55956 50329 -52524 50355
rect -45765 50308 -42163 50366
rect -45765 50305 -45613 50308
rect -45765 50242 -45745 50305
rect -45685 50245 -45613 50305
rect -45553 50305 -42163 50308
rect -45553 50245 -45479 50305
rect -45685 50242 -45479 50245
rect -45419 50242 -42163 50305
rect -45765 50216 -42163 50242
rect -24201 50312 -17340 50366
rect -24201 50309 -24037 50312
rect -24201 50246 -24169 50309
rect -24109 50249 -24037 50309
rect -23977 50309 -17340 50312
rect -23977 50249 -23903 50309
rect -24109 50246 -23903 50249
rect -23843 50246 -17340 50309
rect -7921 50365 -3236 50422
rect -7921 50362 -7751 50365
rect -7921 50299 -7883 50362
rect -7823 50302 -7751 50362
rect -7691 50362 -3236 50365
rect -7691 50302 -7617 50362
rect -7823 50299 -7617 50302
rect -7557 50299 -3236 50362
rect -7921 50272 -3236 50299
rect 14637 50297 18484 50366
rect 14637 50294 14792 50297
rect -24201 50216 -17340 50246
rect 14637 50231 14660 50294
rect 14720 50234 14792 50294
rect 14852 50294 18484 50297
rect 14852 50234 14926 50294
rect 14720 50231 14926 50234
rect 14986 50231 18484 50294
rect 14637 50219 18484 50231
rect 14637 50216 14738 50219
rect 14912 50216 18484 50219
rect -53272 50091 -53149 50105
rect -53272 50012 -53252 50091
rect -53161 50012 -53149 50091
rect -53272 49977 -53149 50012
rect -50932 50009 -50767 50055
rect -3907 50004 -3784 50018
rect -42893 49984 -42770 49998
rect -53874 49939 -53043 49977
rect -53874 49895 -53256 49939
rect -53272 49860 -53256 49895
rect -53165 49895 -53043 49939
rect -42893 49905 -42873 49984
rect -42782 49914 -42770 49984
rect -17998 49967 -17875 49981
rect -42782 49905 -42723 49914
rect -53165 49860 -53149 49895
rect -42893 49864 -42723 49905
rect -17998 49888 -17978 49967
rect -17887 49888 -17875 49967
rect -3907 49925 -3887 50004
rect -3796 49925 -3784 50004
rect -1659 49952 -1449 49998
rect -3907 49920 -3784 49925
rect -17998 49864 -17875 49888
rect -53272 49848 -53149 49860
rect -43513 49832 -42682 49864
rect -43513 49782 -42877 49832
rect -42893 49753 -42877 49782
rect -42786 49782 -42682 49832
rect -18690 49815 -17859 49864
rect -4586 49852 -3755 49920
rect -4586 49838 -3891 49852
rect -18690 49782 -17982 49815
rect -42786 49762 -42723 49782
rect -42786 49760 -42728 49762
rect -42786 49753 -42770 49760
rect -42893 49741 -42770 49753
rect -17998 49736 -17982 49782
rect -17891 49782 -17859 49815
rect -17891 49736 -17875 49782
rect -3907 49773 -3891 49838
rect -3800 49838 -3755 49852
rect 16526 49916 16634 49968
rect 16526 49846 16552 49916
rect 16623 49864 16634 49916
rect 20074 49896 20246 49942
rect 16623 49846 17965 49864
rect -3800 49773 -3784 49838
rect -3907 49761 -3784 49773
rect 16526 49782 17965 49846
rect -17998 49724 -17875 49736
rect 16526 49745 16634 49782
rect 16526 49675 16549 49745
rect 16620 49675 16634 49745
rect 16526 49645 16634 49675
rect -66401 49625 -59425 49628
rect -67807 49606 -59425 49625
rect -67807 49599 -66090 49606
rect -67807 49597 -66220 49599
rect -67807 49539 -66361 49597
rect -66296 49541 -66220 49597
rect -66155 49548 -66090 49599
rect -66025 49548 -59425 49606
rect -66155 49541 -59425 49548
rect -66296 49539 -59425 49541
rect -67807 49514 -59425 49539
rect -67807 49511 -65978 49514
rect -71215 49251 -68664 49276
rect -71215 49170 -68599 49251
rect -71215 49145 -68664 49170
rect -67907 49140 -59442 49245
rect -57490 49231 -57438 49248
rect -58622 49184 -57438 49231
rect -67826 48920 -65272 48924
rect -67826 48887 -59420 48920
rect -67826 48885 -65393 48887
rect -67826 48827 -65668 48885
rect -65603 48883 -65393 48885
rect -65603 48827 -65525 48883
rect -67826 48825 -65525 48827
rect -65460 48829 -65393 48883
rect -65328 48829 -59420 48887
rect -65460 48825 -59420 48829
rect -67826 48810 -59420 48825
rect -65708 48806 -59420 48810
rect -67806 48140 -65978 48193
rect -67806 48120 -59368 48140
rect -67806 48079 -66365 48120
rect -66380 48062 -66365 48079
rect -66300 48119 -59368 48120
rect -66300 48062 -66223 48119
rect -66380 48061 -66223 48062
rect -66158 48061 -66078 48119
rect -66013 48061 -59368 48119
rect -66380 48026 -59368 48061
rect -71239 47823 -68636 47847
rect -71239 47742 -68600 47823
rect -71239 47717 -68636 47742
rect -67891 47710 -59412 47818
rect -57781 47738 -57735 47742
rect -58593 47691 -57735 47738
rect -67804 47418 -65272 47490
rect -67804 47416 -59372 47418
rect -67804 47415 -65377 47416
rect -67804 47376 -65661 47415
rect -65698 47357 -65661 47376
rect -65596 47412 -65377 47415
rect -65596 47357 -65522 47412
rect -65698 47354 -65522 47357
rect -65457 47358 -65377 47412
rect -65312 47358 -59372 47416
rect -65457 47354 -59372 47358
rect -65698 47304 -59372 47354
rect -67742 46683 -65978 46743
rect -67742 46663 -66086 46683
rect -67742 46654 -66232 46663
rect -67742 46629 -66365 46654
rect -66390 46596 -66365 46629
rect -66300 46605 -66232 46654
rect -66167 46625 -66086 46663
rect -66021 46662 -65978 46683
rect -66021 46625 -59294 46662
rect -66167 46605 -59294 46625
rect -66300 46596 -59294 46605
rect -66390 46548 -59294 46596
rect -71123 46378 -68594 46404
rect -71123 46297 -68542 46378
rect -71123 46270 -68594 46297
rect -67838 46266 -59384 46372
rect -58593 46218 -57999 46265
rect -67742 45969 -65278 46043
rect -67742 45960 -65383 45969
rect -67742 45959 -65526 45960
rect -67742 45929 -65667 45959
rect -65708 45901 -65667 45929
rect -65602 45902 -65526 45959
rect -65461 45911 -65383 45960
rect -65318 45965 -65278 45969
rect -65318 45911 -59252 45965
rect -65461 45902 -59252 45911
rect -65602 45901 -59252 45902
rect -65708 45851 -59252 45901
rect -68490 43508 -66212 43622
rect -66326 43301 -66212 43508
rect -66386 43235 -62472 43301
rect -66386 43230 -66069 43235
rect -66386 43148 -66357 43230
rect -66293 43225 -66069 43230
rect -66293 43148 -66216 43225
rect -66386 43143 -66216 43148
rect -66152 43153 -66069 43225
rect -66005 43153 -62472 43235
rect -66152 43143 -62472 43153
rect -66386 43110 -62472 43143
rect -58055 42986 -57999 46218
rect -69864 42955 -69744 42956
rect -69866 42878 -69260 42955
rect -67809 42944 -67621 42974
rect -69864 42137 -69744 42878
rect -67809 42874 -67772 42944
rect -67706 42874 -67621 42944
rect -67809 42856 -67621 42874
rect -66730 42896 -66440 42940
rect -58729 42930 -57999 42986
rect -66730 42860 -62813 42896
rect -66520 42852 -62813 42860
rect -66520 42756 -62654 42852
rect -57781 42832 -57735 47691
rect -58846 42786 -57735 42832
rect -66520 42713 -62813 42756
rect -57490 42697 -57438 49184
rect -54509 49008 -54387 49042
rect -54509 48965 -53039 49008
rect -54509 48888 -54492 48965
rect -54412 48934 -53039 48965
rect -43959 48973 -43868 48998
rect -54412 48888 -54387 48934
rect -54509 48777 -54387 48888
rect -54509 48700 -54492 48777
rect -54412 48700 -54387 48777
rect -54509 48667 -54387 48700
rect -43959 48913 -43940 48973
rect -43888 48913 -43868 48973
rect -4975 48951 -4851 49035
rect -4975 48936 -3751 48951
rect -43959 48895 -43868 48913
rect -43959 48854 -42678 48895
rect -19394 48895 -19274 48918
rect -43959 48794 -43938 48854
rect -43886 48821 -42678 48854
rect -19394 48853 -17855 48895
rect -43886 48794 -43868 48821
rect -43959 48666 -43868 48794
rect -19394 48785 -19370 48853
rect -19289 48821 -17855 48853
rect -4975 48861 -4950 48936
rect -4873 48877 -3751 48936
rect 15329 48912 15710 48942
rect 15329 48909 15482 48912
rect 15329 48895 15350 48909
rect -4873 48861 -4851 48877
rect -19289 48785 -19274 48821
rect -35401 48779 -31921 48785
rect -35401 48776 -35248 48779
rect -35401 48713 -35380 48776
rect -35320 48716 -35248 48776
rect -35188 48776 -31921 48779
rect -35188 48716 -35114 48776
rect -35320 48713 -35114 48716
rect -35054 48713 -31921 48776
rect -35401 48703 -31921 48713
rect -19394 48713 -19274 48785
rect -19394 48645 -19377 48713
rect -19296 48645 -19274 48713
rect -4975 48763 -4851 48861
rect 15316 48846 15350 48895
rect 15410 48849 15482 48909
rect 15542 48909 15710 48912
rect 15542 48849 15616 48909
rect 15410 48846 15616 48849
rect 15676 48895 15710 48909
rect 15676 48846 17969 48895
rect 15316 48821 17969 48846
rect -4975 48688 -4951 48763
rect -4874 48688 -4851 48763
rect -4975 48661 -4851 48688
rect 4067 48740 6925 48745
rect 4067 48737 4212 48740
rect 4067 48674 4080 48737
rect 4140 48677 4212 48737
rect 4272 48737 6925 48740
rect 4272 48677 4346 48737
rect 4140 48674 4346 48677
rect 4406 48674 6925 48737
rect 4067 48663 6925 48674
rect -19394 48623 -19274 48645
rect -10233 48139 -8342 48170
rect -10233 48136 -8419 48139
rect -55275 48051 -54901 48076
rect -55275 48048 -55127 48051
rect -55275 48036 -55259 48048
rect -55295 47985 -55259 48036
rect -55199 47988 -55127 48048
rect -55067 48048 -54901 48051
rect -55067 47988 -54993 48048
rect -55199 47985 -54993 47988
rect -54933 48036 -54901 48048
rect -10233 48039 -8564 48136
rect -8508 48042 -8419 48136
rect -8363 48042 -8342 48139
rect -8508 48039 -8342 48042
rect -54933 47985 -53043 48036
rect -55295 47958 -53043 47985
rect -10233 48021 -8342 48039
rect -44938 47938 -44557 47954
rect -44938 47935 -44783 47938
rect -44938 47923 -44915 47935
rect -44955 47872 -44915 47923
rect -44855 47875 -44783 47935
rect -44723 47935 -44557 47938
rect -44723 47875 -44649 47935
rect -44855 47872 -44649 47875
rect -44589 47923 -44557 47935
rect -23393 47933 -23006 47954
rect -23393 47930 -23249 47933
rect -23393 47923 -23381 47930
rect -44589 47872 -42682 47923
rect -44955 47845 -42682 47872
rect -23399 47867 -23381 47923
rect -23321 47870 -23249 47930
rect -23189 47930 -23006 47933
rect -23189 47870 -23115 47930
rect -23321 47867 -23115 47870
rect -23055 47923 -23006 47930
rect -23055 47867 -17859 47923
rect -23399 47845 -17859 47867
rect -44688 47760 -44588 47845
rect -55305 47672 -50656 47704
rect -55305 47669 -55139 47672
rect -55305 47606 -55271 47669
rect -55211 47609 -55139 47669
rect -55079 47669 -50656 47672
rect -55079 47609 -55005 47669
rect -55211 47606 -55005 47609
rect -54945 47606 -50656 47669
rect -46556 47660 -44588 47760
rect -30735 47721 -30689 47818
rect -55305 47587 -50656 47606
rect -44688 47591 -44588 47660
rect -10867 47647 -10383 47674
rect -44937 47567 -40295 47591
rect -44937 47564 -44776 47567
rect -44937 47501 -44908 47564
rect -44848 47504 -44776 47564
rect -44716 47564 -40295 47567
rect -44716 47504 -44642 47564
rect -44848 47501 -44642 47504
rect -44582 47501 -40295 47564
rect -36195 47547 -34305 47647
rect -10919 47601 -10383 47647
rect -23402 47561 -15472 47591
rect -10867 47574 -10383 47601
rect -23402 47558 -23251 47561
rect -44937 47474 -40295 47501
rect -53825 47213 -53188 47281
rect -53953 46870 -53843 46884
rect -53953 46793 -53933 46870
rect -53856 46793 -53843 46870
rect -53953 46754 -53843 46793
rect -53953 46731 -53180 46754
rect -53953 46650 -53936 46731
rect -53855 46677 -53180 46731
rect -53051 46714 -46132 46786
rect -53855 46650 -53843 46677
rect -53953 46634 -53843 46650
rect -44693 46150 -44553 47474
rect -43479 47197 -43171 47213
rect -43479 47168 -43454 47197
rect -43495 47100 -43454 47168
rect -43479 47097 -43454 47100
rect -43354 47196 -43171 47197
rect -43354 47098 -43282 47196
rect -43184 47168 -43171 47196
rect -43184 47100 -42827 47168
rect -43184 47098 -43171 47100
rect -43354 47097 -43171 47098
rect -43479 47079 -43171 47097
rect -43767 46629 -43510 46641
rect -43401 46629 -42819 46641
rect -43767 46555 -43752 46629
rect -43678 46555 -43597 46629
rect -43523 46564 -42819 46629
rect -42690 46601 -35771 46673
rect -43523 46555 -43283 46564
rect -43767 46539 -43510 46555
rect -34622 46370 -34424 47547
rect -23402 47495 -23383 47558
rect -23323 47498 -23251 47558
rect -23191 47558 -15472 47561
rect -23191 47498 -23117 47558
rect -23323 47495 -23117 47498
rect -23057 47495 -15472 47558
rect -23402 47474 -15472 47495
rect -18993 47188 -18665 47226
rect -18993 47187 -18775 47188
rect -18993 47089 -18960 47187
rect -18862 47089 -18775 47187
rect -18993 47088 -18775 47089
rect -18675 47088 -18001 47188
rect -18993 47053 -18665 47088
rect -10483 47046 -10383 47574
rect -10233 47399 -10084 48021
rect 16771 48012 16849 48051
rect -7142 47985 -6762 48003
rect -7142 47982 -6990 47985
rect -7142 47979 -7122 47982
rect -7147 47919 -7122 47979
rect -7062 47922 -6990 47982
rect -6930 47982 -6762 47985
rect -6930 47922 -6856 47982
rect -7062 47919 -6856 47922
rect -6796 47979 -6762 47982
rect -6796 47919 -3755 47979
rect -7147 47901 -3755 47919
rect 16771 47952 16787 48012
rect 16840 47952 16849 48012
rect 16771 47923 16849 47952
rect 16771 47869 17965 47923
rect 16771 47809 16781 47869
rect 16834 47845 17965 47869
rect 16834 47809 16849 47845
rect 16771 47795 16849 47809
rect -9075 47700 -7507 47726
rect -9075 47697 -7741 47700
rect -9075 47634 -7873 47697
rect -7813 47637 -7741 47697
rect -7681 47697 -7507 47700
rect -7681 47637 -7607 47697
rect -7813 47634 -7607 47637
rect -7547 47634 -7507 47697
rect 2732 47688 5232 47703
rect 2732 47685 4979 47688
rect -9075 47613 -7507 47634
rect -7150 47612 -1368 47647
rect -7150 47609 -6991 47612
rect -7150 47546 -7123 47609
rect -7063 47549 -6991 47609
rect -6931 47609 -1368 47612
rect -6931 47549 -6857 47609
rect -7063 47546 -6857 47549
rect -6797 47546 -1368 47609
rect 2732 47616 4844 47685
rect 4902 47619 4979 47685
rect 5037 47686 5232 47688
rect 5037 47619 5128 47686
rect 4902 47617 5128 47619
rect 5186 47617 5232 47686
rect 8111 47683 8157 47788
rect 4902 47616 5232 47617
rect 2732 47603 5232 47616
rect 24452 47642 26426 47647
rect 24452 47638 26306 47642
rect -7150 47530 -1368 47546
rect 15312 47557 20352 47591
rect 15312 47554 15474 47557
rect 15312 47491 15342 47554
rect 15402 47494 15474 47554
rect 15534 47554 20352 47557
rect 15534 47494 15608 47554
rect 15402 47491 15608 47494
rect 15668 47491 20352 47554
rect 24452 47556 26026 47638
rect 26085 47556 26164 47638
rect 26223 47560 26306 47638
rect 26365 47560 26426 47642
rect 26223 47556 26426 47560
rect 24452 47547 26426 47556
rect 15312 47474 20352 47491
rect -8615 47442 -8384 47459
rect -10233 47365 -9969 47399
rect -8615 47388 -8599 47442
rect -8546 47440 -8384 47442
rect -8546 47388 -8468 47440
rect -9172 47386 -8468 47388
rect -8415 47388 -8384 47440
rect -8415 47386 -8383 47388
rect -10233 47284 -9873 47365
rect -9172 47300 -8383 47386
rect -9172 47298 -8464 47300
rect -10233 47250 -9969 47284
rect -9172 47245 -8594 47298
rect -8615 47244 -8594 47245
rect -8541 47246 -8464 47298
rect -8411 47246 -8383 47300
rect -8541 47245 -8383 47246
rect -8541 47244 -8384 47245
rect -8615 47228 -8384 47244
rect -4499 47156 -3900 47224
rect -10483 46946 -9777 47046
rect -9058 47001 -6741 47026
rect -9058 46998 -6986 47001
rect -9058 46935 -7118 46998
rect -7058 46938 -6986 46998
rect -6926 46998 -6741 47001
rect -6926 46938 -6852 46998
rect -7058 46935 -6852 46938
rect -6792 46935 -6741 46998
rect -9058 46913 -6741 46935
rect -31914 46704 -31714 46716
rect -4661 46713 -4350 46727
rect -32095 46703 -31785 46704
rect -32095 46648 -31908 46703
rect -31853 46648 -31785 46703
rect -32095 46647 -31785 46648
rect -31728 46647 -31439 46704
rect -31914 46636 -31714 46647
rect -18454 46645 -18175 46668
rect -18454 46641 -18434 46645
rect -18578 46564 -18434 46641
rect -18454 46556 -18434 46564
rect -18345 46644 -18175 46645
rect -18345 46557 -18276 46644
rect -18189 46641 -18175 46644
rect -18189 46564 -17996 46641
rect -17867 46601 -10948 46673
rect -4661 46618 -4647 46713
rect -4552 46712 -4350 46713
rect -4552 46619 -4457 46712
rect -4364 46697 -4350 46712
rect -4364 46620 -3892 46697
rect -3763 46657 3156 46729
rect 6967 46664 7166 46678
rect 6751 46663 7407 46664
rect -4364 46619 -4350 46620
rect -4552 46618 -4350 46619
rect -4661 46607 -4350 46618
rect 6751 46608 6977 46663
rect 7032 46608 7098 46663
rect 7153 46608 7407 46663
rect 6751 46607 7407 46608
rect 6967 46597 7166 46607
rect -18189 46557 -18175 46564
rect -18345 46556 -18175 46557
rect -18454 46540 -18175 46556
rect -34707 46337 -31310 46370
rect -34707 46334 -34550 46337
rect -34707 46271 -34682 46334
rect -34622 46274 -34550 46334
rect -34490 46334 -31310 46337
rect -34490 46274 -34416 46334
rect -34622 46271 -34416 46274
rect -34356 46271 -31310 46334
rect -34707 46257 -31310 46271
rect -24768 46342 -22997 46364
rect -24768 46265 -23383 46342
rect -23320 46341 -22997 46342
rect -23320 46265 -23240 46341
rect -24768 46264 -23240 46265
rect -23177 46264 -23101 46341
rect -23038 46264 -22997 46341
rect -46476 46010 -44540 46150
rect -34585 46030 -34462 46257
rect -24768 46253 -22997 46264
rect 4817 46294 7536 46330
rect 15447 46329 15578 47474
rect 17221 47100 17820 47168
rect 16994 46829 17122 46852
rect 16994 46737 17013 46829
rect 17105 46737 17122 46829
rect 16994 46668 17122 46737
rect 16994 46574 17012 46668
rect 17106 46641 17122 46668
rect 17106 46574 17828 46641
rect 17957 46601 24876 46673
rect 16994 46564 17828 46574
rect 16994 46560 17122 46564
rect 4817 46291 4981 46294
rect 4817 46228 4849 46291
rect 4909 46231 4981 46291
rect 5041 46291 7536 46294
rect 5041 46231 5115 46291
rect 4909 46228 5115 46231
rect 5175 46228 7536 46291
rect 4817 46217 7536 46228
rect 4933 46104 5236 46217
rect 14068 46198 15724 46329
rect -36106 45907 -34462 46030
rect -32085 45973 -31005 46067
rect -11511 46006 -6738 46036
rect -11511 46003 -6836 46006
rect -11511 45906 -7129 46003
rect -7059 45999 -6836 46003
rect -7059 45906 -6984 45999
rect -11511 45902 -6984 45906
rect -6914 45909 -6836 45999
rect -6766 45909 -6738 46006
rect 2801 45944 5236 46104
rect 6761 45933 7841 46027
rect 24433 46002 26418 46031
rect 24433 46000 26174 46002
rect -6914 45902 -6738 45909
rect -11511 45877 -6738 45902
rect 24433 45918 26034 46000
rect 26093 45920 26174 46000
rect 26233 46001 26418 46002
rect 26233 45920 26325 46001
rect 26093 45919 26325 45920
rect 26384 45919 26418 46001
rect 26093 45918 26418 45919
rect 24433 45900 26418 45918
rect -4975 45266 -4851 45404
rect -4975 45190 -4954 45266
rect -4870 45190 -4851 45266
rect -4975 45155 -4851 45190
rect 16254 45155 16393 45174
rect -4996 45105 16393 45155
rect -4996 45091 16282 45105
rect -4996 45015 -4949 45091
rect -4865 45017 16282 45091
rect 16382 45017 16393 45105
rect -4865 45015 16393 45017
rect -4996 44988 16393 45015
rect -4975 44983 -4851 44988
rect 16254 44907 16393 44988
rect -43973 44795 -43853 44849
rect 16254 44819 16272 44907
rect 16372 44819 16393 44907
rect 16254 44798 16393 44819
rect -43973 44733 -43938 44795
rect -43884 44733 -43853 44795
rect -43973 44665 -43853 44733
rect -33980 44672 -33860 44717
rect -33980 44665 -33957 44672
rect -43973 44653 -33957 44665
rect -43973 44591 -43941 44653
rect -43887 44612 -33957 44653
rect -33884 44612 -33860 44672
rect -43887 44591 -33860 44612
rect -43973 44545 -33860 44591
rect -33980 44527 -33860 44545
rect -33980 44467 -33959 44527
rect -33886 44467 -33860 44527
rect -19394 44610 -19274 44711
rect -19394 44543 -19373 44610
rect -19296 44543 -19274 44610
rect -19394 44483 -19274 44543
rect -5153 44578 -5020 44627
rect -5153 44515 -5125 44578
rect -5047 44515 -5020 44578
rect -5153 44483 -5020 44515
rect -33980 44441 -33860 44467
rect -31939 44415 -31828 44464
rect -31939 44345 -31905 44415
rect -31844 44345 -31828 44415
rect -19400 44449 -5020 44483
rect -19400 44382 -19373 44449
rect -19296 44412 -5020 44449
rect -19296 44382 -5129 44412
rect -19400 44350 -5129 44382
rect -43648 44256 -43256 44272
rect -31939 44256 -31828 44345
rect -5153 44349 -5129 44350
rect -5051 44349 -5020 44412
rect -5153 44329 -5020 44349
rect -43648 44145 -43630 44256
rect -43519 44255 -30823 44256
rect -43519 44146 -43378 44255
rect -43268 44236 -30823 44255
rect -43268 44166 -31915 44236
rect -31854 44166 -30823 44236
rect -43268 44146 -30823 44166
rect -43519 44145 -30823 44146
rect -43648 44134 -43256 44145
rect -30934 44015 -30823 44145
rect -30945 43996 -30823 44015
rect -43394 43936 -43015 43953
rect -31602 43936 -31461 43941
rect -43394 43825 -43380 43936
rect -43269 43935 -31461 43936
rect -43269 43826 -43132 43935
rect -43023 43906 -31461 43935
rect -43023 43826 -31577 43906
rect -43269 43825 -31577 43826
rect -43394 43813 -43015 43825
rect -31602 43797 -31577 43825
rect -31468 43797 -31461 43906
rect -31602 43693 -31461 43797
rect -30945 43913 -30930 43996
rect -30847 43966 -30823 43996
rect -18983 44132 -18856 44155
rect -18983 44043 -18962 44132
rect -18880 44126 -18856 44132
rect -4191 44126 -3830 44141
rect 7012 44126 7225 44147
rect -18880 44043 -4168 44126
rect -18983 44042 -4168 44043
rect -4084 44042 -3928 44126
rect -3844 44118 7225 44126
rect -3844 44117 7145 44118
rect -3844 44062 7031 44117
rect 7083 44063 7145 44117
rect 7197 44063 7225 44118
rect 7083 44062 7225 44063
rect -3844 44042 7225 44062
rect -30847 43913 -30827 43966
rect -30945 43817 -30827 43913
rect -30945 43736 -30928 43817
rect -30847 43736 -30827 43817
rect -18983 43890 -18856 44042
rect -4191 44015 -3830 44042
rect 7012 44035 7225 44042
rect -18983 43806 -18963 43890
rect -18879 43806 -18856 43890
rect -18983 43792 -18856 43806
rect 7807 43946 7945 43964
rect 7807 43868 7834 43946
rect 7910 43868 7945 43946
rect -30945 43721 -30827 43736
rect -18496 43757 -18336 43788
rect -4884 43757 -4404 43783
rect 7807 43762 7945 43868
rect 7807 43757 7842 43762
rect -18496 43756 -4553 43757
rect -31602 43692 -31459 43693
rect -31602 43581 -31579 43692
rect -31468 43581 -31459 43692
rect -31602 43580 -31459 43581
rect -18496 43647 -18472 43756
rect -18363 43750 -4857 43756
rect -18361 43647 -4857 43750
rect -4748 43647 -4553 43756
rect -18496 43641 -18470 43647
rect -18361 43646 -4553 43647
rect -4437 43684 7842 43757
rect 7918 43684 7945 43762
rect -4437 43646 7945 43684
rect -18361 43641 -18336 43646
rect -31602 43551 -31461 43580
rect -31993 43365 -30852 43439
rect -18496 43398 -18336 43641
rect -4884 43622 -4404 43646
rect 7807 43640 7945 43646
rect -18496 43287 -18472 43398
rect -18361 43287 -18336 43398
rect -18496 43267 -18336 43287
rect -3939 43497 -3831 43510
rect -3939 43423 -3921 43497
rect -3847 43423 -3831 43497
rect -3939 43364 -3831 43423
rect -3939 43363 -3611 43364
rect -3939 43291 -3920 43363
rect -3848 43291 -3611 43363
rect -3939 43290 -3611 43291
rect -3939 43271 -3831 43290
rect -35829 43097 -34300 43106
rect -35829 43093 -34392 43097
rect -35829 43092 -34537 43093
rect -55306 43046 -40305 43058
rect -55306 43045 -54984 43046
rect -55306 43044 -55133 43045
rect -55306 42963 -55281 43044
rect -55217 42964 -55133 43044
rect -55069 42965 -54984 43045
rect -54920 43041 -40305 43046
rect -54920 43040 -44635 43041
rect -54920 43039 -44782 43040
rect -54920 42965 -44931 43039
rect -44870 42966 -44782 43039
rect -44721 42967 -44635 43040
rect -44574 42967 -40305 43041
rect -35829 43015 -34690 43092
rect -34620 43016 -34537 43092
rect -34467 43020 -34392 43093
rect -34322 43020 -34300 43097
rect -34467 43016 -34300 43020
rect -34620 43015 -34300 43016
rect -35829 43001 -34300 43015
rect -24699 43078 -22958 43105
rect -24699 43076 -23244 43078
rect -24699 42994 -23387 43076
rect -23321 42996 -23244 43076
rect -23178 43076 -22958 43078
rect -23178 42996 -23090 43076
rect -23321 42994 -23090 42996
rect -23024 43002 -22958 43076
rect 3488 43020 9983 43032
rect 3488 43010 4980 43020
rect -23024 42994 -15027 43002
rect -24699 42980 -15027 42994
rect -44721 42966 -40305 42967
rect -44870 42965 -40305 42966
rect -55069 42964 -40305 42965
rect -55217 42963 -40305 42964
rect -55306 42953 -40305 42963
rect -40410 42851 -40305 42953
rect -31592 42863 -31451 42901
rect -23083 42877 -15027 42980
rect -10670 42953 -6742 42967
rect -10670 42951 -6989 42953
rect -10670 42935 -7135 42951
rect -10749 42889 -7135 42935
rect -31592 42752 -31579 42863
rect -31470 42752 -31451 42863
rect -10670 42871 -7135 42889
rect -7074 42873 -6989 42951
rect -6928 42873 -6840 42953
rect -6779 42873 -6742 42953
rect 3488 42920 4840 43010
rect 4920 42930 4980 43010
rect 5060 43010 9983 43020
rect 5060 42930 5120 43010
rect 4920 42920 5120 42930
rect 5200 42920 9983 43010
rect 3488 42908 9983 42920
rect 14199 42945 20614 42965
rect 14199 42943 15464 42945
rect -7074 42871 -6742 42873
rect -10670 42858 -6742 42871
rect 14199 42872 15330 42943
rect 15389 42874 15464 42943
rect 15523 42874 15601 42945
rect 15660 42874 20614 42945
rect 26027 42881 31528 42986
rect 15389 42872 20614 42874
rect 14199 42860 20614 42872
rect 20424 42807 20614 42860
rect 24852 42872 31528 42881
rect 24852 42866 26419 42872
rect 24852 42861 26169 42866
rect 24852 42786 26028 42861
rect 26087 42791 26169 42861
rect 26228 42865 26419 42866
rect 26228 42791 26323 42865
rect 26087 42790 26323 42791
rect 26382 42790 26419 42865
rect 26087 42786 26419 42790
rect 24852 42776 26419 42786
rect -31592 42738 -31451 42752
rect -59197 42645 -57435 42697
rect -31990 42627 -31451 42738
rect -31592 42625 -31451 42627
rect -65696 42502 -62555 42523
rect -31592 42514 -31580 42625
rect -31469 42514 -31451 42625
rect -4589 42663 -4184 42697
rect -4589 42552 -4553 42663
rect -4442 42662 -3515 42663
rect -4442 42553 -4311 42662
rect -4202 42553 -3515 42662
rect -4442 42552 -3515 42553
rect -4589 42524 -4184 42552
rect -31592 42511 -31451 42514
rect -65696 42501 -65415 42502
rect -65696 42498 -65547 42501
rect -65696 42425 -65689 42498
rect -65623 42428 -65547 42498
rect -65481 42429 -65415 42501
rect -65349 42429 -62555 42502
rect -65481 42428 -62555 42429
rect -65623 42425 -62555 42428
rect -65696 42410 -62555 42425
rect -65696 42388 -65296 42410
rect -68388 42258 -65296 42388
rect -66443 42137 -62617 42166
rect -69864 42104 -62617 42137
rect -69864 42017 -62491 42104
rect -66443 41988 -62491 42017
rect -55936 42094 -52516 42147
rect -55936 42090 -55633 42094
rect -55936 42086 -55769 42090
rect -55936 42015 -55907 42086
rect -55849 42019 -55769 42086
rect -55711 42023 -55633 42090
rect -55575 42023 -52516 42094
rect -45775 42139 -42210 42195
rect -45775 42131 -45591 42139
rect -45775 42075 -45731 42131
rect -45679 42083 -45591 42131
rect -45539 42130 -42210 42139
rect -45539 42083 -45462 42130
rect -45679 42075 -45462 42083
rect -45775 42074 -45462 42075
rect -45410 42074 -42210 42130
rect -45775 42045 -42210 42074
rect -55711 42019 -52516 42023
rect -55849 42015 -52516 42019
rect -55936 41997 -52516 42015
rect -24204 42016 -17163 42054
rect -24204 42003 -24043 42016
rect -24204 41947 -24173 42003
rect -24121 41960 -24043 42003
rect -23991 42003 -17163 42016
rect -23991 41960 -23920 42003
rect -24121 41947 -23920 41960
rect -23868 41947 -17163 42003
rect -24204 41904 -17163 41947
rect 4060 41998 6623 42054
rect 4060 41995 4208 41998
rect 4060 41939 4087 41995
rect 4139 41942 4208 41995
rect 4260 41942 4322 41998
rect 4374 41942 6623 41998
rect 25319 42019 28312 42071
rect 25319 42016 25485 42019
rect 4139 41939 6623 41942
rect 4060 41904 6623 41939
rect 14619 41904 17370 41970
rect 25319 41953 25353 42016
rect 25413 41956 25485 42016
rect 25545 42016 28312 42019
rect 25545 41956 25619 42016
rect 25413 41953 25619 41956
rect 25679 41953 28312 42016
rect 25319 41921 28312 41953
rect 14619 41900 14923 41904
rect 14619 41899 14802 41900
rect -68498 41790 -65981 41834
rect -68498 41703 -66364 41790
rect -66303 41703 -66233 41790
rect -66172 41784 -65981 41790
rect -66172 41703 -66077 41784
rect -68498 41697 -66077 41703
rect -66016 41697 -65981 41784
rect -68498 41682 -65981 41697
rect -63314 41805 -62482 41893
rect 14619 41843 14659 41899
rect 14711 41844 14802 41899
rect 14854 41848 14923 41900
rect 14975 41848 17370 41904
rect 14854 41844 17370 41848
rect 14711 41843 17370 41844
rect 14619 41820 17370 41843
rect -63314 41726 -62488 41805
rect -42874 41787 -42751 41801
rect -53195 41757 -53072 41771
rect -63314 41637 -63147 41726
rect -53195 41678 -53175 41757
rect -53084 41678 -53072 41757
rect -42874 41708 -42854 41787
rect -42763 41708 -42751 41787
rect -40602 41725 -40470 41771
rect -42874 41693 -42751 41708
rect -53195 41645 -53072 41678
rect -65600 41470 -63147 41637
rect -53866 41605 -53035 41645
rect -43560 41635 -42729 41693
rect 28791 41689 28914 41703
rect -43560 41611 -42858 41635
rect -53866 41563 -53179 41605
rect -53195 41526 -53179 41563
rect -53088 41563 -53035 41605
rect -53088 41526 -53072 41563
rect -42874 41556 -42858 41611
rect -42767 41611 -42729 41635
rect -17825 41655 -17702 41669
rect -42767 41556 -42751 41611
rect -42874 41544 -42751 41556
rect -17825 41576 -17805 41655
rect -17714 41576 -17702 41655
rect 9441 41584 9548 41630
rect 28791 41610 28811 41689
rect 28902 41610 28914 41689
rect -17825 41552 -17702 41576
rect -53195 41514 -53072 41526
rect -18513 41503 -17682 41552
rect -18513 41470 -17809 41503
rect -65600 41161 -65433 41470
rect -17825 41424 -17809 41470
rect -17718 41470 -17682 41503
rect 7109 41542 7296 41554
rect 7109 41541 7232 41542
rect 7109 41487 7119 41541
rect 7173 41487 7232 41541
rect 7109 41486 7232 41487
rect 7288 41537 7296 41542
rect 7288 41494 7318 41537
rect 16528 41532 16632 41566
rect 7288 41486 7384 41494
rect 7109 41471 7384 41486
rect -17718 41424 -17702 41470
rect 7272 41448 7384 41471
rect 16528 41459 16546 41532
rect 16617 41468 16632 41532
rect 17838 41565 17961 41579
rect 17838 41486 17858 41565
rect 17949 41486 17961 41565
rect 16617 41459 17242 41468
rect -17825 41412 -17702 41424
rect 16528 41386 17242 41459
rect 17838 41413 17961 41486
rect 28791 41537 28914 41610
rect 31055 41601 31183 41647
rect 28791 41458 28807 41537
rect 28898 41458 28914 41537
rect 28791 41446 28914 41458
rect 16528 41362 16632 41386
rect 16528 41289 16541 41362
rect 16612 41289 16632 41362
rect 17838 41334 17854 41413
rect 17945 41334 17961 41413
rect 17838 41322 17961 41334
rect 16528 41267 16632 41289
rect -66601 41133 -65433 41161
rect -69420 41120 -69330 41121
rect -69420 41107 -69215 41120
rect -69420 41042 -69407 41107
rect -69346 41042 -69215 41107
rect -69420 41029 -69215 41042
rect -69419 41027 -69215 41029
rect -66835 41021 -65433 41133
rect -66601 40994 -65433 41021
rect -63615 40954 -62748 40988
rect -63615 40847 -63590 40954
rect -63479 40847 -62748 40954
rect -63615 40829 -62748 40847
rect -63615 40821 -63448 40829
rect -44020 40786 -43854 40804
rect -54190 40754 -54017 40769
rect -54190 40702 -54168 40754
rect -54040 40702 -54017 40754
rect -54190 40676 -54017 40702
rect -44020 40732 -44003 40786
rect -43874 40732 -43854 40786
rect -44020 40724 -43854 40732
rect -54190 40630 -53031 40676
rect -44020 40667 -42725 40724
rect -19720 40738 -19576 40765
rect -54190 40578 -54168 40630
rect -54040 40602 -53031 40630
rect -44020 40613 -44003 40667
rect -43874 40650 -42725 40667
rect -19720 40664 -19690 40738
rect -19616 40664 -19576 40738
rect -43874 40613 -43854 40650
rect -54040 40578 -54017 40602
rect -68436 40534 -65296 40565
rect -68436 40529 -65549 40534
rect -68436 40444 -65678 40529
rect -65617 40449 -65549 40529
rect -65488 40531 -65296 40534
rect -65488 40449 -65389 40531
rect -65617 40446 -65389 40449
rect -65328 40446 -65296 40531
rect -65617 40444 -65296 40446
rect -68436 40425 -65296 40444
rect -54190 40487 -54017 40578
rect -54190 40435 -54167 40487
rect -54039 40435 -54017 40487
rect -54190 40416 -54017 40435
rect -44020 40553 -43854 40613
rect -19720 40608 -19576 40664
rect -44020 40499 -44004 40553
rect -43875 40499 -43854 40553
rect -44020 40399 -43854 40499
rect -35408 40573 -31837 40580
rect -35408 40570 -35099 40573
rect -35408 40568 -35248 40570
rect -35408 40512 -35369 40568
rect -35317 40514 -35248 40568
rect -35196 40517 -35099 40570
rect -35047 40517 -31837 40573
rect -35196 40514 -31837 40517
rect -35317 40512 -31837 40514
rect -35408 40498 -31837 40512
rect -19720 40534 -19689 40608
rect -19615 40583 -19576 40608
rect -19615 40534 -17678 40583
rect 4836 40595 5185 40618
rect 4836 40588 4972 40595
rect 4836 40583 4855 40588
rect -19720 40509 -17678 40534
rect 4830 40532 4855 40583
rect 4907 40539 4972 40588
rect 5024 40592 5185 40595
rect 5024 40539 5089 40592
rect 4907 40536 5089 40539
rect 5141 40583 5185 40592
rect 27286 40613 27390 40627
rect 5141 40536 6591 40583
rect 27286 40558 27306 40613
rect 27364 40600 27390 40613
rect 27364 40558 28326 40600
rect 4907 40532 6591 40536
rect 4830 40509 6591 40532
rect 16277 40529 16379 40545
rect -19720 40472 -19576 40509
rect -19720 40398 -19689 40472
rect -19615 40398 -19576 40472
rect -7944 40490 -3746 40505
rect -7944 40434 -7900 40490
rect -7848 40434 -7768 40490
rect -7716 40489 -3746 40490
rect -7716 40434 -7647 40489
rect -7944 40433 -7647 40434
rect -7595 40433 -3746 40489
rect -7944 40423 -3746 40433
rect 16277 40463 16299 40529
rect 16363 40499 16379 40529
rect 27286 40526 28326 40558
rect 16363 40463 17265 40499
rect 16277 40425 17265 40463
rect 27286 40469 27390 40526
rect -19720 40378 -19576 40398
rect 16277 40391 16379 40425
rect 16277 40325 16301 40391
rect 16365 40325 16379 40391
rect 16277 40239 16379 40325
rect 27286 40414 27311 40469
rect 27369 40414 27390 40469
rect 27286 40343 27390 40414
rect 27286 40288 27309 40343
rect 27367 40288 27390 40343
rect 27286 40262 27390 40288
rect 16277 40173 16289 40239
rect 16353 40173 16379 40239
rect 16277 40150 16379 40173
rect -68614 40006 -65978 40054
rect -68614 39919 -66359 40006
rect -66299 40002 -65978 40006
rect -66299 39919 -66224 40002
rect -68614 39915 -66224 39919
rect -66164 40001 -65978 40002
rect -66164 39915 -66089 40001
rect -68614 39914 -66089 39915
rect -66029 39914 -65978 40001
rect -68614 39893 -65978 39914
rect -65421 40019 -62932 40034
rect -65421 39877 -62857 40019
rect -65421 39863 -62932 39877
rect -65421 39396 -65250 39863
rect -44933 39752 -44585 39771
rect -44943 39750 -44669 39752
rect -55284 39724 -54906 39741
rect -55284 39723 -54996 39724
rect -55284 39721 -55137 39723
rect -55284 39704 -55273 39721
rect -55299 39650 -55273 39704
rect -55215 39652 -55137 39721
rect -55079 39653 -54996 39723
rect -54938 39704 -54906 39724
rect -54938 39653 -53035 39704
rect -44943 39694 -44918 39750
rect -44866 39694 -44788 39750
rect -44736 39696 -44669 39750
rect -44617 39696 -42729 39752
rect 28461 39732 28584 39746
rect -44736 39694 -42729 39696
rect -44943 39674 -42729 39694
rect 6210 39694 6288 39728
rect -55079 39652 -53035 39653
rect -55215 39650 -53035 39652
rect -55299 39626 -53035 39650
rect -30651 39531 -30605 39615
rect -23393 39613 -23028 39635
rect -23393 39611 -23244 39613
rect -23402 39607 -23244 39611
rect -23402 39551 -23377 39607
rect -23325 39557 -23244 39607
rect -23192 39557 -23108 39613
rect -23056 39611 -23028 39613
rect 6210 39631 6222 39694
rect 6275 39631 6288 39694
rect 6210 39611 6288 39631
rect 16745 39643 16868 39657
rect -23056 39557 -17682 39611
rect -23325 39551 -17682 39557
rect -23402 39533 -17682 39551
rect 6210 39556 6649 39611
rect -36242 39467 -34303 39476
rect -36242 39464 -34393 39467
rect -66601 39361 -65250 39396
rect -46548 39420 -44762 39428
rect -46548 39379 -40342 39420
rect -46548 39377 -44659 39379
rect -67917 39335 -67684 39360
rect -69533 39299 -69355 39309
rect -69533 39225 -69513 39299
rect -69434 39225 -69355 39299
rect -67917 39268 -67893 39335
rect -67820 39268 -67684 39335
rect -67917 39242 -67684 39268
rect -66813 39259 -65250 39361
rect -66601 39225 -65250 39259
rect -55292 39346 -50648 39372
rect -55292 39345 -55003 39346
rect -55292 39343 -55144 39345
rect -55292 39272 -55280 39343
rect -55222 39274 -55144 39343
rect -55086 39275 -55003 39345
rect -54945 39275 -50648 39346
rect -46548 39328 -44908 39377
rect -44970 39321 -44908 39328
rect -44856 39321 -44778 39377
rect -44726 39323 -44659 39377
rect -44607 39323 -40342 39379
rect -36242 39387 -34694 39464
rect -34624 39387 -34544 39464
rect -34474 39390 -34393 39464
rect -34323 39390 -34303 39467
rect -34474 39387 -34303 39390
rect -36242 39376 -34303 39387
rect -44726 39321 -40342 39323
rect -44970 39303 -40342 39321
rect -23224 39279 -23077 39533
rect -2464 39438 -2418 39534
rect 6210 39493 6223 39556
rect 6276 39533 6649 39556
rect 16745 39564 16765 39643
rect 16856 39564 16868 39643
rect 6276 39493 6288 39533
rect 6210 39482 6288 39493
rect 16745 39527 16868 39564
rect 28461 39653 28481 39732
rect 28572 39653 28584 39732
rect 28461 39580 28584 39653
rect 16745 39491 17284 39527
rect 16745 39412 16761 39491
rect 16852 39449 17284 39491
rect 28461 39501 28477 39580
rect 28568 39501 28584 39580
rect 28461 39489 28584 39501
rect 16852 39412 16868 39449
rect 16745 39400 16868 39412
rect -55086 39274 -50648 39275
rect -55222 39272 -50648 39274
rect -55292 39255 -50648 39272
rect -23411 39245 -15295 39279
rect -23411 39239 -23243 39245
rect -69533 39210 -69355 39225
rect -23411 39183 -23376 39239
rect -23324 39189 -23243 39239
rect -23191 39189 -23107 39245
rect -23055 39189 -15295 39245
rect -11195 39235 -6884 39335
rect -23324 39183 -15295 39189
rect -23411 39162 -15295 39183
rect -63020 39051 -61629 39058
rect -63128 39031 -61629 39051
rect -63128 39017 -61581 39031
rect -63128 38910 -63103 39017
rect -62992 38920 -61581 39017
rect -62992 38910 -61629 38920
rect -63128 38893 -61629 38910
rect -63128 38884 -62961 38893
rect -53779 38881 -53180 38949
rect -43473 38929 -42874 38997
rect -68488 38754 -65297 38785
rect -68488 38746 -65373 38754
rect -68488 38659 -65682 38746
rect -65622 38745 -65373 38746
rect -65622 38659 -65525 38745
rect -68488 38658 -65525 38659
rect -65465 38667 -65373 38745
rect -65313 38667 -65297 38754
rect -65465 38658 -65297 38667
rect -68488 38648 -65297 38658
rect -67412 38450 -65981 38492
rect -43755 38470 -43481 38491
rect -43755 38459 -42866 38470
rect -43755 38454 -43595 38459
rect -67412 38448 -66064 38450
rect -67412 38447 -66225 38448
rect -67412 38343 -66367 38447
rect -66304 38344 -66225 38447
rect -66162 38346 -66064 38448
rect -66001 38346 -65981 38450
rect -66162 38344 -65981 38346
rect -66304 38343 -65981 38344
rect -67412 38326 -65981 38343
rect -53812 38413 -53172 38422
rect -53812 38344 -53804 38413
rect -53741 38345 -53172 38413
rect -53043 38382 -46124 38454
rect -43755 38400 -43728 38454
rect -43673 38405 -43595 38454
rect -43540 38405 -42866 38459
rect -42737 38430 -35818 38502
rect -33720 38499 -33512 38507
rect -33720 38498 -31355 38499
rect -33720 38443 -33700 38498
rect -33645 38443 -33574 38498
rect -33519 38443 -31355 38498
rect -33720 38442 -31355 38443
rect -33720 38429 -33512 38442
rect -43673 38400 -42866 38405
rect -43755 38393 -42866 38400
rect -43755 38368 -43481 38393
rect -53741 38344 -53735 38345
rect -53812 38253 -53735 38344
rect -53812 38184 -53805 38253
rect -53742 38184 -53735 38253
rect -53812 38163 -53735 38184
rect -34720 38133 -31226 38165
rect -23224 38163 -23077 39162
rect -18489 38886 -18167 38908
rect -18489 38775 -18470 38886
rect -18359 38885 -18167 38886
rect -18359 38776 -18296 38885
rect -18187 38856 -18167 38885
rect -18187 38788 -17827 38856
rect -18187 38776 -18167 38788
rect -18359 38775 -18167 38776
rect -18489 38756 -18167 38775
rect -9364 38740 -9133 38766
rect -9364 38670 -9350 38740
rect -9270 38670 -9133 38740
rect -9364 38620 -9133 38670
rect -9364 38550 -9250 38620
rect -9170 38550 -9133 38620
rect -9364 38535 -9133 38550
rect -19001 38331 -18631 38367
rect -19001 38247 -18963 38331
rect -18879 38247 -18731 38331
rect -18647 38329 -18356 38331
rect -18647 38252 -17819 38329
rect -17690 38289 -10771 38361
rect -18647 38247 -18356 38252
rect -19001 38224 -18631 38247
rect -34720 38131 -34405 38133
rect -34720 38125 -34538 38131
rect -65585 38072 -63352 38107
rect -65585 37968 -63175 38072
rect -34720 38069 -34669 38125
rect -34617 38075 -34538 38125
rect -34486 38077 -34405 38131
rect -34353 38077 -31226 38133
rect -34486 38075 -31226 38077
rect -34617 38069 -31226 38075
rect -34720 38052 -31226 38069
rect -65585 37933 -63352 37968
rect -65585 37813 -65411 37933
rect -34525 37869 -34404 38052
rect -24722 38016 -22992 38163
rect -6984 38090 -6884 39235
rect 4817 39244 6734 39279
rect 4817 39237 4973 39244
rect 4817 39181 4856 39237
rect 4908 39188 4973 39237
rect 5025 39241 6734 39244
rect 5025 39188 5090 39241
rect 4908 39185 5090 39188
rect 5142 39185 6734 39241
rect 13807 39235 15575 39335
rect 26010 39265 28399 39296
rect 26010 39262 26181 39265
rect 26010 39251 26049 39262
rect 4908 39181 6734 39185
rect 4817 39162 6734 39181
rect 15225 39195 15575 39235
rect 24258 39199 26049 39251
rect 26109 39202 26181 39262
rect 26241 39262 28399 39265
rect 26241 39202 26315 39262
rect 26109 39199 26315 39202
rect 26375 39199 28399 39262
rect 15225 39172 17365 39195
rect -5386 38430 -5204 38442
rect -5386 38428 -5266 38430
rect -5386 38372 -5374 38428
rect -5322 38374 -5266 38428
rect -5214 38424 -5204 38430
rect -5214 38374 -3675 38424
rect -5322 38372 -3675 38374
rect -5386 38367 -3675 38372
rect -5386 38359 -5204 38367
rect -7147 38053 -3705 38090
rect 4989 38081 5110 39162
rect 15225 39157 15353 39172
rect 15292 39116 15353 39157
rect 15405 39166 17365 39172
rect 15405 39162 15594 39166
rect 15405 39116 15470 39162
rect 15292 39106 15470 39116
rect 15522 39110 15594 39162
rect 15646 39110 17365 39166
rect 24258 39179 28399 39199
rect 24258 39151 26264 39179
rect 15522 39106 17365 39110
rect 15292 39078 17365 39106
rect 15448 39019 15575 39078
rect 6421 38967 6528 39015
rect 6421 38892 6437 38967
rect 6512 38892 6528 38967
rect 6421 38887 6528 38892
rect 6421 38796 7202 38887
rect 6421 38721 6435 38796
rect 6510 38780 7202 38796
rect 6510 38721 6528 38780
rect 6421 38711 6528 38721
rect 6666 38523 6775 38541
rect 6666 38431 6674 38523
rect 6766 38431 6775 38523
rect 6666 38346 6775 38431
rect 6664 38345 6776 38346
rect 6664 38251 6673 38345
rect 6767 38251 6776 38345
rect 8036 38289 8240 38361
rect 6664 38250 6776 38251
rect 6666 38235 6775 38250
rect -7147 38048 -6870 38053
rect -7147 38045 -6991 38048
rect -7147 37989 -7122 38045
rect -7070 37992 -6991 38045
rect -6939 37997 -6870 38048
rect -6818 37997 -3705 38053
rect -6939 37992 -3705 37997
rect -7070 37989 -3705 37992
rect -7147 37977 -3705 37989
rect -67256 37774 -65411 37813
rect -67547 37678 -65411 37774
rect -67256 37639 -65411 37678
rect -46466 37771 -44541 37811
rect -46466 37768 -44645 37771
rect -46466 37694 -44930 37768
rect -44869 37766 -44645 37768
rect -44869 37694 -44795 37766
rect -46466 37692 -44795 37694
rect -44734 37697 -44645 37766
rect -44584 37697 -44541 37771
rect -36152 37748 -34404 37869
rect -33313 37850 -30921 37862
rect -33313 37845 -33157 37850
rect -33313 37788 -33290 37845
rect -33230 37793 -33157 37845
rect -33097 37793 -30921 37850
rect -33230 37788 -30921 37793
rect -33313 37768 -30921 37788
rect -6960 37712 -6832 37977
rect 3498 37960 5110 38081
rect -44734 37692 -44541 37697
rect -46466 37675 -44541 37692
rect -11109 37584 -6832 37712
rect -5057 37753 -3705 37787
rect -5057 37701 -5049 37753
rect -4997 37701 -4936 37753
rect -4884 37701 -3705 37753
rect -5057 37693 -3705 37701
rect 15448 37678 15562 39019
rect 16996 38419 17117 38435
rect 16996 38327 17013 38419
rect 17105 38327 17117 38419
rect 16996 38260 17117 38327
rect 16996 38166 17012 38260
rect 17106 38245 17117 38260
rect 17106 38168 17411 38245
rect 18740 38205 20540 38277
rect 17106 38166 17117 38168
rect 16996 38144 17117 38166
rect 13899 37564 15562 37678
rect 26111 37618 26264 39151
rect 27929 38873 28138 38892
rect 27929 38805 27946 38873
rect 28014 38872 28338 38873
rect 28014 38806 28070 38872
rect 28136 38806 28338 38872
rect 28014 38805 28338 38806
rect 27929 38783 28138 38805
rect 28287 38346 28405 38348
rect 28287 38345 28550 38346
rect 28287 38270 28308 38345
rect 28383 38270 28550 38345
rect 29796 38306 31064 38378
rect 28287 38269 28550 38270
rect 28287 38197 28405 38269
rect 28287 38120 28307 38197
rect 28384 38120 28405 38197
rect 28287 38109 28405 38120
rect 24531 37465 26264 37618
rect -67465 37197 -65296 37225
rect -67465 37192 -65375 37197
rect -67465 37101 -65682 37192
rect -65614 37101 -65528 37192
rect -65460 37106 -65375 37192
rect -65307 37106 -65296 37197
rect -65460 37101 -65296 37106
rect -67465 37082 -65296 37101
rect -54508 36947 -54384 37025
rect -54508 36856 -54477 36947
rect -54406 36856 -54384 36947
rect -64663 36755 -64523 36758
rect -54508 36755 -54384 36856
rect -64663 36665 -54487 36755
rect -64663 36585 -64629 36665
rect -64549 36664 -54487 36665
rect -54416 36664 -54384 36755
rect -64549 36631 -54384 36664
rect -64549 36585 -64523 36631
rect -64663 36486 -64523 36585
rect -64663 36406 -64628 36486
rect -64548 36406 -64523 36486
rect -64663 36370 -64523 36406
rect -53821 36507 -53726 36519
rect -53821 36434 -53800 36507
rect -53729 36434 -53726 36507
rect -53821 36337 -53726 36434
rect -64384 36335 -53726 36337
rect -64388 36297 -53806 36335
rect -64388 36225 -64379 36297
rect -64303 36262 -53806 36297
rect -53735 36262 -53726 36335
rect -64303 36242 -53726 36262
rect -53258 36287 -53155 36296
rect -64303 36225 -64295 36242
rect -64388 36132 -64295 36225
rect -53258 36215 -53242 36287
rect -53165 36215 -53155 36287
rect -53258 36141 -53155 36215
rect -64125 36137 -53150 36141
rect -64388 36060 -64380 36132
rect -64304 36060 -64295 36132
rect -64388 36047 -64295 36060
rect -64142 36119 -53150 36137
rect -64142 36040 -64121 36119
rect -64046 36047 -53246 36119
rect -53169 36047 -53150 36119
rect -64046 36040 -53150 36047
rect -64142 36034 -53150 36040
rect -64142 35943 -64035 36034
rect -64142 35864 -64126 35943
rect -64051 35864 -64035 35943
rect -64142 35847 -64035 35864
rect 16258 35984 16384 36028
rect 16258 35921 16285 35984
rect 16365 35921 16384 35984
rect 16258 35818 16384 35921
rect 16258 35813 16281 35818
rect 6455 35767 16281 35813
rect 6455 35709 6484 35767
rect 6549 35755 16281 35767
rect 16361 35755 16384 35818
rect 6549 35726 16384 35755
rect 6549 35709 6563 35726
rect 6455 35640 6563 35709
rect 6455 35582 6480 35640
rect 6545 35582 6563 35640
rect 6455 35553 6563 35582
rect 27263 35598 27398 35633
rect 27263 35524 27309 35598
rect 27388 35524 27398 35598
rect -4643 35514 -4427 35517
rect -4688 35466 -4427 35514
rect -4688 35377 -4653 35466
rect -4575 35451 -4427 35466
rect 27263 35451 27398 35524
rect -4575 35415 27404 35451
rect -4575 35377 27308 35415
rect -4688 35341 27308 35377
rect 27387 35341 27404 35415
rect -4688 35316 27404 35341
rect -4688 35276 -4549 35316
rect -4688 35187 -4654 35276
rect -4576 35187 -4549 35276
rect -4688 35153 -4549 35187
rect 2036 34956 16677 35057
rect -25604 34941 16677 34956
rect -34022 34878 -33847 34879
rect -25604 34878 2152 34941
rect -34022 34871 2152 34878
rect -34022 34817 -33992 34871
rect -33863 34840 2152 34871
rect 16561 34867 16585 34941
rect 16649 34867 16677 34941
rect -33863 34817 -25488 34840
rect -34022 34762 -25488 34817
rect 16561 34797 16677 34867
rect -34022 34758 -33847 34762
rect -34022 34704 -33993 34758
rect -33864 34704 -33847 34758
rect -34022 34650 -33847 34704
rect 16561 34723 16589 34797
rect 16653 34723 16677 34797
rect 16561 34703 16677 34723
rect -65702 34613 -60638 34629
rect -65702 34610 -65386 34613
rect -65702 34510 -65680 34610
rect -65606 34510 -65534 34610
rect -65460 34513 -65386 34610
rect -65312 34513 -60638 34613
rect -65460 34510 -60638 34513
rect -65702 34499 -60638 34510
rect -56334 34598 -50381 34621
rect -56334 34595 -55156 34598
rect -56334 34520 -55284 34595
rect -55225 34523 -55156 34595
rect -55097 34597 -50381 34598
rect -55097 34523 -55027 34597
rect -55225 34522 -55027 34523
rect -54968 34522 -50381 34597
rect -55225 34520 -50381 34522
rect -56334 34507 -50381 34520
rect -46167 34593 -40008 34609
rect -46167 34520 -44928 34593
rect -44866 34592 -40008 34593
rect -44866 34520 -44802 34592
rect -46167 34519 -44802 34520
rect -44740 34519 -44647 34592
rect -44585 34519 -40008 34592
rect -34022 34596 -33992 34650
rect -33863 34596 -33847 34650
rect -46167 34506 -40008 34519
rect -35792 34573 -34299 34589
rect -35792 34572 -34545 34573
rect -35792 34483 -34693 34572
rect -34623 34484 -34545 34572
rect -34475 34572 -34299 34573
rect -34475 34484 -34401 34572
rect -34623 34483 -34401 34484
rect -34331 34483 -34299 34572
rect -35792 34472 -34299 34483
rect -34416 34278 -34299 34472
rect -34022 34539 -33847 34596
rect -34022 34485 -33999 34539
rect -33870 34485 -33847 34539
rect -34022 34466 -33847 34485
rect 3067 34494 9825 34516
rect 3067 34492 5137 34494
rect -10911 34435 -1335 34451
rect -24736 34379 -15284 34401
rect -29256 34365 -29139 34366
rect -29256 34278 -29113 34365
rect -24736 34301 -23382 34379
rect -23321 34378 -15284 34379
rect -23321 34301 -23242 34378
rect -24736 34300 -23242 34301
rect -23181 34377 -15284 34378
rect -23181 34300 -23081 34377
rect -24736 34299 -23081 34300
rect -23020 34299 -15284 34377
rect -10911 34360 -7133 34435
rect -7080 34434 -1335 34435
rect -7080 34431 -6869 34434
rect -7080 34360 -7003 34431
rect -10911 34356 -7003 34360
rect -6950 34359 -6869 34431
rect -6816 34359 -1335 34434
rect 3067 34423 4841 34492
rect 4906 34423 4991 34492
rect 5056 34425 5137 34492
rect 5202 34425 9825 34494
rect 5056 34423 9825 34425
rect 3067 34413 9825 34423
rect 14048 34440 20740 34454
rect 14048 34439 15622 34440
rect -6950 34356 -1335 34359
rect -10911 34349 -1335 34356
rect 14048 34362 15327 34439
rect 15402 34362 15478 34439
rect 15553 34363 15622 34439
rect 15697 34363 20740 34440
rect 15553 34362 20740 34363
rect 14048 34353 20740 34362
rect 24927 34406 31452 34420
rect -24736 34289 -15284 34299
rect -34416 34161 -29113 34278
rect -15453 34218 -15284 34289
rect -1498 34256 -1335 34349
rect 24927 34311 26028 34406
rect 26101 34311 26176 34406
rect 26249 34311 26330 34406
rect 26403 34311 31452 34406
rect 24927 34302 31452 34311
rect -1498 34255 -1396 34256
rect 31334 34188 31452 34302
rect -66381 33652 -63898 33706
rect -66381 33649 -66221 33652
rect -66381 33586 -66353 33649
rect -66293 33589 -66221 33649
rect -66161 33649 -63898 33652
rect -66161 33589 -66087 33649
rect -66293 33586 -66087 33589
rect -66027 33586 -63898 33649
rect -66381 33556 -63898 33586
rect -55937 33662 -53660 33699
rect -55937 33658 -55639 33662
rect -55937 33577 -55922 33658
rect -55854 33577 -55779 33658
rect -55711 33581 -55639 33658
rect -55571 33581 -53660 33662
rect -55711 33577 -53660 33581
rect -66277 32081 -66129 33556
rect -55937 33549 -53660 33577
rect -45763 33630 -43425 33672
rect -45763 33629 -45469 33630
rect -45763 33548 -45755 33629
rect -45685 33628 -45469 33629
rect -45685 33548 -45621 33628
rect -45763 33547 -45621 33548
rect -45551 33549 -45469 33628
rect -45399 33549 -43425 33630
rect -45551 33547 -43425 33549
rect -45763 33522 -43425 33547
rect -7912 33552 -4486 33606
rect -7912 33542 -7615 33552
rect -24190 33501 -18347 33542
rect -24190 33497 -23912 33501
rect -24190 33495 -24038 33497
rect -35391 33448 -32296 33487
rect -35391 33444 -35112 33448
rect -35391 33440 -35237 33444
rect -35391 33357 -35379 33440
rect -35309 33361 -35237 33440
rect -35167 33365 -35112 33444
rect -35042 33365 -32296 33448
rect -24190 33412 -24174 33495
rect -24104 33414 -24038 33495
rect -23968 33418 -23912 33497
rect -23842 33418 -18347 33501
rect -7912 33534 -7749 33542
rect -7912 33474 -7902 33534
rect -7848 33482 -7749 33534
rect -7695 33492 -7615 33542
rect -7561 33492 -4486 33552
rect -7695 33482 -4486 33492
rect -7848 33474 -4486 33482
rect -7912 33456 -4486 33474
rect 4069 33485 6502 33545
rect 25325 33512 28265 33574
rect 25325 33509 25488 33512
rect -23968 33414 -18347 33418
rect -24104 33412 -18347 33414
rect -24190 33392 -18347 33412
rect 4069 33421 4082 33485
rect 4138 33421 4220 33485
rect 4276 33484 6502 33485
rect 4276 33421 4360 33484
rect 4069 33420 4360 33421
rect 4416 33420 6502 33484
rect 4069 33395 6502 33420
rect 14619 33437 17466 33503
rect 14619 33433 14768 33437
rect -35167 33361 -32296 33365
rect -35309 33357 -32296 33361
rect -35391 33337 -32296 33357
rect 14619 33377 14655 33433
rect 14707 33381 14768 33433
rect 14820 33433 17466 33437
rect 14820 33381 14881 33433
rect 14707 33377 14881 33381
rect 14933 33377 17466 33433
rect 25325 33446 25356 33509
rect 25416 33449 25488 33509
rect 25548 33509 28265 33512
rect 25548 33449 25622 33509
rect 25416 33446 25622 33449
rect 25682 33446 28265 33509
rect 25325 33424 28265 33446
rect 14619 33353 17466 33377
rect -63376 33288 -63253 33302
rect -63376 33209 -63356 33288
rect -63265 33209 -63253 33288
rect -63376 33136 -63253 33209
rect -63376 33057 -63360 33136
rect -63269 33057 -63253 33136
rect -63376 33045 -63253 33057
rect -53204 33293 -53081 33307
rect -53204 33214 -53184 33293
rect -53093 33214 -53081 33293
rect -53204 33141 -53081 33214
rect -53204 33062 -53188 33141
rect -53097 33062 -53081 33141
rect -53204 33050 -53081 33062
rect -42810 33264 -42687 33278
rect -42810 33185 -42790 33264
rect -42699 33185 -42687 33264
rect -42810 33112 -42687 33185
rect -3974 33195 -3851 33209
rect -17936 33150 -17813 33164
rect -42810 33033 -42794 33112
rect -42703 33033 -42687 33112
rect -42810 33021 -42687 33033
rect -31751 33108 -31628 33122
rect -31751 33029 -31731 33108
rect -31640 33029 -31628 33108
rect -31751 32956 -31628 33029
rect -31751 32877 -31735 32956
rect -31644 32877 -31628 32956
rect -17936 33071 -17916 33150
rect -17825 33071 -17813 33150
rect -17936 32998 -17813 33071
rect -17936 32919 -17920 32998
rect -17829 32919 -17813 32998
rect -3974 33116 -3954 33195
rect -3863 33116 -3851 33195
rect -3974 33043 -3851 33116
rect -3974 32964 -3958 33043
rect -3867 32964 -3851 33043
rect -3974 32952 -3851 32964
rect 7002 33192 7125 33206
rect 7002 33113 7022 33192
rect 7113 33113 7125 33192
rect 7002 33040 7125 33113
rect 17889 33195 18012 33209
rect 17889 33116 17909 33195
rect 18000 33116 18012 33195
rect 7002 32961 7018 33040
rect 7109 32961 7125 33040
rect 7002 32949 7125 32961
rect 16847 33071 16953 33109
rect 16847 33000 16873 33071
rect 16940 33001 16953 33071
rect 17889 33043 18012 33116
rect 16940 33000 17350 33001
rect -17936 32907 -17813 32919
rect 16847 32919 17350 33000
rect 17889 32964 17905 33043
rect 17996 32964 18012 33043
rect 17889 32952 18012 32964
rect 28805 33195 28928 33209
rect 28805 33116 28825 33195
rect 28916 33116 28928 33195
rect 28805 33043 28928 33116
rect 28805 32964 28821 33043
rect 28912 32964 28928 33043
rect 28805 32952 28928 32964
rect -31751 32865 -31628 32877
rect 16847 32888 16953 32919
rect 16847 32817 16864 32888
rect 16931 32817 16953 32888
rect 16847 32800 16953 32817
rect -4682 32351 -4557 32472
rect -54190 32327 -54017 32350
rect -64663 32263 -64523 32326
rect -64663 32148 -64642 32263
rect -64555 32235 -64523 32263
rect -54190 32270 -54170 32327
rect -54034 32270 -54017 32327
rect -64555 32161 -63904 32235
rect -54190 32228 -54017 32270
rect -44020 32262 -43854 32274
rect -54190 32181 -53801 32228
rect -64555 32148 -64523 32161
rect -66824 31933 -65980 32081
rect -64663 32030 -64523 32148
rect -64663 31915 -64637 32030
rect -64550 31915 -64523 32030
rect -54190 32124 -54169 32181
rect -54033 32154 -53801 32181
rect -44020 32203 -44000 32262
rect -43873 32203 -43854 32262
rect -19708 32255 -19583 32317
rect -44020 32201 -43854 32203
rect -54033 32124 -54017 32154
rect -54190 32060 -54017 32124
rect -54190 32003 -54169 32060
rect -54033 32003 -54017 32060
rect -54190 31983 -54017 32003
rect -44020 32150 -43404 32201
rect -44020 32091 -44001 32150
rect -43874 32127 -43404 32150
rect -34022 32194 -33847 32214
rect -34022 32128 -34001 32194
rect -33863 32128 -33847 32194
rect -43874 32091 -43854 32127
rect -44020 32024 -43854 32091
rect -44020 31965 -44004 32024
rect -43877 31965 -43854 32024
rect -44020 31950 -43854 31965
rect -34022 32016 -33847 32128
rect -19708 32173 -19684 32255
rect -19601 32173 -19583 32255
rect -19708 32071 -19583 32173
rect -4682 32265 -4661 32351
rect -4574 32265 -4557 32351
rect -4682 32152 -4557 32265
rect -34022 32011 -32374 32016
rect -64663 31873 -64523 31915
rect -34022 31945 -34006 32011
rect -33868 31945 -32374 32011
rect -19708 31989 -19685 32071
rect -19602 31997 -18501 32071
rect -4682 32066 -4663 32152
rect -4576 32066 -4557 32152
rect -4682 32036 -4557 32066
rect 6455 32201 6563 32270
rect 6455 32129 6477 32201
rect 6543 32129 6563 32201
rect 6455 32044 6563 32129
rect -19602 31989 -19583 31997
rect -19708 31963 -19583 31989
rect 6455 31972 6478 32044
rect 6544 31972 6563 32044
rect 6455 31951 6563 31972
rect 16564 32171 16681 32237
rect 16564 32101 16584 32171
rect 16661 32101 16681 32171
rect 16564 32032 16681 32101
rect 27537 32161 27700 32190
rect 27537 32083 27573 32161
rect 27664 32103 27700 32161
rect 27664 32083 28215 32103
rect 16564 32007 17359 32032
rect -34022 31942 -32374 31945
rect -34022 31862 -33847 31942
rect 16564 31937 16583 32007
rect 16660 31958 17359 32007
rect 27537 32029 28215 32083
rect 16660 31937 16681 31958
rect 16564 31913 16681 31937
rect 27537 31954 27700 32029
rect -34022 31796 -34008 31862
rect -33870 31796 -33847 31862
rect 27537 31876 27582 31954
rect 27673 31876 27700 31954
rect 27537 31820 27700 31876
rect -34022 31780 -33847 31796
rect -63789 31350 -63666 31364
rect -63789 31294 -63769 31350
rect -63865 31271 -63769 31294
rect -63678 31271 -63666 31350
rect -68341 31187 -68170 31198
rect -68341 31130 -68318 31187
rect -68237 31130 -68170 31187
rect -68341 31113 -68170 31130
rect -66733 31186 -66583 31229
rect -66733 31115 -66690 31186
rect -66620 31115 -66583 31186
rect -63865 31198 -63666 31271
rect -63865 31154 -63773 31198
rect -66733 31079 -66583 31115
rect -63789 31119 -63773 31154
rect -63682 31119 -63666 31198
rect -63789 31107 -63666 31119
rect -53503 31350 -53380 31364
rect -53503 31271 -53483 31350
rect -53392 31271 -53380 31350
rect -53503 31198 -53380 31271
rect -53503 31119 -53487 31198
rect -53396 31119 -53380 31198
rect -53503 31107 -53380 31119
rect -43129 31319 -43006 31333
rect -43129 31240 -43109 31319
rect -43018 31240 -43006 31319
rect -43129 31167 -43006 31240
rect -4270 31225 -4147 31239
rect -43129 31088 -43113 31167
rect -43022 31088 -43006 31167
rect -18227 31174 -18104 31188
rect -43129 31076 -43006 31088
rect -32055 31134 -31932 31148
rect -32055 31055 -32035 31134
rect -31944 31055 -31932 31134
rect -65695 30906 -63845 30931
rect -65695 30903 -65547 30906
rect -65695 30840 -65679 30903
rect -65619 30843 -65547 30903
rect -65487 30903 -63845 30906
rect -65487 30843 -65413 30903
rect -65619 30840 -65413 30843
rect -65353 30840 -63845 30903
rect -56735 30924 -54913 30987
rect -32055 30982 -31932 31055
rect -56735 30914 -53619 30924
rect -56735 30910 -54990 30914
rect -56735 30907 -55127 30910
rect -56735 30887 -55272 30907
rect -65695 30814 -63845 30840
rect -55294 30826 -55272 30887
rect -55204 30829 -55127 30907
rect -55059 30833 -54990 30910
rect -54922 30833 -53619 30914
rect -46559 30897 -44611 30980
rect -46559 30880 -43339 30897
rect -55059 30829 -53619 30833
rect -55204 30826 -53619 30829
rect -65567 30573 -65419 30814
rect -55294 30807 -53619 30826
rect -44940 30875 -43339 30880
rect -44940 30872 -44651 30875
rect -44940 30871 -44805 30872
rect -67009 30425 -65294 30573
rect -64383 30033 -64306 30076
rect -64383 29974 -64374 30033
rect -64315 29981 -64306 30033
rect -64315 29974 -63672 29981
rect -64383 29904 -63672 29974
rect -61729 29941 -61138 30013
rect -64383 29884 -64306 29904
rect -64383 29825 -64376 29884
rect -64317 29825 -64306 29884
rect -64383 29810 -64306 29825
rect -55046 29373 -54889 30807
rect -44940 30798 -44932 30871
rect -44866 30799 -44805 30871
rect -44739 30802 -44651 30872
rect -44585 30802 -43339 30875
rect -36385 30853 -34420 30953
rect -32055 30903 -32039 30982
rect -31948 30903 -31932 30982
rect -18227 31095 -18207 31174
rect -18116 31095 -18104 31174
rect -18227 31022 -18104 31095
rect -18227 30943 -18211 31022
rect -18120 30943 -18104 31022
rect -4270 31146 -4250 31225
rect -4159 31146 -4147 31225
rect 28530 31229 28653 31243
rect -4270 31073 -4147 31146
rect -4270 30994 -4254 31073
rect -4163 30994 -4147 31073
rect -4270 30982 -4147 30994
rect 6690 31174 6813 31188
rect 6690 31095 6710 31174
rect 6801 31095 6813 31174
rect 28530 31150 28550 31229
rect 28641 31150 28653 31229
rect 6690 31022 6813 31095
rect -18227 30931 -18104 30943
rect 6690 30943 6706 31022
rect 6797 30943 6813 31022
rect 6690 30931 6813 30943
rect 17160 31119 17283 31133
rect 17160 31040 17180 31119
rect 17271 31040 17283 31119
rect 17160 30967 17283 31040
rect 28530 31077 28653 31150
rect 28530 30998 28546 31077
rect 28637 30998 28653 31077
rect 28530 30986 28653 30998
rect -32055 30891 -31932 30903
rect 17160 30888 17176 30967
rect 17267 30888 17283 30967
rect -44739 30799 -43339 30802
rect -44866 30798 -43339 30799
rect -44940 30780 -43339 30798
rect -53898 29974 -53800 29983
rect -53898 29973 -53640 29974
rect -53898 29898 -53884 29973
rect -53809 29898 -53640 29973
rect -51821 29934 -51099 30006
rect -53898 29897 -53640 29898
rect -53898 29796 -53800 29897
rect -53898 29795 -53798 29796
rect -53898 29718 -53884 29795
rect -53807 29718 -53798 29795
rect -53898 29717 -53798 29718
rect -53898 29708 -53800 29717
rect -56663 29216 -54889 29373
rect -44757 29342 -44633 30780
rect -34520 30712 -34420 30853
rect -7145 30823 -4298 30831
rect -11299 30792 -4298 30823
rect -25121 30767 -23102 30768
rect -25121 30752 -18374 30767
rect -25121 30750 -23091 30752
rect -34701 30708 -32073 30712
rect -34701 30698 -34550 30708
rect -34701 30615 -34681 30698
rect -34611 30625 -34550 30698
rect -34480 30706 -32073 30708
rect -34480 30625 -34422 30706
rect -34611 30623 -34422 30625
rect -34352 30623 -32073 30706
rect -25121 30668 -23377 30750
rect -23397 30667 -23377 30668
rect -23307 30667 -23227 30750
rect -23157 30669 -23091 30750
rect -23021 30669 -18374 30752
rect -11299 30732 -7140 30792
rect -7086 30789 -6869 30792
rect -7086 30732 -7002 30789
rect -11299 30729 -7002 30732
rect -6948 30732 -6869 30789
rect -6815 30732 -4298 30792
rect 2673 30809 4848 30887
rect 17160 30876 17283 30888
rect 2673 30787 5180 30809
rect -6948 30729 -4298 30732
rect -11299 30723 -4298 30729
rect -7145 30714 -4298 30723
rect 4748 30770 5180 30787
rect 4748 30740 6587 30770
rect 4748 30739 5127 30740
rect 4748 30736 4971 30739
rect -23157 30667 -18374 30669
rect -23397 30650 -18374 30667
rect -34611 30615 -32073 30623
rect -34701 30595 -32073 30615
rect -43726 29947 -43530 29959
rect -43726 29932 -43063 29947
rect -43726 29871 -43708 29932
rect -43648 29871 -43596 29932
rect -43537 29871 -43063 29932
rect -41183 29907 -40563 29979
rect -43726 29870 -43063 29871
rect -43726 29840 -43530 29870
rect -46471 29218 -44633 29342
rect -34534 29300 -34441 30595
rect -32322 29776 -31960 29809
rect -32322 29770 -32106 29776
rect -32322 29704 -32283 29770
rect -32222 29710 -32106 29770
rect -32045 29710 -31960 29776
rect -30082 29722 -29492 29794
rect -32222 29704 -31960 29710
rect -32322 29670 -31960 29704
rect -36081 29207 -34441 29300
rect -43404 29155 -43296 29171
rect -43404 29075 -43389 29155
rect -43309 29075 -43296 29155
rect -43404 29000 -43296 29075
rect -31849 29000 -31737 29279
rect -23249 29136 -23125 30650
rect -18480 30372 -18152 30389
rect -18480 30261 -18470 30372
rect -18359 30371 -18152 30372
rect -18359 30262 -18285 30371
rect -18176 30262 -18152 30371
rect -18359 30261 -18152 30262
rect -18480 30245 -18152 30261
rect -18994 29819 -18656 29852
rect -18994 29735 -18963 29819
rect -18879 29735 -18763 29819
rect -18679 29735 -18398 29819
rect -15442 29777 -14340 29849
rect -18994 29712 -18656 29735
rect -6988 29210 -6872 30714
rect 4748 30709 4839 30736
rect 4833 30672 4839 30709
rect 4895 30675 4971 30736
rect 5027 30676 5127 30739
rect 5183 30676 6587 30740
rect 13647 30728 15692 30826
rect 26010 30784 28484 30799
rect 24542 30765 28484 30784
rect 24542 30762 26181 30765
rect 13647 30726 17544 30728
rect 5027 30675 6587 30676
rect 4895 30672 6587 30675
rect 4833 30653 6587 30672
rect 15304 30696 17544 30726
rect 15304 30690 15459 30696
rect -4538 29908 -4222 29931
rect -4538 29824 -4486 29908
rect -4402 29907 -4222 29908
rect -4402 29825 -4322 29907
rect -4240 29825 -4222 29907
rect -2687 29841 -1724 29913
rect -4402 29824 -4222 29825
rect -4538 29801 -4222 29824
rect 4962 29277 5122 30653
rect 15304 30634 15339 30690
rect 15391 30640 15459 30690
rect 15511 30640 15595 30696
rect 15647 30640 17544 30696
rect 24542 30699 26049 30762
rect 26109 30702 26181 30762
rect 26241 30762 28484 30765
rect 26241 30702 26315 30762
rect 26109 30699 26315 30702
rect 26375 30699 28484 30762
rect 24542 30684 28484 30699
rect 26010 30682 28484 30684
rect 15391 30634 17544 30640
rect 15304 30611 17544 30634
rect 6045 30367 6502 30406
rect 6045 30256 6064 30367
rect 6175 30366 6502 30367
rect 6175 30257 6367 30366
rect 6476 30257 6502 30366
rect 6175 30256 6502 30257
rect 6045 30244 6502 30256
rect 6409 29838 6753 29857
rect 6409 29837 6631 29838
rect 6409 29735 6427 29837
rect 6529 29735 6631 29837
rect 6409 29734 6631 29735
rect 6735 29734 6753 29838
rect 8487 29780 9560 29852
rect 6409 29713 6753 29734
rect -25033 29012 -23125 29136
rect -11207 29094 -6872 29210
rect 2742 29117 5122 29277
rect 15391 29210 15534 30611
rect 17440 30304 17538 30329
rect 17440 30238 17459 30304
rect 17525 30238 17538 30304
rect 17440 30138 17538 30238
rect 17440 30070 17458 30138
rect 17526 30070 17538 30138
rect 17440 30055 17538 30070
rect 17636 29778 17749 29810
rect 17258 29701 17413 29778
rect 17636 29701 17655 29778
rect 17732 29701 17749 29778
rect 19283 29738 20166 29810
rect 17636 29632 17749 29701
rect 17636 29555 17646 29632
rect 17724 29555 17749 29632
rect 17636 29532 17749 29555
rect 13725 29067 15534 29210
rect 26174 29169 26323 30682
rect 27918 30555 28036 30569
rect 27918 30469 27932 30555
rect 28018 30469 28036 30555
rect 27918 30393 28036 30469
rect 27918 30305 27936 30393
rect 28024 30305 28291 30393
rect 27918 30282 28036 30305
rect 28441 29848 28564 29865
rect 28441 29773 28460 29848
rect 28540 29773 28564 29848
rect 30643 29809 31566 29881
rect 28441 29684 28564 29773
rect 28441 29607 28462 29684
rect 28539 29607 28564 29684
rect 28441 29587 28564 29607
rect 24617 29020 29248 29169
rect -43404 28987 -31737 29000
rect -43654 28969 -43544 28983
rect -43654 28887 -43642 28969
rect -43560 28887 -43544 28969
rect -43404 28905 -43390 28987
rect -43308 28905 -31737 28987
rect -43404 28888 -31737 28905
rect -43654 28778 -43544 28887
rect 17427 28832 17529 28836
rect 28731 28833 28849 28856
rect 28731 28832 28754 28833
rect 17423 28824 28754 28832
rect -32436 28778 -32074 28792
rect -43654 28777 -32207 28778
rect -43654 28759 -32427 28777
rect -43654 28677 -43642 28759
rect -43560 28677 -32427 28759
rect -43654 28667 -32427 28677
rect -32317 28667 -32207 28777
rect -43654 28666 -32207 28667
rect -32095 28666 -32074 28778
rect -32436 28653 -32074 28666
rect -4055 28742 -3896 28762
rect -4055 28631 -4030 28742
rect -3919 28631 -3896 28742
rect 17423 28741 17439 28824
rect 17522 28749 28754 28824
rect 28820 28749 28849 28833
rect 17522 28741 28849 28749
rect 17423 28732 28849 28741
rect -18489 28532 -18088 28550
rect -4055 28532 -3896 28631
rect 17427 28677 17529 28732
rect 17427 28590 17439 28677
rect 17522 28590 17529 28677
rect 17427 28578 17529 28590
rect 28731 28696 28849 28732
rect 28731 28612 28756 28696
rect 28822 28612 28849 28696
rect 28731 28579 28849 28612
rect -18489 28421 -18470 28532
rect -18359 28421 -18221 28532
rect -18110 28531 -3896 28532
rect -18110 28422 -4030 28531
rect -3921 28422 -3896 28531
rect -18110 28421 -3896 28422
rect -18489 28406 -18088 28421
rect -4055 28402 -3896 28421
rect 6411 28470 6782 28486
rect 18511 28470 18650 28480
rect 6411 28469 6658 28470
rect 6049 28351 6188 28369
rect 6411 28367 6432 28469
rect 6534 28367 6658 28469
rect 6411 28366 6658 28367
rect 6762 28460 18650 28470
rect 6762 28366 18531 28460
rect 6411 28351 6782 28366
rect 18511 28356 18531 28366
rect 18635 28356 18650 28460
rect 6049 28240 6064 28351
rect 6175 28240 6188 28351
rect -4497 28170 -4388 28187
rect -4497 28086 -4486 28170
rect -4402 28086 -4388 28170
rect -18981 28006 -18651 28021
rect -4497 28006 -4388 28086
rect -18981 27922 -18963 28006
rect -18879 27922 -18739 28006
rect -18655 28005 -4388 28006
rect -18655 27923 -4485 28005
rect -4403 27923 -4388 28005
rect 6049 28100 6188 28240
rect 18511 28277 18650 28356
rect 18511 28175 18532 28277
rect 18634 28175 18650 28277
rect 18511 28158 18650 28175
rect 17881 28100 18025 28105
rect 6049 28099 18025 28100
rect 6049 27990 6065 28099
rect 6174 28036 18025 28099
rect 6174 27990 17899 28036
rect 6049 27989 17899 27990
rect 6049 27972 6188 27989
rect -18655 27922 -4388 27923
rect -18981 27901 -18651 27922
rect -4497 27906 -4388 27922
rect 17881 27925 17899 27989
rect 18010 27925 18025 28036
rect 17881 27787 18025 27925
rect -19720 27625 -19576 27734
rect 17881 27678 17900 27787
rect 18009 27678 18025 27787
rect 17881 27658 18025 27678
rect 27539 27809 27685 27894
rect 27539 27714 27567 27809
rect 27650 27714 27685 27809
rect -19720 27552 -19700 27625
rect -19604 27552 -19576 27625
rect -19720 27513 -19576 27552
rect 27539 27576 27685 27714
rect 27539 27513 27571 27576
rect -19720 27486 27571 27513
rect -19720 27458 -5692 27486
rect -19720 27385 -19696 27458
rect -19600 27405 -5692 27458
rect -5591 27481 27571 27486
rect 27654 27481 27685 27576
rect -5591 27405 27685 27481
rect -19600 27385 27685 27405
rect -19720 27367 27685 27385
rect -19720 27362 -19576 27367
rect -5715 27251 -5569 27367
rect -5715 27170 -5692 27251
rect -5591 27170 -5569 27251
rect -5715 27142 -5569 27170
rect 28441 27292 28566 27323
rect 28441 27197 28462 27292
rect 28557 27197 28566 27292
rect 17619 27140 17734 27152
rect 17619 27137 17631 27140
rect 17724 27137 17734 27140
rect 28441 27137 28566 27197
rect 17619 27042 17630 27137
rect 17725 27136 28566 27137
rect 17725 27043 28463 27136
rect 28556 27043 28566 27136
rect 17725 27042 28566 27043
rect 17619 26970 17734 27042
rect 28441 27009 28566 27042
rect 17619 26875 17630 26970
rect 17725 26875 17734 26970
rect 17619 26867 17734 26875
rect -10810 26764 -9132 26791
rect -10810 26761 -9213 26764
rect -10810 26695 -9349 26761
rect -9295 26698 -9213 26761
rect -9159 26698 -9132 26764
rect -9295 26695 -9132 26698
rect -10810 26667 -9132 26695
rect -64377 26583 -64305 26608
rect -64377 26581 -64367 26583
rect -64381 26530 -64367 26581
rect -64313 26581 -64305 26583
rect -64313 26530 -63781 26581
rect -64381 26507 -63781 26530
rect -53898 26515 -53804 26526
rect -64381 26476 -64305 26507
rect -64381 26423 -64368 26476
rect -64314 26423 -64305 26476
rect -64381 26368 -64305 26423
rect -64381 26315 -64370 26368
rect -64316 26315 -64305 26368
rect -64381 26295 -64305 26315
rect -53898 26443 -53886 26515
rect -53814 26503 -53804 26515
rect -53814 26443 -53475 26503
rect -53898 26429 -53475 26443
rect -53898 26379 -53804 26429
rect -53898 26307 -53886 26379
rect -53814 26307 -53804 26379
rect -53898 26297 -53804 26307
rect -64381 26293 -64307 26295
rect -56702 26230 -54888 26253
rect -56702 26129 -55284 26230
rect -55214 26229 -54888 26230
rect -55214 26227 -55004 26229
rect -55214 26129 -55150 26227
rect -56702 26126 -55150 26129
rect -55080 26128 -55004 26227
rect -54934 26128 -54888 26229
rect -55080 26126 -54888 26128
rect -56702 26118 -54888 26126
rect -46328 26144 -40201 26182
rect -46328 26054 -44927 26144
rect -44861 26142 -44645 26144
rect -44861 26054 -44783 26142
rect -46328 26052 -44783 26054
rect -44717 26054 -44645 26142
rect -44579 26054 -40201 26144
rect -44717 26052 -40201 26054
rect -46328 26025 -40201 26052
rect -35987 26140 -34297 26169
rect -35987 26138 -34391 26140
rect -35987 26063 -34687 26138
rect -34625 26135 -34391 26138
rect -34625 26063 -34553 26135
rect -35987 26060 -34553 26063
rect -34491 26065 -34391 26135
rect -34329 26065 -34297 26140
rect -34491 26060 -34297 26065
rect -35987 26045 -34297 26060
rect -33717 26134 -33408 26152
rect -33717 26133 -33502 26134
rect -33717 26061 -33703 26133
rect -33631 26061 -33502 26133
rect -33717 26060 -33502 26061
rect -33428 26060 -32657 26134
rect -33717 26045 -33408 26060
rect -64110 25880 -64040 25930
rect -10810 25885 -10686 26667
rect 14069 26441 15726 26460
rect -5360 26380 -5270 26430
rect -5389 26361 -5113 26380
rect 14069 26365 15331 26441
rect 15402 26365 15484 26441
rect 15555 26438 15726 26441
rect 15555 26365 15637 26438
rect 14069 26362 15637 26365
rect 15708 26362 15726 26438
rect 18530 26390 18630 26610
rect 28166 26494 28576 26510
rect 28166 26493 28441 26494
rect -5389 26360 -5197 26361
rect -5389 26288 -5373 26360
rect -5301 26288 -5197 26360
rect -5389 26287 -5197 26288
rect -5123 26287 -4657 26361
rect 14069 26348 15726 26362
rect 28166 26376 28178 26493
rect 28295 26376 28441 26493
rect 28166 26375 28441 26376
rect 28560 26375 28576 26494
rect 28166 26361 28576 26375
rect -5389 26274 -5113 26287
rect -5360 26260 -5270 26274
rect -9708 26211 -7503 26245
rect -9708 26205 -7615 26211
rect -9708 26200 -7764 26205
rect -9708 26147 -7904 26200
rect -7852 26152 -7764 26200
rect -7712 26158 -7615 26205
rect -7563 26158 -7503 26211
rect -7712 26152 -7503 26158
rect -7852 26147 -7503 26152
rect 24767 26165 29113 26209
rect 24767 26162 26165 26165
rect -9708 26132 -7503 26147
rect 9095 26057 9603 26150
rect 24767 26087 26025 26162
rect 26084 26090 26165 26162
rect 26224 26090 26312 26165
rect 26371 26090 29113 26165
rect 26084 26087 29113 26090
rect 24767 26075 29113 26087
rect 2379 26025 9603 26057
rect 2379 26021 5134 26025
rect -9420 25965 -9188 25978
rect -9420 25961 -9271 25965
rect -9420 25907 -9399 25961
rect -9345 25909 -9271 25961
rect -9215 25909 -9188 25965
rect -9345 25907 -9188 25909
rect -9420 25904 -9188 25907
rect 2379 25923 4846 26021
rect 4915 26020 5134 26021
rect 4915 25923 4986 26020
rect 2379 25922 4986 25923
rect 5055 25927 5134 26020
rect 5203 25998 9603 26025
rect 5203 25927 9247 25998
rect 5055 25922 9247 25927
rect 2379 25905 9247 25922
rect 17881 25964 18020 26001
rect -64144 25870 -63833 25880
rect -64144 25813 -64112 25870
rect -64054 25813 -63833 25870
rect -64144 25769 -63833 25813
rect -10810 25842 -10477 25885
rect -9757 25854 -9188 25904
rect -9757 25849 -9269 25854
rect -53595 25781 -53134 25802
rect -53595 25775 -53446 25781
rect -64144 25758 -64033 25769
rect -64144 25701 -64113 25758
rect -64055 25701 -64033 25758
rect -64144 25645 -64033 25701
rect -53595 25717 -53594 25775
rect -53536 25723 -53446 25775
rect -53388 25723 -53134 25781
rect -53536 25717 -53134 25723
rect -53595 25691 -53134 25717
rect -25548 25787 -16062 25808
rect -25548 25785 -23087 25787
rect -25548 25782 -23236 25785
rect -25548 25670 -23387 25782
rect -23311 25673 -23236 25782
rect -23160 25675 -23087 25785
rect -23011 25675 -16062 25787
rect -10810 25761 -10465 25842
rect -9757 25825 -9399 25849
rect -9679 25803 -9399 25825
rect -9420 25793 -9399 25803
rect -9343 25800 -9269 25849
rect -9215 25800 -9188 25854
rect 17881 25855 17897 25964
rect 18006 25855 18020 25964
rect -9343 25793 -9188 25800
rect -9420 25788 -9188 25793
rect 17490 25729 17688 25840
rect 17881 25750 18020 25855
rect -23160 25673 -16062 25675
rect -23311 25670 -16062 25673
rect -25548 25659 -16062 25670
rect -25548 25658 -16049 25659
rect -64144 25588 -64114 25645
rect -64056 25588 -64033 25645
rect -16135 25613 -16049 25658
rect -64144 25552 -64033 25588
rect -4766 25549 -4485 25660
rect 17881 25639 17896 25750
rect 18007 25639 18020 25750
rect 17881 25616 18020 25639
rect 28572 25924 28712 25948
rect 28572 25815 28588 25924
rect 28697 25815 28712 25924
rect 28572 25654 28712 25815
rect -11464 25503 -6734 25545
rect -11464 25450 -7118 25503
rect -7066 25450 -6985 25503
rect -6933 25498 -6734 25503
rect -6933 25450 -6844 25498
rect -11464 25445 -6844 25450
rect -6792 25445 -6734 25498
rect -32835 25322 -32445 25433
rect -11464 25431 -6734 25445
rect 4061 25499 6607 25546
rect 28572 25543 28587 25654
rect 28698 25543 28712 25654
rect 28572 25536 28712 25543
rect 4061 25496 4374 25499
rect 4061 25493 4224 25496
rect -11458 25380 -11344 25431
rect 4061 25427 4084 25493
rect 4150 25430 4224 25493
rect 4290 25433 4374 25496
rect 4440 25433 6607 25499
rect 4290 25430 6607 25433
rect 4150 25427 6607 25430
rect 4061 25396 6607 25427
rect -24190 25270 -19145 25310
rect -45756 25206 -43545 25249
rect -45756 25205 -45608 25206
rect -45756 25127 -45746 25205
rect -45674 25128 -45608 25205
rect -45536 25128 -45474 25206
rect -45402 25128 -43545 25206
rect -24190 25180 -24150 25270
rect -24060 25186 -23920 25270
rect -23829 25186 -19145 25270
rect -24060 25180 -19145 25186
rect -24190 25160 -19145 25180
rect -45674 25127 -43545 25128
rect -45756 25099 -43545 25127
rect 7039 25142 7162 25156
rect 7039 25063 7059 25142
rect 7150 25063 7162 25142
rect 7039 24990 7162 25063
rect 7039 24911 7055 24990
rect 7146 24911 7162 24990
rect -18635 24891 -18512 24905
rect 7039 24899 7162 24911
rect -43024 24853 -42901 24867
rect -43024 24774 -43004 24853
rect -42913 24774 -42901 24853
rect -43024 24701 -42901 24774
rect -43024 24622 -43008 24701
rect -42917 24622 -42901 24701
rect -18635 24812 -18615 24891
rect -18524 24812 -18512 24891
rect -18635 24739 -18512 24812
rect -18635 24660 -18619 24739
rect -18528 24660 -18512 24739
rect -18635 24648 -18512 24660
rect -43024 24610 -42901 24622
rect -5056 24230 -4677 24244
rect -5056 24119 -5043 24230
rect -4932 24229 -4291 24230
rect -4932 24120 -4794 24229
rect -4685 24120 -4291 24229
rect -4932 24119 -4291 24120
rect -5056 24106 -4677 24119
rect 5556 24101 5745 24109
rect 5556 24044 5684 24101
rect 5737 24075 5745 24101
rect 5737 24044 6430 24075
rect 5556 24035 6430 24044
rect -32970 24003 -32599 24028
rect -32970 23892 -32950 24003
rect -32839 24002 -32213 24003
rect -32839 23893 -32723 24002
rect -32614 23893 -32213 24002
rect -32839 23892 -32213 23893
rect 5556 23978 5571 24035
rect 5624 24001 6430 24035
rect 5624 23978 5745 24001
rect 5556 23948 5745 23978
rect -32970 23872 -32599 23892
rect 5556 23891 5678 23948
rect 5731 23891 5745 23948
rect -43681 23806 -43519 23849
rect -66371 23723 -66012 23728
rect -66371 23722 -66231 23723
rect -66380 23720 -66231 23722
rect -66380 23702 -66363 23720
rect -66831 23657 -66363 23702
rect -66303 23660 -66231 23720
rect -66171 23722 -66012 23723
rect -66171 23720 -63957 23722
rect -66171 23660 -66097 23720
rect -66303 23657 -66097 23660
rect -66037 23657 -63957 23720
rect -66831 23640 -63957 23657
rect -43681 23694 -43648 23806
rect -43539 23694 -43519 23806
rect -66831 23554 -66096 23640
rect -55937 23636 -53572 23644
rect -55937 23633 -55653 23636
rect -55937 23630 -55787 23633
rect -55937 23572 -55922 23630
rect -55864 23575 -55787 23630
rect -55729 23578 -55653 23633
rect -55595 23578 -53572 23636
rect -55729 23575 -53572 23578
rect -55864 23572 -53572 23575
rect -55937 23562 -53572 23572
rect -43681 23569 -43519 23694
rect -43681 23457 -43656 23569
rect -43547 23457 -43519 23569
rect -19635 23839 -19480 23883
rect 5556 23870 5745 23891
rect -19635 23815 -19268 23839
rect -19635 23758 -19606 23815
rect -19517 23765 -19268 23815
rect 5556 23813 5574 23870
rect 5627 23813 5745 23870
rect 5556 23799 5745 23813
rect -19517 23758 -19480 23765
rect -19635 23695 -19480 23758
rect -19635 23638 -19605 23695
rect -19516 23638 -19480 23695
rect -19635 23586 -19480 23638
rect 14617 23673 17515 23682
rect 14617 23617 14654 23673
rect 14706 23672 17515 23673
rect 14706 23617 14782 23672
rect 14617 23616 14782 23617
rect 14834 23671 17515 23672
rect 14834 23616 14921 23671
rect 14617 23615 14921 23616
rect 14973 23615 17515 23671
rect 14617 23600 17515 23615
rect 25325 23614 28213 23620
rect 25325 23611 25480 23614
rect -19635 23529 -19606 23586
rect -19517 23529 -19480 23586
rect 25325 23548 25348 23611
rect 25408 23551 25480 23611
rect 25540 23611 28213 23614
rect 25540 23551 25614 23611
rect 25408 23548 25614 23551
rect 25674 23548 28213 23611
rect 25325 23538 28213 23548
rect -19635 23510 -19480 23529
rect -43681 23420 -43519 23457
rect -7914 23493 -4853 23502
rect -7914 23490 -7640 23493
rect -7914 23486 -7776 23490
rect -7914 23429 -7897 23486
rect -7845 23433 -7776 23486
rect -7724 23436 -7640 23490
rect -7588 23436 -4853 23493
rect -7724 23433 -4853 23436
rect -7845 23429 -4853 23433
rect -7914 23420 -4853 23429
rect -35391 23261 -32795 23275
rect -35391 23260 -35240 23261
rect -35391 23200 -35376 23260
rect -35316 23201 -35240 23260
rect -35180 23201 -35086 23261
rect -35026 23201 -32795 23261
rect -35316 23200 -32795 23201
rect -35391 23193 -32795 23200
rect 6708 23211 6831 23225
rect 6708 23132 6728 23211
rect 6819 23132 6831 23211
rect 6708 23059 6831 23132
rect 6708 22980 6724 23059
rect 6815 22980 6831 23059
rect -19049 22965 -18926 22979
rect 6708 22968 6831 22980
rect -62649 22870 -62603 22961
rect -43323 22913 -43200 22927
rect -66722 22822 -66566 22858
rect -68368 22803 -68034 22819
rect -68368 22714 -68348 22803
rect -68263 22714 -68034 22803
rect -68368 22696 -68034 22714
rect -66722 22748 -66681 22822
rect -66602 22748 -66566 22822
rect -66722 22702 -66566 22748
rect -43323 22834 -43303 22913
rect -43212 22834 -43200 22913
rect -43323 22761 -43200 22834
rect -43323 22682 -43307 22761
rect -43216 22682 -43200 22761
rect -19049 22886 -19029 22965
rect -18938 22886 -18926 22965
rect -19049 22813 -18926 22886
rect -19049 22734 -19033 22813
rect -18942 22734 -18926 22813
rect -19049 22722 -18926 22734
rect 4837 22739 6655 22771
rect 4837 22738 5132 22739
rect 4837 22737 4991 22738
rect -43323 22670 -43200 22682
rect 4837 22675 4847 22737
rect 4911 22676 4991 22737
rect 5055 22677 5132 22738
rect 5196 22677 6655 22739
rect 13683 22727 15620 22827
rect 5055 22676 6655 22677
rect 4911 22675 6655 22676
rect -52264 22590 -52218 22669
rect 4837 22654 6655 22675
rect -23377 22535 -23260 22543
rect -23136 22535 -23019 22547
rect -23397 22530 -18824 22535
rect -44937 22441 -43478 22474
rect -44937 22439 -44681 22441
rect -44937 22437 -44806 22439
rect -44937 22381 -44926 22437
rect -44874 22383 -44806 22437
rect -44754 22385 -44681 22439
rect -44629 22385 -43478 22441
rect -36385 22430 -34294 22530
rect -23397 22526 -23124 22530
rect -23397 22436 -23365 22526
rect -23275 22440 -23124 22526
rect -23034 22440 -18824 22530
rect -12009 22490 -6879 22590
rect -23275 22436 -18824 22440
rect -44754 22383 -43478 22385
rect -44874 22381 -43478 22383
rect -44937 22357 -43478 22381
rect -67016 22046 -65432 22194
rect -65580 21307 -65432 22046
rect -56308 21619 -56195 21642
rect -56308 21547 -56286 21619
rect -56214 21547 -56195 21619
rect -65696 21294 -63890 21307
rect -65696 21291 -65540 21294
rect -65696 21228 -65672 21291
rect -65612 21231 -65540 21291
rect -65480 21291 -63890 21294
rect -65480 21231 -65406 21291
rect -65612 21228 -65406 21231
rect -65346 21228 -63890 21291
rect -65696 21194 -63890 21228
rect -67610 21171 -67487 21188
rect -66929 21171 -66806 21188
rect -67610 21081 -67592 21171
rect -67502 21170 -66806 21171
rect -67502 21082 -66912 21170
rect -66824 21082 -66806 21170
rect -67502 21081 -66806 21082
rect -67610 21058 -67487 21081
rect -66929 21058 -66806 21081
rect -63021 20680 -62787 21016
rect -56308 21004 -56195 21547
rect -53370 21562 -53180 21571
rect -53370 21507 -53361 21562
rect -53306 21507 -53250 21562
rect -53195 21507 -53180 21562
rect -53370 21498 -53180 21507
rect -44771 21245 -44618 22357
rect -55292 21195 -53297 21229
rect -55292 21193 -54999 21195
rect -55292 21192 -55145 21193
rect -55292 21137 -55278 21192
rect -55223 21138 -55145 21192
rect -55090 21140 -54999 21193
rect -54944 21140 -53297 21195
rect -55090 21138 -53297 21140
rect -55223 21137 -53297 21138
rect -55292 21116 -53297 21137
rect -46318 21092 -44618 21245
rect -53902 21004 -53803 21024
rect -56308 20990 -53803 21004
rect -56308 20935 -53876 20990
rect -53821 20935 -53803 20990
rect -56308 20891 -53803 20935
rect -53902 20857 -53803 20891
rect -53902 20802 -53875 20857
rect -53820 20802 -53803 20857
rect -53902 20776 -53803 20802
rect -53694 20724 -53597 20755
rect -53694 20680 -53675 20724
rect -63021 20669 -53675 20680
rect -53620 20669 -53597 20724
rect -63021 20591 -53597 20669
rect -63021 20567 -53674 20591
rect -53694 20536 -53674 20567
rect -53619 20536 -53597 20591
rect -43344 20560 -43231 21528
rect -41668 21484 -40444 21556
rect -34476 20909 -34376 22430
rect -23397 22418 -18824 22436
rect -31487 22208 -31441 22298
rect -32637 21201 -32400 21211
rect -32637 21194 -32602 21201
rect -32847 21148 -32602 21194
rect -32550 21194 -32400 21201
rect -32550 21148 -32487 21194
rect -32847 21141 -32487 21148
rect -32435 21141 -32400 21194
rect -32847 21137 -32400 21141
rect -32637 21120 -32400 21137
rect -36282 20860 -34376 20909
rect -36282 20831 -32677 20860
rect -23223 20857 -23110 22418
rect -19224 21575 -18883 21612
rect -19224 21571 -18989 21575
rect -19224 21499 -19197 21571
rect -19131 21503 -18989 21571
rect -18923 21503 -18883 21575
rect -16493 21545 -15939 21617
rect -19131 21499 -18883 21503
rect -19224 21452 -18883 21499
rect -6979 21087 -6879 22490
rect -3559 22456 -3513 22537
rect -4829 21413 -4509 21470
rect -4829 21408 -4636 21413
rect -4829 21344 -4813 21408
rect -4751 21349 -4636 21408
rect -4574 21349 -4509 21413
rect -4751 21344 -4509 21349
rect -4829 21294 -4509 21344
rect -7143 21058 -4434 21087
rect 4978 21059 5096 22654
rect 6063 22348 6174 22354
rect 6063 22347 6658 22348
rect 6063 22281 6085 22347
rect 6151 22281 6658 22347
rect 6063 22280 6658 22281
rect 6063 22192 6174 22280
rect 6063 22124 6084 22192
rect 6152 22124 6174 22192
rect 6063 22118 6174 22124
rect 6418 21824 6751 21850
rect 6418 21720 6426 21824
rect 6530 21823 6751 21824
rect 6530 21721 6637 21823
rect 6739 21721 6751 21823
rect 8940 21781 9830 21853
rect 6530 21720 6751 21721
rect 6418 21704 6751 21720
rect 15520 21267 15620 22727
rect 18820 22616 18866 22720
rect 29516 22551 29562 22662
rect 17638 21601 17856 21611
rect 17638 21600 17790 21601
rect 17638 21545 17650 21600
rect 17705 21545 17790 21600
rect 17638 21544 17790 21545
rect 17847 21544 17856 21601
rect 17638 21535 17856 21544
rect 28479 21538 28564 21552
rect 28479 21483 28493 21538
rect 28548 21483 28564 21538
rect 28479 21419 28564 21483
rect 28479 21364 28493 21419
rect 28548 21364 28564 21419
rect 28479 21343 28564 21364
rect 13729 21232 17792 21267
rect 13729 21228 15443 21232
rect 13729 21172 15336 21228
rect 15388 21176 15443 21228
rect 15495 21228 17792 21232
rect 15495 21176 15568 21228
rect 15388 21172 15568 21176
rect 15620 21172 17792 21228
rect 13729 21154 17792 21172
rect 24780 21180 28313 21205
rect 24780 21177 26174 21180
rect 24780 21114 26042 21177
rect 26102 21117 26174 21177
rect 26234 21177 28313 21180
rect 26234 21117 26308 21177
rect 26102 21114 26308 21117
rect 26368 21114 28313 21177
rect 24780 21092 28313 21114
rect -7143 21054 -6859 21058
rect -7143 21000 -7120 21054
rect -7064 21000 -6990 21054
rect -6934 21004 -6859 21054
rect -6803 21004 -4434 21058
rect -6934 21000 -4434 21004
rect -7143 20989 -4434 21000
rect -36282 20827 -34399 20831
rect -36282 20824 -34543 20827
rect -36282 20815 -34682 20824
rect -34698 20762 -34682 20815
rect -34623 20765 -34543 20824
rect -34484 20769 -34399 20827
rect -34340 20769 -32677 20831
rect -34484 20765 -32677 20769
rect -34623 20762 -32677 20765
rect -34698 20747 -32677 20762
rect -25521 20744 -23110 20857
rect -11929 20974 -4434 20989
rect -11929 20848 -6757 20974
rect 2404 20941 5096 21059
rect 6052 21019 6189 21040
rect 6052 20907 6064 21019
rect 6175 20907 6189 21019
rect 6052 20793 6189 20907
rect -33718 20650 -33607 20670
rect -33718 20590 -33690 20650
rect -33630 20590 -33607 20650
rect -33718 20560 -33607 20590
rect -53694 20504 -53597 20536
rect -53209 20538 -33607 20560
rect -53209 20481 -53173 20538
rect -53113 20481 -53058 20538
rect -52998 20510 -33607 20538
rect -52998 20481 -33690 20510
rect -53209 20450 -33690 20481
rect -33630 20450 -33607 20510
rect -53209 20447 -33607 20450
rect -33718 20430 -33607 20447
rect -33253 20530 -33142 20570
rect -4941 20557 -4785 20782
rect -3870 20680 -3670 20790
rect 6052 20679 6064 20793
rect 6175 20792 6189 20793
rect 28153 20863 28487 20902
rect 28153 20792 28942 20863
rect 6175 20681 28942 20792
rect 6175 20679 6189 20681
rect 6052 20668 6189 20679
rect -33253 20470 -33230 20530
rect -33170 20470 -33142 20530
rect -33253 20410 -33142 20470
rect -43092 20351 -42762 20362
rect -33253 20351 -33230 20410
rect -52615 20350 -42887 20351
rect -52615 20336 -43080 20350
rect -52615 20279 -52583 20336
rect -52523 20279 -52468 20336
rect -52408 20279 -43080 20336
rect -52615 20239 -43080 20279
rect -42969 20239 -42887 20350
rect -52615 20238 -42887 20239
rect -42774 20350 -33230 20351
rect -33170 20350 -33142 20410
rect -32840 20533 -4785 20557
rect -32840 20530 -22103 20533
rect -32840 20463 -22292 20530
rect -22216 20466 -22103 20530
rect -22027 20466 -4785 20533
rect -22216 20463 -4785 20466
rect -32840 20401 -4785 20463
rect 6416 20584 6543 20595
rect 6416 20480 6426 20584
rect 6530 20532 6543 20584
rect 28455 20532 28838 20546
rect 6530 20531 28838 20532
rect 6530 20480 28464 20531
rect 6416 20422 28464 20480
rect 28573 20422 28713 20531
rect 28822 20422 28838 20531
rect 6416 20421 28838 20422
rect -42774 20330 -33142 20350
rect 6416 20346 6543 20421
rect 28455 20408 28838 20421
rect -42774 20238 -33148 20330
rect 6416 20244 6427 20346
rect 6529 20244 6543 20346
rect -43092 20230 -42762 20238
rect -32642 20231 -32358 20243
rect -42888 20229 -42773 20230
rect -32642 20228 -32446 20231
rect -32642 20175 -32610 20228
rect -32558 20178 -32446 20228
rect -32394 20221 -32358 20231
rect -4832 20221 -4521 20241
rect 6416 20231 6543 20244
rect -32394 20179 -4521 20221
rect -32394 20178 -21949 20179
rect -32558 20175 -21949 20178
rect -32642 20112 -21949 20175
rect -21873 20112 -21783 20179
rect -21707 20177 -4521 20179
rect -21707 20124 -4796 20177
rect -4740 20175 -4521 20177
rect -4740 20124 -4649 20175
rect -21707 20122 -4649 20124
rect -4593 20122 -4521 20175
rect -21707 20112 -4521 20122
rect -32642 20085 -4521 20112
rect -4832 20053 -4521 20085
rect 18270 19864 18676 19877
rect -18839 19863 18527 19864
rect -18839 19820 18278 19863
rect -18839 19817 -18672 19820
rect -18839 19761 -18824 19817
rect -18767 19764 -18672 19817
rect -18615 19764 18278 19820
rect -18767 19761 18278 19764
rect -18839 19748 18278 19761
rect -18839 19728 -5026 19748
rect -5053 19668 -5026 19728
rect -4954 19729 18278 19748
rect 18412 19729 18527 19863
rect -4954 19728 18527 19729
rect 18663 19728 18676 19864
rect -4954 19668 -4924 19728
rect 18270 19716 18676 19728
rect -5377 19538 -5248 19572
rect -5377 19523 -5347 19538
rect -19113 19479 -5347 19523
rect -19113 19476 -18946 19479
rect -19113 19420 -19098 19476
rect -19041 19423 -18946 19476
rect -18889 19458 -5347 19479
rect -5275 19523 -5248 19538
rect -5053 19547 -4924 19668
rect -5275 19458 -5246 19523
rect -18889 19423 -5246 19458
rect -5053 19467 -5023 19547
rect -4951 19467 -4924 19547
rect 17632 19539 17768 19578
rect 17632 19536 17656 19539
rect -5053 19438 -4924 19467
rect -4674 19459 17656 19536
rect 17738 19459 17768 19539
rect -19041 19420 -5246 19423
rect -19113 19387 -5246 19420
rect -5382 19330 -5246 19387
rect -4674 19400 17768 19459
rect -4674 19330 -4538 19400
rect -5382 19325 -4538 19330
rect -5382 19245 -5344 19325
rect -5272 19245 -4538 19325
rect 17632 19367 17768 19400
rect 17632 19287 17656 19367
rect 17738 19287 17768 19367
rect -19637 19199 -19478 19241
rect -19637 19093 -19604 19199
rect -19511 19093 -19478 19199
rect -5382 19194 -4538 19245
rect 5563 19200 5741 19259
rect 17632 19256 17768 19287
rect 5563 19116 5587 19200
rect 5719 19116 5741 19200
rect 5563 19112 5741 19116
rect -19637 19022 -19478 19093
rect -19637 18954 -19603 19022
rect -19508 18954 -19478 19022
rect -19637 18916 -19478 18954
rect -54131 18906 -19478 18916
rect -54190 18875 -19478 18906
rect -54190 18808 -54148 18875
rect -54063 18859 -19478 18875
rect -54063 18808 -19596 18859
rect -54190 18769 -19596 18808
rect -19505 18769 -19478 18859
rect -54190 18757 -19478 18769
rect -54190 18744 -54017 18757
rect -54190 18635 -54150 18744
rect -54048 18635 -54017 18744
rect -19637 18743 -19478 18757
rect -19111 18919 -5718 19097
rect -54190 18505 -54017 18635
rect -54190 18396 -54158 18505
rect -54056 18396 -54017 18505
rect -19111 18482 -18933 18919
rect -5896 18827 -5718 18919
rect -4233 19046 5741 19112
rect -4233 18962 5591 19046
rect 5723 18962 5741 19046
rect -4233 18934 5741 18962
rect -4233 18827 -4055 18934
rect -5896 18649 -4055 18827
rect -72156 18176 -72081 18374
rect -54190 18354 -54017 18396
rect -43412 18423 -43229 18450
rect -43412 18322 -43384 18423
rect -43283 18322 -43229 18423
rect -43412 18231 -43229 18322
rect -43412 18130 -43367 18231
rect -43266 18130 -43229 18231
rect -43412 18083 -43229 18130
rect -64604 18077 -43229 18083
rect -64663 18056 -43229 18077
rect -64663 17955 -43377 18056
rect -43276 17955 -43229 18056
rect -64663 17925 -43229 17955
rect -64663 17820 -64639 17925
rect -64565 17900 -43229 17925
rect -42919 18304 -18933 18482
rect -64565 17820 -64523 17900
rect -64663 17708 -64523 17820
rect -64663 17603 -64633 17708
rect -64559 17603 -64523 17708
rect -64663 17565 -64523 17603
rect -42919 17586 -42741 18304
rect 27209 17778 27413 17842
rect 27209 17660 27251 17778
rect 27369 17660 27413 17778
rect 27209 17606 27413 17660
rect -43841 17585 -42741 17586
rect -43913 17557 -42741 17585
rect -43913 17498 -43887 17557
rect -43780 17498 -42741 17557
rect -43913 17430 -42741 17498
rect 12849 17543 27413 17606
rect 12849 17495 27246 17543
rect 5831 17485 27246 17495
rect -43913 17371 -43883 17430
rect -43776 17408 -42741 17430
rect 5719 17462 27246 17485
rect -43776 17371 -43747 17408
rect -46187 17307 -44539 17325
rect -46187 17229 -44933 17307
rect -44868 17305 -44539 17307
rect -44868 17229 -44796 17305
rect -46187 17227 -44796 17229
rect -44731 17227 -44650 17305
rect -44585 17227 -44539 17305
rect -46187 17217 -44539 17227
rect -43913 17307 -43747 17371
rect -43913 17248 -43886 17307
rect -43779 17248 -43747 17307
rect -65699 17034 -60594 17052
rect -65699 17029 -65523 17034
rect -65699 16946 -65684 17029
rect -65623 16951 -65523 17029
rect -65462 17029 -60594 17034
rect -65462 16951 -65391 17029
rect -65623 16946 -65391 16951
rect -65330 16946 -60594 17029
rect -65699 16936 -60594 16946
rect -56304 17035 -50854 17054
rect -56304 17034 -55138 17035
rect -56304 16945 -55282 17034
rect -55223 16946 -55138 17034
rect -55079 17034 -50854 17035
rect -55079 16946 -54982 17034
rect -55223 16945 -54982 16946
rect -54923 17027 -50854 17034
rect -54923 16945 -50641 17027
rect -56304 16934 -50641 16945
rect -50974 16907 -50641 16934
rect -44650 17017 -44542 17217
rect -43913 17186 -43747 17248
rect 5719 17386 5770 17462
rect 5852 17425 27246 17462
rect 27364 17425 27413 17543
rect 5852 17402 27413 17425
rect 5852 17386 13053 17402
rect 5719 17296 13053 17386
rect 5719 17220 5773 17296
rect 5855 17291 13053 17296
rect 5855 17220 5911 17291
rect -25592 17163 -22995 17175
rect -25592 17158 -23091 17163
rect -25592 17074 -23382 17158
rect -23325 17156 -23091 17158
rect -23325 17074 -23236 17156
rect -25592 17072 -23236 17074
rect -23179 17079 -23091 17156
rect -23034 17079 -22995 17163
rect -23179 17072 -22995 17079
rect -25592 17059 -22995 17072
rect 5719 17128 5911 17220
rect 5719 17052 5779 17128
rect 5861 17052 5911 17128
rect -7147 17019 -1139 17041
rect -44650 16909 -40198 17017
rect -7147 17016 -6987 17019
rect -35948 16970 -30051 16990
rect -35948 16969 -34391 16970
rect -50974 16859 -50854 16907
rect -35948 16892 -34687 16969
rect -34625 16968 -34391 16969
rect -34625 16892 -34540 16968
rect -35948 16891 -34540 16892
rect -34478 16893 -34391 16968
rect -34329 16893 -30051 16970
rect -7147 16935 -7137 17016
rect -7066 16938 -6987 17016
rect -6916 17014 -1139 17019
rect -6916 16938 -6831 17014
rect -7066 16935 -6831 16938
rect -7147 16933 -6831 16935
rect -6760 16933 -1139 17014
rect -7147 16918 -1139 16933
rect 3243 17012 5238 17039
rect 5719 17033 5911 17052
rect 3243 17011 5081 17012
rect 3243 16940 4841 17011
rect 4898 16940 4961 17011
rect 5018 16941 5081 17011
rect 5138 16941 5238 17012
rect 25901 16974 31441 16978
rect 24945 16954 31441 16974
rect 24945 16951 26319 16954
rect 24945 16946 26180 16951
rect 5018 16940 5238 16941
rect 3243 16924 5238 16940
rect -34478 16891 -30051 16893
rect -35948 16876 -30051 16891
rect 5123 16870 5238 16924
rect 13876 16920 20479 16941
rect 5123 16755 9437 16870
rect 13876 16842 15334 16920
rect 15388 16917 20479 16920
rect 15388 16842 15475 16917
rect 13876 16839 15475 16842
rect 15529 16916 20479 16917
rect 15529 16839 15626 16916
rect 13876 16838 15626 16839
rect 15680 16838 20479 16916
rect 24945 16873 26025 16946
rect 26082 16878 26180 16946
rect 26237 16881 26319 16951
rect 26376 16881 31441 16954
rect 26237 16878 31441 16881
rect 26082 16873 31441 16878
rect 24945 16858 31441 16873
rect 25901 16855 31441 16858
rect 13876 16827 20479 16838
rect 9358 16712 9426 16755
rect -10849 16413 -10795 16521
rect -55937 16379 -53631 16413
rect -55937 16288 -55926 16379
rect -55850 16378 -55633 16379
rect -55850 16288 -55784 16378
rect -55937 16287 -55784 16288
rect -55708 16288 -55633 16378
rect -55557 16288 -53631 16379
rect -55708 16287 -53631 16288
rect -55937 16263 -53631 16287
rect -35385 16206 -32895 16259
rect -35385 16201 -35081 16206
rect -35385 16200 -35217 16201
rect -35385 16144 -35367 16200
rect -35314 16145 -35217 16200
rect -35164 16150 -35081 16201
rect -35028 16150 -32895 16206
rect -35164 16145 -32895 16150
rect -35314 16144 -32895 16145
rect -66381 16081 -63861 16136
rect -35385 16109 -32895 16144
rect -66381 16078 -66231 16081
rect -66381 16015 -66363 16078
rect -66303 16018 -66231 16078
rect -66171 16078 -63861 16081
rect -66171 16018 -66097 16078
rect -66303 16015 -66097 16018
rect -66037 16015 -63861 16078
rect -66381 15986 -63861 16015
rect -45779 16037 -43499 16075
rect -66282 14625 -66134 15986
rect -53179 15933 -53092 15954
rect -53179 15877 -53166 15933
rect -53110 15877 -53092 15933
rect -45779 15951 -45752 16037
rect -45682 16036 -43499 16037
rect -45682 15951 -45608 16036
rect -45779 15950 -45608 15951
rect -45538 15950 -45479 16036
rect -45409 15950 -43499 16036
rect -9151 16017 -9065 16304
rect -7913 16078 -4255 16123
rect -7913 16077 -7622 16078
rect -7913 16014 -7892 16077
rect -7830 16014 -7758 16077
rect -7696 16015 -7622 16077
rect -7560 16015 -4255 16078
rect -7696 16014 -4255 16015
rect -45779 15925 -43499 15950
rect -20784 15942 -20361 15975
rect -7913 15973 -4255 16014
rect 4061 15982 6345 16026
rect 4061 15980 4372 15982
rect -20784 15941 -20524 15942
rect -53179 15822 -53092 15877
rect -53179 15766 -53170 15822
rect -53114 15766 -53092 15822
rect -20784 15816 -20770 15941
rect -20644 15816 -20524 15941
rect -20784 15815 -20524 15816
rect -20397 15815 -20361 15942
rect 4061 15914 4083 15980
rect 4144 15979 4372 15980
rect 4144 15914 4230 15979
rect 4061 15913 4230 15914
rect 4291 15916 4372 15979
rect 4433 15916 6345 15982
rect 4291 15913 6345 15916
rect 4061 15876 6345 15913
rect 14619 15993 17573 16058
rect 14619 15990 14896 15993
rect 14619 15934 14661 15990
rect 14713 15934 14775 15990
rect 14827 15937 14896 15990
rect 14948 15937 17573 15993
rect 14827 15934 17573 15937
rect 14619 15908 17573 15934
rect 25328 15988 28287 16052
rect 25328 15985 25480 15988
rect 25328 15922 25348 15985
rect 25408 15925 25480 15985
rect 25540 15985 28287 15988
rect 25540 15925 25614 15985
rect 25408 15922 25614 15925
rect 25674 15922 28287 15985
rect 25328 15902 28287 15922
rect -20784 15794 -20361 15815
rect -53179 15751 -53092 15766
rect -32606 15760 -32519 15781
rect -63334 15703 -63247 15724
rect -63334 15647 -63321 15703
rect -63265 15647 -63247 15703
rect -63334 15592 -63247 15647
rect -32606 15704 -32593 15760
rect -32537 15704 -32519 15760
rect -32606 15649 -32519 15704
rect -63334 15536 -63325 15592
rect -63269 15536 -63247 15592
rect -63334 15521 -63247 15536
rect -42976 15622 -42889 15643
rect -42976 15566 -42963 15622
rect -42907 15566 -42889 15622
rect -32606 15593 -32597 15649
rect -32541 15593 -32519 15649
rect -32606 15578 -32519 15593
rect -3768 15668 -3681 15689
rect -3768 15612 -3755 15668
rect -3699 15612 -3681 15668
rect -42976 15511 -42889 15566
rect -42976 15455 -42967 15511
rect -42911 15455 -42889 15511
rect -3768 15557 -3681 15612
rect -3768 15501 -3759 15557
rect -3703 15501 -3681 15557
rect -3768 15486 -3681 15501
rect 6877 15582 6964 15603
rect 6877 15526 6890 15582
rect 6946 15526 6964 15582
rect -42976 15440 -42889 15455
rect 6877 15471 6964 15526
rect 6877 15415 6886 15471
rect 6942 15415 6964 15471
rect 6877 15400 6964 15415
rect 17940 15592 18027 15613
rect 17940 15536 17953 15592
rect 18009 15536 18027 15592
rect 17940 15481 18027 15536
rect 17940 15425 17949 15481
rect 18005 15425 18027 15481
rect 17940 15410 18027 15425
rect 28851 15585 28938 15606
rect 28851 15529 28864 15585
rect 28920 15529 28938 15585
rect 28851 15474 28938 15529
rect 28851 15418 28860 15474
rect 28916 15418 28938 15474
rect 28851 15403 28938 15418
rect -54114 14968 -54017 15035
rect -54114 14901 -54097 14968
rect -54033 14942 -54017 14968
rect -54033 14901 -53481 14942
rect -54114 14868 -53481 14901
rect -54114 14795 -54017 14868
rect -64624 14728 -64524 14763
rect -64624 14668 -64608 14728
rect -64544 14668 -64524 14728
rect -54114 14728 -54100 14795
rect -54036 14728 -54017 14795
rect -54114 14696 -54017 14728
rect -33946 14830 -33847 14863
rect -33946 14760 -33934 14830
rect -33866 14788 -33847 14830
rect -33866 14760 -32959 14788
rect -33946 14714 -32959 14760
rect -54097 14695 -54023 14696
rect -64624 14665 -64524 14668
rect -66847 14477 -65979 14625
rect -64624 14591 -63835 14665
rect -43882 14626 -43776 14677
rect -64624 14560 -64524 14591
rect -64624 14500 -64607 14560
rect -64543 14500 -64524 14560
rect -64624 14486 -64524 14500
rect -43882 14559 -43866 14626
rect -43794 14604 -43776 14626
rect -33946 14654 -33847 14714
rect -43794 14559 -43551 14604
rect -33946 14584 -33934 14654
rect -33866 14584 -33847 14654
rect -5670 14669 -5569 14742
rect -33946 14576 -33847 14584
rect -43882 14530 -43551 14559
rect -43882 14434 -43776 14530
rect -10834 14493 -10780 14607
rect -5670 14602 -5653 14669
rect -5582 14652 -5569 14669
rect -5582 14602 -4354 14652
rect -9723 14538 -9508 14584
rect -5670 14578 -4354 14602
rect 26028 14600 26409 14621
rect 26028 14597 26195 14600
rect 16988 14587 17071 14589
rect -5670 14493 -5569 14578
rect -43882 14367 -43869 14434
rect -43797 14367 -43776 14434
rect -5670 14426 -5658 14493
rect -5587 14426 -5569 14493
rect -5670 14411 -5569 14426
rect 5811 14555 5908 14585
rect 16988 14566 17591 14587
rect 26028 14581 26063 14597
rect 5811 14497 6332 14555
rect 5811 14431 5833 14497
rect 5892 14481 6332 14497
rect 16988 14511 17004 14566
rect 17059 14513 17591 14566
rect 26007 14534 26063 14581
rect 26123 14537 26195 14597
rect 26255 14597 26409 14600
rect 26255 14537 26329 14597
rect 26123 14534 26329 14537
rect 26389 14581 26409 14597
rect 26389 14534 28464 14581
rect 17059 14511 17071 14513
rect 5892 14431 5908 14481
rect -43882 14351 -43776 14367
rect -9523 14266 -9467 14399
rect 5811 14318 5908 14431
rect 16988 14424 17071 14511
rect 26007 14507 28464 14534
rect 16988 14369 17000 14424
rect 17055 14369 17071 14424
rect 16988 14358 17071 14369
rect 5811 14252 5826 14318
rect 5885 14252 5908 14318
rect 5811 14232 5908 14252
rect 5828 14231 5902 14232
rect 9033 14140 9431 14238
rect -24196 14096 -23787 14126
rect -24196 14094 -23950 14096
rect -53474 14035 -53387 14056
rect -53474 13979 -53461 14035
rect -53405 13979 -53387 14035
rect -24196 14008 -24175 14094
rect -24069 14010 -23950 14094
rect -23844 14010 -23787 14096
rect -24069 14008 -23787 14010
rect -24196 13984 -23787 14008
rect -53474 13924 -53387 13979
rect -53474 13868 -53465 13924
rect -53409 13868 -53387 13924
rect -53474 13853 -53387 13868
rect -32944 13852 -32857 13873
rect -32944 13796 -32931 13852
rect -32875 13796 -32857 13852
rect -63624 13763 -63537 13784
rect -68360 13716 -68233 13749
rect -68360 13646 -68333 13716
rect -68258 13646 -68233 13716
rect -68360 13622 -68233 13646
rect -66723 13709 -66590 13747
rect -66723 13646 -66686 13709
rect -66620 13646 -66590 13709
rect -66723 13614 -66590 13646
rect -63624 13707 -63611 13763
rect -63555 13707 -63537 13763
rect -63624 13652 -63537 13707
rect -32944 13741 -32857 13796
rect -63624 13596 -63615 13652
rect -63559 13596 -63537 13652
rect -63624 13581 -63537 13596
rect -55295 13631 -53639 13638
rect -55295 13540 -55278 13631
rect -55202 13629 -53639 13631
rect -55202 13540 -55146 13629
rect -55295 13538 -55146 13540
rect -55070 13538 -55006 13629
rect -54930 13538 -53639 13629
rect -46767 13594 -44667 13694
rect -32944 13685 -32935 13741
rect -32879 13685 -32857 13741
rect -55295 13521 -53639 13538
rect -55133 13417 -54985 13521
rect -65692 13338 -63830 13361
rect -65692 13335 -65540 13338
rect -65692 13272 -65672 13335
rect -65612 13275 -65540 13335
rect -65480 13335 -63830 13338
rect -65480 13275 -65406 13335
rect -65612 13272 -65406 13275
rect -65346 13272 -63830 13335
rect -56716 13317 -54985 13417
rect -65692 13244 -63830 13272
rect -65573 13117 -65425 13244
rect -72220 12969 -65293 13117
rect -72220 12907 -72072 12969
rect -72843 12790 -72071 12907
rect -72843 12787 -72176 12790
rect -72115 12726 -71891 12743
rect -72115 12722 -72089 12726
rect -72585 12676 -72089 12722
rect -72115 12672 -72089 12676
rect -72035 12672 -71966 12726
rect -71912 12672 -71891 12726
rect -72115 12654 -71891 12672
rect -72589 12584 -72405 12630
rect -72494 12565 -72405 12584
rect -72494 12476 -71259 12565
rect -72006 12357 -71735 12369
rect -72006 12356 -71464 12357
rect -72006 12268 -71988 12356
rect -71900 12268 -71829 12356
rect -71741 12268 -71464 12356
rect -72006 12267 -71464 12268
rect -72006 12244 -71735 12267
rect -71554 12224 -71464 12267
rect -71348 12314 -71259 12476
rect -71348 12263 -71333 12314
rect -71275 12263 -71259 12314
rect -71348 12251 -71259 12263
rect -73245 12149 -72621 12180
rect -71554 12176 -71539 12224
rect -71480 12176 -71464 12224
rect -71554 12173 -71464 12176
rect -71554 12162 -71465 12173
rect -73245 12147 -72885 12149
rect -73245 12012 -73140 12147
rect -72991 12014 -72885 12147
rect -72736 12014 -72621 12149
rect -72991 12012 -72621 12014
rect -73245 11991 -72621 12012
rect -71774 11948 -71605 12068
rect -71774 11335 -71588 11948
rect -71432 11947 -71382 12065
rect -71226 12048 -65978 12064
rect -71226 11976 -66370 12048
rect -66308 11976 -66255 12048
rect -66193 11976 -66141 12048
rect -66079 11976 -65978 12048
rect -71226 11963 -65978 11976
rect -71226 11948 -71103 11963
rect -71204 11885 -71103 11948
rect -71538 11733 -71370 11752
rect -71234 11750 -71091 11885
rect -71538 11633 -71510 11733
rect -71399 11633 -71370 11733
rect -71538 11619 -71370 11633
rect -71271 11735 -71091 11750
rect -71271 11635 -71253 11735
rect -71142 11733 -71091 11735
rect -71104 11719 -71091 11733
rect -65573 11743 -65425 12969
rect -64381 12450 -64304 12488
rect -64381 12389 -64372 12450
rect -64311 12411 -64304 12450
rect -64311 12389 -63804 12411
rect -64381 12334 -63804 12389
rect -61554 12371 -60577 12443
rect -64381 12315 -64304 12334
rect -64381 12254 -64373 12315
rect -64312 12254 -64304 12315
rect -64381 12243 -64304 12254
rect -55133 11743 -54985 13317
rect -44767 13300 -44667 13594
rect -43281 13664 -43194 13685
rect -32944 13670 -32857 13685
rect -4111 13741 -4024 13762
rect -4111 13685 -4098 13741
rect -4042 13685 -4024 13741
rect -43281 13608 -43268 13664
rect -43212 13608 -43194 13664
rect -43281 13553 -43194 13608
rect -4111 13630 -4024 13685
rect -4111 13574 -4102 13630
rect -4046 13574 -4024 13630
rect -4111 13559 -4024 13574
rect 6631 13730 6718 13751
rect 6631 13674 6644 13730
rect 6700 13674 6718 13730
rect 28527 13723 28614 13744
rect 6631 13619 6718 13674
rect 6631 13563 6640 13619
rect 6696 13563 6718 13619
rect -43281 13497 -43272 13553
rect -43216 13497 -43194 13553
rect 6631 13548 6718 13563
rect 17627 13700 17714 13721
rect 17627 13644 17640 13700
rect 17696 13644 17714 13700
rect 17627 13589 17714 13644
rect -43281 13482 -43194 13497
rect -25990 13531 -20740 13540
rect -25990 13526 -23242 13531
rect -34700 13448 -33032 13484
rect -34700 13447 -34400 13448
rect -34700 13409 -34685 13447
rect -34704 13394 -34685 13409
rect -34630 13446 -34400 13447
rect -34630 13394 -34546 13446
rect -34704 13393 -34546 13394
rect -34491 13395 -34400 13446
rect -34345 13395 -33032 13448
rect -25990 13448 -23387 13526
rect -23320 13453 -23242 13526
rect -23175 13529 -20740 13531
rect -23175 13453 -23103 13529
rect -23320 13451 -23103 13453
rect -23036 13451 -20740 13529
rect 17627 13533 17636 13589
rect 17692 13533 17714 13589
rect 28527 13667 28540 13723
rect 28596 13667 28614 13723
rect 28527 13612 28614 13667
rect 28527 13556 28536 13612
rect 28592 13556 28614 13612
rect 28527 13541 28614 13556
rect 17627 13518 17714 13533
rect -23320 13448 -20740 13451
rect -25990 13440 -20740 13448
rect -34491 13393 -33032 13395
rect -34704 13367 -33032 13393
rect -34704 13356 -34420 13367
rect -44941 13276 -43304 13300
rect -44941 13275 -44679 13276
rect -44941 13271 -44810 13275
rect -44941 13207 -44931 13271
rect -44876 13211 -44810 13271
rect -44755 13212 -44679 13275
rect -44624 13212 -43304 13276
rect -36360 13256 -34420 13356
rect -20840 13263 -20740 13440
rect -44755 13211 -43304 13212
rect -44876 13207 -43304 13211
rect -44941 13183 -43304 13207
rect -53899 12850 -53793 12863
rect -53899 12773 -53885 12850
rect -53808 12773 -53793 12850
rect -53899 12688 -53793 12773
rect -53899 12687 -53666 12688
rect -53899 12612 -53885 12687
rect -53810 12612 -53666 12687
rect -51472 12648 -50569 12720
rect -53899 12611 -53666 12612
rect -53899 12599 -53793 12611
rect -71271 11634 -71203 11635
rect -71104 11634 -71073 11719
rect -71271 11621 -71073 11634
rect -71216 11580 -71073 11621
rect -65573 11595 -54985 11743
rect -71216 11486 -71185 11580
rect -71100 11486 -71073 11580
rect -71216 11460 -71073 11486
rect -53880 11520 -53794 12599
rect -44761 12103 -44608 13183
rect -43386 12349 -43136 12366
rect -43386 12274 -43377 12349
rect -43302 12274 -43224 12349
rect -43149 12274 -43136 12349
rect -41234 12310 -40346 12382
rect -43386 12264 -43136 12274
rect -46493 11950 -44608 12103
rect -53266 11852 -53180 11861
rect -53266 11794 -53255 11852
rect -53197 11794 -53180 11852
rect -43053 11827 -42967 11867
rect -53266 11741 -53180 11794
rect -43058 11741 -42967 11827
rect -34574 11750 -34420 13256
rect -13450 12749 -13287 12837
rect -33735 12549 -33276 12575
rect -33735 12438 -33718 12549
rect -33607 12438 -33410 12549
rect -33299 12536 -33276 12549
rect -33299 12459 -32938 12536
rect -30962 12494 -30086 12566
rect -33299 12438 -33276 12459
rect -33735 12420 -33276 12438
rect -19376 11945 -19243 12032
rect -32533 11794 -20847 11838
rect -32533 11750 -23383 11794
rect -53266 11716 -42967 11741
rect -53266 11660 -53254 11716
rect -53198 11660 -42967 11716
rect -53266 11655 -42967 11660
rect -36287 11709 -23383 11750
rect -36287 11705 -34416 11709
rect -53255 11651 -53197 11655
rect -36287 11614 -34688 11705
rect -34621 11614 -34545 11705
rect -34478 11618 -34416 11705
rect -34349 11703 -23383 11709
rect -23316 11792 -20847 11794
rect -23316 11703 -23227 11792
rect -34349 11701 -23227 11703
rect -23160 11701 -23095 11792
rect -23028 11701 -20847 11792
rect -17390 11785 -17332 11903
rect -34349 11684 -20847 11701
rect -34349 11618 -32379 11684
rect -34478 11614 -32379 11618
rect -36287 11596 -32379 11614
rect -13992 11592 -13775 11689
rect -43488 11520 -43177 11535
rect -53880 11519 -43278 11520
rect -53880 11435 -43482 11519
rect -43398 11435 -43278 11519
rect -53880 11434 -43278 11435
rect -43192 11434 -43177 11520
rect -43488 11422 -43177 11434
rect -71933 11310 -71466 11335
rect -14403 11325 -14353 11453
rect -71933 11197 -71904 11310
rect -71787 11307 -71466 11310
rect -71787 11197 -71610 11307
rect -71933 11194 -71610 11197
rect -71493 11194 -71466 11307
rect -71933 11012 -71466 11194
rect -71933 10899 -71907 11012
rect -71790 10899 -71617 11012
rect -71500 10899 -71466 11012
rect -71933 10868 -71466 10899
rect -18209 10583 -18068 10629
rect -66380 10444 -62955 10472
rect -66380 10443 -66095 10444
rect -66380 10387 -66361 10443
rect -66308 10387 -66251 10443
rect -66198 10388 -66095 10443
rect -66042 10401 -62955 10444
rect -66042 10388 -62983 10401
rect -66198 10387 -62983 10388
rect -66380 10361 -62983 10387
rect -35397 10398 -33487 10434
rect -18907 10404 -18860 10509
rect -35397 10392 -35095 10398
rect -35397 10339 -35373 10392
rect -35318 10339 -35242 10392
rect -35187 10345 -35095 10392
rect -35040 10389 -33487 10398
rect -35040 10345 -33403 10389
rect -35187 10339 -33403 10345
rect -35397 10318 -33403 10339
rect -18058 10303 -18012 10399
rect -71457 10112 -62990 10138
rect -71457 10031 -62886 10112
rect -71457 10005 -62990 10031
rect -62314 9999 -33591 10108
rect -32849 9976 -24643 10055
rect -65697 9763 -65290 9801
rect -65697 9761 -65402 9763
rect -65710 9757 -65534 9761
rect -65710 9701 -65679 9757
rect -65626 9705 -65534 9757
rect -65481 9707 -65402 9761
rect -65349 9761 -65290 9763
rect -65349 9707 -62979 9761
rect -33558 9708 -33502 9734
rect -65481 9705 -62979 9707
rect -65626 9701 -62979 9705
rect -65710 9692 -62979 9701
rect -34703 9695 -33490 9708
rect -34703 9692 -34560 9695
rect -65697 9682 -65290 9692
rect -34703 9639 -34690 9692
rect -34635 9642 -34560 9692
rect -34505 9693 -33490 9695
rect -34505 9642 -34411 9693
rect -34635 9640 -34411 9642
rect -34356 9640 -33490 9693
rect -34635 9639 -33490 9640
rect -34703 9629 -33490 9639
rect -66387 9528 -62962 9564
rect -66387 9527 -66110 9528
rect -66387 9471 -66359 9527
rect -66306 9526 -66110 9527
rect -66306 9471 -66231 9526
rect -66387 9470 -66231 9471
rect -66178 9472 -66110 9526
rect -66057 9472 -62962 9528
rect -66178 9470 -62962 9472
rect -66387 9453 -62962 9470
rect -35405 9506 -33411 9550
rect -35405 9505 -35101 9506
rect -35405 9500 -35239 9505
rect -35405 9447 -35378 9500
rect -35323 9452 -35239 9500
rect -35184 9453 -35101 9505
rect -35046 9453 -33411 9506
rect -35184 9452 -33411 9453
rect -35323 9447 -33411 9452
rect -35405 9434 -33411 9447
rect -71446 9095 -63001 9220
rect -62327 9083 -33600 9196
rect -32873 9078 -25096 9153
rect -65702 8844 -65295 8876
rect -65702 8840 -65529 8844
rect -65702 8837 -65671 8840
rect -65706 8784 -65671 8837
rect -65618 8788 -65529 8840
rect -65476 8843 -65295 8844
rect -65476 8788 -65391 8843
rect -65618 8787 -65391 8788
rect -65338 8837 -65295 8843
rect -65338 8787 -62975 8837
rect -65618 8784 -62975 8787
rect -65706 8768 -62975 8784
rect -34709 8804 -33496 8815
rect -34709 8800 -34542 8804
rect -65702 8757 -65295 8768
rect -34709 8747 -34687 8800
rect -34632 8751 -34542 8800
rect -34487 8802 -33496 8804
rect -34487 8751 -34412 8802
rect -34632 8749 -34412 8751
rect -34357 8749 -33496 8802
rect -34632 8747 -33496 8749
rect -34709 8736 -33496 8747
rect -66387 8621 -62962 8648
rect -66387 8619 -66077 8621
rect -66387 8617 -66224 8619
rect -66387 8561 -66360 8617
rect -66307 8563 -66224 8617
rect -66171 8565 -66077 8619
rect -66024 8565 -62962 8621
rect -66171 8563 -62962 8565
rect -66307 8561 -62962 8563
rect -66387 8537 -62962 8561
rect -35405 8566 -33411 8599
rect -35405 8562 -35117 8566
rect -35405 8555 -35249 8562
rect -35405 8502 -35372 8555
rect -35317 8509 -35249 8555
rect -35194 8513 -35117 8562
rect -35062 8513 -33411 8566
rect -35194 8509 -33411 8513
rect -35317 8502 -33411 8509
rect -35405 8483 -33411 8502
rect -71417 8179 -62988 8308
rect -62302 8236 -33595 8275
rect -62302 8176 -33543 8236
rect -33739 8155 -33543 8176
rect -32855 8139 -25393 8215
rect -65698 7921 -65291 7950
rect -65698 7919 -65388 7921
rect -65698 7917 -65538 7919
rect -65706 7861 -65672 7917
rect -65619 7863 -65538 7917
rect -65485 7865 -65388 7919
rect -65335 7917 -65291 7921
rect -65335 7865 -62975 7917
rect -65485 7863 -62975 7865
rect -65619 7861 -62975 7863
rect -65706 7848 -62975 7861
rect -34704 7858 -33491 7873
rect -34704 7857 -34544 7858
rect -65698 7831 -65291 7848
rect -34704 7804 -34683 7857
rect -34628 7805 -34544 7857
rect -34489 7805 -34398 7858
rect -34343 7805 -33491 7858
rect -34628 7804 -33491 7805
rect -34704 7794 -33491 7804
rect -66391 7703 -62966 7739
rect -66391 7696 -66199 7703
rect -66391 7640 -66357 7696
rect -66304 7647 -66199 7696
rect -66146 7701 -62966 7703
rect -66146 7647 -66063 7701
rect -66304 7645 -66063 7647
rect -66010 7645 -62966 7701
rect -66304 7640 -62966 7645
rect -66391 7628 -62966 7640
rect -35392 7685 -33398 7721
rect -35392 7678 -35125 7685
rect -35392 7671 -35256 7678
rect -35392 7618 -35382 7671
rect -35327 7625 -35256 7671
rect -35201 7632 -35125 7678
rect -35070 7632 -33398 7685
rect -35201 7625 -33398 7632
rect -35327 7618 -33398 7625
rect -35392 7605 -33398 7618
rect -71398 7273 -62990 7399
rect -62335 7374 -61542 7495
rect -62335 7354 -33575 7374
rect -62328 7263 -33575 7354
rect -32869 7256 -25670 7337
rect -65701 7032 -65294 7061
rect -65701 7023 -65554 7032
rect -65717 7022 -65554 7023
rect -65717 6966 -65673 7022
rect -65620 6976 -65554 7022
rect -65501 6976 -65408 7032
rect -65355 7023 -65294 7032
rect -65355 6976 -62986 7023
rect -65620 6966 -62986 6976
rect -65717 6954 -62986 6966
rect -34704 6991 -33491 6999
rect -34704 6985 -34416 6991
rect -34704 6984 -34552 6985
rect -65701 6942 -65294 6954
rect -34704 6931 -34685 6984
rect -34630 6932 -34552 6984
rect -34497 6938 -34416 6985
rect -34361 6938 -33491 6991
rect -34497 6932 -33491 6938
rect -34630 6931 -33491 6932
rect -34704 6920 -33491 6931
rect -66391 6793 -62966 6826
rect -66391 6792 -66090 6793
rect -66391 6786 -66232 6792
rect -66391 6730 -66365 6786
rect -66312 6736 -66232 6786
rect -66179 6737 -66090 6792
rect -66037 6737 -62966 6793
rect -66179 6736 -62966 6737
rect -66312 6730 -62966 6736
rect -66391 6715 -62966 6730
rect -35405 6770 -33411 6804
rect -35405 6765 -35244 6770
rect -35405 6712 -35371 6765
rect -35316 6717 -35244 6765
rect -35189 6769 -33411 6770
rect -35189 6717 -35117 6769
rect -35316 6716 -35117 6717
rect -35062 6716 -33411 6769
rect -35316 6712 -33411 6716
rect -35405 6688 -33411 6712
rect -25756 6668 -25670 7256
rect -25465 6933 -25393 8139
rect -25177 7235 -25096 9078
rect -24724 7493 -24643 9976
rect -18282 9828 -17819 9832
rect -18282 9776 -18261 9828
rect -18209 9826 -17819 9828
rect -18209 9776 -18155 9826
rect -18282 9774 -18155 9776
rect -18095 9817 -17819 9826
rect -18095 9774 -17901 9817
rect -18282 9770 -17901 9774
rect -17829 9770 -17819 9817
rect -18282 9764 -17819 9770
rect -18150 9763 -17820 9764
rect -17901 9761 -17820 9763
rect -17901 9756 -17827 9761
rect -17123 9718 -17076 9821
rect -19275 9460 -19229 9560
rect -18327 9466 -18272 9561
rect -17790 9454 -17737 9557
rect -17458 9462 -17406 9594
rect -16920 9590 -16869 9685
rect -17129 9470 -17004 9527
rect -16595 9519 -16532 9614
rect -17129 9269 -17072 9470
rect -16921 9378 -16870 9477
rect -18158 9154 -18068 9203
rect -15850 9162 -15799 9251
rect -12896 9127 -12587 13377
rect -7145 13309 -4130 13348
rect -7145 13307 -6894 13309
rect -7145 13305 -7011 13307
rect -7145 13249 -7130 13305
rect -7077 13251 -7011 13305
rect -6958 13253 -6894 13307
rect -6841 13253 -4130 13309
rect 2647 13304 4841 13404
rect -6958 13251 -4130 13253
rect -7077 13249 -4130 13251
rect -7145 13231 -4130 13249
rect 4741 13299 4841 13304
rect 4741 13251 5201 13299
rect 13497 13283 15411 13307
rect -7020 12668 -6839 13231
rect 4741 13220 6430 13251
rect 4741 13215 4981 13220
rect 4741 13199 4848 13215
rect 4835 13151 4848 13199
rect 4910 13156 4981 13215
rect 5043 13156 5121 13220
rect 5183 13156 6430 13220
rect 13497 13245 17663 13283
rect 13497 13238 15595 13245
rect 13497 13236 15459 13238
rect 13497 13207 15341 13236
rect 15304 13180 15341 13207
rect 15393 13182 15459 13236
rect 15511 13189 15595 13238
rect 15647 13189 17663 13245
rect 24554 13277 26225 13331
rect 24554 13245 28405 13277
rect 24554 13242 26187 13245
rect 24554 13231 26055 13242
rect 15511 13182 17663 13189
rect 15393 13180 17663 13182
rect 15304 13166 17663 13180
rect 26010 13179 26055 13231
rect 26115 13182 26187 13242
rect 26247 13242 28405 13245
rect 26247 13182 26321 13242
rect 26115 13179 26321 13182
rect 26381 13179 28405 13242
rect 26010 13160 28405 13179
rect 4910 13151 6430 13156
rect 4835 13134 6430 13151
rect -8994 12487 -6839 12668
rect 6043 12849 6195 12876
rect 6043 12721 6064 12849
rect 6175 12832 6195 12849
rect 27804 12854 27909 12874
rect 27804 12849 28313 12854
rect 6175 12721 6364 12832
rect 27804 12783 27828 12849
rect 27894 12786 28313 12849
rect 27894 12783 27909 12786
rect 6043 12652 6195 12721
rect 6043 12543 6065 12652
rect 6174 12543 6195 12652
rect 27804 12694 27909 12783
rect 27804 12628 27828 12694
rect 27894 12628 27909 12694
rect 27804 12615 27909 12628
rect 6043 12527 6195 12543
rect -7020 11727 -6839 12487
rect -4385 12413 -4074 12463
rect -4385 12405 -4183 12413
rect -4385 12342 -4360 12405
rect -4303 12350 -4183 12405
rect -4126 12350 -4074 12413
rect -2052 12358 -1148 12430
rect -4303 12342 -4074 12350
rect -4385 12311 -4074 12342
rect 17355 12333 17605 12350
rect 6227 12302 6544 12317
rect 6227 12301 6426 12302
rect 6227 12199 6254 12301
rect 6356 12199 6426 12301
rect 6227 12198 6426 12199
rect 6530 12198 6544 12302
rect 8611 12261 9531 12333
rect 17355 12332 17522 12333
rect 17355 12257 17365 12332
rect 17441 12257 17522 12332
rect 17355 12256 17522 12257
rect 17599 12256 17605 12333
rect 19663 12293 20700 12365
rect 28107 12327 28204 12349
rect 28107 12326 28362 12327
rect 17355 12246 17605 12256
rect 28107 12251 28119 12326
rect 28194 12251 28362 12326
rect 30582 12287 31443 12359
rect 28107 12250 28362 12251
rect 6227 12184 6544 12198
rect 28107 12152 28204 12250
rect 28107 12075 28118 12152
rect 28195 12075 28204 12152
rect 28107 12067 28204 12075
rect -7147 11706 6201 11727
rect -7147 11700 -6988 11706
rect -7147 11601 -7136 11700
rect -7068 11607 -6988 11700
rect -6920 11698 6201 11706
rect -6920 11607 -6843 11698
rect -7068 11601 -6843 11607
rect -7147 11599 -6843 11601
rect -6775 11694 6201 11698
rect -6775 11693 4983 11694
rect -6775 11605 4843 11693
rect 4904 11606 4983 11693
rect 5044 11688 6201 11694
rect 5044 11606 5124 11688
rect 4904 11605 5124 11606
rect -6775 11600 5124 11605
rect 5185 11600 6201 11688
rect -6775 11599 6201 11600
rect -7147 11582 6201 11599
rect 6056 11568 6201 11582
rect 6056 11531 35638 11568
rect 6056 11530 15493 11531
rect 6056 11452 15340 11530
rect 15394 11453 15493 11530
rect 15547 11526 35638 11531
rect 15547 11522 26173 11526
rect 15547 11453 15626 11522
rect 15394 11452 15626 11453
rect 6056 11444 15626 11452
rect 15680 11521 26173 11522
rect 15680 11448 26033 11521
rect 26090 11453 26173 11521
rect 26230 11525 35638 11526
rect 26230 11453 26325 11525
rect 26090 11452 26325 11453
rect 26382 11452 35638 11525
rect 26090 11448 35638 11452
rect 15680 11444 35638 11448
rect 6056 11423 35638 11444
rect -9037 9233 -6738 9278
rect -9037 9230 -6832 9233
rect -9037 9226 -6984 9230
rect -9037 9144 -7125 9226
rect -7059 9148 -6984 9226
rect -6918 9151 -6832 9230
rect -6766 9151 -6738 9233
rect -6918 9148 -6738 9151
rect -7059 9144 -6738 9148
rect -15563 8810 -15200 8842
rect -12961 8810 -12023 9127
rect -9037 9103 -6738 9144
rect -23395 8799 -12023 8810
rect -23395 8792 -23225 8799
rect -23395 8718 -23371 8792
rect -23304 8725 -23225 8792
rect -23158 8725 -23080 8799
rect -23013 8759 -12023 8799
rect -23013 8725 -12047 8759
rect -23304 8718 -12047 8725
rect -23395 8658 -12047 8718
rect -23395 8650 -23077 8658
rect -23395 8646 -23220 8650
rect -23395 8572 -23370 8646
rect -23303 8576 -23220 8646
rect -23153 8584 -23077 8650
rect -23010 8584 -12047 8658
rect -23153 8576 -12047 8584
rect -23303 8572 -12047 8576
rect -23395 8545 -12047 8572
rect -23396 8498 -12047 8545
rect -23396 8494 -23116 8498
rect -23396 8400 -23367 8494
rect -23280 8404 -23116 8494
rect -23029 8404 -12047 8498
rect -23280 8400 -12047 8404
rect -23396 8354 -12047 8400
rect -23395 8329 -12047 8354
rect -15563 8248 -12047 8329
rect -15563 8173 -12042 8248
rect -15563 8169 -15200 8173
rect -15391 8161 -15200 8169
rect -24189 7832 -21414 7866
rect -24189 7738 -24167 7832
rect -24080 7738 -23917 7832
rect -23830 7738 -21414 7832
rect -24189 7728 -21414 7738
rect -15867 7632 -15782 7717
rect -24724 7412 -21326 7493
rect -16037 7425 -15866 7493
rect -25177 7154 -21769 7235
rect -25465 6861 -22064 6933
rect -25756 6582 -22332 6668
rect -71427 6357 -62999 6487
rect -62329 6343 -33583 6465
rect -32880 6333 -26130 6432
rect -26215 6297 -26130 6333
rect -26215 6212 -22598 6297
rect -65697 6093 -65290 6128
rect -65697 6091 -65403 6093
rect -65697 6089 -65539 6091
rect -65697 6088 -65664 6089
rect -65710 6033 -65664 6088
rect -65611 6035 -65539 6089
rect -65486 6037 -65403 6091
rect -65350 6088 -65290 6093
rect -65350 6037 -62979 6088
rect -65486 6035 -62979 6037
rect -65611 6033 -62979 6035
rect -65710 6019 -62979 6033
rect -34706 6075 -33493 6085
rect -34706 6073 -34403 6075
rect -34706 6070 -34545 6073
rect -65697 6009 -65290 6019
rect -34706 6017 -34686 6070
rect -34631 6020 -34545 6070
rect -34490 6022 -34403 6073
rect -34348 6022 -33493 6075
rect -34490 6020 -33493 6022
rect -34631 6017 -33493 6020
rect -34706 6006 -33493 6017
rect -66387 5868 -62962 5899
rect -66387 5812 -66355 5868
rect -66302 5866 -62962 5868
rect -66302 5865 -66084 5866
rect -66302 5812 -66221 5865
rect -66387 5809 -66221 5812
rect -66168 5810 -66084 5865
rect -66031 5810 -62962 5866
rect -66168 5809 -62962 5810
rect -66387 5788 -62962 5809
rect -35401 5858 -33407 5896
rect -35401 5852 -35243 5858
rect -35401 5799 -35369 5852
rect -35314 5805 -35243 5852
rect -35188 5856 -33407 5858
rect -35188 5805 -35103 5856
rect -35314 5803 -35103 5805
rect -35048 5803 -33407 5856
rect -35314 5799 -33407 5803
rect -35401 5780 -33407 5799
rect -24400 5877 -22866 5960
rect -71430 5425 -63003 5562
rect -62337 5413 -33583 5537
rect -24400 5526 -24300 5877
rect -32890 5426 -24300 5526
rect -65699 5178 -65292 5210
rect -65699 5175 -65537 5178
rect -65699 5171 -65678 5175
rect -65702 5119 -65678 5171
rect -65625 5122 -65537 5175
rect -65484 5122 -65390 5178
rect -65337 5171 -65292 5178
rect -62757 5171 -60759 5189
rect -65337 5122 -60759 5171
rect -65625 5119 -60759 5122
rect -65702 5102 -60759 5119
rect -65699 5091 -65292 5102
rect -62757 5083 -60759 5102
rect -34696 5160 -33483 5176
rect -34696 5159 -34400 5160
rect -34696 5158 -34551 5159
rect -34696 5105 -34679 5158
rect -34624 5106 -34551 5158
rect -34496 5107 -34400 5159
rect -34345 5107 -33483 5160
rect -34496 5106 -33483 5107
rect -34624 5105 -33483 5106
rect -34696 5097 -33483 5105
rect -60865 4619 -60759 5083
rect -56331 4728 -50596 4736
rect -56331 4720 -54966 4728
rect -56331 4715 -55124 4720
rect -56331 4641 -55285 4715
rect -55229 4646 -55124 4715
rect -55068 4654 -54966 4720
rect -54910 4654 -50596 4728
rect -55068 4646 -50596 4654
rect -55229 4641 -50596 4646
rect -56331 4628 -50596 4641
rect -50704 4354 -50596 4628
rect -46181 4379 -40176 4399
rect -46181 4377 -44798 4379
rect -46181 4302 -44929 4377
rect -44877 4304 -44798 4377
rect -44746 4374 -40176 4379
rect -44746 4304 -44652 4374
rect -44877 4302 -44652 4304
rect -46181 4299 -44652 4302
rect -44600 4299 -40176 4374
rect -46181 4287 -40176 4299
rect -40288 4097 -40176 4287
rect -35637 4167 -29944 4192
rect -35637 4165 -34392 4167
rect -35637 4077 -34680 4165
rect -34610 4161 -34392 4165
rect -34610 4077 -34544 4161
rect -35637 4073 -34544 4077
rect -34474 4079 -34392 4161
rect -34322 4079 -29944 4167
rect -22949 4188 -22866 5877
rect -22683 4391 -22598 6212
rect -22418 4909 -22332 6582
rect -22136 5756 -22064 6861
rect -21850 6625 -21769 7154
rect -15923 6775 -15826 6839
rect -21850 6544 -21378 6625
rect -16008 6564 -15856 6633
rect -14435 6063 -14387 6167
rect -22136 5684 -21370 5756
rect -16012 5709 -15860 5771
rect -12502 5352 -12042 8173
rect -22418 4823 -21424 4909
rect -16101 4842 -15999 4896
rect -12949 4773 -12880 4906
rect 14265 4522 21256 4564
rect 14265 4519 15584 4522
rect 14265 4463 15344 4519
rect 15396 4463 15472 4519
rect 15524 4466 15584 4519
rect 15636 4466 21256 4522
rect 15524 4463 21256 4466
rect -22683 4306 -21446 4391
rect 5040 4358 9629 4366
rect 3291 4338 9629 4358
rect 3291 4332 5142 4338
rect 3291 4328 4990 4332
rect 3291 4259 4842 4328
rect 4897 4263 4990 4328
rect 5045 4269 5142 4332
rect 5197 4269 9629 4338
rect 14265 4330 21256 4463
rect 25106 4421 34733 4453
rect 25106 4411 26319 4421
rect 25106 4406 26174 4411
rect 25106 4336 26031 4406
rect 26099 4341 26174 4406
rect 26242 4351 26319 4411
rect 26387 4351 34733 4421
rect 26242 4341 34733 4351
rect 26099 4336 34733 4341
rect 5045 4263 9629 4269
rect 4897 4259 9629 4263
rect 3291 4240 9629 4259
rect 5040 4232 9629 4240
rect 25106 4266 34733 4336
rect 25106 4263 26327 4266
rect 25106 4193 26032 4263
rect 26100 4193 26176 4263
rect 26244 4196 26327 4263
rect 26395 4196 34733 4266
rect 26244 4193 34733 4196
rect -22949 4105 -21334 4188
rect 25106 4178 34733 4193
rect -11797 4112 -1177 4132
rect -34474 4073 -29944 4079
rect -35637 3984 -29944 4073
rect -35637 3977 -34528 3984
rect -35637 3889 -34685 3977
rect -34615 3896 -34528 3977
rect -34458 3896 -34388 3984
rect -34318 3896 -29944 3984
rect -34615 3889 -29944 3896
rect -35637 3870 -29944 3889
rect -11991 4059 -1177 4112
rect -11991 3962 -7124 4059
rect -7056 3962 -6971 4059
rect -6903 3962 -6827 4059
rect -6759 3962 -1177 4059
rect -30003 3843 -29957 3870
rect -11991 3862 -1177 3962
rect -11991 3858 -6826 3862
rect -66381 3775 -63917 3824
rect -66381 3772 -66221 3775
rect -66381 3709 -66353 3772
rect -66293 3712 -66221 3772
rect -66161 3772 -63917 3775
rect -66161 3712 -66087 3772
rect -66293 3709 -66087 3712
rect -66027 3709 -63917 3772
rect -11991 3761 -7135 3858
rect -7067 3855 -6826 3858
rect -7067 3761 -6970 3855
rect -11991 3758 -6970 3761
rect -6902 3765 -6826 3855
rect -6758 3765 -1177 3862
rect -6902 3758 -1177 3765
rect -11991 3742 -1177 3758
rect -66381 3674 -63917 3709
rect -25320 3692 -22994 3737
rect -25320 3689 -23100 3692
rect -25320 3684 -23241 3689
rect -25320 3616 -23380 3684
rect -23325 3621 -23241 3684
rect -23186 3624 -23100 3689
rect -23045 3624 -22994 3692
rect -23186 3621 -22994 3624
rect -23325 3616 -22994 3621
rect -11530 3620 -11407 3742
rect -25320 3503 -22994 3616
rect 4063 3601 6527 3654
rect 4063 3599 4360 3601
rect 4063 3529 4084 3599
rect 4156 3529 4235 3599
rect 4307 3531 4360 3599
rect 4432 3531 6527 3601
rect 4307 3529 6527 3531
rect 4063 3504 6527 3529
rect -25320 3498 -23244 3503
rect -55936 3439 -53752 3485
rect -55936 3435 -55642 3439
rect -63342 3380 -63255 3401
rect -63342 3324 -63329 3380
rect -63273 3324 -63255 3380
rect -55936 3358 -55918 3435
rect -55853 3358 -55783 3435
rect -55718 3362 -55642 3435
rect -55577 3362 -53752 3439
rect -25320 3430 -23388 3498
rect -23333 3435 -23244 3498
rect -23189 3435 -23086 3503
rect -23031 3435 -22994 3503
rect 14619 3468 17394 3531
rect 14619 3463 14923 3468
rect 14619 3456 14798 3463
rect -23333 3430 -22994 3435
rect -25320 3418 -22994 3430
rect -55718 3358 -53752 3362
rect -55936 3335 -53752 3358
rect -7914 3394 -4155 3441
rect -7914 3392 -7610 3394
rect -7914 3390 -7746 3392
rect -63342 3269 -63255 3324
rect -63342 3213 -63333 3269
rect -63277 3213 -63255 3269
rect -35391 3288 -32901 3339
rect -7914 3317 -7895 3390
rect -7828 3319 -7746 3390
rect -7679 3321 -7610 3392
rect -7543 3321 -4155 3394
rect 14619 3400 14651 3456
rect 14703 3407 14798 3456
rect 14850 3412 14923 3463
rect 14975 3412 17394 3468
rect 14850 3407 17394 3412
rect 14703 3400 17394 3407
rect 14619 3381 17394 3400
rect -7679 3319 -4155 3321
rect -7828 3317 -4155 3319
rect -7914 3291 -4155 3317
rect -35391 3287 -35080 3288
rect -35391 3284 -35226 3287
rect -63342 3198 -63255 3213
rect -45766 3214 -43419 3257
rect -45766 3212 -45473 3214
rect -45766 3138 -45753 3212
rect -45681 3138 -45618 3212
rect -45546 3140 -45473 3212
rect -45401 3140 -43419 3214
rect -35391 3228 -35368 3284
rect -35314 3231 -35226 3284
rect -35172 3232 -35080 3287
rect -35026 3232 -32901 3288
rect -35172 3231 -32901 3232
rect -35314 3228 -32901 3231
rect -35391 3189 -32901 3228
rect 25328 3251 28081 3308
rect 25328 3248 25486 3251
rect -45546 3138 -43419 3140
rect -45766 3107 -43419 3138
rect 7103 3168 7190 3189
rect 7103 3112 7116 3168
rect 7172 3112 7190 3168
rect 25328 3185 25354 3248
rect 25414 3188 25486 3248
rect 25546 3248 28081 3251
rect 25546 3188 25620 3248
rect 25414 3185 25620 3188
rect 25680 3185 28081 3248
rect 25328 3158 28081 3185
rect -53207 3049 -53120 3070
rect -53207 2993 -53194 3049
rect -53138 2993 -53120 3049
rect 7103 3057 7190 3112
rect 7103 3001 7112 3057
rect 7168 3001 7190 3057
rect -53207 2938 -53120 2993
rect -53207 2882 -53198 2938
rect -53142 2882 -53120 2938
rect -53207 2867 -53120 2882
rect -3720 2975 -3633 2996
rect 7103 2986 7190 3001
rect 17949 3088 18036 3109
rect 17949 3032 17962 3088
rect 18018 3032 18036 3088
rect -3720 2919 -3707 2975
rect -3651 2919 -3633 2975
rect -3720 2864 -3633 2919
rect 17949 2977 18036 3032
rect 17949 2921 17958 2977
rect 18014 2921 18036 2977
rect 17949 2906 18036 2921
rect -42791 2816 -42704 2837
rect -42791 2760 -42778 2816
rect -42722 2760 -42704 2816
rect -42791 2705 -42704 2760
rect -42791 2649 -42782 2705
rect -42726 2649 -42704 2705
rect -42791 2634 -42704 2649
rect -32487 2818 -32400 2839
rect -32487 2762 -32474 2818
rect -32418 2762 -32400 2818
rect -3720 2808 -3711 2864
rect -3655 2808 -3633 2864
rect -32487 2707 -32400 2762
rect -32487 2651 -32478 2707
rect -32422 2651 -32400 2707
rect -32487 2636 -32400 2651
rect -24190 2746 -18866 2796
rect -3720 2793 -3633 2808
rect 28609 2863 28696 2884
rect 28609 2807 28622 2863
rect 28678 2807 28696 2863
rect -24190 2742 -23866 2746
rect -24190 2736 -24005 2742
rect -24190 2659 -24146 2736
rect -24088 2665 -24005 2736
rect -23947 2669 -23866 2742
rect -23808 2669 -18866 2746
rect 28609 2752 28696 2807
rect 28609 2696 28618 2752
rect 28674 2696 28696 2752
rect 28609 2681 28696 2696
rect -23947 2665 -18866 2669
rect -24088 2659 -18866 2665
rect -24190 2568 -18866 2659
rect -24190 2561 -24014 2568
rect -64616 2456 -64528 2513
rect -24190 2484 -24173 2561
rect -24115 2491 -24014 2561
rect -23956 2566 -18866 2568
rect -23956 2491 -23870 2566
rect -24115 2489 -23870 2491
rect -23812 2489 -18866 2566
rect -24115 2484 -18866 2489
rect -24190 2461 -18866 2484
rect -64616 2391 -64601 2456
rect -64545 2391 -64528 2456
rect -64616 2353 -64528 2391
rect -64616 2293 -63807 2353
rect -64616 2228 -64600 2293
rect -64544 2279 -63807 2293
rect 5813 2335 5910 2370
rect -64544 2228 -64528 2279
rect -64616 2216 -64528 2228
rect 5813 2266 5832 2335
rect 5896 2266 5910 2335
rect -54117 2167 -54017 2211
rect -54117 2098 -54104 2167
rect -54036 2098 -54017 2167
rect 5813 2183 5910 2266
rect 16987 2211 17070 2267
rect 5813 2169 6450 2183
rect -66853 2027 -65981 2057
rect -66853 2021 -66223 2027
rect -66853 1926 -66367 2021
rect -66301 1932 -66223 2021
rect -66157 1932 -66064 2027
rect -65998 1932 -65981 2027
rect -54117 2026 -54017 2098
rect -54117 1957 -54106 2026
rect -54038 2014 -54017 2026
rect -34093 2104 -33928 2116
rect -34093 2041 -33848 2104
rect -18289 2079 -18065 2149
rect -5672 2080 -5568 2121
rect 5813 2100 5831 2169
rect 5895 2109 6450 2169
rect 16987 2151 17002 2211
rect 17058 2151 17070 2211
rect 5895 2100 5910 2109
rect 5813 2086 5910 2100
rect -54038 1957 -53733 2014
rect -54117 1941 -53733 1957
rect -54110 1940 -53733 1941
rect -43883 1951 -43780 1988
rect -66301 1926 -65981 1932
rect -66853 1909 -65981 1926
rect -43883 1888 -43868 1951
rect -43800 1888 -43780 1951
rect -34093 1971 -33928 2041
rect -33868 1971 -33848 2041
rect -34093 1947 -33848 1971
rect -5672 2008 -5650 2080
rect -5581 2008 -5568 2080
rect -5672 1970 -5568 2008
rect 16987 2060 17070 2151
rect 16987 2036 17422 2060
rect 16987 1976 16999 2036
rect 17055 1986 17422 2036
rect 17055 1976 17070 1986
rect -43883 1786 -43780 1888
rect -35148 1878 -33841 1947
rect -35148 1808 -33928 1878
rect -33868 1868 -33841 1878
rect -5672 1907 -4153 1970
rect 16987 1956 17070 1976
rect -33868 1808 -33005 1868
rect -5672 1835 -5656 1907
rect -5587 1896 -4153 1907
rect -5587 1835 -5568 1896
rect 26027 1858 26409 1879
rect 26027 1855 26198 1858
rect 26027 1837 26066 1855
rect -5672 1818 -5568 1835
rect -35148 1794 -33005 1808
rect -43883 1723 -43869 1786
rect -43801 1723 -43387 1786
rect -43883 1712 -43387 1723
rect -35148 1782 -33841 1794
rect -43883 1704 -43780 1712
rect -63755 1410 -63668 1431
rect -63755 1354 -63742 1410
rect -63686 1354 -63668 1410
rect -63755 1299 -63668 1354
rect -63755 1243 -63746 1299
rect -63690 1243 -63668 1299
rect -63755 1228 -63668 1243
rect -68362 1157 -68225 1175
rect -68362 1064 -68328 1157
rect -68246 1064 -68225 1157
rect -68362 1038 -68225 1064
rect -66754 1148 -66624 1178
rect -66754 1083 -66723 1148
rect -66653 1083 -66624 1148
rect -66754 1052 -66624 1083
rect -65695 1025 -63792 1049
rect -65695 1022 -65530 1025
rect -65695 959 -65662 1022
rect -65602 962 -65530 1022
rect -65470 1022 -63792 1025
rect -65470 962 -65396 1022
rect -65602 959 -65396 962
rect -65336 959 -63792 1022
rect -56734 999 -55024 1099
rect -65695 932 -63792 959
rect -55124 710 -55024 999
rect -53640 1094 -53553 1115
rect -53640 1038 -53627 1094
rect -53571 1038 -53553 1094
rect -53640 983 -53553 1038
rect -53640 927 -53631 983
rect -53575 927 -53553 983
rect -53640 912 -53553 927
rect -43147 907 -43060 928
rect -43147 851 -43134 907
rect -43078 851 -43060 907
rect -43147 796 -43060 851
rect -55292 693 -53600 710
rect -55292 690 -54997 693
rect -55292 685 -55150 690
rect -55292 608 -55280 685
rect -55215 613 -55150 685
rect -55085 616 -54997 690
rect -54932 616 -53600 693
rect -46590 666 -44699 766
rect -43147 740 -43138 796
rect -43082 740 -43060 796
rect -43147 725 -43060 740
rect -55085 613 -53600 616
rect -55215 608 -53600 613
rect -55292 593 -53600 608
rect -67033 504 -65288 549
rect -67033 502 -65402 504
rect -67033 423 -65682 502
rect -65622 423 -65546 502
rect -65486 425 -65402 502
rect -65342 425 -65288 504
rect -44799 482 -44699 666
rect -65486 423 -65288 425
rect -67033 401 -65288 423
rect -44955 449 -43304 482
rect -44955 389 -44930 449
rect -44864 448 -44679 449
rect -44864 389 -44809 448
rect -44955 388 -44809 389
rect -44743 389 -44679 448
rect -44613 389 -43304 449
rect -44743 388 -43304 389
rect -44955 365 -43304 388
rect -64375 240 -64298 299
rect -64375 183 -64360 240
rect -64306 183 -64298 240
rect -64375 99 -64298 183
rect -64375 93 -63832 99
rect -64375 36 -64364 93
rect -64310 36 -63832 93
rect -61431 59 -60328 131
rect -64375 22 -63832 36
rect -54009 -239 -53698 -226
rect -54009 -241 -53826 -239
rect -54009 -316 -53994 -241
rect -53919 -316 -53826 -241
rect -53749 -240 -53698 -239
rect -53749 -316 -53634 -240
rect -51478 -280 -50660 -208
rect -54009 -317 -53634 -316
rect -54009 -322 -53698 -317
rect -53827 -325 -53748 -322
rect -43185 -468 -43106 -467
rect -43347 -469 -43270 -468
rect -43347 -544 -43346 -469
rect -43271 -544 -43270 -469
rect -43347 -545 -43270 -544
rect -43185 -545 -43184 -468
rect -43107 -545 -43106 -468
rect -41075 -508 -40210 -436
rect -43185 -546 -43106 -545
rect -65713 -684 -54875 -642
rect -65713 -688 -65385 -684
rect -65713 -695 -65518 -688
rect -65713 -808 -65671 -695
rect -65594 -801 -65518 -695
rect -65441 -797 -65385 -688
rect -65308 -693 -54875 -684
rect -65308 -770 -55282 -693
rect -55225 -770 -55151 -693
rect -55094 -694 -54875 -693
rect -55094 -770 -55022 -694
rect -65308 -771 -55022 -770
rect -54965 -771 -54875 -694
rect -65308 -797 -54875 -771
rect -65441 -801 -54875 -797
rect -65594 -808 -54875 -801
rect -65713 -831 -54875 -808
rect -46528 -875 -44538 -832
rect -46528 -877 -44631 -875
rect -46528 -879 -44782 -877
rect -46528 -969 -44917 -879
rect -44861 -967 -44782 -879
rect -44726 -965 -44631 -877
rect -44575 -965 -44538 -875
rect -44726 -967 -44538 -965
rect -44861 -969 -44538 -967
rect -46528 -1008 -44538 -969
rect -43497 -1017 -43397 -998
rect -43497 -1076 -43474 -1017
rect -43417 -1076 -43397 -1017
rect -43497 -1121 -43397 -1076
rect -54023 -1140 -43397 -1121
rect -54023 -1146 -43473 -1140
rect -54023 -1205 -54003 -1146
rect -53937 -1199 -43473 -1146
rect -43416 -1199 -43397 -1140
rect -53937 -1205 -43397 -1199
rect -54023 -1224 -43397 -1205
rect -43292 -1149 -43217 -1137
rect -43292 -1204 -43282 -1149
rect -43229 -1204 -43217 -1149
rect -43292 -1221 -43217 -1204
rect -54019 -1262 -53924 -1224
rect -54019 -1321 -54005 -1262
rect -53939 -1321 -53924 -1262
rect -43291 -1259 -43217 -1221
rect -43291 -1305 -43281 -1259
rect -54019 -1346 -53924 -1321
rect -53761 -1314 -43281 -1305
rect -43228 -1314 -43217 -1259
rect -53761 -1330 -43217 -1314
rect -53761 -1390 -53743 -1330
rect -53678 -1337 -43217 -1330
rect -53678 -1390 -43219 -1337
rect -53761 -1408 -43219 -1390
rect -53759 -1446 -53662 -1408
rect -53759 -1506 -53742 -1446
rect -53677 -1506 -53662 -1446
rect -53759 -1529 -53662 -1506
rect -35148 -2860 -34983 1782
rect -17385 1724 -17202 1807
rect 26018 1792 26066 1837
rect 26126 1795 26198 1855
rect 26258 1855 26409 1858
rect 26258 1795 26332 1855
rect 26126 1792 26332 1795
rect 26392 1837 26409 1855
rect 26392 1792 28052 1837
rect 26018 1763 28052 1792
rect 6759 1266 6846 1287
rect 6759 1210 6772 1266
rect 6828 1210 6846 1266
rect 6759 1155 6846 1210
rect 6759 1099 6768 1155
rect 6824 1099 6846 1155
rect 6759 1084 6846 1099
rect 17564 1148 17651 1169
rect 17564 1092 17577 1148
rect 17633 1092 17651 1148
rect -4084 1040 -3997 1061
rect -32846 967 -32759 988
rect -32846 911 -32833 967
rect -32777 911 -32759 967
rect -32846 856 -32759 911
rect -4084 984 -4071 1040
rect -4015 984 -3997 1040
rect -4084 929 -3997 984
rect 17564 1037 17651 1092
rect 17564 981 17573 1037
rect 17629 981 17651 1037
rect 17564 966 17651 981
rect 28335 951 28422 972
rect -4084 873 -4075 929
rect -4019 873 -3997 929
rect -4084 858 -3997 873
rect -32846 800 -32837 856
rect -32781 800 -32759 856
rect -32846 785 -32759 800
rect 4835 844 6619 879
rect 4835 841 4977 844
rect 4835 799 4848 841
rect 4716 781 4848 799
rect 4910 784 4977 841
rect 5039 784 5110 844
rect 5172 784 6619 844
rect 13711 833 15676 933
rect 15300 830 15590 833
rect 15300 821 15350 830
rect 4910 781 6619 784
rect 4716 762 6619 781
rect 15302 774 15350 821
rect 15402 774 15478 830
rect 15530 777 15590 830
rect 15642 777 15676 833
rect 28335 895 28348 951
rect 28404 895 28422 951
rect 28335 840 28422 895
rect 15530 774 15676 777
rect 4716 722 5181 762
rect 15302 756 15676 774
rect 15302 731 17627 756
rect 2880 699 5181 722
rect 15304 722 17627 731
rect 15304 719 15591 722
rect -7144 638 -4097 666
rect -7144 636 -6980 638
rect -34695 531 -32979 564
rect -34695 528 -34398 531
rect -34695 527 -34529 528
rect -34695 474 -34686 527
rect -34632 475 -34529 527
rect -34475 478 -34398 528
rect -34344 478 -32979 531
rect -25882 520 -23111 620
rect -7144 568 -7126 636
rect -7065 570 -6980 636
rect -6919 570 -6841 638
rect -6780 570 -4097 638
rect 2880 622 4816 699
rect 15304 663 15351 719
rect 15403 663 15479 719
rect 15531 666 15591 719
rect 15643 666 17627 722
rect 24554 697 26311 797
rect 28335 784 28344 840
rect 28400 784 28422 840
rect 28335 769 28422 784
rect 15531 663 17627 666
rect 15304 639 17627 663
rect -7065 568 -4097 570
rect -7144 549 -4097 568
rect 26211 533 26311 697
rect -34475 475 -32979 478
rect -34632 474 -32979 475
rect -34695 447 -32979 474
rect -23211 -94 -23111 520
rect 26013 508 28213 533
rect 26013 505 26187 508
rect 26013 442 26055 505
rect 26115 445 26187 505
rect 26247 505 28213 508
rect 26247 445 26321 505
rect 26115 442 26321 445
rect 26381 442 28213 505
rect 26013 416 28213 442
rect 27808 111 27903 136
rect 27808 43 27820 111
rect 27888 110 27903 111
rect 27888 43 28072 110
rect 27808 42 28072 43
rect -18831 -94 -18533 -66
rect -23398 -123 -18533 -94
rect -23398 -125 -23092 -123
rect -23398 -193 -23386 -125
rect -23332 -126 -23092 -125
rect -23332 -193 -23235 -126
rect -23398 -194 -23235 -193
rect -23181 -191 -23092 -126
rect -23038 -138 -18533 -123
rect -23038 -191 -18813 -138
rect -23181 -194 -18813 -191
rect -23398 -204 -18813 -194
rect -18831 -223 -18813 -204
rect -18748 -223 -18638 -138
rect -18573 -223 -18533 -138
rect -18831 -255 -18533 -223
rect -4388 -240 -3891 -216
rect -33203 -361 -32800 -342
rect -33203 -470 -33186 -361
rect -33077 -470 -32936 -361
rect -33203 -472 -32936 -470
rect -32825 -472 -32800 -361
rect -30753 -426 -29917 -354
rect -4388 -378 -4368 -240
rect -4230 -241 -3891 -240
rect -4230 -377 -4045 -241
rect -3909 -377 -3891 -241
rect -2006 -324 -1031 -252
rect -4230 -378 -3891 -377
rect -4388 -392 -3891 -378
rect -33203 -493 -32800 -472
rect -7148 -1078 5240 -1023
rect -7148 -1083 5158 -1078
rect -7148 -1084 4997 -1083
rect -34722 -1127 -22932 -1110
rect -34722 -1132 -23103 -1127
rect -34722 -1134 -23254 -1132
rect -34722 -1171 -23389 -1134
rect -34722 -1181 -34391 -1171
rect -34722 -1281 -34687 -1181
rect -34614 -1183 -34391 -1181
rect -34614 -1281 -34536 -1183
rect -34722 -1283 -34536 -1281
rect -34463 -1271 -34391 -1183
rect -34318 -1202 -23389 -1171
rect -23334 -1200 -23254 -1134
rect -23199 -1195 -23103 -1132
rect -23048 -1195 -22932 -1127
rect -7148 -1153 4847 -1084
rect 4902 -1152 4997 -1084
rect 5052 -1147 5158 -1083
rect 5213 -1147 5240 -1078
rect 5052 -1152 5240 -1147
rect 4902 -1153 5240 -1152
rect -7148 -1182 5240 -1153
rect -7148 -1194 -6733 -1182
rect -23199 -1200 -22932 -1195
rect -23334 -1202 -22932 -1200
rect -34318 -1271 -22932 -1202
rect -34463 -1272 -23104 -1271
rect -34463 -1274 -23251 -1272
rect -34463 -1283 -23392 -1274
rect -34722 -1342 -23392 -1283
rect -23337 -1340 -23251 -1274
rect -23196 -1339 -23104 -1272
rect -23049 -1339 -22932 -1271
rect -11539 -1212 -6733 -1194
rect -11539 -1214 -6989 -1212
rect -11539 -1293 -7133 -1214
rect -7071 -1291 -6989 -1214
rect -6927 -1213 -6733 -1212
rect -6927 -1291 -6857 -1213
rect -7071 -1292 -6857 -1291
rect -6795 -1283 -6733 -1213
rect 6670 -1218 6800 -77
rect 8820 -111 9629 -39
rect 27808 -75 27903 42
rect 27808 -141 27821 -75
rect 27887 -141 27903 -75
rect 16681 -194 16793 -182
rect 16681 -195 17557 -194
rect 16681 -270 16703 -195
rect 16778 -270 17557 -195
rect 19630 -234 20455 -162
rect 27808 -164 27903 -141
rect 16681 -271 17557 -270
rect 16681 -409 16793 -271
rect 16681 -486 16702 -409
rect 16779 -486 16793 -409
rect 16681 -499 16793 -486
rect 28107 -418 28206 -399
rect 28107 -493 28121 -418
rect 28197 -493 28206 -418
rect 30343 -457 31144 -385
rect 6967 -536 7097 -533
rect 6920 -663 7097 -536
rect 28107 -563 28206 -493
rect 13767 -656 15721 -628
rect 13767 -658 15606 -656
rect 6920 -923 7050 -663
rect 13767 -733 15332 -658
rect 15395 -662 15606 -658
rect 15395 -733 15474 -662
rect 13767 -737 15474 -733
rect 15537 -731 15606 -662
rect 15669 -731 15721 -656
rect 28107 -640 28118 -563
rect 28195 -640 28206 -563
rect 28107 -659 28206 -640
rect 15537 -737 15721 -731
rect 13767 -752 15721 -737
rect 17006 -688 17108 -671
rect 17006 -765 17013 -688
rect 17091 -694 17108 -688
rect 17091 -758 17928 -694
rect 17091 -765 17108 -758
rect 17006 -852 17108 -765
rect 17006 -923 17018 -852
rect 6920 -929 17018 -923
rect 17096 -923 17108 -852
rect 24604 -780 26427 -750
rect 24604 -793 26454 -780
rect 24604 -795 26319 -793
rect 24604 -799 26183 -795
rect 24604 -898 26033 -799
rect 26100 -894 26183 -799
rect 26250 -892 26319 -795
rect 26386 -892 26454 -793
rect 26250 -894 26454 -892
rect 26100 -898 26454 -894
rect 24604 -914 26454 -898
rect 17096 -929 17109 -923
rect 6920 -1053 17109 -929
rect 26282 -1091 26454 -914
rect 6650 -1246 16796 -1218
rect -6795 -1292 -6744 -1283
rect -7071 -1293 -6744 -1292
rect -11539 -1319 -6744 -1293
rect -23196 -1340 -22932 -1339
rect -23337 -1342 -22932 -1340
rect -34722 -1351 -22932 -1342
rect 6650 -1323 16700 -1246
rect 16778 -1323 16796 -1246
rect 26282 -1263 35418 -1091
rect 6650 -1348 16796 -1323
rect 16693 -1410 16795 -1348
rect -18720 -1530 -18500 -1410
rect 16693 -1487 16705 -1410
rect 16783 -1487 16795 -1410
rect 16693 -1509 16795 -1487
rect -18750 -1770 -18530 -1650
rect -43765 -2861 -34983 -2860
rect -43801 -2965 -34983 -2861
rect -43801 -3122 -43764 -2965
rect -43673 -3025 -34983 -2965
rect -43673 -3122 -43647 -3025
rect -54371 -3259 -54203 -3198
rect -54371 -3396 -54337 -3259
rect -54234 -3396 -54203 -3259
rect -54371 -3511 -54203 -3396
rect -43801 -3245 -43647 -3122
rect -43801 -3402 -43772 -3245
rect -43681 -3402 -43647 -3245
rect -43801 -3431 -43647 -3402
rect -64581 -3528 -54346 -3511
rect -64606 -3648 -54346 -3528
rect -54243 -3648 -54203 -3511
rect -64606 -3659 -54203 -3648
rect -64606 -3793 -64576 -3659
rect -64498 -3679 -54203 -3659
rect -64498 -3793 -64482 -3679
rect -64606 -3861 -64482 -3793
rect -64606 -3995 -64578 -3861
rect -64500 -3995 -64482 -3861
rect -64606 -4025 -64482 -3995
rect -19364 -3937 -3483 -3892
rect -19364 -3940 -3584 -3937
rect -19364 -3993 -3711 -3940
rect -3659 -3990 -3584 -3940
rect -3532 -3990 -3483 -3937
rect -3659 -3993 -3483 -3990
rect -19364 -4020 -3483 -3993
rect -19364 -4110 -19319 -4020
rect -19229 -4042 -3483 -4020
rect -19229 -4110 -19200 -4042
rect -33055 -4142 -32542 -4116
rect -19364 -4142 -19200 -4110
rect -33055 -4292 -33023 -4142
rect -32873 -4143 -19200 -4142
rect -32873 -4291 -32705 -4143
rect -32557 -4179 -19200 -4143
rect -32557 -4186 -21740 -4179
rect -32557 -4262 -21964 -4186
rect -21877 -4255 -21740 -4186
rect -21653 -4184 -19200 -4179
rect -21653 -4255 -19319 -4184
rect -21877 -4262 -19319 -4255
rect -32557 -4274 -19319 -4262
rect -19229 -4274 -19200 -4184
rect -32557 -4291 -19200 -4274
rect -32873 -4292 -19200 -4291
rect -33055 -4311 -32542 -4292
rect -18841 -4334 -3761 -4184
rect -54018 -4403 -53920 -4390
rect -54018 -4404 -53469 -4403
rect -54018 -4476 -54002 -4404
rect -53930 -4476 -53469 -4404
rect -54018 -4477 -53469 -4476
rect -18841 -4422 -18823 -4334
rect -18735 -4422 -18691 -4334
rect -54018 -4553 -53920 -4477
rect -18841 -4515 -18691 -4422
rect -18841 -4541 -18823 -4515
rect -54018 -4627 -54003 -4553
rect -53929 -4627 -53920 -4553
rect -54018 -4641 -53920 -4627
rect -33401 -4574 -18823 -4541
rect -33401 -4579 -22080 -4574
rect -33401 -4655 -22308 -4579
rect -22221 -4650 -22080 -4579
rect -21993 -4603 -18823 -4574
rect -18735 -4603 -18691 -4515
rect -21993 -4650 -18691 -4603
rect -22221 -4655 -18691 -4650
rect -33401 -4691 -18691 -4655
rect -3911 -4549 -3761 -4334
rect 16684 -4364 16787 -4353
rect 16684 -4365 17722 -4364
rect 16684 -4437 16703 -4365
rect 16775 -4437 17722 -4365
rect 16684 -4438 17722 -4437
rect 28098 -4423 28444 -4397
rect 16684 -4528 16787 -4438
rect 28098 -4488 28133 -4423
rect 28197 -4426 28444 -4423
rect 28197 -4488 28315 -4426
rect 28098 -4491 28315 -4488
rect 28379 -4491 28444 -4426
rect 28098 -4515 28444 -4491
rect -55069 -4759 -52866 -4727
rect -56184 -4777 -52866 -4759
rect -56184 -4781 -54975 -4777
rect -65695 -4824 -65313 -4816
rect -65695 -4829 -65400 -4824
rect -65695 -4832 -65551 -4829
rect -65695 -4833 -65684 -4832
rect -65698 -4911 -65684 -4833
rect -65618 -4908 -65551 -4832
rect -65485 -4903 -65400 -4829
rect -65334 -4833 -65313 -4824
rect -65334 -4903 -60835 -4833
rect -65485 -4908 -60835 -4903
rect -65618 -4911 -60835 -4908
rect -65698 -4968 -60835 -4911
rect -65698 -4969 -65393 -4968
rect -65698 -5048 -65686 -4969
rect -65620 -5048 -65541 -4969
rect -65475 -5047 -65393 -4969
rect -65327 -5047 -60835 -4968
rect -56184 -4852 -55281 -4781
rect -55224 -4783 -54975 -4781
rect -55224 -4852 -55137 -4783
rect -56184 -4854 -55137 -4852
rect -55080 -4848 -54975 -4783
rect -54918 -4848 -52866 -4777
rect -55080 -4854 -52866 -4848
rect -56184 -4868 -52866 -4854
rect -46284 -4754 -37053 -4704
rect -46284 -4851 -44927 -4754
rect -44863 -4851 -44778 -4754
rect -44714 -4851 -44630 -4754
rect -44566 -4851 -37053 -4754
rect -56184 -4940 -54889 -4868
rect -46284 -4879 -37053 -4851
rect -35812 -4915 -34453 -4789
rect -33401 -4905 -32220 -4691
rect -3911 -4699 -2734 -4549
rect 16684 -4602 16702 -4528
rect 16776 -4602 16787 -4528
rect 16684 -4615 16787 -4602
rect 26237 -4681 29080 -4669
rect 24890 -4746 29080 -4681
rect 24890 -4824 26022 -4746
rect 26093 -4747 29080 -4746
rect 26093 -4824 26177 -4747
rect 24890 -4825 26177 -4824
rect 26248 -4750 29080 -4747
rect 26248 -4825 26330 -4750
rect 24890 -4828 26330 -4825
rect 26401 -4774 29080 -4750
rect 26401 -4828 26415 -4774
rect 24890 -4843 26415 -4828
rect -56184 -4944 -54971 -4940
rect -56184 -5015 -55283 -4944
rect -55226 -4945 -54971 -4944
rect -55226 -5015 -55139 -4945
rect -56184 -5016 -55139 -5015
rect -55082 -5011 -54971 -4945
rect -54914 -5011 -54889 -4940
rect -55082 -5016 -54889 -5011
rect -56184 -5027 -54889 -5016
rect -65475 -5048 -60835 -5047
rect -65698 -5059 -60835 -5048
rect -34579 -5099 -34453 -4915
rect -16940 -5068 -16786 -4916
rect -12195 -4924 -3611 -4891
rect -12195 -4925 -6992 -4924
rect -12195 -4980 -7128 -4925
rect -7073 -4979 -6992 -4925
rect -6937 -4925 -3611 -4924
rect -6937 -4979 -6838 -4925
rect -7073 -4980 -6838 -4979
rect -6783 -4980 -3611 -4925
rect -12195 -5004 -3611 -4980
rect 3435 -4899 13056 -4863
rect 3435 -5001 4843 -4899
rect 4922 -4900 5139 -4899
rect 4922 -5001 4993 -4900
rect 3435 -5002 4993 -5001
rect 5072 -5001 5139 -4900
rect 5218 -5001 13056 -4899
rect 27801 -4956 27912 -4888
rect 5072 -5002 13056 -5001
rect 3435 -5022 13056 -5002
rect 14228 -5009 15736 -4994
rect 14228 -5013 15462 -5009
rect 9636 -5068 13039 -5022
rect -53775 -5127 -53304 -5104
rect -53775 -5128 -53571 -5127
rect -53775 -5186 -53741 -5128
rect -53685 -5185 -53571 -5128
rect -53515 -5185 -53304 -5127
rect -53685 -5186 -53304 -5185
rect -53775 -5215 -53304 -5186
rect -34699 -5123 -33217 -5099
rect -34699 -5126 -34531 -5123
rect -34699 -5193 -34685 -5126
rect -34621 -5190 -34531 -5126
rect -34467 -5125 -33217 -5123
rect -34467 -5190 -34397 -5125
rect -34621 -5192 -34397 -5190
rect -34333 -5192 -33217 -5125
rect -34621 -5193 -33217 -5192
rect -34699 -5212 -33217 -5193
rect -26093 -5119 -16786 -5068
rect -26093 -5192 -23384 -5119
rect -23313 -5124 -16786 -5119
rect -23313 -5192 -23227 -5124
rect -26093 -5197 -23227 -5192
rect -23156 -5128 -16786 -5124
rect -23156 -5197 -23074 -5128
rect -26093 -5201 -23074 -5197
rect -23003 -5201 -16786 -5128
rect 14228 -5084 15330 -5013
rect 15396 -5080 15462 -5013
rect 15528 -5012 15736 -5009
rect 15528 -5080 15623 -5012
rect 15396 -5083 15623 -5080
rect 15689 -5083 15736 -5012
rect 15396 -5084 15736 -5083
rect -26093 -5222 -16786 -5201
rect -3577 -5175 -3487 -5162
rect -3577 -5228 -3552 -5175
rect -3500 -5228 -3487 -5175
rect -3577 -5290 -3487 -5228
rect 14228 -5196 15736 -5084
rect 17183 -5076 17659 -5029
rect 17183 -5077 17541 -5076
rect 17183 -5135 17262 -5077
rect 17318 -5083 17541 -5077
rect 17318 -5135 17380 -5083
rect 17183 -5141 17380 -5135
rect 17436 -5134 17541 -5083
rect 17597 -5134 17659 -5076
rect 17436 -5141 17659 -5134
rect 17183 -5192 17659 -5141
rect 27801 -5031 27820 -4956
rect 27892 -5031 27912 -4956
rect 27801 -5120 27912 -5031
rect 27801 -5133 28390 -5120
rect 14228 -5198 15632 -5196
rect 14228 -5269 15328 -5198
rect 15394 -5200 15632 -5198
rect 15394 -5269 15478 -5200
rect 14228 -5271 15478 -5269
rect 15544 -5267 15632 -5200
rect 15698 -5267 15736 -5196
rect 27801 -5208 27815 -5133
rect 27887 -5208 28390 -5133
rect 27801 -5231 28390 -5208
rect 27810 -5240 27880 -5231
rect 15544 -5271 15736 -5267
rect 14228 -5282 15736 -5271
rect -3577 -5343 -3566 -5290
rect -3514 -5343 -3487 -5290
rect -33082 -5379 -32956 -5355
rect -3577 -5358 -3487 -5343
rect -33082 -5434 -33042 -5379
rect -32987 -5434 -32956 -5379
rect -33082 -5490 -32956 -5434
rect -33082 -5545 -33041 -5490
rect -32986 -5545 -32956 -5490
rect -33082 -5567 -32956 -5545
rect -66381 -5738 -63920 -5688
rect -66381 -5741 -66224 -5738
rect -66381 -5804 -66356 -5741
rect -66296 -5801 -66224 -5741
rect -66164 -5741 -63920 -5738
rect -66164 -5801 -66090 -5741
rect -66296 -5804 -66090 -5801
rect -66030 -5804 -63920 -5741
rect -66381 -5838 -63920 -5804
rect -45768 -5761 -43443 -5710
rect -45768 -5763 -45478 -5761
rect -45768 -5764 -45614 -5763
rect -45768 -5826 -45752 -5764
rect -45687 -5825 -45614 -5764
rect -45549 -5823 -45478 -5763
rect -45413 -5823 -43443 -5761
rect -45549 -5825 -43443 -5823
rect -45687 -5826 -43443 -5825
rect -45768 -5860 -43443 -5826
rect -24189 -5855 -19896 -5824
rect -24189 -5858 -23919 -5855
rect -24189 -5943 -24154 -5858
rect -24071 -5940 -23919 -5858
rect -23836 -5940 -19896 -5855
rect -24071 -5943 -19896 -5940
rect -24189 -5974 -19896 -5943
rect 4056 -5977 6539 -5933
rect 4056 -5979 4369 -5977
rect 4056 -6052 4082 -5979
rect 4161 -5980 4369 -5979
rect 4161 -6052 4231 -5980
rect 4056 -6053 4231 -6052
rect 4310 -6050 4369 -5980
rect 4448 -6050 6539 -5977
rect 4310 -6053 6539 -6050
rect 4056 -6083 6539 -6053
rect -63351 -6122 -63264 -6101
rect -63351 -6178 -63338 -6122
rect -63282 -6178 -63264 -6122
rect -63351 -6233 -63264 -6178
rect -63351 -6289 -63342 -6233
rect -63286 -6289 -63264 -6233
rect -63351 -6304 -63264 -6289
rect -42812 -6147 -42725 -6126
rect -42812 -6203 -42799 -6147
rect -42743 -6203 -42725 -6147
rect -42812 -6258 -42725 -6203
rect -42812 -6314 -42803 -6258
rect -42747 -6314 -42725 -6258
rect -42812 -6329 -42725 -6314
rect -19347 -6183 -19260 -6162
rect -19347 -6239 -19334 -6183
rect -19278 -6239 -19260 -6183
rect -19347 -6294 -19260 -6239
rect -19347 -6350 -19338 -6294
rect -19282 -6350 -19260 -6294
rect -19347 -6365 -19260 -6350
rect 7086 -6370 7173 -6349
rect 7086 -6426 7099 -6370
rect 7155 -6426 7173 -6370
rect 7086 -6481 7173 -6426
rect 7086 -6537 7095 -6481
rect 7151 -6537 7173 -6481
rect -32038 -6653 -31992 -6554
rect -2552 -6631 -2506 -6548
rect 7086 -6552 7173 -6537
rect -66699 -7084 -65981 -7054
rect -66699 -7088 -66070 -7084
rect -66699 -7093 -66225 -7088
rect -66699 -7181 -66367 -7093
rect -66302 -7176 -66225 -7093
rect -66160 -7172 -66070 -7088
rect -66005 -7172 -65981 -7084
rect -66160 -7176 -65981 -7172
rect -66302 -7181 -65981 -7176
rect -66699 -7196 -65981 -7181
rect -64587 -7141 -64502 -7091
rect -64587 -7205 -64572 -7141
rect -64513 -7159 -64502 -7141
rect -43769 -7123 -43663 -7105
rect -64513 -7205 -63960 -7159
rect -64587 -7233 -63960 -7205
rect -43769 -7205 -43750 -7123
rect -43682 -7181 -43663 -7123
rect -20587 -7178 -20448 -7167
rect -43682 -7205 -43115 -7181
rect -64587 -7309 -64502 -7233
rect -43769 -7255 -43115 -7205
rect -20587 -7249 -20561 -7178
rect -20476 -7249 -20448 -7178
rect -64587 -7373 -64575 -7309
rect -64516 -7373 -64502 -7309
rect -55935 -7272 -53567 -7262
rect -55935 -7273 -55668 -7272
rect -55935 -7277 -55794 -7273
rect -55935 -7329 -55922 -7277
rect -55865 -7325 -55794 -7277
rect -55737 -7324 -55668 -7273
rect -55611 -7324 -53567 -7272
rect -55737 -7325 -53567 -7324
rect -55865 -7329 -53567 -7325
rect -55935 -7344 -53567 -7329
rect -43769 -7315 -43663 -7255
rect -64587 -7389 -64502 -7373
rect -43769 -7397 -43750 -7315
rect -43682 -7397 -43663 -7315
rect -43769 -7415 -43663 -7397
rect -20587 -7295 -20448 -7249
rect 14606 -7236 17587 -7223
rect 14606 -7237 14900 -7236
rect 14606 -7238 14766 -7237
rect 14606 -7294 14647 -7238
rect 14699 -7293 14766 -7238
rect 14818 -7292 14900 -7237
rect 14952 -7292 17587 -7236
rect 25346 -7278 25705 -7275
rect 14818 -7293 17587 -7292
rect 14699 -7294 17587 -7293
rect -20587 -7319 -19884 -7295
rect 14606 -7305 17587 -7294
rect 25325 -7280 28228 -7278
rect 25325 -7283 25486 -7280
rect -20587 -7390 -20563 -7319
rect -20478 -7369 -19884 -7319
rect -7911 -7344 -3818 -7337
rect -20478 -7390 -20448 -7369
rect -20587 -7458 -20448 -7390
rect -7911 -7410 -7898 -7344
rect -7838 -7345 -3818 -7344
rect -7838 -7410 -7743 -7345
rect -7911 -7411 -7743 -7410
rect -7683 -7411 -7610 -7345
rect -7550 -7411 -3818 -7345
rect 25325 -7346 25354 -7283
rect 25414 -7343 25486 -7283
rect 25546 -7283 28228 -7280
rect 25546 -7343 25620 -7283
rect 25414 -7346 25620 -7343
rect 25680 -7346 28228 -7283
rect 4854 -7379 5199 -7356
rect 25325 -7360 28228 -7346
rect 4854 -7383 5123 -7379
rect 4854 -7384 4996 -7383
rect 4854 -7404 4869 -7384
rect -7911 -7419 -3818 -7411
rect -20587 -7529 -20568 -7458
rect -20483 -7529 -20448 -7458
rect 4825 -7438 4869 -7404
rect 4926 -7437 4996 -7384
rect 5053 -7433 5123 -7383
rect 5180 -7404 5199 -7379
rect 5180 -7433 6641 -7404
rect 5053 -7437 6641 -7433
rect 4926 -7438 6641 -7437
rect 4825 -7478 6641 -7438
rect -35403 -7552 -33300 -7545
rect -35403 -7554 -35076 -7552
rect -35403 -7616 -35376 -7554
rect -35316 -7616 -35231 -7554
rect -35171 -7614 -35076 -7554
rect -35016 -7614 -33300 -7552
rect -20587 -7553 -20448 -7529
rect -35171 -7616 -33300 -7614
rect -35403 -7627 -33300 -7616
rect -68390 -7945 -68177 -7937
rect -68390 -8020 -68368 -7945
rect -68292 -8020 -68177 -7945
rect -68390 -8060 -68177 -8020
rect -66725 -7948 -66595 -7924
rect -66725 -8026 -66691 -7948
rect -66618 -8026 -66595 -7948
rect -66725 -8046 -66595 -8026
rect -64345 -8080 -64254 -8026
rect -64345 -8086 -64327 -8080
rect -64345 -8142 -64331 -8086
rect -64270 -8131 -64254 -8080
rect -43130 -8034 -42977 -8009
rect -43130 -8116 -43097 -8034
rect -43015 -8116 -42977 -8034
rect -64270 -8135 -63806 -8131
rect -64275 -8142 -63806 -8135
rect -64345 -8197 -63806 -8142
rect -64345 -8253 -64335 -8197
rect -64279 -8206 -63806 -8197
rect -64277 -8209 -63806 -8206
rect -43130 -8199 -42977 -8116
rect -64345 -8261 -64334 -8253
rect -64277 -8261 -64254 -8209
rect -64345 -8277 -64254 -8261
rect -52296 -8326 -52250 -8240
rect -43130 -8281 -43097 -8199
rect -43015 -8281 -42977 -8199
rect -43130 -8294 -42977 -8281
rect -19863 -8232 -19578 -8199
rect -19863 -8314 -19850 -8232
rect -19768 -8314 -19685 -8232
rect -19603 -8314 -19578 -8232
rect 18852 -8284 18898 -8197
rect -19863 -8352 -19578 -8314
rect 6460 -8328 6745 -8295
rect -56753 -8427 -54888 -8407
rect -56753 -8429 -54987 -8427
rect -65700 -8481 -63786 -8463
rect -65700 -8484 -65533 -8481
rect -65700 -8547 -65665 -8484
rect -65605 -8544 -65533 -8484
rect -65473 -8484 -63786 -8481
rect -65473 -8544 -65399 -8484
rect -65605 -8547 -65399 -8544
rect -65339 -8547 -63786 -8484
rect -56753 -8495 -55285 -8429
rect -55233 -8432 -54987 -8429
rect -55233 -8495 -55149 -8432
rect -56753 -8498 -55149 -8495
rect -55097 -8493 -54987 -8432
rect -54935 -8493 -54888 -8427
rect 6460 -8410 6473 -8328
rect 6555 -8410 6638 -8328
rect 6720 -8410 6745 -8328
rect 29536 -8334 29582 -8255
rect -36203 -8445 -34301 -8429
rect -36203 -8447 -34553 -8445
rect -55097 -8498 -54888 -8493
rect -56753 -8507 -54888 -8498
rect -65700 -8561 -63786 -8547
rect -66685 -8562 -63786 -8561
rect -66678 -8580 -63786 -8562
rect -44953 -8515 -43347 -8485
rect -44953 -8517 -44654 -8515
rect -44953 -8518 -44795 -8517
rect -44953 -8579 -44930 -8518
rect -44874 -8578 -44795 -8518
rect -44739 -8576 -44654 -8517
rect -44598 -8576 -43347 -8515
rect -36203 -8512 -34692 -8447
rect -34629 -8510 -34553 -8447
rect -34490 -8447 -34301 -8445
rect -34490 -8510 -34397 -8447
rect -34629 -8512 -34397 -8510
rect -34334 -8512 -34301 -8447
rect 6460 -8448 6745 -8410
rect -36203 -8529 -34301 -8512
rect -44739 -8578 -43347 -8576
rect -44874 -8579 -43347 -8578
rect -66678 -8708 -65422 -8580
rect -44953 -8602 -43347 -8579
rect -12732 -8557 -6739 -8543
rect -12732 -8565 -6841 -8557
rect -23396 -8613 -19640 -8599
rect -23396 -8618 -23115 -8613
rect -23396 -8703 -23378 -8618
rect -23292 -8698 -23115 -8618
rect -23029 -8698 -19640 -8613
rect -12732 -8631 -7135 -8565
rect -7074 -8631 -6998 -8565
rect -6937 -8623 -6841 -8565
rect -6780 -8623 -6739 -8557
rect -6937 -8631 -6739 -8623
rect -12732 -8643 -6739 -8631
rect -23292 -8703 -19640 -8698
rect -23396 -8716 -19640 -8703
rect 13690 -8676 15720 -8652
rect 4808 -8742 6670 -8708
rect 4808 -8746 5100 -8742
rect 4808 -8747 4973 -8746
rect 4808 -8801 4846 -8747
rect 4903 -8800 4973 -8747
rect 5030 -8796 5100 -8746
rect 5157 -8796 6670 -8742
rect 13690 -8736 15330 -8676
rect 15384 -8736 15461 -8676
rect 15515 -8678 15720 -8676
rect 15515 -8736 15602 -8678
rect 13690 -8738 15602 -8736
rect 15656 -8738 15720 -8678
rect 13690 -8752 15720 -8738
rect 5030 -8800 6670 -8796
rect 4903 -8801 6670 -8800
rect 4808 -8825 6670 -8801
rect -64134 -8908 -63744 -8886
rect -64134 -8970 -64126 -8908
rect -64070 -8954 -63744 -8908
rect -64070 -8970 -64066 -8954
rect -64134 -9048 -64066 -8970
rect -64134 -9110 -64125 -9048
rect -64069 -9110 -64066 -9048
rect -64134 -9128 -64066 -9110
rect 17304 -9304 17503 -9291
rect -53483 -9344 -53237 -9336
rect -63892 -9417 -63805 -9406
rect -63892 -9471 -63872 -9417
rect -63818 -9471 -63805 -9417
rect -61667 -9453 -60732 -9381
rect -53483 -9399 -53466 -9344
rect -53411 -9399 -53323 -9344
rect -53268 -9399 -53237 -9344
rect 17304 -9361 17316 -9304
rect 17373 -9359 17437 -9304
rect 17492 -9359 17653 -9304
rect 17373 -9361 17653 -9359
rect 28503 -9359 28587 -9341
rect 17304 -9368 17503 -9361
rect -53483 -9409 -53237 -9399
rect -43482 -9445 -43135 -9435
rect -63892 -9547 -63805 -9471
rect -43482 -9502 -43466 -9445
rect -43414 -9446 -43135 -9445
rect -43414 -9502 -43341 -9446
rect -43482 -9503 -43341 -9502
rect -43289 -9503 -43135 -9446
rect -41081 -9475 -40591 -9403
rect 28503 -9416 28516 -9359
rect 28573 -9416 28587 -9359
rect -4102 -9451 -3692 -9449
rect -4102 -9471 -3674 -9451
rect -43482 -9512 -43135 -9503
rect -4102 -9481 -3827 -9471
rect -63892 -9601 -63873 -9547
rect -63819 -9601 -63805 -9547
rect -63892 -9631 -63805 -9601
rect -55294 -9703 -53227 -9677
rect -55294 -9767 -55274 -9703
rect -55203 -9704 -53227 -9703
rect -55203 -9767 -55134 -9704
rect -55294 -9768 -55134 -9767
rect -55063 -9708 -53227 -9704
rect -55063 -9768 -54991 -9708
rect -55294 -9772 -54991 -9768
rect -54920 -9772 -53227 -9708
rect -55294 -9790 -53227 -9772
rect -46282 -9706 -44532 -9668
rect -46282 -9712 -44788 -9706
rect -55144 -10010 -55021 -9790
rect -46282 -9791 -44928 -9712
rect -44868 -9785 -44788 -9712
rect -44728 -9785 -44634 -9706
rect -44574 -9785 -44532 -9706
rect -44868 -9791 -44532 -9785
rect -46282 -9807 -44532 -9791
rect -33374 -9674 -32936 -9649
rect -33374 -9785 -33319 -9674
rect -33208 -9675 -32936 -9674
rect -33208 -9784 -33092 -9675
rect -32981 -9784 -32936 -9675
rect -33208 -9785 -32936 -9784
rect -65708 -10167 -62971 -10082
rect -56664 -10133 -55021 -10010
rect -44757 -10091 -44566 -9807
rect -33374 -9843 -32936 -9785
rect -26009 -10059 -22984 -10002
rect -44757 -10103 -34301 -10091
rect -65708 -10171 -65389 -10167
rect -65708 -10247 -65680 -10171
rect -65618 -10247 -65539 -10171
rect -65477 -10243 -65389 -10171
rect -65327 -10243 -62971 -10167
rect -65477 -10247 -62971 -10243
rect -65708 -10267 -62971 -10247
rect -44757 -10165 -32409 -10103
rect -26009 -10132 -23386 -10059
rect -23315 -10062 -22984 -10059
rect -23315 -10132 -23233 -10062
rect -26009 -10135 -23233 -10132
rect -23162 -10135 -23078 -10062
rect -23007 -10135 -22984 -10062
rect -26009 -10158 -22984 -10135
rect -44757 -10172 -34394 -10165
rect -44757 -10255 -34688 -10172
rect -34632 -10176 -34394 -10172
rect -34632 -10255 -34544 -10176
rect -44757 -10259 -34544 -10255
rect -34488 -10248 -34394 -10176
rect -34338 -10248 -32409 -10165
rect -34488 -10259 -32409 -10248
rect -44757 -10282 -34301 -10259
rect -33491 -10412 -33162 -10411
rect -19941 -10412 -19776 -9549
rect -17613 -9589 -16737 -9517
rect -4102 -9571 -4065 -9481
rect -3984 -9561 -3827 -9481
rect -3746 -9480 -3674 -9471
rect -3746 -9561 -3630 -9480
rect -3984 -9571 -3630 -9561
rect 28503 -9484 28587 -9416
rect 28503 -9543 28518 -9484
rect 28577 -9543 28587 -9484
rect 28503 -9570 28587 -9543
rect -4102 -9580 -3630 -9571
rect -4102 -9588 -3674 -9580
rect -4091 -9589 -3674 -9588
rect 3431 -9856 5232 -9819
rect 3431 -9858 5133 -9856
rect 3431 -9932 4844 -9858
rect 4899 -9860 5133 -9858
rect 4899 -9932 4983 -9860
rect 3431 -9934 4983 -9932
rect 5038 -9930 5133 -9860
rect 5188 -9930 5232 -9856
rect 5038 -9934 5232 -9930
rect 3431 -9951 5232 -9934
rect -12577 -10190 -6740 -10153
rect -12577 -10197 -6861 -10190
rect -12577 -10198 -7002 -10197
rect -12577 -10276 -7136 -10198
rect -7081 -10275 -7002 -10198
rect -6947 -10268 -6861 -10197
rect -6806 -10268 -6740 -10190
rect -6947 -10275 -6740 -10268
rect -7081 -10276 -6740 -10275
rect -12577 -10298 -6740 -10276
rect -4297 -10176 -3738 -10162
rect 6473 -10168 6603 -9657
rect 8809 -9698 9654 -9626
rect 15318 -9669 17709 -9638
rect 15318 -9672 15585 -9669
rect 15318 -9681 15463 -9672
rect 15318 -9737 15334 -9681
rect 15386 -9728 15463 -9681
rect 15515 -9725 15585 -9672
rect 15637 -9725 17709 -9669
rect 15515 -9728 17709 -9725
rect 15386 -9737 17709 -9728
rect 15318 -9751 17709 -9737
rect 24704 -9723 28295 -9693
rect 24704 -9726 26183 -9723
rect 6176 -10176 6613 -10168
rect -4297 -10177 6613 -10176
rect -4297 -10204 6184 -10177
rect -4297 -10205 -4047 -10204
rect -4297 -10277 -4274 -10205
rect -4202 -10277 -4047 -10205
rect -4297 -10278 -4047 -10277
rect -3973 -10205 6184 -10204
rect -3973 -10277 -3844 -10205
rect -3772 -10277 6184 -10205
rect -3973 -10278 6184 -10277
rect -4297 -10305 6184 -10278
rect 6312 -10305 6474 -10177
rect 6602 -10305 6613 -10177
rect -4297 -10306 6613 -10305
rect -4297 -10307 -3738 -10306
rect 6176 -10319 6613 -10306
rect -53363 -10455 -19776 -10412
rect -53363 -10458 -33282 -10455
rect -53363 -10467 -33437 -10458
rect -53363 -10543 -53325 -10467
rect -53248 -10470 -33437 -10467
rect -53248 -10539 -53170 -10470
rect -53103 -10527 -33437 -10470
rect -33371 -10523 -33282 -10458
rect -33205 -10523 -19776 -10455
rect 6918 -10523 7082 -10135
rect 15386 -10238 15573 -9751
rect 24704 -9789 26051 -9726
rect 26111 -9786 26183 -9726
rect 26243 -9726 28295 -9723
rect 26243 -9786 26317 -9726
rect 26111 -9789 26317 -9786
rect 26377 -9789 28295 -9726
rect 24704 -9806 28295 -9789
rect 13870 -10425 15573 -10238
rect 17517 -10523 17681 -9940
rect -33371 -10527 -19776 -10523
rect -53103 -10539 -19776 -10527
rect -53248 -10543 -19776 -10539
rect -53363 -10577 -19776 -10543
rect -3497 -10561 17681 -10523
rect -3497 -10577 -3179 -10561
rect -3497 -10662 -3402 -10577
rect -3304 -10646 -3179 -10577
rect -3081 -10646 -2936 -10561
rect -2838 -10646 17681 -10561
rect -3304 -10662 17681 -10646
rect -3497 -10687 17681 -10662
rect -33087 -10828 -32662 -10817
rect -20036 -10827 -19434 -10787
rect -20036 -10828 -20018 -10827
rect -52701 -10859 -20018 -10828
rect -52701 -10860 -33063 -10859
rect -52701 -10936 -52653 -10860
rect -52576 -10863 -33063 -10860
rect -52576 -10932 -52498 -10863
rect -52431 -10932 -33063 -10863
rect -52576 -10936 -33063 -10932
rect -52701 -10970 -33063 -10936
rect -32952 -10968 -32797 -10859
rect -32688 -10968 -20018 -10859
rect -32952 -10970 -20018 -10968
rect -52701 -10982 -20018 -10970
rect -19863 -10829 -19434 -10827
rect -19863 -10982 -19686 -10829
rect -19533 -10982 -19434 -10829
rect 17282 -10865 17758 -10855
rect 17282 -10866 17294 -10865
rect -52701 -10983 -19434 -10982
rect -33087 -10988 -32662 -10983
rect -20036 -11012 -19434 -10983
rect 6459 -10880 17294 -10866
rect 6459 -10992 6474 -10880
rect 6586 -10881 17294 -10880
rect 6586 -10991 6747 -10881
rect 6857 -10991 17294 -10881
rect 6586 -10992 17294 -10991
rect 6459 -11004 17294 -10992
rect 17433 -10867 17758 -10865
rect 17433 -11004 17605 -10867
rect 17742 -11004 17758 -10867
rect 6753 -11005 17758 -11004
rect 17282 -11018 17758 -11005
rect 29200 -11130 29374 -10992
rect 29200 -11230 29254 -11130
rect 29339 -11230 29374 -11130
rect 29200 -11284 29374 -11230
rect 16985 -11301 29377 -11284
rect -20587 -11439 -20448 -11363
rect 16985 -11437 16996 -11301
rect 17131 -11306 29377 -11301
rect 17131 -11406 29243 -11306
rect 29328 -11406 29377 -11306
rect 17131 -11437 29377 -11406
rect 16039 -11439 16215 -11438
rect -20587 -11503 16215 -11439
rect -20587 -11618 -20562 -11503
rect -20476 -11530 16215 -11503
rect -20476 -11606 16091 -11530
rect 16172 -11606 16215 -11530
rect -20476 -11613 16215 -11606
rect 16985 -11458 29377 -11437
rect -20476 -11618 -20448 -11613
rect -20587 -11704 -20448 -11618
rect -20587 -11819 -20565 -11704
rect -20479 -11819 -20448 -11704
rect -20587 -11849 -20448 -11819
rect 16039 -11738 16215 -11613
rect 16039 -11814 16087 -11738
rect 16168 -11814 16215 -11738
rect 16039 -11855 16215 -11814
rect 16663 -11623 16822 -11607
rect 16663 -11759 16675 -11623
rect 16810 -11759 16822 -11623
rect 16039 -11858 16213 -11855
rect 16663 -11977 16822 -11759
rect 16985 -11634 17147 -11458
rect 16985 -11770 16996 -11634
rect 17131 -11770 17147 -11634
rect 16985 -11785 17147 -11770
rect 6238 -12002 6393 -11997
rect -18615 -12006 6393 -12002
rect -18626 -12060 6393 -12006
rect -18626 -12176 -18597 -12060
rect -18509 -12133 6271 -12060
rect 6370 -12133 6393 -12060
rect 16663 -12113 16675 -11977
rect 16810 -11982 16822 -11977
rect 28489 -11974 28601 -11925
rect 28489 -11982 28521 -11974
rect 16810 -12026 28521 -11982
rect 28576 -11982 28601 -11974
rect 28576 -12026 28617 -11982
rect 16810 -12109 28617 -12026
rect 16810 -12113 28512 -12109
rect 16663 -12125 28512 -12113
rect -18509 -12176 6393 -12133
rect 16671 -12156 28512 -12125
rect -18626 -12193 6393 -12176
rect 28489 -12161 28512 -12156
rect 28567 -12156 28617 -12109
rect 28567 -12161 28601 -12156
rect 28489 -12182 28601 -12161
rect -18626 -12289 -18480 -12193
rect -64587 -12362 -64502 -12343
rect -64587 -12450 -64575 -12362
rect -64516 -12450 -64502 -12362
rect -18626 -12405 -18596 -12289
rect -18508 -12405 -18480 -12289
rect -64587 -12536 -64502 -12450
rect -64587 -12624 -64573 -12536
rect -64514 -12557 -64502 -12536
rect -43801 -12447 -43647 -12424
rect -18626 -12434 -18480 -12405
rect 6238 -12216 6393 -12193
rect 6238 -12289 6271 -12216
rect 6370 -12289 6393 -12216
rect 6238 -12372 6393 -12289
rect -64514 -12584 -54219 -12557
rect -64514 -12624 -54294 -12584
rect -64587 -12643 -54294 -12624
rect -64587 -12644 -64502 -12643
rect -54305 -12674 -54294 -12643
rect -54231 -12674 -54219 -12584
rect -54305 -12779 -54219 -12674
rect -43801 -12607 -43772 -12447
rect -43666 -12607 -43647 -12447
rect 6238 -12445 6266 -12372
rect 6365 -12445 6393 -12372
rect 6238 -12479 6393 -12445
rect -43801 -12718 -43647 -12607
rect -34043 -12718 -33918 -12712
rect -54305 -12869 -54295 -12779
rect -54232 -12869 -54219 -12779
rect -54305 -12884 -54219 -12869
rect -43804 -12727 -33918 -12718
rect -32608 -12724 -5517 -12723
rect -43804 -12887 -43777 -12727
rect -43671 -12765 -33918 -12727
rect -43671 -12869 -34022 -12765
rect -33936 -12869 -33918 -12765
rect -43671 -12887 -33918 -12869
rect -43804 -12915 -33918 -12887
rect -34043 -13019 -33918 -12915
rect -34043 -13123 -34025 -13019
rect -33939 -13123 -33918 -13019
rect -32624 -12772 -5517 -12724
rect -32624 -12876 -32602 -12772
rect -32524 -12870 -5637 -12772
rect -5540 -12870 -5517 -12772
rect -32524 -12872 -5517 -12870
rect -32524 -12876 -32507 -12872
rect -32624 -12973 -32507 -12876
rect -32624 -13077 -32608 -12973
rect -32530 -13077 -32507 -12973
rect -32624 -13093 -32507 -13077
rect -5666 -13002 -5517 -12872
rect -5666 -13100 -5645 -13002
rect -5548 -13100 -5517 -13002
rect -5666 -13119 -5517 -13100
rect -34043 -13148 -33918 -13123
rect -53775 -13188 -53370 -13171
rect -53775 -13293 -53761 -13188
rect -53656 -13291 -53489 -13188
rect -53386 -13291 -53370 -13188
rect -53656 -13293 -53370 -13291
rect -53775 -13308 -53370 -13293
rect -56214 -13497 -53302 -13469
rect -56214 -13499 -55000 -13497
rect -56214 -13500 -55137 -13499
rect -65699 -13570 -60761 -13554
rect -65699 -13643 -65682 -13570
rect -65611 -13571 -60761 -13570
rect -65611 -13643 -65551 -13571
rect -65699 -13644 -65551 -13643
rect -65480 -13576 -60761 -13571
rect -65480 -13644 -65395 -13576
rect -65699 -13649 -65395 -13644
rect -65324 -13649 -60761 -13576
rect -56214 -13568 -55276 -13500
rect -55214 -13567 -55137 -13500
rect -55075 -13565 -55000 -13499
rect -54938 -13565 -53302 -13497
rect -55075 -13567 -53302 -13565
rect -55214 -13568 -53302 -13567
rect -56214 -13582 -53302 -13568
rect -46207 -13492 -40640 -13430
rect -46207 -13494 -44803 -13492
rect -46207 -13563 -44924 -13494
rect -44870 -13561 -44803 -13494
rect -44749 -13561 -44652 -13492
rect -44598 -13561 -40640 -13492
rect -44870 -13563 -40640 -13561
rect -46207 -13594 -40640 -13563
rect -65699 -13755 -60761 -13649
rect -40804 -13604 -40640 -13594
rect -65699 -13761 -65534 -13755
rect -65699 -13834 -65685 -13761
rect -65614 -13828 -65534 -13761
rect -65463 -13756 -60761 -13755
rect -65463 -13828 -65392 -13756
rect -65614 -13829 -65392 -13828
rect -65321 -13829 -60761 -13756
rect -65614 -13834 -60761 -13829
rect -65699 -13847 -60761 -13834
rect -54012 -13738 -53926 -13730
rect -54012 -13795 -53999 -13738
rect -53942 -13795 -53926 -13738
rect -40804 -13768 -37994 -13604
rect -24860 -13606 -11760 -13578
rect -24860 -13611 -23091 -13606
rect -24860 -13614 -23248 -13611
rect -29397 -13714 -29343 -13673
rect -24860 -13695 -23388 -13614
rect -23327 -13692 -23248 -13614
rect -23187 -13687 -23091 -13611
rect -23030 -13687 -11760 -13606
rect -1236 -13659 -1118 -13529
rect 3345 -13533 9653 -13512
rect 3345 -13536 5122 -13533
rect 3345 -13610 4844 -13536
rect 4907 -13539 5122 -13536
rect 4907 -13610 5001 -13539
rect 3345 -13613 5001 -13610
rect 5064 -13607 5122 -13539
rect 5185 -13607 9653 -13533
rect 25122 -13571 31184 -13544
rect 25122 -13579 26180 -13571
rect 5064 -13613 9653 -13607
rect 3345 -13624 9653 -13613
rect -23187 -13692 -11760 -13687
rect -23327 -13695 -11760 -13692
rect -24860 -13707 -11760 -13695
rect -10867 -13688 -1118 -13659
rect -35815 -13749 -29341 -13714
rect -35815 -13755 -34539 -13749
rect -54012 -13859 -53926 -13795
rect -35815 -13820 -34681 -13755
rect -34623 -13814 -34539 -13755
rect -34481 -13757 -29341 -13749
rect -34481 -13814 -34394 -13757
rect -34623 -13820 -34394 -13814
rect -35815 -13822 -34394 -13820
rect -34336 -13822 -29341 -13757
rect -10867 -13752 -7132 -13688
rect -7080 -13692 -6827 -13688
rect -7080 -13752 -6994 -13692
rect -10867 -13756 -6994 -13752
rect -6942 -13752 -6827 -13692
rect -6775 -13752 -1118 -13688
rect -6942 -13756 -1118 -13752
rect -10867 -13777 -1118 -13756
rect 9541 -13763 9653 -13624
rect 14265 -13597 14373 -13594
rect 14265 -13626 14380 -13597
rect 15098 -13626 20464 -13615
rect 14265 -13652 20464 -13626
rect 14265 -13654 15467 -13652
rect 14265 -13727 15328 -13654
rect 15382 -13725 15467 -13654
rect 15521 -13654 20464 -13652
rect 15521 -13725 15611 -13654
rect 15382 -13727 15611 -13725
rect 15665 -13727 20464 -13654
rect 25122 -13657 26027 -13579
rect 26088 -13649 26180 -13579
rect 26241 -13572 31184 -13571
rect 26241 -13649 26339 -13572
rect 26088 -13650 26339 -13649
rect 26400 -13650 31184 -13572
rect 26088 -13657 31184 -13650
rect 25122 -13669 31184 -13657
rect 14265 -13741 20464 -13727
rect 14272 -13744 14380 -13741
rect 15098 -13750 20464 -13741
rect 31059 -13800 31184 -13669
rect -54012 -13860 -53466 -13859
rect -54012 -13915 -53999 -13860
rect -53944 -13915 -53466 -13860
rect -54012 -13916 -53466 -13915
rect -35815 -13916 -29341 -13822
rect -54012 -13923 -53926 -13916
rect -35815 -13924 -34387 -13916
rect -35815 -13927 -34547 -13924
rect -35815 -13992 -34693 -13927
rect -34635 -13989 -34547 -13927
rect -34489 -13981 -34387 -13924
rect -34329 -13981 -29341 -13916
rect -34489 -13989 -29341 -13981
rect -34635 -13992 -29341 -13989
rect -35815 -14000 -29341 -13992
rect -7914 -14459 -4087 -14426
rect -66381 -14518 -63937 -14464
rect -66381 -14521 -66217 -14518
rect -66381 -14584 -66349 -14521
rect -66289 -14581 -66217 -14521
rect -66157 -14521 -63937 -14518
rect -66157 -14581 -66083 -14521
rect -66289 -14584 -66083 -14581
rect -66023 -14584 -63937 -14521
rect -66381 -14614 -63937 -14584
rect -35391 -14543 -32453 -14501
rect -35391 -14544 -35093 -14543
rect -35391 -14547 -35245 -14544
rect -35391 -14627 -35385 -14547
rect -35314 -14624 -35245 -14547
rect -35174 -14623 -35093 -14544
rect -35022 -14623 -32453 -14543
rect -7914 -14546 -7903 -14459
rect -7831 -14546 -7762 -14459
rect -7690 -14460 -4087 -14459
rect -7690 -14546 -7624 -14460
rect -7914 -14547 -7624 -14546
rect -7552 -14547 -4087 -14460
rect -7914 -14576 -4087 -14547
rect 4069 -14435 6522 -14400
rect 4069 -14436 4214 -14435
rect 4069 -14531 4077 -14436
rect 4149 -14530 4214 -14436
rect 4286 -14530 4359 -14435
rect 4431 -14530 6522 -14435
rect 4149 -14531 6522 -14530
rect 4069 -14550 6522 -14531
rect 14607 -14527 17358 -14465
rect -35174 -14624 -32453 -14623
rect -35314 -14627 -32453 -14624
rect -45762 -14674 -43501 -14633
rect -35391 -14651 -32453 -14627
rect -24189 -14610 -18303 -14576
rect -24189 -14613 -23911 -14610
rect -24189 -14614 -24046 -14613
rect -45762 -14675 -45492 -14674
rect -45762 -14678 -45627 -14675
rect -45762 -14744 -45753 -14678
rect -45681 -14741 -45627 -14678
rect -45555 -14740 -45492 -14675
rect -45420 -14740 -43501 -14674
rect -24189 -14699 -24181 -14614
rect -24108 -14698 -24046 -14614
rect -23973 -14695 -23911 -14613
rect -23838 -14695 -18303 -14610
rect 14607 -14583 14645 -14527
rect 14697 -14583 14761 -14527
rect 14813 -14531 17358 -14527
rect 14813 -14583 14876 -14531
rect 14607 -14587 14876 -14583
rect 14928 -14587 17358 -14531
rect 14607 -14615 17358 -14587
rect 25328 -14490 27997 -14440
rect 25328 -14493 25492 -14490
rect 25328 -14556 25360 -14493
rect 25420 -14553 25492 -14493
rect 25552 -14493 27997 -14490
rect 25552 -14553 25626 -14493
rect 25420 -14556 25626 -14553
rect 25686 -14556 27997 -14493
rect 25328 -14590 27997 -14556
rect -23973 -14698 -18303 -14695
rect -24108 -14699 -18303 -14698
rect -24189 -14726 -18303 -14699
rect -45555 -14741 -43501 -14740
rect -45681 -14744 -43501 -14741
rect -45762 -14783 -43501 -14744
rect -5302 -14862 -5188 -14822
rect -63347 -14909 -63260 -14888
rect -63347 -14965 -63334 -14909
rect -63278 -14965 -63260 -14909
rect -63347 -15020 -63260 -14965
rect -5302 -14941 -5277 -14862
rect -5207 -14928 -5188 -14862
rect -3682 -14879 -3595 -14858
rect -5207 -14941 -4067 -14928
rect -63347 -15076 -63338 -15020
rect -63282 -15076 -63260 -15020
rect -63347 -15091 -63260 -15076
rect -31868 -14996 -31781 -14975
rect -31868 -15052 -31855 -14996
rect -31799 -15052 -31781 -14996
rect -5302 -15010 -4067 -14941
rect -3682 -14935 -3669 -14879
rect -3613 -14935 -3595 -14879
rect -3682 -14990 -3595 -14935
rect -5302 -15045 -5188 -15010
rect -42985 -15099 -42898 -15078
rect -42985 -15155 -42972 -15099
rect -42916 -15155 -42898 -15099
rect -52249 -15245 -52203 -15158
rect -42985 -15210 -42898 -15155
rect -31868 -15107 -31781 -15052
rect -31868 -15163 -31859 -15107
rect -31803 -15163 -31781 -15107
rect -31868 -15178 -31781 -15163
rect -17864 -15072 -17777 -15051
rect -17864 -15128 -17851 -15072
rect -17795 -15128 -17777 -15072
rect -42985 -15266 -42976 -15210
rect -42920 -15266 -42898 -15210
rect -17864 -15183 -17777 -15128
rect -5302 -15124 -5281 -15045
rect -5211 -15124 -5188 -15045
rect -3682 -15046 -3673 -14990
rect -3617 -15046 -3595 -14990
rect 7092 -14862 7179 -14841
rect 7092 -14918 7105 -14862
rect 7161 -14918 7179 -14862
rect 7092 -14973 7179 -14918
rect 7092 -15029 7101 -14973
rect 7157 -15029 7179 -14973
rect 7092 -15044 7179 -15029
rect 17933 -14910 18020 -14889
rect 17933 -14966 17946 -14910
rect 18002 -14966 18020 -14910
rect 17933 -15021 18020 -14966
rect -3682 -15061 -3595 -15046
rect 17933 -15077 17942 -15021
rect 17998 -15077 18020 -15021
rect 17933 -15092 18020 -15077
rect 28638 -14904 28725 -14883
rect 28638 -14960 28651 -14904
rect 28707 -14960 28725 -14904
rect 28638 -15015 28725 -14960
rect 28638 -15071 28647 -15015
rect 28703 -15071 28725 -15015
rect 28638 -15086 28725 -15071
rect -5302 -15137 -5188 -15124
rect -17864 -15239 -17855 -15183
rect -17799 -15239 -17777 -15183
rect -17864 -15254 -17777 -15239
rect -42985 -15281 -42898 -15266
rect -32618 -15769 -32515 -15657
rect -32618 -15868 -32597 -15769
rect -32527 -15868 -32515 -15769
rect -64604 -15912 -64505 -15877
rect -64604 -15982 -64593 -15912
rect -64520 -15935 -64505 -15912
rect -55941 -15924 -53557 -15915
rect -55941 -15925 -55624 -15924
rect -64520 -15982 -63988 -15935
rect -64604 -16009 -63988 -15982
rect -55941 -15983 -55915 -15925
rect -55862 -15983 -55771 -15925
rect -55718 -15982 -55624 -15925
rect -55571 -15982 -53557 -15924
rect -55718 -15983 -53557 -15982
rect -55941 -15997 -53557 -15983
rect -32618 -15949 -32515 -15868
rect -64604 -16094 -64505 -16009
rect -64604 -16164 -64593 -16094
rect -64520 -16164 -64505 -16094
rect -64604 -16181 -64505 -16164
rect -43849 -16048 -43697 -16005
rect -43849 -16137 -43829 -16048
rect -43717 -16104 -43697 -16048
rect -32618 -16048 -32602 -15949
rect -32532 -16048 -32515 -15949
rect -32618 -16071 -32515 -16048
rect -18626 -15808 -18480 -15630
rect -18626 -15909 -18605 -15808
rect -18507 -15909 -18480 -15808
rect -18626 -16003 -18480 -15909
rect -18626 -16104 -18600 -16003
rect -18502 -16104 -18480 -16003
rect -43717 -16137 -43582 -16104
rect -18626 -16133 -18480 -16104
rect -5606 -15818 -5520 -15777
rect -5606 -15871 -5589 -15818
rect -5532 -15871 -5520 -15818
rect -5606 -15897 -5520 -15871
rect 6272 -15840 6361 -15742
rect -5606 -15937 -4052 -15897
rect -5606 -15990 -5594 -15937
rect -5537 -15971 -4052 -15937
rect 6272 -15919 6286 -15840
rect 6347 -15871 6361 -15840
rect 6347 -15919 6447 -15871
rect 6272 -15945 6447 -15919
rect 16367 -15936 16458 -15889
rect 26019 -15897 26394 -15882
rect 26019 -15900 26173 -15897
rect 26019 -15911 26041 -15900
rect -5537 -15990 -5520 -15971
rect -5606 -16050 -5520 -15990
rect -5606 -16103 -5592 -16050
rect -5535 -16103 -5520 -16050
rect -5606 -16121 -5520 -16103
rect 6272 -16023 6361 -15945
rect 6272 -16102 6285 -16023
rect 6346 -16102 6361 -16023
rect 6272 -16121 6361 -16102
rect 16367 -15950 17315 -15936
rect 16367 -16020 16378 -15950
rect 16441 -16010 17315 -15950
rect 26014 -15963 26041 -15911
rect 26101 -15960 26173 -15900
rect 26233 -15900 26394 -15897
rect 26233 -15960 26307 -15900
rect 26101 -15963 26307 -15960
rect 26367 -15911 26394 -15900
rect 26367 -15963 28036 -15911
rect 26014 -15985 28036 -15963
rect 16441 -16020 16458 -16010
rect -5598 -16123 -5524 -16121
rect -43849 -16178 -43582 -16137
rect 16367 -16138 16458 -16020
rect -43849 -16278 -43697 -16178
rect 16367 -16208 16380 -16138
rect 16443 -16208 16458 -16138
rect 16367 -16223 16458 -16208
rect 16378 -16225 16452 -16223
rect -43849 -16367 -43832 -16278
rect -43720 -16367 -43697 -16278
rect -43849 -16393 -43697 -16367
rect -64349 -16760 -64248 -16748
rect -64349 -16838 -64337 -16760
rect -64259 -16838 -64248 -16760
rect -4046 -16754 -3896 -16730
rect -64349 -16907 -64248 -16838
rect -32218 -16809 -32087 -16789
rect -63669 -16879 -63582 -16858
rect -64349 -16908 -63923 -16907
rect -64349 -16984 -64336 -16908
rect -64260 -16984 -63923 -16908
rect -64349 -16985 -63923 -16984
rect -63669 -16935 -63656 -16879
rect -63600 -16935 -63582 -16879
rect -64349 -17004 -64248 -16985
rect -63669 -16990 -63582 -16935
rect -32218 -16887 -32183 -16809
rect -32114 -16887 -32087 -16809
rect -63669 -17046 -63660 -16990
rect -63604 -17046 -63582 -16990
rect -63669 -17061 -63582 -17046
rect -43337 -16972 -43250 -16951
rect -43337 -17028 -43324 -16972
rect -43268 -17028 -43250 -16972
rect -43337 -17083 -43250 -17028
rect -32218 -16991 -32087 -16887
rect -4931 -16795 -4841 -16778
rect -4931 -16859 -4920 -16795
rect -4856 -16859 -4841 -16795
rect -4931 -16869 -4841 -16859
rect -4046 -16819 -4002 -16754
rect -3932 -16819 -3896 -16754
rect -32218 -17069 -32183 -16991
rect -32114 -17069 -32087 -16991
rect -32218 -17083 -32087 -17069
rect -18454 -16969 -18169 -16936
rect -18454 -17051 -18441 -16969
rect -18359 -17051 -18276 -16969
rect -18194 -17051 -18169 -16969
rect -4931 -16943 -4074 -16869
rect -4931 -17007 -4923 -16943
rect -4859 -16947 -4074 -16943
rect -4046 -16913 -3896 -16819
rect -4859 -17007 -4841 -16947
rect -4046 -16978 -4008 -16913
rect -3938 -16978 -3896 -16913
rect -4046 -16995 -3896 -16978
rect 6633 -16765 6771 -16748
rect 6633 -16836 6667 -16765
rect 6738 -16836 6771 -16765
rect 28305 -16761 28443 -16744
rect 6633 -16941 6771 -16836
rect -4931 -17022 -4841 -17007
rect 6633 -17012 6663 -16941
rect 6734 -17012 6771 -16941
rect 6633 -17022 6771 -17012
rect 17414 -16820 17552 -16803
rect 17414 -16891 17448 -16820
rect 17519 -16891 17552 -16820
rect 17414 -16996 17552 -16891
rect -43337 -17139 -43328 -17083
rect -43272 -17139 -43250 -17083
rect -18454 -17089 -18169 -17051
rect 17414 -17067 17444 -16996
rect 17515 -17067 17552 -16996
rect 28305 -16832 28339 -16761
rect 28410 -16832 28443 -16761
rect 28305 -16937 28443 -16832
rect 28305 -17008 28335 -16937
rect 28406 -17008 28443 -16937
rect 28305 -17018 28443 -17008
rect 17414 -17077 17552 -17067
rect -43337 -17154 -43250 -17139
rect 2932 -17175 5232 -17145
rect -56753 -17196 -54894 -17183
rect -56753 -17198 -54986 -17196
rect -65695 -17265 -63716 -17239
rect -65695 -17268 -65540 -17265
rect -65695 -17331 -65672 -17268
rect -65612 -17328 -65540 -17268
rect -65480 -17268 -63716 -17265
rect -65480 -17328 -65406 -17268
rect -65612 -17331 -65406 -17328
rect -65346 -17331 -63716 -17268
rect -56753 -17266 -55285 -17198
rect -55233 -17266 -55152 -17198
rect -55100 -17264 -54986 -17198
rect -54934 -17264 -54894 -17196
rect 2932 -17196 6678 -17175
rect 2932 -17199 4966 -17196
rect -55100 -17266 -54894 -17264
rect -56753 -17283 -54894 -17266
rect -65695 -17356 -63716 -17331
rect -34701 -17307 -32284 -17276
rect -34701 -17309 -34438 -17307
rect -34701 -17311 -34572 -17309
rect -34701 -17352 -34694 -17311
rect -36365 -17378 -34694 -17352
rect -34636 -17376 -34572 -17311
rect -34514 -17374 -34438 -17309
rect -34380 -17374 -32284 -17307
rect -25269 -17320 -23457 -17220
rect -7145 -17226 -4097 -17201
rect -7145 -17229 -6871 -17226
rect -7145 -17230 -7005 -17229
rect -7145 -17295 -7135 -17230
rect -7080 -17294 -7005 -17230
rect -6950 -17291 -6871 -17229
rect -6816 -17291 -4097 -17226
rect 2932 -17245 4843 -17199
rect -6950 -17294 -4097 -17291
rect 4834 -17269 4843 -17245
rect 4901 -17266 4966 -17199
rect 5024 -17197 6678 -17196
rect 5024 -17266 5105 -17197
rect 4901 -17267 5105 -17266
rect 5163 -17267 6678 -17197
rect 13698 -17219 15671 -17119
rect 4901 -17269 6678 -17267
rect 4834 -17292 6678 -17269
rect 15286 -17240 15671 -17219
rect 24542 -17215 26130 -17184
rect 15286 -17266 17579 -17240
rect 15286 -17273 15588 -17266
rect 15286 -17278 15472 -17273
rect 15304 -17280 15472 -17278
rect -7080 -17295 -4097 -17294
rect -34514 -17376 -32284 -17374
rect -34636 -17378 -32284 -17376
rect -36365 -17393 -32284 -17378
rect -23557 -17330 -23457 -17320
rect -11256 -17318 -4097 -17295
rect -23557 -17351 -23015 -17330
rect -23557 -17377 -18280 -17351
rect -23557 -17382 -23120 -17377
rect -44940 -17444 -43264 -17408
rect -44940 -17502 -44930 -17444
rect -44876 -17445 -44652 -17444
rect -44876 -17502 -44802 -17445
rect -44940 -17503 -44802 -17502
rect -44748 -17502 -44652 -17445
rect -44598 -17502 -43264 -17444
rect -36365 -17452 -34434 -17393
rect -23557 -17430 -23388 -17382
rect -23396 -17444 -23388 -17430
rect -23331 -17444 -23268 -17382
rect -23211 -17439 -23120 -17382
rect -23063 -17439 -18280 -17377
rect -11256 -17395 -6770 -17318
rect 15304 -17336 15331 -17280
rect 15383 -17329 15472 -17280
rect 15524 -17322 15588 -17273
rect 15640 -17322 17579 -17266
rect 24542 -17246 28295 -17215
rect 24542 -17249 26173 -17246
rect 24542 -17284 26041 -17249
rect 15524 -17329 17579 -17322
rect 15383 -17336 17579 -17329
rect 26010 -17312 26041 -17284
rect 26101 -17309 26173 -17249
rect 26233 -17249 28295 -17246
rect 26233 -17309 26307 -17249
rect 26101 -17312 26307 -17309
rect 26367 -17312 28295 -17249
rect 26010 -17332 28295 -17312
rect 15304 -17357 17579 -17336
rect -23211 -17444 -18280 -17439
rect -23396 -17468 -18280 -17444
rect -44748 -17503 -43264 -17502
rect -44940 -17525 -43264 -17503
rect 17007 -17509 17122 -17491
rect 17007 -17575 17042 -17509
rect 17108 -17575 17122 -17509
rect -64133 -17685 -63916 -17662
rect -64133 -17747 -64123 -17685
rect -64070 -17730 -63916 -17685
rect 17007 -17663 17122 -17575
rect 27805 -17638 27909 -17616
rect 27805 -17639 28096 -17638
rect 17007 -17698 17516 -17663
rect -64070 -17747 -64065 -17730
rect -64133 -17822 -64065 -17747
rect 17007 -17764 17042 -17698
rect 17108 -17731 17516 -17698
rect 27805 -17705 27827 -17639
rect 27893 -17705 28096 -17639
rect 27805 -17706 28096 -17705
rect 17108 -17764 17122 -17731
rect 17007 -17787 17122 -17764
rect -64133 -17884 -64123 -17822
rect -64070 -17884 -64065 -17822
rect -64133 -17906 -64065 -17884
rect 27805 -17804 27909 -17706
rect 27805 -17872 27826 -17804
rect 27894 -17872 27909 -17804
rect 27805 -17892 27909 -17872
rect 16683 -18022 16795 -17995
rect -53675 -18065 -53342 -18044
rect -53675 -18140 -53634 -18065
rect -53560 -18070 -53342 -18065
rect -53560 -18134 -53451 -18070
rect -53377 -18134 -53290 -18070
rect -53560 -18140 -53290 -18134
rect -63894 -18200 -63798 -18152
rect -53675 -18155 -53342 -18140
rect -4047 -18152 -3949 -18142
rect -63894 -18254 -63867 -18200
rect -63815 -18254 -63798 -18200
rect -61638 -18229 -60691 -18157
rect -32294 -18226 -32192 -18212
rect -32294 -18227 -32110 -18226
rect -63894 -18332 -63798 -18254
rect -32294 -18302 -32277 -18227
rect -32202 -18302 -32110 -18227
rect -30159 -18266 -29281 -18194
rect -4047 -18227 -4042 -18152
rect -3966 -18227 -3949 -18152
rect -1972 -18191 -1041 -18119
rect 6712 -18133 6791 -18122
rect -18323 -18285 -18198 -18284
rect -32294 -18303 -32110 -18302
rect -63894 -18386 -63868 -18332
rect -63816 -18386 -63798 -18332
rect -63894 -18407 -63798 -18386
rect -46238 -18416 -44539 -18383
rect -46238 -18417 -44640 -18416
rect -46238 -18419 -44785 -18417
rect -46238 -18503 -44929 -18419
rect -44866 -18501 -44785 -18419
rect -44722 -18500 -44640 -18417
rect -44577 -18500 -44539 -18416
rect -44722 -18501 -44539 -18500
rect -44866 -18503 -44539 -18501
rect -46238 -18526 -44539 -18503
rect -54006 -18782 -53911 -18773
rect -54006 -18783 -53396 -18782
rect -56596 -18836 -54888 -18789
rect -56596 -18845 -54983 -18836
rect -56596 -18848 -55139 -18845
rect -63905 -18983 -63795 -18901
rect -56596 -18934 -55280 -18848
rect -55214 -18931 -55139 -18848
rect -55073 -18922 -54983 -18845
rect -54917 -18922 -54888 -18836
rect -55073 -18931 -54888 -18922
rect -55214 -18934 -54888 -18931
rect -56596 -18950 -54888 -18934
rect -54006 -18855 -53991 -18783
rect -53919 -18855 -53396 -18783
rect -54006 -18856 -53396 -18855
rect -54006 -18925 -53911 -18856
rect -54006 -18946 -53907 -18925
rect -63905 -19056 -63886 -18983
rect -63807 -19056 -63795 -18983
rect -54006 -19016 -53992 -18946
rect -63905 -19076 -63795 -19056
rect -54019 -19020 -53992 -19016
rect -53918 -19020 -53907 -18946
rect -54019 -19076 -53907 -19020
rect -63905 -19169 -53907 -19076
rect -63905 -19242 -63889 -19169
rect -63810 -19170 -53907 -19169
rect -63810 -19242 -63795 -19170
rect -63905 -19270 -63795 -19242
rect -53765 -19238 -53660 -19187
rect -53765 -19331 -53748 -19238
rect -53671 -19331 -53660 -19238
rect -64167 -19368 -64043 -19366
rect -53765 -19368 -53660 -19331
rect -64167 -19387 -53660 -19368
rect -64167 -19403 -53751 -19387
rect -64167 -19471 -64144 -19403
rect -64064 -19471 -53751 -19403
rect -64167 -19480 -53751 -19471
rect -53674 -19480 -53660 -19387
rect -64167 -19494 -53660 -19480
rect -64167 -19589 -64041 -19494
rect -53765 -19501 -53660 -19494
rect -64167 -19657 -64145 -19589
rect -64065 -19657 -64041 -19589
rect -64167 -19680 -64041 -19657
rect -43363 -19621 -43256 -18355
rect -41258 -18398 -40472 -18326
rect -32294 -18394 -32192 -18303
rect -18423 -18319 -18107 -18285
rect -18423 -18320 -18206 -18319
rect -18423 -18381 -18383 -18320
rect -18329 -18380 -18206 -18320
rect -18152 -18380 -18107 -18319
rect -16130 -18341 -15397 -18269
rect -4047 -18315 -3949 -18227
rect -18329 -18381 -18107 -18380
rect -32294 -18395 -32191 -18394
rect -32294 -18472 -32277 -18395
rect -32200 -18472 -32191 -18395
rect -18423 -18410 -18107 -18381
rect -4047 -18390 -4033 -18315
rect -3958 -18390 -3949 -18315
rect 6712 -18194 6721 -18133
rect 6780 -18194 6791 -18133
rect 8784 -18165 9653 -18093
rect 16683 -18099 16702 -18022
rect 16779 -18099 16795 -18022
rect 6712 -18261 6791 -18194
rect 6712 -18322 6724 -18261
rect 6783 -18322 6791 -18261
rect 16683 -18190 16795 -18099
rect 28109 -18017 28214 -18000
rect 28109 -18094 28123 -18017
rect 28200 -18094 28214 -18017
rect 16683 -18191 17483 -18190
rect 16683 -18266 16703 -18191
rect 16778 -18266 17483 -18191
rect 19648 -18230 20167 -18158
rect 28109 -18165 28214 -18094
rect 28109 -18166 28280 -18165
rect 16683 -18267 17483 -18266
rect 28109 -18241 28124 -18166
rect 28199 -18241 28280 -18166
rect 30349 -18205 31163 -18133
rect 28109 -18242 28280 -18241
rect 16683 -18290 16795 -18267
rect 28109 -18278 28214 -18242
rect 6712 -18359 6791 -18322
rect -18322 -18412 -18197 -18410
rect -4047 -18413 -3949 -18390
rect -32294 -18473 -32191 -18472
rect -32294 -18486 -32192 -18473
rect -43091 -19318 -42989 -18842
rect -36202 -18983 -34286 -18956
rect -31727 -18983 -22982 -18966
rect -36202 -19009 -22982 -18983
rect -36202 -19011 -23101 -19009
rect -36202 -19015 -23259 -19011
rect -36202 -19034 -23384 -19015
rect -36202 -19099 -34688 -19034
rect -34630 -19036 -23384 -19034
rect -34630 -19037 -34399 -19036
rect -34630 -19099 -34555 -19037
rect -36202 -19102 -34555 -19099
rect -34497 -19101 -34399 -19037
rect -34341 -19097 -23384 -19036
rect -23321 -19093 -23259 -19015
rect -23196 -19091 -23101 -19011
rect -23038 -19091 -22982 -19009
rect -23196 -19093 -22982 -19091
rect -23321 -19097 -22982 -19093
rect -34341 -19101 -22982 -19097
rect -34497 -19102 -22982 -19101
rect -36202 -19112 -22982 -19102
rect -36202 -19124 -34286 -19112
rect -17969 -19318 -17867 -18786
rect -11162 -18950 35409 -18881
rect -11162 -18955 -6833 -18950
rect -11162 -18963 -6992 -18955
rect -11162 -19027 -7129 -18963
rect -7077 -19019 -6992 -18963
rect -6940 -19014 -6833 -18955
rect -6781 -18951 35409 -18950
rect -6781 -18959 26321 -18951
rect -6781 -18961 5148 -18959
rect -6781 -19014 4848 -18961
rect -6940 -19019 4848 -19014
rect -7077 -19027 4848 -19019
rect -11162 -19035 4848 -19027
rect 4911 -19035 4986 -18961
rect 5049 -19033 5148 -18961
rect 5211 -18961 26321 -18959
rect 5211 -18970 26187 -18961
rect 5211 -18973 26035 -18970
rect 5211 -18974 15628 -18973
rect 5211 -19033 15336 -18974
rect 5049 -19035 15336 -19033
rect -11162 -19047 15336 -19035
rect 15390 -18975 15628 -18974
rect 15390 -19047 15472 -18975
rect -11162 -19048 15472 -19047
rect 15526 -19046 15628 -18975
rect 15682 -19046 26035 -18973
rect 15526 -19048 26035 -19046
rect 26096 -19039 26187 -18970
rect 26248 -19029 26321 -18961
rect 26382 -19029 35409 -18951
rect 26248 -19039 35409 -19029
rect 26096 -19048 35409 -19039
rect -11162 -19067 35409 -19048
rect -43091 -19337 -17867 -19318
rect -43091 -19393 -31960 -19337
rect -31904 -19393 -17867 -19337
rect -43091 -19420 -17867 -19393
rect -31978 -19459 -31879 -19420
rect -32298 -19528 -32195 -19513
rect -32298 -19589 -32280 -19528
rect -32218 -19589 -32195 -19528
rect -31978 -19515 -31954 -19459
rect -31898 -19515 -31879 -19459
rect -31978 -19543 -31879 -19515
rect -32298 -19621 -32195 -19589
rect -18352 -19620 -18003 -19604
rect -18352 -19621 -18124 -19620
rect -43363 -19622 -18124 -19621
rect -43363 -19656 -18343 -19622
rect -64167 -19681 -64043 -19680
rect -43363 -19717 -32282 -19656
rect -32220 -19717 -18343 -19656
rect -43363 -19727 -18343 -19717
rect -18238 -19727 -18124 -19622
rect -18017 -19727 -18003 -19620
rect -43363 -19728 -18003 -19727
rect -18352 -19741 -18003 -19728
rect -5606 -20120 -5520 -20045
rect -5606 -20172 -5590 -20120
rect -5533 -20172 -5520 -20120
rect -5606 -20240 -5520 -20172
rect 5825 -20218 5924 -20140
rect 5825 -20240 5842 -20218
rect -5606 -20256 5842 -20240
rect -5606 -20308 -5593 -20256
rect -5536 -20282 5842 -20256
rect 5908 -20282 5924 -20218
rect -5536 -20308 5924 -20282
rect -5606 -20326 5924 -20308
rect 5825 -20374 5924 -20326
rect 5408 -20448 5502 -20420
rect -3763 -20486 -3688 -20472
rect -18588 -20558 -18225 -20537
rect -3763 -20539 -3750 -20486
rect -3697 -20539 -3688 -20486
rect -3763 -20558 -3688 -20539
rect 5408 -20504 5431 -20448
rect 5486 -20504 5502 -20448
rect 5825 -20438 5842 -20374
rect 5908 -20438 5924 -20374
rect 6271 -20166 6362 -20125
rect 6271 -20226 6286 -20166
rect 6343 -20177 6362 -20166
rect 6343 -20217 17173 -20177
rect 6343 -20226 17089 -20217
rect 6271 -20277 17089 -20226
rect 6271 -20312 6362 -20277
rect 6271 -20372 6284 -20312
rect 6341 -20372 6362 -20312
rect 6271 -20388 6362 -20372
rect 17073 -20325 17089 -20277
rect 17158 -20325 17173 -20217
rect 5825 -20458 5924 -20438
rect 6988 -20452 7077 -20428
rect 5408 -20558 5502 -20504
rect 6988 -20505 7005 -20452
rect 7063 -20505 7077 -20452
rect 6988 -20558 7077 -20505
rect 17073 -20463 17173 -20325
rect -18588 -20559 -18336 -20558
rect -18588 -20651 -18560 -20559
rect -18468 -20651 -18336 -20559
rect -18588 -20652 -18336 -20651
rect -18242 -20575 7084 -20558
rect -18242 -20578 7004 -20575
rect -18242 -20594 5426 -20578
rect -18242 -20647 -3751 -20594
rect -3698 -20634 5426 -20594
rect 5481 -20628 7004 -20578
rect 7062 -20628 7084 -20575
rect 17073 -20571 17089 -20463
rect 17158 -20571 17173 -20463
rect 17073 -20592 17173 -20571
rect 5481 -20634 7084 -20628
rect -3698 -20647 7084 -20634
rect -18242 -20652 7084 -20647
rect -18588 -20667 -18225 -20652
rect -3763 -20659 -3688 -20652
rect 6988 -20657 7077 -20652
rect -34046 -20871 -33918 -20783
rect 5581 -20796 5675 -20766
rect -34046 -20965 -34026 -20871
rect -33939 -20965 -33918 -20871
rect -34046 -21044 -33918 -20965
rect -18881 -20839 -18754 -20809
rect -4056 -20839 -3941 -20836
rect 5581 -20839 5597 -20796
rect -18881 -20840 5597 -20839
rect -18881 -20932 -18864 -20840
rect -18772 -20851 5597 -20840
rect 5655 -20839 5675 -20796
rect 6527 -20839 6800 -20827
rect 5655 -20851 6800 -20839
rect -18772 -20925 -4037 -20851
rect -3963 -20855 6800 -20851
rect -3963 -20911 6573 -20855
rect 6637 -20862 6800 -20855
rect 6637 -20911 6714 -20862
rect -3963 -20918 6714 -20911
rect 6778 -20918 6800 -20862
rect -3963 -20925 6800 -20918
rect -18772 -20932 6800 -20925
rect -18881 -20933 6800 -20932
rect -19162 -21044 -19067 -21042
rect -34046 -21063 -19067 -21044
rect -34046 -21157 -34027 -21063
rect -33940 -21066 -19067 -21063
rect -33940 -21136 -19142 -21066
rect -19087 -21136 -19067 -21066
rect -33940 -21157 -19067 -21136
rect -34046 -21191 -19067 -21157
rect -18881 -21064 -18754 -20933
rect -18881 -21158 -18865 -21064
rect -18771 -21158 -18754 -21064
rect -18881 -21179 -18754 -21158
rect -4056 -21071 -3941 -20933
rect 5581 -20939 5675 -20933
rect 5581 -20994 5597 -20939
rect 5655 -20994 5675 -20939
rect 6527 -20965 6800 -20933
rect 5581 -21009 5675 -20994
rect -4056 -21145 -4037 -21071
rect -3963 -21145 -3941 -21071
rect -34046 -21192 -33918 -21191
rect -19162 -21229 -19067 -21191
rect -32299 -21307 -32200 -21286
rect -19162 -21299 -19140 -21229
rect -19085 -21299 -19067 -21229
rect -32299 -21308 -31744 -21307
rect -32299 -21380 -32282 -21308
rect -32210 -21380 -31744 -21308
rect -19162 -21333 -19067 -21299
rect -4056 -21262 -3941 -21145
rect -4056 -21263 -3776 -21262
rect -4056 -21335 -4036 -21263
rect -3964 -21335 -3776 -21263
rect -4056 -21336 -3776 -21335
rect -3641 -21336 -3566 -21262
rect -4056 -21372 -3941 -21336
rect -32299 -21381 -31744 -21380
rect -32299 -21494 -32200 -21381
rect -32299 -21568 -32283 -21494
rect -32209 -21568 -32200 -21494
rect -32299 -21579 -32200 -21568
rect -46038 -21619 -36670 -21586
rect -46038 -21621 -44610 -21619
rect -65698 -21648 -60846 -21627
rect -65698 -21655 -65545 -21648
rect -65698 -21752 -65679 -21655
rect -65617 -21745 -65545 -21655
rect -65483 -21657 -60846 -21648
rect -65483 -21745 -65410 -21657
rect -65617 -21752 -65410 -21745
rect -65698 -21754 -65410 -21752
rect -65348 -21754 -60846 -21657
rect -65698 -21848 -60846 -21754
rect -56384 -21673 -50667 -21645
rect -56384 -21677 -55004 -21673
rect -56384 -21749 -55288 -21677
rect -55226 -21749 -55155 -21677
rect -55093 -21745 -55004 -21677
rect -54942 -21745 -50667 -21673
rect -46038 -21688 -44932 -21621
rect -44878 -21622 -44610 -21621
rect -44878 -21688 -44775 -21622
rect -46038 -21689 -44775 -21688
rect -44721 -21686 -44610 -21622
rect -44556 -21686 -36670 -21619
rect -44721 -21689 -36670 -21686
rect -46038 -21705 -36670 -21689
rect -35822 -21644 -34295 -21619
rect 3432 -21627 13395 -21599
rect 3432 -21631 4996 -21627
rect -35822 -21649 -34377 -21644
rect -35822 -21652 -34539 -21649
rect -35822 -21721 -34695 -21652
rect -34637 -21718 -34539 -21652
rect -34481 -21713 -34377 -21649
rect -34319 -21713 -34295 -21644
rect -34481 -21718 -34295 -21713
rect -34637 -21721 -34295 -21718
rect -35822 -21734 -34295 -21721
rect -24737 -21674 -15153 -21631
rect -55093 -21749 -50667 -21745
rect -56384 -21762 -50667 -21749
rect -65698 -21945 -65683 -21848
rect -65621 -21945 -65535 -21848
rect -65473 -21851 -60846 -21848
rect -65473 -21945 -65388 -21851
rect -65698 -21948 -65388 -21945
rect -65326 -21948 -60846 -21851
rect -50784 -21875 -50667 -21762
rect -24737 -21766 -23388 -21674
rect -23320 -21679 -15153 -21674
rect -23320 -21766 -23233 -21679
rect -24737 -21771 -23233 -21766
rect -23165 -21680 -15153 -21679
rect -23165 -21771 -23086 -21680
rect -24737 -21772 -23086 -21771
rect -23018 -21772 -15153 -21680
rect -24737 -21786 -15153 -21772
rect -10762 -21670 -6736 -21641
rect -10762 -21677 -6828 -21670
rect -10762 -21679 -6975 -21677
rect -10762 -21759 -7139 -21679
rect -7079 -21757 -6975 -21679
rect -6915 -21750 -6828 -21677
rect -6768 -21750 -6736 -21670
rect 3432 -21726 4842 -21631
rect 4915 -21722 4996 -21631
rect 5069 -21629 13395 -21627
rect 5069 -21722 5143 -21629
rect 4915 -21724 5143 -21722
rect 5216 -21724 13395 -21629
rect 24943 -21624 34979 -21593
rect 24943 -21627 26307 -21624
rect 4915 -21726 13395 -21724
rect 3432 -21748 13395 -21726
rect 14233 -21704 20470 -21664
rect 14233 -21705 15612 -21704
rect -6915 -21757 -6736 -21750
rect -7079 -21759 -6736 -21757
rect -10762 -21774 -6736 -21759
rect 14233 -21777 15332 -21705
rect 15388 -21708 15612 -21705
rect 15388 -21777 15472 -21708
rect 14233 -21780 15472 -21777
rect 15528 -21776 15612 -21708
rect 15668 -21776 20470 -21704
rect 24943 -21708 26028 -21627
rect 26084 -21708 26172 -21627
rect 26228 -21705 26307 -21627
rect 26363 -21705 34979 -21624
rect 26228 -21708 34979 -21705
rect 24943 -21722 34979 -21708
rect 15528 -21780 20470 -21776
rect 14233 -21797 20470 -21780
rect -31976 -21859 -31865 -21813
rect -65698 -21960 -60846 -21948
rect -31976 -21922 -31954 -21859
rect -31889 -21922 -31865 -21859
rect -31976 -22008 -31865 -21922
rect -3767 -21882 -3670 -21861
rect -3767 -21940 -3754 -21882
rect -3696 -21940 -3670 -21882
rect 20337 -21884 20470 -21797
rect -3767 -21963 -3670 -21940
rect -3847 -21996 -3595 -21963
rect -31976 -22031 -31654 -22008
rect -31976 -22094 -31959 -22031
rect -31894 -22094 -31654 -22031
rect -3847 -22054 -3756 -21996
rect -3698 -22054 -3595 -21996
rect -3847 -22074 -3595 -22054
rect -3767 -22086 -3670 -22074
rect -31976 -22119 -31654 -22094
rect -68464 -22562 -66006 -22517
rect -55937 -22527 -53703 -22501
rect -55937 -22528 -55630 -22527
rect -68464 -22611 -63952 -22562
rect -68464 -22614 -66231 -22611
rect -68464 -22665 -66363 -22614
rect -66387 -22677 -66363 -22665
rect -66303 -22674 -66231 -22614
rect -66171 -22614 -63952 -22611
rect -66171 -22674 -66097 -22614
rect -66303 -22677 -66097 -22674
rect -66037 -22677 -63952 -22614
rect -55937 -22631 -55917 -22528
rect -55837 -22529 -55630 -22528
rect -55837 -22631 -55769 -22529
rect -55937 -22632 -55769 -22631
rect -55689 -22630 -55630 -22529
rect -55550 -22630 -53703 -22527
rect -55689 -22632 -53703 -22630
rect -55937 -22651 -53703 -22632
rect -45768 -22605 -43338 -22535
rect -45768 -22608 -45464 -22605
rect -45768 -22615 -45624 -22608
rect -66387 -22712 -63952 -22677
rect -45768 -22671 -45752 -22615
rect -45700 -22664 -45624 -22615
rect -45572 -22661 -45464 -22608
rect -45412 -22661 -43338 -22605
rect -45572 -22664 -43338 -22661
rect -45700 -22671 -43338 -22664
rect -45768 -22685 -43338 -22671
rect -24192 -22593 -18456 -22564
rect 14632 -22571 17358 -22516
rect 14632 -22578 14765 -22571
rect -24192 -22600 -23895 -22593
rect -24192 -22603 -24039 -22600
rect -24192 -22690 -24172 -22603
rect -24112 -22687 -24039 -22603
rect -23979 -22680 -23895 -22600
rect -23835 -22680 -18456 -22593
rect -23979 -22687 -18456 -22680
rect -24112 -22690 -18456 -22687
rect -24192 -22714 -18456 -22690
rect 4054 -22657 6723 -22589
rect 4054 -22659 4361 -22657
rect 4054 -22662 4232 -22659
rect 4054 -22718 4094 -22662
rect 4146 -22715 4232 -22662
rect 4284 -22713 4361 -22659
rect 4413 -22713 6723 -22657
rect 14632 -22634 14652 -22578
rect 14704 -22627 14765 -22578
rect 14817 -22627 14888 -22571
rect 14940 -22627 17358 -22571
rect 14704 -22634 17358 -22627
rect 14632 -22666 17358 -22634
rect 25328 -22616 28494 -22551
rect 25328 -22619 25485 -22616
rect 25328 -22682 25353 -22619
rect 25413 -22679 25485 -22619
rect 25545 -22619 28494 -22616
rect 25545 -22679 25619 -22619
rect 25413 -22682 25619 -22679
rect 25679 -22682 28494 -22619
rect 25328 -22701 28494 -22682
rect 4284 -22715 6723 -22713
rect 4146 -22718 6723 -22715
rect 4054 -22739 6723 -22718
rect -53204 -22980 -53117 -22959
rect -63396 -23012 -63309 -22991
rect -63396 -23068 -63383 -23012
rect -63327 -23068 -63309 -23012
rect -63396 -23123 -63309 -23068
rect -63396 -23179 -63387 -23123
rect -63331 -23179 -63309 -23123
rect -53204 -23036 -53191 -22980
rect -53135 -23036 -53117 -22980
rect -53204 -23091 -53117 -23036
rect -53204 -23147 -53195 -23091
rect -53139 -23147 -53117 -23091
rect -53204 -23162 -53117 -23147
rect -42813 -22989 -42726 -22968
rect -42813 -23045 -42800 -22989
rect -42744 -23045 -42726 -22989
rect -42813 -23100 -42726 -23045
rect -42813 -23156 -42804 -23100
rect -42748 -23156 -42726 -23100
rect -42813 -23171 -42726 -23156
rect -17905 -23001 -17818 -22980
rect -17905 -23057 -17892 -23001
rect -17836 -23057 -17818 -23001
rect 14642 -23006 14999 -22986
rect 14642 -23013 14771 -23006
rect 14642 -23018 14658 -23013
rect -17905 -23112 -17818 -23057
rect 14626 -23069 14658 -23018
rect 14710 -23062 14771 -23013
rect 14823 -23062 14894 -23006
rect 14946 -23018 14999 -23006
rect 14946 -23062 17563 -23018
rect 25338 -23042 25706 -23029
rect 25338 -23045 25486 -23042
rect 25338 -23053 25354 -23045
rect 14710 -23069 17563 -23062
rect 4074 -23091 4446 -23069
rect -17905 -23168 -17896 -23112
rect -17840 -23168 -17818 -23112
rect -63396 -23194 -63309 -23179
rect -17905 -23183 -17818 -23168
rect 4043 -23094 6678 -23091
rect 4043 -23096 4360 -23094
rect 4043 -23099 4231 -23096
rect 4043 -23155 4093 -23099
rect 4145 -23152 4231 -23099
rect 4283 -23150 4360 -23096
rect 4412 -23150 6678 -23094
rect 14626 -23100 17563 -23069
rect 25325 -23108 25354 -23053
rect 25414 -23105 25486 -23045
rect 25546 -23045 25706 -23042
rect 25546 -23105 25620 -23045
rect 25414 -23108 25620 -23105
rect 25680 -23053 25706 -23045
rect 25680 -23108 28329 -23053
rect 25325 -23135 28329 -23108
rect 4283 -23152 6678 -23150
rect 4145 -23155 6678 -23152
rect 4043 -23173 6678 -23155
rect -68544 -23421 -68408 -23396
rect -68544 -23497 -68519 -23421
rect -68436 -23497 -68408 -23421
rect -68544 -23522 -68408 -23497
rect -66896 -23417 -66736 -23397
rect -66896 -23497 -66855 -23417
rect -66759 -23497 -66736 -23417
rect -66896 -23523 -66736 -23497
rect 17073 -23782 17172 -23765
rect 5823 -23940 5925 -23869
rect -68274 -24173 -65295 -24025
rect -64374 -24026 -64283 -23957
rect -64374 -24084 -64355 -24026
rect -64297 -24033 -64283 -24026
rect -54239 -23972 -54158 -23962
rect -54239 -24001 -53818 -23972
rect -64297 -24084 -63952 -24033
rect -64374 -24107 -63952 -24084
rect -54239 -24059 -54223 -24001
rect -54171 -24046 -53818 -24001
rect -19162 -23981 -19070 -23949
rect -43805 -24018 -43377 -24006
rect -54171 -24059 -54157 -24046
rect -65607 -25337 -65459 -24173
rect -64374 -24207 -64283 -24107
rect -64374 -24265 -64361 -24207
rect -64303 -24265 -64283 -24207
rect -54239 -24171 -54157 -24059
rect -54239 -24229 -54228 -24171
rect -54176 -24229 -54157 -24171
rect -54239 -24240 -54157 -24229
rect -43805 -24082 -43793 -24018
rect -43740 -24080 -43377 -24018
rect -19162 -24048 -19149 -23981
rect -19082 -24035 -19070 -23981
rect 5823 -24003 5833 -23940
rect 5909 -24003 5925 -23940
rect -19082 -24048 -18315 -24035
rect -43740 -24082 -43731 -24080
rect -43805 -24200 -43731 -24082
rect -19162 -24109 -18315 -24048
rect 5823 -24060 5925 -24003
rect 17073 -23870 17087 -23782
rect 17153 -23870 17172 -23782
rect 17073 -23957 17172 -23870
rect 17073 -24045 17086 -23957
rect 17152 -23987 17172 -23957
rect 17152 -24045 17284 -23987
rect 26027 -24007 26395 -23994
rect 26027 -24010 26175 -24007
rect 26027 -24022 26043 -24010
rect 5823 -24097 6587 -24060
rect 17073 -24061 17284 -24045
rect 26009 -24073 26043 -24022
rect 26103 -24070 26175 -24010
rect 26235 -24010 26395 -24007
rect 26235 -24070 26309 -24010
rect 26103 -24073 26309 -24070
rect 26369 -24022 26395 -24010
rect 26369 -24073 28318 -24022
rect 26009 -24096 28318 -24073
rect -64374 -24279 -64283 -24265
rect -43805 -24264 -43796 -24200
rect -43743 -24264 -43731 -24200
rect -35395 -24179 -31967 -24166
rect -35395 -24235 -35377 -24179
rect -35325 -24180 -31967 -24179
rect -35325 -24181 -35104 -24180
rect -35325 -24235 -35251 -24181
rect -35395 -24237 -35251 -24235
rect -35199 -24236 -35104 -24181
rect -35052 -24236 -31967 -24180
rect -35199 -24237 -31967 -24236
rect -35395 -24248 -31967 -24237
rect -19162 -24171 -19070 -24109
rect -19162 -24238 -19154 -24171
rect -19087 -24238 -19070 -24171
rect -7918 -24134 -3816 -24121
rect -7918 -24190 -7900 -24134
rect -7848 -24135 -7663 -24134
rect -7848 -24190 -7785 -24135
rect -7918 -24191 -7785 -24190
rect -7733 -24190 -7663 -24135
rect -7611 -24190 -3816 -24134
rect 5823 -24160 5834 -24097
rect 5910 -24134 6587 -24097
rect 5910 -24160 5925 -24134
rect 5823 -24171 5925 -24160
rect -7733 -24191 -3816 -24190
rect -7918 -24203 -3816 -24191
rect -19162 -24251 -19070 -24238
rect -43805 -24281 -43731 -24264
rect -18293 -24854 -18140 -24841
rect -53554 -24909 -53409 -24882
rect -63739 -24952 -63652 -24931
rect -63739 -25008 -63726 -24952
rect -63670 -25008 -63652 -24952
rect -63739 -25063 -63652 -25008
rect -63739 -25119 -63730 -25063
rect -63674 -25119 -63652 -25063
rect -63739 -25127 -63652 -25119
rect -53554 -24971 -53526 -24909
rect -53467 -24971 -53409 -24909
rect -53554 -25047 -53409 -24971
rect -18293 -24936 -18255 -24854
rect -18173 -24936 -18140 -24854
rect -53554 -25109 -53543 -25047
rect -53484 -25109 -53409 -25047
rect -53554 -25124 -53409 -25109
rect -43355 -25037 -43028 -24974
rect -43355 -25050 -43186 -25037
rect -43355 -25117 -43341 -25050
rect -43267 -25104 -43186 -25050
rect -43112 -25104 -43028 -25037
rect -43267 -25117 -43028 -25104
rect -43355 -25126 -43028 -25117
rect -18293 -25019 -18140 -24936
rect -18293 -25101 -18255 -25019
rect -18173 -25101 -18140 -25019
rect 6656 -24974 6999 -24908
rect 6656 -24990 6880 -24974
rect 6656 -25067 6666 -24990
rect 6734 -25051 6880 -24990
rect 6948 -25051 6999 -24974
rect 6734 -25067 6999 -25051
rect -18293 -25126 -18140 -25101
rect -55289 -25280 -53594 -25276
rect -55289 -25284 -55272 -25280
rect -65695 -25368 -63698 -25337
rect -65695 -25371 -65540 -25368
rect -65695 -25434 -65672 -25371
rect -65612 -25431 -65540 -25371
rect -65480 -25371 -63698 -25368
rect -65480 -25431 -65406 -25371
rect -65612 -25434 -65406 -25431
rect -65346 -25434 -63698 -25371
rect -56785 -25383 -55272 -25284
rect -55192 -25281 -54983 -25280
rect -55192 -25383 -55120 -25281
rect -56785 -25384 -55120 -25383
rect -55040 -25383 -54983 -25281
rect -54903 -25383 -53594 -25280
rect -46596 -25310 -44565 -25220
rect -30674 -25223 -30628 -25131
rect -2508 -25191 -2462 -25095
rect 6656 -25121 6999 -25067
rect 17320 -24952 17731 -24878
rect 17320 -24962 17593 -24952
rect 17320 -25055 17338 -24962
rect 17421 -25045 17593 -24962
rect 17676 -25045 17731 -24952
rect 17421 -25055 17731 -25045
rect 17320 -25100 17731 -25055
rect 28308 -24912 28480 -24908
rect 28308 -24969 28407 -24912
rect 28463 -24969 28480 -24912
rect 28308 -25015 28480 -24969
rect 28308 -25072 28314 -25015
rect 28370 -25072 28480 -25015
rect 28308 -25084 28480 -25072
rect -36214 -25271 -34292 -25254
rect -36214 -25273 -34430 -25271
rect -36214 -25274 -34558 -25273
rect -46596 -25320 -43209 -25310
rect -55040 -25384 -53594 -25383
rect -55289 -25393 -53594 -25384
rect -44944 -25352 -43209 -25320
rect -44944 -25354 -44693 -25352
rect -44944 -25360 -44810 -25354
rect -44944 -25416 -44926 -25360
rect -44874 -25410 -44810 -25360
rect -44758 -25408 -44693 -25354
rect -44641 -25408 -43209 -25352
rect -36214 -25343 -34692 -25274
rect -34634 -25342 -34558 -25274
rect -34500 -25340 -34430 -25273
rect -34372 -25340 -34292 -25271
rect -11302 -25305 -6737 -25283
rect -11302 -25308 -6840 -25305
rect -34500 -25342 -34292 -25340
rect -34634 -25343 -34292 -25342
rect -36214 -25354 -34292 -25343
rect -23401 -25351 -18356 -25339
rect -44758 -25410 -43209 -25408
rect -44874 -25416 -43209 -25410
rect -44944 -25427 -43209 -25416
rect -23401 -25358 -23106 -25351
rect -23401 -25361 -23250 -25358
rect -65695 -25454 -63698 -25434
rect -23401 -25448 -23383 -25361
rect -23323 -25445 -23250 -25361
rect -23190 -25438 -23106 -25358
rect -23046 -25438 -18356 -25351
rect -11302 -25370 -7135 -25308
rect -7078 -25310 -6840 -25308
rect -7078 -25370 -6999 -25310
rect -11302 -25372 -6999 -25370
rect -6942 -25367 -6840 -25310
rect -6783 -25367 -6737 -25305
rect 15324 -25311 17459 -25291
rect 13822 -25325 17459 -25311
rect 13822 -25336 15457 -25325
rect -6942 -25372 -6737 -25367
rect -11302 -25383 -6737 -25372
rect -23190 -25445 -18356 -25438
rect -23323 -25448 -18356 -25445
rect -23401 -25456 -18356 -25448
rect 4832 -25402 6723 -25364
rect 4832 -25406 5117 -25402
rect 4832 -25462 4859 -25406
rect 4911 -25407 5117 -25406
rect 4911 -25462 5002 -25407
rect 4832 -25463 5002 -25462
rect 5054 -25458 5117 -25407
rect 5169 -25458 6723 -25402
rect 13822 -25392 15341 -25336
rect 15393 -25381 15457 -25336
rect 15509 -25330 17459 -25325
rect 15509 -25381 15582 -25330
rect 15393 -25386 15582 -25381
rect 15634 -25386 17459 -25330
rect 24530 -25326 26294 -25235
rect 24530 -25335 28186 -25326
rect 15393 -25392 17459 -25386
rect 13822 -25408 17459 -25392
rect 26013 -25352 28186 -25335
rect 26013 -25355 26177 -25352
rect 13822 -25411 15489 -25408
rect 26013 -25418 26045 -25355
rect 26105 -25415 26177 -25355
rect 26237 -25355 28186 -25352
rect 26237 -25415 26311 -25355
rect 26105 -25418 26311 -25415
rect 26371 -25418 28186 -25355
rect 26013 -25443 28186 -25418
rect 5054 -25463 6723 -25458
rect 4832 -25481 6723 -25463
rect -66934 -25615 -65974 -25570
rect -66934 -25618 -66204 -25615
rect -66934 -25702 -66369 -25618
rect -66299 -25699 -66204 -25618
rect -66134 -25699 -66063 -25615
rect -65993 -25699 -65974 -25615
rect -66299 -25702 -65974 -25699
rect -66934 -25717 -65974 -25702
rect -64137 -25692 -64058 -25669
rect -64137 -25758 -64119 -25692
rect -64066 -25758 -64058 -25692
rect 27808 -25702 27908 -25686
rect -64137 -25760 -64058 -25758
rect -64137 -25818 -63922 -25760
rect -64137 -25884 -64127 -25818
rect -64074 -25828 -63922 -25818
rect 6406 -25772 6508 -25749
rect -64074 -25884 -64058 -25828
rect -64137 -25903 -64058 -25884
rect 6406 -25848 6419 -25772
rect 6495 -25787 6508 -25772
rect 27808 -25770 27825 -25702
rect 27893 -25749 27908 -25702
rect 27893 -25770 28110 -25749
rect 6495 -25848 6780 -25787
rect 6406 -25854 6424 -25848
rect 6490 -25854 6780 -25848
rect 6406 -25855 6780 -25854
rect 27808 -25817 28110 -25770
rect 6406 -25962 6508 -25855
rect 27808 -25877 27908 -25817
rect 27808 -25943 27826 -25877
rect 27892 -25943 27908 -25877
rect 27808 -25961 27908 -25943
rect -54014 -26041 -53903 -26026
rect 6406 -26030 6423 -25962
rect 6491 -26030 6508 -25962
rect 6406 -26040 6508 -26030
rect -54014 -26118 -53999 -26041
rect -53922 -26118 -53903 -26041
rect -4607 -26064 -4503 -26043
rect -63882 -26184 -63802 -26168
rect -63882 -26238 -63865 -26184
rect -63812 -26238 -63802 -26184
rect -63882 -26287 -63802 -26238
rect -54014 -26226 -53903 -26118
rect -33384 -26115 -33297 -26095
rect -33384 -26172 -33372 -26115
rect -33315 -26172 -33297 -26115
rect -54014 -26227 -53672 -26226
rect -63882 -26292 -63687 -26287
rect -63882 -26347 -63860 -26292
rect -63807 -26347 -63687 -26292
rect -61668 -26327 -60883 -26255
rect -54014 -26302 -53999 -26227
rect -53924 -26302 -53672 -26227
rect -51484 -26266 -50630 -26194
rect -54014 -26303 -53672 -26302
rect -43625 -26282 -43314 -26260
rect -54014 -26325 -53903 -26303
rect -63882 -26364 -63687 -26347
rect -43625 -26338 -43616 -26282
rect -43555 -26337 -43314 -26282
rect -41119 -26300 -40184 -26228
rect -33384 -26247 -33297 -26172
rect -18879 -26115 -18765 -26094
rect -18879 -26192 -18858 -26115
rect -18781 -26192 -18765 -26115
rect -33384 -26248 -31908 -26247
rect -33384 -26303 -33366 -26248
rect -33311 -26303 -31908 -26248
rect -33384 -26304 -31908 -26303
rect -18879 -26289 -18765 -26192
rect -4607 -26121 -4581 -26064
rect -4524 -26121 -4503 -26064
rect -4607 -26202 -4503 -26121
rect 28095 -26122 28222 -26099
rect 28095 -26197 28123 -26122
rect 28198 -26197 28222 -26122
rect -4607 -26203 -3758 -26202
rect -18879 -26290 -18360 -26289
rect -33384 -26313 -33297 -26304
rect -43555 -26338 -43548 -26337
rect -43625 -26406 -43548 -26338
rect -18879 -26365 -18858 -26290
rect -18783 -26365 -18360 -26290
rect -16192 -26329 -15348 -26257
rect -4607 -26258 -4581 -26203
rect -4526 -26258 -3758 -26203
rect -4607 -26259 -3758 -26258
rect -4607 -26275 -4503 -26259
rect 6696 -26315 6813 -26290
rect -18879 -26366 -18360 -26365
rect -18879 -26393 -18765 -26366
rect 6696 -26390 6710 -26315
rect 6785 -26390 6813 -26315
rect 8937 -26354 9745 -26282
rect -68616 -26477 -68488 -26457
rect -68616 -26561 -68598 -26477
rect -68504 -26561 -68488 -26477
rect -68616 -26585 -68488 -26561
rect -66964 -26469 -66815 -26427
rect -66964 -26559 -66935 -26469
rect -66854 -26559 -66815 -26469
rect -43625 -26462 -43618 -26406
rect -43557 -26462 -43548 -26406
rect -43625 -26476 -43548 -26462
rect 6696 -26481 6813 -26390
rect -66964 -26588 -66815 -26559
rect -7147 -26567 -3667 -26536
rect -34696 -26614 -31783 -26581
rect -34696 -26619 -34407 -26614
rect -34696 -26627 -34552 -26619
rect -34696 -26683 -34684 -26627
rect -34632 -26675 -34552 -26627
rect -34500 -26670 -34407 -26619
rect -34355 -26670 -31783 -26614
rect -34500 -26675 -31783 -26670
rect -34632 -26683 -31783 -26675
rect -34696 -26694 -31783 -26683
rect -24727 -26606 -18360 -26568
rect -34611 -26757 -34464 -26694
rect -24727 -26698 -23390 -26606
rect -23322 -26613 -18360 -26606
rect -23322 -26698 -23225 -26613
rect -24727 -26705 -23225 -26698
rect -23157 -26705 -23080 -26613
rect -23012 -26705 -18360 -26613
rect -7147 -26572 -6866 -26567
rect -7147 -26581 -6996 -26572
rect -7147 -26637 -7135 -26581
rect -7083 -26628 -6996 -26581
rect -6944 -26623 -6866 -26572
rect -6814 -26623 -3667 -26567
rect -6944 -26628 -3667 -26623
rect -7083 -26637 -3667 -26628
rect -7147 -26649 -3667 -26637
rect 3441 -26564 5230 -26530
rect 3441 -26565 4985 -26564
rect -24727 -26718 -18360 -26705
rect -34611 -26826 -34568 -26757
rect -34510 -26826 -34464 -26757
rect -34611 -26917 -34464 -26826
rect -53346 -26949 -34464 -26917
rect -53346 -26968 -34568 -26949
rect -53346 -26969 -44792 -26968
rect -53346 -26999 -44934 -26969
rect -63580 -27046 -44934 -26999
rect -63580 -27058 -54971 -27046
rect -63580 -27079 -55286 -27058
rect -66972 -27116 -55286 -27079
rect -66972 -27118 -65522 -27116
rect -66972 -27209 -65682 -27118
rect -65616 -27207 -65522 -27118
rect -65456 -27118 -55286 -27116
rect -65456 -27207 -65380 -27118
rect -65616 -27209 -65380 -27207
rect -65314 -27130 -55286 -27118
rect -55224 -27130 -55145 -27058
rect -55083 -27118 -54971 -27058
rect -54909 -27047 -44934 -27046
rect -44876 -27046 -44792 -26969
rect -44734 -26971 -34568 -26968
rect -44734 -27046 -44625 -26971
rect -44876 -27047 -44625 -27046
rect -54909 -27049 -44625 -27047
rect -44567 -27018 -34568 -26971
rect -34510 -27018 -34464 -26949
rect -44567 -27049 -34464 -27018
rect -54909 -27064 -34464 -27049
rect -33055 -26862 -32958 -26838
rect -33055 -26919 -33031 -26862
rect -32973 -26884 -32958 -26862
rect -32973 -26919 -31776 -26884
rect -33055 -26978 -31776 -26919
rect -33055 -26984 -32958 -26978
rect -33055 -27041 -33034 -26984
rect -32976 -27041 -32958 -26984
rect -54909 -27118 -52917 -27064
rect -33055 -27079 -32958 -27041
rect -18510 -27010 -18360 -26718
rect -7049 -27010 -6899 -26649
rect 3441 -26658 4840 -26565
rect 4913 -26657 4985 -26565
rect 5058 -26567 5230 -26564
rect 5058 -26657 5131 -26567
rect 4913 -26658 5131 -26657
rect 3441 -26660 5131 -26658
rect 5204 -26660 5230 -26567
rect 6696 -26558 6709 -26481
rect 6786 -26558 6813 -26481
rect 6696 -26576 6813 -26558
rect 3441 -26676 5230 -26660
rect -4318 -26839 -4069 -26828
rect -4318 -26857 -3697 -26839
rect -4318 -26860 -4151 -26857
rect -4318 -26915 -4282 -26860
rect -4227 -26912 -4151 -26860
rect -4096 -26912 -3697 -26857
rect -4227 -26915 -3697 -26912
rect -4318 -26933 -3697 -26915
rect -4318 -26957 -4069 -26933
rect 13880 -26949 15727 -26900
rect 13880 -26951 15480 -26949
rect -55083 -27130 -52917 -27118
rect -65314 -27146 -52917 -27130
rect -65314 -27209 -63433 -27146
rect -18510 -27160 -6899 -27010
rect 13880 -27044 15336 -26951
rect 15401 -27042 15480 -26951
rect 15545 -26951 15727 -26949
rect 15545 -27042 15622 -26951
rect 15401 -27044 15622 -27042
rect 15687 -27044 15727 -26951
rect 6687 -27136 6814 -27079
rect 13880 -27082 15727 -27044
rect -66972 -27226 -63433 -27209
rect 6687 -27221 6707 -27136
rect 6785 -27221 6814 -27136
rect 6687 -27289 6814 -27221
rect 17425 -27289 17550 -26224
rect 19646 -26281 20507 -26209
rect 28095 -26276 28222 -26197
rect 28095 -26277 28321 -26276
rect 28095 -26352 28119 -26277
rect 28195 -26352 28321 -26277
rect 30370 -26316 31178 -26244
rect 28095 -26353 28321 -26352
rect 28095 -26389 28222 -26353
rect 6684 -27296 17550 -27289
rect 6684 -27381 6709 -27296
rect 6787 -27381 17550 -27296
rect 6684 -27414 17550 -27381
rect 6687 -27416 6814 -27414
rect 6392 -27521 6516 -27469
rect 6392 -27601 6418 -27521
rect 6498 -27601 6516 -27521
rect 6392 -27659 6516 -27601
rect 17804 -27659 17929 -26728
rect 24590 -26878 27930 -26824
rect 24590 -26979 26027 -26878
rect 26103 -26880 27930 -26878
rect 26103 -26882 26333 -26880
rect 26103 -26979 26184 -26882
rect 24590 -26983 26184 -26979
rect 26260 -26981 26333 -26882
rect 26409 -26981 27930 -26880
rect 26260 -26983 27930 -26981
rect 24590 -27003 27930 -26983
rect 27751 -27021 27930 -27003
rect 28854 -27021 35408 -27016
rect 27751 -27200 35408 -27021
rect 6387 -27678 17929 -27659
rect 6387 -27758 6415 -27678
rect 6495 -27758 17929 -27678
rect -43815 -27798 -43727 -27763
rect 6387 -27784 17929 -27758
rect 6392 -27789 6516 -27784
rect -43815 -27856 -43801 -27798
rect -43741 -27856 -43727 -27798
rect -43815 -27921 -43727 -27856
rect -19162 -27877 -19070 -27858
rect -43815 -27936 -43021 -27921
rect -43815 -27994 -43803 -27936
rect -43743 -27994 -43021 -27936
rect -43815 -28009 -43021 -27994
rect -54240 -28060 -54157 -28019
rect -54240 -28121 -54225 -28060
rect -54170 -28121 -54157 -28060
rect -54240 -28212 -54157 -28121
rect -43901 -28172 -43816 -28151
rect -43901 -28212 -43887 -28172
rect -54241 -28224 -43887 -28212
rect -54241 -28285 -54229 -28224
rect -54174 -28233 -43887 -28224
rect -43827 -28233 -43816 -28172
rect -54174 -28285 -43816 -28233
rect -54241 -28297 -43816 -28285
rect -43901 -28337 -43816 -28297
rect -43901 -28398 -43891 -28337
rect -43831 -28398 -43816 -28337
rect -43109 -28291 -43021 -28009
rect -19162 -27939 -19151 -27877
rect -19083 -27939 -19070 -27877
rect -19162 -28027 -19070 -27939
rect -4591 -28027 -4476 -27977
rect -19163 -28030 -4476 -28027
rect -19163 -28043 -4570 -28030
rect -19163 -28105 -19151 -28043
rect -19083 -28105 -4570 -28043
rect -19163 -28106 -4570 -28105
rect -4499 -28106 -4476 -28030
rect -19163 -28118 -4476 -28106
rect -19401 -28215 -19313 -28180
rect -19401 -28274 -19388 -28215
rect -19326 -28274 -19313 -28215
rect -19401 -28291 -19313 -28274
rect -43109 -28379 -19313 -28291
rect -4591 -28255 -4476 -28118
rect -4591 -28331 -4569 -28255
rect -4498 -28331 -4476 -28255
rect -4591 -28358 -4476 -28331
rect -43901 -28408 -43816 -28398
rect -19401 -28380 -19313 -28379
rect -64376 -28449 -64281 -28425
rect -64376 -28505 -64357 -28449
rect -64291 -28505 -64281 -28449
rect -19401 -28439 -19391 -28380
rect -19329 -28439 -19313 -28380
rect -19401 -28451 -19313 -28439
rect -64376 -28585 -64281 -28505
rect -43637 -28498 -43528 -28464
rect -43637 -28562 -43607 -28498
rect -54131 -28564 -43607 -28562
rect -43551 -28562 -43528 -28498
rect -18982 -28505 -18873 -28486
rect -18982 -28562 -18955 -28505
rect -43551 -28564 -18955 -28562
rect -54131 -28580 -18955 -28564
rect -18890 -28580 -18873 -28505
rect -64377 -28608 -54326 -28585
rect -64377 -28664 -64364 -28608
rect -64298 -28621 -54326 -28608
rect -64298 -28664 -54400 -28621
rect -64377 -28676 -54400 -28664
rect -54342 -28676 -54326 -28621
rect -64377 -28680 -54326 -28676
rect -54421 -28784 -54326 -28680
rect -54421 -28839 -54406 -28784
rect -54348 -28839 -54326 -28784
rect -54421 -28857 -54326 -28839
rect -54131 -28586 -18873 -28580
rect -54131 -28596 -32650 -28586
rect -54131 -28654 -54099 -28596
rect -54037 -28651 -32650 -28596
rect -54037 -28654 -43616 -28651
rect -54131 -28671 -43616 -28654
rect -54131 -28751 -54022 -28671
rect -43637 -28717 -43616 -28671
rect -43560 -28652 -32650 -28651
rect -32581 -28652 -18873 -28586
rect -43560 -28671 -18873 -28652
rect -43560 -28717 -43528 -28671
rect -43637 -28744 -43528 -28717
rect -32665 -28706 -32568 -28671
rect -54131 -28809 -54098 -28751
rect -54036 -28809 -54022 -28751
rect -32665 -28772 -32652 -28706
rect -32583 -28772 -32568 -28706
rect -32665 -28788 -32568 -28772
rect -18982 -28699 -18873 -28671
rect -18982 -28774 -18961 -28699
rect -18896 -28774 -18873 -28699
rect -18982 -28802 -18873 -28774
rect -54131 -28866 -54022 -28809
rect -53845 -28848 -32851 -28830
rect -53845 -28852 -32932 -28848
rect -66963 -29010 -56216 -28886
rect -66963 -29093 -56389 -29010
rect -56423 -29119 -56389 -29093
rect -56253 -29119 -56216 -29010
rect -56423 -29259 -56216 -29119
rect -53845 -28941 -53823 -28852
rect -53745 -28909 -32932 -28852
rect -32873 -28909 -32851 -28848
rect -53745 -28920 -32851 -28909
rect -53745 -28941 -43332 -28920
rect -53845 -28942 -43332 -28941
rect -53845 -29057 -53733 -28942
rect -53845 -29146 -53819 -29057
rect -53741 -29146 -53733 -29057
rect -53845 -29203 -53733 -29146
rect -43361 -29004 -43332 -28942
rect -43262 -28924 -32851 -28920
rect -43262 -28942 -18590 -28924
rect -43262 -29004 -43249 -28942
rect -43361 -29076 -43249 -29004
rect -32963 -28964 -18590 -28942
rect -32963 -29025 -32939 -28964
rect -32880 -28987 -18590 -28964
rect -32880 -29025 -18667 -28987
rect -32963 -29036 -18667 -29025
rect -32953 -29037 -32858 -29036
rect -43361 -29160 -43340 -29076
rect -43270 -29160 -43249 -29076
rect -43361 -29181 -43249 -29160
rect -18702 -29054 -18667 -29036
rect -18602 -29054 -18590 -28987
rect -18702 -29175 -18590 -29054
rect -56423 -29368 -56397 -29259
rect -56261 -29368 -56216 -29259
rect -18702 -29242 -18681 -29175
rect -18616 -29242 -18590 -29175
rect -18702 -29271 -18590 -29242
rect -56423 -29406 -56216 -29368
rect -32675 -29432 -32550 -29396
rect -32675 -29506 -32649 -29432
rect -32575 -29506 -32550 -29432
rect -32675 -29605 -32550 -29506
rect -32675 -29606 -31410 -29605
rect -32675 -29678 -32648 -29606
rect -32576 -29678 -31410 -29606
rect 6690 -29611 6791 -29596
rect -32675 -29679 -31410 -29678
rect -32675 -29697 -32550 -29679
rect -10942 -29684 2593 -29652
rect -10942 -29685 -6879 -29684
rect -10942 -29686 -7009 -29685
rect -55307 -29739 -50573 -29727
rect -55307 -29745 -55142 -29739
rect -55307 -29823 -55284 -29745
rect -55223 -29817 -55142 -29745
rect -55081 -29742 -50573 -29739
rect -55081 -29817 -54974 -29742
rect -55223 -29820 -54974 -29817
rect -54913 -29820 -50573 -29742
rect -55223 -29823 -50573 -29820
rect -55307 -29832 -50573 -29823
rect -50663 -29834 -50573 -29832
rect -46153 -29752 -36389 -29725
rect -46153 -29756 -44626 -29752
rect -46153 -29827 -44931 -29756
rect -44876 -29757 -44626 -29756
rect -44876 -29827 -44788 -29757
rect -46153 -29828 -44788 -29827
rect -44733 -29823 -44626 -29757
rect -44571 -29823 -36389 -29752
rect -44733 -29828 -36389 -29823
rect -46153 -29843 -36389 -29828
rect -35616 -29733 -34304 -29703
rect -35616 -29734 -34424 -29733
rect -35616 -29738 -34562 -29734
rect -35616 -29818 -34684 -29738
rect -34627 -29814 -34562 -29738
rect -34505 -29813 -34424 -29734
rect -34367 -29813 -34304 -29733
rect -10942 -29783 -7135 -29686
rect -7069 -29782 -7009 -29686
rect -6943 -29781 -6879 -29685
rect -6813 -29781 2593 -29684
rect 6690 -29667 6708 -29611
rect 6764 -29667 6791 -29611
rect 6690 -29724 6791 -29667
rect -6943 -29782 2593 -29781
rect -7069 -29783 2593 -29782
rect -10942 -29797 2593 -29783
rect 3431 -29790 5244 -29761
rect 3431 -29793 4991 -29790
rect -34505 -29814 -34304 -29813
rect -34627 -29818 -34304 -29814
rect -35616 -29843 -34304 -29818
rect -998 -29821 2559 -29797
rect 3431 -29869 4844 -29793
rect 4918 -29866 4991 -29793
rect 5065 -29791 5244 -29790
rect 5065 -29866 5139 -29791
rect 4918 -29867 5139 -29866
rect 5213 -29867 5244 -29791
rect 6690 -29780 6708 -29724
rect 6764 -29727 6791 -29724
rect 6764 -29780 6988 -29727
rect 6690 -29799 6988 -29780
rect 6699 -29801 6988 -29799
rect 24984 -29772 26429 -29748
rect 24984 -29775 26318 -29772
rect 24984 -29845 26023 -29775
rect 26089 -29776 26318 -29775
rect 26089 -29845 26175 -29776
rect 24984 -29846 26175 -29845
rect 26241 -29842 26318 -29776
rect 26384 -29842 26429 -29772
rect 26241 -29846 26429 -29842
rect 24984 -29858 26429 -29846
rect 4918 -29869 5244 -29867
rect 3431 -29886 5244 -29869
rect -24703 -29982 -15406 -29935
rect -24703 -29984 -23092 -29982
rect -24703 -29990 -23232 -29984
rect -66387 -30037 -63178 -30019
rect -66387 -30044 -66217 -30037
rect -66387 -30126 -66366 -30044
rect -66289 -30119 -66217 -30044
rect -66140 -30038 -63178 -30037
rect -66140 -30119 -66067 -30038
rect -66289 -30120 -66067 -30119
rect -65990 -30120 -63178 -30038
rect -32962 -30075 -32851 -30014
rect -66289 -30126 -63178 -30120
rect -66387 -30137 -63178 -30126
rect -32965 -30135 -32851 -30075
rect -24703 -30075 -23386 -29990
rect -23320 -30069 -23232 -29990
rect -23166 -30067 -23092 -29984
rect -23026 -30067 -15406 -29982
rect -23166 -30069 -15406 -30067
rect -23320 -30075 -15406 -30069
rect -24703 -30092 -15406 -30075
rect -32965 -30207 -32935 -30135
rect -32865 -30207 -32851 -30135
rect 14111 -30094 20518 -30053
rect 14111 -30098 15636 -30094
rect 14111 -30101 15479 -30098
rect 14111 -30191 15334 -30101
rect 15405 -30188 15479 -30101
rect 15550 -30184 15636 -30098
rect 15707 -30184 20518 -30094
rect 15550 -30188 20518 -30184
rect 15405 -30191 20518 -30188
rect 14111 -30204 20518 -30191
rect -32965 -30289 -32851 -30207
rect -32965 -30361 -32943 -30289
rect -32873 -30306 -32851 -30289
rect -32873 -30361 -31818 -30306
rect -32965 -30417 -31818 -30361
rect 6397 -30446 7122 -30428
rect -59814 -30528 -56575 -30452
rect -59814 -30571 -56668 -30528
rect -56694 -30592 -56668 -30571
rect -56587 -30592 -56575 -30528
rect 6397 -30527 6412 -30446
rect 6492 -30527 7122 -30446
rect 6397 -30539 7122 -30527
rect -56694 -30679 -56575 -30592
rect -24203 -30639 -18489 -30583
rect -24203 -30642 -24024 -30639
rect -56694 -30743 -56677 -30679
rect -56596 -30743 -56575 -30679
rect -56694 -30762 -56575 -30743
rect -55946 -30701 -53673 -30642
rect -55946 -30704 -55781 -30701
rect -55946 -30767 -55913 -30704
rect -55853 -30764 -55781 -30704
rect -55721 -30704 -53673 -30701
rect -55721 -30764 -55647 -30704
rect -55853 -30767 -55647 -30764
rect -55587 -30767 -53673 -30704
rect -55946 -30792 -53673 -30767
rect -45764 -30705 -43273 -30642
rect -45764 -30708 -45603 -30705
rect -45764 -30771 -45735 -30708
rect -45675 -30768 -45603 -30708
rect -45543 -30708 -43273 -30705
rect -45543 -30768 -45469 -30708
rect -45675 -30771 -45469 -30768
rect -45409 -30771 -43273 -30708
rect -24203 -30705 -24156 -30642
rect -24096 -30702 -24024 -30642
rect -23964 -30642 -18489 -30639
rect -23964 -30702 -23890 -30642
rect -24096 -30705 -23890 -30702
rect -23830 -30705 -18489 -30642
rect 6397 -30587 6508 -30539
rect 6397 -30668 6415 -30587
rect 6495 -30668 6508 -30587
rect -24203 -30733 -18489 -30705
rect -45764 -30792 -43273 -30771
rect -7929 -30739 -4140 -30682
rect -7929 -30742 -7765 -30739
rect -7929 -30805 -7897 -30742
rect -7837 -30802 -7765 -30742
rect -7705 -30742 -4140 -30739
rect -7705 -30802 -7631 -30742
rect -7837 -30805 -7631 -30802
rect -7571 -30805 -4140 -30742
rect 6397 -30763 6508 -30668
rect 14636 -30719 17395 -30661
rect 14636 -30722 14792 -30719
rect -7929 -30832 -4140 -30805
rect 14636 -30785 14660 -30722
rect 14720 -30782 14792 -30722
rect 14852 -30722 17395 -30719
rect 14852 -30782 14926 -30722
rect 14720 -30785 14926 -30782
rect 14986 -30785 17395 -30722
rect 14636 -30811 17395 -30785
rect -68616 -31091 -67614 -30986
rect -66971 -31013 -65969 -30991
rect -66971 -31015 -66108 -31013
rect -66971 -31018 -66256 -31015
rect -66971 -31079 -66369 -31018
rect -66310 -31076 -66256 -31018
rect -66197 -31074 -66108 -31015
rect -66049 -31074 -65969 -31013
rect -66197 -31076 -65969 -31074
rect -66310 -31079 -65969 -31076
rect -66971 -31096 -65969 -31079
rect -24180 -31074 -23805 -31042
rect -24180 -31077 -24024 -31074
rect -24180 -31085 -24156 -31077
rect -45753 -31115 -45381 -31091
rect -55931 -31137 -55557 -31115
rect -55931 -31140 -55781 -31137
rect -55931 -31144 -55913 -31140
rect -59990 -31228 -56888 -31176
rect -55939 -31203 -55913 -31144
rect -55853 -31200 -55781 -31140
rect -55721 -31140 -55557 -31137
rect -55721 -31200 -55647 -31140
rect -55853 -31203 -55647 -31200
rect -55587 -31144 -55557 -31140
rect -45753 -31118 -45597 -31115
rect -45753 -31144 -45729 -31118
rect -55587 -31203 -53532 -31144
rect -55939 -31226 -53532 -31203
rect -45765 -31181 -45729 -31144
rect -45669 -31178 -45597 -31118
rect -45537 -31118 -45381 -31115
rect -45537 -31178 -45463 -31118
rect -45669 -31181 -45463 -31178
rect -45403 -31144 -45381 -31118
rect -24194 -31140 -24156 -31085
rect -24096 -31137 -24024 -31077
rect -23964 -31077 -23805 -31074
rect -23964 -31137 -23890 -31077
rect -24096 -31140 -23890 -31137
rect -23830 -31085 -23805 -31077
rect -23830 -31140 -18401 -31085
rect -45403 -31181 -43137 -31144
rect -24194 -31167 -18401 -31140
rect -45765 -31226 -43137 -31181
rect -7912 -31175 -7532 -31148
rect 14639 -31150 15018 -31132
rect 14639 -31153 14792 -31150
rect 14639 -31163 14660 -31153
rect -7912 -31178 -7765 -31175
rect -7912 -31183 -7897 -31178
rect -71037 -31444 -69405 -31342
rect -64242 -31364 -63942 -31278
rect -59990 -31300 -57009 -31228
rect -56906 -31300 -56888 -31228
rect -7920 -31241 -7897 -31183
rect -7837 -31238 -7765 -31178
rect -7705 -31178 -7532 -31175
rect -7705 -31238 -7631 -31178
rect -7837 -31241 -7631 -31238
rect -7571 -31183 -7532 -31178
rect -7571 -31241 -3995 -31183
rect -7920 -31266 -3995 -31241
rect 14628 -31216 14660 -31163
rect 14720 -31213 14792 -31153
rect 14852 -31153 15018 -31150
rect 14852 -31213 14926 -31153
rect 14720 -31216 14926 -31213
rect 14986 -31163 15018 -31153
rect 14986 -31216 17522 -31163
rect 14628 -31245 17522 -31216
rect -59990 -31324 -56888 -31300
rect -68728 -31455 -67712 -31367
rect -66995 -31371 -63942 -31364
rect -66995 -31457 -64149 -31371
rect -57036 -31408 -56888 -31324
rect -60010 -31544 -57253 -31414
rect -57036 -31480 -57019 -31408
rect -56916 -31480 -56888 -31408
rect -57036 -31500 -56888 -31480
rect -59900 -31584 -57253 -31544
rect -59900 -31620 -57382 -31584
rect -57459 -31663 -57382 -31620
rect -57283 -31663 -57253 -31584
rect -68622 -31806 -67620 -31701
rect -66938 -31714 -65275 -31698
rect -66938 -31717 -65522 -31714
rect -66938 -31778 -65665 -31717
rect -65606 -31775 -65522 -31717
rect -65463 -31719 -65275 -31714
rect -65463 -31775 -65397 -31719
rect -65606 -31778 -65397 -31775
rect -66938 -31780 -65397 -31778
rect -65338 -31780 -65275 -31719
rect -66938 -31803 -65275 -31780
rect -57459 -31751 -57253 -31663
rect -57459 -31830 -57379 -31751
rect -57280 -31830 -57253 -31751
rect -57459 -31854 -57253 -31830
rect 16368 -31906 16470 -31873
rect -54425 -31953 -54328 -31930
rect -54425 -32019 -54411 -31953
rect -54345 -32019 -54328 -31953
rect -54425 -32113 -54328 -32019
rect -43907 -31995 -43812 -31952
rect -43907 -32051 -43893 -31995
rect -43827 -32051 -43812 -31995
rect -43907 -32113 -43812 -32051
rect -19400 -31953 -19310 -31926
rect -19400 -32014 -19382 -31953
rect -19329 -32014 -19310 -31953
rect -19400 -32054 -19310 -32014
rect -4585 -31993 -4481 -31963
rect -19400 -32112 -18331 -32054
rect -54425 -32138 -53579 -32113
rect -54425 -32204 -54410 -32138
rect -54344 -32187 -53579 -32138
rect -43907 -32154 -43401 -32113
rect -54344 -32204 -54328 -32187
rect -54425 -32220 -54328 -32204
rect -43907 -32210 -43895 -32154
rect -43829 -32187 -43401 -32154
rect -19400 -32173 -19384 -32112
rect -19331 -32128 -18331 -32112
rect -4585 -32060 -4562 -31993
rect -4493 -32060 -4481 -31993
rect -19331 -32173 -19310 -32128
rect -43829 -32210 -43812 -32187
rect -19400 -32190 -19310 -32173
rect -4585 -32153 -4481 -32060
rect 16368 -31985 16383 -31906
rect 16454 -31985 16470 -31906
rect 16368 -32112 16470 -31985
rect -4585 -32170 -4152 -32153
rect -43907 -32230 -43812 -32210
rect -4585 -32237 -4568 -32170
rect -4499 -32227 -4152 -32170
rect 16368 -32191 16384 -32112
rect 16455 -32132 16470 -32112
rect 16455 -32191 17352 -32132
rect 16368 -32206 17352 -32191
rect -4499 -32237 -4481 -32227
rect -4585 -32257 -4481 -32237
rect -64569 -32400 -63786 -32293
rect -59558 -32338 -57585 -32326
rect -68649 -32575 -67647 -32470
rect -66965 -32494 -65963 -32480
rect -66965 -32507 -66098 -32494
rect -66965 -32509 -66231 -32507
rect -66965 -32570 -66371 -32509
rect -66312 -32568 -66231 -32509
rect -66172 -32555 -66098 -32507
rect -66039 -32555 -65963 -32494
rect -66172 -32568 -65963 -32555
rect -66312 -32570 -65963 -32568
rect -66965 -32585 -65963 -32570
rect -71062 -32928 -69429 -32827
rect -64569 -32843 -64462 -32400
rect -59647 -32415 -57585 -32338
rect -59647 -32486 -57715 -32415
rect -59558 -32497 -57715 -32486
rect -57756 -32502 -57715 -32497
rect -57596 -32502 -57585 -32415
rect -35383 -32464 -35024 -32462
rect -57756 -32637 -57585 -32502
rect -35394 -32467 -31987 -32464
rect -35394 -32470 -35243 -32467
rect -35394 -32533 -35375 -32470
rect -35315 -32530 -35243 -32470
rect -35183 -32470 -31987 -32467
rect -35183 -32530 -35109 -32470
rect -35315 -32533 -35109 -32530
rect -35049 -32533 -31987 -32470
rect -35394 -32546 -31987 -32533
rect -57756 -32724 -57733 -32637
rect -57614 -32724 -57585 -32637
rect 4071 -32591 6864 -32586
rect 4071 -32594 4220 -32591
rect 4071 -32657 4088 -32594
rect 4148 -32654 4220 -32594
rect 4280 -32594 6864 -32591
rect 4280 -32654 4354 -32594
rect 4148 -32657 4354 -32654
rect 4414 -32657 6864 -32594
rect 4071 -32668 6864 -32657
rect -57756 -32739 -57585 -32724
rect -68735 -32941 -67699 -32850
rect -66993 -32950 -64462 -32843
rect -53649 -33085 -53369 -33030
rect -53649 -33086 -53468 -33085
rect -53649 -33162 -53632 -33086
rect -53556 -33162 -53468 -33086
rect -53649 -33163 -53468 -33162
rect -53390 -33163 -53369 -33085
rect -68653 -33291 -67651 -33186
rect -66968 -33205 -65281 -33184
rect -66968 -33208 -65384 -33205
rect -66968 -33210 -65532 -33208
rect -66968 -33271 -65676 -33210
rect -65617 -33269 -65532 -33210
rect -65473 -33266 -65384 -33208
rect -65325 -33266 -65281 -33205
rect -53649 -33213 -53369 -33163
rect -43142 -33085 -42954 -33053
rect -43142 -33088 -43020 -33085
rect -43142 -33147 -43133 -33088
rect -43077 -33144 -43020 -33088
rect -42964 -33144 -42954 -33085
rect -43077 -33147 -42954 -33144
rect -43142 -33176 -42954 -33147
rect -18454 -33079 -18146 -33026
rect -18454 -33081 -18259 -33079
rect -18454 -33149 -18438 -33081
rect -18377 -33147 -18259 -33081
rect -18198 -33147 -18146 -33079
rect -18377 -33149 -18146 -33147
rect -18454 -33177 -18146 -33149
rect -4136 -33092 -3864 -33047
rect -4136 -33114 -3968 -33092
rect -4136 -33175 -4122 -33114
rect -4054 -33153 -3968 -33114
rect -3900 -33153 -3864 -33092
rect -4054 -33175 -3864 -33153
rect -4136 -33200 -3864 -33175
rect 17512 -33091 17772 -33037
rect 17512 -33093 17683 -33091
rect 17512 -33157 17525 -33093
rect 17583 -33155 17683 -33093
rect 17741 -33155 17772 -33091
rect 17583 -33157 17772 -33155
rect 17512 -33184 17772 -33157
rect -65473 -33269 -65281 -33266
rect -65617 -33271 -65281 -33269
rect -66968 -33289 -65281 -33271
rect -59563 -33293 -57936 -33273
rect -64657 -33371 -63561 -33325
rect -68659 -33753 -67657 -33648
rect -66974 -33681 -65972 -33652
rect -66974 -33683 -66078 -33681
rect -66974 -33744 -66369 -33683
rect -66310 -33744 -66216 -33683
rect -66157 -33742 -66078 -33683
rect -66019 -33742 -65972 -33681
rect -66157 -33744 -65972 -33742
rect -66974 -33757 -65972 -33744
rect -71037 -34090 -69458 -34000
rect -64657 -34006 -64544 -33371
rect -59652 -33392 -57936 -33293
rect -59652 -33422 -58055 -33392
rect -59563 -33440 -58055 -33422
rect -58103 -33473 -58055 -33440
rect -57975 -33473 -57936 -33392
rect -46563 -33417 -44568 -33361
rect -36175 -33379 -34303 -33361
rect -36175 -33382 -34393 -33379
rect -58103 -33592 -57936 -33473
rect -55297 -33443 -53609 -33417
rect -55297 -33446 -55126 -33443
rect -55297 -33509 -55258 -33446
rect -55198 -33506 -55126 -33446
rect -55066 -33446 -53609 -33443
rect -55066 -33506 -54992 -33446
rect -55198 -33509 -54992 -33506
rect -54932 -33509 -53609 -33446
rect -46563 -33447 -43160 -33417
rect -46563 -33450 -44789 -33447
rect -46563 -33461 -44921 -33450
rect -55297 -33534 -53609 -33509
rect -44945 -33513 -44921 -33461
rect -44861 -33510 -44789 -33450
rect -44729 -33450 -43160 -33447
rect -44729 -33510 -44655 -33450
rect -44861 -33513 -44655 -33510
rect -44595 -33513 -43160 -33450
rect -36175 -33450 -34697 -33382
rect -34640 -33450 -34562 -33382
rect -34505 -33447 -34393 -33382
rect -34336 -33447 -34303 -33379
rect -23398 -33381 -18342 -33358
rect -23398 -33384 -23248 -33381
rect -34505 -33450 -34303 -33447
rect -36175 -33461 -34303 -33450
rect -44945 -33534 -43160 -33513
rect -30639 -33519 -30593 -33425
rect -23398 -33447 -23380 -33384
rect -23320 -33444 -23248 -33384
rect -23188 -33384 -18342 -33381
rect -23188 -33444 -23114 -33384
rect -23320 -33447 -23114 -33444
rect -23054 -33447 -18342 -33384
rect -11345 -33402 -7180 -33302
rect 24579 -33395 26426 -33380
rect 24579 -33399 26311 -33395
rect -23398 -33475 -18342 -33447
rect -7280 -33424 -7180 -33402
rect 3017 -33417 5239 -33401
rect 3017 -33419 4998 -33417
rect -7280 -33457 -6812 -33424
rect -7280 -33485 -4019 -33457
rect -7280 -33488 -6996 -33485
rect -7280 -33524 -7128 -33488
rect -7144 -33551 -7128 -33524
rect -7068 -33548 -6996 -33488
rect -6936 -33488 -4019 -33485
rect -6936 -33548 -6862 -33488
rect -7068 -33551 -6862 -33548
rect -6802 -33551 -4019 -33488
rect 3017 -33486 4841 -33419
rect 4907 -33484 4998 -33419
rect 5064 -33418 5239 -33417
rect 5064 -33484 5135 -33418
rect 4907 -33485 5135 -33484
rect 5201 -33485 5239 -33418
rect 4907 -33486 5239 -33485
rect 3017 -33501 5239 -33486
rect 15315 -33462 17591 -33436
rect 15315 -33465 15480 -33462
rect -7144 -33574 -4019 -33551
rect 15315 -33528 15348 -33465
rect 15408 -33525 15480 -33465
rect 15540 -33465 17591 -33462
rect 15540 -33525 15614 -33465
rect 15408 -33528 15614 -33525
rect 15674 -33528 17591 -33465
rect 24579 -33469 26028 -33399
rect 26094 -33469 26162 -33399
rect 26228 -33465 26311 -33399
rect 26377 -33465 26426 -33395
rect 26228 -33469 26426 -33465
rect 24579 -33480 26426 -33469
rect 15315 -33553 17591 -33528
rect -58103 -33673 -58069 -33592
rect -57989 -33673 -57936 -33592
rect 8172 -33658 8218 -33557
rect -58103 -33692 -57936 -33673
rect -68765 -34108 -67705 -34018
rect -66993 -34119 -64544 -34006
rect -54118 -34227 -54041 -34188
rect -58450 -34264 -58287 -34259
rect -68650 -34457 -67678 -34348
rect -66962 -34379 -65275 -34353
rect -66962 -34382 -65545 -34379
rect -66962 -34443 -65683 -34382
rect -65624 -34440 -65545 -34382
rect -65486 -34440 -65399 -34379
rect -65340 -34440 -65275 -34379
rect -60923 -34399 -58287 -34264
rect -60923 -34401 -58410 -34399
rect -65624 -34443 -65275 -34440
rect -66962 -34458 -65275 -34443
rect -58450 -34481 -58410 -34401
rect -58313 -34481 -58287 -34399
rect -54118 -34289 -54103 -34227
rect -54050 -34289 -54041 -34227
rect -18970 -34196 -18893 -34184
rect -54118 -34355 -54041 -34289
rect -43622 -34255 -43545 -34228
rect -43622 -34308 -43609 -34255
rect -43554 -34308 -43545 -34255
rect -54118 -34417 -54109 -34355
rect -54056 -34367 -54041 -34355
rect -54056 -34417 -53664 -34367
rect -51475 -34407 -50479 -34335
rect -43622 -34367 -43545 -34308
rect -18970 -34257 -18964 -34196
rect -18901 -34257 -18893 -34196
rect -18970 -34308 -18893 -34257
rect -18970 -34316 -18398 -34308
rect -43622 -34381 -43273 -34367
rect -54118 -34444 -53664 -34417
rect -43622 -34434 -43614 -34381
rect -43559 -34434 -43273 -34381
rect -41054 -34407 -40218 -34335
rect -18970 -34377 -18963 -34316
rect -18900 -34377 -18398 -34316
rect -16242 -34348 -15411 -34276
rect -32293 -34404 -32203 -34378
rect -18970 -34385 -18398 -34377
rect -18970 -34393 -18893 -34385
rect -43622 -34444 -43273 -34434
rect -58450 -34579 -58287 -34481
rect -58450 -34661 -58415 -34579
rect -58318 -34661 -58287 -34579
rect -32293 -34461 -32275 -34404
rect -32218 -34461 -32203 -34404
rect -32293 -34545 -32203 -34461
rect -4198 -34404 -3878 -34379
rect -4198 -34415 -4001 -34404
rect -4198 -34513 -4166 -34415
rect -4075 -34502 -4001 -34415
rect -3910 -34502 -3878 -34404
rect -1866 -34447 -962 -34375
rect 17352 -34405 17660 -34373
rect 17352 -34469 17381 -34405
rect 17446 -34469 17499 -34405
rect 17564 -34469 17660 -34405
rect 19701 -34426 20490 -34354
rect 17352 -34500 17660 -34469
rect -4075 -34513 -3878 -34502
rect -4198 -34540 -3878 -34513
rect 5587 -34522 5674 -34509
rect -32293 -34546 -31877 -34545
rect -58450 -34689 -58287 -34661
rect -57159 -34745 -56769 -34597
rect -32293 -34601 -32275 -34546
rect -32220 -34601 -31877 -34546
rect -32293 -34602 -31877 -34601
rect 5587 -34579 5606 -34522
rect 5663 -34579 5674 -34522
rect -32293 -34609 -32203 -34602
rect 5587 -34667 5674 -34579
rect 5587 -34668 7070 -34667
rect 5587 -34723 5607 -34668
rect 5662 -34723 7070 -34668
rect 5587 -34724 7070 -34723
rect 5587 -34731 5674 -34724
rect -57159 -34999 -57011 -34745
rect -34713 -34905 -31856 -34879
rect -34864 -34909 -31856 -34905
rect -34864 -34912 -34553 -34909
rect -46416 -35006 -44535 -34945
rect -59151 -35223 -58258 -35209
rect -59200 -35348 -58258 -35223
rect -59151 -35360 -58258 -35348
rect -58409 -35555 -58258 -35360
rect -57084 -35539 -56886 -35473
rect -65695 -35605 -63173 -35577
rect -65695 -35610 -65411 -35605
rect -65695 -35613 -65544 -35610
rect -65695 -35679 -65687 -35613
rect -65624 -35676 -65544 -35613
rect -65481 -35671 -65411 -35610
rect -65348 -35671 -63173 -35605
rect -65481 -35676 -63173 -35671
rect -58409 -35643 -58002 -35555
rect -57209 -35591 -56886 -35539
rect -55389 -35492 -54317 -35480
rect -55389 -35544 -54305 -35492
rect -58409 -35675 -58258 -35643
rect -57209 -35657 -56966 -35591
rect -55389 -35603 -54413 -35544
rect -54443 -35604 -54413 -35603
rect -54350 -35604 -54305 -35544
rect -54443 -35630 -54305 -35604
rect -65624 -35679 -63173 -35676
rect -65695 -35690 -63173 -35679
rect -52974 -36105 -52826 -35057
rect -46416 -35077 -44922 -35006
rect -44867 -35010 -44535 -35006
rect -44867 -35077 -44782 -35010
rect -46416 -35081 -44782 -35077
rect -44727 -35021 -44535 -35010
rect -44727 -35081 -44632 -35021
rect -46416 -35092 -44632 -35081
rect -44577 -35066 -44535 -35021
rect -34864 -34975 -34685 -34912
rect -34625 -34972 -34553 -34912
rect -34493 -34912 -31856 -34909
rect -34493 -34972 -34419 -34912
rect -34625 -34975 -34419 -34972
rect -34359 -34975 -31856 -34912
rect -34864 -34992 -31856 -34975
rect -24695 -34906 -18747 -34860
rect -24695 -34909 -23087 -34906
rect -24695 -34911 -23236 -34909
rect -34864 -35050 -34300 -34992
rect -24695 -34995 -23389 -34911
rect -23317 -34993 -23236 -34911
rect -23164 -34990 -23087 -34909
rect -23015 -34976 -18747 -34906
rect -23015 -34990 -4715 -34976
rect -23164 -34993 -4715 -34990
rect -23317 -34995 -4715 -34993
rect -24695 -35017 -4715 -34995
rect -18904 -35021 -6842 -35017
rect -18904 -35025 -6984 -35021
rect -34864 -35066 -34719 -35050
rect -44577 -35092 -34719 -35066
rect -46416 -35137 -34719 -35092
rect -18904 -35114 -7137 -35025
rect -7071 -35110 -6984 -35025
rect -6918 -35106 -6842 -35021
rect -6776 -35100 -4715 -35017
rect 4828 -35027 7030 -35001
rect 4828 -35030 4985 -35027
rect 4828 -35093 4853 -35030
rect 4913 -35090 4985 -35030
rect 5045 -35030 7030 -35027
rect 5045 -35090 5119 -35030
rect 4913 -35093 5119 -35090
rect 5179 -35093 7030 -35030
rect 4828 -35100 7030 -35093
rect -6776 -35106 7030 -35100
rect -6918 -35110 7030 -35106
rect -7071 -35114 7030 -35110
rect 14117 -35017 15724 -34985
rect 14117 -35021 15601 -35017
rect 14117 -35111 15333 -35021
rect 15404 -35111 15470 -35021
rect 15541 -35107 15601 -35021
rect 15672 -35061 15724 -35017
rect 15672 -35083 26428 -35061
rect 15672 -35085 26175 -35083
rect 15672 -35107 26033 -35085
rect 15541 -35111 26033 -35107
rect -18904 -35133 5198 -35114
rect -44626 -35211 -34719 -35137
rect -32094 -35182 -32000 -35150
rect -32094 -35207 -31823 -35182
rect -32094 -35260 -32072 -35207
rect -32010 -35260 -31823 -35207
rect -4872 -35257 5198 -35133
rect 14117 -35139 26033 -35111
rect 15459 -35155 26033 -35139
rect 26099 -35153 26175 -35085
rect 26241 -35088 26428 -35083
rect 26241 -35153 26315 -35088
rect 26099 -35155 26315 -35153
rect 15459 -35158 26315 -35155
rect 26381 -35158 26428 -35088
rect 15459 -35172 26428 -35158
rect 5408 -35236 5502 -35226
rect -32094 -35276 -31823 -35260
rect -32094 -35355 -32000 -35276
rect -32094 -35408 -32075 -35355
rect -32013 -35408 -32000 -35355
rect -32094 -35425 -32000 -35408
rect 5408 -35299 5426 -35236
rect 5486 -35299 5502 -35236
rect 5408 -35304 5502 -35299
rect 5408 -35369 7098 -35304
rect 17853 -35340 17965 -35337
rect 5408 -35432 5426 -35369
rect 5486 -35398 7098 -35369
rect 5486 -35432 5502 -35398
rect 5408 -35451 5502 -35432
rect 17852 -35419 17989 -35340
rect 17852 -35499 17882 -35419
rect 17963 -35499 17989 -35419
rect -3701 -35547 -3399 -35541
rect 6122 -35545 6536 -35533
rect 6122 -35547 6399 -35545
rect -3701 -35558 6399 -35547
rect -3701 -35567 6128 -35558
rect -3701 -35569 -3515 -35567
rect -56741 -36150 -52826 -36105
rect -56741 -36228 -55277 -36150
rect -55219 -36228 -55148 -36150
rect -55090 -36156 -52826 -36150
rect -55090 -36228 -55002 -36156
rect -56741 -36234 -55002 -36228
rect -54944 -36234 -52826 -36156
rect -56741 -36253 -52826 -36234
rect -50450 -35802 -12770 -35649
rect -57408 -36485 -57252 -36414
rect -57408 -36552 -57382 -36485
rect -57288 -36543 -57252 -36485
rect -50450 -36543 -50297 -35802
rect -57288 -36552 -50297 -36543
rect -57408 -36623 -50297 -36552
rect -57408 -36690 -57382 -36623
rect -57288 -36690 -50297 -36623
rect -57408 -36696 -50297 -36690
rect -49934 -36204 -28283 -36044
rect -57408 -36718 -57252 -36696
rect -58103 -36892 -57936 -36811
rect -58103 -36963 -58065 -36892
rect -57992 -36963 -57936 -36892
rect -58103 -36989 -57936 -36963
rect -49934 -36989 -49774 -36204
rect -48612 -36553 -48204 -36405
rect -47480 -36418 -45350 -36405
rect -47480 -36426 -45463 -36418
rect -47480 -36524 -45753 -36426
rect -45695 -36524 -45595 -36426
rect -45537 -36516 -45463 -36426
rect -45405 -36516 -45350 -36418
rect -45537 -36524 -45350 -36516
rect -47480 -36553 -45350 -36524
rect -48612 -36768 -48464 -36553
rect -58103 -37049 -49774 -36989
rect -58103 -37120 -58062 -37049
rect -57989 -37120 -49774 -37049
rect -28443 -36906 -28283 -36204
rect -26925 -36142 -26516 -35994
rect -25183 -36034 -23791 -35994
rect -25183 -36035 -24036 -36034
rect -25183 -36120 -24177 -36035
rect -24120 -36119 -24036 -36035
rect -23979 -36035 -23791 -36034
rect -23979 -36119 -23891 -36035
rect -24120 -36120 -23891 -36119
rect -23834 -36120 -23791 -36035
rect -25183 -36142 -23791 -36120
rect -26925 -36270 -26777 -36142
rect -28443 -36933 -28059 -36906
rect -28443 -37038 -27731 -36933
rect -26825 -36936 -26605 -36875
rect -19584 -36877 -19260 -36830
rect -26885 -36993 -26605 -36936
rect -25127 -36884 -19260 -36877
rect -25127 -36895 -19388 -36884
rect -25127 -36980 -19550 -36895
rect -19493 -36969 -19388 -36895
rect -19331 -36969 -19260 -36884
rect -19493 -36980 -19260 -36969
rect -28443 -37066 -28059 -37038
rect -26885 -37054 -26707 -36993
rect -25127 -37000 -19260 -36980
rect -19584 -37033 -19260 -37000
rect -12923 -37036 -12770 -35802
rect -4005 -35693 -3852 -35596
rect -3701 -35637 -3675 -35569
rect -3605 -35635 -3515 -35569
rect -3445 -35635 6128 -35567
rect -3605 -35637 6128 -35635
rect -3701 -35648 6128 -35637
rect 6218 -35648 6399 -35558
rect -3701 -35659 6399 -35648
rect -3701 -35667 -3399 -35659
rect 6122 -35661 6399 -35659
rect 6495 -35547 6536 -35545
rect 17852 -35547 17989 -35499
rect 6495 -35559 17989 -35547
rect 6495 -35639 17881 -35559
rect 17962 -35639 17989 -35559
rect 6495 -35659 17989 -35639
rect 6495 -35661 6536 -35659
rect 6122 -35681 6536 -35661
rect 17852 -35667 17989 -35659
rect -4005 -35770 -3975 -35693
rect -3883 -35770 -3852 -35693
rect -4005 -35837 -3852 -35770
rect 6366 -35837 6828 -35815
rect -4005 -35838 17657 -35837
rect -4005 -35935 -3985 -35838
rect -3866 -35839 17657 -35838
rect -3866 -35844 6687 -35839
rect -3866 -35931 6418 -35844
rect 6526 -35931 6687 -35844
rect -3866 -35935 6687 -35931
rect -4005 -35936 6687 -35935
rect 6811 -35857 17657 -35839
rect 6811 -35861 17557 -35857
rect 6811 -35936 17255 -35861
rect -4005 -35938 17255 -35936
rect 17337 -35862 17557 -35861
rect 17337 -35938 17403 -35862
rect -4005 -35939 17403 -35938
rect 17485 -35934 17557 -35862
rect 17639 -35934 17657 -35857
rect 17485 -35939 17657 -35934
rect -4005 -35958 17657 -35939
rect -4005 -35959 -3852 -35958
rect 6366 -35982 6828 -35958
rect -11295 -36140 -7505 -36104
rect -11295 -36146 -7611 -36140
rect -11295 -36150 -7758 -36146
rect -11295 -36231 -7898 -36150
rect -7842 -36227 -7758 -36150
rect -7702 -36221 -7611 -36146
rect -7555 -36221 -7505 -36140
rect -7702 -36227 -7505 -36221
rect -7842 -36231 -7505 -36227
rect -11295 -36252 -7505 -36231
rect 1495 -36216 4472 -36168
rect -11295 -36440 -11147 -36252
rect 1495 -36297 4082 -36216
rect 4138 -36297 4243 -36216
rect 4299 -36218 4472 -36216
rect 4299 -36297 4400 -36218
rect 1495 -36299 4400 -36297
rect 4456 -36299 4472 -36218
rect 1495 -36316 4472 -36299
rect 1495 -36469 1643 -36316
rect 12644 -36435 13149 -36287
rect 13721 -36289 15036 -36287
rect 13721 -36328 20617 -36289
rect 13721 -36332 14793 -36328
rect 13721 -36414 14656 -36332
rect 14723 -36410 14793 -36332
rect 14860 -36332 20617 -36328
rect 14860 -36410 14935 -36332
rect 14723 -36414 14935 -36410
rect 15002 -36414 20617 -36332
rect 13721 -36435 20617 -36414
rect 12644 -36632 12792 -36435
rect 14877 -36437 20617 -36435
rect 20469 -36639 20617 -36437
rect -4742 -36979 -4410 -36958
rect -9324 -36987 -4410 -36979
rect -58103 -37149 -49774 -37120
rect -58103 -37152 -57936 -37149
rect -26796 -37167 -26750 -37054
rect -12923 -37067 -12413 -37036
rect -11200 -37046 -10992 -37000
rect -12923 -37157 -12118 -37067
rect -11339 -37096 -10992 -37046
rect -9511 -37031 -4410 -36987
rect -9511 -37038 -4584 -37031
rect -12923 -37189 -12413 -37157
rect -11339 -37164 -11151 -37096
rect -9511 -37110 -4705 -37038
rect -9324 -37117 -4705 -37110
rect -4742 -37121 -4705 -37117
rect -4648 -37114 -4584 -37038
rect -4527 -37114 -4410 -37031
rect 5764 -37051 6006 -37027
rect 1620 -37110 1804 -37065
rect -4648 -37121 -4410 -37114
rect -4742 -37153 -4410 -37121
rect -377 -37171 378 -37118
rect 1471 -37151 1804 -37110
rect 3306 -37071 6006 -37051
rect 3306 -37076 5919 -37071
rect -377 -37252 703 -37171
rect 1471 -37228 1716 -37151
rect 3306 -37158 5792 -37076
rect 5848 -37153 5919 -37076
rect 5975 -37153 6006 -37071
rect 5848 -37158 6006 -37153
rect 3306 -37174 6006 -37158
rect 5764 -37188 6006 -37174
rect 14538 -37199 16483 -37170
rect 14538 -37205 16357 -37199
rect 1641 -37232 1716 -37228
rect 11183 -37233 11648 -37208
rect -43941 -37288 -43741 -37267
rect -58448 -37406 -49415 -37375
rect -58448 -37459 -58410 -37406
rect -58341 -37459 -49415 -37406
rect -48525 -37410 -48301 -37305
rect -46815 -37312 -43741 -37288
rect -46815 -37313 -43808 -37312
rect -46815 -37411 -43923 -37313
rect -43865 -37410 -43808 -37313
rect -43750 -37410 -43741 -37312
rect -43865 -37411 -43741 -37410
rect -43941 -37443 -43741 -37411
rect -377 -37307 378 -37252
rect -58448 -37472 -49415 -37459
rect -26460 -37536 -22991 -37502
rect -26460 -37538 -23089 -37536
rect -26460 -37548 -23229 -37538
rect -26460 -37633 -23380 -37548
rect -23323 -37623 -23229 -37548
rect -23172 -37621 -23089 -37538
rect -23032 -37621 -22991 -37536
rect -23172 -37623 -22991 -37621
rect -23323 -37633 -22991 -37623
rect -26460 -37650 -22991 -37633
rect -10844 -37649 -6739 -37612
rect -10844 -37658 -6858 -37649
rect -10844 -37663 -6982 -37658
rect -10844 -37744 -7132 -37663
rect -7076 -37739 -6982 -37663
rect -6926 -37730 -6858 -37658
rect -6802 -37730 -6739 -37649
rect -6926 -37739 -6739 -37730
rect -7076 -37744 -6739 -37739
rect -10844 -37760 -6739 -37744
rect -48148 -37948 -44540 -37913
rect -48148 -37953 -44623 -37948
rect -57756 -38058 -57585 -38014
rect -57756 -38116 -57731 -38058
rect -57631 -38116 -57585 -38058
rect -48148 -38051 -44929 -37953
rect -44871 -38051 -44782 -37953
rect -44724 -38046 -44623 -37953
rect -44565 -38046 -44540 -37948
rect -44724 -38051 -44540 -38046
rect -48148 -38061 -44540 -38051
rect -57756 -38186 -57585 -38116
rect -57756 -38244 -57732 -38186
rect -57632 -38193 -57585 -38186
rect -377 -38193 -188 -37307
rect 11183 -37356 11947 -37233
rect 12874 -37318 13059 -37205
rect 14538 -37266 16226 -37205
rect 16291 -37260 16357 -37205
rect 16422 -37260 16483 -37199
rect 16291 -37266 16483 -37260
rect 14538 -37293 16483 -37266
rect 16799 -37172 17156 -37162
rect 16799 -37200 18756 -37172
rect 16799 -37202 17067 -37200
rect 16799 -37209 16950 -37202
rect 16799 -37283 16823 -37209
rect 16883 -37276 16950 -37209
rect 17010 -37274 17067 -37202
rect 17127 -37274 18756 -37200
rect 17010 -37276 18756 -37274
rect 16883 -37283 18756 -37276
rect 16799 -37295 18756 -37283
rect 20259 -37231 20402 -37203
rect 16799 -37301 17156 -37295
rect 20259 -37314 20599 -37231
rect 21655 -37244 22052 -37201
rect 20371 -37349 20599 -37314
rect 21360 -37351 22052 -37244
rect 11183 -37383 11648 -37356
rect 1973 -37714 5251 -37676
rect 1973 -37716 5125 -37714
rect 1973 -37804 4856 -37716
rect 4919 -37804 4998 -37716
rect 5061 -37802 5125 -37716
rect 5188 -37802 5251 -37714
rect 5061 -37804 5251 -37802
rect 1973 -37824 5251 -37804
rect -57632 -38244 -188 -38193
rect -57756 -38296 -188 -38244
rect -57756 -38354 -57731 -38296
rect -57631 -38354 -188 -38296
rect -57756 -38382 -188 -38354
rect -57756 -38383 -57585 -38382
rect -56707 -38680 -56561 -38595
rect -56707 -38730 -56683 -38680
rect -56708 -38745 -56683 -38730
rect -56580 -38730 -56561 -38680
rect 11183 -38730 11358 -37383
rect 21655 -37396 22052 -37351
rect 13205 -37797 15724 -37795
rect 13205 -37840 20064 -37797
rect 13205 -37841 15617 -37840
rect 13205 -37923 15331 -37841
rect 15398 -37923 15466 -37841
rect 15533 -37922 15617 -37841
rect 15684 -37922 20064 -37840
rect 15533 -37923 20064 -37922
rect 13205 -37943 20064 -37923
rect 15531 -37945 20064 -37943
rect -56580 -38745 11358 -38730
rect -56708 -38816 11358 -38745
rect -56708 -38881 -56690 -38816
rect -56587 -38881 11358 -38816
rect -56708 -38905 11358 -38881
rect -56707 -38906 -56561 -38905
rect -57036 -39064 -56888 -38988
rect -57036 -39128 -57012 -39064
rect -56931 -39128 -56888 -39064
rect -57036 -39190 -56888 -39128
rect -57036 -39237 -57008 -39190
rect -57059 -39254 -57008 -39237
rect -56927 -39237 -56888 -39190
rect 21857 -39237 22052 -37396
rect -56927 -39254 22052 -39237
rect -57059 -39315 22052 -39254
rect -57059 -39379 -57010 -39315
rect -56929 -39379 22052 -39315
rect -57059 -39432 22052 -39379
<< via1 >>
rect -66351 60691 -66237 60795
rect -66142 60696 -66028 60800
rect -66354 60526 -66240 60630
rect -66141 60525 -66027 60629
rect -66351 60000 -66237 60104
rect -66128 60000 -66014 60104
rect -66350 59843 -66236 59947
rect -66128 59844 -66014 59948
rect -70897 57087 -70844 57140
rect -70742 57088 -70689 57141
rect -70584 57088 -70531 57141
rect -70895 56981 -70842 57034
rect -70738 56978 -70685 57031
rect -70585 56978 -70532 57031
rect -70896 56872 -70843 56925
rect -70738 56873 -70685 56926
rect -70586 56871 -70533 56924
rect -70893 56763 -70840 56816
rect -70737 56762 -70684 56815
rect -70584 56762 -70531 56815
rect -70210 57086 -70157 57139
rect -70055 57087 -70002 57140
rect -69897 57087 -69844 57140
rect -70208 56980 -70155 57033
rect -70051 56977 -69998 57030
rect -69898 56977 -69845 57030
rect -70209 56871 -70156 56924
rect -70051 56872 -69998 56925
rect -69899 56870 -69846 56923
rect -70206 56762 -70153 56815
rect -70050 56761 -69997 56814
rect -69897 56761 -69844 56814
rect -66369 57122 -66316 57175
rect -66214 57123 -66161 57176
rect -66056 57123 -66003 57176
rect -66367 57016 -66314 57069
rect -66210 57013 -66157 57066
rect -66057 57013 -66004 57066
rect -66368 56907 -66315 56960
rect -66210 56908 -66157 56961
rect -66058 56906 -66005 56959
rect -66365 56798 -66312 56851
rect -66209 56797 -66156 56850
rect -66056 56797 -66003 56850
rect -65683 57118 -65630 57171
rect -65528 57119 -65475 57172
rect -65370 57119 -65317 57172
rect -65681 57012 -65628 57065
rect -65524 57009 -65471 57062
rect -65371 57009 -65318 57062
rect -65682 56903 -65629 56956
rect -65524 56904 -65471 56957
rect -65372 56902 -65319 56955
rect -65679 56794 -65626 56847
rect -65523 56793 -65470 56846
rect -65370 56793 -65317 56846
rect -8560 56713 -8508 56766
rect -8423 56712 -8371 56765
rect -8555 56567 -8503 56620
rect -8409 56567 -8357 56620
rect -43752 52520 -43678 52594
rect -53932 52343 -53860 52415
rect -43752 52341 -43678 52415
rect -32393 52342 -32319 52416
rect -32152 52342 -32078 52416
rect -18434 52336 -18347 52423
rect -4639 52373 -4563 52449
rect 6516 52372 6594 52450
rect 6681 52372 6759 52450
rect 16664 52362 16763 52461
rect 16857 52363 16954 52460
rect -53933 52120 -53859 52194
rect -53671 52067 -53573 52165
rect -43453 52067 -43355 52165
rect -32642 52066 -32542 52166
rect -32415 52066 -32315 52166
rect -18775 52067 -18677 52165
rect -18434 52132 -18345 52221
rect -4640 52173 -4562 52251
rect -53672 51887 -53572 51987
rect -43454 51851 -43354 51951
rect -18776 51828 -18676 51928
rect -4366 52090 -4261 52195
rect 6370 52089 6477 52196
rect 17284 52090 17389 52195
rect -4366 51863 -4259 51970
rect 6371 51884 6476 51989
rect 17283 51886 17390 51993
rect -32152 51743 -32078 51817
rect -46588 51638 -46533 51694
rect 6681 51692 6759 51770
rect -46382 51499 -46327 51555
rect -36227 51525 -36172 51581
rect -32151 51571 -32079 51643
rect 2700 51581 2755 51637
rect 6682 51530 6758 51606
rect 24420 51525 24475 51581
rect 2906 51442 2961 51498
rect -36021 51386 -35966 51442
rect 24626 51386 24681 51442
rect -44929 51306 -44876 51363
rect -44814 51306 -44761 51363
rect -44678 51305 -44625 51362
rect -34692 51187 -34618 51258
rect -34546 51190 -34472 51261
rect -34395 51193 -34321 51264
rect -23385 51196 -23314 51271
rect -23234 51198 -23163 51273
rect -23089 51197 -23018 51272
rect -7131 51185 -7078 51261
rect -7009 51184 -6956 51260
rect -6869 51187 -6816 51263
rect 4845 51240 4907 51316
rect 4973 51239 5035 51315
rect 5158 51243 5220 51319
rect -32421 51057 -32310 51168
rect 15334 51153 15395 51242
rect 15482 51152 15543 51241
rect 15644 51152 15705 51241
rect 26024 51178 26083 51260
rect 26161 51180 26220 51262
rect 26325 51183 26384 51265
rect 6368 51018 6479 51129
rect -32421 50833 -32312 50942
rect 6369 50793 6478 50902
rect -55901 50355 -55841 50418
rect -55769 50358 -55709 50421
rect -55635 50355 -55575 50418
rect -45745 50242 -45685 50305
rect -45613 50245 -45553 50308
rect -45479 50242 -45419 50305
rect -24169 50246 -24109 50309
rect -24037 50249 -23977 50312
rect -23903 50246 -23843 50309
rect -7883 50299 -7823 50362
rect -7751 50302 -7691 50365
rect -7617 50299 -7557 50362
rect 14660 50231 14720 50294
rect 14792 50234 14852 50297
rect 14926 50231 14986 50294
rect -53252 50012 -53161 50091
rect -53256 49860 -53165 49939
rect -42873 49905 -42782 49984
rect -17978 49888 -17887 49967
rect -3887 49925 -3796 50004
rect -42877 49753 -42786 49832
rect -17982 49736 -17891 49815
rect -3891 49773 -3800 49852
rect 16552 49846 16623 49916
rect 16549 49675 16620 49745
rect -66361 49539 -66296 49597
rect -66220 49541 -66155 49599
rect -66090 49548 -66025 49606
rect -65668 48827 -65603 48885
rect -65525 48825 -65460 48883
rect -65393 48829 -65328 48887
rect -66365 48062 -66300 48120
rect -66223 48061 -66158 48119
rect -66078 48061 -66013 48119
rect -65661 47357 -65596 47415
rect -65522 47354 -65457 47412
rect -65377 47358 -65312 47416
rect -66365 46596 -66300 46654
rect -66232 46605 -66167 46663
rect -66086 46625 -66021 46683
rect -65667 45901 -65602 45959
rect -65526 45902 -65461 45960
rect -65383 45911 -65318 45969
rect -66357 43148 -66293 43230
rect -66216 43143 -66152 43225
rect -66069 43153 -66005 43235
rect -68358 42888 -68297 42954
rect -67772 42874 -67706 42944
rect -50866 48978 -50812 49032
rect -54492 48888 -54412 48965
rect -54492 48700 -54412 48777
rect -43940 48913 -43888 48973
rect -40505 48865 -40451 48919
rect -43938 48794 -43886 48854
rect -15682 48865 -15628 48919
rect -19370 48785 -19289 48853
rect -4950 48861 -4873 48936
rect -1578 48921 -1524 48975
rect -35380 48713 -35320 48776
rect -35248 48716 -35188 48779
rect -35114 48713 -35054 48776
rect -19377 48645 -19296 48713
rect 15350 48846 15410 48909
rect 15482 48849 15542 48912
rect 15616 48846 15676 48909
rect 20142 48865 20196 48919
rect -4951 48688 -4874 48763
rect 4080 48674 4140 48737
rect 4212 48677 4272 48740
rect 4346 48674 4406 48737
rect -55259 47985 -55199 48048
rect -55127 47988 -55067 48051
rect -54993 47985 -54933 48048
rect -8564 48039 -8508 48136
rect -8419 48042 -8363 48139
rect -44915 47872 -44855 47935
rect -44783 47875 -44723 47938
rect -44649 47872 -44589 47935
rect -23381 47867 -23321 47930
rect -23249 47870 -23189 47933
rect -23115 47867 -23055 47930
rect -55271 47606 -55211 47669
rect -55139 47609 -55079 47672
rect -55005 47606 -54945 47669
rect -44908 47501 -44848 47564
rect -44776 47504 -44716 47567
rect -44642 47501 -44582 47564
rect -53933 46793 -53856 46870
rect -53936 46650 -53855 46731
rect -50819 46471 -50764 46530
rect -43454 47097 -43354 47197
rect -43282 47098 -43184 47196
rect -43752 46555 -43678 46629
rect -43597 46555 -43523 46629
rect -40458 46358 -40403 46417
rect -23383 47495 -23323 47558
rect -23251 47498 -23191 47561
rect -23117 47495 -23057 47558
rect -18960 47089 -18862 47187
rect -18775 47088 -18675 47188
rect -7122 47919 -7062 47982
rect -6990 47922 -6930 47985
rect -6856 47919 -6796 47982
rect 16787 47952 16840 48012
rect 16781 47809 16834 47869
rect -7873 47634 -7813 47697
rect -7741 47637 -7681 47700
rect -7607 47634 -7547 47697
rect -7123 47546 -7063 47609
rect -6991 47549 -6931 47612
rect -6857 47546 -6797 47609
rect 4844 47616 4902 47685
rect 4979 47619 5037 47688
rect 5128 47617 5186 47686
rect 15342 47491 15402 47554
rect 15474 47494 15534 47557
rect 15608 47491 15668 47554
rect 26026 47556 26085 47638
rect 26164 47556 26223 47638
rect 26306 47560 26365 47642
rect -8599 47388 -8546 47442
rect -8468 47386 -8415 47440
rect -8594 47244 -8541 47298
rect -8464 47246 -8411 47300
rect -7118 46935 -7058 46998
rect -6986 46938 -6926 47001
rect -6852 46935 -6792 46998
rect -31908 46648 -31853 46703
rect -31785 46647 -31728 46704
rect -18434 46556 -18345 46645
rect -18276 46557 -18189 46644
rect -4647 46618 -4552 46713
rect -4457 46619 -4364 46712
rect 6977 46608 7032 46663
rect 7098 46608 7153 46663
rect -34682 46271 -34622 46334
rect -34550 46274 -34490 46337
rect -34416 46271 -34356 46334
rect -15635 46358 -15580 46417
rect -1531 46414 -1476 46473
rect -23383 46265 -23320 46342
rect -23240 46264 -23177 46341
rect -23101 46264 -23038 46341
rect 17013 46737 17105 46829
rect 17012 46574 17106 46668
rect 20189 46358 20244 46417
rect 4849 46228 4909 46291
rect 4981 46231 5041 46294
rect 5115 46228 5175 46291
rect -7129 45906 -7059 46003
rect -6984 45902 -6914 45999
rect -6836 45909 -6766 46006
rect 26034 45918 26093 46000
rect 26174 45920 26233 46002
rect 26325 45919 26384 46001
rect -4954 45190 -4870 45266
rect -4949 45015 -4865 45091
rect 16282 45017 16382 45105
rect 16272 44819 16372 44907
rect -43938 44733 -43884 44795
rect -43941 44591 -43887 44653
rect -33957 44612 -33884 44672
rect -33959 44467 -33886 44527
rect -19373 44543 -19296 44610
rect -5125 44515 -5047 44578
rect -31905 44345 -31844 44415
rect -19373 44382 -19296 44449
rect -5129 44349 -5051 44412
rect -43630 44145 -43519 44256
rect -43378 44146 -43268 44255
rect -31915 44166 -31854 44236
rect -43380 43825 -43269 43936
rect -43132 43826 -43023 43935
rect -31577 43797 -31468 43906
rect -30930 43913 -30847 43996
rect -18962 44043 -18880 44132
rect -4168 44042 -4084 44126
rect -3928 44042 -3844 44126
rect 7031 44062 7083 44117
rect 7145 44063 7197 44118
rect -30928 43736 -30847 43817
rect -18963 43806 -18879 43890
rect 7834 43868 7910 43946
rect -31579 43581 -31468 43692
rect -18472 43750 -18363 43756
rect -18472 43647 -18361 43750
rect -4857 43647 -4748 43756
rect -18470 43641 -18361 43647
rect -4553 43646 -4437 43757
rect 7842 43684 7918 43762
rect -46580 43306 -46525 43362
rect -36274 43354 -36219 43410
rect -18472 43287 -18361 43398
rect -46374 43167 -46319 43223
rect -36068 43215 -36013 43271
rect -3921 43423 -3847 43497
rect -3920 43291 -3848 43363
rect -11227 43213 -11172 43269
rect -55281 42963 -55217 43044
rect -55133 42964 -55069 43045
rect -54984 42965 -54920 43046
rect -44931 42965 -44870 43039
rect -44782 42966 -44721 43040
rect -44635 42967 -44574 43041
rect -34690 43015 -34620 43092
rect -34537 43016 -34467 43093
rect -34392 43020 -34322 43097
rect -23387 42994 -23321 43076
rect -23244 42996 -23178 43078
rect -23090 42994 -23024 43076
rect -11021 43074 -10966 43130
rect -31579 42752 -31470 42863
rect -7135 42871 -7074 42951
rect -6989 42873 -6928 42953
rect -6840 42873 -6779 42953
rect 4840 42920 4920 43010
rect 4980 42930 5060 43020
rect 5120 42920 5200 43010
rect 15330 42872 15389 42943
rect 15464 42874 15523 42945
rect 15601 42874 15660 42945
rect 26028 42786 26087 42861
rect 26169 42791 26228 42866
rect 26323 42790 26382 42865
rect -31580 42514 -31469 42625
rect -4553 42552 -4442 42663
rect -4311 42553 -4202 42662
rect -65689 42425 -65623 42498
rect -65547 42428 -65481 42501
rect -65415 42429 -65349 42502
rect -55907 42015 -55849 42086
rect -55769 42019 -55711 42090
rect -55633 42023 -55575 42094
rect -45731 42075 -45679 42131
rect -45591 42083 -45539 42139
rect -45462 42074 -45410 42130
rect -24173 41947 -24121 42003
rect -24043 41960 -23991 42016
rect -23920 41947 -23868 42003
rect 4087 41939 4139 41995
rect 4208 41942 4260 41998
rect 4322 41942 4374 41998
rect 25353 41953 25413 42016
rect 25485 41956 25545 42019
rect 25619 41953 25679 42016
rect -66364 41703 -66303 41790
rect -66233 41703 -66172 41790
rect -66077 41697 -66016 41784
rect 14659 41843 14711 41899
rect 14802 41844 14854 41900
rect 14923 41848 14975 41904
rect -53175 41678 -53084 41757
rect -42854 41708 -42763 41787
rect -53179 41526 -53088 41605
rect -42858 41556 -42767 41635
rect -17805 41576 -17714 41655
rect 28811 41610 28902 41689
rect -17809 41424 -17718 41503
rect 7119 41487 7173 41541
rect 7232 41486 7288 41542
rect 16546 41459 16617 41532
rect 17858 41486 17949 41565
rect 28807 41458 28898 41537
rect 16541 41289 16612 41362
rect 17854 41334 17945 41413
rect -69407 41042 -69346 41107
rect -68334 41063 -68276 41115
rect -67788 41042 -67719 41107
rect -63590 40847 -63479 40954
rect -54168 40702 -54040 40754
rect -44003 40732 -43874 40786
rect -50858 40646 -50804 40700
rect -40552 40694 -40498 40748
rect -54168 40578 -54040 40630
rect -44003 40613 -43874 40667
rect -19690 40664 -19616 40738
rect -65678 40444 -65617 40529
rect -65549 40449 -65488 40534
rect -65389 40446 -65328 40531
rect -54167 40435 -54039 40487
rect -44004 40499 -43875 40553
rect -35369 40512 -35317 40568
rect -35248 40514 -35196 40570
rect -35099 40517 -35047 40573
rect -19689 40534 -19615 40608
rect -15505 40553 -15451 40607
rect 4855 40532 4907 40588
rect 4972 40539 5024 40595
rect 5089 40536 5141 40592
rect 27306 40558 27364 40613
rect -19689 40398 -19615 40472
rect -7900 40434 -7848 40490
rect -7768 40434 -7716 40490
rect -7647 40433 -7595 40489
rect 16299 40463 16363 40529
rect 16301 40325 16365 40391
rect 27311 40414 27369 40469
rect 27309 40288 27367 40343
rect 16289 40173 16353 40239
rect -66359 39919 -66299 40006
rect -66224 39915 -66164 40002
rect -66089 39914 -66029 40001
rect -55273 39650 -55215 39721
rect -55137 39652 -55079 39723
rect -54996 39653 -54938 39724
rect -44918 39694 -44866 39750
rect -44788 39694 -44736 39750
rect -44669 39696 -44617 39752
rect -23377 39551 -23325 39607
rect -23244 39557 -23192 39613
rect -23108 39557 -23056 39613
rect 6222 39631 6275 39694
rect -69513 39225 -69434 39299
rect -68433 39252 -68370 39315
rect -67893 39268 -67820 39335
rect -55280 39272 -55222 39343
rect -55144 39274 -55086 39345
rect -55003 39275 -54945 39346
rect -44908 39321 -44856 39377
rect -44778 39321 -44726 39377
rect -44659 39323 -44607 39379
rect -34694 39387 -34624 39464
rect -34544 39387 -34474 39464
rect -34393 39390 -34323 39467
rect 6223 39493 6276 39556
rect 16765 39564 16856 39643
rect 28481 39653 28572 39732
rect 16761 39412 16852 39491
rect 28477 39501 28568 39580
rect -23376 39183 -23324 39239
rect -23243 39189 -23191 39245
rect -23107 39189 -23055 39245
rect -63103 38910 -62992 39017
rect -65682 38659 -65622 38746
rect -65525 38658 -65465 38745
rect -65373 38667 -65313 38754
rect -66367 38343 -66304 38447
rect -66225 38344 -66162 38448
rect -66064 38346 -66001 38450
rect -53804 38344 -53741 38413
rect -43728 38400 -43673 38454
rect -43595 38405 -43540 38459
rect -33700 38443 -33645 38498
rect -33574 38443 -33519 38498
rect -53805 38184 -53742 38253
rect -50811 38139 -50756 38198
rect -40505 38187 -40450 38246
rect -18470 38775 -18359 38886
rect -18296 38776 -18187 38885
rect -9350 38670 -9270 38740
rect -9250 38550 -9170 38620
rect -18963 38247 -18879 38331
rect -18731 38247 -18647 38331
rect -34669 38069 -34617 38125
rect -34538 38075 -34486 38131
rect -34405 38077 -34353 38133
rect -15458 38046 -15403 38105
rect 4856 39181 4908 39237
rect 4973 39188 5025 39244
rect 5090 39185 5142 39241
rect 26049 39199 26109 39262
rect 26181 39202 26241 39265
rect 26315 39199 26375 39262
rect -5374 38372 -5322 38428
rect -5266 38374 -5214 38430
rect 15353 39116 15405 39172
rect 15470 39106 15522 39162
rect 15594 39110 15646 39166
rect 6437 38892 6512 38967
rect 6435 38721 6510 38796
rect 6674 38431 6766 38523
rect 6673 38251 6767 38345
rect -7122 37989 -7070 38045
rect -6991 37992 -6939 38048
rect -6870 37997 -6818 38053
rect -68507 37695 -68437 37774
rect -44930 37694 -44869 37768
rect -44795 37692 -44734 37766
rect -44645 37697 -44584 37771
rect -33290 37788 -33230 37845
rect -33157 37793 -33097 37850
rect -5049 37701 -4997 37753
rect -4936 37701 -4884 37753
rect 17013 38327 17105 38419
rect 17012 38166 17106 38260
rect 27946 38805 28014 38873
rect 28070 38806 28136 38872
rect 28308 38270 28383 38345
rect 28307 38120 28384 38197
rect -65682 37101 -65614 37192
rect -65528 37101 -65460 37192
rect -65375 37106 -65307 37197
rect -54477 36856 -54406 36947
rect -64629 36585 -64549 36665
rect -54487 36664 -54416 36755
rect -64628 36406 -64548 36486
rect -53800 36434 -53729 36507
rect -64379 36225 -64303 36297
rect -53806 36262 -53735 36335
rect -53242 36215 -53165 36287
rect -64380 36060 -64304 36132
rect -64121 36040 -64046 36119
rect -53246 36047 -53169 36119
rect -64126 35864 -64051 35943
rect 16285 35921 16365 35984
rect 6484 35709 6549 35767
rect 16281 35755 16361 35818
rect 6480 35582 6545 35640
rect 27309 35524 27388 35598
rect -4653 35377 -4575 35466
rect 27308 35341 27387 35415
rect -4654 35187 -4576 35276
rect -33992 34817 -33863 34871
rect 16585 34867 16649 34941
rect -33993 34704 -33864 34758
rect 16589 34723 16653 34797
rect -65680 34510 -65606 34610
rect -65534 34510 -65460 34610
rect -65386 34513 -65312 34613
rect -55284 34520 -55225 34595
rect -55156 34523 -55097 34598
rect -55027 34522 -54968 34597
rect -44928 34520 -44866 34593
rect -44802 34519 -44740 34592
rect -44647 34519 -44585 34592
rect -33992 34596 -33863 34650
rect -34693 34483 -34623 34572
rect -34545 34484 -34475 34573
rect -34401 34483 -34331 34572
rect -33999 34485 -33870 34539
rect -23382 34301 -23321 34379
rect -23242 34300 -23181 34378
rect -23081 34299 -23020 34377
rect -7133 34360 -7080 34435
rect -7003 34356 -6950 34431
rect -6869 34359 -6816 34434
rect 4841 34423 4906 34492
rect 4991 34423 5056 34492
rect 5137 34425 5202 34494
rect 15327 34362 15402 34439
rect 15478 34362 15553 34439
rect 15622 34363 15697 34440
rect 26028 34311 26101 34406
rect 26176 34311 26249 34406
rect 26330 34311 26403 34406
rect -66353 33586 -66293 33649
rect -66221 33589 -66161 33652
rect -66087 33586 -66027 33649
rect -55922 33577 -55854 33658
rect -55779 33577 -55711 33658
rect -55639 33581 -55571 33662
rect -45755 33548 -45685 33629
rect -45621 33547 -45551 33628
rect -45469 33549 -45399 33630
rect -35379 33357 -35309 33440
rect -35237 33361 -35167 33444
rect -35112 33365 -35042 33448
rect -24174 33412 -24104 33495
rect -24038 33414 -23968 33497
rect -23912 33418 -23842 33501
rect -7902 33474 -7848 33534
rect -7749 33482 -7695 33542
rect -7615 33492 -7561 33552
rect 4082 33421 4138 33485
rect 4220 33421 4276 33485
rect 4360 33420 4416 33484
rect 14655 33377 14707 33433
rect 14768 33381 14820 33437
rect 14881 33377 14933 33433
rect 25356 33446 25416 33509
rect 25488 33449 25548 33512
rect 25622 33446 25682 33509
rect -63356 33209 -63265 33288
rect -63360 33057 -63269 33136
rect -53184 33214 -53093 33293
rect -53188 33062 -53097 33141
rect -42790 33185 -42699 33264
rect -42794 33033 -42703 33112
rect -31731 33029 -31640 33108
rect -31735 32877 -31644 32956
rect -17916 33071 -17825 33150
rect -17920 32919 -17829 32998
rect -3954 33116 -3863 33195
rect -3958 32964 -3867 33043
rect 7022 33113 7113 33192
rect 17909 33116 18000 33195
rect 7018 32961 7109 33040
rect 16873 33000 16940 33071
rect 17905 32964 17996 33043
rect 28825 33116 28916 33195
rect 28821 32964 28912 33043
rect 16864 32817 16931 32888
rect -64642 32148 -64555 32263
rect -54170 32270 -54034 32327
rect -64637 31915 -64550 32030
rect -54169 32124 -54033 32181
rect -44000 32203 -43873 32262
rect -54169 32003 -54033 32060
rect -44001 32091 -43874 32150
rect -34001 32128 -33863 32194
rect -44004 31965 -43877 32024
rect -19684 32173 -19601 32255
rect -4661 32265 -4574 32351
rect -34006 31945 -33868 32011
rect -19685 31989 -19602 32071
rect -4663 32066 -4576 32152
rect 6477 32129 6543 32201
rect 6478 31972 6544 32044
rect 16584 32101 16661 32171
rect 27573 32083 27664 32161
rect 16583 31937 16660 32007
rect -34008 31796 -33870 31862
rect 27582 31876 27673 31954
rect -63769 31271 -63678 31350
rect -68318 31130 -68237 31187
rect -66690 31115 -66620 31186
rect -63773 31119 -63682 31198
rect -53483 31271 -53392 31350
rect -53487 31119 -53396 31198
rect -43109 31240 -43018 31319
rect -43113 31088 -43022 31167
rect -32035 31055 -31944 31134
rect -65679 30840 -65619 30903
rect -65547 30843 -65487 30906
rect -65413 30840 -65353 30903
rect -55272 30826 -55204 30907
rect -55127 30829 -55059 30910
rect -54990 30833 -54922 30914
rect -64374 29974 -64315 30033
rect -64376 29825 -64317 29884
rect -44932 30798 -44866 30871
rect -44805 30799 -44739 30872
rect -44651 30802 -44585 30875
rect -32039 30903 -31948 30982
rect -18207 31095 -18116 31174
rect -18211 30943 -18120 31022
rect -4250 31146 -4159 31225
rect -4254 30994 -4163 31073
rect 6710 31095 6801 31174
rect 28550 31150 28641 31229
rect 6706 30943 6797 31022
rect 17180 31040 17271 31119
rect 28546 30998 28637 31077
rect 17176 30888 17267 30967
rect -53884 29898 -53809 29973
rect -53884 29718 -53807 29795
rect -34681 30615 -34611 30698
rect -34550 30625 -34480 30708
rect -34422 30623 -34352 30706
rect -23377 30667 -23307 30750
rect -23227 30667 -23157 30750
rect -23091 30669 -23021 30752
rect -7140 30732 -7086 30792
rect -7002 30729 -6948 30789
rect -6869 30732 -6815 30792
rect -43708 29871 -43648 29932
rect -43596 29871 -43537 29932
rect -32283 29704 -32222 29770
rect -32106 29710 -32045 29776
rect -43389 29075 -43309 29155
rect -18470 30261 -18359 30372
rect -18285 30262 -18176 30371
rect -18963 29735 -18879 29819
rect -18763 29735 -18679 29819
rect 4839 30672 4895 30736
rect 4971 30675 5027 30739
rect 5127 30676 5183 30740
rect -4486 29824 -4402 29908
rect -4322 29825 -4240 29907
rect 15339 30634 15391 30690
rect 15459 30640 15511 30696
rect 15595 30640 15647 30696
rect 26049 30699 26109 30762
rect 26181 30702 26241 30765
rect 26315 30699 26375 30762
rect 6064 30256 6175 30367
rect 6367 30257 6476 30366
rect 6427 29735 6529 29837
rect 6631 29734 6735 29838
rect 17459 30238 17525 30304
rect 17458 30070 17526 30138
rect 17655 29701 17732 29778
rect 17646 29555 17724 29632
rect 27932 30469 28018 30555
rect 27936 30305 28024 30393
rect 28460 29773 28540 29848
rect 28462 29607 28539 29684
rect -43642 28887 -43560 28969
rect -43390 28905 -43308 28987
rect -43642 28677 -43560 28759
rect -32427 28667 -32317 28777
rect -32207 28666 -32095 28778
rect -4030 28631 -3919 28742
rect 17439 28741 17522 28824
rect 28754 28749 28820 28833
rect 17439 28590 17522 28677
rect 28756 28612 28822 28696
rect -18470 28421 -18359 28532
rect -18221 28421 -18110 28532
rect -4030 28422 -3921 28531
rect 6432 28367 6534 28469
rect 6658 28366 6762 28470
rect 18531 28356 18635 28460
rect 6064 28240 6175 28351
rect -4486 28086 -4402 28170
rect -18963 27922 -18879 28006
rect -18739 27922 -18655 28006
rect -4485 27923 -4403 28005
rect 18532 28175 18634 28277
rect 6065 27990 6174 28099
rect 17899 27925 18010 28036
rect 17900 27678 18009 27787
rect 27567 27714 27650 27809
rect -19700 27552 -19604 27625
rect -19696 27385 -19600 27458
rect -5692 27405 -5591 27486
rect 27571 27481 27654 27576
rect -5692 27170 -5591 27251
rect 28462 27197 28557 27292
rect 17631 27137 17724 27140
rect 17630 27042 17725 27137
rect 28463 27043 28556 27136
rect 17630 26875 17725 26970
rect -9349 26695 -9295 26761
rect -9213 26698 -9159 26764
rect -64367 26530 -64313 26583
rect -64368 26423 -64314 26476
rect -64370 26315 -64316 26368
rect -53886 26443 -53814 26515
rect -53886 26307 -53814 26379
rect -55284 26129 -55214 26230
rect -55150 26126 -55080 26227
rect -55004 26128 -54934 26229
rect -44927 26054 -44861 26144
rect -44783 26052 -44717 26142
rect -44645 26054 -44579 26144
rect -34687 26063 -34625 26138
rect -34553 26060 -34491 26135
rect -34391 26065 -34329 26140
rect -33703 26061 -33631 26133
rect -33502 26060 -33428 26134
rect 15331 26365 15402 26441
rect 15484 26365 15555 26441
rect 15637 26362 15708 26438
rect -5373 26288 -5301 26360
rect -5197 26287 -5123 26361
rect 28178 26376 28295 26493
rect 28441 26375 28560 26494
rect -7904 26147 -7852 26200
rect -7764 26152 -7712 26205
rect -7615 26158 -7563 26211
rect 26025 26087 26084 26162
rect 26165 26090 26224 26165
rect 26312 26090 26371 26165
rect -9399 25907 -9345 25961
rect -9271 25909 -9215 25965
rect 4846 25923 4915 26021
rect 4986 25922 5055 26020
rect 5134 25927 5203 26025
rect -64112 25813 -64054 25870
rect -64113 25701 -64055 25758
rect -53594 25717 -53536 25775
rect -53446 25723 -53388 25781
rect -23387 25670 -23311 25782
rect -23236 25673 -23160 25785
rect -23087 25675 -23011 25787
rect -9399 25793 -9343 25849
rect -9269 25800 -9215 25854
rect 17897 25855 18006 25964
rect -64114 25588 -64056 25645
rect 17896 25639 18007 25750
rect 28588 25815 28697 25924
rect -7118 25450 -7066 25503
rect -6985 25450 -6933 25503
rect -6844 25445 -6792 25498
rect 28587 25543 28698 25654
rect 4084 25427 4150 25493
rect 4224 25430 4290 25496
rect 4374 25433 4440 25499
rect -45746 25127 -45674 25205
rect -45608 25128 -45536 25206
rect -45474 25128 -45402 25206
rect -24150 25180 -24060 25270
rect -23920 25186 -23829 25270
rect 7059 25063 7150 25142
rect 7055 24911 7146 24990
rect -43004 24774 -42913 24853
rect -43008 24622 -42917 24701
rect -18615 24812 -18524 24891
rect -18619 24660 -18528 24739
rect -5043 24119 -4932 24230
rect -4794 24120 -4685 24229
rect 5684 24044 5737 24101
rect -32950 23892 -32839 24003
rect -32723 23893 -32614 24002
rect 5571 23978 5624 24035
rect 5678 23891 5731 23948
rect -66363 23657 -66303 23720
rect -66231 23660 -66171 23723
rect -66097 23657 -66037 23720
rect -43648 23694 -43539 23806
rect -55922 23572 -55864 23630
rect -55787 23575 -55729 23633
rect -55653 23578 -55595 23636
rect -43656 23457 -43547 23569
rect -19606 23758 -19517 23815
rect 5574 23813 5627 23870
rect -19605 23638 -19516 23695
rect 14654 23617 14706 23673
rect 14782 23616 14834 23672
rect 14921 23615 14973 23671
rect -19606 23529 -19517 23586
rect 25348 23548 25408 23611
rect 25480 23551 25540 23614
rect 25614 23548 25674 23611
rect -7897 23429 -7845 23486
rect -7776 23433 -7724 23490
rect -7640 23436 -7588 23493
rect -35376 23200 -35316 23260
rect -35240 23201 -35180 23261
rect -35086 23201 -35026 23261
rect 6728 23132 6819 23211
rect 6724 22980 6815 23059
rect -68348 22714 -68263 22803
rect -66681 22748 -66602 22822
rect -43303 22834 -43212 22913
rect -43307 22682 -43216 22761
rect -19029 22886 -18938 22965
rect -19033 22734 -18942 22813
rect 4847 22675 4911 22737
rect 4991 22676 5055 22738
rect 5132 22677 5196 22739
rect -44926 22381 -44874 22437
rect -44806 22383 -44754 22439
rect -44681 22385 -44629 22441
rect -23365 22436 -23275 22526
rect -23124 22440 -23034 22530
rect -65672 21228 -65612 21291
rect -65540 21231 -65480 21294
rect -65406 21228 -65346 21291
rect -67592 21081 -67502 21171
rect -66912 21082 -66824 21170
rect -53361 21507 -53306 21562
rect -53250 21507 -53195 21562
rect -55278 21137 -55223 21192
rect -55145 21138 -55090 21193
rect -54999 21140 -54944 21195
rect -53876 20935 -53821 20990
rect -53875 20802 -53820 20857
rect -53675 20669 -53620 20724
rect -53674 20536 -53619 20591
rect -32602 21148 -32550 21201
rect -32487 21141 -32435 21194
rect -19197 21499 -19131 21571
rect -18989 21503 -18923 21575
rect -4813 21344 -4751 21408
rect -4636 21349 -4574 21413
rect 6085 22281 6151 22347
rect 6084 22124 6152 22192
rect 6426 21720 6530 21824
rect 6637 21721 6739 21823
rect 17650 21545 17705 21600
rect 17790 21544 17847 21601
rect 28493 21483 28548 21538
rect 28493 21364 28548 21419
rect 15336 21172 15388 21228
rect 15443 21176 15495 21232
rect 15568 21172 15620 21228
rect 26042 21114 26102 21177
rect 26174 21117 26234 21180
rect 26308 21114 26368 21177
rect -7120 21000 -7064 21054
rect -6990 21000 -6934 21054
rect -6859 21004 -6803 21058
rect -34682 20762 -34623 20824
rect -34543 20765 -34484 20827
rect -34399 20769 -34340 20831
rect 6064 20907 6175 21019
rect -33690 20590 -33630 20650
rect -53173 20481 -53113 20538
rect -53058 20481 -52998 20538
rect -33690 20450 -33630 20510
rect 6064 20679 6175 20793
rect -33230 20470 -33170 20530
rect -52583 20279 -52523 20336
rect -52468 20279 -52408 20336
rect -43080 20239 -42969 20350
rect -42887 20238 -42774 20351
rect -33230 20350 -33170 20410
rect -22292 20463 -22216 20530
rect -22103 20466 -22027 20533
rect 6426 20480 6530 20584
rect 28464 20422 28573 20531
rect 28713 20422 28822 20531
rect 6427 20244 6529 20346
rect -32610 20175 -32558 20228
rect -32446 20178 -32394 20231
rect -21949 20112 -21873 20179
rect -21783 20112 -21707 20179
rect -4796 20124 -4740 20177
rect -4649 20122 -4593 20175
rect -18824 19761 -18767 19817
rect -18672 19764 -18615 19820
rect -5026 19668 -4954 19748
rect 18278 19729 18412 19863
rect 18527 19728 18663 19864
rect -19098 19420 -19041 19476
rect -18946 19423 -18889 19479
rect -5347 19458 -5275 19538
rect -5023 19467 -4951 19547
rect 17656 19459 17738 19539
rect -5344 19245 -5272 19325
rect 17656 19287 17738 19367
rect -19604 19093 -19511 19199
rect 5587 19116 5719 19200
rect -19603 18954 -19508 19022
rect -54148 18808 -54063 18875
rect -19596 18769 -19505 18859
rect -54150 18635 -54048 18744
rect -54158 18396 -54056 18505
rect 5591 18962 5723 19046
rect -43384 18322 -43283 18423
rect -43367 18130 -43266 18231
rect -43377 17955 -43276 18056
rect -64639 17820 -64565 17925
rect -64633 17603 -64559 17708
rect 27251 17660 27369 17778
rect -43887 17498 -43780 17557
rect -43883 17371 -43776 17430
rect -44933 17229 -44868 17307
rect -44796 17227 -44731 17305
rect -44650 17227 -44585 17305
rect -43886 17248 -43779 17307
rect -65684 16946 -65623 17029
rect -65523 16951 -65462 17034
rect -65391 16946 -65330 17029
rect -55282 16945 -55223 17034
rect -55138 16946 -55079 17035
rect -54982 16945 -54923 17034
rect 5770 17386 5852 17462
rect 27246 17425 27364 17543
rect 5773 17220 5855 17296
rect -23382 17074 -23325 17158
rect -23236 17072 -23179 17156
rect -23091 17079 -23034 17163
rect 5779 17052 5861 17128
rect -34687 16892 -34625 16969
rect -34540 16891 -34478 16968
rect -34391 16893 -34329 16970
rect -7137 16935 -7066 17016
rect -6987 16938 -6916 17019
rect -6831 16933 -6760 17014
rect 4841 16940 4898 17011
rect 4961 16940 5018 17011
rect 5081 16941 5138 17012
rect 15334 16842 15388 16920
rect 15475 16839 15529 16917
rect 15626 16838 15680 16916
rect 26025 16873 26082 16946
rect 26180 16878 26237 16951
rect 26319 16881 26376 16954
rect -55926 16288 -55850 16379
rect -55784 16287 -55708 16378
rect -55633 16288 -55557 16379
rect -35367 16144 -35314 16200
rect -35217 16145 -35164 16201
rect -35081 16150 -35028 16206
rect -66363 16015 -66303 16078
rect -66231 16018 -66171 16081
rect -66097 16015 -66037 16078
rect -53166 15877 -53110 15933
rect -45752 15951 -45682 16037
rect -45608 15950 -45538 16036
rect -45479 15950 -45409 16036
rect -7892 16014 -7830 16077
rect -7758 16014 -7696 16077
rect -7622 16015 -7560 16078
rect -53170 15766 -53114 15822
rect -20770 15816 -20644 15941
rect -20524 15815 -20397 15942
rect 4083 15914 4144 15980
rect 4230 15913 4291 15979
rect 4372 15916 4433 15982
rect 14661 15934 14713 15990
rect 14775 15934 14827 15990
rect 14896 15937 14948 15993
rect 25348 15922 25408 15985
rect 25480 15925 25540 15988
rect 25614 15922 25674 15985
rect -63321 15647 -63265 15703
rect -32593 15704 -32537 15760
rect -63325 15536 -63269 15592
rect -42963 15566 -42907 15622
rect -32597 15593 -32541 15649
rect -3755 15612 -3699 15668
rect -42967 15455 -42911 15511
rect -3759 15501 -3703 15557
rect 6890 15526 6946 15582
rect 6886 15415 6942 15471
rect 17953 15536 18009 15592
rect 17949 15425 18005 15481
rect 28864 15529 28920 15585
rect 28860 15418 28916 15474
rect -54097 14901 -54033 14968
rect -64608 14668 -64544 14728
rect -54100 14728 -54036 14795
rect -33934 14760 -33866 14830
rect -64607 14500 -64543 14560
rect -43866 14559 -43794 14626
rect -33934 14584 -33866 14654
rect -5653 14602 -5582 14669
rect -43869 14367 -43797 14434
rect -5658 14426 -5587 14493
rect 5833 14431 5892 14497
rect 17004 14511 17059 14566
rect 26063 14534 26123 14597
rect 26195 14537 26255 14600
rect 26329 14534 26389 14597
rect 17000 14369 17055 14424
rect 5826 14252 5885 14318
rect -53461 13979 -53405 14035
rect -24175 14008 -24069 14094
rect -23950 14010 -23844 14096
rect -53465 13868 -53409 13924
rect -32931 13796 -32875 13852
rect -68333 13646 -68258 13716
rect -66686 13646 -66620 13709
rect -63611 13707 -63555 13763
rect -63615 13596 -63559 13652
rect -55278 13540 -55202 13631
rect -55146 13538 -55070 13629
rect -55006 13538 -54930 13629
rect -32935 13685 -32879 13741
rect -65672 13272 -65612 13335
rect -65540 13275 -65480 13338
rect -65406 13272 -65346 13335
rect -72089 12672 -72035 12726
rect -71966 12672 -71912 12726
rect -71988 12268 -71900 12356
rect -71829 12268 -71741 12356
rect -73140 12012 -72991 12147
rect -72885 12014 -72736 12149
rect -66370 11976 -66308 12048
rect -66255 11976 -66193 12048
rect -66141 11976 -66079 12048
rect -71203 11635 -71142 11733
rect -71142 11635 -71104 11733
rect -64372 12389 -64311 12450
rect -64373 12254 -64312 12315
rect -4098 13685 -4042 13741
rect -43268 13608 -43212 13664
rect -4102 13574 -4046 13630
rect 6644 13674 6700 13730
rect 6640 13563 6696 13619
rect -43272 13497 -43216 13553
rect 17640 13644 17696 13700
rect -34685 13394 -34630 13447
rect -34546 13393 -34491 13446
rect -34400 13395 -34345 13448
rect -23387 13448 -23320 13526
rect -23242 13453 -23175 13531
rect -23103 13451 -23036 13529
rect 17636 13533 17692 13589
rect 28540 13667 28596 13723
rect 28536 13556 28592 13612
rect -44931 13207 -44876 13271
rect -44810 13211 -44755 13275
rect -44679 13212 -44624 13276
rect -53885 12773 -53808 12850
rect -53885 12612 -53810 12687
rect -71203 11634 -71104 11635
rect -71185 11486 -71100 11580
rect -43377 12274 -43302 12349
rect -43224 12274 -43149 12349
rect -53255 11794 -53197 11852
rect -33718 12438 -33607 12549
rect -33410 12438 -33299 12549
rect -53254 11660 -53198 11716
rect -34688 11614 -34621 11705
rect -34545 11614 -34478 11705
rect -34416 11618 -34349 11709
rect -23383 11703 -23316 11794
rect -23227 11701 -23160 11792
rect -23095 11701 -23028 11792
rect -43482 11435 -43398 11519
rect -43278 11434 -43192 11520
rect -71904 11197 -71787 11310
rect -71610 11194 -71493 11307
rect -71907 10899 -71790 11012
rect -71617 10899 -71500 11012
rect -66361 10387 -66308 10443
rect -66251 10387 -66198 10443
rect -66095 10388 -66042 10444
rect -35373 10339 -35318 10392
rect -35242 10339 -35187 10392
rect -35095 10345 -35040 10398
rect -65679 9701 -65626 9757
rect -65534 9705 -65481 9761
rect -65402 9707 -65349 9763
rect -34690 9639 -34635 9692
rect -34560 9642 -34505 9695
rect -34411 9640 -34356 9693
rect -66359 9471 -66306 9527
rect -66231 9470 -66178 9526
rect -66110 9472 -66057 9528
rect -35378 9447 -35323 9500
rect -35239 9452 -35184 9505
rect -35101 9453 -35046 9506
rect -65671 8784 -65618 8840
rect -65529 8788 -65476 8844
rect -65391 8787 -65338 8843
rect -34687 8747 -34632 8800
rect -34542 8751 -34487 8804
rect -34412 8749 -34357 8802
rect -66360 8561 -66307 8617
rect -66224 8563 -66171 8619
rect -66077 8565 -66024 8621
rect -35372 8502 -35317 8555
rect -35249 8509 -35194 8562
rect -35117 8513 -35062 8566
rect -65672 7861 -65619 7917
rect -65538 7863 -65485 7919
rect -65388 7865 -65335 7921
rect -34683 7804 -34628 7857
rect -34544 7805 -34489 7858
rect -34398 7805 -34343 7858
rect -66357 7640 -66304 7696
rect -66199 7647 -66146 7703
rect -66063 7645 -66010 7701
rect -35382 7618 -35327 7671
rect -35256 7625 -35201 7678
rect -35125 7632 -35070 7685
rect -65673 6966 -65620 7022
rect -65554 6976 -65501 7032
rect -65408 6976 -65355 7032
rect -34685 6931 -34630 6984
rect -34552 6932 -34497 6985
rect -34416 6938 -34361 6991
rect -66365 6730 -66312 6786
rect -66232 6736 -66179 6792
rect -66090 6737 -66037 6793
rect -35371 6712 -35316 6765
rect -35244 6717 -35189 6770
rect -35117 6716 -35062 6769
rect -18261 9776 -18209 9828
rect -18155 9774 -18095 9826
rect -7130 13249 -7077 13305
rect -7011 13251 -6958 13307
rect -6894 13253 -6841 13309
rect 4848 13151 4910 13215
rect 4981 13156 5043 13220
rect 5121 13156 5183 13220
rect 15341 13180 15393 13236
rect 15459 13182 15511 13238
rect 15595 13189 15647 13245
rect 26055 13179 26115 13242
rect 26187 13182 26247 13245
rect 26321 13179 26381 13242
rect 6064 12721 6175 12849
rect 27828 12783 27894 12849
rect 6065 12543 6174 12652
rect 27828 12628 27894 12694
rect -4360 12342 -4303 12405
rect -4183 12350 -4126 12413
rect 6254 12199 6356 12301
rect 6426 12198 6530 12302
rect 17365 12257 17441 12332
rect 17522 12256 17599 12333
rect 28119 12251 28194 12326
rect 28118 12075 28195 12152
rect -7136 11601 -7068 11700
rect -6988 11607 -6920 11706
rect -6843 11599 -6775 11698
rect 4843 11605 4904 11693
rect 4983 11606 5044 11694
rect 5124 11600 5185 11688
rect 15340 11452 15394 11530
rect 15493 11453 15547 11531
rect 15626 11444 15680 11522
rect 26033 11448 26090 11521
rect 26173 11453 26230 11526
rect 26325 11452 26382 11525
rect -7125 9144 -7059 9226
rect -6984 9148 -6918 9230
rect -6832 9151 -6766 9233
rect -23371 8718 -23304 8792
rect -23225 8725 -23158 8799
rect -23080 8725 -23013 8799
rect -23370 8572 -23303 8646
rect -23220 8576 -23153 8650
rect -23077 8584 -23010 8658
rect -23367 8400 -23280 8494
rect -23116 8404 -23029 8498
rect -24167 7738 -24080 7832
rect -23917 7738 -23830 7832
rect -65664 6033 -65611 6089
rect -65539 6035 -65486 6091
rect -65403 6037 -65350 6093
rect -34686 6017 -34631 6070
rect -34545 6020 -34490 6073
rect -34403 6022 -34348 6075
rect -66355 5812 -66302 5868
rect -66221 5809 -66168 5865
rect -66084 5810 -66031 5866
rect -35369 5799 -35314 5852
rect -35243 5805 -35188 5858
rect -35103 5803 -35048 5856
rect -65678 5119 -65625 5175
rect -65537 5122 -65484 5178
rect -65390 5122 -65337 5178
rect -34679 5105 -34624 5158
rect -34551 5106 -34496 5159
rect -34400 5107 -34345 5160
rect -55285 4641 -55229 4715
rect -55124 4646 -55068 4720
rect -54966 4654 -54910 4728
rect -44929 4302 -44877 4377
rect -44798 4304 -44746 4379
rect -44652 4299 -44600 4374
rect -34680 4077 -34610 4165
rect -34544 4073 -34474 4161
rect -34392 4079 -34322 4167
rect 15344 4463 15396 4519
rect 15472 4463 15524 4519
rect 15584 4466 15636 4522
rect 4842 4259 4897 4328
rect 4990 4263 5045 4332
rect 5142 4269 5197 4338
rect 26031 4336 26099 4406
rect 26174 4341 26242 4411
rect 26319 4351 26387 4421
rect 26032 4193 26100 4263
rect 26176 4193 26244 4263
rect 26327 4196 26395 4266
rect -34685 3889 -34615 3977
rect -34528 3896 -34458 3984
rect -34388 3896 -34318 3984
rect -7124 3962 -7056 4059
rect -6971 3962 -6903 4059
rect -6827 3962 -6759 4059
rect -66353 3709 -66293 3772
rect -66221 3712 -66161 3775
rect -66087 3709 -66027 3772
rect -7135 3761 -7067 3858
rect -6970 3758 -6902 3855
rect -6826 3765 -6758 3862
rect -23380 3616 -23325 3684
rect -23241 3621 -23186 3689
rect -23100 3624 -23045 3692
rect 4084 3529 4156 3599
rect 4235 3529 4307 3599
rect 4360 3531 4432 3601
rect -63329 3324 -63273 3380
rect -55918 3358 -55853 3435
rect -55783 3358 -55718 3435
rect -55642 3362 -55577 3439
rect -23388 3430 -23333 3498
rect -23244 3435 -23189 3503
rect -23086 3435 -23031 3503
rect -63333 3213 -63277 3269
rect -7895 3317 -7828 3390
rect -7746 3319 -7679 3392
rect -7610 3321 -7543 3394
rect 14651 3400 14703 3456
rect 14798 3407 14850 3463
rect 14923 3412 14975 3468
rect -45753 3138 -45681 3212
rect -45618 3138 -45546 3212
rect -45473 3140 -45401 3214
rect -35368 3228 -35314 3284
rect -35226 3231 -35172 3287
rect -35080 3232 -35026 3288
rect 7116 3112 7172 3168
rect 25354 3185 25414 3248
rect 25486 3188 25546 3251
rect 25620 3185 25680 3248
rect -53194 2993 -53138 3049
rect 7112 3001 7168 3057
rect -53198 2882 -53142 2938
rect 17962 3032 18018 3088
rect -3707 2919 -3651 2975
rect 17958 2921 18014 2977
rect -42778 2760 -42722 2816
rect -42782 2649 -42726 2705
rect -32474 2762 -32418 2818
rect -3711 2808 -3655 2864
rect -32478 2651 -32422 2707
rect 28622 2807 28678 2863
rect -24146 2659 -24088 2736
rect -24005 2665 -23947 2742
rect -23866 2669 -23808 2746
rect 28618 2696 28674 2752
rect -24173 2484 -24115 2561
rect -24014 2491 -23956 2568
rect -23870 2489 -23812 2566
rect -64601 2391 -64545 2456
rect -64600 2228 -64544 2293
rect 5832 2266 5896 2335
rect -54104 2098 -54036 2167
rect -66367 1926 -66301 2021
rect -66223 1932 -66157 2027
rect -66064 1932 -65998 2027
rect -54106 1957 -54038 2026
rect 5831 2100 5895 2169
rect 17002 2151 17058 2211
rect -43868 1888 -43800 1951
rect -33928 1971 -33868 2041
rect -5650 2008 -5581 2080
rect 16999 1976 17055 2036
rect -33928 1808 -33868 1878
rect -5656 1835 -5587 1907
rect -43869 1723 -43801 1786
rect -63742 1354 -63686 1410
rect -63746 1243 -63690 1299
rect -68328 1064 -68246 1157
rect -66723 1083 -66653 1148
rect -65662 959 -65602 1022
rect -65530 962 -65470 1025
rect -65396 959 -65336 1022
rect -53627 1038 -53571 1094
rect -53631 927 -53575 983
rect -43134 851 -43078 907
rect -55280 608 -55215 685
rect -55150 613 -55085 690
rect -54997 616 -54932 693
rect -43138 740 -43082 796
rect -65682 423 -65622 502
rect -65546 423 -65486 502
rect -65402 425 -65342 504
rect -44930 389 -44864 449
rect -44809 388 -44743 448
rect -44679 389 -44613 449
rect -64360 183 -64306 240
rect -64364 36 -64310 93
rect -53994 -316 -53919 -241
rect -53826 -316 -53749 -239
rect -43346 -544 -43271 -469
rect -43184 -545 -43107 -468
rect -65671 -808 -65594 -695
rect -65518 -801 -65441 -688
rect -65385 -797 -65308 -684
rect -55282 -770 -55225 -693
rect -55151 -770 -55094 -693
rect -55022 -771 -54965 -694
rect -44917 -969 -44861 -879
rect -44782 -967 -44726 -877
rect -44631 -965 -44575 -875
rect -43474 -1076 -43417 -1017
rect -54003 -1205 -53937 -1146
rect -43473 -1199 -43416 -1140
rect -43282 -1204 -43229 -1149
rect -54005 -1321 -53939 -1262
rect -43281 -1314 -43228 -1259
rect -53743 -1390 -53678 -1330
rect -53742 -1506 -53677 -1446
rect 26066 1792 26126 1855
rect 26198 1795 26258 1858
rect 26332 1792 26392 1855
rect 6772 1210 6828 1266
rect 6768 1099 6824 1155
rect 17577 1092 17633 1148
rect -32833 911 -32777 967
rect -4071 984 -4015 1040
rect 17573 981 17629 1037
rect -4075 873 -4019 929
rect -32837 800 -32781 856
rect 4848 781 4910 841
rect 4977 784 5039 844
rect 5110 784 5172 844
rect 15350 774 15402 830
rect 15478 774 15530 830
rect 15590 777 15642 833
rect 28348 895 28404 951
rect -34686 474 -34632 527
rect -34529 475 -34475 528
rect -34398 478 -34344 531
rect -7126 568 -7065 636
rect -6980 570 -6919 638
rect -6841 570 -6780 638
rect 15351 663 15403 719
rect 15479 663 15531 719
rect 15591 666 15643 722
rect 28344 784 28400 840
rect 26055 442 26115 505
rect 26187 445 26247 508
rect 26321 442 26381 505
rect 27820 43 27888 111
rect -23386 -193 -23332 -125
rect -23235 -194 -23181 -126
rect -23092 -191 -23038 -123
rect -18813 -223 -18748 -138
rect -18638 -223 -18573 -138
rect -33186 -470 -33077 -361
rect -32936 -472 -32825 -361
rect -4368 -378 -4230 -240
rect -4045 -377 -3909 -241
rect -34687 -1281 -34614 -1181
rect -34536 -1283 -34463 -1183
rect -34391 -1271 -34318 -1171
rect -23389 -1202 -23334 -1134
rect -23254 -1200 -23199 -1132
rect -23103 -1195 -23048 -1127
rect 4847 -1153 4902 -1084
rect 4997 -1152 5052 -1083
rect 5158 -1147 5213 -1078
rect -23392 -1342 -23337 -1274
rect -23251 -1340 -23196 -1272
rect -23104 -1339 -23049 -1271
rect -7133 -1293 -7071 -1214
rect -6989 -1291 -6927 -1212
rect -6857 -1292 -6795 -1213
rect 27821 -141 27887 -75
rect 16703 -270 16778 -195
rect 16702 -486 16779 -409
rect 28121 -493 28197 -418
rect 15332 -733 15395 -658
rect 15474 -737 15537 -662
rect 15606 -731 15669 -656
rect 28118 -640 28195 -563
rect 17013 -765 17091 -688
rect 17018 -929 17096 -852
rect 26033 -898 26100 -799
rect 26183 -894 26250 -795
rect 26319 -892 26386 -793
rect 16700 -1323 16778 -1246
rect 16705 -1487 16783 -1410
rect -43764 -3122 -43673 -2965
rect -54337 -3396 -54234 -3259
rect -43772 -3402 -43681 -3245
rect -54346 -3648 -54243 -3511
rect -64576 -3793 -64498 -3659
rect -64578 -3995 -64500 -3861
rect -3711 -3993 -3659 -3940
rect -3584 -3990 -3532 -3937
rect -19319 -4110 -19229 -4020
rect -33023 -4292 -32873 -4142
rect -32705 -4291 -32557 -4143
rect -21964 -4262 -21877 -4186
rect -21740 -4255 -21653 -4179
rect -19319 -4274 -19229 -4184
rect -54002 -4476 -53930 -4404
rect -18823 -4422 -18735 -4334
rect -54003 -4627 -53929 -4553
rect -22308 -4655 -22221 -4579
rect -22080 -4650 -21993 -4574
rect -18823 -4603 -18735 -4515
rect 16703 -4437 16775 -4365
rect 28133 -4488 28197 -4423
rect 28315 -4491 28379 -4426
rect -65684 -4911 -65618 -4832
rect -65551 -4908 -65485 -4829
rect -65400 -4903 -65334 -4824
rect -65686 -5048 -65620 -4969
rect -65541 -5048 -65475 -4969
rect -65393 -5047 -65327 -4968
rect -55281 -4852 -55224 -4781
rect -55137 -4854 -55080 -4783
rect -54975 -4848 -54918 -4777
rect -44927 -4851 -44863 -4754
rect -44778 -4851 -44714 -4754
rect -44630 -4851 -44566 -4754
rect 16702 -4602 16776 -4528
rect 26022 -4824 26093 -4746
rect 26177 -4825 26248 -4747
rect 26330 -4828 26401 -4750
rect -55283 -5015 -55226 -4944
rect -55139 -5016 -55082 -4945
rect -54971 -5011 -54914 -4940
rect -7128 -4980 -7073 -4925
rect -6992 -4979 -6937 -4924
rect -6838 -4980 -6783 -4925
rect 4843 -5001 4922 -4899
rect 4993 -5002 5072 -4900
rect 5139 -5001 5218 -4899
rect -53741 -5186 -53685 -5128
rect -53571 -5185 -53515 -5127
rect -34685 -5193 -34621 -5126
rect -34531 -5190 -34467 -5123
rect -34397 -5192 -34333 -5125
rect -23384 -5192 -23313 -5119
rect -23227 -5197 -23156 -5124
rect -23074 -5201 -23003 -5128
rect 15330 -5084 15396 -5013
rect 15462 -5080 15528 -5009
rect 15623 -5083 15689 -5012
rect -3552 -5228 -3500 -5175
rect 17262 -5135 17318 -5077
rect 17380 -5141 17436 -5083
rect 17541 -5134 17597 -5076
rect 27820 -5031 27892 -4956
rect 15328 -5269 15394 -5198
rect 15478 -5271 15544 -5200
rect 15632 -5267 15698 -5196
rect 27815 -5208 27887 -5133
rect -3566 -5343 -3514 -5290
rect -33042 -5434 -32987 -5379
rect -33041 -5545 -32986 -5490
rect -66356 -5804 -66296 -5741
rect -66224 -5801 -66164 -5738
rect -66090 -5804 -66030 -5741
rect -45752 -5826 -45687 -5764
rect -45614 -5825 -45549 -5763
rect -45478 -5823 -45413 -5761
rect -24154 -5943 -24071 -5858
rect -23919 -5940 -23836 -5855
rect 4082 -6052 4161 -5979
rect 4231 -6053 4310 -5980
rect 4369 -6050 4448 -5977
rect -63338 -6178 -63282 -6122
rect -63342 -6289 -63286 -6233
rect -42799 -6203 -42743 -6147
rect -42803 -6314 -42747 -6258
rect -19334 -6239 -19278 -6183
rect -19338 -6350 -19282 -6294
rect 7099 -6426 7155 -6370
rect 7095 -6537 7151 -6481
rect -66367 -7181 -66302 -7093
rect -66225 -7176 -66160 -7088
rect -66070 -7172 -66005 -7084
rect -64572 -7205 -64513 -7141
rect -43750 -7205 -43682 -7123
rect -20561 -7249 -20476 -7178
rect -64575 -7373 -64516 -7309
rect -55922 -7329 -55865 -7277
rect -55794 -7325 -55737 -7273
rect -55668 -7324 -55611 -7272
rect -43750 -7397 -43682 -7315
rect 14647 -7294 14699 -7238
rect 14766 -7293 14818 -7237
rect 14900 -7292 14952 -7236
rect -20563 -7390 -20478 -7319
rect -7898 -7410 -7838 -7344
rect -7743 -7411 -7683 -7345
rect -7610 -7411 -7550 -7345
rect 25354 -7346 25414 -7283
rect 25486 -7343 25546 -7280
rect 25620 -7346 25680 -7283
rect -20568 -7529 -20483 -7458
rect 4869 -7438 4926 -7384
rect 4996 -7437 5053 -7383
rect 5123 -7433 5180 -7379
rect -35376 -7616 -35316 -7554
rect -35231 -7616 -35171 -7554
rect -35076 -7614 -35016 -7552
rect -68368 -8020 -68292 -7945
rect -66691 -8026 -66618 -7948
rect -64327 -8086 -64270 -8080
rect -64331 -8135 -64270 -8086
rect -43097 -8116 -43015 -8034
rect -64331 -8142 -64275 -8135
rect -64335 -8206 -64279 -8197
rect -64335 -8253 -64277 -8206
rect -64334 -8261 -64277 -8253
rect -43097 -8281 -43015 -8199
rect -19850 -8314 -19768 -8232
rect -19685 -8314 -19603 -8232
rect -65665 -8547 -65605 -8484
rect -65533 -8544 -65473 -8481
rect -65399 -8547 -65339 -8484
rect -55285 -8495 -55233 -8429
rect -55149 -8498 -55097 -8432
rect -54987 -8493 -54935 -8427
rect 6473 -8410 6555 -8328
rect 6638 -8410 6720 -8328
rect -44930 -8579 -44874 -8518
rect -44795 -8578 -44739 -8517
rect -44654 -8576 -44598 -8515
rect -34692 -8512 -34629 -8447
rect -34553 -8510 -34490 -8445
rect -34397 -8512 -34334 -8447
rect -23378 -8703 -23292 -8618
rect -23115 -8698 -23029 -8613
rect -7135 -8631 -7074 -8565
rect -6998 -8631 -6937 -8565
rect -6841 -8623 -6780 -8557
rect 4846 -8801 4903 -8747
rect 4973 -8800 5030 -8746
rect 5100 -8796 5157 -8742
rect 15330 -8736 15384 -8676
rect 15461 -8736 15515 -8676
rect 15602 -8738 15656 -8678
rect -64126 -8970 -64070 -8908
rect -64125 -9110 -64069 -9048
rect -63872 -9471 -63818 -9417
rect -53466 -9399 -53411 -9344
rect -53323 -9399 -53268 -9344
rect 17316 -9361 17373 -9304
rect 17437 -9359 17492 -9304
rect -43466 -9502 -43414 -9445
rect -43341 -9503 -43289 -9446
rect 28516 -9416 28573 -9359
rect -63873 -9601 -63819 -9547
rect -55274 -9767 -55203 -9703
rect -55134 -9768 -55063 -9704
rect -54991 -9772 -54920 -9708
rect -44928 -9791 -44868 -9712
rect -44788 -9785 -44728 -9706
rect -44634 -9785 -44574 -9706
rect -33319 -9785 -33208 -9674
rect -33092 -9784 -32981 -9675
rect -65680 -10247 -65618 -10171
rect -65539 -10247 -65477 -10171
rect -65389 -10243 -65327 -10167
rect -23386 -10132 -23315 -10059
rect -23233 -10135 -23162 -10062
rect -23078 -10135 -23007 -10062
rect -34688 -10255 -34632 -10172
rect -34544 -10259 -34488 -10176
rect -34394 -10248 -34338 -10165
rect -4065 -9571 -3984 -9481
rect -3827 -9561 -3746 -9471
rect 28518 -9543 28577 -9484
rect 4844 -9932 4899 -9858
rect 4983 -9934 5038 -9860
rect 5133 -9930 5188 -9856
rect -7136 -10276 -7081 -10198
rect -7002 -10275 -6947 -10197
rect -6861 -10268 -6806 -10190
rect 15334 -9737 15386 -9681
rect 15463 -9728 15515 -9672
rect 15585 -9725 15637 -9669
rect -4274 -10277 -4202 -10205
rect -4047 -10278 -3973 -10204
rect -3844 -10277 -3772 -10205
rect 6184 -10305 6312 -10177
rect 6474 -10305 6602 -10177
rect -53325 -10543 -53248 -10467
rect -53170 -10539 -53103 -10470
rect -33437 -10527 -33371 -10458
rect -33282 -10523 -33205 -10455
rect 26051 -9789 26111 -9726
rect 26183 -9786 26243 -9723
rect 26317 -9789 26377 -9726
rect -3402 -10662 -3304 -10577
rect -3179 -10646 -3081 -10561
rect -2936 -10646 -2838 -10561
rect -52653 -10936 -52576 -10860
rect -52498 -10932 -52431 -10863
rect -33063 -10970 -32952 -10859
rect -32797 -10968 -32688 -10859
rect -20018 -10982 -19863 -10827
rect -19686 -10982 -19533 -10829
rect 6474 -10992 6586 -10880
rect 6747 -10991 6857 -10881
rect 17294 -11004 17433 -10865
rect 17605 -11004 17742 -10867
rect 29254 -11230 29339 -11130
rect 16996 -11437 17131 -11301
rect 29243 -11406 29328 -11306
rect -20562 -11618 -20476 -11503
rect 16091 -11606 16172 -11530
rect -20565 -11819 -20479 -11704
rect 16087 -11814 16168 -11738
rect 16675 -11759 16810 -11623
rect 16996 -11770 17131 -11634
rect -18597 -12176 -18509 -12060
rect 6271 -12133 6370 -12060
rect 16675 -12113 16810 -11977
rect 28521 -12026 28576 -11974
rect 28512 -12161 28567 -12109
rect -64575 -12450 -64516 -12362
rect -18596 -12405 -18508 -12289
rect -64573 -12624 -64514 -12536
rect 6271 -12289 6370 -12216
rect -54294 -12674 -54231 -12584
rect -43772 -12607 -43666 -12447
rect 6266 -12445 6365 -12372
rect -54295 -12869 -54232 -12779
rect -43777 -12887 -43671 -12727
rect -34022 -12869 -33936 -12765
rect -34025 -13123 -33939 -13019
rect -32602 -12876 -32524 -12772
rect -5637 -12870 -5540 -12772
rect -32608 -13077 -32530 -12973
rect -5645 -13100 -5548 -13002
rect -53761 -13293 -53656 -13188
rect -53489 -13291 -53386 -13188
rect -65682 -13643 -65611 -13570
rect -65551 -13644 -65480 -13571
rect -65395 -13649 -65324 -13576
rect -55276 -13568 -55214 -13500
rect -55137 -13567 -55075 -13499
rect -55000 -13565 -54938 -13497
rect -44924 -13563 -44870 -13494
rect -44803 -13561 -44749 -13492
rect -44652 -13561 -44598 -13492
rect -65685 -13834 -65614 -13761
rect -65534 -13828 -65463 -13755
rect -65392 -13829 -65321 -13756
rect -53999 -13795 -53942 -13738
rect -23388 -13695 -23327 -13614
rect -23248 -13692 -23187 -13611
rect -23091 -13687 -23030 -13606
rect 4844 -13610 4907 -13536
rect 5001 -13613 5064 -13539
rect 5122 -13607 5185 -13533
rect -34681 -13820 -34623 -13755
rect -34539 -13814 -34481 -13749
rect -34394 -13822 -34336 -13757
rect -7132 -13752 -7080 -13688
rect -6994 -13756 -6942 -13692
rect -6827 -13752 -6775 -13688
rect 15328 -13727 15382 -13654
rect 15467 -13725 15521 -13652
rect 15611 -13727 15665 -13654
rect 26027 -13657 26088 -13579
rect 26180 -13649 26241 -13571
rect 26339 -13650 26400 -13572
rect -53999 -13915 -53944 -13860
rect -34693 -13992 -34635 -13927
rect -34547 -13989 -34489 -13924
rect -34387 -13981 -34329 -13916
rect -66349 -14584 -66289 -14521
rect -66217 -14581 -66157 -14518
rect -66083 -14584 -66023 -14521
rect -35385 -14627 -35314 -14547
rect -35245 -14624 -35174 -14544
rect -35093 -14623 -35022 -14543
rect -7903 -14546 -7831 -14459
rect -7762 -14546 -7690 -14459
rect -7624 -14547 -7552 -14460
rect 4077 -14531 4149 -14436
rect 4214 -14530 4286 -14435
rect 4359 -14530 4431 -14435
rect -45753 -14744 -45681 -14678
rect -45627 -14741 -45555 -14675
rect -45492 -14740 -45420 -14674
rect -24181 -14699 -24108 -14614
rect -24046 -14698 -23973 -14613
rect -23911 -14695 -23838 -14610
rect 14645 -14583 14697 -14527
rect 14761 -14583 14813 -14527
rect 14876 -14587 14928 -14531
rect 25360 -14556 25420 -14493
rect 25492 -14553 25552 -14490
rect 25626 -14556 25686 -14493
rect -63334 -14965 -63278 -14909
rect -5277 -14941 -5207 -14862
rect -63338 -15076 -63282 -15020
rect -31855 -15052 -31799 -14996
rect -3669 -14935 -3613 -14879
rect -42972 -15155 -42916 -15099
rect -31859 -15163 -31803 -15107
rect -17851 -15128 -17795 -15072
rect -42976 -15266 -42920 -15210
rect -5281 -15124 -5211 -15045
rect -3673 -15046 -3617 -14990
rect 7105 -14918 7161 -14862
rect 7101 -15029 7157 -14973
rect 17946 -14966 18002 -14910
rect 17942 -15077 17998 -15021
rect 28651 -14960 28707 -14904
rect 28647 -15071 28703 -15015
rect -17855 -15239 -17799 -15183
rect -32597 -15868 -32527 -15769
rect -64593 -15982 -64520 -15912
rect -55915 -15983 -55862 -15925
rect -55771 -15983 -55718 -15925
rect -55624 -15982 -55571 -15924
rect -64593 -16164 -64520 -16094
rect -43829 -16137 -43717 -16048
rect -32602 -16048 -32532 -15949
rect -18605 -15909 -18507 -15808
rect -18600 -16104 -18502 -16003
rect -5589 -15871 -5532 -15818
rect -5594 -15990 -5537 -15937
rect 6286 -15919 6347 -15840
rect -5592 -16103 -5535 -16050
rect 6285 -16102 6346 -16023
rect 16378 -16020 16441 -15950
rect 26041 -15963 26101 -15900
rect 26173 -15960 26233 -15897
rect 26307 -15963 26367 -15900
rect 16380 -16208 16443 -16138
rect -43832 -16367 -43720 -16278
rect -64337 -16838 -64259 -16760
rect -64336 -16984 -64260 -16908
rect -63656 -16935 -63600 -16879
rect -32183 -16887 -32114 -16809
rect -63660 -17046 -63604 -16990
rect -43324 -17028 -43268 -16972
rect -4920 -16859 -4856 -16795
rect -4002 -16819 -3932 -16754
rect -32183 -17069 -32114 -16991
rect -18441 -17051 -18359 -16969
rect -18276 -17051 -18194 -16969
rect -4923 -17007 -4859 -16943
rect -4008 -16978 -3938 -16913
rect 6667 -16836 6738 -16765
rect 6663 -17012 6734 -16941
rect 17448 -16891 17519 -16820
rect -43328 -17139 -43272 -17083
rect 17444 -17067 17515 -16996
rect 28339 -16832 28410 -16761
rect 28335 -17008 28406 -16937
rect -65672 -17331 -65612 -17268
rect -65540 -17328 -65480 -17265
rect -65406 -17331 -65346 -17268
rect -55285 -17266 -55233 -17198
rect -55152 -17266 -55100 -17198
rect -54986 -17264 -54934 -17196
rect -34694 -17378 -34636 -17311
rect -34572 -17376 -34514 -17309
rect -34438 -17374 -34380 -17307
rect -7135 -17295 -7080 -17230
rect -7005 -17294 -6950 -17229
rect -6871 -17291 -6816 -17226
rect 4843 -17269 4901 -17199
rect 4966 -17266 5024 -17196
rect 5105 -17267 5163 -17197
rect -44930 -17502 -44876 -17444
rect -44802 -17503 -44748 -17445
rect -44652 -17502 -44598 -17444
rect -23388 -17444 -23331 -17382
rect -23268 -17444 -23211 -17382
rect -23120 -17439 -23063 -17377
rect 15331 -17336 15383 -17280
rect 15472 -17329 15524 -17273
rect 15588 -17322 15640 -17266
rect 26041 -17312 26101 -17249
rect 26173 -17309 26233 -17246
rect 26307 -17312 26367 -17249
rect 17042 -17575 17108 -17509
rect -64123 -17747 -64070 -17685
rect 17042 -17764 17108 -17698
rect 27827 -17705 27893 -17639
rect -64123 -17884 -64070 -17822
rect 27826 -17872 27894 -17804
rect -53634 -18140 -53560 -18065
rect -53451 -18134 -53377 -18070
rect -63867 -18254 -63815 -18200
rect -32277 -18302 -32202 -18227
rect -4042 -18227 -3966 -18152
rect -63868 -18386 -63816 -18332
rect -44929 -18503 -44866 -18419
rect -44785 -18501 -44722 -18417
rect -44640 -18500 -44577 -18416
rect -55280 -18934 -55214 -18848
rect -55139 -18931 -55073 -18845
rect -54983 -18922 -54917 -18836
rect -53991 -18855 -53919 -18783
rect -63886 -19056 -63807 -18983
rect -53992 -19020 -53918 -18946
rect -63889 -19242 -63810 -19169
rect -53748 -19331 -53671 -19238
rect -64144 -19471 -64064 -19403
rect -53751 -19480 -53674 -19387
rect -64145 -19657 -64065 -19589
rect -18383 -18381 -18329 -18320
rect -18206 -18380 -18152 -18319
rect -32277 -18472 -32200 -18395
rect -4033 -18390 -3958 -18315
rect 6721 -18194 6780 -18133
rect 16702 -18099 16779 -18022
rect 6724 -18322 6783 -18261
rect 28123 -18094 28200 -18017
rect 16703 -18266 16778 -18191
rect 28124 -18241 28199 -18166
rect -34688 -19099 -34630 -19034
rect -34555 -19102 -34497 -19037
rect -34399 -19101 -34341 -19036
rect -23384 -19097 -23321 -19015
rect -23259 -19093 -23196 -19011
rect -23101 -19091 -23038 -19009
rect -7129 -19027 -7077 -18963
rect -6992 -19019 -6940 -18955
rect -6833 -19014 -6781 -18950
rect 4848 -19035 4911 -18961
rect 4986 -19035 5049 -18961
rect 5148 -19033 5211 -18959
rect 15336 -19047 15390 -18974
rect 15472 -19048 15526 -18975
rect 15628 -19046 15682 -18973
rect 26035 -19048 26096 -18970
rect 26187 -19039 26248 -18961
rect 26321 -19029 26382 -18951
rect -31960 -19393 -31904 -19337
rect -32280 -19589 -32218 -19528
rect -31954 -19515 -31898 -19459
rect -32282 -19717 -32220 -19656
rect -18343 -19727 -18238 -19622
rect -18124 -19727 -18017 -19620
rect -5590 -20172 -5533 -20120
rect -5593 -20308 -5536 -20256
rect 5842 -20282 5908 -20218
rect -3750 -20539 -3697 -20486
rect 5431 -20504 5486 -20448
rect 5842 -20438 5908 -20374
rect 6286 -20226 6343 -20166
rect 6284 -20372 6341 -20312
rect 17089 -20325 17158 -20217
rect 7005 -20505 7063 -20452
rect -18560 -20651 -18468 -20559
rect -18336 -20652 -18242 -20558
rect -3751 -20647 -3698 -20594
rect 5426 -20634 5481 -20578
rect 7004 -20628 7062 -20575
rect 17089 -20571 17158 -20463
rect -34026 -20965 -33939 -20871
rect -18864 -20932 -18772 -20840
rect 5597 -20851 5655 -20796
rect -4037 -20925 -3963 -20851
rect 6573 -20911 6637 -20855
rect 6714 -20918 6778 -20862
rect -34027 -21157 -33940 -21063
rect -19142 -21136 -19087 -21066
rect -18865 -21158 -18771 -21064
rect 5597 -20994 5655 -20939
rect -4037 -21145 -3963 -21071
rect -19140 -21299 -19085 -21229
rect -32282 -21380 -32210 -21308
rect -4036 -21335 -3964 -21263
rect -32283 -21568 -32209 -21494
rect -65679 -21752 -65617 -21655
rect -65545 -21745 -65483 -21648
rect -65410 -21754 -65348 -21657
rect -55288 -21749 -55226 -21677
rect -55155 -21749 -55093 -21677
rect -55004 -21745 -54942 -21673
rect -44932 -21688 -44878 -21621
rect -44775 -21689 -44721 -21622
rect -44610 -21686 -44556 -21619
rect -34695 -21721 -34637 -21652
rect -34539 -21718 -34481 -21649
rect -34377 -21713 -34319 -21644
rect -65683 -21945 -65621 -21848
rect -65535 -21945 -65473 -21848
rect -65388 -21948 -65326 -21851
rect -23388 -21766 -23320 -21674
rect -23233 -21771 -23165 -21679
rect -23086 -21772 -23018 -21680
rect -7139 -21759 -7079 -21679
rect -6975 -21757 -6915 -21677
rect -6828 -21750 -6768 -21670
rect 4842 -21726 4915 -21631
rect 4996 -21722 5069 -21627
rect 5143 -21724 5216 -21629
rect 15332 -21777 15388 -21705
rect 15472 -21780 15528 -21708
rect 15612 -21776 15668 -21704
rect 26028 -21708 26084 -21627
rect 26172 -21708 26228 -21627
rect 26307 -21705 26363 -21624
rect -31954 -21922 -31889 -21859
rect -3754 -21940 -3696 -21882
rect -31959 -22094 -31894 -22031
rect -3756 -22054 -3698 -21996
rect -66363 -22677 -66303 -22614
rect -66231 -22674 -66171 -22611
rect -66097 -22677 -66037 -22614
rect -55917 -22631 -55837 -22528
rect -55769 -22632 -55689 -22529
rect -55630 -22630 -55550 -22527
rect -45752 -22671 -45700 -22615
rect -45624 -22664 -45572 -22608
rect -45464 -22661 -45412 -22605
rect -24172 -22690 -24112 -22603
rect -24039 -22687 -23979 -22600
rect -23895 -22680 -23835 -22593
rect 4094 -22718 4146 -22662
rect 4232 -22715 4284 -22659
rect 4361 -22713 4413 -22657
rect 14652 -22634 14704 -22578
rect 14765 -22627 14817 -22571
rect 14888 -22627 14940 -22571
rect 25353 -22682 25413 -22619
rect 25485 -22679 25545 -22616
rect 25619 -22682 25679 -22619
rect -63383 -23068 -63327 -23012
rect -63387 -23179 -63331 -23123
rect -53191 -23036 -53135 -22980
rect -53195 -23147 -53139 -23091
rect -42800 -23045 -42744 -22989
rect -42804 -23156 -42748 -23100
rect -17892 -23057 -17836 -23001
rect 14658 -23069 14710 -23013
rect 14771 -23062 14823 -23006
rect 14894 -23062 14946 -23006
rect -17896 -23168 -17840 -23112
rect 4093 -23155 4145 -23099
rect 4231 -23152 4283 -23096
rect 4360 -23150 4412 -23094
rect 25354 -23108 25414 -23045
rect 25486 -23105 25546 -23042
rect 25620 -23108 25680 -23045
rect -68519 -23497 -68436 -23421
rect -66855 -23497 -66759 -23417
rect -64355 -24084 -64297 -24026
rect -54223 -24059 -54171 -24001
rect -64361 -24265 -64303 -24207
rect -54228 -24229 -54176 -24171
rect -43793 -24082 -43740 -24018
rect -19149 -24048 -19082 -23981
rect 5833 -24003 5909 -23940
rect 17087 -23870 17153 -23782
rect 17086 -24045 17152 -23957
rect 26043 -24073 26103 -24010
rect 26175 -24070 26235 -24007
rect 26309 -24073 26369 -24010
rect -43796 -24264 -43743 -24200
rect -35377 -24235 -35325 -24179
rect -35251 -24237 -35199 -24181
rect -35104 -24236 -35052 -24180
rect -19154 -24238 -19087 -24171
rect -7900 -24190 -7848 -24134
rect -7785 -24191 -7733 -24135
rect -7663 -24190 -7611 -24134
rect 5834 -24160 5910 -24097
rect -63726 -25008 -63670 -24952
rect -63730 -25119 -63674 -25063
rect -53526 -24971 -53467 -24909
rect -18255 -24936 -18173 -24854
rect -53543 -25109 -53484 -25047
rect -43341 -25117 -43267 -25050
rect -43186 -25104 -43112 -25037
rect -18255 -25101 -18173 -25019
rect 6666 -25067 6734 -24990
rect 6880 -25051 6948 -24974
rect -65672 -25434 -65612 -25371
rect -65540 -25431 -65480 -25368
rect -65406 -25434 -65346 -25371
rect -55272 -25383 -55192 -25280
rect -55120 -25384 -55040 -25281
rect -54983 -25383 -54903 -25280
rect 17338 -25055 17421 -24962
rect 17593 -25045 17676 -24952
rect 28407 -24969 28463 -24912
rect 28314 -25072 28370 -25015
rect -44926 -25416 -44874 -25360
rect -44810 -25410 -44758 -25354
rect -44693 -25408 -44641 -25352
rect -34692 -25343 -34634 -25274
rect -34558 -25342 -34500 -25273
rect -34430 -25340 -34372 -25271
rect -23383 -25448 -23323 -25361
rect -23250 -25445 -23190 -25358
rect -23106 -25438 -23046 -25351
rect -7135 -25370 -7078 -25308
rect -6999 -25372 -6942 -25310
rect -6840 -25367 -6783 -25305
rect 4859 -25462 4911 -25406
rect 5002 -25463 5054 -25407
rect 5117 -25458 5169 -25402
rect 15341 -25392 15393 -25336
rect 15457 -25381 15509 -25325
rect 15582 -25386 15634 -25330
rect 26045 -25418 26105 -25355
rect 26177 -25415 26237 -25352
rect 26311 -25418 26371 -25355
rect -66369 -25702 -66299 -25618
rect -66204 -25699 -66134 -25615
rect -66063 -25699 -65993 -25615
rect -64119 -25758 -64066 -25692
rect -64127 -25884 -64074 -25818
rect 6419 -25848 6495 -25772
rect 27825 -25770 27893 -25702
rect 6424 -25854 6490 -25848
rect 27826 -25943 27892 -25877
rect 6423 -26030 6491 -25962
rect -53999 -26118 -53922 -26041
rect -63865 -26238 -63812 -26184
rect -33372 -26172 -33315 -26115
rect -63860 -26347 -63807 -26292
rect -53999 -26302 -53924 -26227
rect -43616 -26338 -43555 -26282
rect -18858 -26192 -18781 -26115
rect -33366 -26303 -33311 -26248
rect -4581 -26121 -4524 -26064
rect 28123 -26197 28198 -26122
rect -18858 -26365 -18783 -26290
rect -4581 -26258 -4526 -26203
rect 6710 -26390 6785 -26315
rect -68598 -26561 -68504 -26477
rect -66935 -26559 -66854 -26469
rect -43618 -26462 -43557 -26406
rect -34684 -26683 -34632 -26627
rect -34552 -26675 -34500 -26619
rect -34407 -26670 -34355 -26614
rect -23390 -26698 -23322 -26606
rect -23225 -26705 -23157 -26613
rect -23080 -26705 -23012 -26613
rect -7135 -26637 -7083 -26581
rect -6996 -26628 -6944 -26572
rect -6866 -26623 -6814 -26567
rect -34568 -26826 -34510 -26757
rect -65682 -27209 -65616 -27118
rect -65522 -27207 -65456 -27116
rect -65380 -27209 -65314 -27118
rect -55286 -27130 -55224 -27058
rect -55145 -27130 -55083 -27058
rect -54971 -27118 -54909 -27046
rect -44934 -27047 -44876 -26969
rect -44792 -27046 -44734 -26968
rect -44625 -27049 -44567 -26971
rect -34568 -27018 -34510 -26949
rect -33031 -26919 -32973 -26862
rect -33034 -27041 -32976 -26984
rect 4840 -26658 4913 -26565
rect 4985 -26657 5058 -26564
rect 5131 -26660 5204 -26567
rect 6709 -26558 6786 -26481
rect -4282 -26915 -4227 -26860
rect -4151 -26912 -4096 -26857
rect 15336 -27044 15401 -26951
rect 15480 -27042 15545 -26949
rect 15622 -27044 15687 -26951
rect 6707 -27221 6785 -27136
rect 28119 -26352 28195 -26277
rect 6709 -27381 6787 -27296
rect 6418 -27601 6498 -27521
rect 26027 -26979 26103 -26878
rect 26184 -26983 26260 -26882
rect 26333 -26981 26409 -26880
rect 6415 -27758 6495 -27678
rect -43801 -27856 -43741 -27798
rect -43803 -27994 -43743 -27936
rect -54225 -28121 -54170 -28060
rect -54229 -28285 -54174 -28224
rect -43887 -28233 -43827 -28172
rect -43891 -28398 -43831 -28337
rect -19151 -27939 -19083 -27877
rect -19151 -28105 -19083 -28043
rect -4570 -28106 -4499 -28030
rect -19388 -28274 -19326 -28215
rect -4569 -28331 -4498 -28255
rect -64357 -28505 -64291 -28449
rect -19391 -28439 -19329 -28380
rect -43607 -28564 -43551 -28498
rect -18955 -28580 -18890 -28505
rect -64364 -28664 -64298 -28608
rect -54400 -28676 -54342 -28621
rect -54406 -28839 -54348 -28784
rect -54099 -28654 -54037 -28596
rect -43616 -28717 -43560 -28651
rect -32650 -28652 -32581 -28586
rect -54098 -28809 -54036 -28751
rect -32652 -28772 -32583 -28706
rect -18961 -28774 -18896 -28699
rect -56389 -29119 -56253 -29010
rect -53823 -28941 -53745 -28852
rect -32932 -28909 -32873 -28848
rect -53819 -29146 -53741 -29057
rect -43332 -29004 -43262 -28920
rect -32939 -29025 -32880 -28964
rect -43340 -29160 -43270 -29076
rect -18667 -29054 -18602 -28987
rect -56397 -29368 -56261 -29259
rect -18681 -29242 -18616 -29175
rect -32649 -29506 -32575 -29432
rect -32648 -29678 -32576 -29606
rect -55284 -29823 -55223 -29745
rect -55142 -29817 -55081 -29739
rect -54974 -29820 -54913 -29742
rect -44931 -29827 -44876 -29756
rect -44788 -29828 -44733 -29757
rect -44626 -29823 -44571 -29752
rect -34684 -29818 -34627 -29738
rect -34562 -29814 -34505 -29734
rect -34424 -29813 -34367 -29733
rect -7135 -29783 -7069 -29686
rect -7009 -29782 -6943 -29685
rect -6879 -29781 -6813 -29684
rect 6708 -29667 6764 -29611
rect 4844 -29869 4918 -29793
rect 4991 -29866 5065 -29790
rect 5139 -29867 5213 -29791
rect 6708 -29780 6764 -29724
rect 26023 -29845 26089 -29775
rect 26175 -29846 26241 -29776
rect 26318 -29842 26384 -29772
rect -66366 -30126 -66289 -30044
rect -66217 -30119 -66140 -30037
rect -66067 -30120 -65990 -30038
rect -23386 -30075 -23320 -29990
rect -23232 -30069 -23166 -29984
rect -23092 -30067 -23026 -29982
rect -32935 -30207 -32865 -30135
rect 15334 -30191 15405 -30101
rect 15479 -30188 15550 -30098
rect 15636 -30184 15707 -30094
rect -32943 -30361 -32873 -30289
rect -56668 -30592 -56587 -30528
rect 6412 -30527 6492 -30446
rect -56677 -30743 -56596 -30679
rect -55913 -30767 -55853 -30704
rect -55781 -30764 -55721 -30701
rect -55647 -30767 -55587 -30704
rect -45735 -30771 -45675 -30708
rect -45603 -30768 -45543 -30705
rect -45469 -30771 -45409 -30708
rect -24156 -30705 -24096 -30642
rect -24024 -30702 -23964 -30639
rect -23890 -30705 -23830 -30642
rect 6415 -30668 6495 -30587
rect -7897 -30805 -7837 -30742
rect -7765 -30802 -7705 -30739
rect -7631 -30805 -7571 -30742
rect 14660 -30785 14720 -30722
rect 14792 -30782 14852 -30719
rect 14926 -30785 14986 -30722
rect -66369 -31079 -66310 -31018
rect -66256 -31076 -66197 -31015
rect -66108 -31074 -66049 -31013
rect -55913 -31203 -55853 -31140
rect -55781 -31200 -55721 -31137
rect -55647 -31203 -55587 -31140
rect -45729 -31181 -45669 -31118
rect -45597 -31178 -45537 -31115
rect -45463 -31181 -45403 -31118
rect -24156 -31140 -24096 -31077
rect -24024 -31137 -23964 -31074
rect -23890 -31140 -23830 -31077
rect -57009 -31300 -56906 -31228
rect -7897 -31241 -7837 -31178
rect -7765 -31238 -7705 -31175
rect -7631 -31241 -7571 -31178
rect 14660 -31216 14720 -31153
rect 14792 -31213 14852 -31150
rect 14926 -31216 14986 -31153
rect -57019 -31480 -56916 -31408
rect -57382 -31663 -57283 -31584
rect -65665 -31778 -65606 -31717
rect -65522 -31775 -65463 -31714
rect -65397 -31780 -65338 -31719
rect -57379 -31830 -57280 -31751
rect -54411 -32019 -54345 -31953
rect -43893 -32051 -43827 -31995
rect -19382 -32014 -19329 -31953
rect -54410 -32204 -54344 -32138
rect -43895 -32210 -43829 -32154
rect -19384 -32173 -19331 -32112
rect -4562 -32060 -4493 -31993
rect 16383 -31985 16454 -31906
rect -4568 -32237 -4499 -32170
rect 16384 -32191 16455 -32112
rect -66371 -32570 -66312 -32509
rect -66231 -32568 -66172 -32507
rect -66098 -32555 -66039 -32494
rect -57715 -32502 -57596 -32415
rect -35375 -32533 -35315 -32470
rect -35243 -32530 -35183 -32467
rect -35109 -32533 -35049 -32470
rect -57733 -32724 -57614 -32637
rect 4088 -32657 4148 -32594
rect 4220 -32654 4280 -32591
rect 4354 -32657 4414 -32594
rect -53632 -33162 -53556 -33086
rect -53468 -33163 -53390 -33085
rect -65676 -33271 -65617 -33210
rect -65532 -33269 -65473 -33208
rect -65384 -33266 -65325 -33205
rect -43133 -33147 -43077 -33088
rect -43020 -33144 -42964 -33085
rect -18438 -33149 -18377 -33081
rect -18259 -33147 -18198 -33079
rect -4122 -33175 -4054 -33114
rect -3968 -33153 -3900 -33092
rect 17525 -33157 17583 -33093
rect 17683 -33155 17741 -33091
rect -66369 -33744 -66310 -33683
rect -66216 -33744 -66157 -33683
rect -66078 -33742 -66019 -33681
rect -58055 -33473 -57975 -33392
rect -55258 -33509 -55198 -33446
rect -55126 -33506 -55066 -33443
rect -54992 -33509 -54932 -33446
rect -44921 -33513 -44861 -33450
rect -44789 -33510 -44729 -33447
rect -44655 -33513 -44595 -33450
rect -34697 -33450 -34640 -33382
rect -34562 -33450 -34505 -33382
rect -34393 -33447 -34336 -33379
rect -23380 -33447 -23320 -33384
rect -23248 -33444 -23188 -33381
rect -23114 -33447 -23054 -33384
rect -7128 -33551 -7068 -33488
rect -6996 -33548 -6936 -33485
rect -6862 -33551 -6802 -33488
rect 4841 -33486 4907 -33419
rect 4998 -33484 5064 -33417
rect 5135 -33485 5201 -33418
rect 15348 -33528 15408 -33465
rect 15480 -33525 15540 -33462
rect 15614 -33528 15674 -33465
rect 26028 -33469 26094 -33399
rect 26162 -33469 26228 -33399
rect 26311 -33465 26377 -33395
rect -58069 -33673 -57989 -33592
rect -65683 -34443 -65624 -34382
rect -65545 -34440 -65486 -34379
rect -65399 -34440 -65340 -34379
rect -58410 -34481 -58313 -34399
rect -54103 -34289 -54050 -34227
rect -43609 -34308 -43554 -34255
rect -54109 -34417 -54056 -34355
rect -18964 -34257 -18901 -34196
rect -43614 -34434 -43559 -34381
rect -18963 -34377 -18900 -34316
rect -58415 -34661 -58318 -34579
rect -32275 -34461 -32218 -34404
rect -4166 -34513 -4075 -34415
rect -4001 -34502 -3910 -34404
rect 17381 -34469 17446 -34405
rect 17499 -34469 17564 -34405
rect -32275 -34601 -32220 -34546
rect 5606 -34579 5663 -34522
rect -55924 -34727 -55864 -34645
rect -55798 -34731 -55738 -34649
rect -55659 -34724 -55599 -34642
rect 5607 -34723 5662 -34668
rect -65687 -35679 -65624 -35613
rect -65544 -35676 -65481 -35610
rect -65411 -35671 -65348 -35605
rect -54413 -35604 -54350 -35544
rect -44922 -35077 -44867 -35006
rect -44782 -35081 -44727 -35010
rect -44632 -35092 -44577 -35021
rect -34685 -34975 -34625 -34912
rect -34553 -34972 -34493 -34909
rect -34419 -34975 -34359 -34912
rect -23389 -34995 -23317 -34911
rect -23236 -34993 -23164 -34909
rect -23087 -34990 -23015 -34906
rect -7137 -35114 -7071 -35025
rect -6984 -35110 -6918 -35021
rect -6842 -35106 -6776 -35017
rect 4853 -35093 4913 -35030
rect 4985 -35090 5045 -35027
rect 5119 -35093 5179 -35030
rect 15333 -35111 15404 -35021
rect 15470 -35111 15541 -35021
rect 15601 -35107 15672 -35017
rect -32072 -35260 -32010 -35207
rect 26033 -35155 26099 -35085
rect 26175 -35153 26241 -35083
rect 26315 -35158 26381 -35088
rect -32075 -35408 -32013 -35355
rect 5426 -35299 5486 -35236
rect 5426 -35432 5486 -35369
rect 17882 -35499 17963 -35419
rect -55277 -36228 -55219 -36150
rect -55148 -36228 -55090 -36150
rect -55002 -36234 -54944 -36156
rect -57382 -36552 -57288 -36485
rect -57382 -36690 -57288 -36623
rect -58065 -36963 -57992 -36892
rect -45753 -36524 -45695 -36426
rect -45595 -36524 -45537 -36426
rect -45463 -36516 -45405 -36418
rect -58062 -37120 -57989 -37049
rect -24177 -36120 -24120 -36035
rect -24036 -36119 -23979 -36034
rect -23891 -36120 -23834 -36035
rect -19550 -36980 -19493 -36895
rect -19388 -36969 -19331 -36884
rect -3675 -35637 -3605 -35569
rect -3515 -35635 -3445 -35567
rect 6128 -35648 6218 -35558
rect 6399 -35661 6495 -35545
rect 17881 -35639 17962 -35559
rect -3975 -35770 -3883 -35693
rect -3985 -35935 -3866 -35838
rect 6418 -35931 6526 -35844
rect 6687 -35936 6811 -35839
rect 17255 -35938 17337 -35861
rect 17403 -35939 17485 -35862
rect 17557 -35934 17639 -35857
rect -7898 -36231 -7842 -36150
rect -7758 -36227 -7702 -36146
rect -7611 -36221 -7555 -36140
rect 4082 -36297 4138 -36216
rect 4243 -36297 4299 -36216
rect 4400 -36299 4456 -36218
rect 14656 -36414 14723 -36332
rect 14793 -36410 14860 -36328
rect 14935 -36414 15002 -36332
rect -4705 -37121 -4648 -37038
rect -4584 -37114 -4527 -37031
rect 5792 -37158 5848 -37076
rect 5919 -37153 5975 -37071
rect -58410 -37459 -58341 -37406
rect -43923 -37411 -43865 -37313
rect -43808 -37410 -43750 -37312
rect -23380 -37633 -23323 -37548
rect -23229 -37623 -23172 -37538
rect -23089 -37621 -23032 -37536
rect -7132 -37744 -7076 -37663
rect -6982 -37739 -6926 -37658
rect -6858 -37730 -6802 -37649
rect -57731 -38116 -57631 -38058
rect -44929 -38051 -44871 -37953
rect -44782 -38051 -44724 -37953
rect -44623 -38046 -44565 -37948
rect -57732 -38244 -57632 -38186
rect 16226 -37266 16291 -37205
rect 16357 -37260 16422 -37199
rect 16823 -37283 16883 -37209
rect 16950 -37276 17010 -37202
rect 17067 -37274 17127 -37200
rect 4856 -37804 4919 -37716
rect 4998 -37804 5061 -37716
rect 5125 -37802 5188 -37714
rect -57731 -38354 -57631 -38296
rect -56683 -38745 -56580 -38680
rect 15331 -37923 15398 -37841
rect 15466 -37923 15533 -37841
rect 15617 -37922 15684 -37840
rect -56690 -38881 -56587 -38816
rect -57012 -39128 -56931 -39064
rect -57008 -39254 -56927 -39190
rect -57010 -39379 -56929 -39315
<< metal2 >>
rect -66381 60800 -65982 60875
rect -66381 60795 -66142 60800
rect -66381 60691 -66351 60795
rect -66237 60696 -66142 60795
rect -66028 60696 -65982 60800
rect -66237 60691 -65982 60696
rect -66381 60630 -65982 60691
rect -66381 60526 -66354 60630
rect -66240 60629 -65982 60630
rect -66240 60526 -66141 60629
rect -66381 60525 -66141 60526
rect -66027 60525 -65982 60629
rect -66381 60104 -65982 60525
rect -66381 60000 -66351 60104
rect -66237 60000 -66128 60104
rect -66014 60000 -65982 60104
rect -66381 59948 -65982 60000
rect -66381 59947 -66128 59948
rect -66381 59843 -66350 59947
rect -66236 59844 -66128 59947
rect -66014 59844 -65982 59948
rect -66236 59843 -65982 59844
rect -66381 57176 -65982 59843
rect -66381 57175 -66214 57176
rect -70909 57141 -70510 57148
rect -70909 57140 -70742 57141
rect -70909 57087 -70897 57140
rect -70844 57088 -70742 57140
rect -70689 57088 -70584 57141
rect -70531 57088 -70510 57141
rect -70844 57087 -70510 57088
rect -70909 57034 -70510 57087
rect -70909 56981 -70895 57034
rect -70842 57031 -70510 57034
rect -70842 56981 -70738 57031
rect -70909 56978 -70738 56981
rect -70685 56978 -70585 57031
rect -70532 56978 -70510 57031
rect -70909 56926 -70510 56978
rect -70909 56925 -70738 56926
rect -70909 56872 -70896 56925
rect -70843 56873 -70738 56925
rect -70685 56924 -70510 56926
rect -70685 56873 -70586 56924
rect -70843 56872 -70586 56873
rect -70909 56871 -70586 56872
rect -70533 56871 -70510 56924
rect -70909 56816 -70510 56871
rect -70909 56763 -70893 56816
rect -70840 56815 -70510 56816
rect -70840 56763 -70737 56815
rect -70909 56762 -70737 56763
rect -70684 56762 -70584 56815
rect -70531 56762 -70510 56815
rect -70909 52578 -70510 56762
rect -70915 52576 -70510 52578
rect -70223 57140 -69824 57148
rect -70223 57139 -70055 57140
rect -70223 57086 -70210 57139
rect -70157 57087 -70055 57139
rect -70002 57087 -69897 57140
rect -69844 57087 -69824 57140
rect -70157 57086 -69824 57087
rect -70223 57033 -69824 57086
rect -70223 56980 -70208 57033
rect -70155 57030 -69824 57033
rect -70155 56980 -70051 57030
rect -70223 56977 -70051 56980
rect -69998 56977 -69898 57030
rect -69845 56977 -69824 57030
rect -70223 56925 -69824 56977
rect -70223 56924 -70051 56925
rect -70223 56871 -70209 56924
rect -70156 56872 -70051 56924
rect -69998 56923 -69824 56925
rect -69998 56872 -69899 56923
rect -70156 56871 -69899 56872
rect -70223 56870 -69899 56871
rect -69846 56870 -69824 56923
rect -70223 56815 -69824 56870
rect -70223 56762 -70206 56815
rect -70153 56814 -69824 56815
rect -70153 56762 -70050 56814
rect -70223 56761 -70050 56762
rect -69997 56761 -69897 56814
rect -69844 56761 -69824 56814
rect -70223 53624 -69824 56761
rect -66381 57122 -66369 57175
rect -66316 57123 -66214 57175
rect -66161 57123 -66056 57176
rect -66003 57123 -65982 57176
rect -66316 57122 -65982 57123
rect -66381 57069 -65982 57122
rect -66381 57016 -66367 57069
rect -66314 57066 -65982 57069
rect -66314 57016 -66210 57066
rect -66381 57013 -66210 57016
rect -66157 57013 -66057 57066
rect -66004 57013 -65982 57066
rect -66381 56961 -65982 57013
rect -66381 56960 -66210 56961
rect -66381 56907 -66368 56960
rect -66315 56908 -66210 56960
rect -66157 56959 -65982 56961
rect -66157 56908 -66058 56959
rect -66315 56907 -66058 56908
rect -66381 56906 -66058 56907
rect -66005 56906 -65982 56959
rect -66381 56851 -65982 56906
rect -66381 56798 -66365 56851
rect -66312 56850 -65982 56851
rect -66312 56798 -66209 56850
rect -66381 56797 -66209 56798
rect -66156 56797 -66056 56850
rect -66003 56797 -65982 56850
rect -66381 54811 -65982 56797
rect -65695 57172 -65296 57182
rect -65695 57171 -65528 57172
rect -65695 57118 -65683 57171
rect -65630 57119 -65528 57171
rect -65475 57119 -65370 57172
rect -65317 57119 -65296 57172
rect -65630 57118 -65296 57119
rect -65695 57065 -65296 57118
rect -65695 57012 -65681 57065
rect -65628 57062 -65296 57065
rect -65628 57012 -65524 57062
rect -65695 57009 -65524 57012
rect -65471 57009 -65371 57062
rect -65318 57009 -65296 57062
rect -65695 56957 -65296 57009
rect -65695 56956 -65524 56957
rect -65695 56903 -65682 56956
rect -65629 56904 -65524 56956
rect -65471 56955 -65296 56957
rect -65471 56904 -65372 56955
rect -65629 56903 -65372 56904
rect -65695 56902 -65372 56903
rect -65319 56902 -65296 56955
rect -65695 56847 -65296 56902
rect -65695 56794 -65679 56847
rect -65626 56846 -65296 56847
rect -65626 56794 -65523 56846
rect -65695 56793 -65523 56794
rect -65470 56793 -65370 56846
rect -65317 56793 -65296 56846
rect -65695 55849 -65296 56793
rect -8574 56766 -8343 56775
rect -8574 56713 -8560 56766
rect -8508 56765 -8343 56766
rect -8508 56713 -8423 56765
rect -8574 56712 -8423 56713
rect -8371 56712 -8343 56765
rect -8574 56620 -8343 56712
rect -8574 56567 -8555 56620
rect -8503 56567 -8409 56620
rect -8357 56567 -8343 56620
rect -65695 55832 -65284 55849
rect -65695 55829 -65367 55832
rect -65695 55824 -65516 55829
rect -65695 55729 -65675 55824
rect -65598 55734 -65516 55824
rect -65439 55737 -65367 55829
rect -65290 55737 -65284 55832
rect -65439 55734 -65284 55737
rect -65598 55729 -65284 55734
rect -65695 55656 -65284 55729
rect -65695 55653 -65370 55656
rect -65695 55648 -65519 55653
rect -65695 55553 -65678 55648
rect -65601 55558 -65519 55648
rect -65442 55561 -65370 55653
rect -65293 55561 -65284 55656
rect -65442 55558 -65284 55561
rect -65601 55553 -65284 55558
rect -65695 55497 -65284 55553
rect -65695 55494 -65368 55497
rect -65695 55489 -65517 55494
rect -65695 55394 -65676 55489
rect -65599 55399 -65517 55489
rect -65440 55402 -65368 55494
rect -65291 55402 -65284 55497
rect -65440 55399 -65284 55402
rect -65599 55394 -65284 55399
rect -65695 55339 -65284 55394
rect -65695 55336 -65369 55339
rect -65695 55331 -65518 55336
rect -65695 55236 -65677 55331
rect -65600 55241 -65518 55331
rect -65441 55244 -65369 55336
rect -65292 55244 -65284 55339
rect -65441 55241 -65284 55244
rect -65600 55236 -65284 55241
rect -65695 55224 -65284 55236
rect -66381 54794 -65971 54811
rect -66381 54791 -66054 54794
rect -66381 54786 -66203 54791
rect -66381 54691 -66362 54786
rect -66285 54696 -66203 54786
rect -66126 54699 -66054 54791
rect -65977 54699 -65971 54794
rect -66126 54696 -65971 54699
rect -66285 54691 -65971 54696
rect -66381 54618 -65971 54691
rect -66381 54615 -66057 54618
rect -66381 54610 -66206 54615
rect -66381 54515 -66365 54610
rect -66288 54520 -66206 54610
rect -66129 54523 -66057 54615
rect -65980 54523 -65971 54618
rect -66129 54520 -65971 54523
rect -66288 54515 -65971 54520
rect -66381 54459 -65971 54515
rect -66381 54456 -66055 54459
rect -66381 54451 -66204 54456
rect -66381 54356 -66363 54451
rect -66286 54361 -66204 54451
rect -66127 54364 -66055 54456
rect -65978 54364 -65971 54459
rect -66127 54361 -65971 54364
rect -66286 54356 -65971 54361
rect -66381 54301 -65971 54356
rect -66381 54298 -66056 54301
rect -66381 54293 -66205 54298
rect -66381 54198 -66364 54293
rect -66287 54203 -66205 54293
rect -66128 54206 -66056 54298
rect -65979 54206 -65971 54301
rect -66128 54203 -65971 54206
rect -66287 54198 -65971 54203
rect -66381 54186 -65971 54198
rect -70223 53607 -69812 53624
rect -70223 53604 -69895 53607
rect -70223 53599 -70044 53604
rect -70223 53504 -70203 53599
rect -70126 53509 -70044 53599
rect -69967 53512 -69895 53604
rect -69818 53512 -69812 53607
rect -69967 53509 -69812 53512
rect -70126 53504 -69812 53509
rect -70223 53431 -69812 53504
rect -70223 53428 -69898 53431
rect -70223 53423 -70047 53428
rect -70223 53328 -70206 53423
rect -70129 53333 -70047 53423
rect -69970 53336 -69898 53428
rect -69821 53336 -69812 53431
rect -69970 53333 -69812 53336
rect -70129 53328 -69812 53333
rect -70223 53272 -69812 53328
rect -70223 53269 -69896 53272
rect -70223 53264 -70045 53269
rect -70223 53169 -70204 53264
rect -70127 53174 -70045 53264
rect -69968 53177 -69896 53269
rect -69819 53177 -69812 53272
rect -69968 53174 -69812 53177
rect -70127 53169 -69812 53174
rect -70223 53114 -69812 53169
rect -70223 53111 -69897 53114
rect -70223 53106 -70046 53111
rect -70223 53011 -70205 53106
rect -70128 53016 -70046 53106
rect -69969 53019 -69897 53111
rect -69820 53019 -69812 53114
rect -69969 53016 -69812 53019
rect -70128 53011 -69812 53016
rect -70223 52999 -69812 53011
rect -70915 52559 -70508 52576
rect -70915 52556 -70591 52559
rect -70915 52551 -70740 52556
rect -70915 52456 -70899 52551
rect -70822 52461 -70740 52551
rect -70663 52464 -70591 52556
rect -70514 52464 -70508 52559
rect -70663 52461 -70508 52464
rect -70822 52456 -70508 52461
rect -70915 52383 -70508 52456
rect -70915 52380 -70594 52383
rect -70915 52375 -70743 52380
rect -70915 52280 -70902 52375
rect -70825 52285 -70743 52375
rect -70666 52288 -70594 52380
rect -70517 52288 -70508 52383
rect -70666 52285 -70508 52288
rect -70825 52280 -70508 52285
rect -70915 52224 -70508 52280
rect -70915 52221 -70592 52224
rect -70915 52216 -70741 52221
rect -70915 52121 -70900 52216
rect -70823 52126 -70741 52216
rect -70664 52129 -70592 52221
rect -70515 52129 -70508 52224
rect -70664 52126 -70508 52129
rect -70823 52121 -70508 52126
rect -70915 52066 -70508 52121
rect -70915 52063 -70593 52066
rect -70915 52058 -70742 52063
rect -70915 51963 -70901 52058
rect -70824 51968 -70742 52058
rect -70665 51971 -70593 52063
rect -70516 51971 -70508 52066
rect -70665 51968 -70508 51971
rect -70824 51963 -70508 51968
rect -70915 51951 -70508 51963
rect -70915 51950 -70510 51951
rect -70909 44208 -70510 51950
rect -70911 44206 -70510 44208
rect -70223 45249 -69824 52999
rect -66381 49606 -65982 54186
rect -66381 49599 -66090 49606
rect -66381 49597 -66220 49599
rect -66381 49539 -66361 49597
rect -66296 49541 -66220 49597
rect -66155 49548 -66090 49599
rect -66025 49548 -65982 49606
rect -66155 49541 -65982 49548
rect -66296 49539 -65982 49541
rect -66381 48120 -65982 49539
rect -66381 48062 -66365 48120
rect -66300 48119 -65982 48120
rect -66300 48062 -66223 48119
rect -66381 48061 -66223 48062
rect -66158 48061 -66078 48119
rect -66013 48061 -65982 48119
rect -66381 46683 -65982 48061
rect -66381 46663 -66086 46683
rect -66381 46654 -66232 46663
rect -66381 46596 -66365 46654
rect -66300 46605 -66232 46654
rect -66167 46625 -66086 46663
rect -66021 46625 -65982 46683
rect -66167 46605 -65982 46625
rect -66300 46596 -65982 46605
rect -70223 45232 -69812 45249
rect -70223 45229 -69895 45232
rect -70223 45224 -70044 45229
rect -70223 45129 -70203 45224
rect -70126 45134 -70044 45224
rect -69967 45137 -69895 45229
rect -69818 45137 -69812 45232
rect -69967 45134 -69812 45137
rect -70126 45129 -69812 45134
rect -70223 45056 -69812 45129
rect -70223 45053 -69898 45056
rect -70223 45048 -70047 45053
rect -70223 44953 -70206 45048
rect -70129 44958 -70047 45048
rect -69970 44961 -69898 45053
rect -69821 44961 -69812 45056
rect -69970 44958 -69812 44961
rect -70129 44953 -69812 44958
rect -70223 44897 -69812 44953
rect -70223 44894 -69896 44897
rect -70223 44889 -70045 44894
rect -70223 44794 -70204 44889
rect -70127 44799 -70045 44889
rect -69968 44802 -69896 44894
rect -69819 44802 -69812 44897
rect -69968 44799 -69812 44802
rect -70127 44794 -69812 44799
rect -70223 44739 -69812 44794
rect -70223 44736 -69897 44739
rect -70223 44731 -70046 44736
rect -70223 44636 -70205 44731
rect -70128 44641 -70046 44731
rect -69969 44644 -69897 44736
rect -69820 44644 -69812 44739
rect -69969 44641 -69812 44644
rect -70128 44636 -69812 44641
rect -70223 44624 -69812 44636
rect -70911 44189 -70504 44206
rect -70911 44186 -70587 44189
rect -70911 44181 -70736 44186
rect -70911 44086 -70895 44181
rect -70818 44091 -70736 44181
rect -70659 44094 -70587 44186
rect -70510 44094 -70504 44189
rect -70659 44091 -70504 44094
rect -70818 44086 -70504 44091
rect -70911 44013 -70504 44086
rect -70911 44010 -70590 44013
rect -70911 44005 -70739 44010
rect -70911 43910 -70898 44005
rect -70821 43915 -70739 44005
rect -70662 43918 -70590 44010
rect -70513 43918 -70504 44013
rect -70662 43915 -70504 43918
rect -70821 43910 -70504 43915
rect -70911 43854 -70504 43910
rect -70911 43851 -70588 43854
rect -70911 43846 -70737 43851
rect -70911 43751 -70896 43846
rect -70819 43756 -70737 43846
rect -70660 43759 -70588 43851
rect -70511 43759 -70504 43854
rect -70660 43756 -70504 43759
rect -70819 43751 -70504 43756
rect -70911 43696 -70504 43751
rect -70911 43693 -70589 43696
rect -70911 43688 -70738 43693
rect -70911 43593 -70897 43688
rect -70820 43598 -70738 43688
rect -70661 43601 -70589 43693
rect -70512 43601 -70504 43696
rect -70661 43598 -70504 43601
rect -70820 43593 -70504 43598
rect -70911 43581 -70504 43593
rect -70911 43580 -70510 43581
rect -70909 35781 -70510 43580
rect -70223 37032 -69824 44624
rect -66381 43235 -65982 46596
rect -66381 43230 -66069 43235
rect -66381 43148 -66357 43230
rect -66293 43225 -66069 43230
rect -66293 43148 -66216 43225
rect -66381 43143 -66216 43148
rect -66152 43153 -66069 43225
rect -66005 43153 -65982 43235
rect -66152 43143 -65982 43153
rect -68379 42979 -68275 42986
rect -68379 42954 -68061 42979
rect -68379 42888 -68358 42954
rect -68297 42888 -68061 42954
rect -68379 42874 -68061 42888
rect -68379 42869 -68275 42874
rect -68166 42622 -68061 42874
rect -67816 42944 -66649 43004
rect -67816 42874 -67772 42944
rect -67706 42874 -66649 42944
rect -67816 42821 -66649 42874
rect -67211 42622 -67082 42634
rect -68166 42517 -67082 42622
rect -69420 41107 -69330 41121
rect -69420 41042 -69407 41107
rect -69346 41042 -69330 41107
rect -69420 41029 -69330 41042
rect -68355 41118 -68262 41140
rect -68355 41115 -68067 41118
rect -68355 41063 -68334 41115
rect -68276 41063 -68067 41115
rect -68355 41042 -68067 41063
rect -68355 41031 -68262 41042
rect -68143 40855 -68067 41042
rect -67806 41111 -67694 41133
rect -67806 41107 -67654 41111
rect -67806 41042 -67788 41107
rect -67719 41102 -67654 41107
rect -67462 41102 -67365 41111
rect -67719 41042 -67365 41102
rect -67806 41022 -67365 41042
rect -67806 41021 -67694 41022
rect -68150 40765 -67615 40855
rect -67705 39583 -67615 40765
rect -67462 39790 -67365 41022
rect -67211 40050 -67082 42517
rect -66832 40688 -66649 42821
rect -66381 41790 -65982 43143
rect -66381 41703 -66364 41790
rect -66303 41703 -66233 41790
rect -66172 41784 -65982 41790
rect -66172 41703 -66077 41784
rect -66381 41697 -66077 41703
rect -66016 41697 -65982 41784
rect -67211 39921 -66978 40050
rect -67462 39693 -67265 39790
rect -67705 39493 -67502 39583
rect -67917 39339 -67799 39360
rect -67917 39335 -67716 39339
rect -69535 39299 -69394 39328
rect -69535 39225 -69513 39299
rect -69434 39225 -69394 39299
rect -68449 39326 -68358 39328
rect -68449 39315 -68064 39326
rect -68449 39252 -68433 39315
rect -68370 39252 -68064 39315
rect -68449 39237 -68064 39252
rect -67917 39268 -67893 39335
rect -67820 39268 -67716 39335
rect -67917 39242 -67716 39268
rect -68449 39232 -68358 39237
rect -69535 39187 -69394 39225
rect -68153 39095 -68064 39237
rect -67862 39236 -67716 39242
rect -67862 39201 -67713 39236
rect -68153 39006 -67922 39095
rect -68526 37782 -68407 37793
rect -68526 37774 -68187 37782
rect -68526 37695 -68507 37774
rect -68437 37695 -68187 37774
rect -68526 37692 -68187 37695
rect -68526 37682 -68407 37692
rect -70223 37015 -69812 37032
rect -70223 37012 -69895 37015
rect -70223 37007 -70044 37012
rect -70223 36912 -70203 37007
rect -70126 36917 -70044 37007
rect -69967 36920 -69895 37012
rect -69818 36920 -69812 37015
rect -69967 36917 -69812 36920
rect -70126 36912 -69812 36917
rect -70223 36839 -69812 36912
rect -70223 36836 -69898 36839
rect -70223 36831 -70047 36836
rect -70223 36736 -70206 36831
rect -70129 36741 -70047 36831
rect -69970 36744 -69898 36836
rect -69821 36744 -69812 36839
rect -69970 36741 -69812 36744
rect -70129 36736 -69812 36741
rect -70223 36680 -69812 36736
rect -70223 36677 -69896 36680
rect -70223 36672 -70045 36677
rect -70223 36577 -70204 36672
rect -70127 36582 -70045 36672
rect -69968 36585 -69896 36677
rect -69819 36585 -69812 36680
rect -69968 36582 -69812 36585
rect -70127 36577 -69812 36582
rect -70223 36522 -69812 36577
rect -70223 36519 -69897 36522
rect -70223 36514 -70046 36519
rect -70223 36419 -70205 36514
rect -70128 36424 -70046 36514
rect -69969 36427 -69897 36519
rect -69820 36427 -69812 36522
rect -69969 36424 -69812 36427
rect -70128 36419 -69812 36424
rect -70223 36407 -69812 36419
rect -70909 35764 -70500 35781
rect -70909 35761 -70583 35764
rect -70909 35756 -70732 35761
rect -70909 35661 -70891 35756
rect -70814 35666 -70732 35756
rect -70655 35669 -70583 35761
rect -70506 35669 -70500 35764
rect -70655 35666 -70500 35669
rect -70814 35661 -70500 35666
rect -70909 35588 -70500 35661
rect -70909 35585 -70586 35588
rect -70909 35580 -70735 35585
rect -70909 35485 -70894 35580
rect -70817 35490 -70735 35580
rect -70658 35493 -70586 35585
rect -70509 35493 -70500 35588
rect -70658 35490 -70500 35493
rect -70817 35485 -70500 35490
rect -70909 35429 -70500 35485
rect -70909 35426 -70584 35429
rect -70909 35421 -70733 35426
rect -70909 35326 -70892 35421
rect -70815 35331 -70733 35421
rect -70656 35334 -70584 35426
rect -70507 35334 -70500 35429
rect -70656 35331 -70500 35334
rect -70815 35326 -70500 35331
rect -70909 35271 -70500 35326
rect -70909 35268 -70585 35271
rect -70909 35263 -70734 35268
rect -70909 35168 -70893 35263
rect -70816 35173 -70734 35263
rect -70657 35176 -70585 35268
rect -70508 35176 -70500 35271
rect -70657 35173 -70500 35176
rect -70816 35168 -70500 35173
rect -70909 35156 -70500 35168
rect -70909 27365 -70510 35156
rect -70223 28475 -69824 36407
rect -69455 34452 -69327 34471
rect -68277 34452 -68187 37692
rect -69455 34362 -68187 34452
rect -70223 28458 -69816 28475
rect -70223 28455 -69899 28458
rect -70223 28450 -70048 28455
rect -70223 28355 -70207 28450
rect -70130 28360 -70048 28450
rect -69971 28363 -69899 28455
rect -69822 28363 -69816 28458
rect -69971 28360 -69816 28363
rect -70130 28355 -69816 28360
rect -70223 28282 -69816 28355
rect -70223 28279 -69902 28282
rect -70223 28274 -70051 28279
rect -70223 28179 -70210 28274
rect -70133 28184 -70051 28274
rect -69974 28187 -69902 28279
rect -69825 28187 -69816 28282
rect -69974 28184 -69816 28187
rect -70133 28179 -69816 28184
rect -70223 28123 -69816 28179
rect -70223 28120 -69900 28123
rect -70223 28115 -70049 28120
rect -70223 28020 -70208 28115
rect -70131 28025 -70049 28115
rect -69972 28028 -69900 28120
rect -69823 28028 -69816 28123
rect -69972 28025 -69816 28028
rect -70131 28020 -69816 28025
rect -70223 27965 -69816 28020
rect -70223 27962 -69901 27965
rect -70223 27957 -70050 27962
rect -70223 27862 -70209 27957
rect -70132 27867 -70050 27957
rect -69973 27870 -69901 27962
rect -69824 27870 -69816 27965
rect -69973 27867 -69816 27870
rect -70132 27862 -69816 27867
rect -70223 27850 -69816 27862
rect -70909 27348 -70500 27365
rect -70909 27345 -70583 27348
rect -70909 27340 -70732 27345
rect -70909 27245 -70891 27340
rect -70814 27250 -70732 27340
rect -70655 27253 -70583 27345
rect -70506 27253 -70500 27348
rect -70655 27250 -70500 27253
rect -70814 27245 -70500 27250
rect -70909 27172 -70500 27245
rect -70909 27169 -70586 27172
rect -70909 27164 -70735 27169
rect -70909 27069 -70894 27164
rect -70817 27074 -70735 27164
rect -70658 27077 -70586 27169
rect -70509 27077 -70500 27172
rect -70658 27074 -70500 27077
rect -70817 27069 -70500 27074
rect -70909 27013 -70500 27069
rect -70909 27010 -70584 27013
rect -70909 27005 -70733 27010
rect -70909 26910 -70892 27005
rect -70815 26915 -70733 27005
rect -70656 26918 -70584 27010
rect -70507 26918 -70500 27013
rect -70656 26915 -70500 26918
rect -70815 26910 -70500 26915
rect -70909 26855 -70500 26910
rect -70909 26852 -70585 26855
rect -70909 26847 -70734 26852
rect -70909 26752 -70893 26847
rect -70816 26757 -70734 26847
rect -70657 26760 -70585 26852
rect -70508 26760 -70500 26855
rect -70657 26757 -70500 26760
rect -70816 26752 -70500 26757
rect -70909 26740 -70500 26752
rect -70909 18338 -70510 26740
rect -70911 18336 -70510 18338
rect -70223 19417 -69824 27850
rect -70223 19400 -69812 19417
rect -70223 19397 -69895 19400
rect -70223 19392 -70044 19397
rect -70223 19297 -70203 19392
rect -70126 19302 -70044 19392
rect -69967 19305 -69895 19397
rect -69818 19305 -69812 19400
rect -69967 19302 -69812 19305
rect -70126 19297 -69812 19302
rect -70223 19224 -69812 19297
rect -70223 19221 -69898 19224
rect -70223 19216 -70047 19221
rect -70223 19121 -70206 19216
rect -70129 19126 -70047 19216
rect -69970 19129 -69898 19221
rect -69821 19129 -69812 19224
rect -69970 19126 -69812 19129
rect -70129 19121 -69812 19126
rect -70223 19065 -69812 19121
rect -70223 19062 -69896 19065
rect -70223 19057 -70045 19062
rect -70223 18962 -70204 19057
rect -70127 18967 -70045 19057
rect -69968 18970 -69896 19062
rect -69819 18970 -69812 19065
rect -69968 18967 -69812 18970
rect -70127 18962 -69812 18967
rect -70223 18907 -69812 18962
rect -70223 18904 -69897 18907
rect -70223 18899 -70046 18904
rect -70223 18804 -70205 18899
rect -70128 18809 -70046 18899
rect -69969 18812 -69897 18904
rect -69820 18812 -69812 18907
rect -69969 18809 -69812 18812
rect -70128 18804 -69812 18809
rect -70223 18792 -69812 18804
rect -70911 18319 -70504 18336
rect -70911 18316 -70587 18319
rect -70911 18311 -70736 18316
rect -72241 18178 -72081 18251
rect -70911 18216 -70895 18311
rect -70818 18221 -70736 18311
rect -70659 18224 -70587 18316
rect -70510 18224 -70504 18319
rect -70659 18221 -70504 18224
rect -70818 18216 -70504 18221
rect -70911 18143 -70504 18216
rect -70911 18140 -70590 18143
rect -70911 18135 -70739 18140
rect -70911 18040 -70898 18135
rect -70821 18045 -70739 18135
rect -70662 18048 -70590 18140
rect -70513 18048 -70504 18143
rect -70662 18045 -70504 18048
rect -70821 18040 -70504 18045
rect -70911 17984 -70504 18040
rect -70911 17981 -70588 17984
rect -70911 17976 -70737 17981
rect -70911 17881 -70896 17976
rect -70819 17886 -70737 17976
rect -70660 17889 -70588 17981
rect -70511 17889 -70504 17984
rect -70660 17886 -70504 17889
rect -70819 17881 -70504 17886
rect -70911 17826 -70504 17881
rect -70911 17823 -70589 17826
rect -70911 17818 -70738 17823
rect -70911 17723 -70897 17818
rect -70820 17728 -70738 17818
rect -70661 17731 -70589 17823
rect -70512 17731 -70504 17826
rect -70661 17728 -70504 17731
rect -70820 17723 -70504 17728
rect -70911 17711 -70504 17723
rect -70911 17710 -70510 17711
rect -72115 12726 -71891 12743
rect -72115 12672 -72089 12726
rect -72035 12672 -71966 12726
rect -71912 12672 -71891 12726
rect -72115 12654 -71891 12672
rect -71989 12369 -71899 12654
rect -72006 12356 -71735 12369
rect -72006 12268 -71988 12356
rect -71900 12268 -71829 12356
rect -71741 12268 -71735 12356
rect -72006 12244 -71735 12268
rect -73201 12149 -72652 12161
rect -73201 12147 -72885 12149
rect -73201 12012 -73140 12147
rect -72991 12014 -72885 12147
rect -72736 12014 -72652 12149
rect -72991 12012 -72652 12014
rect -73201 11993 -72652 12012
rect -72835 11801 -72654 11993
rect -72835 11733 -71072 11801
rect -72835 11634 -71203 11733
rect -71104 11634 -71072 11733
rect -72835 11620 -71072 11634
rect -71216 11580 -71073 11620
rect -71216 11486 -71185 11580
rect -71100 11486 -71073 11580
rect -71216 11460 -71073 11486
rect -71933 11310 -71466 11335
rect -71933 11197 -71904 11310
rect -71787 11307 -71466 11310
rect -71787 11197 -71610 11307
rect -71933 11194 -71610 11197
rect -71493 11194 -71466 11307
rect -71933 11012 -71466 11194
rect -71933 10899 -71907 11012
rect -71790 10899 -71617 11012
rect -71500 10899 -71466 11012
rect -71933 10868 -71466 10899
rect -70909 6169 -70510 17710
rect -70915 6167 -70510 6169
rect -70223 7397 -69824 18792
rect -70223 7380 -69812 7397
rect -70223 7377 -69895 7380
rect -70223 7372 -70044 7377
rect -70223 7277 -70203 7372
rect -70126 7282 -70044 7372
rect -69967 7285 -69895 7377
rect -69818 7285 -69812 7380
rect -69967 7282 -69812 7285
rect -70126 7277 -69812 7282
rect -70223 7204 -69812 7277
rect -70223 7201 -69898 7204
rect -70223 7196 -70047 7201
rect -70223 7101 -70206 7196
rect -70129 7106 -70047 7196
rect -69970 7109 -69898 7201
rect -69821 7109 -69812 7204
rect -69970 7106 -69812 7109
rect -70129 7101 -69812 7106
rect -70223 7045 -69812 7101
rect -70223 7042 -69896 7045
rect -70223 7037 -70045 7042
rect -70223 6942 -70204 7037
rect -70127 6947 -70045 7037
rect -69968 6950 -69896 7042
rect -69819 6950 -69812 7045
rect -69968 6947 -69812 6950
rect -70127 6942 -69812 6947
rect -70223 6887 -69812 6942
rect -70223 6884 -69897 6887
rect -70223 6879 -70046 6884
rect -70223 6784 -70205 6879
rect -70128 6789 -70046 6879
rect -69969 6792 -69897 6884
rect -69820 6792 -69812 6887
rect -69969 6789 -69812 6792
rect -70128 6784 -69812 6789
rect -70223 6772 -69812 6784
rect -70915 6150 -70508 6167
rect -70915 6147 -70591 6150
rect -70915 6142 -70740 6147
rect -70915 6047 -70899 6142
rect -70822 6052 -70740 6142
rect -70663 6055 -70591 6147
rect -70514 6055 -70508 6150
rect -70663 6052 -70508 6055
rect -70822 6047 -70508 6052
rect -70915 5974 -70508 6047
rect -70915 5971 -70594 5974
rect -70915 5966 -70743 5971
rect -70915 5871 -70902 5966
rect -70825 5876 -70743 5966
rect -70666 5879 -70594 5971
rect -70517 5879 -70508 5974
rect -70666 5876 -70508 5879
rect -70825 5871 -70508 5876
rect -70915 5815 -70508 5871
rect -70915 5812 -70592 5815
rect -70915 5807 -70741 5812
rect -70915 5712 -70900 5807
rect -70823 5717 -70741 5807
rect -70664 5720 -70592 5812
rect -70515 5720 -70508 5815
rect -70664 5717 -70508 5720
rect -70823 5712 -70508 5717
rect -70915 5657 -70508 5712
rect -70915 5654 -70593 5657
rect -70915 5649 -70742 5654
rect -70915 5554 -70901 5649
rect -70824 5559 -70742 5649
rect -70665 5562 -70593 5654
rect -70516 5562 -70508 5657
rect -70665 5559 -70508 5562
rect -70824 5554 -70508 5559
rect -70915 5542 -70508 5554
rect -70915 5541 -70510 5542
rect -70909 -3525 -70510 5541
rect -70223 -2444 -69824 6772
rect -70223 -2461 -69812 -2444
rect -70223 -2464 -69895 -2461
rect -70223 -2469 -70044 -2464
rect -70223 -2564 -70203 -2469
rect -70126 -2559 -70044 -2469
rect -69967 -2556 -69895 -2464
rect -69818 -2556 -69812 -2461
rect -69967 -2559 -69812 -2556
rect -70126 -2564 -69812 -2559
rect -70223 -2637 -69812 -2564
rect -70223 -2640 -69898 -2637
rect -70223 -2645 -70047 -2640
rect -70223 -2740 -70206 -2645
rect -70129 -2735 -70047 -2645
rect -69970 -2732 -69898 -2640
rect -69821 -2732 -69812 -2637
rect -69970 -2735 -69812 -2732
rect -70129 -2740 -69812 -2735
rect -70223 -2796 -69812 -2740
rect -70223 -2799 -69896 -2796
rect -70223 -2804 -70045 -2799
rect -70223 -2899 -70204 -2804
rect -70127 -2894 -70045 -2804
rect -69968 -2891 -69896 -2799
rect -69819 -2891 -69812 -2796
rect -69968 -2894 -69812 -2891
rect -70127 -2899 -69812 -2894
rect -70223 -2954 -69812 -2899
rect -70223 -2957 -69897 -2954
rect -70223 -2962 -70046 -2957
rect -70223 -3057 -70205 -2962
rect -70128 -3052 -70046 -2962
rect -69969 -3049 -69897 -2957
rect -69820 -3049 -69812 -2954
rect -69969 -3052 -69812 -3049
rect -70128 -3057 -69812 -3052
rect -70223 -3069 -69812 -3057
rect -70909 -3542 -70500 -3525
rect -70909 -3545 -70583 -3542
rect -70909 -3550 -70732 -3545
rect -70909 -3645 -70891 -3550
rect -70814 -3640 -70732 -3550
rect -70655 -3637 -70583 -3545
rect -70506 -3637 -70500 -3542
rect -70655 -3640 -70500 -3637
rect -70814 -3645 -70500 -3640
rect -70909 -3718 -70500 -3645
rect -70909 -3721 -70586 -3718
rect -70909 -3726 -70735 -3721
rect -70909 -3821 -70894 -3726
rect -70817 -3816 -70735 -3726
rect -70658 -3813 -70586 -3721
rect -70509 -3813 -70500 -3718
rect -70658 -3816 -70500 -3813
rect -70817 -3821 -70500 -3816
rect -70909 -3877 -70500 -3821
rect -70909 -3880 -70584 -3877
rect -70909 -3885 -70733 -3880
rect -70909 -3980 -70892 -3885
rect -70815 -3975 -70733 -3885
rect -70656 -3972 -70584 -3880
rect -70507 -3972 -70500 -3877
rect -70656 -3975 -70500 -3972
rect -70815 -3980 -70500 -3975
rect -70909 -4035 -70500 -3980
rect -70909 -4038 -70585 -4035
rect -70909 -4043 -70734 -4038
rect -70909 -4138 -70893 -4043
rect -70816 -4133 -70734 -4043
rect -70657 -4130 -70585 -4038
rect -70508 -4130 -70500 -4035
rect -70657 -4133 -70500 -4130
rect -70816 -4138 -70500 -4133
rect -70909 -4150 -70500 -4138
rect -70909 -12411 -70510 -4150
rect -70223 -11367 -69824 -3069
rect -70223 -11369 -69820 -11367
rect -70223 -11386 -69808 -11369
rect -70223 -11389 -69891 -11386
rect -70223 -11394 -70040 -11389
rect -70223 -11489 -70199 -11394
rect -70122 -11484 -70040 -11394
rect -69963 -11481 -69891 -11389
rect -69814 -11481 -69808 -11386
rect -69963 -11484 -69808 -11481
rect -70122 -11489 -69808 -11484
rect -70223 -11562 -69808 -11489
rect -70223 -11565 -69894 -11562
rect -70223 -11570 -70043 -11565
rect -70223 -11665 -70202 -11570
rect -70125 -11660 -70043 -11570
rect -69966 -11657 -69894 -11565
rect -69817 -11657 -69808 -11562
rect -69966 -11660 -69808 -11657
rect -70125 -11665 -69808 -11660
rect -70223 -11721 -69808 -11665
rect -70223 -11724 -69892 -11721
rect -70223 -11729 -70041 -11724
rect -70223 -11824 -70200 -11729
rect -70123 -11819 -70041 -11729
rect -69964 -11816 -69892 -11724
rect -69815 -11816 -69808 -11721
rect -69964 -11819 -69808 -11816
rect -70123 -11824 -69808 -11819
rect -70223 -11879 -69808 -11824
rect -70223 -11882 -69893 -11879
rect -70223 -11887 -70042 -11882
rect -70223 -11982 -70201 -11887
rect -70124 -11977 -70042 -11887
rect -69965 -11974 -69893 -11882
rect -69816 -11974 -69808 -11879
rect -69965 -11977 -69808 -11974
rect -70124 -11982 -69808 -11977
rect -70223 -11994 -69808 -11982
rect -70223 -11995 -69820 -11994
rect -70909 -12413 -70508 -12411
rect -70909 -12430 -70496 -12413
rect -70909 -12433 -70579 -12430
rect -70909 -12438 -70728 -12433
rect -70909 -12533 -70887 -12438
rect -70810 -12528 -70728 -12438
rect -70651 -12525 -70579 -12433
rect -70502 -12525 -70496 -12430
rect -70651 -12528 -70496 -12525
rect -70810 -12533 -70496 -12528
rect -70909 -12606 -70496 -12533
rect -70909 -12609 -70582 -12606
rect -70909 -12614 -70731 -12609
rect -70909 -12709 -70890 -12614
rect -70813 -12704 -70731 -12614
rect -70654 -12701 -70582 -12609
rect -70505 -12701 -70496 -12606
rect -70654 -12704 -70496 -12701
rect -70813 -12709 -70496 -12704
rect -70909 -12765 -70496 -12709
rect -70909 -12768 -70580 -12765
rect -70909 -12773 -70729 -12768
rect -70909 -12868 -70888 -12773
rect -70811 -12863 -70729 -12773
rect -70652 -12860 -70580 -12768
rect -70503 -12860 -70496 -12765
rect -70652 -12863 -70496 -12860
rect -70811 -12868 -70496 -12863
rect -70909 -12923 -70496 -12868
rect -70909 -12926 -70581 -12923
rect -70909 -12931 -70730 -12926
rect -70909 -13026 -70889 -12931
rect -70812 -13021 -70730 -12931
rect -70653 -13018 -70581 -12926
rect -70504 -13018 -70496 -12923
rect -70653 -13021 -70496 -13018
rect -70812 -13026 -70496 -13021
rect -70909 -13038 -70496 -13026
rect -70909 -13039 -70508 -13038
rect -70909 -20496 -70510 -13039
rect -70911 -20498 -70510 -20496
rect -70223 -19458 -69824 -11995
rect -70223 -19475 -69812 -19458
rect -70223 -19478 -69895 -19475
rect -70223 -19483 -70044 -19478
rect -70223 -19578 -70203 -19483
rect -70126 -19573 -70044 -19483
rect -69967 -19570 -69895 -19478
rect -69818 -19570 -69812 -19475
rect -69967 -19573 -69812 -19570
rect -70126 -19578 -69812 -19573
rect -70223 -19651 -69812 -19578
rect -70223 -19654 -69898 -19651
rect -70223 -19659 -70047 -19654
rect -70223 -19754 -70206 -19659
rect -70129 -19749 -70047 -19659
rect -69970 -19746 -69898 -19654
rect -69821 -19746 -69812 -19651
rect -69970 -19749 -69812 -19746
rect -70129 -19754 -69812 -19749
rect -70223 -19810 -69812 -19754
rect -70223 -19813 -69896 -19810
rect -70223 -19818 -70045 -19813
rect -70223 -19913 -70204 -19818
rect -70127 -19908 -70045 -19818
rect -69968 -19905 -69896 -19813
rect -69819 -19905 -69812 -19810
rect -69968 -19908 -69812 -19905
rect -70127 -19913 -69812 -19908
rect -70223 -19968 -69812 -19913
rect -70223 -19971 -69897 -19968
rect -70223 -19976 -70046 -19971
rect -70223 -20071 -70205 -19976
rect -70128 -20066 -70046 -19976
rect -69969 -20063 -69897 -19971
rect -69820 -20063 -69812 -19968
rect -69969 -20066 -69812 -20063
rect -70128 -20071 -69812 -20066
rect -70223 -20083 -69812 -20071
rect -70911 -20515 -70504 -20498
rect -70911 -20518 -70587 -20515
rect -70911 -20523 -70736 -20518
rect -70911 -20618 -70895 -20523
rect -70818 -20613 -70736 -20523
rect -70659 -20610 -70587 -20518
rect -70510 -20610 -70504 -20515
rect -70659 -20613 -70504 -20610
rect -70818 -20618 -70504 -20613
rect -70911 -20691 -70504 -20618
rect -70911 -20694 -70590 -20691
rect -70911 -20699 -70739 -20694
rect -70911 -20794 -70898 -20699
rect -70821 -20789 -70739 -20699
rect -70662 -20786 -70590 -20694
rect -70513 -20786 -70504 -20691
rect -70662 -20789 -70504 -20786
rect -70821 -20794 -70504 -20789
rect -70911 -20850 -70504 -20794
rect -70911 -20853 -70588 -20850
rect -70911 -20858 -70737 -20853
rect -70911 -20953 -70896 -20858
rect -70819 -20948 -70737 -20858
rect -70660 -20945 -70588 -20853
rect -70511 -20945 -70504 -20850
rect -70660 -20948 -70504 -20945
rect -70819 -20953 -70504 -20948
rect -70911 -21008 -70504 -20953
rect -70911 -21011 -70589 -21008
rect -70911 -21016 -70738 -21011
rect -70911 -21111 -70897 -21016
rect -70820 -21106 -70738 -21016
rect -70661 -21103 -70589 -21011
rect -70512 -21103 -70504 -21008
rect -70661 -21106 -70504 -21103
rect -70820 -21111 -70504 -21106
rect -70911 -21123 -70504 -21111
rect -70911 -21124 -70510 -21123
rect -70909 -28535 -70510 -21124
rect -70223 -27506 -69824 -20083
rect -69455 -26457 -69327 34362
rect -68341 31187 -68170 31198
rect -68341 31130 -68318 31187
rect -68237 31130 -68170 31187
rect -68341 31113 -68170 31130
rect -68368 22803 -68245 22819
rect -68368 22714 -68348 22803
rect -68263 22714 -68245 22803
rect -68368 22696 -68245 22714
rect -68360 13716 -68233 13749
rect -68360 13646 -68333 13716
rect -68258 13646 -68233 13716
rect -68360 13622 -68233 13646
rect -68362 1157 -68225 1175
rect -68362 1064 -68328 1157
rect -68246 1064 -68225 1157
rect -68362 1038 -68225 1064
rect -68415 -7936 -68380 -7856
rect -68289 -7936 -68244 -7856
rect -68415 -7945 -68244 -7936
rect -68415 -8020 -68368 -7945
rect -68292 -8020 -68244 -7945
rect -68415 -8031 -68244 -8020
rect -68415 -8111 -68379 -8031
rect -68288 -8111 -68244 -8031
rect -68415 -16634 -68244 -8111
rect -68415 -16749 -68375 -16634
rect -68295 -16749 -68244 -16634
rect -68415 -16891 -68244 -16749
rect -68415 -17006 -68377 -16891
rect -68297 -17006 -68244 -16891
rect -68415 -17023 -68244 -17006
rect -68544 -23421 -68408 -23396
rect -68544 -23497 -68519 -23421
rect -68436 -23433 -68408 -23421
rect -68011 -23433 -67922 39006
rect -67798 20108 -67713 39201
rect -67592 21188 -67502 39493
rect -67362 21811 -67265 39693
rect -67107 30001 -66978 39921
rect -66815 31229 -66665 40688
rect -66381 40006 -65982 41697
rect -66381 39919 -66359 40006
rect -66299 40002 -65982 40006
rect -66299 39919 -66224 40002
rect -66381 39915 -66224 39919
rect -66164 40001 -65982 40002
rect -66164 39915 -66089 40001
rect -66381 39914 -66089 39915
rect -66029 39914 -65982 40001
rect -66381 38450 -65982 39914
rect -66381 38448 -66064 38450
rect -66381 38447 -66225 38448
rect -66381 38343 -66367 38447
rect -66304 38344 -66225 38447
rect -66162 38346 -66064 38448
rect -66001 38346 -65982 38450
rect -66162 38344 -65982 38346
rect -66304 38343 -65982 38344
rect -66381 33652 -65982 38343
rect -66381 33649 -66221 33652
rect -66381 33586 -66353 33649
rect -66293 33589 -66221 33649
rect -66161 33649 -65982 33652
rect -66161 33589 -66087 33649
rect -66293 33586 -66087 33589
rect -66027 33586 -65982 33649
rect -66815 31186 -66583 31229
rect -66815 31115 -66690 31186
rect -66620 31115 -66583 31186
rect -66815 31079 -66583 31115
rect -66897 30001 -66741 30014
rect -67107 29872 -66741 30001
rect -66897 22858 -66741 29872
rect -66381 23723 -65982 33586
rect -66381 23720 -66231 23723
rect -66381 23657 -66363 23720
rect -66303 23660 -66231 23720
rect -66171 23720 -65982 23723
rect -66171 23660 -66097 23720
rect -66303 23657 -66097 23660
rect -66037 23657 -65982 23720
rect -66897 22822 -66566 22858
rect -66897 22748 -66681 22822
rect -66602 22748 -66566 22822
rect -66897 22702 -66566 22748
rect -67362 21714 -67123 21811
rect -67610 21171 -67487 21188
rect -67610 21081 -67592 21171
rect -67502 21081 -67487 21171
rect -67610 21058 -67487 21081
rect -67220 20508 -67123 21714
rect -67345 20478 -67123 20508
rect -67385 20411 -67123 20478
rect -66929 21170 -66806 21188
rect -66929 21082 -66912 21170
rect -66824 21082 -66806 21170
rect -67798 20072 -67613 20108
rect -67798 20023 -67585 20072
rect -67725 -248 -67585 20023
rect -67385 12113 -67206 20411
rect -66929 13755 -66806 21082
rect -66381 16081 -65982 23657
rect -66381 16078 -66231 16081
rect -66381 16015 -66363 16078
rect -66303 16018 -66231 16078
rect -66171 16078 -65982 16081
rect -66171 16018 -66097 16078
rect -66303 16015 -66097 16018
rect -66037 16015 -65982 16078
rect -66929 13747 -66761 13755
rect -66929 13709 -66590 13747
rect -66929 13646 -66686 13709
rect -66620 13646 -66590 13709
rect -66929 13616 -66590 13646
rect -66770 13614 -66590 13616
rect -67385 11934 -66783 12113
rect -66962 1229 -66783 11934
rect -66381 12048 -65982 16015
rect -66381 11976 -66370 12048
rect -66308 11976 -66255 12048
rect -66193 11976 -66141 12048
rect -66079 11976 -65982 12048
rect -66381 10444 -65982 11976
rect -66381 10443 -66095 10444
rect -66381 10387 -66361 10443
rect -66308 10387 -66251 10443
rect -66198 10388 -66095 10443
rect -66042 10388 -65982 10444
rect -66198 10387 -65982 10388
rect -66381 9528 -65982 10387
rect -66381 9527 -66110 9528
rect -66381 9471 -66359 9527
rect -66306 9526 -66110 9527
rect -66306 9471 -66231 9526
rect -66381 9470 -66231 9471
rect -66178 9472 -66110 9526
rect -66057 9472 -65982 9528
rect -66178 9470 -65982 9472
rect -66381 8621 -65982 9470
rect -66381 8619 -66077 8621
rect -66381 8617 -66224 8619
rect -66381 8561 -66360 8617
rect -66307 8563 -66224 8617
rect -66171 8565 -66077 8619
rect -66024 8565 -65982 8621
rect -66171 8563 -65982 8565
rect -66307 8561 -65982 8563
rect -66381 7703 -65982 8561
rect -66381 7696 -66199 7703
rect -66381 7640 -66357 7696
rect -66304 7647 -66199 7696
rect -66146 7701 -65982 7703
rect -66146 7647 -66063 7701
rect -66304 7645 -66063 7647
rect -66010 7645 -65982 7701
rect -66304 7640 -65982 7645
rect -66381 6793 -65982 7640
rect -66381 6792 -66090 6793
rect -66381 6786 -66232 6792
rect -66381 6730 -66365 6786
rect -66312 6736 -66232 6786
rect -66179 6737 -66090 6792
rect -66037 6737 -65982 6793
rect -66179 6736 -65982 6737
rect -66312 6730 -65982 6736
rect -66381 5868 -65982 6730
rect -66381 5812 -66355 5868
rect -66302 5866 -65982 5868
rect -66302 5865 -66084 5866
rect -66302 5812 -66221 5865
rect -66381 5809 -66221 5812
rect -66168 5810 -66084 5865
rect -66031 5810 -65982 5866
rect -66168 5809 -65982 5810
rect -66381 3775 -65982 5809
rect -66381 3772 -66221 3775
rect -66381 3709 -66353 3772
rect -66293 3712 -66221 3772
rect -66161 3772 -65982 3775
rect -66161 3712 -66087 3772
rect -66293 3709 -66087 3712
rect -66027 3709 -65982 3772
rect -66381 2027 -65982 3709
rect -66381 2021 -66223 2027
rect -66381 1926 -66367 2021
rect -66301 1932 -66223 2021
rect -66157 1932 -66064 2027
rect -65998 1932 -65982 2027
rect -66301 1926 -65982 1932
rect -66962 1148 -66576 1229
rect -66962 1083 -66723 1148
rect -66653 1083 -66576 1148
rect -66962 1050 -66576 1083
rect -66947 -248 -66756 -222
rect -67725 -388 -66756 -248
rect -66947 -7893 -66756 -388
rect -66381 -5738 -65982 1926
rect -66381 -5741 -66224 -5738
rect -66381 -5804 -66356 -5741
rect -66296 -5801 -66224 -5741
rect -66164 -5741 -65982 -5738
rect -66164 -5801 -66090 -5741
rect -66296 -5804 -66090 -5801
rect -66030 -5804 -65982 -5741
rect -66381 -7084 -65982 -5804
rect -66381 -7088 -66070 -7084
rect -66381 -7093 -66225 -7088
rect -66381 -7181 -66367 -7093
rect -66302 -7176 -66225 -7093
rect -66160 -7172 -66070 -7088
rect -66005 -7172 -65982 -7084
rect -66160 -7176 -65982 -7172
rect -66302 -7181 -65982 -7176
rect -66947 -7948 -66582 -7893
rect -66947 -8026 -66691 -7948
rect -66618 -8026 -66582 -7948
rect -66947 -8084 -66582 -8026
rect -66381 -14518 -65982 -7181
rect -66381 -14521 -66217 -14518
rect -66381 -14584 -66349 -14521
rect -66289 -14581 -66217 -14521
rect -66157 -14521 -65982 -14518
rect -66157 -14581 -66083 -14521
rect -66289 -14584 -66083 -14581
rect -66023 -14584 -65982 -14521
rect -66381 -22611 -65982 -14584
rect -66381 -22614 -66231 -22611
rect -66381 -22677 -66363 -22614
rect -66303 -22674 -66231 -22614
rect -66171 -22614 -65982 -22611
rect -66171 -22674 -66097 -22614
rect -66303 -22677 -66097 -22674
rect -66037 -22677 -65982 -22614
rect -68436 -23497 -67922 -23433
rect -68544 -23522 -67922 -23497
rect -66896 -23417 -66736 -23397
rect -66896 -23497 -66855 -23417
rect -66759 -23497 -66736 -23417
rect -66896 -23523 -66736 -23497
rect -66381 -25615 -65982 -22677
rect -66381 -25618 -66204 -25615
rect -66381 -25702 -66369 -25618
rect -66299 -25699 -66204 -25618
rect -66134 -25699 -66063 -25615
rect -65993 -25699 -65982 -25615
rect -66299 -25702 -65982 -25699
rect -66964 -26434 -66815 -26427
rect -69455 -26477 -68488 -26457
rect -69455 -26561 -68598 -26477
rect -68504 -26561 -68488 -26477
rect -69455 -26585 -68488 -26561
rect -66964 -26469 -66756 -26434
rect -66964 -26559 -66935 -26469
rect -66854 -26559 -66756 -26469
rect -66964 -26588 -66756 -26559
rect -70223 -27523 -69812 -27506
rect -70223 -27526 -69895 -27523
rect -70223 -27531 -70044 -27526
rect -70223 -27626 -70203 -27531
rect -70126 -27621 -70044 -27531
rect -69967 -27618 -69895 -27526
rect -69818 -27618 -69812 -27523
rect -69967 -27621 -69812 -27618
rect -70126 -27626 -69812 -27621
rect -70223 -27699 -69812 -27626
rect -70223 -27702 -69898 -27699
rect -70223 -27707 -70047 -27702
rect -70223 -27802 -70206 -27707
rect -70129 -27797 -70047 -27707
rect -69970 -27794 -69898 -27702
rect -69821 -27794 -69812 -27699
rect -69970 -27797 -69812 -27794
rect -70129 -27802 -69812 -27797
rect -70223 -27858 -69812 -27802
rect -70223 -27861 -69896 -27858
rect -70223 -27866 -70045 -27861
rect -70223 -27961 -70204 -27866
rect -70127 -27956 -70045 -27866
rect -69968 -27953 -69896 -27861
rect -69819 -27953 -69812 -27858
rect -69968 -27956 -69812 -27953
rect -70127 -27961 -69812 -27956
rect -70223 -28016 -69812 -27961
rect -70223 -28019 -69897 -28016
rect -70223 -28024 -70046 -28019
rect -70223 -28119 -70205 -28024
rect -70128 -28114 -70046 -28024
rect -69969 -28111 -69897 -28019
rect -69820 -28111 -69812 -28016
rect -69969 -28114 -69812 -28111
rect -70128 -28119 -69812 -28114
rect -70223 -28131 -69812 -28119
rect -70909 -28537 -70508 -28535
rect -70909 -28554 -70496 -28537
rect -70909 -28557 -70579 -28554
rect -70909 -28562 -70728 -28557
rect -70909 -28657 -70887 -28562
rect -70810 -28652 -70728 -28562
rect -70651 -28649 -70579 -28557
rect -70502 -28649 -70496 -28554
rect -70651 -28652 -70496 -28649
rect -70810 -28657 -70496 -28652
rect -70909 -28730 -70496 -28657
rect -70909 -28733 -70582 -28730
rect -70909 -28738 -70731 -28733
rect -70909 -28833 -70890 -28738
rect -70813 -28828 -70731 -28738
rect -70654 -28825 -70582 -28733
rect -70505 -28825 -70496 -28730
rect -70654 -28828 -70496 -28825
rect -70813 -28833 -70496 -28828
rect -70909 -28889 -70496 -28833
rect -70909 -28892 -70580 -28889
rect -70909 -28897 -70729 -28892
rect -70909 -28992 -70888 -28897
rect -70811 -28987 -70729 -28897
rect -70652 -28984 -70580 -28892
rect -70503 -28984 -70496 -28889
rect -70652 -28987 -70496 -28984
rect -70811 -28992 -70496 -28987
rect -70909 -29047 -70496 -28992
rect -70909 -29050 -70581 -29047
rect -70909 -29055 -70730 -29050
rect -70909 -29150 -70889 -29055
rect -70812 -29145 -70730 -29055
rect -70653 -29142 -70581 -29050
rect -70504 -29142 -70496 -29047
rect -70653 -29145 -70496 -29142
rect -70812 -29150 -70496 -29145
rect -70909 -29162 -70496 -29150
rect -70909 -29163 -70508 -29162
rect -70909 -38193 -70510 -29163
rect -70223 -38193 -69824 -28131
rect -66963 -29093 -66756 -26588
rect -66381 -30037 -65982 -25702
rect -66381 -30044 -66217 -30037
rect -66381 -30126 -66366 -30044
rect -66289 -30119 -66217 -30044
rect -66140 -30038 -65982 -30037
rect -66140 -30119 -66067 -30038
rect -66289 -30120 -66067 -30119
rect -65990 -30120 -65982 -30038
rect -66289 -30126 -65982 -30120
rect -66381 -31013 -65982 -30126
rect -66381 -31015 -66108 -31013
rect -66381 -31018 -66256 -31015
rect -66381 -31079 -66369 -31018
rect -66310 -31076 -66256 -31018
rect -66197 -31074 -66108 -31015
rect -66049 -31074 -65982 -31013
rect -66197 -31076 -65982 -31074
rect -66310 -31079 -65982 -31076
rect -66381 -32494 -65982 -31079
rect -66381 -32507 -66098 -32494
rect -66381 -32509 -66231 -32507
rect -66381 -32570 -66371 -32509
rect -66312 -32568 -66231 -32509
rect -66172 -32555 -66098 -32507
rect -66039 -32555 -65982 -32494
rect -66172 -32568 -65982 -32555
rect -66312 -32570 -65982 -32568
rect -66381 -33681 -65982 -32570
rect -66381 -33683 -66078 -33681
rect -66381 -33744 -66369 -33683
rect -66310 -33744 -66216 -33683
rect -66157 -33742 -66078 -33683
rect -66019 -33742 -65982 -33681
rect -66157 -33744 -65982 -33742
rect -66381 -37536 -65982 -33744
rect -65695 48887 -65296 55224
rect -55938 54813 -55539 55873
rect -55294 55848 -54895 55873
rect -55294 55831 -54883 55848
rect -55294 55828 -54966 55831
rect -55294 55823 -55115 55828
rect -55294 55728 -55274 55823
rect -55197 55733 -55115 55823
rect -55038 55736 -54966 55828
rect -54889 55736 -54883 55831
rect -55038 55733 -54883 55736
rect -55197 55728 -54883 55733
rect -55294 55655 -54883 55728
rect -55294 55652 -54969 55655
rect -55294 55647 -55118 55652
rect -55294 55552 -55277 55647
rect -55200 55557 -55118 55647
rect -55041 55560 -54969 55652
rect -54892 55560 -54883 55655
rect -55041 55557 -54883 55560
rect -55200 55552 -54883 55557
rect -55294 55496 -54883 55552
rect -55294 55493 -54967 55496
rect -55294 55488 -55116 55493
rect -55294 55393 -55275 55488
rect -55198 55398 -55116 55488
rect -55039 55401 -54967 55493
rect -54890 55401 -54883 55496
rect -55039 55398 -54883 55401
rect -55198 55393 -54883 55398
rect -55294 55338 -54883 55393
rect -55294 55335 -54968 55338
rect -55294 55330 -55117 55335
rect -55294 55235 -55276 55330
rect -55199 55240 -55117 55330
rect -55040 55243 -54968 55335
rect -54891 55243 -54883 55338
rect -55040 55240 -54883 55243
rect -55199 55235 -54883 55240
rect -55294 55223 -54883 55235
rect -55941 54796 -55531 54813
rect -55941 54793 -55614 54796
rect -55941 54788 -55763 54793
rect -55941 54693 -55922 54788
rect -55845 54698 -55763 54788
rect -55686 54701 -55614 54793
rect -55537 54701 -55531 54796
rect -55686 54698 -55531 54701
rect -55845 54693 -55531 54698
rect -55941 54620 -55531 54693
rect -55941 54617 -55617 54620
rect -55941 54612 -55766 54617
rect -55941 54517 -55925 54612
rect -55848 54522 -55766 54612
rect -55689 54525 -55617 54617
rect -55540 54525 -55531 54620
rect -55689 54522 -55531 54525
rect -55848 54517 -55531 54522
rect -55941 54461 -55531 54517
rect -55941 54458 -55615 54461
rect -55941 54453 -55764 54458
rect -55941 54358 -55923 54453
rect -55846 54363 -55764 54453
rect -55687 54366 -55615 54458
rect -55538 54366 -55531 54461
rect -55687 54363 -55531 54366
rect -55846 54358 -55531 54363
rect -55941 54303 -55531 54358
rect -55941 54300 -55616 54303
rect -55941 54295 -55765 54300
rect -55941 54200 -55924 54295
rect -55847 54205 -55765 54295
rect -55688 54208 -55616 54300
rect -55539 54208 -55531 54303
rect -55688 54205 -55531 54208
rect -55847 54200 -55531 54205
rect -55941 54188 -55531 54200
rect -65695 48885 -65393 48887
rect -65695 48827 -65668 48885
rect -65603 48883 -65393 48885
rect -65603 48827 -65525 48883
rect -65695 48825 -65525 48827
rect -65460 48829 -65393 48883
rect -65328 48829 -65296 48887
rect -65460 48825 -65296 48829
rect -65695 47416 -65296 48825
rect -65695 47415 -65377 47416
rect -65695 47357 -65661 47415
rect -65596 47412 -65377 47415
rect -65596 47357 -65522 47412
rect -65695 47354 -65522 47357
rect -65457 47358 -65377 47412
rect -65312 47358 -65296 47416
rect -65457 47354 -65296 47358
rect -65695 45969 -65296 47354
rect -65695 45960 -65383 45969
rect -65695 45959 -65526 45960
rect -65695 45901 -65667 45959
rect -65602 45902 -65526 45959
rect -65461 45911 -65383 45960
rect -65318 45911 -65296 45969
rect -65461 45902 -65296 45911
rect -65602 45901 -65296 45902
rect -65695 42502 -65296 45901
rect -65695 42501 -65415 42502
rect -65695 42498 -65547 42501
rect -65695 42425 -65689 42498
rect -65623 42428 -65547 42498
rect -65481 42429 -65415 42501
rect -65349 42429 -65296 42502
rect -65481 42428 -65296 42429
rect -65623 42425 -65296 42428
rect -65695 40534 -65296 42425
rect -55938 50421 -55539 54188
rect -55938 50418 -55769 50421
rect -55938 50355 -55901 50418
rect -55841 50358 -55769 50418
rect -55709 50418 -55539 50421
rect -55709 50358 -55635 50418
rect -55841 50355 -55635 50358
rect -55575 50355 -55539 50418
rect -55938 42094 -55539 50355
rect -55938 42090 -55633 42094
rect -55938 42086 -55769 42090
rect -55938 42015 -55907 42086
rect -55849 42019 -55769 42086
rect -55711 42023 -55633 42090
rect -55575 42023 -55539 42094
rect -55711 42019 -55539 42023
rect -55849 42015 -55539 42019
rect -63615 40954 -63448 40988
rect -63615 40847 -63590 40954
rect -63479 40847 -63448 40954
rect -63615 40821 -63448 40847
rect -65695 40529 -65549 40534
rect -65695 40444 -65678 40529
rect -65617 40449 -65549 40529
rect -65488 40531 -65296 40534
rect -65488 40449 -65389 40531
rect -65617 40446 -65389 40449
rect -65328 40446 -65296 40531
rect -65617 40444 -65296 40446
rect -65695 38754 -65296 40444
rect -63128 39017 -62961 39051
rect -63128 38910 -63103 39017
rect -62992 38910 -62961 39017
rect -63128 38884 -62961 38910
rect -65695 38746 -65373 38754
rect -65695 38659 -65682 38746
rect -65622 38745 -65373 38746
rect -65622 38659 -65525 38745
rect -65695 38658 -65525 38659
rect -65465 38667 -65373 38745
rect -65313 38667 -65296 38754
rect -65465 38658 -65296 38667
rect -65695 37197 -65296 38658
rect -65695 37192 -65375 37197
rect -65695 37101 -65682 37192
rect -65614 37101 -65528 37192
rect -65460 37106 -65375 37192
rect -65307 37106 -65296 37197
rect -65460 37101 -65296 37106
rect -65695 34613 -65296 37101
rect -56592 37020 -56484 37054
rect -56592 36925 -56569 37020
rect -56492 36925 -56484 37020
rect -56592 36844 -56484 36925
rect -65695 34610 -65386 34613
rect -65695 34510 -65680 34610
rect -65606 34510 -65534 34610
rect -65460 34513 -65386 34610
rect -65312 34513 -65296 34613
rect -65460 34510 -65296 34513
rect -65695 30906 -65296 34510
rect -65695 30903 -65547 30906
rect -65695 30840 -65679 30903
rect -65619 30843 -65547 30903
rect -65487 30903 -65296 30906
rect -65487 30843 -65413 30903
rect -65619 30840 -65413 30843
rect -65353 30840 -65296 30903
rect -65695 21294 -65296 30840
rect -65695 21291 -65540 21294
rect -65695 21228 -65672 21291
rect -65612 21231 -65540 21291
rect -65480 21291 -65296 21294
rect -65480 21231 -65406 21291
rect -65612 21228 -65406 21231
rect -65346 21228 -65296 21291
rect -65695 17034 -65296 21228
rect -65695 17029 -65523 17034
rect -65695 16946 -65684 17029
rect -65623 16951 -65523 17029
rect -65462 17029 -65296 17034
rect -65462 16951 -65391 17029
rect -65623 16946 -65391 16951
rect -65330 16946 -65296 17029
rect -65695 13338 -65296 16946
rect -65695 13335 -65540 13338
rect -65695 13272 -65672 13335
rect -65612 13275 -65540 13335
rect -65480 13335 -65296 13338
rect -65480 13275 -65406 13335
rect -65612 13272 -65406 13275
rect -65346 13272 -65296 13335
rect -65695 9763 -65296 13272
rect -65695 9761 -65402 9763
rect -65695 9757 -65534 9761
rect -65695 9701 -65679 9757
rect -65626 9705 -65534 9757
rect -65481 9707 -65402 9761
rect -65349 9707 -65296 9763
rect -65481 9705 -65296 9707
rect -65626 9701 -65296 9705
rect -65695 8844 -65296 9701
rect -65695 8840 -65529 8844
rect -65695 8784 -65671 8840
rect -65618 8788 -65529 8840
rect -65476 8843 -65296 8844
rect -65476 8788 -65391 8843
rect -65618 8787 -65391 8788
rect -65338 8787 -65296 8843
rect -65618 8784 -65296 8787
rect -65695 7921 -65296 8784
rect -65695 7919 -65388 7921
rect -65695 7917 -65538 7919
rect -65695 7861 -65672 7917
rect -65619 7863 -65538 7917
rect -65485 7865 -65388 7919
rect -65335 7865 -65296 7921
rect -65485 7863 -65296 7865
rect -65619 7861 -65296 7863
rect -65695 7032 -65296 7861
rect -65695 7022 -65554 7032
rect -65695 6966 -65673 7022
rect -65620 6976 -65554 7022
rect -65501 6976 -65408 7032
rect -65355 6976 -65296 7032
rect -65620 6966 -65296 6976
rect -65695 6093 -65296 6966
rect -65695 6091 -65403 6093
rect -65695 6089 -65539 6091
rect -65695 6033 -65664 6089
rect -65611 6035 -65539 6089
rect -65486 6037 -65403 6091
rect -65350 6037 -65296 6093
rect -65486 6035 -65296 6037
rect -65611 6033 -65296 6035
rect -65695 5178 -65296 6033
rect -65695 5175 -65537 5178
rect -65695 5119 -65678 5175
rect -65625 5122 -65537 5175
rect -65484 5122 -65390 5178
rect -65337 5122 -65296 5178
rect -65625 5119 -65296 5122
rect -65695 1025 -65296 5119
rect -65695 1022 -65530 1025
rect -65695 959 -65662 1022
rect -65602 962 -65530 1022
rect -65470 1022 -65296 1025
rect -65470 962 -65396 1022
rect -65602 959 -65396 962
rect -65336 959 -65296 1022
rect -65695 504 -65296 959
rect -65695 502 -65402 504
rect -65695 423 -65682 502
rect -65622 423 -65546 502
rect -65486 425 -65402 502
rect -65342 425 -65296 504
rect -65486 423 -65296 425
rect -65695 -684 -65296 423
rect -65695 -688 -65385 -684
rect -65695 -695 -65518 -688
rect -65695 -808 -65671 -695
rect -65594 -801 -65518 -695
rect -65441 -797 -65385 -688
rect -65308 -797 -65296 -684
rect -65441 -801 -65296 -797
rect -65594 -808 -65296 -801
rect -65695 -4824 -65296 -808
rect -64663 36665 -64523 36758
rect -64663 36585 -64629 36665
rect -64549 36585 -64523 36665
rect -64663 36486 -64523 36585
rect -64663 36406 -64628 36486
rect -64548 36406 -64523 36486
rect -64663 32263 -64523 36406
rect -56592 36749 -56572 36844
rect -56495 36749 -56484 36844
rect -56592 36685 -56484 36749
rect -56592 36590 -56570 36685
rect -56493 36590 -56484 36685
rect -56592 36527 -56484 36590
rect -56592 36432 -56571 36527
rect -56494 36432 -56484 36527
rect -64663 32148 -64642 32263
rect -64555 32148 -64523 32263
rect -64663 32030 -64523 32148
rect -64663 31915 -64637 32030
rect -64550 31915 -64523 32030
rect -64663 17925 -64523 31915
rect -64663 17820 -64639 17925
rect -64565 17820 -64523 17925
rect -64663 17708 -64523 17820
rect -64663 17603 -64633 17708
rect -64559 17603 -64523 17708
rect -64663 14728 -64523 17603
rect -64663 14668 -64608 14728
rect -64544 14668 -64523 14728
rect -64663 14560 -64523 14668
rect -64663 14500 -64607 14560
rect -64543 14500 -64523 14560
rect -64663 2522 -64523 14500
rect -64388 36297 -64295 36335
rect -64388 36225 -64379 36297
rect -64303 36225 -64295 36297
rect -64388 36132 -64295 36225
rect -64388 36060 -64380 36132
rect -64304 36060 -64295 36132
rect -64388 30033 -64295 36060
rect -64388 29974 -64374 30033
rect -64315 29974 -64295 30033
rect -64388 29884 -64295 29974
rect -64388 29825 -64376 29884
rect -64317 29825 -64295 29884
rect -64388 26583 -64295 29825
rect -64388 26530 -64367 26583
rect -64313 26530 -64295 26583
rect -64388 26476 -64295 26530
rect -64388 26423 -64368 26476
rect -64314 26423 -64295 26476
rect -64388 26368 -64295 26423
rect -64388 26315 -64370 26368
rect -64316 26315 -64295 26368
rect -64388 12450 -64295 26315
rect -64388 12389 -64372 12450
rect -64311 12389 -64295 12450
rect -64388 12315 -64295 12389
rect -64388 12254 -64373 12315
rect -64312 12254 -64295 12315
rect -64663 2456 -64521 2522
rect -64663 2391 -64601 2456
rect -64545 2391 -64521 2456
rect -64663 2293 -64521 2391
rect -64663 2228 -64600 2293
rect -64544 2228 -64521 2293
rect -64663 2095 -64521 2228
rect -64663 -1543 -64530 2095
rect -64388 240 -64295 12254
rect -64142 36119 -64035 36137
rect -64142 36040 -64121 36119
rect -64046 36040 -64035 36119
rect -64142 35943 -64035 36040
rect -64142 35864 -64126 35943
rect -64051 35864 -64035 35943
rect -64142 30524 -64035 35864
rect -56795 35763 -56690 35807
rect -56795 35668 -56777 35763
rect -56700 35668 -56690 35763
rect -56795 35587 -56690 35668
rect -56795 35492 -56780 35587
rect -56703 35492 -56690 35587
rect -56795 35428 -56690 35492
rect -56795 35333 -56778 35428
rect -56701 35333 -56690 35428
rect -56795 35270 -56690 35333
rect -56795 35175 -56779 35270
rect -56702 35175 -56690 35270
rect -56795 34204 -56690 35175
rect -56592 34188 -56484 36432
rect -55938 33662 -55539 42015
rect -55938 33658 -55639 33662
rect -55938 33577 -55922 33658
rect -55854 33577 -55779 33658
rect -55711 33581 -55639 33658
rect -55571 33581 -55539 33662
rect -55711 33577 -55539 33581
rect -63376 33288 -63253 33302
rect -63376 33209 -63356 33288
rect -63265 33209 -63253 33288
rect -63376 33136 -63253 33209
rect -63376 33057 -63360 33136
rect -63269 33057 -63253 33136
rect -63376 33045 -63253 33057
rect -61049 32709 -60993 32928
rect -61038 32026 -60982 32271
rect -63789 31350 -63666 31364
rect -63789 31271 -63769 31350
rect -63678 31271 -63666 31350
rect -63789 31198 -63666 31271
rect -63789 31119 -63773 31198
rect -63682 31119 -63666 31198
rect -63789 31107 -63666 31119
rect -64142 30417 -63349 30524
rect -64142 25870 -64035 30417
rect -60997 29686 -60940 29932
rect -64142 25813 -64112 25870
rect -64054 25813 -64035 25870
rect -64142 25758 -64035 25813
rect -64142 25701 -64113 25758
rect -64055 25701 -64035 25758
rect -64142 25645 -64035 25701
rect -64142 25588 -64114 25645
rect -64056 25588 -64035 25645
rect -64142 12972 -64035 25588
rect -62655 24045 -62599 24203
rect -55938 23636 -55539 33577
rect -55938 23633 -55653 23636
rect -55938 23630 -55787 23633
rect -55938 23572 -55922 23630
rect -55864 23575 -55787 23630
rect -55729 23578 -55653 23633
rect -55595 23578 -55539 23636
rect -55729 23575 -55539 23578
rect -55864 23572 -55539 23575
rect -63269 22892 -63213 23004
rect -62205 21806 -62149 21941
rect -56573 19435 -56465 19449
rect -56575 19409 -56465 19435
rect -56575 19314 -56557 19409
rect -56480 19314 -56465 19409
rect -56575 19233 -56465 19314
rect -56575 19138 -56560 19233
rect -56483 19138 -56465 19233
rect -56575 19074 -56465 19138
rect -56575 18979 -56558 19074
rect -56481 18979 -56465 19074
rect -56575 18916 -56465 18979
rect -56575 18821 -56559 18916
rect -56482 18821 -56465 18916
rect -56575 18798 -56465 18821
rect -56776 18352 -56671 18371
rect -56776 18326 -56669 18352
rect -56776 18231 -56752 18326
rect -56675 18231 -56669 18326
rect -56776 18150 -56669 18231
rect -56776 18055 -56755 18150
rect -56678 18055 -56669 18150
rect -56776 17991 -56669 18055
rect -56776 17896 -56753 17991
rect -56676 17896 -56669 17991
rect -56776 17833 -56669 17896
rect -56776 17738 -56754 17833
rect -56677 17738 -56669 17833
rect -56776 17715 -56669 17738
rect -56776 16725 -56671 17715
rect -56573 16660 -56465 18798
rect -55938 16379 -55539 23572
rect -55938 16288 -55926 16379
rect -55850 16378 -55633 16379
rect -55850 16288 -55784 16378
rect -55938 16287 -55784 16288
rect -55708 16288 -55633 16378
rect -55557 16288 -55539 16379
rect -55708 16287 -55539 16288
rect -63334 15703 -63247 15724
rect -63334 15647 -63321 15703
rect -63265 15647 -63247 15703
rect -63334 15592 -63247 15647
rect -63334 15536 -63325 15592
rect -63269 15536 -63247 15592
rect -63334 15521 -63247 15536
rect -61030 14972 -60974 15210
rect -61027 14468 -60971 14696
rect -63624 13763 -63537 13784
rect -63624 13707 -63611 13763
rect -63555 13707 -63537 13763
rect -63624 13652 -63537 13707
rect -63624 13596 -63615 13652
rect -63559 13596 -63537 13652
rect -63624 13581 -63537 13596
rect -64142 12865 -63325 12972
rect -64142 635 -64035 12865
rect -60978 12120 -60921 12368
rect -56591 7396 -56483 7432
rect -56591 7301 -56569 7396
rect -56492 7301 -56483 7396
rect -56591 7220 -56483 7301
rect -56591 7125 -56572 7220
rect -56495 7125 -56483 7220
rect -56591 7061 -56483 7125
rect -56591 6966 -56570 7061
rect -56493 6966 -56483 7061
rect -56591 6903 -56483 6966
rect -56591 6808 -56571 6903
rect -56494 6808 -56483 6903
rect -56794 6157 -56689 6202
rect -56794 6062 -56773 6157
rect -56696 6062 -56689 6157
rect -56794 5981 -56689 6062
rect -56794 5886 -56776 5981
rect -56699 5886 -56689 5981
rect -56794 5822 -56689 5886
rect -56794 5727 -56774 5822
rect -56697 5727 -56689 5822
rect -56794 5664 -56689 5727
rect -56794 5569 -56775 5664
rect -56698 5569 -56689 5664
rect -56794 4456 -56689 5569
rect -56591 4379 -56483 6808
rect -55938 3439 -55539 16287
rect -55938 3435 -55642 3439
rect -63342 3380 -63255 3401
rect -63342 3324 -63329 3380
rect -63273 3324 -63255 3380
rect -63342 3269 -63255 3324
rect -63342 3213 -63333 3269
rect -63277 3213 -63255 3269
rect -63342 3198 -63255 3213
rect -55938 3358 -55918 3435
rect -55853 3358 -55783 3435
rect -55718 3362 -55642 3435
rect -55577 3362 -55539 3439
rect -55718 3358 -55539 3362
rect -61048 2635 -60992 2855
rect -61045 2154 -60989 2379
rect -63755 1410 -63668 1431
rect -63755 1354 -63742 1410
rect -63686 1354 -63668 1410
rect -63755 1299 -63668 1354
rect -63755 1243 -63746 1299
rect -63690 1243 -63668 1299
rect -63755 1228 -63668 1243
rect -64142 528 -63346 635
rect -64388 183 -64360 240
rect -64306 183 -64295 240
rect -64388 93 -64295 183
rect -64388 36 -64364 93
rect -64310 36 -64295 93
rect -64388 8 -64295 36
rect -60996 -195 -60939 55
rect -65695 -4829 -65400 -4824
rect -65695 -4832 -65551 -4829
rect -65695 -4911 -65684 -4832
rect -65618 -4908 -65551 -4832
rect -65485 -4903 -65400 -4829
rect -65334 -4903 -65296 -4824
rect -65485 -4908 -65296 -4903
rect -65618 -4911 -65296 -4908
rect -65695 -4968 -65296 -4911
rect -65695 -4969 -65393 -4968
rect -65695 -5048 -65686 -4969
rect -65620 -5048 -65541 -4969
rect -65475 -5047 -65393 -4969
rect -65327 -5047 -65296 -4968
rect -65475 -5048 -65296 -5047
rect -65695 -8481 -65296 -5048
rect -65695 -8484 -65533 -8481
rect -65695 -8547 -65665 -8484
rect -65605 -8544 -65533 -8484
rect -65473 -8484 -65296 -8481
rect -65473 -8544 -65399 -8484
rect -65605 -8547 -65399 -8544
rect -65339 -8547 -65296 -8484
rect -65695 -10167 -65296 -8547
rect -65695 -10171 -65389 -10167
rect -65695 -10247 -65680 -10171
rect -65618 -10247 -65539 -10171
rect -65477 -10243 -65389 -10171
rect -65327 -10243 -65296 -10167
rect -65477 -10247 -65296 -10243
rect -65695 -13570 -65296 -10247
rect -65695 -13643 -65682 -13570
rect -65611 -13571 -65296 -13570
rect -65611 -13643 -65551 -13571
rect -65695 -13644 -65551 -13643
rect -65480 -13576 -65296 -13571
rect -65480 -13644 -65395 -13576
rect -65695 -13649 -65395 -13644
rect -65324 -13649 -65296 -13576
rect -65695 -13755 -65296 -13649
rect -65695 -13761 -65534 -13755
rect -65695 -13834 -65685 -13761
rect -65614 -13828 -65534 -13761
rect -65463 -13756 -65296 -13755
rect -65463 -13828 -65392 -13756
rect -65614 -13829 -65392 -13828
rect -65321 -13829 -65296 -13756
rect -65614 -13834 -65296 -13829
rect -65695 -17265 -65296 -13834
rect -65088 -1676 -64530 -1543
rect -65088 -15878 -64955 -1676
rect -56610 -2455 -56502 -2392
rect -56610 -2550 -56591 -2455
rect -56514 -2550 -56502 -2455
rect -56610 -2631 -56502 -2550
rect -56610 -2726 -56594 -2631
rect -56517 -2726 -56502 -2631
rect -56610 -2790 -56502 -2726
rect -56610 -2885 -56592 -2790
rect -56515 -2885 -56502 -2790
rect -56610 -2948 -56502 -2885
rect -56610 -3043 -56593 -2948
rect -56516 -3043 -56502 -2948
rect -56813 -3526 -56708 -3480
rect -64606 -3659 -64482 -3528
rect -64606 -3793 -64576 -3659
rect -64498 -3793 -64482 -3659
rect -64606 -3861 -64482 -3793
rect -64606 -3995 -64578 -3861
rect -64500 -3995 -64482 -3861
rect -64606 -7141 -64482 -3995
rect -56813 -3621 -56794 -3526
rect -56717 -3621 -56708 -3526
rect -56813 -3702 -56708 -3621
rect -56813 -3797 -56797 -3702
rect -56720 -3797 -56708 -3702
rect -56813 -3861 -56708 -3797
rect -56813 -3956 -56795 -3861
rect -56718 -3956 -56708 -3861
rect -56813 -4019 -56708 -3956
rect -56813 -4114 -56796 -4019
rect -56719 -4114 -56708 -4019
rect -56813 -5165 -56708 -4114
rect -56610 -5082 -56502 -3043
rect -63351 -6122 -63264 -6101
rect -63351 -6178 -63338 -6122
rect -63282 -6178 -63264 -6122
rect -63351 -6186 -63264 -6178
rect -63351 -6233 -63107 -6186
rect -63351 -6289 -63342 -6233
rect -63286 -6266 -63107 -6233
rect -63286 -6289 -63264 -6266
rect -63351 -6304 -63264 -6289
rect -64606 -7205 -64572 -7141
rect -64513 -7205 -64482 -7141
rect -64606 -7309 -64482 -7205
rect -64606 -7373 -64575 -7309
rect -64516 -7373 -64482 -7309
rect -64606 -7521 -64482 -7373
rect -64587 -12362 -64502 -7521
rect -64587 -12450 -64575 -12362
rect -64516 -12450 -64502 -12362
rect -64587 -12536 -64502 -12450
rect -64587 -12624 -64573 -12536
rect -64514 -12624 -64502 -12536
rect -64587 -12644 -64502 -12624
rect -64350 -8080 -64249 -8023
rect -64350 -8086 -64327 -8080
rect -64350 -8142 -64331 -8086
rect -64270 -8135 -64249 -8080
rect -64275 -8142 -64249 -8135
rect -64350 -8197 -64249 -8142
rect -64350 -8253 -64335 -8197
rect -64279 -8206 -64249 -8197
rect -64350 -8261 -64334 -8253
rect -64277 -8261 -64249 -8206
rect -64604 -15878 -64506 -15871
rect -65088 -15912 -64506 -15878
rect -65088 -15982 -64593 -15912
rect -64520 -15982 -64506 -15912
rect -65088 -16011 -64506 -15982
rect -65695 -17268 -65540 -17265
rect -65695 -17331 -65672 -17268
rect -65612 -17328 -65540 -17268
rect -65480 -17268 -65296 -17265
rect -65480 -17328 -65406 -17268
rect -65612 -17331 -65406 -17328
rect -65346 -17331 -65296 -17268
rect -65695 -21648 -65296 -17331
rect -65695 -21655 -65545 -21648
rect -65695 -21752 -65679 -21655
rect -65617 -21745 -65545 -21655
rect -65483 -21657 -65296 -21648
rect -65483 -21745 -65410 -21657
rect -65617 -21752 -65410 -21745
rect -65695 -21754 -65410 -21752
rect -65348 -21754 -65296 -21657
rect -65695 -21848 -65296 -21754
rect -65695 -21945 -65683 -21848
rect -65621 -21945 -65535 -21848
rect -65473 -21851 -65296 -21848
rect -65473 -21945 -65388 -21851
rect -65695 -21948 -65388 -21945
rect -65326 -21948 -65296 -21851
rect -65695 -25368 -65296 -21948
rect -64604 -16094 -64506 -16011
rect -64604 -16164 -64593 -16094
rect -64520 -16164 -64506 -16094
rect -64604 -23960 -64506 -16164
rect -64350 -16748 -64249 -8261
rect -64136 -8908 -64061 -8875
rect -64136 -8970 -64126 -8908
rect -64070 -8970 -64061 -8908
rect -63187 -8961 -63107 -6266
rect -61067 -6876 -61011 -6656
rect -61063 -7368 -61007 -7120
rect -55938 -7272 -55539 3358
rect -55938 -7273 -55668 -7272
rect -55938 -7277 -55794 -7273
rect -55938 -7329 -55922 -7277
rect -55865 -7325 -55794 -7277
rect -55737 -7324 -55668 -7273
rect -55611 -7324 -55539 -7272
rect -55737 -7325 -55539 -7324
rect -55865 -7329 -55539 -7325
rect -64136 -9048 -64061 -8970
rect -64136 -9110 -64125 -9048
rect -64069 -9110 -64061 -9048
rect -64350 -16760 -64248 -16748
rect -64350 -16763 -64337 -16760
rect -64349 -16838 -64337 -16763
rect -64259 -16838 -64248 -16760
rect -64349 -16908 -64248 -16838
rect -64349 -16984 -64336 -16908
rect -64260 -16984 -64248 -16908
rect -64349 -17004 -64248 -16984
rect -64136 -17685 -64061 -9110
rect -63247 -9041 -63107 -8961
rect -64136 -17747 -64123 -17685
rect -64070 -17747 -64061 -17685
rect -64136 -17822 -64061 -17747
rect -64136 -17884 -64123 -17822
rect -64070 -17884 -64061 -17822
rect -64136 -19366 -64061 -17884
rect -63896 -9417 -63797 -9391
rect -63896 -9471 -63872 -9417
rect -63818 -9471 -63797 -9417
rect -63896 -9547 -63797 -9471
rect -63896 -9601 -63873 -9547
rect -63819 -9601 -63797 -9547
rect -63896 -18200 -63797 -9601
rect -63247 -14882 -63167 -9041
rect -61015 -9717 -60958 -9459
rect -56610 -11381 -56502 -11345
rect -56610 -11476 -56585 -11381
rect -56508 -11476 -56502 -11381
rect -56610 -11557 -56502 -11476
rect -56610 -11652 -56588 -11557
rect -56511 -11652 -56502 -11557
rect -56610 -11716 -56502 -11652
rect -56610 -11811 -56586 -11716
rect -56509 -11811 -56502 -11716
rect -56610 -11874 -56502 -11811
rect -56610 -11969 -56587 -11874
rect -56510 -11969 -56502 -11874
rect -56813 -12421 -56708 -12369
rect -56813 -12516 -56792 -12421
rect -56715 -12516 -56708 -12421
rect -56813 -12597 -56708 -12516
rect -56813 -12692 -56795 -12597
rect -56718 -12692 -56708 -12597
rect -56813 -12756 -56708 -12692
rect -56813 -12851 -56793 -12756
rect -56716 -12851 -56708 -12756
rect -56813 -12914 -56708 -12851
rect -56813 -13009 -56794 -12914
rect -56717 -13009 -56708 -12914
rect -56813 -13971 -56708 -13009
rect -56610 -13899 -56502 -11969
rect -63330 -14888 -63167 -14882
rect -63347 -14909 -63167 -14888
rect -63347 -14965 -63334 -14909
rect -63278 -14962 -63167 -14909
rect -63278 -14965 -63260 -14962
rect -63347 -15020 -63260 -14965
rect -63347 -15076 -63338 -15020
rect -63282 -15076 -63260 -15020
rect -63347 -15091 -63260 -15076
rect -61067 -15688 -61011 -15515
rect -61064 -16134 -61008 -15900
rect -55938 -15924 -55539 -7329
rect -55938 -15925 -55624 -15924
rect -55938 -15983 -55915 -15925
rect -55862 -15983 -55771 -15925
rect -55718 -15982 -55624 -15925
rect -55571 -15982 -55539 -15924
rect -55718 -15983 -55539 -15982
rect -63669 -16879 -63582 -16858
rect -63669 -16935 -63656 -16879
rect -63600 -16935 -63582 -16879
rect -63669 -16990 -63582 -16935
rect -63669 -17046 -63660 -16990
rect -63604 -17046 -63582 -16990
rect -63669 -17061 -63582 -17046
rect -63896 -18254 -63867 -18200
rect -63815 -18254 -63797 -18200
rect -63896 -18332 -63797 -18254
rect -63896 -18386 -63868 -18332
rect -63816 -18386 -63797 -18332
rect -63896 -18901 -63797 -18386
rect -61015 -18483 -60958 -18241
rect -63905 -18983 -63795 -18901
rect -63905 -19056 -63886 -18983
rect -63807 -19056 -63795 -18983
rect -63905 -19169 -63795 -19056
rect -63905 -19242 -63889 -19169
rect -63810 -19242 -63795 -19169
rect -63905 -19270 -63795 -19242
rect -64167 -19403 -64043 -19366
rect -64167 -19471 -64144 -19403
rect -64064 -19471 -64043 -19403
rect -64167 -19589 -64043 -19471
rect -64167 -19657 -64145 -19589
rect -64065 -19657 -64043 -19589
rect -64167 -19681 -64043 -19657
rect -64376 -23960 -64281 -23959
rect -64604 -24026 -64281 -23960
rect -64604 -24084 -64355 -24026
rect -64297 -24084 -64281 -24026
rect -64604 -24207 -64281 -24084
rect -64604 -24265 -64361 -24207
rect -64303 -24265 -64281 -24207
rect -64604 -24287 -64281 -24265
rect -65695 -25371 -65540 -25368
rect -65695 -25434 -65672 -25371
rect -65612 -25431 -65540 -25371
rect -65480 -25371 -65296 -25368
rect -65480 -25431 -65406 -25371
rect -65612 -25434 -65406 -25431
rect -65346 -25434 -65296 -25371
rect -65695 -27116 -65296 -25434
rect -65695 -27118 -65522 -27116
rect -65695 -27209 -65682 -27118
rect -65616 -27207 -65522 -27118
rect -65456 -27118 -65296 -27116
rect -65456 -27207 -65380 -27118
rect -65616 -27209 -65380 -27207
rect -65314 -27209 -65296 -27118
rect -65695 -31714 -65296 -27209
rect -64376 -28449 -64281 -24287
rect -64136 -25669 -64061 -19681
rect -64137 -25692 -64058 -25669
rect -64137 -25758 -64119 -25692
rect -64066 -25758 -64058 -25692
rect -64137 -25818 -64058 -25758
rect -64137 -25884 -64127 -25818
rect -64074 -25884 -64058 -25818
rect -64137 -25903 -64058 -25884
rect -63896 -26184 -63797 -19270
rect -56642 -19450 -56534 -19434
rect -56645 -19476 -56534 -19450
rect -56645 -19571 -56627 -19476
rect -56550 -19571 -56534 -19476
rect -56645 -19652 -56534 -19571
rect -56645 -19747 -56630 -19652
rect -56553 -19747 -56534 -19652
rect -56645 -19811 -56534 -19747
rect -56645 -19906 -56628 -19811
rect -56551 -19906 -56534 -19811
rect -56645 -19969 -56534 -19906
rect -56645 -20064 -56629 -19969
rect -56552 -20064 -56534 -19969
rect -56645 -20087 -56534 -20064
rect -56845 -20487 -56740 -20452
rect -56849 -20513 -56740 -20487
rect -56849 -20608 -56831 -20513
rect -56754 -20608 -56740 -20513
rect -56849 -20689 -56740 -20608
rect -56849 -20784 -56834 -20689
rect -56757 -20784 -56740 -20689
rect -56849 -20848 -56740 -20784
rect -56849 -20943 -56832 -20848
rect -56755 -20943 -56740 -20848
rect -56849 -21006 -56740 -20943
rect -56849 -21101 -56833 -21006
rect -56756 -21101 -56740 -21006
rect -56849 -21124 -56740 -21101
rect -56845 -22011 -56740 -21124
rect -56642 -21957 -56534 -20087
rect -55938 -22527 -55539 -15983
rect -55938 -22528 -55630 -22527
rect -55938 -22631 -55917 -22528
rect -55837 -22529 -55630 -22528
rect -55837 -22631 -55769 -22529
rect -55938 -22632 -55769 -22631
rect -55689 -22630 -55630 -22529
rect -55550 -22630 -55539 -22527
rect -55689 -22632 -55539 -22630
rect -63396 -23012 -63309 -22991
rect -63396 -23068 -63383 -23012
rect -63327 -23068 -63309 -23012
rect -63396 -23123 -63309 -23068
rect -63396 -23179 -63387 -23123
rect -63331 -23179 -63309 -23123
rect -63396 -23194 -63309 -23179
rect -61099 -23802 -61043 -23599
rect -61096 -24242 -61040 -24041
rect -63739 -24952 -63652 -24931
rect -63739 -25008 -63726 -24952
rect -63670 -25008 -63652 -24952
rect -63739 -25063 -63652 -25008
rect -63739 -25119 -63730 -25063
rect -63674 -25119 -63652 -25063
rect -63739 -25127 -63652 -25119
rect -63896 -26238 -63865 -26184
rect -63812 -26238 -63797 -26184
rect -63896 -26292 -63797 -26238
rect -63896 -26347 -63860 -26292
rect -63807 -26347 -63797 -26292
rect -63896 -26367 -63797 -26347
rect -61047 -26580 -60990 -26332
rect -64376 -28505 -64357 -28449
rect -64291 -28505 -64281 -28449
rect -64376 -28608 -64281 -28505
rect -64376 -28664 -64364 -28608
rect -64298 -28664 -64281 -28608
rect -64376 -28679 -64281 -28664
rect -56423 -29010 -56216 -28892
rect -56423 -29119 -56389 -29010
rect -56253 -29119 -56216 -29010
rect -56423 -29259 -56216 -29119
rect -56423 -29368 -56397 -29259
rect -56261 -29368 -56216 -29259
rect -56707 -30528 -56561 -30443
rect -56707 -30592 -56668 -30528
rect -56587 -30592 -56561 -30528
rect -56707 -30679 -56561 -30592
rect -56707 -30743 -56677 -30679
rect -56596 -30743 -56561 -30679
rect -57036 -31228 -56888 -31172
rect -57036 -31300 -57009 -31228
rect -56906 -31300 -56888 -31228
rect -57036 -31408 -56888 -31300
rect -65695 -31717 -65522 -31714
rect -65695 -31778 -65665 -31717
rect -65606 -31775 -65522 -31717
rect -65463 -31719 -65296 -31714
rect -65463 -31775 -65397 -31719
rect -65606 -31778 -65397 -31775
rect -65695 -31780 -65397 -31778
rect -65338 -31780 -65296 -31719
rect -65695 -33205 -65296 -31780
rect -57408 -31584 -57252 -31410
rect -57408 -31663 -57382 -31584
rect -57283 -31663 -57252 -31584
rect -57408 -31751 -57252 -31663
rect -57408 -31830 -57379 -31751
rect -57280 -31830 -57252 -31751
rect -65695 -33208 -65384 -33205
rect -65695 -33210 -65532 -33208
rect -65695 -33271 -65676 -33210
rect -65617 -33269 -65532 -33210
rect -65473 -33266 -65384 -33208
rect -65325 -33266 -65296 -33205
rect -65473 -33269 -65296 -33266
rect -57756 -32415 -57585 -32325
rect -57756 -32502 -57715 -32415
rect -57596 -32502 -57585 -32415
rect -57756 -32637 -57585 -32502
rect -57756 -32724 -57733 -32637
rect -57614 -32724 -57585 -32637
rect -65617 -33271 -65296 -33269
rect -65695 -34379 -65296 -33271
rect -58103 -33392 -57936 -33269
rect -58103 -33473 -58055 -33392
rect -57975 -33473 -57936 -33392
rect -58103 -33592 -57936 -33473
rect -58103 -33673 -58069 -33592
rect -57989 -33673 -57936 -33592
rect -65695 -34382 -65545 -34379
rect -65695 -34443 -65683 -34382
rect -65624 -34440 -65545 -34382
rect -65486 -34440 -65399 -34379
rect -65340 -34440 -65296 -34379
rect -65624 -34443 -65296 -34440
rect -65695 -35605 -65296 -34443
rect -65695 -35610 -65411 -35605
rect -65695 -35613 -65544 -35610
rect -65695 -35679 -65687 -35613
rect -65624 -35676 -65544 -35613
rect -65481 -35671 -65411 -35610
rect -65348 -35671 -65296 -35605
rect -65481 -35676 -65296 -35671
rect -65624 -35679 -65296 -35676
rect -65695 -36504 -65296 -35679
rect -58450 -34399 -58287 -34259
rect -58450 -34481 -58410 -34399
rect -58313 -34481 -58287 -34399
rect -58450 -34579 -58287 -34481
rect -58450 -34661 -58415 -34579
rect -58318 -34661 -58287 -34579
rect -65695 -36521 -65284 -36504
rect -65695 -36524 -65367 -36521
rect -65695 -36529 -65516 -36524
rect -65695 -36624 -65675 -36529
rect -65598 -36619 -65516 -36529
rect -65439 -36616 -65367 -36524
rect -65290 -36616 -65284 -36521
rect -65439 -36619 -65284 -36616
rect -65598 -36624 -65284 -36619
rect -65695 -36697 -65284 -36624
rect -65695 -36700 -65370 -36697
rect -65695 -36705 -65519 -36700
rect -65695 -36800 -65678 -36705
rect -65601 -36795 -65519 -36705
rect -65442 -36792 -65370 -36700
rect -65293 -36792 -65284 -36697
rect -65442 -36795 -65284 -36792
rect -65601 -36800 -65284 -36795
rect -65695 -36856 -65284 -36800
rect -65695 -36859 -65368 -36856
rect -65695 -36864 -65517 -36859
rect -65695 -36959 -65676 -36864
rect -65599 -36954 -65517 -36864
rect -65440 -36951 -65368 -36859
rect -65291 -36951 -65284 -36856
rect -65440 -36954 -65284 -36951
rect -65599 -36959 -65284 -36954
rect -65695 -37014 -65284 -36959
rect -65695 -37017 -65369 -37014
rect -65695 -37022 -65518 -37017
rect -65695 -37117 -65677 -37022
rect -65600 -37112 -65518 -37022
rect -65441 -37109 -65369 -37017
rect -65292 -37109 -65284 -37014
rect -65441 -37112 -65284 -37109
rect -65600 -37117 -65284 -37112
rect -65695 -37129 -65284 -37117
rect -66390 -37553 -65980 -37536
rect -66390 -37556 -66063 -37553
rect -66390 -37561 -66212 -37556
rect -66390 -37656 -66371 -37561
rect -66294 -37651 -66212 -37561
rect -66135 -37648 -66063 -37556
rect -65986 -37648 -65980 -37553
rect -66135 -37651 -65980 -37648
rect -66294 -37656 -65980 -37651
rect -66390 -37729 -65980 -37656
rect -66390 -37732 -66066 -37729
rect -66390 -37737 -66215 -37732
rect -66390 -37832 -66374 -37737
rect -66297 -37827 -66215 -37737
rect -66138 -37824 -66066 -37732
rect -65989 -37824 -65980 -37729
rect -66138 -37827 -65980 -37824
rect -66297 -37832 -65980 -37827
rect -66390 -37888 -65980 -37832
rect -66390 -37891 -66064 -37888
rect -66390 -37896 -66213 -37891
rect -66390 -37991 -66372 -37896
rect -66295 -37986 -66213 -37896
rect -66136 -37983 -66064 -37891
rect -65987 -37983 -65980 -37888
rect -66136 -37986 -65980 -37983
rect -66295 -37991 -65980 -37986
rect -66390 -38046 -65980 -37991
rect -66390 -38049 -66065 -38046
rect -66390 -38054 -66214 -38049
rect -66390 -38149 -66373 -38054
rect -66296 -38144 -66214 -38054
rect -66137 -38141 -66065 -38049
rect -65988 -38141 -65980 -38046
rect -66137 -38144 -65980 -38141
rect -66296 -38149 -65980 -38144
rect -66390 -38161 -65980 -38149
rect -66381 -38193 -65982 -38161
rect -65695 -38193 -65296 -37129
rect -58450 -37359 -58287 -34661
rect -58103 -36892 -57936 -33673
rect -58103 -36963 -58065 -36892
rect -57992 -36963 -57936 -36892
rect -58103 -37049 -57936 -36963
rect -58103 -37120 -58062 -37049
rect -57989 -37120 -57936 -37049
rect -58103 -37152 -57936 -37120
rect -58449 -37406 -58287 -37359
rect -58449 -37459 -58410 -37406
rect -58341 -37459 -58287 -37406
rect -58449 -37475 -58287 -37459
rect -57756 -38058 -57585 -32724
rect -57408 -36485 -57252 -31830
rect -57408 -36552 -57382 -36485
rect -57288 -36552 -57252 -36485
rect -57408 -36623 -57252 -36552
rect -57408 -36690 -57382 -36623
rect -57288 -36690 -57252 -36623
rect -57408 -36718 -57252 -36690
rect -57036 -31480 -57019 -31408
rect -56916 -31480 -56888 -31408
rect -57756 -38116 -57731 -38058
rect -57631 -38116 -57585 -38058
rect -57756 -38186 -57585 -38116
rect -57756 -38244 -57732 -38186
rect -57632 -38244 -57585 -38186
rect -57756 -38296 -57585 -38244
rect -57756 -38354 -57731 -38296
rect -57631 -38354 -57585 -38296
rect -57756 -38383 -57585 -38354
rect -57036 -39064 -56888 -31480
rect -56707 -38680 -56561 -30743
rect -56423 -32893 -56216 -29368
rect -56423 -32969 -56365 -32893
rect -56276 -32969 -56216 -32893
rect -56423 -33084 -56216 -32969
rect -56423 -33160 -56370 -33084
rect -56281 -33160 -56216 -33084
rect -56423 -33234 -56216 -33160
rect -55938 -30701 -55539 -22632
rect -55938 -30704 -55781 -30701
rect -55938 -30767 -55913 -30704
rect -55853 -30764 -55781 -30704
rect -55721 -30704 -55539 -30701
rect -55721 -30764 -55647 -30704
rect -55853 -30767 -55647 -30764
rect -55587 -30767 -55539 -30704
rect -55938 -31137 -55539 -30767
rect -55938 -31140 -55781 -31137
rect -55938 -31203 -55913 -31140
rect -55853 -31200 -55781 -31140
rect -55721 -31140 -55539 -31137
rect -55721 -31200 -55647 -31140
rect -55853 -31203 -55647 -31200
rect -55587 -31203 -55539 -31140
rect -55938 -34642 -55539 -31203
rect -55938 -34645 -55659 -34642
rect -55938 -34727 -55924 -34645
rect -55864 -34649 -55659 -34645
rect -55864 -34727 -55798 -34649
rect -55938 -34731 -55798 -34727
rect -55738 -34724 -55659 -34649
rect -55599 -34724 -55539 -34642
rect -55738 -34731 -55539 -34724
rect -55938 -37539 -55539 -34731
rect -55294 48051 -54895 55223
rect -45764 54837 -45365 55873
rect -44941 55852 -44542 55873
rect -44941 55834 -44529 55852
rect -44941 55831 -44612 55834
rect -44941 55826 -44761 55831
rect -44941 55731 -44920 55826
rect -44843 55736 -44761 55826
rect -44684 55739 -44612 55831
rect -44535 55739 -44529 55834
rect -44684 55736 -44529 55739
rect -44843 55731 -44529 55736
rect -44941 55658 -44529 55731
rect -44941 55655 -44615 55658
rect -44941 55650 -44764 55655
rect -44941 55555 -44923 55650
rect -44846 55560 -44764 55650
rect -44687 55563 -44615 55655
rect -44538 55563 -44529 55658
rect -44687 55560 -44529 55563
rect -44846 55555 -44529 55560
rect -44941 55499 -44529 55555
rect -44941 55496 -44613 55499
rect -44941 55491 -44762 55496
rect -44941 55396 -44921 55491
rect -44844 55401 -44762 55491
rect -44685 55404 -44613 55496
rect -44536 55404 -44529 55499
rect -44685 55401 -44529 55404
rect -44844 55396 -44529 55401
rect -44941 55341 -44529 55396
rect -44941 55338 -44614 55341
rect -44941 55333 -44763 55338
rect -44941 55238 -44922 55333
rect -44845 55243 -44763 55333
rect -44686 55246 -44614 55338
rect -44537 55246 -44529 55341
rect -44686 55243 -44529 55246
rect -44845 55238 -44529 55243
rect -44941 55226 -44529 55238
rect -45764 54809 -45349 54837
rect -45764 54806 -45434 54809
rect -45764 54801 -45583 54806
rect -45764 54706 -45742 54801
rect -45665 54711 -45583 54801
rect -45506 54714 -45434 54806
rect -45357 54714 -45349 54809
rect -45506 54711 -45349 54714
rect -45665 54706 -45349 54711
rect -45764 54633 -45349 54706
rect -45764 54630 -45437 54633
rect -45764 54625 -45586 54630
rect -45764 54530 -45745 54625
rect -45668 54535 -45586 54625
rect -45509 54538 -45437 54630
rect -45360 54538 -45349 54633
rect -45509 54535 -45349 54538
rect -45668 54530 -45349 54535
rect -45764 54474 -45349 54530
rect -45764 54471 -45435 54474
rect -45764 54466 -45584 54471
rect -45764 54371 -45743 54466
rect -45666 54376 -45584 54466
rect -45507 54379 -45435 54471
rect -45358 54379 -45349 54474
rect -45507 54376 -45349 54379
rect -45666 54371 -45349 54376
rect -45764 54316 -45349 54371
rect -45764 54313 -45436 54316
rect -45764 54308 -45585 54313
rect -45764 54213 -45744 54308
rect -45667 54218 -45585 54308
rect -45508 54221 -45436 54313
rect -45359 54221 -45349 54316
rect -45508 54218 -45349 54221
rect -45667 54213 -45349 54218
rect -45764 54199 -45349 54213
rect -46413 53602 -46305 53633
rect -46413 53507 -46395 53602
rect -46318 53507 -46305 53602
rect -46413 53426 -46305 53507
rect -46413 53331 -46398 53426
rect -46321 53331 -46305 53426
rect -46413 53267 -46305 53331
rect -46413 53172 -46396 53267
rect -46319 53172 -46305 53267
rect -46413 53109 -46305 53172
rect -46413 53014 -46397 53109
rect -46320 53014 -46305 53109
rect -46616 52572 -46511 52586
rect -46616 52477 -46599 52572
rect -46522 52477 -46511 52572
rect -53949 52415 -53842 52442
rect -53949 52343 -53932 52415
rect -53860 52343 -53842 52415
rect -53949 52194 -53842 52343
rect -53949 52120 -53933 52194
rect -53859 52120 -53842 52194
rect -46616 52369 -46511 52477
rect -46616 52274 -46600 52369
rect -46523 52274 -46511 52369
rect -53949 52105 -53842 52120
rect -53685 52165 -53551 52183
rect -55294 48048 -55127 48051
rect -55294 47985 -55259 48048
rect -55199 47988 -55127 48048
rect -55067 48048 -54895 48051
rect -55067 47988 -54993 48048
rect -55199 47985 -54993 47988
rect -54933 47985 -54895 48048
rect -55294 47672 -54895 47985
rect -55294 47669 -55139 47672
rect -55294 47606 -55271 47669
rect -55211 47609 -55139 47669
rect -55079 47669 -54895 47672
rect -55079 47609 -55005 47669
rect -55211 47606 -55005 47609
rect -54945 47606 -54895 47669
rect -55294 43046 -54895 47606
rect -55294 43045 -54984 43046
rect -55294 43044 -55133 43045
rect -55294 42963 -55281 43044
rect -55217 42964 -55133 43044
rect -55069 42965 -54984 43045
rect -54920 42965 -54895 43046
rect -55069 42964 -54895 42965
rect -55217 42963 -54895 42964
rect -55294 39724 -54895 42963
rect -55294 39723 -54996 39724
rect -55294 39721 -55137 39723
rect -55294 39650 -55273 39721
rect -55215 39652 -55137 39721
rect -55079 39653 -54996 39723
rect -54938 39653 -54895 39724
rect -55079 39652 -54895 39653
rect -55215 39650 -54895 39652
rect -55294 39346 -54895 39650
rect -55294 39345 -55003 39346
rect -55294 39343 -55144 39345
rect -55294 39272 -55280 39343
rect -55222 39274 -55144 39343
rect -55086 39275 -55003 39345
rect -54945 39275 -54895 39346
rect -55086 39274 -54895 39275
rect -55222 39272 -54895 39274
rect -55294 34598 -54895 39272
rect -54509 48965 -54387 49041
rect -54509 48888 -54492 48965
rect -54412 48888 -54387 48965
rect -54509 48777 -54387 48888
rect -54509 48700 -54492 48777
rect -54412 48700 -54387 48777
rect -54509 37025 -54387 48700
rect -53936 46884 -53855 52105
rect -53685 52067 -53671 52165
rect -53573 52067 -53551 52165
rect -53685 51987 -53551 52067
rect -53685 51887 -53672 51987
rect -53572 51887 -53551 51987
rect -53685 51877 -53551 51887
rect -46616 52167 -46511 52274
rect -46616 52072 -46601 52167
rect -46524 52072 -46511 52167
rect -53672 47298 -53572 51877
rect -46616 51694 -46511 52072
rect -46616 51638 -46588 51694
rect -46533 51638 -46511 51694
rect -53272 50091 -53149 50105
rect -53272 50012 -53252 50091
rect -53161 50012 -53149 50091
rect -53272 49939 -53149 50012
rect -50867 49999 -50272 50055
rect -53272 49860 -53256 49939
rect -53165 49860 -53149 49939
rect -53272 49848 -53149 49860
rect -50867 49032 -50811 49051
rect -50867 48978 -50866 49032
rect -50812 48978 -50811 49032
rect -50867 48835 -50811 48978
rect -46616 48169 -46511 51638
rect -46413 51555 -46305 53014
rect -46413 51499 -46382 51555
rect -46327 51499 -46305 51555
rect -46413 50813 -46305 51499
rect -45764 50308 -45365 54199
rect -45764 50305 -45613 50308
rect -45764 50242 -45745 50305
rect -45685 50245 -45613 50305
rect -45553 50305 -45365 50308
rect -45553 50245 -45479 50305
rect -45685 50242 -45479 50245
rect -45419 50242 -45365 50305
rect -53672 47198 -53166 47298
rect -53953 46870 -53843 46884
rect -53953 46793 -53933 46870
rect -53856 46793 -53843 46870
rect -53953 46731 -53843 46793
rect -53953 46650 -53936 46731
rect -53855 46650 -53843 46731
rect -53953 46634 -53843 46650
rect -50818 46530 -50761 46638
rect -50764 46471 -50761 46530
rect -50818 46462 -50761 46471
rect -46405 45228 -46297 45269
rect -46405 45133 -46389 45228
rect -46312 45133 -46297 45228
rect -46405 45052 -46297 45133
rect -46405 44957 -46392 45052
rect -46315 44957 -46297 45052
rect -46405 44893 -46297 44957
rect -46405 44798 -46390 44893
rect -46313 44798 -46297 44893
rect -46405 44735 -46297 44798
rect -46405 44640 -46391 44735
rect -46314 44640 -46297 44735
rect -46608 44191 -46503 44230
rect -46608 44096 -46592 44191
rect -46515 44096 -46503 44191
rect -46608 44015 -46503 44096
rect -46608 43920 -46595 44015
rect -46518 43920 -46503 44015
rect -46608 43856 -46503 43920
rect -46608 43761 -46593 43856
rect -46516 43761 -46503 43856
rect -46608 43698 -46503 43761
rect -46608 43603 -46594 43698
rect -46517 43603 -46503 43698
rect -46608 43362 -46503 43603
rect -46608 43306 -46580 43362
rect -46525 43306 -46503 43362
rect -46608 42738 -46503 43306
rect -46405 43223 -46297 44640
rect -46405 43167 -46374 43223
rect -46319 43167 -46297 43223
rect -46405 42783 -46297 43167
rect -45764 42139 -45365 50242
rect -45764 42131 -45591 42139
rect -45764 42075 -45731 42131
rect -45679 42083 -45591 42131
rect -45539 42130 -45365 42139
rect -45539 42083 -45462 42130
rect -45679 42075 -45462 42083
rect -45764 42074 -45462 42075
rect -45410 42074 -45365 42130
rect -53195 41757 -53072 41771
rect -53195 41678 -53175 41757
rect -53084 41678 -53072 41757
rect -53195 41605 -53072 41678
rect -50859 41667 -50264 41723
rect -53195 41526 -53179 41605
rect -53088 41526 -53072 41605
rect -53195 41514 -53072 41526
rect -50862 41102 -50806 41439
rect -54190 40754 -54017 40769
rect -54190 40702 -54168 40754
rect -54040 40702 -54017 40754
rect -54190 40630 -54017 40702
rect -54190 40578 -54168 40630
rect -54040 40578 -54017 40630
rect -54190 40487 -54017 40578
rect -54190 40435 -54167 40487
rect -54039 40435 -54017 40487
rect -50859 40700 -50803 40719
rect -50859 40646 -50858 40700
rect -50804 40646 -50803 40700
rect -50859 40467 -50803 40646
rect -54509 37021 -54384 37025
rect -54508 36947 -54384 37021
rect -54508 36856 -54477 36947
rect -54406 36856 -54384 36947
rect -54508 36755 -54384 36856
rect -54508 36664 -54487 36755
rect -54416 36664 -54384 36755
rect -54508 36652 -54384 36664
rect -55294 34595 -55156 34598
rect -55294 34520 -55284 34595
rect -55225 34523 -55156 34595
rect -55097 34597 -54895 34598
rect -55097 34523 -55027 34597
rect -55225 34522 -55027 34523
rect -54968 34522 -54895 34597
rect -55225 34520 -54895 34522
rect -55294 30914 -54895 34520
rect -55294 30910 -54990 30914
rect -55294 30907 -55127 30910
rect -55294 30826 -55272 30907
rect -55204 30829 -55127 30907
rect -55059 30833 -54990 30910
rect -54922 30833 -54895 30914
rect -55059 30829 -54895 30833
rect -55204 30826 -54895 30829
rect -55294 26230 -54895 30826
rect -55294 26129 -55284 26230
rect -55214 26229 -54895 26230
rect -55214 26227 -55004 26229
rect -55214 26129 -55150 26227
rect -55294 26126 -55150 26129
rect -55080 26128 -55004 26227
rect -54934 26128 -54895 26229
rect -55080 26126 -54895 26128
rect -55294 21195 -54895 26126
rect -55294 21193 -54999 21195
rect -55294 21192 -55145 21193
rect -55294 21137 -55278 21192
rect -55223 21138 -55145 21192
rect -55090 21140 -54999 21193
rect -54944 21140 -54895 21195
rect -55090 21138 -54895 21140
rect -55223 21137 -54895 21138
rect -55294 17035 -54895 21137
rect -55294 17034 -55138 17035
rect -55294 16945 -55282 17034
rect -55223 16946 -55138 17034
rect -55079 17034 -54895 17035
rect -55079 16946 -54982 17034
rect -55223 16945 -54982 16946
rect -54923 16945 -54895 17034
rect -55294 13631 -54895 16945
rect -55294 13540 -55278 13631
rect -55202 13629 -54895 13631
rect -55202 13540 -55146 13629
rect -55294 13538 -55146 13540
rect -55070 13538 -55006 13629
rect -54930 13538 -54895 13629
rect -55294 4728 -54895 13538
rect -55294 4720 -54966 4728
rect -55294 4715 -55124 4720
rect -55294 4641 -55285 4715
rect -55229 4646 -55124 4715
rect -55068 4654 -54966 4720
rect -54910 4654 -54895 4728
rect -55068 4646 -54895 4654
rect -55229 4641 -54895 4646
rect -55294 693 -54895 4641
rect -54190 32327 -54017 40435
rect -53825 38413 -53722 38421
rect -53825 38344 -53804 38413
rect -53741 38344 -53722 38413
rect -53825 38253 -53722 38344
rect -53825 38184 -53805 38253
rect -53742 38184 -53722 38253
rect -50810 38198 -50753 38379
rect -53825 36507 -53722 38184
rect -50756 38139 -50753 38198
rect -50810 38131 -50753 38139
rect -53236 37915 -53178 38011
rect -53825 36436 -53800 36507
rect -53821 36434 -53800 36436
rect -53729 36436 -53722 36507
rect -53729 36434 -53726 36436
rect -53821 36335 -53726 36434
rect -53821 36262 -53806 36335
rect -53735 36262 -53726 36335
rect -53821 36240 -53726 36262
rect -53258 36287 -53155 37915
rect -53258 36215 -53242 36287
rect -53165 36215 -53155 36287
rect -53258 36119 -53155 36215
rect -53258 36047 -53246 36119
rect -53169 36047 -53155 36119
rect -53258 36032 -53155 36047
rect -46416 37020 -46308 37054
rect -46416 36925 -46396 37020
rect -46319 36925 -46308 37020
rect -46416 36844 -46308 36925
rect -46416 36749 -46399 36844
rect -46322 36749 -46308 36844
rect -46416 36685 -46308 36749
rect -46416 36590 -46397 36685
rect -46320 36590 -46308 36685
rect -46416 36527 -46308 36590
rect -46416 36432 -46398 36527
rect -46321 36432 -46308 36527
rect -46619 35763 -46514 35795
rect -46619 35668 -46601 35763
rect -46524 35668 -46514 35763
rect -46619 35587 -46514 35668
rect -46619 35492 -46604 35587
rect -46527 35492 -46514 35587
rect -46619 35428 -46514 35492
rect -46619 35333 -46602 35428
rect -46525 35333 -46514 35428
rect -46619 35270 -46514 35333
rect -46619 35175 -46603 35270
rect -46526 35175 -46514 35270
rect -46619 34237 -46514 35175
rect -46416 34334 -46308 36432
rect -45764 33630 -45365 42074
rect -45764 33629 -45469 33630
rect -45764 33548 -45755 33629
rect -45685 33628 -45469 33629
rect -45685 33548 -45621 33628
rect -45764 33547 -45621 33548
rect -45551 33549 -45469 33628
rect -45399 33549 -45365 33630
rect -45551 33547 -45365 33549
rect -53204 33293 -53081 33307
rect -53204 33214 -53184 33293
rect -53093 33214 -53081 33293
rect -53204 33141 -53081 33214
rect -53204 33062 -53188 33141
rect -53097 33062 -53081 33141
rect -53204 33050 -53081 33062
rect -50873 32855 -50817 32970
rect -54190 32270 -54170 32327
rect -54034 32270 -54017 32327
rect -54190 32181 -54017 32270
rect -54190 32124 -54169 32181
rect -54033 32124 -54017 32181
rect -54190 32060 -54017 32124
rect -54190 32003 -54169 32060
rect -54033 32003 -54017 32060
rect -50870 32019 -50814 32244
rect -54190 18875 -54017 32003
rect -53503 31350 -53380 31364
rect -53503 31271 -53483 31350
rect -53392 31271 -53380 31350
rect -53503 31198 -53380 31271
rect -53503 31119 -53487 31198
rect -53396 31119 -53380 31198
rect -53503 31107 -53380 31119
rect -54190 18808 -54148 18875
rect -54063 18808 -54017 18875
rect -54190 18744 -54017 18808
rect -54190 18635 -54150 18744
rect -54048 18635 -54017 18744
rect -54190 18505 -54017 18635
rect -54190 18396 -54158 18505
rect -54056 18396 -54017 18505
rect -54190 14968 -54017 18396
rect -54190 14901 -54097 14968
rect -54033 14901 -54017 14968
rect -54190 14795 -54017 14901
rect -54190 14728 -54100 14795
rect -54036 14728 -54017 14795
rect -54190 2246 -54017 14728
rect -53901 29973 -53788 29991
rect -53901 29898 -53884 29973
rect -53809 29898 -53788 29973
rect -53901 29795 -53788 29898
rect -53901 29718 -53884 29795
rect -53807 29718 -53788 29795
rect -53901 26515 -53788 29718
rect -50821 29678 -50764 29921
rect -53901 26443 -53886 26515
rect -53814 26443 -53788 26515
rect -53901 26379 -53788 26443
rect -53901 26307 -53886 26379
rect -53814 26307 -53788 26379
rect -53901 20990 -53788 26307
rect -53901 20935 -53876 20990
rect -53821 20935 -53788 20990
rect -53901 20857 -53788 20935
rect -53901 20802 -53875 20857
rect -53820 20802 -53788 20857
rect -53901 12850 -53788 20802
rect -53699 29370 -53165 29491
rect -53699 25797 -53578 29370
rect -53699 25781 -53379 25797
rect -53699 25775 -53446 25781
rect -53699 25717 -53594 25775
rect -53536 25723 -53446 25775
rect -53388 25723 -53379 25781
rect -53536 25717 -53379 25723
rect -53699 25703 -53379 25717
rect -53699 20724 -53578 25703
rect -45764 25206 -45365 33547
rect -45764 25205 -45608 25206
rect -45764 25127 -45746 25205
rect -45674 25128 -45608 25205
rect -45536 25128 -45474 25206
rect -45402 25128 -45365 25206
rect -45674 25127 -45365 25128
rect -52270 23965 -52214 24111
rect -52884 22859 -52828 22960
rect -51820 21679 -51764 21869
rect -53370 21562 -53180 21571
rect -53370 21507 -53361 21562
rect -53306 21507 -53250 21562
rect -53195 21507 -53180 21562
rect -53370 21498 -53180 21507
rect -53699 20669 -53675 20724
rect -53620 20669 -53578 20724
rect -53699 20591 -53578 20669
rect -53699 20536 -53674 20591
rect -53619 20536 -53578 20591
rect -53699 13223 -53578 20536
rect -53258 20549 -53187 21498
rect -53258 20538 -52985 20549
rect -53258 20481 -53173 20538
rect -53113 20481 -53058 20538
rect -52998 20481 -52985 20538
rect -53258 20463 -52985 20481
rect -53192 20461 -52985 20463
rect -52534 20347 -52463 21010
rect -52602 20336 -52395 20347
rect -52602 20279 -52583 20336
rect -52523 20279 -52468 20336
rect -52408 20279 -52395 20336
rect -52602 20259 -52395 20279
rect -46424 19409 -46316 19437
rect -46424 19314 -46406 19409
rect -46329 19314 -46316 19409
rect -46424 19233 -46316 19314
rect -46424 19138 -46409 19233
rect -46332 19138 -46316 19233
rect -46424 19074 -46316 19138
rect -46424 18979 -46407 19074
rect -46330 18979 -46316 19074
rect -46424 18916 -46316 18979
rect -46424 18821 -46408 18916
rect -46331 18821 -46316 18916
rect -46627 18322 -46522 18360
rect -46627 18227 -46605 18322
rect -46528 18227 -46522 18322
rect -46627 18146 -46522 18227
rect -46627 18051 -46608 18146
rect -46531 18051 -46522 18146
rect -46627 17987 -46522 18051
rect -46627 17892 -46606 17987
rect -46529 17892 -46522 17987
rect -46627 17829 -46522 17892
rect -46627 17734 -46607 17829
rect -46530 17734 -46522 17829
rect -46627 17018 -46522 17734
rect -46424 17046 -46316 18821
rect -45764 16037 -45365 25127
rect -53179 15933 -53092 15954
rect -53179 15877 -53166 15933
rect -53110 15894 -53092 15933
rect -45764 15951 -45752 16037
rect -45682 16036 -45365 16037
rect -45682 15951 -45608 16036
rect -45764 15950 -45608 15951
rect -45538 15950 -45479 16036
rect -45409 15950 -45365 16036
rect -53110 15877 -52909 15894
rect -53179 15822 -52909 15877
rect -53179 15766 -53170 15822
rect -53114 15798 -52909 15822
rect -53114 15766 -53092 15798
rect -53179 15751 -53092 15766
rect -53474 14035 -53387 14056
rect -53474 13979 -53461 14035
rect -53405 13979 -53387 14035
rect -53474 13924 -53387 13979
rect -53474 13868 -53465 13924
rect -53409 13868 -53387 13924
rect -53474 13853 -53387 13868
rect -53699 13102 -53179 13223
rect -53005 13165 -52909 15798
rect -50881 15234 -50825 15429
rect -50878 14751 -50822 14986
rect -53901 12773 -53885 12850
rect -53808 12773 -53788 12850
rect -53901 12687 -53788 12773
rect -53901 12612 -53885 12687
rect -53810 12612 -53788 12687
rect -53901 12594 -53788 12612
rect -53074 13069 -52909 13165
rect -53255 11862 -53197 12341
rect -53266 11852 -53180 11862
rect -53266 11794 -53255 11852
rect -53197 11794 -53180 11852
rect -53266 11716 -53180 11794
rect -53266 11660 -53254 11716
rect -53198 11660 -53180 11716
rect -53266 11651 -53180 11660
rect -53074 3320 -52978 13069
rect -50829 12384 -50772 12638
rect -46447 7422 -46339 7430
rect -46447 7396 -46336 7422
rect -46447 7301 -46419 7396
rect -46342 7301 -46336 7396
rect -46447 7220 -46336 7301
rect -46447 7125 -46422 7220
rect -46345 7125 -46336 7220
rect -46447 7061 -46336 7125
rect -46447 6966 -46420 7061
rect -46343 6966 -46336 7061
rect -46447 6903 -46336 6966
rect -46447 6808 -46421 6903
rect -46344 6808 -46336 6903
rect -46447 6785 -46336 6808
rect -46650 6187 -46545 6198
rect -46650 6161 -46540 6187
rect -46650 6066 -46623 6161
rect -46546 6066 -46540 6161
rect -46650 5985 -46540 6066
rect -46650 5890 -46626 5985
rect -46549 5890 -46540 5985
rect -46650 5826 -46540 5890
rect -46650 5731 -46624 5826
rect -46547 5731 -46540 5826
rect -46650 5668 -46540 5731
rect -46650 5573 -46625 5668
rect -46548 5573 -46540 5668
rect -46650 5550 -46540 5573
rect -46650 4104 -46545 5550
rect -46447 4073 -46339 6785
rect -53074 3224 -52880 3320
rect -53207 3049 -53120 3070
rect -53207 2993 -53194 3049
rect -53138 2993 -53120 3049
rect -53207 2938 -53120 2993
rect -53207 2882 -53198 2938
rect -53142 2882 -53120 2938
rect -53207 2867 -53120 2882
rect -55294 690 -54997 693
rect -55294 685 -55150 690
rect -55294 608 -55280 685
rect -55215 613 -55150 685
rect -55085 616 -54997 690
rect -54932 616 -54895 693
rect -55085 613 -54895 616
rect -55215 608 -54895 613
rect -55294 -693 -54895 608
rect -55294 -770 -55282 -693
rect -55225 -770 -55151 -693
rect -55094 -694 -54895 -693
rect -55094 -770 -55022 -694
rect -55294 -771 -55022 -770
rect -54965 -771 -54895 -694
rect -55294 -4777 -54895 -771
rect -54371 2167 -54017 2246
rect -54371 2098 -54104 2167
rect -54036 2098 -54017 2167
rect -54371 2026 -54017 2098
rect -54371 1957 -54106 2026
rect -54038 1957 -54017 2026
rect -54371 1953 -54017 1957
rect -54371 -3065 -54203 1953
rect -54117 1941 -54017 1953
rect -54114 1938 -54017 1941
rect -53640 1094 -53553 1115
rect -52976 1105 -52880 3224
rect -45764 3214 -45365 15950
rect -45764 3212 -45473 3214
rect -45764 3138 -45753 3212
rect -45681 3138 -45618 3212
rect -45546 3140 -45473 3212
rect -45401 3140 -45365 3214
rect -45546 3138 -45365 3140
rect -50904 2281 -50848 2457
rect -50901 1814 -50845 2059
rect -53640 1038 -53627 1094
rect -53571 1038 -53553 1094
rect -53640 983 -53553 1038
rect -53640 927 -53631 983
rect -53575 927 -53553 983
rect -53035 1073 -52794 1105
rect -53035 1062 -52878 1073
rect -53035 984 -53009 1062
rect -52949 995 -52878 1062
rect -52818 995 -52794 1073
rect -52949 984 -52794 995
rect -53035 970 -52794 984
rect -52976 967 -52880 970
rect -53640 912 -53553 927
rect -54009 -233 -53698 -226
rect -54023 -239 -53698 -233
rect -54023 -241 -53826 -239
rect -54023 -316 -53994 -241
rect -53919 -316 -53826 -241
rect -53749 -316 -53698 -239
rect -54023 -338 -53698 -316
rect -54023 -1146 -53918 -338
rect -50852 -542 -50795 -287
rect -54023 -1205 -54003 -1146
rect -53937 -1205 -53918 -1146
rect -54023 -1262 -53918 -1205
rect -54023 -1321 -54005 -1262
rect -53939 -1321 -53918 -1262
rect -54371 -3199 -54202 -3065
rect -54371 -3259 -54203 -3199
rect -54371 -3396 -54337 -3259
rect -54234 -3396 -54203 -3259
rect -54371 -3511 -54203 -3396
rect -54371 -3648 -54346 -3511
rect -54243 -3648 -54203 -3511
rect -54371 -3677 -54203 -3648
rect -55294 -4781 -54975 -4777
rect -55294 -4852 -55281 -4781
rect -55224 -4783 -54975 -4781
rect -55224 -4852 -55137 -4783
rect -55294 -4854 -55137 -4852
rect -55080 -4848 -54975 -4783
rect -54918 -4848 -54895 -4777
rect -55080 -4854 -54895 -4848
rect -55294 -4940 -54895 -4854
rect -55294 -4944 -54971 -4940
rect -55294 -5015 -55283 -4944
rect -55226 -4945 -54971 -4944
rect -55226 -5015 -55139 -4945
rect -55294 -5016 -55139 -5015
rect -55082 -5011 -54971 -4945
rect -54914 -5011 -54895 -4940
rect -55082 -5016 -54895 -5011
rect -55294 -8427 -54895 -5016
rect -55294 -8429 -54987 -8427
rect -55294 -8495 -55285 -8429
rect -55233 -8432 -54987 -8429
rect -55233 -8495 -55149 -8432
rect -55294 -8498 -55149 -8495
rect -55097 -8493 -54987 -8432
rect -54935 -8493 -54895 -8427
rect -55097 -8498 -54895 -8493
rect -55294 -9703 -54895 -8498
rect -55294 -9767 -55274 -9703
rect -55203 -9704 -54895 -9703
rect -55203 -9767 -55134 -9704
rect -55294 -9768 -55134 -9767
rect -55063 -9708 -54895 -9704
rect -55063 -9768 -54991 -9708
rect -55294 -9772 -54991 -9768
rect -54920 -9772 -54895 -9708
rect -55294 -13497 -54895 -9772
rect -54023 -4404 -53918 -1321
rect -54023 -4476 -54002 -4404
rect -53930 -4476 -53918 -4404
rect -54023 -4553 -53918 -4476
rect -54023 -4627 -54003 -4553
rect -53929 -4627 -53918 -4553
rect -54305 -12584 -54219 -12556
rect -54305 -12674 -54294 -12584
rect -54231 -12674 -54219 -12584
rect -54305 -12779 -54219 -12674
rect -54305 -12869 -54295 -12779
rect -54232 -12869 -54219 -12779
rect -54305 -12876 -54219 -12869
rect -55294 -13499 -55000 -13497
rect -55294 -13500 -55137 -13499
rect -55294 -13568 -55276 -13500
rect -55214 -13567 -55137 -13500
rect -55075 -13565 -55000 -13499
rect -54938 -13565 -54895 -13497
rect -55075 -13567 -54895 -13565
rect -55214 -13568 -54895 -13567
rect -55294 -17196 -54895 -13568
rect -55294 -17198 -54986 -17196
rect -55294 -17266 -55285 -17198
rect -55233 -17266 -55152 -17198
rect -55100 -17264 -54986 -17198
rect -54934 -17264 -54895 -17196
rect -55100 -17266 -54895 -17264
rect -55294 -18836 -54895 -17266
rect -55294 -18845 -54983 -18836
rect -55294 -18848 -55139 -18845
rect -55294 -18934 -55280 -18848
rect -55214 -18931 -55139 -18848
rect -55073 -18922 -54983 -18845
rect -54917 -18922 -54895 -18836
rect -55073 -18931 -54895 -18922
rect -55214 -18934 -54895 -18931
rect -55294 -21673 -54895 -18934
rect -55294 -21677 -55004 -21673
rect -55294 -21749 -55288 -21677
rect -55226 -21749 -55155 -21677
rect -55093 -21745 -55004 -21677
rect -54942 -21745 -54895 -21673
rect -55093 -21749 -54895 -21745
rect -55294 -25280 -54895 -21749
rect -54306 -23962 -54218 -12876
rect -54023 -13738 -53918 -4627
rect -53761 -830 -53199 -725
rect -53761 -1330 -53656 -830
rect -53761 -1390 -53743 -1330
rect -53678 -1390 -53656 -1330
rect -53761 -1446 -53656 -1390
rect -53761 -1506 -53742 -1446
rect -53677 -1506 -53656 -1446
rect -53761 -5104 -53656 -1506
rect -53775 -5127 -53465 -5104
rect -53775 -5128 -53571 -5127
rect -53775 -5186 -53741 -5128
rect -53685 -5185 -53571 -5128
rect -53515 -5185 -53465 -5127
rect -53685 -5186 -53465 -5185
rect -53775 -5215 -53465 -5186
rect -53761 -13171 -53656 -5215
rect -45764 -5761 -45365 3138
rect -45764 -5763 -45478 -5761
rect -45764 -5764 -45614 -5763
rect -45764 -5826 -45752 -5764
rect -45687 -5825 -45614 -5764
rect -45549 -5823 -45478 -5763
rect -45413 -5823 -45365 -5761
rect -45549 -5825 -45365 -5823
rect -45687 -5826 -45365 -5825
rect -52302 -6929 -52246 -6790
rect -52916 -8164 -52860 -8030
rect -51852 -9226 -51796 -9036
rect -53483 -9344 -53237 -9336
rect -53483 -9399 -53466 -9344
rect -53411 -9399 -53323 -9344
rect -53268 -9399 -53237 -9344
rect -53483 -9409 -53237 -9399
rect -53308 -10450 -53237 -9409
rect -53340 -10467 -53057 -10450
rect -53340 -10543 -53325 -10467
rect -53248 -10470 -53057 -10467
rect -53248 -10539 -53170 -10470
rect -53103 -10539 -53057 -10470
rect -53248 -10543 -53057 -10539
rect -53340 -10555 -53057 -10543
rect -52566 -10843 -52495 -9833
rect -52668 -10860 -52385 -10843
rect -52668 -10936 -52653 -10860
rect -52576 -10863 -52385 -10860
rect -52576 -10932 -52498 -10863
rect -52431 -10932 -52385 -10863
rect -52576 -10936 -52385 -10932
rect -52668 -10948 -52385 -10936
rect -53775 -13188 -53370 -13171
rect -53775 -13293 -53761 -13188
rect -53656 -13291 -53489 -13188
rect -53386 -13291 -53370 -13188
rect -53656 -13293 -53370 -13291
rect -53775 -13308 -53370 -13293
rect -54023 -13795 -53999 -13738
rect -53942 -13795 -53918 -13738
rect -54023 -13860 -53918 -13795
rect -54023 -13915 -53999 -13860
rect -53944 -13915 -53918 -13860
rect -54023 -13935 -53918 -13915
rect -51805 -14220 -51749 -14033
rect -45764 -14674 -45365 -5826
rect -45764 -14675 -45492 -14674
rect -45764 -14678 -45627 -14675
rect -45764 -14744 -45753 -14678
rect -45681 -14741 -45627 -14678
rect -45555 -14740 -45492 -14675
rect -45420 -14740 -45365 -14674
rect -45555 -14741 -45365 -14740
rect -45681 -14744 -45365 -14741
rect -52869 -15274 -52813 -15144
rect -52255 -16481 -52199 -16318
rect -53767 -18065 -53342 -18043
rect -53767 -18140 -53634 -18065
rect -53560 -18070 -53342 -18065
rect -53560 -18134 -53451 -18070
rect -53377 -18134 -53290 -18070
rect -53560 -18140 -53290 -18134
rect -53767 -18155 -53342 -18140
rect -54014 -18783 -53902 -18768
rect -54014 -18855 -53991 -18783
rect -53919 -18855 -53902 -18783
rect -54014 -18946 -53902 -18855
rect -54014 -19020 -53992 -18946
rect -53918 -19020 -53902 -18946
rect -54306 -24001 -54157 -23962
rect -54306 -24059 -54223 -24001
rect -54171 -24059 -54157 -24001
rect -54306 -24171 -54157 -24059
rect -54306 -24229 -54228 -24171
rect -54176 -24229 -54157 -24171
rect -54306 -24502 -54157 -24229
rect -55294 -25383 -55272 -25280
rect -55192 -25281 -54983 -25280
rect -55192 -25383 -55120 -25281
rect -55294 -25384 -55120 -25383
rect -55040 -25383 -54983 -25281
rect -54903 -25383 -54895 -25280
rect -55040 -25384 -54895 -25383
rect -55294 -27046 -54895 -25384
rect -55294 -27058 -54971 -27046
rect -55294 -27130 -55286 -27058
rect -55224 -27130 -55145 -27058
rect -55083 -27118 -54971 -27058
rect -54909 -27118 -54895 -27046
rect -55083 -27130 -54895 -27118
rect -55294 -29739 -54895 -27130
rect -54240 -28060 -54157 -24502
rect -54014 -26041 -53902 -19020
rect -53767 -19238 -53655 -18155
rect -53767 -19331 -53748 -19238
rect -53671 -19331 -53655 -19238
rect -53767 -19387 -53655 -19331
rect -53767 -19480 -53751 -19387
rect -53674 -19480 -53655 -19387
rect -53767 -25680 -53655 -19480
rect -46453 -19471 -46345 -19421
rect -46453 -19566 -46430 -19471
rect -46353 -19566 -46345 -19471
rect -46453 -19647 -46345 -19566
rect -46453 -19742 -46433 -19647
rect -46356 -19742 -46345 -19647
rect -46453 -19806 -46345 -19742
rect -46453 -19901 -46431 -19806
rect -46354 -19901 -46345 -19806
rect -46453 -19964 -46345 -19901
rect -46453 -20059 -46432 -19964
rect -46355 -20059 -46345 -19964
rect -46656 -20509 -46551 -20459
rect -46656 -20604 -46636 -20509
rect -46559 -20604 -46551 -20509
rect -46656 -20685 -46551 -20604
rect -46656 -20780 -46639 -20685
rect -46562 -20780 -46551 -20685
rect -46656 -20844 -46551 -20780
rect -46656 -20939 -46637 -20844
rect -46560 -20939 -46551 -20844
rect -46656 -21002 -46551 -20939
rect -46656 -21097 -46638 -21002
rect -46561 -21097 -46551 -21002
rect -46656 -21906 -46551 -21097
rect -46453 -21963 -46345 -20059
rect -45764 -22605 -45365 -14744
rect -45764 -22608 -45464 -22605
rect -45764 -22615 -45624 -22608
rect -45764 -22671 -45752 -22615
rect -45700 -22664 -45624 -22615
rect -45572 -22661 -45464 -22608
rect -45412 -22661 -45365 -22605
rect -45572 -22664 -45365 -22661
rect -45700 -22671 -45365 -22664
rect -53204 -22980 -53117 -22959
rect -53204 -23036 -53191 -22980
rect -53135 -23036 -53117 -22980
rect -53204 -23091 -53117 -23036
rect -53204 -23147 -53195 -23091
rect -53139 -23147 -53117 -23091
rect -53204 -23162 -53117 -23147
rect -50910 -23738 -50854 -23565
rect -50907 -24176 -50851 -24006
rect -53554 -24909 -53409 -24882
rect -53554 -24971 -53526 -24909
rect -53467 -24971 -53409 -24909
rect -53554 -25047 -53409 -24971
rect -53554 -25109 -53543 -25047
rect -53484 -25109 -53409 -25047
rect -53554 -25124 -53409 -25109
rect -53767 -25792 -53210 -25680
rect -54014 -26118 -53999 -26041
rect -53922 -26118 -53902 -26041
rect -54014 -26227 -53902 -26118
rect -54014 -26302 -53999 -26227
rect -53924 -26302 -53902 -26227
rect -54014 -26309 -53902 -26302
rect -54014 -26325 -53903 -26309
rect -50858 -26515 -50801 -26271
rect -54240 -28121 -54225 -28060
rect -54170 -28121 -54157 -28060
rect -54240 -28224 -54157 -28121
rect -54240 -28285 -54229 -28224
rect -54174 -28285 -54157 -28224
rect -54240 -28297 -54157 -28285
rect -46420 -27513 -46312 -27459
rect -46420 -27608 -46396 -27513
rect -46319 -27608 -46312 -27513
rect -46420 -27689 -46312 -27608
rect -46420 -27784 -46399 -27689
rect -46322 -27784 -46312 -27689
rect -46420 -27848 -46312 -27784
rect -46420 -27943 -46397 -27848
rect -46320 -27943 -46312 -27848
rect -46420 -28006 -46312 -27943
rect -46420 -28101 -46398 -28006
rect -46321 -28101 -46312 -28006
rect -46623 -28529 -46518 -28509
rect -46625 -28555 -46518 -28529
rect -55294 -29745 -55142 -29739
rect -55294 -29823 -55284 -29745
rect -55223 -29817 -55142 -29745
rect -55081 -29742 -54895 -29739
rect -55081 -29817 -54974 -29742
rect -55223 -29820 -54974 -29817
rect -54913 -29820 -54895 -29742
rect -55223 -29823 -54895 -29820
rect -55294 -33443 -54895 -29823
rect -54421 -28621 -54326 -28583
rect -54421 -28676 -54400 -28621
rect -54342 -28676 -54326 -28621
rect -54421 -28784 -54326 -28676
rect -54120 -28596 -54025 -28573
rect -54120 -28654 -54099 -28596
rect -54037 -28654 -54025 -28596
rect -54120 -28747 -54025 -28654
rect -54421 -28839 -54406 -28784
rect -54348 -28839 -54326 -28784
rect -54421 -28857 -54326 -28839
rect -54125 -28751 -54025 -28747
rect -54125 -28809 -54098 -28751
rect -54036 -28809 -54025 -28751
rect -54125 -28825 -54025 -28809
rect -46625 -28650 -46607 -28555
rect -46530 -28650 -46518 -28555
rect -46625 -28731 -46518 -28650
rect -54421 -31607 -54328 -28857
rect -55294 -33446 -55126 -33443
rect -55294 -33509 -55258 -33446
rect -55198 -33506 -55126 -33446
rect -55066 -33446 -54895 -33443
rect -55066 -33506 -54992 -33446
rect -55198 -33509 -54992 -33506
rect -54932 -33509 -54895 -33446
rect -55294 -36150 -54895 -33509
rect -54443 -31953 -54305 -31607
rect -54443 -32019 -54411 -31953
rect -54345 -32019 -54305 -31953
rect -54443 -32138 -54305 -32019
rect -54443 -32204 -54410 -32138
rect -54344 -32204 -54305 -32138
rect -54443 -35544 -54305 -32204
rect -54125 -34227 -54030 -28825
rect -46625 -28826 -46610 -28731
rect -46533 -28826 -46518 -28731
rect -53837 -28852 -53736 -28839
rect -53837 -28941 -53823 -28852
rect -53745 -28941 -53736 -28852
rect -53837 -28974 -53736 -28941
rect -53843 -29057 -53736 -28974
rect -53843 -29146 -53819 -29057
rect -53741 -29146 -53736 -29057
rect -53843 -29160 -53736 -29146
rect -46625 -28890 -46518 -28826
rect -46625 -28985 -46608 -28890
rect -46531 -28985 -46518 -28890
rect -46625 -29048 -46518 -28985
rect -46625 -29143 -46609 -29048
rect -46532 -29143 -46518 -29048
rect -53843 -33830 -53742 -29160
rect -46625 -29166 -46518 -29143
rect -46623 -30023 -46518 -29166
rect -46420 -30049 -46312 -28101
rect -45764 -30705 -45365 -22671
rect -45764 -30708 -45603 -30705
rect -45764 -30771 -45735 -30708
rect -45675 -30768 -45603 -30708
rect -45543 -30708 -45365 -30705
rect -45543 -30768 -45469 -30708
rect -45675 -30771 -45469 -30768
rect -45409 -30771 -45365 -30708
rect -45764 -31115 -45365 -30771
rect -45764 -31118 -45597 -31115
rect -45764 -31181 -45729 -31118
rect -45669 -31178 -45597 -31118
rect -45537 -31118 -45365 -31115
rect -45537 -31178 -45463 -31118
rect -45669 -31181 -45463 -31178
rect -45403 -31181 -45365 -31118
rect -50877 -31748 -50821 -31472
rect -50874 -32310 -50818 -32070
rect -53649 -33085 -53369 -33030
rect -53649 -33163 -53633 -33085
rect -53555 -33163 -53468 -33085
rect -53390 -33163 -53369 -33085
rect -53649 -33213 -53369 -33163
rect -53843 -33931 -53186 -33830
rect -54125 -34289 -54103 -34227
rect -54050 -34289 -54030 -34227
rect -54125 -34355 -54030 -34289
rect -54125 -34417 -54109 -34355
rect -54056 -34417 -54030 -34355
rect -54125 -34442 -54030 -34417
rect -50825 -34672 -50768 -34416
rect -54443 -35604 -54413 -35544
rect -54350 -35604 -54305 -35544
rect -54443 -35630 -54305 -35604
rect -55294 -36228 -55277 -36150
rect -55219 -36228 -55148 -36150
rect -55090 -36156 -54895 -36150
rect -55090 -36228 -55002 -36156
rect -55294 -36234 -55002 -36228
rect -54944 -36234 -54895 -36156
rect -55294 -36493 -54895 -36234
rect -45764 -36418 -45365 -31181
rect -45764 -36426 -45463 -36418
rect -55296 -36510 -54886 -36493
rect -55296 -36513 -54969 -36510
rect -55296 -36518 -55118 -36513
rect -55296 -36613 -55277 -36518
rect -55200 -36608 -55118 -36518
rect -55041 -36605 -54969 -36513
rect -54892 -36605 -54886 -36510
rect -55041 -36608 -54886 -36605
rect -55200 -36613 -54886 -36608
rect -55296 -36686 -54886 -36613
rect -55296 -36689 -54972 -36686
rect -55296 -36694 -55121 -36689
rect -55296 -36789 -55280 -36694
rect -55203 -36784 -55121 -36694
rect -55044 -36781 -54972 -36689
rect -54895 -36781 -54886 -36686
rect -55044 -36784 -54886 -36781
rect -55203 -36789 -54886 -36784
rect -55296 -36845 -54886 -36789
rect -55296 -36848 -54970 -36845
rect -55296 -36853 -55119 -36848
rect -55296 -36948 -55278 -36853
rect -55201 -36943 -55119 -36853
rect -55042 -36940 -54970 -36848
rect -54893 -36940 -54886 -36845
rect -55042 -36943 -54886 -36940
rect -55201 -36948 -54886 -36943
rect -55296 -37003 -54886 -36948
rect -55296 -37006 -54971 -37003
rect -55296 -37011 -55120 -37006
rect -55296 -37106 -55279 -37011
rect -55202 -37101 -55120 -37011
rect -55043 -37098 -54971 -37006
rect -54894 -37098 -54886 -37003
rect -55043 -37101 -54886 -37098
rect -55202 -37106 -54886 -37101
rect -55296 -37118 -54886 -37106
rect -45764 -36524 -45753 -36426
rect -45695 -36524 -45595 -36426
rect -45537 -36516 -45463 -36426
rect -45405 -36516 -45365 -36418
rect -45537 -36524 -45365 -36516
rect -55938 -37556 -55528 -37539
rect -55938 -37559 -55611 -37556
rect -55938 -37564 -55760 -37559
rect -55938 -37659 -55919 -37564
rect -55842 -37654 -55760 -37564
rect -55683 -37651 -55611 -37559
rect -55534 -37651 -55528 -37556
rect -55683 -37654 -55528 -37651
rect -55842 -37659 -55528 -37654
rect -55938 -37732 -55528 -37659
rect -55938 -37735 -55614 -37732
rect -55938 -37740 -55763 -37735
rect -55938 -37835 -55922 -37740
rect -55845 -37830 -55763 -37740
rect -55686 -37827 -55614 -37735
rect -55537 -37827 -55528 -37732
rect -55686 -37830 -55528 -37827
rect -55845 -37835 -55528 -37830
rect -55938 -37891 -55528 -37835
rect -55938 -37894 -55612 -37891
rect -55938 -37899 -55761 -37894
rect -55938 -37994 -55920 -37899
rect -55843 -37989 -55761 -37899
rect -55684 -37986 -55612 -37894
rect -55535 -37986 -55528 -37891
rect -55684 -37989 -55528 -37986
rect -55843 -37994 -55528 -37989
rect -55938 -38049 -55528 -37994
rect -55938 -38052 -55613 -38049
rect -55938 -38057 -55762 -38052
rect -55938 -38152 -55921 -38057
rect -55844 -38147 -55762 -38057
rect -55685 -38144 -55613 -38052
rect -55536 -38144 -55528 -38049
rect -55685 -38147 -55528 -38144
rect -55844 -38152 -55528 -38147
rect -55938 -38164 -55528 -38152
rect -55938 -38319 -55539 -38164
rect -55294 -38332 -54895 -37118
rect -45764 -37539 -45365 -36524
rect -44941 51363 -44542 55226
rect -35392 54813 -34993 55873
rect -34702 55848 -34303 55873
rect -34703 55831 -34293 55848
rect -34703 55828 -34376 55831
rect -34703 55823 -34525 55828
rect -34703 55728 -34684 55823
rect -34607 55733 -34525 55823
rect -34448 55736 -34376 55828
rect -34299 55736 -34293 55831
rect -34448 55733 -34293 55736
rect -34607 55728 -34293 55733
rect -34703 55655 -34293 55728
rect -34703 55652 -34379 55655
rect -34703 55647 -34528 55652
rect -34703 55552 -34687 55647
rect -34610 55557 -34528 55647
rect -34451 55560 -34379 55652
rect -34302 55560 -34293 55655
rect -34451 55557 -34293 55560
rect -34610 55552 -34293 55557
rect -34703 55496 -34293 55552
rect -34703 55493 -34377 55496
rect -34703 55488 -34526 55493
rect -34703 55393 -34685 55488
rect -34608 55398 -34526 55488
rect -34449 55401 -34377 55493
rect -34300 55401 -34293 55496
rect -34449 55398 -34293 55401
rect -34608 55393 -34293 55398
rect -34703 55338 -34293 55393
rect -34703 55335 -34378 55338
rect -34703 55330 -34527 55335
rect -34703 55235 -34686 55330
rect -34609 55240 -34527 55330
rect -34450 55243 -34378 55335
rect -34301 55243 -34293 55338
rect -34450 55240 -34293 55243
rect -34609 55235 -34293 55240
rect -34703 55223 -34293 55235
rect -35393 54796 -34983 54813
rect -35393 54793 -35066 54796
rect -35393 54788 -35215 54793
rect -35393 54693 -35374 54788
rect -35297 54698 -35215 54788
rect -35138 54701 -35066 54793
rect -34989 54701 -34983 54796
rect -35138 54698 -34983 54701
rect -35297 54693 -34983 54698
rect -35393 54620 -34983 54693
rect -35393 54617 -35069 54620
rect -35393 54612 -35218 54617
rect -35393 54517 -35377 54612
rect -35300 54522 -35218 54612
rect -35141 54525 -35069 54617
rect -34992 54525 -34983 54620
rect -35141 54522 -34983 54525
rect -35300 54517 -34983 54522
rect -35393 54461 -34983 54517
rect -35393 54458 -35067 54461
rect -35393 54453 -35216 54458
rect -35393 54358 -35375 54453
rect -35298 54363 -35216 54453
rect -35139 54366 -35067 54458
rect -34990 54366 -34983 54461
rect -35139 54363 -34983 54366
rect -35298 54358 -34983 54363
rect -35393 54303 -34983 54358
rect -35393 54300 -35068 54303
rect -35393 54295 -35217 54300
rect -35393 54200 -35376 54295
rect -35299 54205 -35217 54295
rect -35140 54208 -35068 54300
rect -34991 54208 -34983 54303
rect -35140 54205 -34983 54208
rect -35299 54200 -34983 54205
rect -35393 54188 -34983 54200
rect -36027 53631 -35933 53639
rect -36052 53615 -35933 53631
rect -36052 53520 -36016 53615
rect -35939 53520 -35933 53615
rect -36052 53439 -35933 53520
rect -36052 53344 -36019 53439
rect -35942 53344 -35933 53439
rect -36052 53280 -35933 53344
rect -36052 53185 -36017 53280
rect -35940 53185 -35933 53280
rect -36052 53122 -35933 53185
rect -36052 53027 -36018 53122
rect -35941 53027 -35933 53122
rect -36052 53017 -35933 53027
rect -43768 52594 -43665 52615
rect -43768 52520 -43752 52594
rect -43678 52520 -43665 52594
rect -43768 52415 -43665 52520
rect -43768 52341 -43752 52415
rect -43678 52341 -43665 52415
rect -43768 52323 -43665 52341
rect -36255 52563 -36150 52595
rect -36255 52468 -36236 52563
rect -36159 52468 -36150 52563
rect -36255 52387 -36150 52468
rect -44941 51306 -44929 51363
rect -44876 51306 -44814 51363
rect -44761 51362 -44542 51363
rect -44761 51306 -44678 51362
rect -44941 51305 -44678 51306
rect -44625 51305 -44542 51362
rect -44941 47938 -44542 51305
rect -44941 47935 -44783 47938
rect -44941 47872 -44915 47935
rect -44855 47875 -44783 47935
rect -44723 47935 -44542 47938
rect -44723 47875 -44649 47935
rect -44855 47872 -44649 47875
rect -44589 47872 -44542 47935
rect -44941 47567 -44542 47872
rect -44941 47564 -44776 47567
rect -44941 47501 -44908 47564
rect -44848 47504 -44776 47564
rect -44716 47564 -44542 47567
rect -44716 47504 -44642 47564
rect -44848 47501 -44642 47504
rect -44582 47501 -44542 47564
rect -44941 43041 -44542 47501
rect -43959 48973 -43868 48998
rect -43959 48913 -43940 48973
rect -43888 48913 -43868 48973
rect -43959 48854 -43868 48913
rect -43959 48794 -43938 48854
rect -43886 48794 -43868 48854
rect -43959 44795 -43868 48794
rect -43752 46641 -43678 52323
rect -36255 52292 -36239 52387
rect -36162 52292 -36150 52387
rect -36255 52228 -36150 52292
rect -43467 52165 -43344 52179
rect -43467 52067 -43453 52165
rect -43355 52067 -43344 52165
rect -43467 51951 -43344 52067
rect -43467 51851 -43454 51951
rect -43354 51851 -43344 51951
rect -43467 51842 -43344 51851
rect -36255 52133 -36237 52228
rect -36160 52133 -36150 52228
rect -36255 52070 -36150 52133
rect -36255 51975 -36238 52070
rect -36161 51975 -36150 52070
rect -43454 47213 -43354 51842
rect -36255 51581 -36150 51975
rect -36255 51525 -36227 51581
rect -36172 51525 -36150 51581
rect -36255 51035 -36150 51525
rect -36052 51442 -35944 53017
rect -36052 51386 -36021 51442
rect -35966 51386 -35944 51442
rect -36052 51021 -35944 51386
rect -42893 49984 -42770 49998
rect -42893 49905 -42873 49984
rect -42782 49905 -42770 49984
rect -42893 49832 -42770 49905
rect -40506 49886 -39911 49942
rect -42893 49753 -42877 49832
rect -42786 49753 -42770 49832
rect -42893 49741 -42770 49753
rect -40509 49521 -40453 49748
rect -40493 48919 -40437 48925
rect -40451 48865 -40437 48919
rect -40493 48686 -40437 48865
rect -35392 48779 -34993 54188
rect -35392 48776 -35248 48779
rect -35392 48713 -35380 48776
rect -35320 48716 -35248 48776
rect -35188 48776 -34993 48779
rect -35188 48716 -35114 48776
rect -35320 48713 -35114 48716
rect -35054 48713 -34993 48776
rect -43479 47197 -43171 47213
rect -43479 47097 -43454 47197
rect -43354 47196 -43171 47197
rect -43354 47098 -43282 47196
rect -43184 47098 -43171 47196
rect -43354 47097 -43171 47098
rect -43479 47079 -43171 47097
rect -43767 46629 -43510 46641
rect -43767 46555 -43752 46629
rect -43678 46555 -43597 46629
rect -43523 46555 -43510 46629
rect -43767 46539 -43510 46555
rect -40457 46417 -40400 46592
rect -40403 46358 -40400 46417
rect -40457 46355 -40400 46358
rect -43959 44733 -43938 44795
rect -43884 44733 -43868 44795
rect -43959 44653 -43868 44733
rect -43959 44591 -43941 44653
rect -43887 44591 -43868 44653
rect -43959 44568 -43868 44591
rect -36099 45231 -35991 45268
rect -36099 45136 -36083 45231
rect -36006 45136 -35991 45231
rect -36099 45055 -35991 45136
rect -36099 44960 -36086 45055
rect -36009 44960 -35991 45055
rect -36099 44896 -35991 44960
rect -36099 44801 -36084 44896
rect -36007 44801 -35991 44896
rect -36099 44738 -35991 44801
rect -36099 44643 -36085 44738
rect -36008 44643 -35991 44738
rect -43648 44256 -43256 44272
rect -43648 44145 -43630 44256
rect -43519 44255 -43256 44256
rect -43519 44146 -43378 44255
rect -43268 44146 -43256 44255
rect -43519 44145 -43256 44146
rect -43648 44134 -43256 44145
rect -36302 44188 -36197 44234
rect -44941 43040 -44635 43041
rect -44941 43039 -44782 43040
rect -44941 42965 -44931 43039
rect -44870 42966 -44782 43039
rect -44721 42967 -44635 43040
rect -44574 42967 -44542 43041
rect -44721 42966 -44542 42967
rect -44870 42965 -44542 42966
rect -44941 39752 -44542 42965
rect -44941 39750 -44669 39752
rect -44941 39694 -44918 39750
rect -44866 39694 -44788 39750
rect -44736 39696 -44669 39750
rect -44617 39696 -44542 39752
rect -44736 39694 -44542 39696
rect -44941 39379 -44542 39694
rect -44941 39377 -44659 39379
rect -44941 39321 -44908 39377
rect -44856 39321 -44778 39377
rect -44726 39323 -44659 39377
rect -44607 39323 -44542 39379
rect -44726 39321 -44542 39323
rect -44941 37771 -44542 39321
rect -44941 37768 -44645 37771
rect -44941 37694 -44930 37768
rect -44869 37766 -44645 37768
rect -44869 37694 -44795 37766
rect -44941 37692 -44795 37694
rect -44734 37697 -44645 37766
rect -44584 37697 -44542 37771
rect -44734 37692 -44542 37697
rect -44941 34593 -44542 37692
rect -44941 34520 -44928 34593
rect -44866 34592 -44542 34593
rect -44866 34520 -44802 34592
rect -44941 34519 -44802 34520
rect -44740 34519 -44647 34592
rect -44585 34519 -44542 34592
rect -44941 30875 -44542 34519
rect -44941 30872 -44651 30875
rect -44941 30871 -44805 30872
rect -44941 30798 -44932 30871
rect -44866 30799 -44805 30871
rect -44739 30802 -44651 30872
rect -44585 30802 -44542 30875
rect -44739 30799 -44542 30802
rect -44866 30798 -44542 30799
rect -44941 26144 -44542 30798
rect -44941 26054 -44927 26144
rect -44861 26142 -44645 26144
rect -44861 26054 -44783 26142
rect -44941 26052 -44783 26054
rect -44717 26054 -44645 26142
rect -44579 26054 -44542 26144
rect -44717 26052 -44542 26054
rect -44941 22441 -44542 26052
rect -44941 22439 -44681 22441
rect -44941 22437 -44806 22439
rect -44941 22381 -44926 22437
rect -44874 22383 -44806 22437
rect -44754 22385 -44681 22439
rect -44629 22385 -44542 22441
rect -44754 22383 -44542 22385
rect -44874 22381 -44542 22383
rect -44941 17307 -44542 22381
rect -44020 40786 -43854 40804
rect -44020 40732 -44003 40786
rect -43874 40732 -43854 40786
rect -44020 40667 -43854 40732
rect -44020 40613 -44003 40667
rect -43874 40613 -43854 40667
rect -44020 40553 -43854 40613
rect -44020 40499 -44004 40553
rect -43875 40499 -43854 40553
rect -44020 32262 -43854 40499
rect -43642 38491 -43560 44134
rect -36302 44093 -36289 44188
rect -36212 44093 -36197 44188
rect -36302 44012 -36197 44093
rect -43394 43936 -43015 43953
rect -43394 43825 -43380 43936
rect -43269 43935 -43015 43936
rect -43269 43826 -43132 43935
rect -43023 43826 -43015 43935
rect -43269 43825 -43015 43826
rect -43394 43813 -43015 43825
rect -36302 43917 -36292 44012
rect -36215 43917 -36197 44012
rect -36302 43853 -36197 43917
rect -43390 39001 -43308 43813
rect -36302 43758 -36290 43853
rect -36213 43758 -36197 43853
rect -36302 43695 -36197 43758
rect -36302 43600 -36291 43695
rect -36214 43600 -36197 43695
rect -36302 43410 -36197 43600
rect -36302 43354 -36274 43410
rect -36219 43354 -36197 43410
rect -36302 42729 -36197 43354
rect -36099 43271 -35991 44643
rect -36099 43215 -36068 43271
rect -36013 43215 -35991 43271
rect -36099 42802 -35991 43215
rect -42874 41787 -42751 41801
rect -42874 41708 -42854 41787
rect -42763 41708 -42751 41787
rect -42874 41635 -42751 41708
rect -42874 41556 -42858 41635
rect -42767 41556 -42751 41635
rect -42874 41544 -42751 41556
rect -40556 41771 -40500 41777
rect -40556 41715 -39958 41771
rect -40556 41515 -40500 41715
rect -40553 40748 -40497 40763
rect -40553 40694 -40552 40748
rect -40498 40694 -40497 40748
rect -40553 40515 -40497 40694
rect -35392 40573 -34993 48713
rect -35392 40570 -35099 40573
rect -35392 40568 -35248 40570
rect -35392 40512 -35369 40568
rect -35317 40514 -35248 40568
rect -35196 40517 -35099 40570
rect -35047 40517 -34993 40573
rect -35196 40514 -34993 40517
rect -35317 40512 -34993 40514
rect -43390 38919 -42855 39001
rect -43755 38459 -43481 38491
rect -43755 38454 -43595 38459
rect -43755 38400 -43728 38454
rect -43673 38405 -43595 38454
rect -43540 38405 -43481 38459
rect -43673 38400 -43481 38405
rect -43755 38368 -43481 38400
rect -44020 32203 -44000 32262
rect -43873 32203 -43854 32262
rect -44020 32150 -43854 32203
rect -44020 32091 -44001 32150
rect -43874 32091 -43854 32150
rect -44020 32024 -43854 32091
rect -44020 31965 -44004 32024
rect -43877 31965 -43854 32024
rect -44020 21860 -43854 31965
rect -43642 29959 -43560 38368
rect -43390 30472 -43308 38919
rect -40504 38246 -40447 38424
rect -40450 38187 -40447 38246
rect -40504 38176 -40447 38187
rect -36042 37020 -35934 37064
rect -36042 36925 -36023 37020
rect -35946 36925 -35934 37020
rect -36042 36844 -35934 36925
rect -36042 36749 -36026 36844
rect -35949 36749 -35934 36844
rect -36042 36685 -35934 36749
rect -36042 36590 -36024 36685
rect -35947 36590 -35934 36685
rect -36042 36527 -35934 36590
rect -36042 36432 -36025 36527
rect -35948 36432 -35934 36527
rect -36232 35787 -36138 35790
rect -36245 35766 -36138 35787
rect -36245 35671 -36221 35766
rect -36144 35671 -36138 35766
rect -36245 35590 -36138 35671
rect -36245 35495 -36224 35590
rect -36147 35495 -36138 35590
rect -36245 35431 -36138 35495
rect -36245 35336 -36222 35431
rect -36145 35336 -36138 35431
rect -36245 35273 -36138 35336
rect -36245 35178 -36223 35273
rect -36146 35178 -36138 35273
rect -36245 35168 -36138 35178
rect -36245 34112 -36140 35168
rect -36042 34298 -35934 36432
rect -35392 33448 -34993 40512
rect -35392 33444 -35112 33448
rect -35392 33440 -35237 33444
rect -35392 33357 -35379 33440
rect -35309 33361 -35237 33440
rect -35167 33365 -35112 33444
rect -35042 33365 -34993 33448
rect -35167 33361 -34993 33365
rect -35309 33357 -34993 33361
rect -42810 33264 -42687 33278
rect -42810 33185 -42790 33264
rect -42699 33185 -42687 33264
rect -42810 33112 -42687 33185
rect -42810 33033 -42794 33112
rect -42703 33033 -42687 33112
rect -42810 33021 -42687 33033
rect -40499 32608 -40443 32870
rect -40496 31992 -40440 32225
rect -43129 31319 -43006 31333
rect -43129 31240 -43109 31319
rect -43018 31240 -43006 31319
rect -43129 31167 -43006 31240
rect -43129 31088 -43113 31167
rect -43022 31088 -43006 31167
rect -43129 31076 -43006 31088
rect -43390 30390 -42801 30472
rect -43726 29932 -43530 29959
rect -43726 29871 -43708 29932
rect -43648 29871 -43596 29932
rect -43537 29871 -43530 29932
rect -43726 29840 -43530 29871
rect -43642 28983 -43560 29840
rect -43390 29171 -43308 30390
rect -40447 29659 -40390 29902
rect -43404 29155 -43296 29171
rect -43404 29075 -43389 29155
rect -43309 29075 -43296 29155
rect -43404 28987 -43296 29075
rect -43654 28969 -43544 28983
rect -43654 28887 -43642 28969
rect -43560 28887 -43544 28969
rect -43404 28905 -43390 28987
rect -43308 28905 -43296 28987
rect -43404 28888 -43296 28905
rect -43654 28759 -43544 28887
rect -43654 28677 -43642 28759
rect -43560 28677 -43544 28759
rect -43654 28666 -43544 28677
rect -36242 28459 -36134 28494
rect -36242 28364 -36223 28459
rect -36146 28364 -36134 28459
rect -36242 28283 -36134 28364
rect -36242 28188 -36226 28283
rect -36149 28188 -36134 28283
rect -36242 28124 -36134 28188
rect -36242 28029 -36224 28124
rect -36147 28029 -36134 28124
rect -36242 27966 -36134 28029
rect -36242 27871 -36225 27966
rect -36148 27871 -36134 27966
rect -36445 27344 -36340 27398
rect -36445 27249 -36430 27344
rect -36353 27249 -36340 27344
rect -36445 27168 -36340 27249
rect -36445 27073 -36433 27168
rect -36356 27073 -36340 27168
rect -36445 27009 -36340 27073
rect -36445 26914 -36431 27009
rect -36354 26914 -36340 27009
rect -36445 26851 -36340 26914
rect -36445 26756 -36432 26851
rect -36355 26756 -36340 26851
rect -36445 25861 -36340 26756
rect -36242 25870 -36134 27871
rect -43024 24862 -42901 24867
rect -43024 24853 -42898 24862
rect -43024 24774 -43004 24853
rect -42913 24801 -42898 24853
rect -42913 24774 -42755 24801
rect -43024 24701 -42755 24774
rect -43024 24622 -43008 24701
rect -42917 24622 -42755 24701
rect -43024 24610 -42755 24622
rect -43681 23806 -43519 23849
rect -43681 23694 -43648 23806
rect -43539 23694 -43519 23806
rect -43681 23569 -43519 23694
rect -43681 23457 -43656 23569
rect -43547 23457 -43519 23569
rect -43681 22283 -43519 23457
rect -43323 22913 -43200 22927
rect -43323 22834 -43303 22913
rect -43212 22834 -43200 22913
rect -43323 22761 -43200 22834
rect -43323 22682 -43307 22761
rect -43216 22682 -43200 22761
rect -43323 22670 -43200 22682
rect -43681 22121 -43239 22283
rect -44020 21694 -43747 21860
rect -44941 17229 -44933 17307
rect -44868 17305 -44542 17307
rect -44868 17229 -44796 17305
rect -44941 17227 -44796 17229
rect -44731 17227 -44650 17305
rect -44585 17227 -44542 17305
rect -44941 13276 -44542 17227
rect -44941 13275 -44679 13276
rect -44941 13271 -44810 13275
rect -44941 13207 -44931 13271
rect -44876 13211 -44810 13271
rect -44755 13212 -44679 13275
rect -44624 13212 -44542 13276
rect -44755 13211 -44542 13212
rect -44876 13207 -44542 13211
rect -44941 4379 -44542 13207
rect -44941 4377 -44798 4379
rect -44941 4302 -44929 4377
rect -44877 4304 -44798 4377
rect -44746 4374 -44542 4379
rect -44746 4304 -44652 4374
rect -44877 4302 -44652 4304
rect -44941 4299 -44652 4302
rect -44600 4299 -44542 4374
rect -44941 449 -44542 4299
rect -43913 17557 -43747 21694
rect -43401 18624 -43239 22121
rect -43073 21021 -43015 21290
rect -43083 20362 -43005 21021
rect -42865 20701 -42755 24610
rect -40699 24056 -40643 24249
rect -40696 23587 -40640 23822
rect -35392 23261 -34993 33357
rect -35392 23260 -35240 23261
rect -35392 23200 -35376 23260
rect -35316 23201 -35240 23260
rect -35180 23201 -35086 23261
rect -35026 23201 -34993 23261
rect -35316 23200 -34993 23201
rect -40647 21236 -40590 21478
rect -42865 20591 -42531 20701
rect -43092 20351 -42762 20362
rect -43092 20350 -42887 20351
rect -43092 20239 -43080 20350
rect -42969 20239 -42887 20350
rect -43092 20238 -42887 20239
rect -42774 20238 -42762 20351
rect -43092 20230 -42762 20238
rect -43413 18423 -43228 18624
rect -43413 18355 -43384 18423
rect -43412 18322 -43384 18355
rect -43283 18355 -43228 18423
rect -43283 18322 -43229 18355
rect -43412 18231 -43229 18322
rect -43412 18130 -43367 18231
rect -43266 18130 -43229 18231
rect -43412 18056 -43229 18130
rect -43412 17955 -43377 18056
rect -43276 17955 -43229 18056
rect -43412 17905 -43229 17955
rect -43913 17498 -43887 17557
rect -43780 17498 -43747 17557
rect -43913 17430 -43747 17498
rect -43913 17371 -43883 17430
rect -43776 17371 -43747 17430
rect -43913 17307 -43747 17371
rect -43913 17248 -43886 17307
rect -43779 17248 -43747 17307
rect -43913 14626 -43747 17248
rect -42976 15622 -42889 15643
rect -42976 15566 -42963 15622
rect -42907 15566 -42889 15622
rect -42976 15511 -42889 15566
rect -42976 15455 -42967 15511
rect -42911 15455 -42889 15511
rect -42976 15440 -42889 15455
rect -43913 14559 -43866 14626
rect -43794 14559 -43747 14626
rect -43913 14434 -43747 14559
rect -43913 14367 -43869 14434
rect -43797 14367 -43747 14434
rect -43913 1951 -43747 14367
rect -42641 13749 -42531 20591
rect -36212 19437 -36111 19442
rect -36217 19416 -36109 19437
rect -36217 19321 -36194 19416
rect -36117 19321 -36109 19416
rect -36217 19240 -36109 19321
rect -36217 19145 -36197 19240
rect -36120 19145 -36109 19240
rect -36217 19081 -36109 19145
rect -36217 18986 -36195 19081
rect -36118 18986 -36109 19081
rect -36217 18923 -36109 18986
rect -36217 18828 -36196 18923
rect -36119 18828 -36109 18923
rect -36420 18326 -36315 18383
rect -36420 18231 -36400 18326
rect -36323 18231 -36315 18326
rect -36420 18150 -36315 18231
rect -36420 18055 -36403 18150
rect -36326 18055 -36315 18150
rect -36420 17991 -36315 18055
rect -36420 17896 -36401 17991
rect -36324 17896 -36315 17991
rect -36420 17833 -36315 17896
rect -36420 17738 -36402 17833
rect -36325 17738 -36315 17833
rect -36420 16622 -36315 17738
rect -36217 16643 -36109 18828
rect -35392 16206 -34993 23200
rect -35392 16201 -35081 16206
rect -35392 16200 -35217 16201
rect -35392 16144 -35367 16200
rect -35314 16145 -35217 16200
rect -35164 16150 -35081 16201
rect -35028 16150 -34993 16206
rect -35164 16145 -34993 16150
rect -35314 16144 -34993 16145
rect -40674 14843 -40618 15098
rect -40671 14395 -40615 14658
rect -42710 13722 -42466 13749
rect -42710 13718 -42561 13722
rect -43281 13664 -43194 13685
rect -43281 13608 -43268 13664
rect -43212 13608 -43194 13664
rect -42710 13635 -42693 13718
rect -42628 13639 -42561 13718
rect -42496 13639 -42466 13722
rect -42628 13635 -42466 13639
rect -42710 13623 -42466 13635
rect -42641 13622 -42531 13623
rect -43281 13553 -43194 13608
rect -43281 13497 -43272 13553
rect -43216 13497 -43194 13553
rect -43281 13482 -43194 13497
rect -43386 12349 -43136 12366
rect -43386 12274 -43377 12349
rect -43302 12274 -43224 12349
rect -43149 12274 -43136 12349
rect -43386 12264 -43136 12274
rect -43274 11535 -43188 12264
rect -40622 12063 -40565 12307
rect -43488 11520 -43177 11535
rect -43488 11519 -43278 11520
rect -43488 11435 -43482 11519
rect -43398 11435 -43278 11519
rect -43488 11434 -43278 11435
rect -43192 11434 -43177 11520
rect -43488 11422 -43177 11434
rect -35392 10398 -34993 16144
rect -35392 10392 -35095 10398
rect -35392 10339 -35373 10392
rect -35318 10339 -35242 10392
rect -35187 10345 -35095 10392
rect -35040 10345 -34993 10398
rect -35187 10339 -34993 10345
rect -35392 9506 -34993 10339
rect -35392 9505 -35101 9506
rect -35392 9500 -35239 9505
rect -35392 9447 -35378 9500
rect -35323 9452 -35239 9500
rect -35184 9453 -35101 9505
rect -35046 9453 -34993 9506
rect -35184 9452 -34993 9453
rect -35323 9447 -34993 9452
rect -35392 8566 -34993 9447
rect -35392 8562 -35117 8566
rect -35392 8555 -35249 8562
rect -35392 8502 -35372 8555
rect -35317 8509 -35249 8555
rect -35194 8513 -35117 8562
rect -35062 8513 -34993 8566
rect -35194 8509 -34993 8513
rect -35317 8502 -34993 8509
rect -35392 7685 -34993 8502
rect -35392 7678 -35125 7685
rect -35392 7671 -35256 7678
rect -35392 7618 -35382 7671
rect -35327 7625 -35256 7671
rect -35201 7632 -35125 7678
rect -35070 7632 -34993 7685
rect -35201 7625 -34993 7632
rect -35327 7618 -34993 7625
rect -36037 7419 -35929 7430
rect -36037 7393 -35926 7419
rect -36037 7298 -36009 7393
rect -35932 7298 -35926 7393
rect -36037 7217 -35926 7298
rect -36037 7122 -36012 7217
rect -35935 7122 -35926 7217
rect -36037 7058 -35926 7122
rect -36037 6963 -36010 7058
rect -35933 6963 -35926 7058
rect -36037 6900 -35926 6963
rect -36037 6805 -36011 6900
rect -35934 6805 -35926 6900
rect -36037 6782 -35926 6805
rect -36240 6180 -36135 6198
rect -36240 6154 -36134 6180
rect -36240 6059 -36217 6154
rect -36140 6059 -36134 6154
rect -36240 5978 -36134 6059
rect -36240 5883 -36220 5978
rect -36143 5883 -36134 5978
rect -36240 5819 -36134 5883
rect -36240 5724 -36218 5819
rect -36141 5724 -36134 5819
rect -36240 5661 -36134 5724
rect -36240 5566 -36219 5661
rect -36142 5566 -36134 5661
rect -36240 5543 -36134 5566
rect -36240 3878 -36135 5543
rect -36037 3871 -35929 6782
rect -35392 6770 -34993 7618
rect -35392 6765 -35244 6770
rect -35392 6712 -35371 6765
rect -35316 6717 -35244 6765
rect -35189 6769 -34993 6770
rect -35189 6717 -35117 6769
rect -35316 6716 -35117 6717
rect -35062 6716 -34993 6769
rect -35316 6712 -34993 6716
rect -35392 5858 -34993 6712
rect -35392 5852 -35243 5858
rect -35392 5799 -35369 5852
rect -35314 5805 -35243 5852
rect -35188 5856 -34993 5858
rect -35188 5805 -35103 5856
rect -35314 5803 -35103 5805
rect -35048 5803 -34993 5856
rect -35314 5799 -34993 5803
rect -35392 3288 -34993 5799
rect -35392 3287 -35080 3288
rect -35392 3284 -35226 3287
rect -35392 3228 -35368 3284
rect -35314 3231 -35226 3284
rect -35172 3232 -35080 3287
rect -35026 3232 -34993 3288
rect -35172 3231 -34993 3232
rect -35314 3228 -34993 3231
rect -42791 2816 -42704 2837
rect -42791 2760 -42778 2816
rect -42722 2760 -42704 2816
rect -42791 2757 -42704 2760
rect -42791 2705 -42489 2757
rect -42791 2649 -42782 2705
rect -42726 2664 -42489 2705
rect -42726 2649 -42704 2664
rect -42791 2634 -42704 2649
rect -43913 1888 -43868 1951
rect -43800 1888 -43747 1951
rect -43913 1786 -43747 1888
rect -43913 1723 -43869 1786
rect -43801 1723 -43747 1786
rect -43913 1584 -43747 1723
rect -44941 389 -44930 449
rect -44864 448 -44679 449
rect -44864 389 -44809 448
rect -44941 388 -44809 389
rect -44743 389 -44679 448
rect -44613 389 -44542 449
rect -44743 388 -44542 389
rect -44941 -875 -44542 388
rect -44941 -877 -44631 -875
rect -44941 -879 -44782 -877
rect -44941 -969 -44917 -879
rect -44861 -967 -44782 -879
rect -44726 -965 -44631 -877
rect -44575 -965 -44542 -875
rect -44726 -967 -44542 -965
rect -44861 -969 -44542 -967
rect -44941 -4754 -44542 -969
rect -44941 -4851 -44927 -4754
rect -44863 -4851 -44778 -4754
rect -44714 -4851 -44630 -4754
rect -44566 -4851 -44542 -4754
rect -44941 -8515 -44542 -4851
rect -44941 -8517 -44654 -8515
rect -44941 -8518 -44795 -8517
rect -44941 -8579 -44930 -8518
rect -44874 -8578 -44795 -8518
rect -44739 -8576 -44654 -8517
rect -44598 -8576 -44542 -8515
rect -44739 -8578 -44542 -8576
rect -44874 -8579 -44542 -8578
rect -44941 -9706 -44542 -8579
rect -44941 -9712 -44788 -9706
rect -44941 -9791 -44928 -9712
rect -44868 -9785 -44788 -9712
rect -44728 -9785 -44634 -9706
rect -44574 -9785 -44542 -9706
rect -44868 -9791 -44542 -9785
rect -44941 -13492 -44542 -9791
rect -44941 -13494 -44803 -13492
rect -44941 -13563 -44924 -13494
rect -44870 -13561 -44803 -13494
rect -44749 -13561 -44652 -13492
rect -44598 -13561 -44542 -13492
rect -44870 -13563 -44542 -13561
rect -44941 -17444 -44542 -13563
rect -44356 1418 -43747 1584
rect -44356 -15957 -44190 1418
rect -43147 907 -43060 928
rect -43147 851 -43134 907
rect -43078 851 -43060 907
rect -43147 796 -43060 851
rect -43147 740 -43138 796
rect -43082 740 -43060 796
rect -43147 725 -43060 740
rect -42582 21 -42489 2664
rect -40494 2066 -40438 2266
rect -40491 1577 -40435 1814
rect -42678 -72 -42489 21
rect -43498 -468 -43094 -454
rect -43498 -469 -43184 -468
rect -43498 -544 -43346 -469
rect -43271 -544 -43184 -469
rect -43498 -545 -43184 -544
rect -43107 -545 -43094 -468
rect -43498 -558 -43094 -545
rect -43498 -1017 -43394 -558
rect -43498 -1076 -43474 -1017
rect -43417 -1076 -43394 -1017
rect -43498 -1140 -43394 -1076
rect -43498 -1199 -43473 -1140
rect -43416 -1199 -43394 -1140
rect -43801 -2965 -43647 -2861
rect -43801 -3122 -43764 -2965
rect -43673 -3122 -43647 -2965
rect -43801 -3245 -43647 -3122
rect -43801 -3402 -43772 -3245
rect -43681 -3402 -43647 -3245
rect -43801 -7123 -43647 -3402
rect -43801 -7205 -43750 -7123
rect -43682 -7205 -43647 -7123
rect -43801 -7315 -43647 -7205
rect -43801 -7397 -43750 -7315
rect -43682 -7397 -43647 -7315
rect -43801 -12447 -43647 -7397
rect -43498 -9435 -43394 -1199
rect -43300 -1035 -42787 -945
rect -43300 -1149 -43210 -1035
rect -43300 -1204 -43282 -1149
rect -43229 -1204 -43210 -1149
rect -43300 -1259 -43210 -1204
rect -43300 -1314 -43281 -1259
rect -43228 -1314 -43210 -1259
rect -43300 -8901 -43210 -1314
rect -42678 -5912 -42585 -72
rect -40442 -749 -40385 -516
rect -36060 -2455 -35952 -2392
rect -36060 -2550 -36040 -2455
rect -35963 -2550 -35952 -2455
rect -36060 -2631 -35952 -2550
rect -36060 -2726 -36043 -2631
rect -35966 -2726 -35952 -2631
rect -36060 -2790 -35952 -2726
rect -36060 -2885 -36041 -2790
rect -35964 -2885 -35952 -2790
rect -36060 -2948 -35952 -2885
rect -36060 -3043 -36042 -2948
rect -35965 -3043 -35952 -2948
rect -36263 -3503 -36158 -3480
rect -36265 -3529 -36158 -3503
rect -36265 -3624 -36247 -3529
rect -36170 -3624 -36158 -3529
rect -36265 -3705 -36158 -3624
rect -36265 -3800 -36250 -3705
rect -36173 -3800 -36158 -3705
rect -36265 -3864 -36158 -3800
rect -36265 -3959 -36248 -3864
rect -36171 -3959 -36158 -3864
rect -36265 -4022 -36158 -3959
rect -36265 -4117 -36249 -4022
rect -36172 -4117 -36158 -4022
rect -36265 -4140 -36158 -4117
rect -36263 -5177 -36158 -4140
rect -36060 -5094 -35952 -3043
rect -42678 -6005 -42513 -5912
rect -42812 -6147 -42725 -6126
rect -42812 -6203 -42799 -6147
rect -42743 -6203 -42725 -6147
rect -42812 -6258 -42725 -6203
rect -42812 -6314 -42803 -6258
rect -42747 -6314 -42725 -6258
rect -42812 -6329 -42725 -6314
rect -43130 -8034 -42977 -8009
rect -43130 -8116 -43097 -8034
rect -43015 -8116 -42977 -8034
rect -42606 -8102 -42513 -6005
rect -40517 -6917 -40461 -6764
rect -40514 -7389 -40458 -7144
rect -35392 -7552 -34993 3228
rect -35392 -7554 -35076 -7552
rect -35392 -7616 -35376 -7554
rect -35316 -7616 -35231 -7554
rect -35171 -7614 -35076 -7554
rect -35016 -7614 -34993 -7552
rect -35171 -7616 -34993 -7614
rect -43130 -8199 -42977 -8116
rect -43130 -8281 -43097 -8199
rect -43015 -8281 -42977 -8199
rect -42686 -8133 -42426 -8102
rect -42686 -8137 -42509 -8133
rect -42686 -8223 -42673 -8137
rect -42605 -8219 -42509 -8137
rect -42441 -8219 -42426 -8133
rect -42605 -8223 -42426 -8219
rect -42686 -8234 -42426 -8223
rect -42606 -8236 -42513 -8234
rect -43130 -8294 -42977 -8281
rect -43300 -8991 -42817 -8901
rect -42891 -9203 -42833 -8991
rect -43498 -9445 -43224 -9435
rect -43498 -9502 -43466 -9445
rect -43414 -9446 -43224 -9445
rect -43414 -9502 -43341 -9446
rect -43498 -9503 -43341 -9502
rect -43289 -9503 -43224 -9446
rect -43498 -9539 -43224 -9503
rect -40465 -9725 -40408 -9488
rect -36222 -11377 -36114 -11333
rect -36222 -11472 -36198 -11377
rect -36121 -11472 -36114 -11377
rect -36222 -11553 -36114 -11472
rect -36222 -11648 -36201 -11553
rect -36124 -11648 -36114 -11553
rect -36222 -11712 -36114 -11648
rect -36222 -11807 -36199 -11712
rect -36122 -11807 -36114 -11712
rect -36222 -11870 -36114 -11807
rect -36222 -11965 -36200 -11870
rect -36123 -11965 -36114 -11870
rect -43801 -12607 -43772 -12447
rect -43666 -12607 -43647 -12447
rect -43801 -12727 -43647 -12607
rect -43801 -12887 -43777 -12727
rect -43671 -12887 -43647 -12727
rect -43801 -12915 -43647 -12887
rect -36425 -12422 -36320 -12381
rect -36425 -12517 -36403 -12422
rect -36326 -12517 -36320 -12422
rect -36425 -12598 -36320 -12517
rect -36425 -12693 -36406 -12598
rect -36329 -12693 -36320 -12598
rect -36425 -12757 -36320 -12693
rect -36425 -12852 -36404 -12757
rect -36327 -12852 -36320 -12757
rect -36425 -12915 -36320 -12852
rect -36425 -13010 -36405 -12915
rect -36328 -13010 -36320 -12915
rect -36425 -14080 -36320 -13010
rect -36222 -14203 -36114 -11965
rect -35392 -14543 -34993 -7616
rect -35392 -14544 -35093 -14543
rect -35392 -14547 -35245 -14544
rect -35392 -14627 -35385 -14547
rect -35314 -14624 -35245 -14547
rect -35174 -14623 -35093 -14544
rect -35022 -14623 -34993 -14543
rect -35174 -14624 -34993 -14623
rect -35314 -14627 -34993 -14624
rect -42985 -15099 -42898 -15078
rect -42985 -15155 -42972 -15099
rect -42916 -15155 -42898 -15099
rect -42985 -15158 -42898 -15155
rect -42985 -15210 -42730 -15158
rect -42985 -15266 -42976 -15210
rect -42920 -15221 -42730 -15210
rect -42920 -15266 -42898 -15221
rect -42985 -15281 -42898 -15266
rect -44356 -16048 -43695 -15957
rect -44356 -16137 -43829 -16048
rect -43717 -16137 -43695 -16048
rect -44356 -16220 -43695 -16137
rect -43849 -16278 -43695 -16220
rect -43849 -16367 -43832 -16278
rect -43720 -16367 -43695 -16278
rect -43849 -16393 -43695 -16367
rect -44941 -17502 -44930 -17444
rect -44876 -17445 -44652 -17444
rect -44876 -17502 -44802 -17445
rect -44941 -17503 -44802 -17502
rect -44748 -17502 -44652 -17445
rect -44598 -17502 -44542 -17444
rect -44748 -17503 -44542 -17502
rect -44941 -18416 -44542 -17503
rect -44941 -18417 -44640 -18416
rect -44941 -18419 -44785 -18417
rect -44941 -18503 -44929 -18419
rect -44866 -18501 -44785 -18419
rect -44722 -18500 -44640 -18417
rect -44577 -18500 -44542 -18416
rect -44722 -18501 -44542 -18500
rect -44866 -18503 -44542 -18501
rect -44941 -21619 -44542 -18503
rect -44941 -21621 -44610 -21619
rect -44941 -21688 -44932 -21621
rect -44878 -21622 -44610 -21621
rect -44878 -21688 -44775 -21622
rect -44941 -21689 -44775 -21688
rect -44721 -21686 -44610 -21622
rect -44556 -21686 -44542 -21619
rect -44721 -21689 -44542 -21686
rect -44941 -25352 -44542 -21689
rect -43847 -24018 -43695 -16393
rect -43337 -16972 -43250 -16951
rect -43337 -17028 -43324 -16972
rect -43268 -17028 -43250 -16972
rect -43337 -17083 -43250 -17028
rect -43337 -17139 -43328 -17083
rect -43272 -17139 -43250 -17083
rect -43337 -17154 -43250 -17139
rect -42793 -17910 -42730 -15221
rect -40679 -15848 -40623 -15640
rect -40676 -16302 -40620 -16063
rect -42828 -17973 -42730 -17910
rect -42828 -22630 -42765 -17973
rect -40627 -18648 -40570 -18407
rect -36071 -19466 -35963 -19434
rect -36071 -19561 -36053 -19466
rect -35976 -19561 -35963 -19466
rect -36071 -19642 -35963 -19561
rect -36071 -19737 -36056 -19642
rect -35979 -19737 -35963 -19642
rect -36071 -19801 -35963 -19737
rect -36071 -19896 -36054 -19801
rect -35977 -19896 -35963 -19801
rect -36071 -19959 -35963 -19896
rect -36071 -20054 -36055 -19959
rect -35978 -20054 -35963 -19959
rect -36274 -20487 -36169 -20471
rect -36278 -20513 -36169 -20487
rect -36278 -20608 -36260 -20513
rect -36183 -20608 -36169 -20513
rect -36278 -20689 -36169 -20608
rect -36278 -20784 -36263 -20689
rect -36186 -20784 -36169 -20689
rect -36278 -20848 -36169 -20784
rect -36278 -20943 -36261 -20848
rect -36184 -20943 -36169 -20848
rect -36278 -21006 -36169 -20943
rect -36278 -21101 -36262 -21006
rect -36185 -21101 -36169 -21006
rect -36278 -21124 -36169 -21101
rect -36274 -22036 -36169 -21124
rect -36071 -21957 -35963 -20054
rect -42828 -22693 -42566 -22630
rect -42813 -22989 -42726 -22968
rect -42813 -23045 -42800 -22989
rect -42744 -23045 -42726 -22989
rect -42813 -23100 -42726 -23045
rect -42813 -23156 -42804 -23100
rect -42748 -23156 -42726 -23100
rect -42813 -23171 -42726 -23156
rect -43847 -24082 -43793 -24018
rect -43740 -24082 -43695 -24018
rect -43847 -24200 -43695 -24082
rect -43847 -24264 -43796 -24200
rect -43743 -24264 -43695 -24200
rect -43847 -24432 -43695 -24264
rect -44941 -25354 -44693 -25352
rect -44941 -25360 -44810 -25354
rect -44941 -25416 -44926 -25360
rect -44874 -25410 -44810 -25360
rect -44758 -25408 -44693 -25354
rect -44641 -25408 -44542 -25352
rect -44758 -25410 -44542 -25408
rect -44874 -25416 -44542 -25410
rect -44941 -26968 -44542 -25416
rect -44941 -26969 -44792 -26968
rect -44941 -27047 -44934 -26969
rect -44876 -27046 -44792 -26969
rect -44734 -26971 -44542 -26968
rect -44734 -27046 -44625 -26971
rect -44876 -27047 -44625 -27046
rect -44941 -27049 -44625 -27047
rect -44567 -27049 -44542 -26971
rect -44941 -29752 -44542 -27049
rect -43815 -27798 -43727 -24432
rect -42629 -24973 -42566 -22693
rect -40528 -23736 -40472 -23448
rect -40525 -24215 -40469 -24007
rect -35392 -24179 -34993 -14627
rect -35392 -24235 -35377 -24179
rect -35325 -24180 -34993 -24179
rect -35325 -24181 -35104 -24180
rect -35325 -24235 -35251 -24181
rect -35392 -24237 -35251 -24235
rect -35199 -24236 -35104 -24181
rect -35052 -24236 -34993 -24180
rect -35199 -24237 -34993 -24236
rect -43355 -25037 -43028 -24974
rect -43355 -25050 -43186 -25037
rect -43355 -25117 -43341 -25050
rect -43267 -25104 -43186 -25050
rect -43112 -25104 -43028 -25037
rect -43267 -25117 -43028 -25104
rect -43355 -25126 -43028 -25117
rect -42701 -25023 -42445 -24973
rect -42701 -25027 -42538 -25023
rect -42701 -25098 -42676 -25027
rect -42616 -25094 -42538 -25027
rect -42478 -25094 -42445 -25023
rect -42616 -25098 -42445 -25094
rect -42701 -25126 -42445 -25098
rect -43815 -27856 -43801 -27798
rect -43741 -27856 -43727 -27798
rect -43815 -27936 -43727 -27856
rect -43815 -27994 -43803 -27936
rect -43743 -27994 -43727 -27936
rect -43815 -28009 -43727 -27994
rect -43627 -26282 -43546 -26251
rect -43627 -26338 -43616 -26282
rect -43555 -26338 -43546 -26282
rect -43627 -26406 -43546 -26338
rect -43627 -26462 -43618 -26406
rect -43557 -26462 -43546 -26406
rect -44941 -29756 -44626 -29752
rect -44941 -29827 -44931 -29756
rect -44876 -29757 -44626 -29756
rect -44876 -29827 -44788 -29757
rect -44941 -29828 -44788 -29827
rect -44733 -29823 -44626 -29757
rect -44571 -29823 -44542 -29752
rect -44733 -29828 -44542 -29823
rect -44941 -33447 -44542 -29828
rect -43901 -28172 -43816 -28151
rect -43901 -28233 -43887 -28172
rect -43827 -28233 -43816 -28172
rect -43901 -28337 -43816 -28233
rect -43901 -28398 -43891 -28337
rect -43831 -28398 -43816 -28337
rect -43901 -31669 -43816 -28398
rect -43627 -28475 -43546 -26462
rect -40476 -26559 -40419 -26308
rect -43348 -26824 -42817 -26732
rect -43632 -28498 -43538 -28475
rect -43632 -28564 -43607 -28498
rect -43551 -28564 -43538 -28498
rect -43632 -28651 -43538 -28564
rect -43632 -28717 -43616 -28651
rect -43560 -28717 -43538 -28651
rect -43632 -28736 -43538 -28717
rect -44941 -33450 -44789 -33447
rect -44941 -33513 -44921 -33450
rect -44861 -33510 -44789 -33450
rect -44729 -33450 -44542 -33447
rect -44729 -33510 -44655 -33450
rect -44861 -33513 -44655 -33510
rect -44595 -33513 -44542 -33450
rect -44941 -35006 -44542 -33513
rect -44941 -35077 -44922 -35006
rect -44867 -35010 -44542 -35006
rect -44867 -35077 -44782 -35010
rect -44941 -35081 -44782 -35077
rect -44727 -35021 -44542 -35010
rect -44727 -35081 -44632 -35021
rect -44941 -35092 -44632 -35081
rect -44577 -35092 -44542 -35021
rect -44941 -36500 -44542 -35092
rect -43923 -31995 -43792 -31669
rect -43923 -32051 -43893 -31995
rect -43827 -32051 -43792 -31995
rect -43923 -32154 -43792 -32051
rect -43923 -32210 -43895 -32154
rect -43829 -32210 -43792 -32154
rect -44941 -36517 -44529 -36500
rect -44941 -36520 -44612 -36517
rect -44941 -36525 -44761 -36520
rect -44941 -36620 -44920 -36525
rect -44843 -36615 -44761 -36525
rect -44684 -36612 -44612 -36520
rect -44535 -36612 -44529 -36517
rect -44684 -36615 -44529 -36612
rect -44843 -36620 -44529 -36615
rect -44941 -36693 -44529 -36620
rect -44941 -36696 -44615 -36693
rect -44941 -36701 -44764 -36696
rect -44941 -36796 -44923 -36701
rect -44846 -36791 -44764 -36701
rect -44687 -36788 -44615 -36696
rect -44538 -36788 -44529 -36693
rect -44687 -36791 -44529 -36788
rect -44846 -36796 -44529 -36791
rect -44941 -36852 -44529 -36796
rect -44941 -36855 -44613 -36852
rect -44941 -36860 -44762 -36855
rect -44941 -36955 -44921 -36860
rect -44844 -36950 -44762 -36860
rect -44685 -36947 -44613 -36855
rect -44536 -36947 -44529 -36852
rect -44685 -36950 -44529 -36947
rect -44844 -36955 -44529 -36950
rect -44941 -37010 -44529 -36955
rect -44941 -37013 -44614 -37010
rect -44941 -37018 -44763 -37013
rect -44941 -37113 -44922 -37018
rect -44845 -37108 -44763 -37018
rect -44686 -37105 -44614 -37013
rect -44537 -37105 -44529 -37010
rect -44686 -37108 -44529 -37105
rect -44845 -37113 -44529 -37108
rect -44941 -37125 -44529 -37113
rect -45764 -37556 -45351 -37539
rect -45764 -37559 -45434 -37556
rect -45764 -37564 -45583 -37559
rect -45764 -37659 -45742 -37564
rect -45665 -37654 -45583 -37564
rect -45506 -37651 -45434 -37559
rect -45357 -37651 -45351 -37556
rect -45506 -37654 -45351 -37651
rect -45665 -37659 -45351 -37654
rect -45764 -37732 -45351 -37659
rect -45764 -37735 -45437 -37732
rect -45764 -37740 -45586 -37735
rect -45764 -37835 -45745 -37740
rect -45668 -37830 -45586 -37740
rect -45509 -37827 -45437 -37735
rect -45360 -37827 -45351 -37732
rect -45509 -37830 -45351 -37827
rect -45668 -37835 -45351 -37830
rect -45764 -37891 -45351 -37835
rect -45764 -37894 -45435 -37891
rect -45764 -37899 -45584 -37894
rect -45764 -37994 -45743 -37899
rect -45666 -37989 -45584 -37899
rect -45507 -37986 -45435 -37894
rect -45358 -37986 -45351 -37891
rect -45507 -37989 -45351 -37986
rect -45666 -37994 -45351 -37989
rect -45764 -38049 -45351 -37994
rect -45764 -38052 -45436 -38049
rect -45764 -38057 -45585 -38052
rect -45764 -38152 -45744 -38057
rect -45667 -38147 -45585 -38057
rect -45508 -38144 -45436 -38052
rect -45359 -38144 -45351 -38049
rect -45508 -38147 -45351 -38144
rect -45667 -38152 -45351 -38147
rect -45764 -38164 -45351 -38152
rect -44941 -37948 -44542 -37125
rect -43923 -37267 -43792 -32210
rect -43627 -34255 -43546 -28736
rect -43348 -28870 -43256 -26824
rect -36032 -27509 -35924 -27472
rect -36032 -27604 -36007 -27509
rect -35930 -27604 -35924 -27509
rect -36032 -27685 -35924 -27604
rect -36032 -27780 -36010 -27685
rect -35933 -27780 -35924 -27685
rect -36032 -27844 -35924 -27780
rect -36032 -27939 -36008 -27844
rect -35931 -27939 -35924 -27844
rect -36032 -28002 -35924 -27939
rect -36032 -28097 -36009 -28002
rect -35932 -28097 -35924 -28002
rect -43349 -28920 -43256 -28870
rect -43349 -29004 -43332 -28920
rect -43262 -29004 -43256 -28920
rect -43349 -29076 -43256 -29004
rect -43349 -29160 -43340 -29076
rect -43270 -29160 -43256 -29076
rect -43349 -29170 -43256 -29160
rect -43348 -33832 -43256 -29170
rect -36235 -28551 -36130 -28515
rect -36235 -28646 -36214 -28551
rect -36137 -28646 -36130 -28551
rect -36235 -28727 -36130 -28646
rect -36235 -28822 -36217 -28727
rect -36140 -28822 -36130 -28727
rect -36235 -28886 -36130 -28822
rect -36235 -28981 -36215 -28886
rect -36138 -28981 -36130 -28886
rect -36235 -29044 -36130 -28981
rect -36235 -29139 -36216 -29044
rect -36139 -29139 -36130 -29044
rect -36235 -30047 -36130 -29139
rect -36032 -30024 -35924 -28097
rect -40489 -31737 -40433 -31482
rect -40486 -32322 -40430 -32103
rect -35392 -32467 -34993 -24237
rect -35392 -32470 -35243 -32467
rect -35392 -32533 -35375 -32470
rect -35315 -32530 -35243 -32470
rect -35183 -32470 -34993 -32467
rect -35183 -32530 -35109 -32470
rect -35315 -32533 -35109 -32530
rect -35049 -32533 -34993 -32470
rect -43142 -33085 -42954 -33053
rect -43142 -33088 -43020 -33085
rect -43142 -33147 -43133 -33088
rect -43077 -33144 -43020 -33088
rect -42964 -33144 -42954 -33085
rect -43077 -33147 -42954 -33144
rect -43142 -33176 -42954 -33147
rect -43348 -33924 -42792 -33832
rect -43627 -34308 -43609 -34255
rect -43554 -34308 -43546 -34255
rect -43627 -34381 -43546 -34308
rect -43627 -34434 -43614 -34381
rect -43559 -34434 -43546 -34381
rect -43627 -34450 -43546 -34434
rect -40437 -34658 -40380 -34412
rect -43941 -37312 -43741 -37267
rect -43941 -37313 -43808 -37312
rect -43941 -37411 -43923 -37313
rect -43865 -37410 -43808 -37313
rect -43750 -37410 -43741 -37312
rect -43865 -37411 -43741 -37410
rect -43941 -37443 -43741 -37411
rect -44941 -37953 -44623 -37948
rect -44941 -38051 -44929 -37953
rect -44871 -38051 -44782 -37953
rect -44724 -38046 -44623 -37953
rect -44565 -38046 -44542 -37948
rect -44724 -38051 -44542 -38046
rect -45764 -38313 -45365 -38164
rect -44941 -38313 -44542 -38051
rect -35392 -37543 -34993 -32533
rect -34702 51264 -34303 55223
rect -24190 54809 -23791 55873
rect -23397 55848 -22998 55873
rect -23397 55831 -22984 55848
rect -23397 55828 -23067 55831
rect -23397 55823 -23216 55828
rect -23397 55728 -23375 55823
rect -23298 55733 -23216 55823
rect -23139 55736 -23067 55828
rect -22990 55736 -22984 55831
rect -23139 55733 -22984 55736
rect -23298 55728 -22984 55733
rect -23397 55655 -22984 55728
rect -23397 55652 -23070 55655
rect -23397 55647 -23219 55652
rect -23397 55552 -23378 55647
rect -23301 55557 -23219 55647
rect -23142 55560 -23070 55652
rect -22993 55560 -22984 55655
rect -23142 55557 -22984 55560
rect -23301 55552 -22984 55557
rect -23397 55496 -22984 55552
rect -23397 55493 -23068 55496
rect -23397 55488 -23217 55493
rect -23397 55393 -23376 55488
rect -23299 55398 -23217 55488
rect -23140 55401 -23068 55493
rect -22991 55401 -22984 55496
rect -23140 55398 -22984 55401
rect -23299 55393 -22984 55398
rect -23397 55338 -22984 55393
rect -23397 55335 -23069 55338
rect -23397 55330 -23218 55335
rect -23397 55235 -23377 55330
rect -23300 55240 -23218 55330
rect -23141 55243 -23069 55335
rect -22992 55243 -22984 55338
rect -23141 55240 -22984 55243
rect -23300 55235 -22984 55240
rect -23397 55223 -22984 55235
rect -24190 54792 -23779 54809
rect -24190 54789 -23862 54792
rect -24190 54784 -24011 54789
rect -24190 54689 -24170 54784
rect -24093 54694 -24011 54784
rect -23934 54697 -23862 54789
rect -23785 54697 -23779 54792
rect -23934 54694 -23779 54697
rect -24093 54689 -23779 54694
rect -24190 54616 -23779 54689
rect -24190 54613 -23865 54616
rect -24190 54608 -24014 54613
rect -24190 54513 -24173 54608
rect -24096 54518 -24014 54608
rect -23937 54521 -23865 54613
rect -23788 54521 -23779 54616
rect -23937 54518 -23779 54521
rect -24096 54513 -23779 54518
rect -24190 54457 -23779 54513
rect -24190 54454 -23863 54457
rect -24190 54449 -24012 54454
rect -24190 54354 -24171 54449
rect -24094 54359 -24012 54449
rect -23935 54362 -23863 54454
rect -23786 54362 -23779 54457
rect -23935 54359 -23779 54362
rect -24094 54354 -23779 54359
rect -24190 54299 -23779 54354
rect -24190 54296 -23864 54299
rect -24190 54291 -24013 54296
rect -24190 54196 -24172 54291
rect -24095 54201 -24013 54291
rect -23936 54204 -23864 54296
rect -23787 54204 -23779 54299
rect -23936 54201 -23779 54204
rect -24095 54196 -23779 54201
rect -24190 54184 -23779 54196
rect -32412 52416 -32065 52431
rect -32412 52342 -32393 52416
rect -32319 52342 -32152 52416
rect -32078 52342 -32065 52416
rect -32412 52331 -32065 52342
rect -32652 52166 -32293 52180
rect -32652 52066 -32642 52166
rect -32542 52066 -32415 52166
rect -32315 52066 -32293 52166
rect -32652 52052 -32293 52066
rect -34702 51261 -34395 51264
rect -34702 51258 -34546 51261
rect -34702 51187 -34692 51258
rect -34618 51190 -34546 51258
rect -34472 51193 -34395 51261
rect -34321 51193 -34303 51264
rect -34472 51190 -34303 51193
rect -34618 51187 -34303 51190
rect -32415 51188 -32315 52052
rect -32152 51825 -32078 52331
rect -32166 51817 -32065 51825
rect -32166 51743 -32152 51817
rect -32078 51743 -32065 51817
rect -32166 51643 -32065 51743
rect -32166 51571 -32151 51643
rect -32079 51571 -32065 51643
rect -32166 51556 -32065 51571
rect -34702 46337 -34303 51187
rect -32439 51168 -32291 51188
rect -32439 51057 -32421 51168
rect -32310 51057 -32291 51168
rect -32439 50942 -32291 51057
rect -32439 50833 -32421 50942
rect -32312 50833 -32291 50942
rect -32439 50815 -32291 50833
rect -24190 50312 -23791 54184
rect -24190 50309 -24037 50312
rect -24190 50246 -24169 50309
rect -24109 50249 -24037 50309
rect -23977 50309 -23791 50312
rect -23977 50249 -23903 50309
rect -24109 50246 -23903 50249
rect -23843 50246 -23791 50309
rect -32518 50028 -32331 50077
rect -32518 49929 -32478 50028
rect -32359 49929 -32331 50028
rect -32518 49806 -32331 49929
rect -32518 49707 -32484 49806
rect -32365 49707 -32331 49806
rect -32518 49685 -32331 49707
rect -34702 46334 -34550 46337
rect -34702 46271 -34682 46334
rect -34622 46274 -34550 46334
rect -34490 46334 -34303 46337
rect -34490 46274 -34416 46334
rect -34622 46271 -34416 46274
rect -34356 46271 -34303 46334
rect -34702 43097 -34303 46271
rect -34702 43093 -34392 43097
rect -34702 43092 -34537 43093
rect -34702 43015 -34690 43092
rect -34620 43016 -34537 43092
rect -34467 43020 -34392 43093
rect -34322 43020 -34303 43097
rect -34467 43016 -34303 43020
rect -34620 43015 -34303 43016
rect -34702 39467 -34303 43015
rect -34702 39464 -34393 39467
rect -34702 39387 -34694 39464
rect -34624 39387 -34544 39464
rect -34474 39390 -34393 39464
rect -34323 39390 -34303 39467
rect -34474 39387 -34303 39390
rect -34702 38133 -34303 39387
rect -34702 38131 -34405 38133
rect -34702 38125 -34538 38131
rect -34702 38069 -34669 38125
rect -34617 38075 -34538 38125
rect -34486 38077 -34405 38131
rect -34353 38077 -34303 38133
rect -34486 38075 -34303 38077
rect -34617 38069 -34303 38075
rect -34702 34573 -34303 38069
rect -34702 34572 -34545 34573
rect -34702 34483 -34693 34572
rect -34623 34484 -34545 34572
rect -34475 34572 -34303 34573
rect -34475 34484 -34401 34572
rect -34623 34483 -34401 34484
rect -34331 34483 -34303 34572
rect -34702 30708 -34303 34483
rect -34702 30698 -34550 30708
rect -34702 30615 -34681 30698
rect -34611 30625 -34550 30698
rect -34480 30706 -34303 30708
rect -34480 30625 -34422 30706
rect -34611 30623 -34422 30625
rect -34352 30623 -34303 30706
rect -34611 30615 -34303 30623
rect -34702 26140 -34303 30615
rect -34702 26138 -34391 26140
rect -34702 26063 -34687 26138
rect -34625 26135 -34391 26138
rect -34625 26063 -34553 26135
rect -34702 26060 -34553 26063
rect -34491 26065 -34391 26135
rect -34329 26065 -34303 26140
rect -34491 26060 -34303 26065
rect -34702 20831 -34303 26060
rect -34702 20827 -34399 20831
rect -34702 20824 -34543 20827
rect -34702 20762 -34682 20824
rect -34623 20765 -34543 20824
rect -34484 20769 -34399 20827
rect -34340 20769 -34303 20831
rect -34484 20765 -34303 20769
rect -34623 20762 -34303 20765
rect -34702 16970 -34303 20762
rect -34702 16969 -34391 16970
rect -34702 16892 -34687 16969
rect -34625 16968 -34391 16969
rect -34625 16892 -34540 16968
rect -34702 16891 -34540 16892
rect -34478 16893 -34391 16968
rect -34329 16893 -34303 16970
rect -34478 16891 -34303 16893
rect -34702 13448 -34303 16891
rect -34702 13447 -34400 13448
rect -34702 13394 -34685 13447
rect -34630 13446 -34400 13447
rect -34630 13394 -34546 13446
rect -34702 13393 -34546 13394
rect -34491 13395 -34400 13446
rect -34345 13395 -34303 13448
rect -34491 13393 -34303 13395
rect -34702 11709 -34303 13393
rect -34022 44672 -33847 44719
rect -34022 44612 -33957 44672
rect -33884 44612 -33847 44672
rect -34022 44527 -33847 44612
rect -34022 44467 -33959 44527
rect -33886 44467 -33847 44527
rect -34022 34871 -33847 44467
rect -32491 41790 -32377 49685
rect -30741 49098 -30685 49257
rect -31355 47850 -31299 48021
rect -30291 46819 -30235 47020
rect -31939 46704 -31692 46726
rect -31939 46703 -31785 46704
rect -31939 46648 -31908 46703
rect -31853 46648 -31785 46703
rect -31939 46647 -31785 46648
rect -31728 46647 -31692 46704
rect -31939 46615 -31692 46647
rect -31939 44429 -31828 46615
rect -31579 45977 -30892 46088
rect -31938 44415 -31836 44429
rect -31938 44345 -31905 44415
rect -31844 44345 -31836 44415
rect -31938 44236 -31836 44345
rect -31938 44166 -31915 44236
rect -31854 44166 -31836 44236
rect -31938 44153 -31836 44166
rect -31579 43941 -31468 45977
rect -30945 43996 -30827 44015
rect -31602 43906 -31461 43941
rect -30945 43913 -30930 43996
rect -30847 43913 -30827 43996
rect -31602 43797 -31577 43906
rect -31468 43797 -31459 43906
rect -30945 43817 -30827 43913
rect -31602 43692 -31461 43797
rect -30945 43736 -30928 43817
rect -30847 43736 -30827 43817
rect -30945 43721 -30827 43736
rect -31602 43581 -31579 43692
rect -31468 43581 -31461 43692
rect -31602 43551 -31461 43581
rect -31579 42901 -31468 43551
rect -30930 43293 -30847 43721
rect -30917 43196 -30861 43293
rect -31592 42863 -31451 42901
rect -31592 42752 -31579 42863
rect -31470 42752 -31451 42863
rect -31592 42625 -31451 42752
rect -31592 42514 -31580 42625
rect -31469 42514 -31451 42625
rect -31592 42511 -31451 42514
rect -24190 42016 -23791 50246
rect -24190 42003 -24043 42016
rect -24190 41947 -24173 42003
rect -24121 41960 -24043 42003
rect -23991 42003 -23791 42016
rect -23991 41960 -23920 42003
rect -24121 41947 -23920 41960
rect -23868 41947 -23791 42003
rect -32499 41759 -32337 41790
rect -32499 41675 -32467 41759
rect -32362 41685 -32337 41759
rect -32362 41675 -32213 41685
rect -32499 41568 -32213 41675
rect -32499 41484 -32472 41568
rect -32367 41484 -32213 41568
rect -32499 41461 -32213 41484
rect -32391 41453 -32213 41461
rect -33727 38498 -33509 38514
rect -33727 38443 -33700 38498
rect -33645 38443 -33574 38498
rect -33519 38443 -33509 38498
rect -33727 38403 -33509 38443
rect -34022 34817 -33992 34871
rect -33863 34817 -33847 34871
rect -34022 34758 -33847 34817
rect -34022 34704 -33993 34758
rect -33864 34704 -33847 34758
rect -34022 34650 -33847 34704
rect -34022 34596 -33992 34650
rect -33863 34596 -33847 34650
rect -34022 34539 -33847 34596
rect -34022 34485 -33999 34539
rect -33870 34485 -33847 34539
rect -34022 32194 -33847 34485
rect -34022 32128 -34001 32194
rect -33863 32128 -33847 32194
rect -34022 32011 -33847 32128
rect -34022 31945 -34006 32011
rect -33868 31945 -33847 32011
rect -34022 31862 -33847 31945
rect -34022 31796 -34008 31862
rect -33870 31796 -33847 31862
rect -34022 14830 -33847 31796
rect -34022 14760 -33934 14830
rect -33866 14760 -33847 14830
rect -34022 14654 -33847 14760
rect -34022 14584 -33934 14654
rect -33866 14584 -33847 14654
rect -34022 12237 -33847 14584
rect -33718 26152 -33607 38403
rect -33323 37850 -33091 37863
rect -33323 37845 -33157 37850
rect -33323 37788 -33290 37845
rect -33230 37793 -33157 37845
rect -33097 37793 -33091 37850
rect -33230 37788 -33091 37793
rect -33323 37752 -33091 37788
rect -33718 26134 -33408 26152
rect -33718 26133 -33502 26134
rect -33718 26061 -33703 26133
rect -33631 26061 -33502 26133
rect -33718 26060 -33502 26061
rect -33428 26060 -33408 26134
rect -33718 26045 -33408 26060
rect -33718 20650 -33607 26045
rect -33718 20590 -33690 20650
rect -33630 20590 -33607 20650
rect -33718 20510 -33607 20590
rect -33718 20450 -33690 20510
rect -33630 20450 -33607 20510
rect -33718 12575 -33607 20450
rect -33253 23988 -33142 37752
rect -32327 31139 -32213 41453
rect -30657 40897 -30601 41053
rect -31271 39660 -31215 39829
rect -30207 38644 -30151 38818
rect -24978 37020 -24870 37072
rect -24978 36925 -24963 37020
rect -24886 36925 -24870 37020
rect -24978 36844 -24870 36925
rect -24978 36749 -24966 36844
rect -24889 36749 -24870 36844
rect -24978 36685 -24870 36749
rect -24978 36590 -24964 36685
rect -24887 36590 -24870 36685
rect -24978 36527 -24870 36590
rect -24978 36432 -24965 36527
rect -24888 36432 -24870 36527
rect -25181 35760 -25076 35814
rect -25181 35665 -25161 35760
rect -25084 35665 -25076 35760
rect -25181 35584 -25076 35665
rect -25181 35489 -25164 35584
rect -25087 35489 -25076 35584
rect -25181 35425 -25076 35489
rect -25181 35330 -25162 35425
rect -25085 35330 -25076 35425
rect -25181 35267 -25076 35330
rect -25181 35172 -25163 35267
rect -25086 35172 -25076 35267
rect -25181 34065 -25076 35172
rect -24978 33854 -24870 36432
rect -24190 33501 -23791 41947
rect -24190 33497 -23912 33501
rect -24190 33495 -24038 33497
rect -24190 33412 -24174 33495
rect -24104 33414 -24038 33495
rect -23968 33418 -23912 33497
rect -23842 33418 -23791 33501
rect -23968 33414 -23791 33418
rect -24104 33412 -23791 33414
rect -31751 33108 -31628 33122
rect -31751 33029 -31731 33108
rect -31640 33029 -31628 33108
rect -31751 32956 -31628 33029
rect -31751 32877 -31735 32956
rect -31644 32877 -31628 32956
rect -31751 32865 -31628 32877
rect -29435 32551 -29379 32697
rect -29432 31807 -29376 32038
rect -32055 31139 -31932 31148
rect -32327 31134 -31932 31139
rect -32327 31055 -32035 31134
rect -31944 31055 -31932 31134
rect -32327 31025 -31932 31055
rect -32055 30982 -31932 31025
rect -32055 30903 -32039 30982
rect -31948 30903 -31932 30982
rect -32055 30891 -31932 30903
rect -32322 29776 -31960 29809
rect -32322 29770 -32106 29776
rect -32322 29704 -32283 29770
rect -32222 29710 -32106 29770
rect -32045 29710 -31960 29776
rect -32222 29704 -31960 29710
rect -32322 29670 -31960 29704
rect -32199 28792 -32089 29670
rect -29383 29503 -29326 29708
rect -32436 28778 -32074 28792
rect -32436 28777 -32207 28778
rect -32436 28667 -32427 28777
rect -32317 28667 -32207 28777
rect -32436 28666 -32207 28667
rect -32095 28666 -32074 28778
rect -32436 28653 -32074 28666
rect -24190 25270 -23791 33412
rect -23397 51273 -22998 55223
rect -11229 53602 -11121 53640
rect -11229 53507 -11204 53602
rect -11127 53507 -11121 53602
rect -11229 53426 -11121 53507
rect -11229 53331 -11207 53426
rect -11130 53331 -11121 53426
rect -11229 53267 -11121 53331
rect -11229 53172 -11205 53267
rect -11128 53172 -11121 53267
rect -11229 53109 -11121 53172
rect -11229 53014 -11206 53109
rect -11129 53014 -11121 53109
rect -11432 52556 -11327 52598
rect -11432 52461 -11417 52556
rect -11340 52461 -11327 52556
rect -18447 52423 -18336 52439
rect -18447 52336 -18434 52423
rect -18347 52336 -18336 52423
rect -18447 52221 -18336 52336
rect -18790 52165 -18663 52181
rect -18790 52067 -18775 52165
rect -18677 52067 -18663 52165
rect -18447 52132 -18434 52221
rect -18345 52132 -18336 52221
rect -18447 52117 -18336 52132
rect -11432 52380 -11327 52461
rect -11432 52285 -11420 52380
rect -11343 52285 -11327 52380
rect -11432 52221 -11327 52285
rect -11432 52126 -11418 52221
rect -11341 52126 -11327 52221
rect -18790 51928 -18663 52067
rect -18790 51828 -18776 51928
rect -18676 51828 -18663 51928
rect -18790 51814 -18663 51828
rect -23397 51271 -23234 51273
rect -23397 51196 -23385 51271
rect -23314 51198 -23234 51271
rect -23163 51272 -22998 51273
rect -23163 51198 -23089 51272
rect -23314 51197 -23089 51198
rect -23018 51197 -22998 51272
rect -23314 51196 -22998 51197
rect -23397 47933 -22998 51196
rect -23397 47930 -23249 47933
rect -23397 47867 -23381 47930
rect -23321 47870 -23249 47930
rect -23189 47930 -22998 47933
rect -23189 47870 -23115 47930
rect -23321 47867 -23115 47870
rect -23055 47867 -22998 47930
rect -23397 47561 -22998 47867
rect -23397 47558 -23251 47561
rect -23397 47495 -23383 47558
rect -23323 47498 -23251 47558
rect -23191 47558 -22998 47561
rect -23191 47498 -23117 47558
rect -23323 47495 -23117 47498
rect -23057 47495 -22998 47558
rect -23397 46342 -22998 47495
rect -23397 46265 -23383 46342
rect -23320 46341 -22998 46342
rect -23320 46265 -23240 46341
rect -23397 46264 -23240 46265
rect -23177 46264 -23101 46341
rect -23038 46264 -22998 46341
rect -23397 43078 -22998 46264
rect -19394 48853 -19274 48918
rect -19394 48785 -19370 48853
rect -19289 48785 -19274 48853
rect -19394 48713 -19274 48785
rect -19394 48645 -19377 48713
rect -19296 48645 -19274 48713
rect -19394 44610 -19274 48645
rect -18775 47226 -18675 51814
rect -18993 47188 -18665 47226
rect -18993 47187 -18775 47188
rect -18993 47089 -18960 47187
rect -18862 47089 -18775 47187
rect -18993 47088 -18775 47089
rect -18675 47088 -18665 47188
rect -18993 47053 -18665 47088
rect -18434 46668 -18345 52117
rect -11432 52063 -11327 52126
rect -11432 51968 -11419 52063
rect -11342 51968 -11327 52063
rect -11432 50908 -11327 51968
rect -11229 50970 -11121 53014
rect -17998 49967 -17875 49981
rect -17998 49888 -17978 49967
rect -17887 49888 -17875 49967
rect -17998 49815 -17875 49888
rect -15683 49886 -15088 49942
rect -17998 49736 -17982 49815
rect -17891 49736 -17875 49815
rect -17998 49724 -17875 49736
rect -15686 49432 -15630 49745
rect -15683 48865 -15682 48918
rect -15628 48865 -15627 48918
rect -15683 48703 -15627 48865
rect -8574 48139 -8343 56567
rect -7915 54813 -7516 55873
rect -7146 55849 -6747 55873
rect -7146 55832 -6735 55849
rect -7146 55829 -6818 55832
rect -7146 55824 -6967 55829
rect -7146 55729 -7126 55824
rect -7049 55734 -6967 55824
rect -6890 55737 -6818 55829
rect -6741 55737 -6735 55832
rect -6890 55734 -6735 55737
rect -7049 55729 -6735 55734
rect -7146 55656 -6735 55729
rect -7146 55653 -6821 55656
rect -7146 55648 -6970 55653
rect -7146 55553 -7129 55648
rect -7052 55558 -6970 55648
rect -6893 55561 -6821 55653
rect -6744 55561 -6735 55656
rect -6893 55558 -6735 55561
rect -7052 55553 -6735 55558
rect -7146 55497 -6735 55553
rect -7146 55494 -6819 55497
rect -7146 55489 -6968 55494
rect -7146 55394 -7127 55489
rect -7050 55399 -6968 55489
rect -6891 55402 -6819 55494
rect -6742 55402 -6735 55497
rect -6891 55399 -6735 55402
rect -7050 55394 -6735 55399
rect -7146 55339 -6735 55394
rect -7146 55336 -6820 55339
rect -7146 55331 -6969 55336
rect -7146 55236 -7128 55331
rect -7051 55241 -6969 55331
rect -6892 55244 -6820 55336
rect -6743 55244 -6735 55339
rect -6892 55241 -6735 55244
rect -7051 55236 -6735 55241
rect -7146 55224 -6735 55236
rect -7918 54796 -7508 54813
rect -7918 54793 -7591 54796
rect -7918 54788 -7740 54793
rect -7918 54693 -7899 54788
rect -7822 54698 -7740 54788
rect -7663 54701 -7591 54793
rect -7514 54701 -7508 54796
rect -7663 54698 -7508 54701
rect -7822 54693 -7508 54698
rect -7918 54620 -7508 54693
rect -7918 54617 -7594 54620
rect -7918 54612 -7743 54617
rect -7918 54517 -7902 54612
rect -7825 54522 -7743 54612
rect -7666 54525 -7594 54617
rect -7517 54525 -7508 54620
rect -7666 54522 -7508 54525
rect -7825 54517 -7508 54522
rect -7918 54461 -7508 54517
rect -7918 54458 -7592 54461
rect -7918 54453 -7741 54458
rect -7918 54358 -7900 54453
rect -7823 54363 -7741 54453
rect -7664 54366 -7592 54458
rect -7515 54366 -7508 54461
rect -7664 54363 -7508 54366
rect -7823 54358 -7508 54363
rect -7918 54303 -7508 54358
rect -7918 54300 -7593 54303
rect -7918 54295 -7742 54300
rect -7918 54200 -7901 54295
rect -7824 54205 -7742 54295
rect -7665 54208 -7593 54300
rect -7516 54208 -7508 54303
rect -7665 54205 -7508 54208
rect -7824 54200 -7508 54205
rect -7918 54188 -7508 54200
rect -8574 48136 -8419 48139
rect -8574 48039 -8564 48136
rect -8508 48042 -8419 48136
rect -8363 48042 -8343 48139
rect -8508 48039 -8343 48042
rect -8574 48021 -8343 48039
rect -7915 50365 -7516 54188
rect -7915 50362 -7751 50365
rect -7915 50299 -7883 50362
rect -7823 50302 -7751 50362
rect -7691 50362 -7516 50365
rect -7691 50302 -7617 50362
rect -7823 50299 -7617 50302
rect -7557 50299 -7516 50362
rect -7915 47700 -7516 50299
rect -7915 47697 -7741 47700
rect -7915 47634 -7873 47697
rect -7813 47637 -7741 47697
rect -7681 47697 -7516 47700
rect -7681 47637 -7607 47697
rect -7813 47634 -7607 47637
rect -7547 47634 -7516 47697
rect -8615 47442 -8384 47459
rect -8615 47388 -8599 47442
rect -8546 47440 -8384 47442
rect -8546 47388 -8468 47440
rect -8615 47386 -8468 47388
rect -8415 47386 -8384 47440
rect -8615 47300 -8384 47386
rect -8615 47298 -8464 47300
rect -8615 47244 -8594 47298
rect -8541 47246 -8464 47298
rect -8411 47246 -8384 47300
rect -8541 47244 -8384 47246
rect -18454 46645 -18175 46668
rect -18454 46556 -18434 46645
rect -18345 46644 -18175 46645
rect -18345 46557 -18276 46644
rect -18189 46557 -18175 46644
rect -18345 46556 -18175 46557
rect -18454 46540 -18175 46556
rect -8615 46416 -8384 47244
rect -9364 46185 -8384 46416
rect -19394 44543 -19373 44610
rect -19296 44543 -19274 44610
rect -19394 44449 -19274 44543
rect -19394 44382 -19373 44449
rect -19296 44382 -19274 44449
rect -19394 44356 -19274 44382
rect -11052 45231 -10944 45275
rect -11052 45136 -11035 45231
rect -10958 45136 -10944 45231
rect -11052 45055 -10944 45136
rect -11052 44960 -11038 45055
rect -10961 44960 -10944 45055
rect -11052 44896 -10944 44960
rect -11052 44801 -11036 44896
rect -10959 44801 -10944 44896
rect -11052 44738 -10944 44801
rect -11052 44643 -11037 44738
rect -10960 44643 -10944 44738
rect -11255 44188 -11150 44241
rect -18983 44132 -18856 44155
rect -18983 44043 -18962 44132
rect -18880 44043 -18856 44132
rect -18983 43890 -18856 44043
rect -18983 43806 -18963 43890
rect -18879 43806 -18856 43890
rect -18983 43792 -18856 43806
rect -11255 44093 -11241 44188
rect -11164 44093 -11150 44188
rect -11255 44012 -11150 44093
rect -11255 43917 -11244 44012
rect -11167 43917 -11150 44012
rect -11255 43853 -11150 43917
rect -23397 43076 -23244 43078
rect -23397 42994 -23387 43076
rect -23321 42996 -23244 43076
rect -23178 43076 -22998 43078
rect -23178 42996 -23090 43076
rect -23321 42994 -23090 42996
rect -23024 42994 -22998 43076
rect -23397 39613 -22998 42994
rect -23397 39607 -23244 39613
rect -23397 39551 -23377 39607
rect -23325 39557 -23244 39607
rect -23192 39557 -23108 39613
rect -23056 39557 -22998 39613
rect -23325 39551 -22998 39557
rect -23397 39245 -22998 39551
rect -23397 39239 -23243 39245
rect -23397 39183 -23376 39239
rect -23324 39189 -23243 39239
rect -23191 39189 -23107 39245
rect -23055 39189 -22998 39245
rect -23324 39183 -22998 39189
rect -23397 34379 -22998 39183
rect -23397 34301 -23382 34379
rect -23321 34378 -22998 34379
rect -23321 34301 -23242 34378
rect -23397 34300 -23242 34301
rect -23181 34377 -22998 34378
rect -23181 34300 -23081 34377
rect -23397 34299 -23081 34300
rect -23020 34299 -22998 34377
rect -23397 32310 -22998 34299
rect -23400 32140 -22998 32310
rect -24190 25180 -24150 25270
rect -24060 25186 -23920 25270
rect -23829 25186 -23791 25270
rect -24060 25180 -23791 25186
rect -32970 24003 -32599 24028
rect -33253 23986 -33141 23988
rect -32970 23986 -32950 24003
rect -33253 23892 -32950 23986
rect -32839 24002 -32599 24003
rect -32839 23893 -32723 24002
rect -32614 23893 -32599 24002
rect -32839 23892 -32599 23893
rect -33253 23875 -32599 23892
rect -33253 20530 -33142 23875
rect -32970 23872 -32599 23875
rect -31493 23601 -31437 23755
rect -32107 22432 -32051 22527
rect -31043 21309 -30987 21500
rect -32636 21201 -32400 21211
rect -32636 21148 -32602 21201
rect -32550 21194 -32400 21201
rect -32550 21148 -32487 21194
rect -32636 21141 -32487 21148
rect -32435 21141 -32400 21194
rect -32636 21120 -32400 21141
rect -33253 20470 -33230 20530
rect -33170 20470 -33142 20530
rect -33253 20410 -33142 20470
rect -33253 20350 -33230 20410
rect -33170 20350 -33142 20410
rect -33253 13095 -33142 20350
rect -32620 20243 -32564 21120
rect -32642 20231 -32358 20243
rect -32642 20228 -32446 20231
rect -32642 20175 -32610 20228
rect -32558 20178 -32446 20228
rect -32394 20178 -32358 20231
rect -32558 20175 -32358 20178
rect -32642 20085 -32358 20175
rect -25847 19413 -25739 19454
rect -25847 19318 -25823 19413
rect -25746 19318 -25739 19413
rect -25847 19237 -25739 19318
rect -25847 19142 -25826 19237
rect -25749 19142 -25739 19237
rect -25847 19078 -25739 19142
rect -25847 18983 -25824 19078
rect -25747 18983 -25739 19078
rect -25847 18920 -25739 18983
rect -25847 18825 -25825 18920
rect -25748 18825 -25739 18920
rect -26050 18326 -25945 18371
rect -26050 18231 -26029 18326
rect -25952 18231 -25945 18326
rect -26050 18150 -25945 18231
rect -26050 18055 -26032 18150
rect -25955 18055 -25945 18150
rect -26050 17991 -25945 18055
rect -26050 17896 -26030 17991
rect -25953 17896 -25945 17991
rect -26050 17833 -25945 17896
rect -26050 17738 -26031 17833
rect -25954 17738 -25945 17833
rect -26050 16823 -25945 17738
rect -25847 16793 -25739 18825
rect -32606 15760 -32519 15781
rect -32606 15704 -32593 15760
rect -32537 15704 -32519 15760
rect -32606 15649 -32519 15704
rect -32606 15593 -32597 15649
rect -32541 15593 -32519 15649
rect -32606 15578 -32519 15593
rect -30304 15113 -30248 15269
rect -30301 14579 -30245 14822
rect -24190 14096 -23791 25180
rect -24190 14094 -23950 14096
rect -24190 14008 -24175 14094
rect -24069 14010 -23950 14094
rect -23844 14010 -23791 14096
rect -24069 14008 -23791 14010
rect -32944 13852 -32857 13873
rect -32944 13796 -32931 13852
rect -32875 13796 -32857 13852
rect -32944 13741 -32857 13796
rect -32944 13685 -32935 13741
rect -32879 13685 -32857 13741
rect -32944 13670 -32857 13685
rect -33253 12984 -32605 13095
rect -33735 12549 -33276 12575
rect -33735 12438 -33718 12549
rect -33607 12438 -33410 12549
rect -33299 12438 -33276 12549
rect -33735 12420 -33276 12438
rect -30252 12241 -30195 12490
rect -34022 12090 -33799 12237
rect -34702 11705 -34416 11709
rect -34702 11614 -34688 11705
rect -34621 11614 -34545 11705
rect -34478 11618 -34416 11705
rect -34349 11618 -34303 11709
rect -34478 11614 -34303 11618
rect -34702 9695 -34303 11614
rect -34702 9692 -34560 9695
rect -34702 9639 -34690 9692
rect -34635 9642 -34560 9692
rect -34505 9693 -34303 9695
rect -34505 9642 -34411 9693
rect -34635 9640 -34411 9642
rect -34356 9640 -34303 9693
rect -34635 9639 -34303 9640
rect -34702 8804 -34303 9639
rect -34702 8800 -34542 8804
rect -34702 8747 -34687 8800
rect -34632 8751 -34542 8800
rect -34487 8802 -34303 8804
rect -34487 8751 -34412 8802
rect -34632 8749 -34412 8751
rect -34357 8749 -34303 8802
rect -34632 8747 -34303 8749
rect -34702 7858 -34303 8747
rect -34702 7857 -34544 7858
rect -34702 7804 -34683 7857
rect -34628 7805 -34544 7857
rect -34489 7805 -34398 7858
rect -34343 7805 -34303 7858
rect -34628 7804 -34303 7805
rect -34702 6991 -34303 7804
rect -34702 6985 -34416 6991
rect -34702 6984 -34552 6985
rect -34702 6931 -34685 6984
rect -34630 6932 -34552 6984
rect -34497 6938 -34416 6985
rect -34361 6938 -34303 6991
rect -34497 6932 -34303 6938
rect -34630 6931 -34303 6932
rect -34702 6075 -34303 6931
rect -34702 6073 -34403 6075
rect -34702 6070 -34545 6073
rect -34702 6017 -34686 6070
rect -34631 6020 -34545 6070
rect -34490 6022 -34403 6073
rect -34348 6022 -34303 6075
rect -34490 6020 -34303 6022
rect -34631 6017 -34303 6020
rect -34702 5160 -34303 6017
rect -34702 5159 -34400 5160
rect -34702 5158 -34551 5159
rect -34702 5105 -34679 5158
rect -34624 5106 -34551 5158
rect -34496 5107 -34400 5159
rect -34345 5107 -34303 5160
rect -34496 5106 -34303 5107
rect -34624 5105 -34303 5106
rect -34702 4167 -34303 5105
rect -34702 4165 -34392 4167
rect -34702 4077 -34680 4165
rect -34610 4161 -34392 4165
rect -34610 4077 -34544 4161
rect -34702 4073 -34544 4077
rect -34474 4079 -34392 4161
rect -34322 4079 -34303 4167
rect -34474 4073 -34303 4079
rect -34702 3984 -34303 4073
rect -34702 3977 -34528 3984
rect -34702 3889 -34685 3977
rect -34615 3896 -34528 3977
rect -34458 3896 -34388 3984
rect -34318 3896 -34303 3984
rect -34615 3889 -34303 3896
rect -34702 531 -34303 3889
rect -33993 2041 -33799 12090
rect -24190 7832 -23791 14008
rect -24190 7738 -24167 7832
rect -24080 7738 -23917 7832
rect -23830 7738 -23791 7832
rect -27113 7389 -27005 7430
rect -27113 7294 -27090 7389
rect -27013 7294 -27005 7389
rect -27113 7213 -27005 7294
rect -27113 7118 -27093 7213
rect -27016 7118 -27005 7213
rect -27113 7054 -27005 7118
rect -27113 6959 -27091 7054
rect -27014 6959 -27005 7054
rect -27113 6896 -27005 6959
rect -27113 6801 -27092 6896
rect -27015 6801 -27005 6896
rect -27937 6161 -27832 6210
rect -27937 6066 -27916 6161
rect -27839 6066 -27832 6161
rect -27937 5985 -27832 6066
rect -27937 5890 -27919 5985
rect -27842 5890 -27832 5985
rect -27937 5826 -27832 5890
rect -27937 5731 -27917 5826
rect -27840 5731 -27832 5826
rect -27937 5668 -27832 5731
rect -27937 5573 -27918 5668
rect -27841 5573 -27832 5668
rect -27937 4713 -27832 5573
rect -27113 5173 -27005 6801
rect -27113 5065 -25631 5173
rect -27937 4608 -25837 4713
rect -25942 3961 -25837 4608
rect -25739 3960 -25631 5065
rect -32487 2818 -32400 2839
rect -32487 2762 -32474 2818
rect -32418 2762 -32400 2818
rect -32487 2707 -32400 2762
rect -32487 2651 -32478 2707
rect -32422 2651 -32400 2707
rect -32487 2636 -32400 2651
rect -24190 2746 -23791 7738
rect -24190 2742 -23866 2746
rect -24190 2736 -24005 2742
rect -24190 2659 -24146 2736
rect -24088 2665 -24005 2736
rect -23947 2669 -23866 2742
rect -23808 2669 -23791 2746
rect -23947 2665 -23791 2669
rect -24088 2659 -23791 2665
rect -24190 2568 -23791 2659
rect -24190 2561 -24014 2568
rect -24190 2484 -24173 2561
rect -24115 2491 -24014 2561
rect -23956 2566 -23791 2568
rect -23956 2491 -23870 2566
rect -24115 2489 -23870 2491
rect -23812 2489 -23791 2566
rect -24115 2484 -23791 2489
rect -30196 2135 -30140 2369
rect -33993 1971 -33928 2041
rect -33868 1971 -33799 2041
rect -33993 1878 -33799 1971
rect -33993 1808 -33928 1878
rect -33868 1808 -33799 1878
rect -33993 1759 -33799 1808
rect -30193 1668 -30137 1910
rect -32846 967 -32759 988
rect -32846 911 -32833 967
rect -32777 911 -32759 967
rect -32846 856 -32759 911
rect -32846 800 -32837 856
rect -32781 800 -32759 856
rect -32846 785 -32759 800
rect -34702 528 -34398 531
rect -34702 527 -34529 528
rect -34702 474 -34686 527
rect -34632 475 -34529 527
rect -34475 478 -34398 528
rect -34344 478 -34303 531
rect -34475 475 -34303 478
rect -34632 474 -34303 475
rect -34702 -1171 -34303 474
rect -33203 -361 -32800 -342
rect -34702 -1181 -34391 -1171
rect -34702 -1281 -34687 -1181
rect -34614 -1183 -34391 -1181
rect -34614 -1281 -34536 -1183
rect -34702 -1283 -34536 -1281
rect -34463 -1271 -34391 -1183
rect -34318 -1271 -34303 -1171
rect -34463 -1283 -34303 -1271
rect -34702 -5123 -34303 -1283
rect -34702 -5126 -34531 -5123
rect -34702 -5193 -34685 -5126
rect -34621 -5190 -34531 -5126
rect -34467 -5125 -34303 -5123
rect -34467 -5190 -34397 -5125
rect -34621 -5192 -34397 -5190
rect -34333 -5192 -34303 -5125
rect -34621 -5193 -34303 -5192
rect -34702 -8445 -34303 -5193
rect -34702 -8447 -34553 -8445
rect -34702 -8512 -34692 -8447
rect -34629 -8510 -34553 -8447
rect -34490 -8447 -34303 -8445
rect -34490 -8510 -34397 -8447
rect -34629 -8512 -34397 -8510
rect -34334 -8512 -34303 -8447
rect -34702 -10165 -34303 -8512
rect -34702 -10172 -34394 -10165
rect -34702 -10255 -34688 -10172
rect -34632 -10176 -34394 -10172
rect -34632 -10255 -34544 -10176
rect -34702 -10259 -34544 -10255
rect -34488 -10248 -34394 -10176
rect -34338 -10248 -34303 -10165
rect -34488 -10259 -34303 -10248
rect -34702 -13749 -34303 -10259
rect -33805 -470 -33186 -361
rect -33077 -470 -32936 -361
rect -33805 -472 -32936 -470
rect -32825 -472 -32800 -361
rect -33805 -10435 -33694 -472
rect -33203 -493 -32800 -472
rect -30144 -683 -30087 -431
rect -33500 -981 -32481 -870
rect -33500 -9370 -33389 -981
rect -33055 -4142 -32542 -4116
rect -33055 -4147 -33023 -4142
rect -33057 -4292 -33023 -4147
rect -32873 -4143 -32542 -4142
rect -32873 -4291 -32705 -4143
rect -32557 -4291 -32542 -4143
rect -32873 -4292 -32542 -4291
rect -33057 -4311 -32542 -4292
rect -33048 -5355 -32977 -4311
rect -33082 -5379 -32956 -5355
rect -33082 -5434 -33042 -5379
rect -32987 -5434 -32956 -5379
rect -33082 -5490 -32956 -5434
rect -33082 -5545 -33041 -5490
rect -32986 -5545 -32956 -5490
rect -33082 -5567 -32956 -5545
rect -31594 -5868 -31538 -5666
rect -24190 -5855 -23791 2484
rect -24190 -5858 -23919 -5855
rect -24190 -5943 -24154 -5858
rect -24071 -5940 -23919 -5858
rect -23836 -5940 -23791 -5855
rect -24071 -5943 -23791 -5940
rect -32658 -6856 -32602 -6704
rect -32044 -8094 -31988 -7950
rect -33500 -9481 -32952 -9370
rect -33063 -9649 -32952 -9481
rect -33374 -9674 -32936 -9649
rect -33374 -9785 -33319 -9674
rect -33208 -9675 -32936 -9674
rect -33208 -9784 -33092 -9675
rect -32981 -9784 -32936 -9675
rect -33208 -9785 -32936 -9784
rect -33374 -9843 -32936 -9785
rect -33491 -10435 -33162 -10411
rect -33805 -10455 -33162 -10435
rect -33805 -10458 -33282 -10455
rect -33805 -10527 -33437 -10458
rect -33371 -10523 -33282 -10458
rect -33205 -10523 -33162 -10455
rect -33371 -10527 -33162 -10523
rect -33805 -10546 -33162 -10527
rect -33805 -11229 -33694 -10546
rect -33491 -10577 -33162 -10546
rect -33063 -10817 -32952 -9843
rect -33087 -10859 -32662 -10817
rect -33087 -10970 -33063 -10859
rect -32952 -10968 -32797 -10859
rect -32688 -10968 -32662 -10859
rect -32952 -10970 -32662 -10968
rect -33087 -10988 -32662 -10970
rect -33805 -11340 -33277 -11229
rect -34043 -12765 -33918 -12712
rect -34043 -12869 -34022 -12765
rect -33936 -12869 -33918 -12765
rect -34043 -13019 -33918 -12869
rect -34043 -13123 -34025 -13019
rect -33939 -13123 -33918 -13019
rect -34043 -13132 -33918 -13123
rect -34702 -13755 -34539 -13749
rect -34702 -13820 -34681 -13755
rect -34623 -13814 -34539 -13755
rect -34481 -13757 -34303 -13749
rect -34481 -13814 -34394 -13757
rect -34623 -13820 -34394 -13814
rect -34702 -13822 -34394 -13820
rect -34336 -13822 -34303 -13757
rect -34702 -13916 -34303 -13822
rect -34702 -13924 -34387 -13916
rect -34702 -13927 -34547 -13924
rect -34702 -13992 -34693 -13927
rect -34635 -13989 -34547 -13927
rect -34489 -13981 -34387 -13924
rect -34329 -13981 -34303 -13916
rect -34489 -13989 -34303 -13981
rect -34635 -13992 -34303 -13989
rect -34702 -17307 -34303 -13992
rect -34702 -17309 -34438 -17307
rect -34702 -17311 -34572 -17309
rect -34702 -17378 -34694 -17311
rect -34636 -17376 -34572 -17311
rect -34514 -17374 -34438 -17309
rect -34380 -17374 -34303 -17307
rect -34514 -17376 -34303 -17374
rect -34636 -17378 -34303 -17376
rect -34702 -19034 -34303 -17378
rect -34702 -19099 -34688 -19034
rect -34630 -19036 -34303 -19034
rect -34630 -19037 -34399 -19036
rect -34630 -19099 -34555 -19037
rect -34702 -19102 -34555 -19099
rect -34497 -19101 -34399 -19037
rect -34341 -19101 -34303 -19036
rect -34497 -19102 -34303 -19101
rect -34702 -21644 -34303 -19102
rect -34046 -20871 -33918 -13132
rect -34046 -20965 -34026 -20871
rect -33939 -20965 -33918 -20871
rect -34046 -21063 -33918 -20965
rect -34046 -21157 -34027 -21063
rect -33940 -21157 -33918 -21063
rect -34046 -21192 -33918 -21157
rect -34702 -21649 -34377 -21644
rect -34702 -21652 -34539 -21649
rect -34702 -21721 -34695 -21652
rect -34637 -21718 -34539 -21652
rect -34481 -21713 -34377 -21649
rect -34319 -21713 -34303 -21644
rect -34481 -21718 -34303 -21713
rect -34637 -21721 -34303 -21718
rect -34702 -25271 -34303 -21721
rect -34702 -25273 -34430 -25271
rect -34702 -25274 -34558 -25273
rect -34702 -25343 -34692 -25274
rect -34634 -25342 -34558 -25274
rect -34500 -25340 -34430 -25273
rect -34372 -25340 -34303 -25271
rect -34500 -25342 -34303 -25340
rect -34634 -25343 -34303 -25342
rect -34702 -26614 -34303 -25343
rect -33388 -26115 -33277 -11340
rect -33388 -26172 -33372 -26115
rect -33315 -26172 -33277 -26115
rect -33388 -26248 -33277 -26172
rect -33388 -26303 -33366 -26248
rect -33311 -26303 -33277 -26248
rect -33388 -26319 -33277 -26303
rect -34702 -26619 -34407 -26614
rect -34702 -26627 -34552 -26619
rect -34702 -26683 -34684 -26627
rect -34632 -26675 -34552 -26627
rect -34500 -26670 -34407 -26619
rect -34355 -26670 -34303 -26614
rect -34500 -26675 -34303 -26670
rect -34632 -26683 -34303 -26675
rect -34702 -26757 -34303 -26683
rect -34702 -26826 -34568 -26757
rect -34510 -26826 -34303 -26757
rect -34702 -26949 -34303 -26826
rect -34702 -27018 -34568 -26949
rect -34510 -27018 -34303 -26949
rect -34702 -29733 -34303 -27018
rect -33063 -26862 -32952 -10988
rect -25126 -11377 -25018 -11345
rect -25126 -11472 -25102 -11377
rect -25025 -11472 -25018 -11377
rect -25126 -11553 -25018 -11472
rect -25126 -11648 -25105 -11553
rect -25028 -11648 -25018 -11553
rect -25126 -11712 -25018 -11648
rect -25126 -11807 -25103 -11712
rect -25026 -11807 -25018 -11712
rect -25126 -11870 -25018 -11807
rect -25126 -11965 -25104 -11870
rect -25027 -11965 -25018 -11870
rect -25329 -12396 -25224 -12381
rect -25329 -12422 -25220 -12396
rect -25329 -12517 -25303 -12422
rect -25226 -12517 -25220 -12422
rect -25329 -12598 -25220 -12517
rect -25329 -12693 -25306 -12598
rect -25229 -12693 -25220 -12598
rect -32624 -12772 -32507 -12724
rect -32624 -12876 -32602 -12772
rect -32524 -12876 -32507 -12772
rect -32624 -12973 -32507 -12876
rect -32624 -13077 -32608 -12973
rect -32530 -13077 -32507 -12973
rect -32624 -15754 -32507 -13077
rect -25329 -12757 -25220 -12693
rect -25329 -12852 -25304 -12757
rect -25227 -12852 -25220 -12757
rect -25329 -12915 -25220 -12852
rect -25329 -13010 -25305 -12915
rect -25228 -13010 -25220 -12915
rect -25329 -13033 -25220 -13010
rect -25329 -13934 -25224 -13033
rect -25126 -13936 -25018 -11965
rect -24190 -14610 -23791 -5943
rect -24190 -14613 -23911 -14610
rect -24190 -14614 -24046 -14613
rect -24190 -14699 -24181 -14614
rect -24108 -14698 -24046 -14614
rect -23973 -14695 -23911 -14613
rect -23838 -14695 -23791 -14610
rect -23973 -14698 -23791 -14695
rect -24108 -14699 -23791 -14698
rect -31868 -14996 -31781 -14975
rect -31868 -15052 -31855 -14996
rect -31799 -15052 -31781 -14996
rect -31868 -15107 -31781 -15052
rect -31868 -15163 -31859 -15107
rect -31803 -15163 -31781 -15107
rect -31868 -15178 -31781 -15163
rect -29583 -15746 -29527 -15485
rect -32618 -15769 -32515 -15754
rect -32618 -15868 -32597 -15769
rect -32527 -15868 -32515 -15769
rect -32618 -15949 -32515 -15868
rect -32618 -16048 -32602 -15949
rect -32532 -16048 -32515 -15949
rect -32618 -16071 -32515 -16048
rect -29580 -16181 -29524 -15915
rect -32218 -16809 -32087 -16789
rect -32218 -16887 -32183 -16809
rect -32114 -16887 -32087 -16809
rect -32218 -16991 -32087 -16887
rect -32218 -17069 -32183 -16991
rect -32114 -17069 -32087 -16991
rect -32218 -17083 -32087 -17069
rect -33063 -26919 -33031 -26862
rect -32973 -26919 -32952 -26862
rect -33063 -26984 -32952 -26919
rect -33063 -27041 -33034 -26984
rect -32976 -27041 -32952 -26984
rect -33063 -27096 -32952 -27041
rect -32301 -18227 -32191 -18209
rect -32301 -18302 -32277 -18227
rect -32202 -18302 -32191 -18227
rect -32301 -18395 -32191 -18302
rect -32301 -18472 -32277 -18395
rect -32200 -18472 -32191 -18395
rect -32301 -19528 -32191 -18472
rect -29531 -18510 -29474 -18272
rect -31957 -18717 -31899 -18622
rect -32301 -19589 -32280 -19528
rect -32218 -19589 -32191 -19528
rect -32301 -19656 -32191 -19589
rect -32301 -19717 -32282 -19656
rect -32220 -19717 -32191 -19656
rect -32301 -21308 -32191 -19717
rect -32301 -21380 -32282 -21308
rect -32210 -21380 -32191 -21308
rect -32301 -21494 -32191 -21380
rect -32301 -21568 -32283 -21494
rect -32209 -21568 -32191 -21494
rect -32667 -28586 -32557 -28559
rect -32667 -28652 -32650 -28586
rect -32581 -28652 -32557 -28586
rect -32667 -28706 -32557 -28652
rect -32667 -28772 -32652 -28706
rect -32583 -28772 -32557 -28706
rect -34702 -29734 -34424 -29733
rect -34702 -29738 -34562 -29734
rect -34702 -29818 -34684 -29738
rect -34627 -29814 -34562 -29738
rect -34505 -29813 -34424 -29734
rect -34367 -29813 -34303 -29733
rect -34505 -29814 -34303 -29813
rect -34627 -29818 -34303 -29814
rect -34702 -33379 -34303 -29818
rect -32960 -28848 -32850 -28826
rect -32960 -28909 -32932 -28848
rect -32873 -28909 -32850 -28848
rect -32960 -28964 -32850 -28909
rect -32960 -29025 -32939 -28964
rect -32880 -29025 -32850 -28964
rect -32960 -30135 -32850 -29025
rect -32667 -29396 -32557 -28772
rect -32675 -29432 -32550 -29396
rect -32675 -29506 -32649 -29432
rect -32575 -29506 -32550 -29432
rect -32675 -29606 -32550 -29506
rect -32675 -29678 -32648 -29606
rect -32576 -29678 -32550 -29606
rect -32675 -29697 -32550 -29678
rect -32960 -30207 -32935 -30135
rect -32865 -30207 -32850 -30135
rect -32960 -30289 -32850 -30207
rect -32960 -30361 -32943 -30289
rect -32873 -30361 -32850 -30289
rect -32960 -30385 -32850 -30361
rect -32953 -30387 -32858 -30385
rect -34702 -33382 -34393 -33379
rect -34702 -33450 -34697 -33382
rect -34640 -33450 -34562 -33382
rect -34505 -33447 -34393 -33382
rect -34336 -33447 -34303 -33379
rect -34505 -33450 -34303 -33447
rect -34702 -34909 -34303 -33450
rect -32301 -34404 -32191 -21568
rect -31977 -19337 -31878 -18717
rect -31977 -19393 -31960 -19337
rect -31904 -19393 -31878 -19337
rect -31977 -19459 -31878 -19393
rect -31977 -19515 -31954 -19459
rect -31898 -19515 -31878 -19459
rect -31977 -21859 -31878 -19515
rect -31977 -21922 -31954 -21859
rect -31889 -21922 -31878 -21859
rect -31977 -22031 -31878 -21922
rect -31977 -22094 -31959 -22031
rect -31894 -22094 -31878 -22031
rect -31977 -23781 -31878 -22094
rect -24190 -22593 -23791 -14699
rect -24190 -22600 -23895 -22593
rect -24190 -22603 -24039 -22600
rect -24190 -22690 -24172 -22603
rect -24112 -22687 -24039 -22603
rect -23979 -22680 -23895 -22600
rect -23835 -22680 -23791 -22593
rect -23979 -22687 -23791 -22680
rect -24112 -22690 -23791 -22687
rect -32301 -34461 -32275 -34404
rect -32218 -34461 -32191 -34404
rect -32301 -34546 -32191 -34461
rect -32301 -34601 -32275 -34546
rect -32220 -34601 -32191 -34546
rect -32301 -34619 -32191 -34601
rect -32095 -23880 -31878 -23781
rect -30680 -23859 -30624 -23704
rect -34702 -34912 -34553 -34909
rect -34702 -34975 -34685 -34912
rect -34625 -34972 -34553 -34912
rect -34493 -34912 -34303 -34909
rect -34493 -34972 -34419 -34912
rect -34625 -34975 -34419 -34972
rect -34359 -34975 -34303 -34912
rect -34702 -36496 -34303 -34975
rect -32095 -35207 -31996 -23880
rect -31294 -24958 -31238 -24848
rect -30230 -26131 -30174 -25935
rect -24190 -30639 -23791 -22690
rect -24190 -30642 -24024 -30639
rect -24190 -30705 -24156 -30642
rect -24096 -30702 -24024 -30642
rect -23964 -30642 -23791 -30639
rect -23964 -30702 -23890 -30642
rect -24096 -30705 -23890 -30702
rect -23830 -30705 -23791 -30642
rect -24190 -31074 -23791 -30705
rect -24190 -31077 -24024 -31074
rect -24190 -31140 -24156 -31077
rect -24096 -31137 -24024 -31077
rect -23964 -31077 -23791 -31074
rect -23964 -31137 -23890 -31077
rect -24096 -31140 -23890 -31137
rect -23830 -31140 -23791 -31077
rect -30645 -32148 -30589 -32012
rect -31259 -33363 -31203 -33224
rect -30195 -34428 -30139 -34228
rect -32095 -35260 -32072 -35207
rect -32010 -35260 -31996 -35207
rect -32095 -35355 -31996 -35260
rect -32095 -35408 -32075 -35355
rect -32013 -35408 -31996 -35355
rect -32095 -35423 -31996 -35408
rect -24190 -36034 -23791 -31140
rect -24190 -36035 -24036 -36034
rect -24190 -36120 -24177 -36035
rect -24120 -36119 -24036 -36035
rect -23979 -36035 -23791 -36034
rect -23979 -36119 -23891 -36035
rect -24120 -36120 -23891 -36119
rect -23834 -36120 -23791 -36035
rect -34702 -36513 -34290 -36496
rect -34702 -36516 -34373 -36513
rect -34702 -36521 -34522 -36516
rect -34702 -36616 -34681 -36521
rect -34604 -36611 -34522 -36521
rect -34445 -36608 -34373 -36516
rect -34296 -36608 -34290 -36513
rect -34445 -36611 -34290 -36608
rect -34604 -36616 -34290 -36611
rect -34702 -36689 -34290 -36616
rect -34702 -36692 -34376 -36689
rect -34702 -36697 -34525 -36692
rect -34702 -36792 -34684 -36697
rect -34607 -36787 -34525 -36697
rect -34448 -36784 -34376 -36692
rect -34299 -36784 -34290 -36689
rect -34448 -36787 -34290 -36784
rect -34607 -36792 -34290 -36787
rect -34702 -36848 -34290 -36792
rect -34702 -36851 -34374 -36848
rect -34702 -36856 -34523 -36851
rect -34702 -36951 -34682 -36856
rect -34605 -36946 -34523 -36856
rect -34446 -36943 -34374 -36851
rect -34297 -36943 -34290 -36848
rect -34446 -36946 -34290 -36943
rect -34605 -36951 -34290 -36946
rect -34702 -37006 -34290 -36951
rect -34702 -37009 -34375 -37006
rect -34702 -37014 -34524 -37009
rect -34702 -37109 -34683 -37014
rect -34606 -37104 -34524 -37014
rect -34447 -37101 -34375 -37009
rect -34298 -37101 -34290 -37006
rect -34447 -37104 -34290 -37101
rect -34606 -37109 -34290 -37104
rect -34702 -37121 -34290 -37109
rect -35392 -37560 -34980 -37543
rect -35392 -37563 -35063 -37560
rect -35392 -37568 -35212 -37563
rect -35392 -37663 -35371 -37568
rect -35294 -37658 -35212 -37568
rect -35135 -37655 -35063 -37563
rect -34986 -37655 -34980 -37560
rect -35135 -37658 -34980 -37655
rect -35294 -37663 -34980 -37658
rect -35392 -37736 -34980 -37663
rect -35392 -37739 -35066 -37736
rect -35392 -37744 -35215 -37739
rect -35392 -37839 -35374 -37744
rect -35297 -37834 -35215 -37744
rect -35138 -37831 -35066 -37739
rect -34989 -37831 -34980 -37736
rect -35138 -37834 -34980 -37831
rect -35297 -37839 -34980 -37834
rect -35392 -37895 -34980 -37839
rect -35392 -37898 -35064 -37895
rect -35392 -37903 -35213 -37898
rect -35392 -37998 -35372 -37903
rect -35295 -37993 -35213 -37903
rect -35136 -37990 -35064 -37898
rect -34987 -37990 -34980 -37895
rect -35136 -37993 -34980 -37990
rect -35295 -37998 -34980 -37993
rect -35392 -38053 -34980 -37998
rect -35392 -38056 -35065 -38053
rect -35392 -38061 -35214 -38056
rect -35392 -38156 -35373 -38061
rect -35296 -38151 -35214 -38061
rect -35137 -38148 -35065 -38056
rect -34988 -38148 -34980 -38053
rect -35137 -38151 -34980 -38148
rect -35296 -38156 -34980 -38151
rect -35392 -38168 -34980 -38156
rect -35392 -38309 -34993 -38168
rect -34702 -38309 -34303 -37121
rect -24190 -37532 -23791 -36120
rect -23397 30752 -22998 32140
rect -23397 30750 -23091 30752
rect -23397 30667 -23377 30750
rect -23307 30667 -23227 30750
rect -23157 30669 -23091 30750
rect -23021 30669 -22998 30752
rect -23157 30667 -22998 30669
rect -23397 25787 -22998 30667
rect -19720 40738 -19576 40765
rect -19720 40664 -19690 40738
rect -19616 40664 -19576 40738
rect -19720 40608 -19576 40664
rect -19720 40534 -19689 40608
rect -19615 40534 -19576 40608
rect -19720 40472 -19576 40534
rect -19720 40398 -19689 40472
rect -19615 40398 -19576 40472
rect -19720 32255 -19576 40398
rect -18963 38367 -18879 43792
rect -18496 43756 -18336 43788
rect -18496 43647 -18472 43756
rect -18363 43750 -18336 43756
rect -18496 43641 -18470 43647
rect -18361 43641 -18336 43750
rect -18496 43398 -18336 43641
rect -18496 43287 -18472 43398
rect -18361 43287 -18336 43398
rect -18496 43267 -18336 43287
rect -11255 43758 -11242 43853
rect -11165 43758 -11150 43853
rect -11255 43695 -11150 43758
rect -11255 43600 -11243 43695
rect -11166 43600 -11150 43695
rect -11255 43269 -11150 43600
rect -18470 38908 -18359 43267
rect -11255 43213 -11227 43269
rect -11172 43213 -11150 43269
rect -11255 42536 -11150 43213
rect -11052 43130 -10944 44643
rect -11052 43074 -11021 43130
rect -10966 43074 -10944 43130
rect -11052 42717 -10944 43074
rect -17825 41655 -17702 41669
rect -17825 41576 -17805 41655
rect -17714 41576 -17702 41655
rect -17825 41503 -17702 41576
rect -17825 41424 -17809 41503
rect -17718 41424 -17702 41503
rect -17825 41412 -17702 41424
rect -15509 41630 -15453 41635
rect -15509 41574 -14911 41630
rect -15509 41352 -15453 41574
rect -15506 40553 -15505 40604
rect -15451 40553 -15450 40604
rect -15506 40375 -15450 40553
rect -18489 38886 -18167 38908
rect -18489 38775 -18470 38886
rect -18359 38885 -18167 38886
rect -18359 38776 -18296 38885
rect -18187 38776 -18167 38885
rect -18359 38775 -18167 38776
rect -18489 38756 -18167 38775
rect -19001 38331 -18631 38367
rect -19001 38247 -18963 38331
rect -18879 38247 -18731 38331
rect -18647 38247 -18631 38331
rect -19001 38224 -18631 38247
rect -19314 33244 -19162 33285
rect -19314 33156 -19287 33244
rect -19196 33156 -19162 33244
rect -19314 33037 -19162 33156
rect -19314 32949 -19284 33037
rect -19193 32949 -19162 33037
rect -19314 32922 -19162 32949
rect -19720 32173 -19684 32255
rect -19601 32173 -19576 32255
rect -19720 32071 -19576 32173
rect -19720 31989 -19685 32071
rect -19602 31989 -19576 32071
rect -19720 27625 -19576 31989
rect -19720 27552 -19700 27625
rect -19604 27552 -19576 27625
rect -19720 27458 -19576 27552
rect -19720 27385 -19696 27458
rect -19600 27385 -19576 27458
rect -19720 27362 -19576 27385
rect -23397 25785 -23087 25787
rect -23397 25782 -23236 25785
rect -23397 25670 -23387 25782
rect -23311 25673 -23236 25782
rect -23160 25675 -23087 25785
rect -23011 25675 -22998 25787
rect -23160 25673 -22998 25675
rect -23311 25670 -22998 25673
rect -23397 22530 -22998 25670
rect -23397 22526 -23124 22530
rect -23397 22436 -23365 22526
rect -23275 22440 -23124 22526
rect -23034 22440 -22998 22530
rect -23275 22436 -22998 22440
rect -23397 17163 -22998 22436
rect -19635 23815 -19480 23883
rect -19635 23758 -19606 23815
rect -19517 23758 -19480 23815
rect -19635 23695 -19480 23758
rect -19635 23638 -19605 23695
rect -19516 23638 -19480 23695
rect -19635 23586 -19480 23638
rect -19635 23529 -19606 23586
rect -19517 23529 -19480 23586
rect -23397 17158 -23091 17163
rect -23397 17074 -23382 17158
rect -23325 17156 -23091 17158
rect -23325 17074 -23236 17156
rect -23397 17072 -23236 17074
rect -23179 17079 -23091 17156
rect -23034 17079 -22998 17163
rect -23179 17072 -22998 17079
rect -23397 13531 -22998 17072
rect -23397 13526 -23242 13531
rect -23397 13448 -23387 13526
rect -23320 13453 -23242 13526
rect -23175 13529 -22998 13531
rect -23175 13453 -23103 13529
rect -23320 13451 -23103 13453
rect -23036 13451 -22998 13529
rect -23320 13448 -22998 13451
rect -23397 11794 -22998 13448
rect -23397 11703 -23383 11794
rect -23316 11792 -22998 11794
rect -23316 11703 -23227 11792
rect -23397 11701 -23227 11703
rect -23160 11701 -23095 11792
rect -23028 11701 -22998 11792
rect -23397 8799 -22998 11701
rect -23397 8792 -23225 8799
rect -23397 8718 -23371 8792
rect -23304 8725 -23225 8792
rect -23158 8725 -23080 8799
rect -23013 8725 -22998 8799
rect -23304 8718 -22998 8725
rect -23397 8658 -22998 8718
rect -23397 8650 -23077 8658
rect -23397 8646 -23220 8650
rect -23397 8572 -23370 8646
rect -23303 8576 -23220 8646
rect -23153 8584 -23077 8650
rect -23010 8584 -22998 8658
rect -23153 8576 -22998 8584
rect -23303 8572 -22998 8576
rect -23397 8498 -22998 8572
rect -23397 8494 -23116 8498
rect -23397 8400 -23367 8494
rect -23280 8404 -23116 8494
rect -23029 8404 -22998 8498
rect -23280 8400 -22998 8404
rect -23397 3692 -22998 8400
rect -23397 3689 -23100 3692
rect -23397 3684 -23241 3689
rect -23397 3616 -23380 3684
rect -23325 3621 -23241 3684
rect -23186 3624 -23100 3689
rect -23045 3624 -22998 3692
rect -23186 3621 -22998 3624
rect -23325 3616 -22998 3621
rect -23397 3503 -22998 3616
rect -23397 3498 -23244 3503
rect -23397 3430 -23388 3498
rect -23333 3435 -23244 3498
rect -23189 3435 -23086 3503
rect -23031 3435 -22998 3503
rect -23333 3430 -22998 3435
rect -23397 -123 -22998 3430
rect -23397 -125 -23092 -123
rect -23397 -193 -23386 -125
rect -23332 -126 -23092 -125
rect -23332 -193 -23235 -126
rect -23397 -194 -23235 -193
rect -23181 -191 -23092 -126
rect -23038 -191 -22998 -123
rect -23181 -194 -22998 -191
rect -23397 -1127 -22998 -194
rect -23397 -1132 -23103 -1127
rect -23397 -1134 -23254 -1132
rect -23397 -1202 -23389 -1134
rect -23334 -1200 -23254 -1134
rect -23199 -1195 -23103 -1132
rect -23048 -1195 -22998 -1127
rect -23199 -1200 -22998 -1195
rect -23334 -1202 -22998 -1200
rect -23397 -1271 -22998 -1202
rect -23397 -1272 -23104 -1271
rect -23397 -1274 -23251 -1272
rect -23397 -1342 -23392 -1274
rect -23337 -1340 -23251 -1274
rect -23196 -1339 -23104 -1272
rect -23049 -1339 -22998 -1271
rect -23196 -1340 -22998 -1339
rect -23337 -1342 -22998 -1340
rect -23397 -5119 -22998 -1342
rect -22353 20533 -21948 20557
rect -22353 20530 -22103 20533
rect -22353 20463 -22292 20530
rect -22216 20466 -22103 20530
rect -22027 20466 -21948 20533
rect -22216 20463 -21948 20466
rect -22353 20421 -21948 20463
rect -22353 -4555 -22217 20421
rect -22046 20179 -21671 20221
rect -22046 20112 -21949 20179
rect -21873 20112 -21783 20179
rect -21707 20112 -21671 20179
rect -22046 20085 -21671 20112
rect -22046 -4156 -21910 20085
rect -21254 19415 -21069 19444
rect -21254 19320 -21211 19415
rect -21134 19320 -21069 19415
rect -21254 19239 -21069 19320
rect -19635 19243 -19480 23529
rect -19290 22890 -19182 32922
rect -18963 29852 -18879 38224
rect -18470 30389 -18359 38756
rect -9364 38740 -9133 46185
rect -9364 38670 -9350 38740
rect -9270 38670 -9133 38740
rect -9364 38620 -9133 38670
rect -9364 38550 -9250 38620
rect -9170 38550 -9133 38620
rect -15457 38105 -15400 38282
rect -15403 38047 -15400 38105
rect -11156 37020 -11048 37057
rect -11156 36925 -11137 37020
rect -11060 36925 -11048 37020
rect -11156 36844 -11048 36925
rect -11156 36749 -11140 36844
rect -11063 36749 -11048 36844
rect -11156 36685 -11048 36749
rect -11156 36590 -11138 36685
rect -11061 36590 -11048 36685
rect -11156 36527 -11048 36590
rect -11156 36432 -11139 36527
rect -11062 36432 -11048 36527
rect -11359 35770 -11254 35802
rect -11359 35675 -11338 35770
rect -11261 35675 -11254 35770
rect -11359 35594 -11254 35675
rect -11359 35499 -11341 35594
rect -11264 35499 -11254 35594
rect -11359 35435 -11254 35499
rect -11359 35340 -11339 35435
rect -11262 35340 -11254 35435
rect -11359 35277 -11254 35340
rect -11359 35182 -11340 35277
rect -11263 35182 -11254 35277
rect -11359 34087 -11254 35182
rect -11156 34081 -11048 36432
rect -17936 33150 -17813 33164
rect -17936 33071 -17916 33150
rect -17825 33071 -17813 33150
rect -17936 32998 -17813 33071
rect -17936 32919 -17920 32998
rect -17829 32919 -17813 32998
rect -17936 32907 -17813 32919
rect -15613 32558 -15557 32700
rect -15610 31935 -15554 32093
rect -18227 31174 -18104 31188
rect -18227 31095 -18207 31174
rect -18116 31095 -18104 31174
rect -18227 31022 -18104 31095
rect -18227 30943 -18211 31022
rect -18120 30943 -18104 31022
rect -18227 30931 -18104 30943
rect -18480 30372 -18152 30389
rect -18480 30261 -18470 30372
rect -18359 30371 -18152 30372
rect -18359 30262 -18285 30371
rect -18176 30262 -18152 30371
rect -18359 30261 -18152 30262
rect -18480 30245 -18152 30261
rect -18994 29819 -18656 29852
rect -18994 29735 -18963 29819
rect -18879 29735 -18763 29819
rect -18679 29735 -18656 29819
rect -18994 29712 -18656 29735
rect -18963 28021 -18879 29712
rect -18470 28550 -18359 30245
rect -15561 29520 -15504 29770
rect -18489 28532 -18088 28550
rect -18489 28421 -18470 28532
rect -18359 28421 -18221 28532
rect -18110 28421 -18088 28532
rect -18489 28406 -18088 28421
rect -11866 28456 -11758 28514
rect -11866 28361 -11847 28456
rect -11770 28361 -11758 28456
rect -11866 28280 -11758 28361
rect -11866 28185 -11850 28280
rect -11773 28185 -11758 28280
rect -11866 28121 -11758 28185
rect -11866 28026 -11848 28121
rect -11771 28026 -11758 28121
rect -18981 28006 -18651 28021
rect -18981 27922 -18963 28006
rect -18879 27922 -18739 28006
rect -18655 27922 -18651 28006
rect -18981 27901 -18651 27922
rect -11866 27963 -11758 28026
rect -11866 27868 -11849 27963
rect -11772 27868 -11758 27963
rect -12069 27358 -11964 27394
rect -12069 27263 -12047 27358
rect -11970 27263 -11964 27358
rect -12069 27182 -11964 27263
rect -12069 27087 -12050 27182
rect -11973 27087 -11964 27182
rect -12069 27023 -11964 27087
rect -12069 26928 -12048 27023
rect -11971 26928 -11964 27023
rect -12069 26865 -11964 26928
rect -12069 26770 -12049 26865
rect -11972 26770 -11964 26865
rect -12069 25795 -11964 26770
rect -11866 25929 -11758 27868
rect -9364 26764 -9133 38550
rect -9364 26761 -9213 26764
rect -9364 26695 -9349 26761
rect -9295 26698 -9213 26761
rect -9159 26698 -9133 26764
rect -9295 26695 -9133 26698
rect -9364 26662 -9133 26695
rect -7915 40490 -7516 47634
rect -7915 40434 -7900 40490
rect -7848 40434 -7768 40490
rect -7716 40489 -7516 40490
rect -7716 40434 -7647 40489
rect -7915 40433 -7647 40434
rect -7595 40433 -7516 40489
rect -7915 33552 -7516 40433
rect -7915 33542 -7615 33552
rect -7915 33534 -7749 33542
rect -7915 33474 -7902 33534
rect -7848 33482 -7749 33534
rect -7695 33492 -7615 33542
rect -7561 33492 -7516 33552
rect -7695 33482 -7516 33492
rect -7848 33474 -7516 33482
rect -7915 26211 -7516 33474
rect -7915 26205 -7615 26211
rect -7915 26200 -7764 26205
rect -7915 26147 -7904 26200
rect -7852 26152 -7764 26200
rect -7712 26158 -7615 26205
rect -7563 26158 -7516 26211
rect -7712 26152 -7516 26158
rect -7852 26147 -7516 26152
rect -9420 25965 -9188 25978
rect -9420 25961 -9271 25965
rect -9420 25907 -9399 25961
rect -9345 25909 -9271 25961
rect -9215 25909 -9188 25965
rect -9345 25907 -9188 25909
rect -9420 25854 -9188 25907
rect -9420 25849 -9269 25854
rect -9420 25793 -9399 25849
rect -9343 25800 -9269 25849
rect -9215 25800 -9188 25854
rect -9343 25793 -9188 25800
rect -9420 25788 -9188 25793
rect -18635 24891 -18512 24905
rect -18635 24812 -18615 24891
rect -18524 24812 -18512 24891
rect -18635 24739 -18512 24812
rect -18635 24660 -18619 24739
rect -18528 24660 -18512 24739
rect -18635 24648 -18512 24660
rect -16323 24071 -16267 24255
rect -16320 23630 -16264 23884
rect -19049 22965 -18926 22979
rect -19049 22890 -19029 22965
rect -19290 22886 -19029 22890
rect -18938 22886 -18926 22965
rect -19290 22813 -18926 22886
rect -19290 22782 -19033 22813
rect -19049 22734 -19033 22782
rect -18942 22734 -18926 22813
rect -19049 22722 -18926 22734
rect -19217 21575 -18885 21609
rect -19217 21571 -18989 21575
rect -19217 21499 -19197 21571
rect -19131 21503 -18989 21571
rect -18923 21554 -18885 21575
rect -18923 21503 -18882 21554
rect -19131 21499 -18882 21503
rect -19217 21451 -18882 21499
rect -19096 19523 -18993 21451
rect -16271 21287 -16214 21534
rect -18697 21111 -18639 21158
rect -18719 19864 -18616 21111
rect -18839 19820 -18567 19864
rect -18839 19817 -18672 19820
rect -18839 19761 -18824 19817
rect -18767 19764 -18672 19817
rect -18615 19764 -18567 19820
rect -18767 19761 -18567 19764
rect -18839 19728 -18567 19761
rect -19113 19479 -18841 19523
rect -19113 19476 -18946 19479
rect -19113 19420 -19098 19476
rect -19041 19423 -18946 19476
rect -18889 19423 -18841 19479
rect -19041 19420 -18841 19423
rect -19113 19387 -18841 19420
rect -21254 19144 -21214 19239
rect -21137 19144 -21069 19239
rect -21254 19080 -21069 19144
rect -21254 18985 -21212 19080
rect -21135 18985 -21069 19080
rect -21254 18922 -21069 18985
rect -21254 18827 -21213 18922
rect -21136 18827 -21069 18922
rect -21254 14604 -21069 18827
rect -19637 19199 -19478 19243
rect -19637 19093 -19604 19199
rect -19511 19093 -19478 19199
rect -19637 19022 -19478 19093
rect -19637 18954 -19603 19022
rect -19508 18954 -19478 19022
rect -19637 18859 -19478 18954
rect -19637 18769 -19596 18859
rect -19505 18769 -19478 18859
rect -19637 18743 -19478 18769
rect -20750 18363 -20645 18368
rect -20785 18346 -20618 18363
rect -20785 18251 -20728 18346
rect -20651 18251 -20618 18346
rect -20785 18170 -20618 18251
rect -20785 18075 -20731 18170
rect -20654 18075 -20618 18170
rect -20785 18011 -20618 18075
rect -20785 17916 -20729 18011
rect -20652 17916 -20618 18011
rect -20785 17853 -20618 17916
rect -20785 17758 -20730 17853
rect -20653 17758 -20618 17853
rect -20785 15975 -20618 17758
rect -9419 17179 -9188 25788
rect -8429 24913 -8229 25001
rect -8429 24801 -8395 24913
rect -8259 24801 -8229 24913
rect -8429 24643 -8229 24801
rect -8429 24531 -8407 24643
rect -8271 24531 -8229 24643
rect -8429 24503 -8229 24531
rect -9403 17021 -9322 17179
rect -20785 15942 -20361 15975
rect -20785 15941 -20524 15942
rect -20785 15848 -20770 15941
rect -20784 15816 -20770 15848
rect -20644 15816 -20524 15941
rect -20784 15815 -20524 15816
rect -20397 15815 -20361 15942
rect -20784 15794 -20361 15815
rect -20253 15406 -20108 15455
rect -20253 15320 -20225 15406
rect -20135 15320 -20108 15406
rect -20253 15201 -20108 15320
rect -20253 15115 -20229 15201
rect -20139 15153 -20108 15201
rect -20139 15115 -9632 15153
rect -20253 15114 -9632 15115
rect -20253 15113 -9726 15114
rect -20253 15090 -9885 15113
rect -20240 15037 -9885 15090
rect -9818 15038 -9726 15113
rect -9659 15038 -9632 15114
rect -9818 15037 -9632 15038
rect -20240 15021 -9632 15037
rect -21254 14419 -20635 14604
rect -8912 13773 -8567 13774
rect -8413 13773 -8238 24503
rect -20257 13730 -19895 13763
rect -8912 13730 -8238 13773
rect -20257 13729 -8685 13730
rect -20257 13726 -20022 13729
rect -20257 13625 -20237 13726
rect -20151 13628 -20022 13726
rect -19936 13727 -8685 13729
rect -19936 13628 -8891 13727
rect -20151 13626 -8891 13628
rect -20151 13625 -19895 13626
rect -20257 13609 -19895 13625
rect -8912 13624 -8891 13626
rect -8801 13627 -8685 13727
rect -8595 13627 -8238 13730
rect -8801 13624 -8238 13627
rect -8912 13598 -8238 13624
rect -7915 23493 -7516 26147
rect -7915 23490 -7640 23493
rect -7915 23486 -7776 23490
rect -7915 23429 -7897 23486
rect -7845 23433 -7776 23486
rect -7724 23436 -7640 23490
rect -7588 23436 -7516 23493
rect -7724 23433 -7516 23436
rect -7845 23429 -7516 23433
rect -7915 16078 -7516 23429
rect -7915 16077 -7622 16078
rect -7915 16014 -7892 16077
rect -7830 16014 -7758 16077
rect -7696 16015 -7622 16077
rect -7560 16015 -7516 16078
rect -7696 16014 -7516 16015
rect -8912 13590 -8567 13598
rect -19498 12835 -19442 13004
rect -18808 9831 -18709 9847
rect -18808 9756 -18798 9831
rect -18733 9830 -18223 9831
rect -18733 9828 -18072 9830
rect -18733 9776 -18261 9828
rect -18209 9826 -18072 9828
rect -18209 9776 -18155 9826
rect -18733 9774 -18155 9776
rect -18095 9774 -18072 9826
rect -18733 9764 -18072 9774
rect -18733 9756 -18223 9764
rect -18808 9744 -18709 9756
rect -20210 8700 -20145 9281
rect -18818 8703 -18712 8715
rect -18818 8700 -18798 8703
rect -20210 8635 -18798 8700
rect -18733 8635 -18712 8703
rect -18818 8569 -18712 8635
rect -18818 8504 -18798 8569
rect -18733 8504 -18712 8569
rect -18818 8483 -18712 8504
rect -15954 7717 -15785 7718
rect -15954 7632 -15782 7717
rect -16008 5052 -15871 5123
rect -14474 5052 -14341 5117
rect -7915 3394 -7516 16014
rect -7915 3392 -7610 3394
rect -7915 3390 -7746 3392
rect -7915 3317 -7895 3390
rect -7828 3319 -7746 3390
rect -7679 3321 -7610 3392
rect -7543 3321 -7516 3394
rect -7679 3319 -7516 3321
rect -7828 3317 -7516 3319
rect -17047 2982 -16991 3106
rect -17903 705 -17847 790
rect -18527 -60 -18410 54
rect -18829 -138 -18331 -60
rect -18829 -223 -18813 -138
rect -18748 -223 -18638 -138
rect -18573 -180 -18331 -138
rect -18573 -223 -18217 -180
rect -18829 -256 -18217 -223
rect -18527 -297 -18217 -256
rect -19319 -1522 -18197 -1432
rect -19319 -4002 -19229 -1522
rect -18823 -1750 -17846 -1662
rect -19331 -4020 -19200 -4002
rect -19331 -4110 -19319 -4020
rect -19229 -4110 -19200 -4020
rect -22046 -4179 -21602 -4156
rect -22046 -4186 -21740 -4179
rect -22046 -4262 -21964 -4186
rect -21877 -4255 -21740 -4186
rect -21653 -4255 -21602 -4179
rect -21877 -4262 -21602 -4255
rect -22046 -4292 -21602 -4262
rect -19331 -4184 -19200 -4110
rect -19331 -4274 -19319 -4184
rect -19229 -4274 -19200 -4184
rect -19331 -4285 -19200 -4274
rect -18823 -4315 -18735 -1750
rect -12589 -2455 -12479 -2429
rect -12589 -2550 -12562 -2455
rect -12485 -2550 -12479 -2455
rect -12589 -2631 -12479 -2550
rect -12589 -2726 -12565 -2631
rect -12488 -2726 -12479 -2631
rect -12589 -2790 -12479 -2726
rect -12589 -2885 -12563 -2790
rect -12486 -2885 -12479 -2790
rect -12589 -2948 -12479 -2885
rect -12589 -3043 -12564 -2948
rect -12487 -3043 -12479 -2948
rect -12589 -3066 -12479 -3043
rect -12792 -3507 -12687 -3480
rect -12792 -3533 -12685 -3507
rect -12792 -3628 -12768 -3533
rect -12691 -3628 -12685 -3533
rect -12792 -3709 -12685 -3628
rect -12792 -3804 -12771 -3709
rect -12694 -3804 -12685 -3709
rect -12792 -3868 -12685 -3804
rect -12792 -3963 -12769 -3868
rect -12692 -3963 -12685 -3868
rect -12792 -4026 -12685 -3963
rect -12792 -4121 -12770 -4026
rect -12693 -4121 -12685 -4026
rect -12792 -4144 -12685 -4121
rect -18836 -4334 -18723 -4315
rect -18836 -4422 -18823 -4334
rect -18735 -4422 -18723 -4334
rect -18836 -4515 -18723 -4422
rect -22353 -4574 -21893 -4555
rect -22353 -4579 -22080 -4574
rect -22353 -4655 -22308 -4579
rect -22221 -4650 -22080 -4579
rect -21993 -4650 -21893 -4574
rect -18836 -4603 -18823 -4515
rect -18735 -4603 -18723 -4515
rect -18836 -4614 -18723 -4603
rect -22221 -4655 -21893 -4650
rect -22353 -4691 -21893 -4655
rect -23397 -5192 -23384 -5119
rect -23313 -5124 -22998 -5119
rect -23313 -5192 -23227 -5124
rect -23397 -5197 -23227 -5192
rect -23156 -5128 -22998 -5124
rect -23156 -5197 -23074 -5128
rect -23397 -5201 -23074 -5197
rect -23003 -5201 -22998 -5128
rect -12792 -5165 -12687 -4144
rect -23397 -8613 -22998 -5201
rect -12589 -5227 -12481 -3066
rect -19347 -6183 -19260 -6162
rect -19347 -6239 -19334 -6183
rect -19278 -6239 -19260 -6183
rect -19347 -6294 -19260 -6239
rect -19347 -6350 -19338 -6294
rect -19282 -6350 -19260 -6294
rect -19347 -6365 -19260 -6350
rect -17046 -7022 -16990 -6778
rect -23397 -8618 -23115 -8613
rect -23397 -8703 -23378 -8618
rect -23292 -8698 -23115 -8618
rect -23029 -8698 -22998 -8613
rect -23292 -8703 -22998 -8698
rect -23397 -10059 -22998 -8703
rect -23397 -10132 -23386 -10059
rect -23315 -10062 -22998 -10059
rect -23315 -10132 -23233 -10062
rect -23397 -10135 -23233 -10132
rect -23162 -10135 -23078 -10062
rect -23007 -10135 -22998 -10062
rect -23397 -13606 -22998 -10135
rect -20587 -7178 -20448 -7167
rect -20587 -7249 -20561 -7178
rect -20476 -7249 -20448 -7178
rect -20587 -7319 -20448 -7249
rect -20587 -7390 -20563 -7319
rect -20478 -7390 -20448 -7319
rect -20587 -7458 -20448 -7390
rect -20587 -7529 -20568 -7458
rect -20483 -7529 -20448 -7458
rect -17043 -7504 -16987 -7244
rect -7915 -7344 -7516 3317
rect -7915 -7410 -7898 -7344
rect -7838 -7345 -7516 -7344
rect -7838 -7410 -7743 -7345
rect -7915 -7411 -7743 -7410
rect -7683 -7411 -7610 -7345
rect -7550 -7411 -7516 -7345
rect -20587 -11503 -20448 -7529
rect -19863 -8232 -19578 -8199
rect -19863 -8314 -19850 -8232
rect -19768 -8314 -19685 -8232
rect -19603 -8314 -19578 -8232
rect -19863 -8352 -19578 -8314
rect -16994 -9856 -16937 -9593
rect -19420 -10027 -19362 -9917
rect -19456 -10787 -19346 -10027
rect -20036 -10827 -19346 -10787
rect -20036 -10982 -20018 -10827
rect -19863 -10829 -19346 -10827
rect -19863 -10982 -19686 -10829
rect -19533 -10978 -19346 -10829
rect -19533 -10982 -19434 -10978
rect -20036 -11012 -19434 -10982
rect -20587 -11618 -20562 -11503
rect -20476 -11618 -20448 -11503
rect -20587 -11704 -20448 -11618
rect -20587 -11819 -20565 -11704
rect -20479 -11819 -20448 -11704
rect -20587 -11849 -20448 -11819
rect -11113 -11377 -11005 -11321
rect -11113 -11472 -11090 -11377
rect -11013 -11472 -11005 -11377
rect -11113 -11553 -11005 -11472
rect -11113 -11648 -11093 -11553
rect -11016 -11648 -11005 -11553
rect -11113 -11712 -11005 -11648
rect -11113 -11807 -11091 -11712
rect -11014 -11807 -11005 -11712
rect -11113 -11870 -11005 -11807
rect -11113 -11965 -11092 -11870
rect -11015 -11965 -11005 -11870
rect -23397 -13611 -23091 -13606
rect -23397 -13614 -23248 -13611
rect -23397 -13695 -23388 -13614
rect -23327 -13692 -23248 -13614
rect -23187 -13687 -23091 -13611
rect -23030 -13687 -22998 -13606
rect -23187 -13692 -22998 -13687
rect -23327 -13695 -22998 -13692
rect -23397 -17377 -22998 -13695
rect -18626 -12060 -18480 -12006
rect -18626 -12176 -18597 -12060
rect -18509 -12176 -18480 -12060
rect -18626 -12289 -18480 -12176
rect -18626 -12405 -18596 -12289
rect -18508 -12405 -18480 -12289
rect -18626 -15808 -18480 -12405
rect -11316 -12396 -11211 -12381
rect -11316 -12422 -11208 -12396
rect -11316 -12517 -11291 -12422
rect -11214 -12517 -11208 -12422
rect -11316 -12598 -11208 -12517
rect -11316 -12693 -11294 -12598
rect -11217 -12693 -11208 -12598
rect -11316 -12757 -11208 -12693
rect -11316 -12852 -11292 -12757
rect -11215 -12852 -11208 -12757
rect -11316 -12915 -11208 -12852
rect -11316 -13010 -11293 -12915
rect -11216 -13010 -11208 -12915
rect -11316 -13033 -11208 -13010
rect -11316 -14153 -11211 -13033
rect -11113 -14021 -11005 -11965
rect -7915 -14459 -7516 -7411
rect -7915 -14546 -7903 -14459
rect -7831 -14546 -7762 -14459
rect -7690 -14460 -7516 -14459
rect -7690 -14546 -7624 -14460
rect -7915 -14547 -7624 -14546
rect -7552 -14547 -7516 -14460
rect -17864 -15072 -17777 -15051
rect -17864 -15128 -17851 -15072
rect -17795 -15128 -17777 -15072
rect -17864 -15183 -17777 -15128
rect -17864 -15239 -17855 -15183
rect -17799 -15239 -17777 -15183
rect -17864 -15254 -17777 -15239
rect -15570 -15800 -15514 -15533
rect -18626 -15909 -18605 -15808
rect -18507 -15909 -18480 -15808
rect -18626 -16003 -18480 -15909
rect -18626 -16104 -18600 -16003
rect -18502 -16104 -18480 -16003
rect -18626 -16133 -18480 -16104
rect -15567 -16256 -15511 -15989
rect -18454 -16969 -18169 -16936
rect -18454 -17051 -18441 -16969
rect -18359 -17051 -18276 -16969
rect -18194 -17051 -18169 -16969
rect -18454 -17089 -18169 -17051
rect -23397 -17382 -23120 -17377
rect -23397 -17444 -23388 -17382
rect -23331 -17444 -23268 -17382
rect -23211 -17439 -23120 -17382
rect -23063 -17439 -22998 -17377
rect -23211 -17444 -22998 -17439
rect -23397 -19009 -22998 -17444
rect -18423 -18319 -18107 -18285
rect -18423 -18320 -18206 -18319
rect -18423 -18381 -18383 -18320
rect -18329 -18380 -18206 -18320
rect -18152 -18380 -18107 -18319
rect -18329 -18381 -18107 -18380
rect -18423 -18410 -18107 -18381
rect -23397 -19011 -23101 -19009
rect -23397 -19015 -23259 -19011
rect -23397 -19097 -23384 -19015
rect -23321 -19093 -23259 -19015
rect -23196 -19091 -23101 -19011
rect -23038 -19091 -22998 -19009
rect -23196 -19093 -22998 -19091
rect -23321 -19097 -22998 -19093
rect -23397 -21674 -22998 -19097
rect -18232 -19604 -18107 -18410
rect -15518 -18587 -15461 -18354
rect -11159 -19445 -11051 -19415
rect -11160 -19471 -11051 -19445
rect -11160 -19566 -11142 -19471
rect -11065 -19566 -11051 -19471
rect -18352 -19620 -18003 -19604
rect -18352 -19622 -18124 -19620
rect -18352 -19727 -18343 -19622
rect -18238 -19727 -18124 -19622
rect -18017 -19727 -18003 -19620
rect -18352 -19741 -18003 -19727
rect -11160 -19647 -11051 -19566
rect -11160 -19742 -11145 -19647
rect -11068 -19742 -11051 -19647
rect -11160 -19806 -11051 -19742
rect -11160 -19901 -11143 -19806
rect -11066 -19901 -11051 -19806
rect -11160 -19964 -11051 -19901
rect -11160 -20059 -11144 -19964
rect -11067 -20059 -11051 -19964
rect -11160 -20082 -11051 -20059
rect -11362 -20487 -11257 -20459
rect -11363 -20513 -11257 -20487
rect -18588 -20558 -18225 -20537
rect -18588 -20559 -18336 -20558
rect -18588 -20651 -18560 -20559
rect -18468 -20651 -18336 -20559
rect -18588 -20652 -18336 -20651
rect -18242 -20652 -18225 -20558
rect -18588 -20667 -18225 -20652
rect -11363 -20608 -11345 -20513
rect -11268 -20608 -11257 -20513
rect -18881 -20840 -18754 -20809
rect -18881 -20932 -18864 -20840
rect -18772 -20932 -18754 -20840
rect -23397 -21766 -23388 -21674
rect -23320 -21679 -22998 -21674
rect -23320 -21766 -23233 -21679
rect -23397 -21771 -23233 -21766
rect -23165 -21680 -22998 -21679
rect -23165 -21771 -23086 -21680
rect -23397 -21772 -23086 -21771
rect -23018 -21772 -22998 -21680
rect -23397 -25351 -22998 -21772
rect -23397 -25358 -23106 -25351
rect -23397 -25361 -23250 -25358
rect -23397 -25448 -23383 -25361
rect -23323 -25445 -23250 -25361
rect -23190 -25438 -23106 -25358
rect -23046 -25438 -22998 -25351
rect -23190 -25445 -22998 -25438
rect -23323 -25448 -22998 -25445
rect -23397 -26606 -22998 -25448
rect -23397 -26698 -23390 -26606
rect -23322 -26613 -22998 -26606
rect -23322 -26698 -23225 -26613
rect -23397 -26705 -23225 -26698
rect -23157 -26705 -23080 -26613
rect -23012 -26705 -22998 -26613
rect -23397 -29982 -22998 -26705
rect -19162 -21066 -19067 -21042
rect -19162 -21136 -19142 -21066
rect -19087 -21136 -19067 -21066
rect -19162 -21229 -19067 -21136
rect -19162 -21299 -19140 -21229
rect -19085 -21299 -19067 -21229
rect -19162 -21333 -19067 -21299
rect -18881 -21064 -18754 -20932
rect -18881 -21158 -18865 -21064
rect -18771 -21158 -18754 -21064
rect -19162 -23981 -19070 -21333
rect -19162 -24048 -19149 -23981
rect -19082 -24048 -19070 -23981
rect -19162 -24171 -19070 -24048
rect -19162 -24238 -19154 -24171
rect -19087 -24238 -19070 -24171
rect -19162 -27877 -19070 -24238
rect -18881 -26115 -18754 -21158
rect -18577 -25723 -18455 -20667
rect -11363 -20689 -11257 -20608
rect -11363 -20784 -11348 -20689
rect -11271 -20784 -11257 -20689
rect -11363 -20848 -11257 -20784
rect -11363 -20943 -11346 -20848
rect -11269 -20943 -11257 -20848
rect -11363 -21006 -11257 -20943
rect -11363 -21101 -11347 -21006
rect -11270 -21101 -11257 -21006
rect -11363 -21124 -11257 -21101
rect -11362 -21968 -11257 -21124
rect -11159 -21945 -11051 -20082
rect -17905 -23001 -17818 -22980
rect -17905 -23057 -17892 -23001
rect -17836 -23057 -17818 -23001
rect -17905 -23112 -17818 -23057
rect -17905 -23168 -17896 -23112
rect -17840 -23168 -17818 -23112
rect -17905 -23183 -17818 -23168
rect -15616 -23769 -15560 -23538
rect -15606 -24244 -15550 -24031
rect -7915 -24134 -7516 -14547
rect -7915 -24190 -7900 -24134
rect -7848 -24135 -7663 -24134
rect -7848 -24190 -7785 -24135
rect -7915 -24191 -7785 -24190
rect -7733 -24190 -7663 -24135
rect -7611 -24190 -7516 -24134
rect -7733 -24191 -7516 -24190
rect -18293 -24854 -18140 -24841
rect -18293 -24936 -18255 -24854
rect -18173 -24936 -18140 -24854
rect -18293 -25019 -18140 -24936
rect -18293 -25101 -18255 -25019
rect -18173 -25101 -18140 -25019
rect -18293 -25126 -18140 -25101
rect -18577 -25845 -17913 -25723
rect -18881 -26192 -18858 -26115
rect -18781 -26192 -18754 -26115
rect -18881 -26290 -18754 -26192
rect -18881 -26365 -18858 -26290
rect -18783 -26365 -18754 -26290
rect -18881 -26371 -18754 -26365
rect -18879 -26393 -18765 -26371
rect -15564 -26564 -15507 -26333
rect -19162 -27939 -19151 -27877
rect -19083 -27939 -19070 -27877
rect -19162 -28043 -19070 -27939
rect -19162 -28105 -19151 -28043
rect -19083 -28105 -19070 -28043
rect -19162 -28117 -19070 -28105
rect -11202 -27513 -11094 -27447
rect -11202 -27608 -11180 -27513
rect -11103 -27608 -11094 -27513
rect -11202 -27689 -11094 -27608
rect -11202 -27784 -11183 -27689
rect -11106 -27784 -11094 -27689
rect -11202 -27848 -11094 -27784
rect -11202 -27943 -11181 -27848
rect -11104 -27943 -11094 -27848
rect -11202 -28006 -11094 -27943
rect -11202 -28101 -11182 -28006
rect -11105 -28101 -11094 -28006
rect -19407 -28215 -19311 -28168
rect -19407 -28274 -19388 -28215
rect -19326 -28274 -19311 -28215
rect -19407 -28380 -19311 -28274
rect -19407 -28439 -19391 -28380
rect -19329 -28439 -19311 -28380
rect -19407 -28528 -19311 -28439
rect -23397 -29984 -23092 -29982
rect -23397 -29990 -23232 -29984
rect -23397 -30075 -23386 -29990
rect -23320 -30069 -23232 -29990
rect -23166 -30067 -23092 -29984
rect -23026 -30067 -22998 -29982
rect -23166 -30069 -22998 -30067
rect -23320 -30075 -22998 -30069
rect -23397 -33381 -22998 -30075
rect -19400 -31818 -19311 -28528
rect -18977 -28505 -18880 -28494
rect -18977 -28580 -18955 -28505
rect -18890 -28580 -18880 -28505
rect -18977 -28699 -18880 -28580
rect -18977 -28714 -18961 -28699
rect -18979 -28774 -18961 -28714
rect -18896 -28774 -18880 -28699
rect -18979 -28794 -18880 -28774
rect -11405 -28551 -11300 -28509
rect -11405 -28646 -11386 -28551
rect -11309 -28646 -11300 -28551
rect -11405 -28727 -11300 -28646
rect -23397 -33384 -23248 -33381
rect -23397 -33447 -23380 -33384
rect -23320 -33444 -23248 -33384
rect -23188 -33384 -22998 -33381
rect -23188 -33444 -23114 -33384
rect -23320 -33447 -23114 -33444
rect -23054 -33447 -22998 -33384
rect -23397 -34906 -22998 -33447
rect -23397 -34909 -23087 -34906
rect -23397 -34911 -23236 -34909
rect -23397 -34995 -23389 -34911
rect -23317 -34993 -23236 -34911
rect -23164 -34990 -23087 -34909
rect -23015 -34990 -22998 -34906
rect -23164 -34993 -22998 -34990
rect -23317 -34995 -22998 -34993
rect -23397 -36500 -22998 -34995
rect -19419 -31953 -19291 -31818
rect -19419 -32014 -19382 -31953
rect -19329 -32014 -19291 -31953
rect -19419 -32112 -19291 -32014
rect -19419 -32173 -19384 -32112
rect -19331 -32173 -19291 -32112
rect -23400 -36517 -22990 -36500
rect -23400 -36520 -23073 -36517
rect -23400 -36525 -23222 -36520
rect -23400 -36620 -23381 -36525
rect -23304 -36615 -23222 -36525
rect -23145 -36612 -23073 -36520
rect -22996 -36612 -22990 -36517
rect -23145 -36615 -22990 -36612
rect -23304 -36620 -22990 -36615
rect -23400 -36693 -22990 -36620
rect -23400 -36696 -23076 -36693
rect -23400 -36701 -23225 -36696
rect -23400 -36796 -23384 -36701
rect -23307 -36791 -23225 -36701
rect -23148 -36788 -23076 -36696
rect -22999 -36788 -22990 -36693
rect -23148 -36791 -22990 -36788
rect -23307 -36796 -22990 -36791
rect -23400 -36852 -22990 -36796
rect -19419 -36830 -19291 -32173
rect -18979 -34196 -18882 -28794
rect -11405 -28822 -11389 -28727
rect -11312 -28822 -11300 -28727
rect -11405 -28886 -11300 -28822
rect -18692 -28987 -18596 -28960
rect -18692 -29054 -18667 -28987
rect -18602 -29054 -18596 -28987
rect -18692 -29067 -18596 -29054
rect -11405 -28981 -11387 -28886
rect -11310 -28981 -11300 -28886
rect -11405 -29044 -11300 -28981
rect -18692 -29175 -18594 -29067
rect -18692 -29242 -18681 -29175
rect -18616 -29242 -18594 -29175
rect -18692 -29259 -18594 -29242
rect -18690 -33763 -18594 -29259
rect -11405 -29139 -11388 -29044
rect -11311 -29139 -11300 -29044
rect -11405 -29973 -11300 -29139
rect -11202 -29993 -11094 -28101
rect -7915 -30739 -7516 -24191
rect -7915 -30742 -7765 -30739
rect -7915 -30805 -7897 -30742
rect -7837 -30802 -7765 -30742
rect -7705 -30742 -7516 -30739
rect -7705 -30802 -7631 -30742
rect -7837 -30805 -7631 -30802
rect -7571 -30805 -7516 -30742
rect -7915 -31175 -7516 -30805
rect -7915 -31178 -7765 -31175
rect -7915 -31241 -7897 -31178
rect -7837 -31238 -7765 -31178
rect -7705 -31178 -7516 -31175
rect -7705 -31238 -7631 -31178
rect -7837 -31241 -7631 -31238
rect -7571 -31241 -7516 -31178
rect -15659 -31741 -15603 -31504
rect -15656 -32263 -15600 -32022
rect -18454 -33079 -18146 -33026
rect -18454 -33081 -18259 -33079
rect -18454 -33149 -18438 -33081
rect -18377 -33147 -18259 -33081
rect -18198 -33147 -18146 -33079
rect -18377 -33149 -18146 -33147
rect -18454 -33177 -18146 -33149
rect -18690 -33859 -17958 -33763
rect -18979 -34257 -18964 -34196
rect -18901 -34257 -18882 -34196
rect -18979 -34316 -18882 -34257
rect -18979 -34377 -18963 -34316
rect -18900 -34377 -18882 -34316
rect -18979 -34397 -18882 -34377
rect -15607 -34593 -15550 -34353
rect -7915 -36140 -7516 -31241
rect -7915 -36146 -7611 -36140
rect -7915 -36150 -7758 -36146
rect -7915 -36231 -7898 -36150
rect -7842 -36227 -7758 -36150
rect -7702 -36221 -7611 -36146
rect -7555 -36221 -7516 -36140
rect -7702 -36227 -7516 -36221
rect -7842 -36231 -7516 -36227
rect -23400 -36855 -23074 -36852
rect -23400 -36860 -23223 -36855
rect -23400 -36955 -23382 -36860
rect -23305 -36950 -23223 -36860
rect -23146 -36947 -23074 -36855
rect -22997 -36947 -22990 -36852
rect -23146 -36950 -22990 -36947
rect -23305 -36955 -22990 -36950
rect -23400 -37010 -22990 -36955
rect -23400 -37013 -23075 -37010
rect -23400 -37018 -23224 -37013
rect -23400 -37113 -23383 -37018
rect -23306 -37108 -23224 -37018
rect -23147 -37105 -23075 -37013
rect -22998 -37105 -22990 -37010
rect -19584 -36884 -19260 -36830
rect -19584 -36895 -19388 -36884
rect -19584 -36980 -19550 -36895
rect -19493 -36969 -19388 -36895
rect -19331 -36969 -19260 -36884
rect -19493 -36980 -19260 -36969
rect -19584 -37033 -19260 -36980
rect -23147 -37108 -22990 -37105
rect -23306 -37113 -22990 -37108
rect -23400 -37125 -22990 -37113
rect -24190 -37549 -23779 -37532
rect -24190 -37552 -23862 -37549
rect -24190 -37557 -24011 -37552
rect -24190 -37652 -24170 -37557
rect -24093 -37647 -24011 -37557
rect -23934 -37644 -23862 -37552
rect -23785 -37644 -23779 -37549
rect -23934 -37647 -23779 -37644
rect -24093 -37652 -23779 -37647
rect -24190 -37725 -23779 -37652
rect -24190 -37728 -23865 -37725
rect -24190 -37733 -24014 -37728
rect -24190 -37828 -24173 -37733
rect -24096 -37823 -24014 -37733
rect -23937 -37820 -23865 -37728
rect -23788 -37820 -23779 -37725
rect -23937 -37823 -23779 -37820
rect -24096 -37828 -23779 -37823
rect -24190 -37884 -23779 -37828
rect -24190 -37887 -23863 -37884
rect -24190 -37892 -24012 -37887
rect -24190 -37987 -24171 -37892
rect -24094 -37982 -24012 -37892
rect -23935 -37979 -23863 -37887
rect -23786 -37979 -23779 -37884
rect -23935 -37982 -23779 -37979
rect -24094 -37987 -23779 -37982
rect -24190 -38042 -23779 -37987
rect -24190 -38045 -23864 -38042
rect -24190 -38050 -24013 -38045
rect -24190 -38145 -24172 -38050
rect -24095 -38140 -24013 -38050
rect -23936 -38137 -23864 -38045
rect -23787 -38137 -23779 -38042
rect -23936 -38140 -23779 -38137
rect -24095 -38145 -23779 -38140
rect -24190 -38157 -23779 -38145
rect -23397 -37536 -22998 -37125
rect -23397 -37538 -23089 -37536
rect -23397 -37548 -23229 -37538
rect -23397 -37633 -23380 -37548
rect -23323 -37623 -23229 -37548
rect -23172 -37621 -23089 -37538
rect -23032 -37621 -22998 -37536
rect -23172 -37623 -22998 -37621
rect -23323 -37633 -22998 -37623
rect -24190 -38313 -23791 -38157
rect -23397 -38313 -22998 -37633
rect -7915 -37536 -7516 -36231
rect -7146 51263 -6747 55224
rect 4068 54811 4467 55873
rect 4832 55849 5231 55873
rect 4832 55832 5245 55849
rect 4832 55829 5162 55832
rect 4832 55824 5013 55829
rect 4832 55729 4854 55824
rect 4931 55734 5013 55824
rect 5090 55737 5162 55829
rect 5239 55737 5245 55832
rect 5090 55734 5245 55737
rect 4931 55729 5245 55734
rect 4832 55656 5245 55729
rect 4832 55653 5159 55656
rect 4832 55648 5010 55653
rect 4832 55553 4851 55648
rect 4928 55558 5010 55648
rect 5087 55561 5159 55653
rect 5236 55561 5245 55656
rect 5087 55558 5245 55561
rect 4928 55553 5245 55558
rect 4832 55497 5245 55553
rect 4832 55494 5161 55497
rect 4832 55489 5012 55494
rect 4832 55394 4853 55489
rect 4930 55399 5012 55489
rect 5089 55402 5161 55494
rect 5238 55402 5245 55497
rect 5089 55399 5245 55402
rect 4930 55394 5245 55399
rect 4832 55339 5245 55394
rect 4832 55336 5160 55339
rect 4832 55331 5011 55336
rect 4832 55236 4852 55331
rect 4929 55241 5011 55331
rect 5088 55244 5160 55336
rect 5237 55244 5245 55339
rect 5088 55241 5245 55244
rect 4929 55236 5245 55241
rect 4832 55224 5245 55236
rect 4068 54794 4480 54811
rect 4068 54791 4397 54794
rect 4068 54786 4248 54791
rect 4068 54691 4089 54786
rect 4166 54696 4248 54786
rect 4325 54699 4397 54791
rect 4474 54699 4480 54794
rect 4325 54696 4480 54699
rect 4166 54691 4480 54696
rect 4068 54618 4480 54691
rect 4068 54615 4394 54618
rect 4068 54610 4245 54615
rect 4068 54515 4086 54610
rect 4163 54520 4245 54610
rect 4322 54523 4394 54615
rect 4471 54523 4480 54618
rect 4322 54520 4480 54523
rect 4163 54515 4480 54520
rect 4068 54459 4480 54515
rect 4068 54456 4396 54459
rect 4068 54451 4247 54456
rect 4068 54356 4088 54451
rect 4165 54361 4247 54451
rect 4324 54364 4396 54456
rect 4473 54364 4480 54459
rect 4324 54361 4480 54364
rect 4165 54356 4480 54361
rect 4068 54301 4480 54356
rect 4068 54298 4395 54301
rect 4068 54293 4246 54298
rect 4068 54198 4087 54293
rect 4164 54203 4246 54293
rect 4323 54206 4395 54298
rect 4472 54206 4480 54301
rect 4323 54203 4480 54206
rect 4164 54198 4480 54203
rect 4068 54186 4480 54198
rect 2875 53595 2983 53633
rect 2875 53500 2900 53595
rect 2977 53500 2983 53595
rect 2875 53419 2983 53500
rect 2875 53324 2897 53419
rect 2974 53324 2983 53419
rect 2875 53260 2983 53324
rect 2875 53165 2899 53260
rect 2976 53165 2983 53260
rect 2875 53102 2983 53165
rect 2875 53007 2898 53102
rect 2975 53007 2983 53102
rect 2672 52556 2777 52600
rect -4656 52449 -4553 52465
rect -4656 52373 -4639 52449
rect -4563 52373 -4553 52449
rect -4656 52251 -4553 52373
rect -4656 52173 -4640 52251
rect -4562 52173 -4553 52251
rect 2672 52461 2693 52556
rect 2770 52461 2777 52556
rect 2672 52380 2777 52461
rect 2672 52285 2690 52380
rect 2767 52285 2777 52380
rect 2672 52221 2777 52285
rect -4656 52165 -4553 52173
rect -4381 52195 -4248 52213
rect -7146 51261 -6869 51263
rect -7146 51185 -7131 51261
rect -7078 51260 -6869 51261
rect -7078 51185 -7009 51260
rect -7146 51184 -7009 51185
rect -6956 51187 -6869 51260
rect -6816 51187 -6747 51263
rect -6956 51184 -6747 51187
rect -7146 47985 -6747 51184
rect -4647 51131 -4554 52165
rect -4381 52090 -4366 52195
rect -4261 52090 -4248 52195
rect -4381 51970 -4248 52090
rect -4381 51863 -4366 51970
rect -4259 51863 -4248 51970
rect -4381 51851 -4248 51863
rect 2672 52126 2692 52221
rect 2769 52126 2777 52221
rect 2672 52063 2777 52126
rect 2672 51968 2691 52063
rect 2768 51968 2777 52063
rect -7146 47982 -6990 47985
rect -7146 47919 -7122 47982
rect -7062 47922 -6990 47982
rect -6930 47982 -6747 47985
rect -6930 47922 -6856 47982
rect -7062 47919 -6856 47922
rect -6796 47919 -6747 47982
rect -7146 47612 -6747 47919
rect -7146 47609 -6991 47612
rect -7146 47546 -7123 47609
rect -7063 47549 -6991 47609
rect -6931 47609 -6747 47612
rect -6931 47549 -6857 47609
rect -7063 47546 -6857 47549
rect -6797 47546 -6747 47609
rect -7146 47001 -6747 47546
rect -7146 46998 -6986 47001
rect -7146 46935 -7118 46998
rect -7058 46938 -6986 46998
rect -6926 46998 -6747 47001
rect -6926 46938 -6852 46998
rect -7058 46935 -6852 46938
rect -6792 46935 -6747 46998
rect -7146 46006 -6747 46935
rect -7146 46003 -6836 46006
rect -7146 45906 -7129 46003
rect -7059 45999 -6836 46003
rect -7059 45906 -6984 45999
rect -7146 45902 -6984 45906
rect -6914 45909 -6836 45999
rect -6766 45909 -6747 46006
rect -6914 45902 -6747 45909
rect -7146 42953 -6747 45902
rect -4975 48936 -4851 49035
rect -4975 48861 -4950 48936
rect -4873 48861 -4851 48936
rect -4975 48763 -4851 48861
rect -4975 48688 -4951 48763
rect -4874 48688 -4851 48763
rect -4975 45266 -4851 48688
rect -4647 46727 -4552 51131
rect -4366 47242 -4259 51851
rect 2672 51637 2777 51968
rect 2672 51581 2700 51637
rect 2755 51581 2777 51637
rect 2672 51128 2777 51581
rect 2875 51498 2983 53007
rect 2875 51442 2906 51498
rect 2961 51442 2983 51498
rect 2875 50947 2983 51442
rect -3907 50004 -3784 50018
rect -3907 49925 -3887 50004
rect -3796 49925 -3784 50004
rect -3907 49852 -3784 49925
rect -3907 49773 -3891 49852
rect -3800 49773 -3784 49852
rect -3907 49761 -3784 49773
rect -1582 49998 -1526 50000
rect -1582 49942 -1436 49998
rect -1582 49756 -1526 49942
rect -1579 48921 -1578 48975
rect -1524 48921 -1523 48975
rect -1579 48749 -1523 48921
rect 4068 48740 4467 54186
rect 4068 48737 4212 48740
rect 4068 48674 4080 48737
rect 4140 48677 4212 48737
rect 4272 48737 4467 48740
rect 4272 48677 4346 48737
rect 4140 48674 4346 48677
rect 4406 48674 4467 48737
rect -4366 47135 -3882 47242
rect -4661 46713 -4350 46727
rect -4661 46618 -4647 46713
rect -4552 46712 -4350 46713
rect -4552 46619 -4457 46712
rect -4364 46619 -4350 46712
rect -4552 46618 -4350 46619
rect -4661 46607 -4350 46618
rect -4975 45190 -4954 45266
rect -4870 45190 -4851 45266
rect -4975 45091 -4851 45190
rect -4975 45015 -4949 45091
rect -4865 45015 -4851 45091
rect -4975 44983 -4851 45015
rect -7146 42951 -6989 42953
rect -7146 42871 -7135 42951
rect -7074 42873 -6989 42951
rect -6928 42873 -6840 42953
rect -6779 42873 -6747 42953
rect -7074 42871 -6747 42873
rect -7146 38053 -6747 42871
rect -5158 44578 -5019 44623
rect -5158 44515 -5125 44578
rect -5047 44515 -5019 44578
rect -5158 44412 -5019 44515
rect -5158 44349 -5129 44412
rect -5051 44349 -5019 44412
rect -5158 42174 -5019 44349
rect -4191 44126 -3830 44141
rect -4191 44042 -4168 44126
rect -4084 44042 -3928 44126
rect -3844 44042 -3830 44126
rect -4191 44015 -3830 44042
rect -4884 43757 -4404 43783
rect -4884 43756 -4553 43757
rect -4884 43647 -4857 43756
rect -4748 43647 -4553 43756
rect -4884 43646 -4553 43647
rect -4437 43646 -4404 43757
rect -4884 43622 -4404 43646
rect -4553 42697 -4442 43622
rect -3928 43510 -3844 44015
rect -3939 43497 -3831 43510
rect -3939 43423 -3921 43497
rect -3847 43423 -3831 43497
rect -3939 43363 -3831 43423
rect -3939 43291 -3920 43363
rect -3848 43291 -3831 43363
rect -3939 43271 -3831 43291
rect -4589 42663 -4184 42697
rect -4589 42552 -4553 42663
rect -4442 42662 -4184 42663
rect -4442 42553 -4311 42662
rect -4202 42553 -4184 42662
rect -4442 42552 -4184 42553
rect -4589 42524 -4184 42552
rect -5158 42035 -4549 42174
rect -5386 38430 -5204 38442
rect -5386 38428 -5266 38430
rect -5386 38372 -5374 38428
rect -5322 38374 -5266 38428
rect -5214 38374 -5204 38430
rect -5322 38372 -5204 38374
rect -5386 38359 -5204 38372
rect -7146 38048 -6870 38053
rect -7146 38045 -6991 38048
rect -7146 37989 -7122 38045
rect -7070 37992 -6991 38045
rect -6939 37997 -6870 38048
rect -6818 37997 -6747 38053
rect -6939 37992 -6747 37997
rect -7070 37989 -6747 37992
rect -7146 34435 -6747 37989
rect -7146 34360 -7133 34435
rect -7080 34434 -6747 34435
rect -7080 34431 -6869 34434
rect -7080 34360 -7003 34431
rect -7146 34356 -7003 34360
rect -6950 34359 -6869 34431
rect -6816 34359 -6747 34434
rect -6950 34356 -6747 34359
rect -7146 30792 -6747 34356
rect -7146 30732 -7140 30792
rect -7086 30789 -6869 30792
rect -7086 30732 -7002 30789
rect -7146 30729 -7002 30732
rect -6948 30732 -6869 30789
rect -6815 30732 -6747 30792
rect -6948 30729 -6747 30732
rect -7146 25503 -6747 30729
rect -7146 25450 -7118 25503
rect -7066 25450 -6985 25503
rect -6933 25498 -6747 25503
rect -6933 25450 -6844 25498
rect -7146 25445 -6844 25450
rect -6792 25445 -6747 25498
rect -7146 21058 -6747 25445
rect -7146 21054 -6859 21058
rect -7146 21000 -7120 21054
rect -7064 21000 -6990 21054
rect -6934 21004 -6859 21054
rect -6803 21004 -6747 21058
rect -6934 21000 -6747 21004
rect -7146 17019 -6747 21000
rect -7146 17016 -6987 17019
rect -7146 16935 -7137 17016
rect -7066 16938 -6987 17016
rect -6916 17014 -6747 17019
rect -6916 16938 -6831 17014
rect -7066 16935 -6831 16938
rect -7146 16933 -6831 16935
rect -6760 16933 -6747 17014
rect -7146 13309 -6747 16933
rect -7146 13307 -6894 13309
rect -7146 13305 -7011 13307
rect -7146 13249 -7130 13305
rect -7077 13251 -7011 13305
rect -6958 13253 -6894 13307
rect -6841 13253 -6747 13309
rect -6958 13251 -6747 13253
rect -7077 13249 -6747 13251
rect -7146 11706 -6747 13249
rect -5763 27486 -5569 27509
rect -5763 27405 -5692 27486
rect -5591 27405 -5569 27486
rect -5763 27251 -5569 27405
rect -5763 27170 -5692 27251
rect -5591 27170 -5569 27251
rect -5763 14669 -5569 27170
rect -5384 26380 -5246 38359
rect -5057 37753 -4866 37787
rect -5057 37701 -5049 37753
rect -4997 37701 -4936 37753
rect -4884 37701 -4866 37753
rect -5057 37693 -4866 37701
rect -5389 26361 -5113 26380
rect -5389 26360 -5197 26361
rect -5389 26288 -5373 26360
rect -5301 26288 -5197 26360
rect -5389 26287 -5197 26288
rect -5123 26287 -5113 26361
rect -5389 26274 -5113 26287
rect -5763 14602 -5653 14669
rect -5582 14602 -5569 14669
rect -5763 14493 -5569 14602
rect -5763 14426 -5658 14493
rect -5587 14426 -5569 14493
rect -5763 12126 -5569 14426
rect -5384 19538 -5246 26274
rect -5384 19458 -5347 19538
rect -5275 19458 -5246 19538
rect -5384 19325 -5246 19458
rect -5384 19245 -5344 19325
rect -5272 19245 -5246 19325
rect -5384 12462 -5246 19245
rect -5056 24244 -4918 37693
rect -4688 35466 -4549 42035
rect 4068 41998 4467 48674
rect 4068 41995 4208 41998
rect 4068 41939 4087 41995
rect 4139 41942 4208 41995
rect 4260 41942 4322 41998
rect 4374 41942 4467 41998
rect 4139 41939 4467 41942
rect -2470 40818 -2414 40964
rect -3084 39575 -3028 39744
rect -2020 38543 -1964 38732
rect 2816 37020 2924 37046
rect 2816 36925 2839 37020
rect 2916 36925 2924 37020
rect 2816 36844 2924 36925
rect 2816 36749 2836 36844
rect 2913 36749 2924 36844
rect 2816 36685 2924 36749
rect 2816 36590 2838 36685
rect 2915 36590 2924 36685
rect 2816 36527 2924 36590
rect 2816 36432 2837 36527
rect 2914 36432 2924 36527
rect -4688 35377 -4653 35466
rect -4575 35377 -4549 35466
rect -4688 35276 -4549 35377
rect -4688 35187 -4654 35276
rect -4576 35187 -4549 35276
rect -4688 32471 -4549 35187
rect 2613 35760 2718 35799
rect 2613 35665 2631 35760
rect 2708 35665 2718 35760
rect 2613 35584 2718 35665
rect 2613 35489 2628 35584
rect 2705 35489 2718 35584
rect 2613 35425 2718 35489
rect 2613 35330 2630 35425
rect 2707 35330 2718 35425
rect 2613 35267 2718 35330
rect 2613 35172 2629 35267
rect 2706 35172 2718 35267
rect 2613 34165 2718 35172
rect 2816 34164 2924 36432
rect 4068 33485 4467 41939
rect 4068 33421 4082 33485
rect 4138 33421 4220 33485
rect 4276 33484 4467 33485
rect 4276 33421 4360 33484
rect 4068 33420 4360 33421
rect 4416 33420 4467 33484
rect -3974 33195 -3851 33209
rect -3974 33116 -3954 33195
rect -3863 33116 -3851 33195
rect -3974 33043 -3851 33116
rect -3974 32964 -3958 33043
rect -3867 32964 -3851 33043
rect -3974 32952 -3851 32964
rect -4682 32351 -4557 32471
rect -1641 32420 -1585 32633
rect -4682 32265 -4661 32351
rect -4574 32265 -4557 32351
rect -4682 32152 -4557 32265
rect -4682 32066 -4663 32152
rect -4576 32066 -4557 32152
rect -4682 32014 -4557 32066
rect -1638 32002 -1582 32152
rect -4270 31225 -4147 31239
rect -4270 31146 -4250 31225
rect -4159 31146 -4147 31225
rect -4270 31073 -4147 31146
rect -4270 30994 -4254 31073
rect -4163 30994 -4147 31073
rect -4270 30982 -4147 30994
rect -4538 29908 -4222 29931
rect -4538 29824 -4486 29908
rect -4402 29907 -4222 29908
rect -4402 29825 -4322 29907
rect -4240 29825 -4222 29907
rect -4402 29824 -4222 29825
rect -4538 29801 -4222 29824
rect -4486 28187 -4402 29801
rect -1589 29616 -1532 29834
rect -4030 28762 -3919 29397
rect -4055 28742 -3896 28762
rect -4055 28631 -4030 28742
rect -3919 28631 -3896 28742
rect -4055 28531 -3896 28631
rect -4055 28422 -4030 28531
rect -3921 28422 -3896 28531
rect -4055 28402 -3896 28422
rect -4497 28170 -4388 28187
rect -4497 28086 -4486 28170
rect -4402 28086 -4388 28170
rect -4497 28005 -4388 28086
rect -4497 27923 -4485 28005
rect -4403 27923 -4388 28005
rect -4497 27906 -4388 27923
rect 4068 25499 4467 33420
rect 4068 25496 4374 25499
rect 4068 25493 4224 25496
rect 4068 25427 4084 25493
rect 4150 25430 4224 25493
rect 4290 25433 4374 25496
rect 4440 25433 4467 25499
rect 4290 25430 4467 25433
rect 4150 25427 4467 25430
rect -5056 24230 -4677 24244
rect -5056 24119 -5043 24230
rect -4932 24229 -4677 24230
rect -4932 24120 -4794 24229
rect -4685 24120 -4677 24229
rect -4932 24119 -4677 24120
rect -5056 24106 -4677 24119
rect -5056 19748 -4918 24106
rect -3565 23805 -3509 23949
rect -4179 22583 -4123 22701
rect -3115 21539 -3059 21736
rect -4829 21413 -4509 21470
rect -4829 21408 -4636 21413
rect -4829 21344 -4813 21408
rect -4751 21349 -4636 21408
rect -4574 21349 -4509 21413
rect -4751 21344 -4509 21349
rect -4829 21294 -4509 21344
rect -4669 20241 -4533 21294
rect -3870 20680 -3670 20790
rect -4832 20177 -4520 20241
rect -4832 20124 -4796 20177
rect -4740 20175 -4520 20177
rect -4740 20124 -4649 20175
rect -4832 20122 -4649 20124
rect -4593 20122 -4520 20175
rect -4832 20056 -4520 20122
rect -4832 20053 -4521 20056
rect -5056 19668 -5026 19748
rect -4954 19668 -4918 19748
rect -5056 19547 -4918 19668
rect -5056 19467 -5023 19547
rect -4951 19467 -4918 19547
rect -5056 12985 -4918 19467
rect 2990 19416 3098 19446
rect 2990 19321 3012 19416
rect 3089 19321 3098 19416
rect 2990 19240 3098 19321
rect 2990 19145 3009 19240
rect 3086 19145 3098 19240
rect 2990 19081 3098 19145
rect 2990 18986 3011 19081
rect 3088 18986 3098 19081
rect 2990 18923 3098 18986
rect 2990 18828 3010 18923
rect 3087 18828 3098 18923
rect 2787 18359 2892 18368
rect 2787 18333 2893 18359
rect 2787 18238 2810 18333
rect 2887 18238 2893 18333
rect 2787 18157 2893 18238
rect 2787 18062 2807 18157
rect 2884 18062 2893 18157
rect 2787 17998 2893 18062
rect 2787 17903 2809 17998
rect 2886 17903 2893 17998
rect 2787 17840 2893 17903
rect 2787 17745 2808 17840
rect 2885 17745 2893 17840
rect 2787 17722 2893 17745
rect 2787 16744 2892 17722
rect 2990 16678 3098 18828
rect 4068 15982 4467 25427
rect 4068 15980 4372 15982
rect 4068 15914 4083 15980
rect 4144 15979 4372 15980
rect 4144 15914 4230 15979
rect 4068 15913 4230 15914
rect 4291 15916 4372 15979
rect 4433 15916 4467 15982
rect 4291 15913 4467 15916
rect -3768 15668 -3681 15689
rect -3768 15612 -3755 15668
rect -3699 15612 -3681 15668
rect -3768 15557 -3681 15612
rect -3768 15501 -3759 15557
rect -3703 15501 -3681 15557
rect -3768 15486 -3681 15501
rect -1467 14955 -1411 15123
rect -1464 14451 -1408 14703
rect -4111 13741 -4024 13762
rect -4111 13685 -4098 13741
rect -4042 13685 -4024 13741
rect -4111 13630 -4024 13685
rect -4111 13574 -4102 13630
rect -4046 13574 -4024 13630
rect -4111 13559 -4024 13574
rect -5056 12847 -3759 12985
rect -4385 12462 -4074 12463
rect -5384 12413 -4074 12462
rect -5384 12405 -4183 12413
rect -5384 12342 -4360 12405
rect -4303 12350 -4183 12405
rect -4126 12350 -4074 12413
rect -4303 12342 -4074 12350
rect -5384 12324 -4074 12342
rect -4385 12311 -4074 12324
rect -5763 11904 -5524 12126
rect -1415 12110 -1358 12349
rect -7146 11700 -6988 11706
rect -7146 11601 -7136 11700
rect -7068 11607 -6988 11700
rect -6920 11698 -6747 11706
rect -6920 11607 -6843 11698
rect -7068 11601 -6843 11607
rect -7146 11599 -6843 11601
rect -6775 11599 -6747 11698
rect -7146 9233 -6747 11599
rect -7146 9230 -6832 9233
rect -7146 9226 -6984 9230
rect -7146 9144 -7125 9226
rect -7059 9148 -6984 9226
rect -6918 9151 -6832 9230
rect -6766 9151 -6747 9233
rect -6918 9148 -6747 9151
rect -7059 9144 -6747 9148
rect -7146 4059 -6747 9144
rect -7146 3962 -7124 4059
rect -7056 3962 -6971 4059
rect -6903 3962 -6827 4059
rect -6759 3962 -6747 4059
rect -7146 3862 -6747 3962
rect -7146 3858 -6826 3862
rect -7146 3761 -7135 3858
rect -7067 3855 -6826 3858
rect -7067 3761 -6970 3855
rect -7146 3758 -6970 3761
rect -6902 3765 -6826 3855
rect -6758 3765 -6747 3862
rect -6902 3758 -6747 3765
rect -7146 638 -6747 3758
rect -5713 2170 -5524 11904
rect 3030 7417 3131 7418
rect 3023 7392 3131 7417
rect 3023 7297 3048 7392
rect 3125 7297 3131 7392
rect 3023 7216 3131 7297
rect 3023 7121 3045 7216
rect 3122 7121 3131 7216
rect 3023 7057 3131 7121
rect 3023 6962 3047 7057
rect 3124 6962 3131 7057
rect 3023 6899 3131 6962
rect 3023 6804 3046 6899
rect 3123 6804 3131 6899
rect 2820 6181 2925 6185
rect 2820 6155 2926 6181
rect 2820 6060 2843 6155
rect 2920 6060 2926 6155
rect 2820 5979 2926 6060
rect 2820 5884 2840 5979
rect 2917 5884 2926 5979
rect 2820 5820 2926 5884
rect 2820 5725 2842 5820
rect 2919 5725 2926 5820
rect 2820 5662 2926 5725
rect 2820 5567 2841 5662
rect 2918 5567 2926 5662
rect 2820 5544 2926 5567
rect 2820 3989 2925 5544
rect 3023 3904 3131 6804
rect 4068 3601 4467 15913
rect 4068 3599 4360 3601
rect 4068 3529 4084 3599
rect 4156 3529 4235 3599
rect 4307 3531 4360 3599
rect 4432 3531 4467 3601
rect 4307 3529 4467 3531
rect -3720 2975 -3633 2996
rect -3720 2919 -3707 2975
rect -3651 2919 -3633 2975
rect -3720 2864 -3633 2919
rect -3720 2808 -3711 2864
rect -3655 2808 -3633 2864
rect -3720 2793 -3633 2808
rect -1434 2237 -1378 2558
rect -5713 2080 -5520 2170
rect -5713 2008 -5650 2080
rect -5581 2008 -5520 2080
rect -5713 1907 -5520 2008
rect -5713 1835 -5656 1907
rect -5587 1835 -5520 1907
rect -5713 1790 -5520 1835
rect -7146 636 -6980 638
rect -7146 568 -7126 636
rect -7065 570 -6980 636
rect -6919 570 -6841 638
rect -6780 570 -6747 638
rect -7065 568 -6747 570
rect -7146 -1212 -6747 568
rect -7146 -1214 -6989 -1212
rect -7146 -1293 -7133 -1214
rect -7071 -1291 -6989 -1214
rect -6927 -1213 -6747 -1212
rect -6927 -1291 -6857 -1213
rect -7071 -1292 -6857 -1291
rect -6795 -1292 -6747 -1213
rect -7071 -1293 -6747 -1292
rect -7146 -4924 -6747 -1293
rect -7146 -4925 -6992 -4924
rect -7146 -4980 -7128 -4925
rect -7073 -4979 -6992 -4925
rect -6937 -4925 -6747 -4924
rect -6937 -4979 -6838 -4925
rect -7073 -4980 -6838 -4979
rect -6783 -4980 -6747 -4925
rect -7146 -8557 -6747 -4980
rect -7146 -8565 -6841 -8557
rect -7146 -8631 -7135 -8565
rect -7074 -8631 -6998 -8565
rect -6937 -8623 -6841 -8565
rect -6780 -8623 -6747 -8557
rect -6937 -8631 -6747 -8623
rect -7146 -10190 -6747 -8631
rect -7146 -10197 -6861 -10190
rect -7146 -10198 -7002 -10197
rect -7146 -10276 -7136 -10198
rect -7081 -10275 -7002 -10198
rect -6947 -10268 -6861 -10197
rect -6806 -10268 -6747 -10190
rect -6947 -10275 -6747 -10268
rect -7081 -10276 -6747 -10275
rect -7146 -13688 -6747 -10276
rect -7146 -13752 -7132 -13688
rect -7080 -13692 -6827 -13688
rect -7080 -13752 -6994 -13692
rect -7146 -13756 -6994 -13752
rect -6942 -13752 -6827 -13692
rect -6775 -13752 -6747 -13688
rect -6942 -13756 -6747 -13752
rect -7146 -17226 -6747 -13756
rect -5681 -12721 -5520 1790
rect -1431 1761 -1375 2003
rect -4084 1040 -3997 1061
rect -4084 984 -4071 1040
rect -4015 984 -3997 1040
rect -4084 929 -3997 984
rect -4084 873 -4075 929
rect -4019 873 -3997 929
rect -4084 858 -3997 873
rect -4388 -240 -3891 -216
rect -4388 -378 -4368 -240
rect -4230 -241 -3891 -240
rect -4230 -377 -4045 -241
rect -3909 -377 -3891 -241
rect -4230 -378 -3891 -377
rect -4388 -392 -3891 -378
rect -4368 -10143 -4230 -392
rect -1382 -589 -1325 -333
rect -4102 -896 -3727 -758
rect -4102 -9449 -3964 -896
rect -3759 -3926 -3510 -3919
rect -3759 -3937 -3501 -3926
rect -3759 -3940 -3584 -3937
rect -3759 -3993 -3711 -3940
rect -3659 -3990 -3584 -3940
rect -3532 -3990 -3501 -3937
rect -3659 -3993 -3501 -3990
rect -3759 -4025 -3501 -3993
rect -3564 -5158 -3501 -4025
rect -3577 -5175 -3487 -5158
rect -3577 -5228 -3552 -5175
rect -3500 -5228 -3487 -5175
rect -3577 -5290 -3487 -5228
rect -3577 -5343 -3566 -5290
rect -3514 -5343 -3487 -5290
rect -3577 -5354 -3487 -5343
rect -2108 -5645 -2052 -5458
rect 4068 -5977 4467 3529
rect 4068 -5979 4369 -5977
rect 4068 -6052 4082 -5979
rect 4161 -5980 4369 -5979
rect 4161 -6052 4231 -5980
rect 4068 -6053 4231 -6052
rect 4310 -6050 4369 -5980
rect 4448 -6050 4467 -5977
rect 4310 -6053 4467 -6050
rect -3172 -6696 -3116 -6576
rect -2558 -7885 -2502 -7737
rect -4102 -9451 -3692 -9449
rect -4102 -9471 -3434 -9451
rect -4102 -9481 -3827 -9471
rect -4102 -9571 -4065 -9481
rect -3984 -9561 -3827 -9481
rect -3746 -9561 -3434 -9471
rect -3984 -9571 -3434 -9561
rect -4102 -9589 -3434 -9571
rect -4102 -9822 -3964 -9589
rect -4102 -9960 -3300 -9822
rect -4622 -10162 -4230 -10143
rect -4622 -10204 -3738 -10162
rect -4622 -10205 -4047 -10204
rect -4622 -10277 -4274 -10205
rect -4202 -10277 -4047 -10205
rect -4622 -10278 -4047 -10277
rect -3973 -10205 -3738 -10204
rect -3973 -10277 -3844 -10205
rect -3772 -10277 -3738 -10205
rect -3973 -10278 -3738 -10277
rect -4622 -10281 -3738 -10278
rect -5681 -12772 -5517 -12721
rect -5681 -12870 -5637 -12772
rect -5540 -12870 -5517 -12772
rect -5681 -13002 -5517 -12870
rect -5681 -13100 -5645 -13002
rect -5548 -13100 -5517 -13002
rect -5681 -13119 -5517 -13100
rect -5681 -15818 -5520 -13119
rect -5681 -15871 -5589 -15818
rect -5532 -15871 -5520 -15818
rect -5681 -15937 -5520 -15871
rect -5681 -15990 -5594 -15937
rect -5537 -15990 -5520 -15937
rect -5681 -16050 -5520 -15990
rect -5681 -16103 -5592 -16050
rect -5535 -16103 -5520 -16050
rect -5681 -16255 -5520 -16103
rect -7146 -17229 -6871 -17226
rect -7146 -17230 -7005 -17229
rect -7146 -17295 -7135 -17230
rect -7080 -17294 -7005 -17230
rect -6950 -17291 -6871 -17229
rect -6816 -17291 -6747 -17226
rect -6950 -17294 -6747 -17291
rect -7080 -17295 -6747 -17294
rect -7146 -18950 -6747 -17295
rect -7146 -18955 -6833 -18950
rect -7146 -18963 -6992 -18955
rect -7146 -19027 -7129 -18963
rect -7077 -19019 -6992 -18963
rect -6940 -19014 -6833 -18955
rect -6781 -19014 -6747 -18950
rect -6940 -19019 -6747 -19014
rect -7077 -19027 -6747 -19019
rect -7146 -21670 -6747 -19027
rect -5606 -20120 -5520 -16255
rect -5606 -20172 -5590 -20120
rect -5533 -20172 -5520 -20120
rect -5606 -20256 -5520 -20172
rect -5606 -20308 -5593 -20256
rect -5536 -20308 -5520 -20256
rect -5606 -20326 -5520 -20308
rect -5312 -14862 -5178 -14815
rect -5312 -14941 -5277 -14862
rect -5207 -14941 -5178 -14862
rect -5312 -15045 -5178 -14941
rect -5312 -15124 -5281 -15045
rect -5211 -15124 -5178 -15045
rect -7146 -21677 -6828 -21670
rect -7146 -21679 -6975 -21677
rect -7146 -21759 -7139 -21679
rect -7079 -21757 -6975 -21679
rect -6915 -21750 -6828 -21677
rect -6768 -21750 -6747 -21670
rect -6915 -21757 -6747 -21750
rect -7079 -21759 -6747 -21757
rect -7146 -25305 -6747 -21759
rect -5312 -22845 -5178 -15124
rect -5312 -22926 -5294 -22845
rect -5194 -22926 -5178 -22845
rect -5312 -23046 -5178 -22926
rect -5312 -23127 -5295 -23046
rect -5195 -23127 -5178 -23046
rect -5312 -23145 -5178 -23127
rect -4952 -16795 -4814 -16771
rect -4952 -16859 -4920 -16795
rect -4856 -16859 -4814 -16795
rect -4952 -16943 -4814 -16859
rect -4952 -17007 -4923 -16943
rect -4859 -17007 -4814 -16943
rect -4952 -24665 -4814 -17007
rect -4953 -24701 -4802 -24665
rect -4953 -24811 -4927 -24701
rect -4830 -24811 -4802 -24701
rect -4953 -24987 -4802 -24811
rect -4953 -25097 -4929 -24987
rect -4832 -25097 -4802 -24987
rect -4953 -25126 -4802 -25097
rect -7146 -25308 -6840 -25305
rect -7146 -25370 -7135 -25308
rect -7078 -25310 -6840 -25308
rect -7078 -25370 -6999 -25310
rect -7146 -25372 -6999 -25370
rect -6942 -25367 -6840 -25310
rect -6783 -25367 -6747 -25305
rect -6942 -25372 -6747 -25367
rect -7146 -26567 -6747 -25372
rect -4622 -26064 -4484 -10281
rect -4368 -10307 -3738 -10281
rect -3438 -10520 -3300 -9960
rect -3438 -10540 -2756 -10520
rect -4622 -26121 -4581 -26064
rect -4524 -26121 -4484 -26064
rect -4622 -26203 -4484 -26121
rect -4622 -26258 -4581 -26203
rect -4526 -26258 -4484 -26203
rect -4622 -26289 -4484 -26258
rect -4318 -10561 -2756 -10540
rect -4318 -10577 -3179 -10561
rect -4318 -10662 -3402 -10577
rect -3304 -10646 -3179 -10577
rect -3081 -10646 -2936 -10561
rect -2838 -10646 -2756 -10561
rect -3304 -10662 -2756 -10646
rect -4318 -10678 -2756 -10662
rect -7146 -26572 -6866 -26567
rect -7146 -26581 -6996 -26572
rect -7146 -26637 -7135 -26581
rect -7083 -26628 -6996 -26581
rect -6944 -26623 -6866 -26572
rect -6814 -26623 -6747 -26567
rect -6944 -26628 -6747 -26623
rect -7083 -26637 -6747 -26628
rect -7146 -29684 -6747 -26637
rect -4318 -26828 -4180 -10678
rect -3438 -10686 -2756 -10678
rect 3075 -11355 3183 -11345
rect 3073 -11381 3183 -11355
rect 3073 -11476 3091 -11381
rect 3168 -11476 3183 -11381
rect 3073 -11557 3183 -11476
rect 3073 -11652 3088 -11557
rect 3165 -11652 3183 -11557
rect 3073 -11716 3183 -11652
rect 3073 -11811 3090 -11716
rect 3167 -11811 3183 -11716
rect 3073 -11874 3183 -11811
rect 3073 -11969 3089 -11874
rect 3166 -11969 3183 -11874
rect 3073 -11992 3183 -11969
rect 2872 -12396 2977 -12357
rect 2871 -12422 2977 -12396
rect 2871 -12517 2889 -12422
rect 2966 -12517 2977 -12422
rect 2871 -12598 2977 -12517
rect 2871 -12693 2886 -12598
rect 2963 -12693 2977 -12598
rect 2871 -12757 2977 -12693
rect 2871 -12852 2888 -12757
rect 2965 -12852 2977 -12757
rect 2871 -12915 2977 -12852
rect 2871 -13010 2887 -12915
rect 2964 -13010 2977 -12915
rect 2871 -13033 2977 -13010
rect 2872 -13922 2977 -13033
rect 3075 -13887 3183 -11992
rect 4068 -14435 4467 -6053
rect 4068 -14436 4214 -14435
rect 4068 -14531 4077 -14436
rect 4149 -14530 4214 -14436
rect 4286 -14530 4359 -14435
rect 4431 -14530 4467 -14435
rect 4149 -14531 4467 -14530
rect -3682 -14879 -3595 -14858
rect -3682 -14935 -3669 -14879
rect -3613 -14935 -3595 -14879
rect -3682 -14990 -3595 -14935
rect -3682 -15046 -3673 -14990
rect -3617 -15046 -3595 -14990
rect -3682 -15061 -3595 -15046
rect -1382 -15597 -1326 -15412
rect -1379 -16098 -1323 -15855
rect -4046 -16754 -3896 -16730
rect -4046 -16819 -4002 -16754
rect -3932 -16819 -3896 -16754
rect -4046 -16913 -3896 -16819
rect -4046 -16978 -4008 -16913
rect -3938 -16978 -3896 -16913
rect -4046 -16995 -3896 -16978
rect -4048 -18152 -3941 -18139
rect -4048 -18227 -4042 -18152
rect -3966 -18227 -3941 -18152
rect -4048 -18315 -3941 -18227
rect -4048 -18390 -4033 -18315
rect -3958 -18390 -3941 -18315
rect -4048 -20836 -3941 -18390
rect -1330 -18458 -1273 -18203
rect -3756 -20472 -3698 -18501
rect -3763 -20486 -3688 -20472
rect -3763 -20539 -3750 -20486
rect -3697 -20539 -3688 -20486
rect -3763 -20594 -3688 -20539
rect -3763 -20647 -3751 -20594
rect -3698 -20647 -3688 -20594
rect -3763 -20659 -3688 -20647
rect -4056 -20851 -3941 -20836
rect -4056 -20925 -4037 -20851
rect -3963 -20925 -3941 -20851
rect -4056 -21071 -3941 -20925
rect -4056 -21145 -4037 -21071
rect -3963 -21145 -3941 -21071
rect -4056 -21263 -3941 -21145
rect -4056 -21335 -4036 -21263
rect -3964 -21335 -3941 -21263
rect -4056 -21372 -3941 -21335
rect -3756 -21861 -3698 -20659
rect -3767 -21882 -3670 -21861
rect -3767 -21940 -3754 -21882
rect -3696 -21940 -3670 -21882
rect -3767 -21996 -3670 -21940
rect -3767 -22054 -3756 -21996
rect -3698 -22054 -3670 -21996
rect -3767 -22086 -3670 -22054
rect 4068 -22657 4467 -14531
rect 4068 -22659 4361 -22657
rect 4068 -22662 4232 -22659
rect 4068 -22718 4094 -22662
rect 4146 -22715 4232 -22662
rect 4284 -22713 4361 -22659
rect 4413 -22713 4467 -22657
rect 4284 -22715 4467 -22713
rect 4146 -22718 4467 -22715
rect 4068 -23094 4467 -22718
rect 4068 -23096 4360 -23094
rect 4068 -23099 4231 -23096
rect 4068 -23155 4093 -23099
rect 4145 -23152 4231 -23099
rect 4283 -23150 4360 -23096
rect 4412 -23150 4467 -23094
rect 4283 -23152 4467 -23150
rect 4145 -23155 4467 -23152
rect -2514 -23825 -2458 -23663
rect -3128 -25041 -3072 -24887
rect -2064 -26086 -2008 -25903
rect -4318 -26857 -4003 -26828
rect -4318 -26860 -4151 -26857
rect -4318 -26915 -4282 -26860
rect -4227 -26912 -4151 -26860
rect -4096 -26912 -4003 -26857
rect -4227 -26915 -4003 -26912
rect -4318 -26957 -4003 -26915
rect 3160 -27487 3268 -27459
rect 3156 -27513 3268 -27487
rect 3156 -27608 3174 -27513
rect 3251 -27608 3268 -27513
rect 3156 -27689 3268 -27608
rect 3156 -27784 3171 -27689
rect 3248 -27784 3268 -27689
rect 3156 -27848 3268 -27784
rect 3156 -27943 3173 -27848
rect 3250 -27943 3268 -27848
rect -4591 -28030 -4476 -27977
rect -4591 -28106 -4570 -28030
rect -4499 -28106 -4476 -28030
rect -4591 -28255 -4476 -28106
rect 3156 -28006 3268 -27943
rect 3156 -28101 3172 -28006
rect 3249 -28101 3268 -28006
rect 3156 -28124 3268 -28101
rect -4591 -28331 -4569 -28255
rect -4498 -28331 -4476 -28255
rect -4591 -28358 -4476 -28331
rect -7146 -29685 -6879 -29684
rect -7146 -29686 -7009 -29685
rect -7146 -29783 -7135 -29686
rect -7069 -29782 -7009 -29686
rect -6943 -29781 -6879 -29685
rect -6813 -29781 -6747 -29684
rect -6943 -29782 -6747 -29781
rect -7069 -29783 -6747 -29782
rect -7146 -33485 -6747 -29783
rect -4584 -31801 -4479 -28358
rect 2957 -28529 3062 -28515
rect 2957 -28555 3063 -28529
rect 2957 -28650 2980 -28555
rect 3057 -28650 3063 -28555
rect 2957 -28731 3063 -28650
rect 2957 -28826 2977 -28731
rect 3054 -28826 3063 -28731
rect 2957 -28890 3063 -28826
rect 2957 -28985 2979 -28890
rect 3056 -28985 3063 -28890
rect 2957 -29048 3063 -28985
rect 2957 -29143 2978 -29048
rect 3055 -29143 3063 -29048
rect 2957 -29166 3063 -29143
rect 2957 -30060 3062 -29166
rect 3160 -30068 3268 -28124
rect -7146 -33488 -6996 -33485
rect -7146 -33551 -7128 -33488
rect -7068 -33548 -6996 -33488
rect -6936 -33488 -6747 -33485
rect -6936 -33548 -6862 -33488
rect -7068 -33551 -6862 -33548
rect -6802 -33551 -6747 -33488
rect -7146 -35017 -6747 -33551
rect -7146 -35021 -6842 -35017
rect -7146 -35025 -6984 -35021
rect -7146 -35114 -7137 -35025
rect -7071 -35110 -6984 -35025
rect -6918 -35106 -6842 -35021
rect -6776 -35106 -6747 -35017
rect -6918 -35110 -6747 -35106
rect -7071 -35114 -6747 -35110
rect -7146 -36500 -6747 -35114
rect -4608 -31993 -4454 -31801
rect -1297 -31841 -1241 -31551
rect -4608 -32060 -4562 -31993
rect -4493 -32060 -4454 -31993
rect -4608 -32170 -4454 -32060
rect -4608 -32237 -4568 -32170
rect -4499 -32237 -4454 -32170
rect -7146 -36517 -6734 -36500
rect -7146 -36520 -6817 -36517
rect -7146 -36525 -6966 -36520
rect -7146 -36620 -7125 -36525
rect -7048 -36615 -6966 -36525
rect -6889 -36612 -6817 -36520
rect -6740 -36612 -6734 -36517
rect -6889 -36615 -6734 -36612
rect -7048 -36620 -6734 -36615
rect -7146 -36693 -6734 -36620
rect -7146 -36696 -6820 -36693
rect -7146 -36701 -6969 -36696
rect -7146 -36796 -7128 -36701
rect -7051 -36791 -6969 -36701
rect -6892 -36788 -6820 -36696
rect -6743 -36788 -6734 -36693
rect -6892 -36791 -6734 -36788
rect -7051 -36796 -6734 -36791
rect -7146 -36852 -6734 -36796
rect -7146 -36855 -6818 -36852
rect -7146 -36860 -6967 -36855
rect -7146 -36955 -7126 -36860
rect -7049 -36950 -6967 -36860
rect -6890 -36947 -6818 -36855
rect -6741 -36947 -6734 -36852
rect -6890 -36950 -6734 -36947
rect -7049 -36955 -6734 -36950
rect -7146 -37010 -6734 -36955
rect -4608 -36958 -4454 -32237
rect -1294 -32354 -1238 -32164
rect 4068 -32591 4467 -23155
rect 4068 -32594 4220 -32591
rect 4068 -32657 4088 -32594
rect 4148 -32654 4220 -32594
rect 4280 -32594 4467 -32591
rect 4280 -32654 4354 -32594
rect 4148 -32657 4354 -32654
rect 4414 -32657 4467 -32594
rect -4136 -33092 -3864 -33047
rect -4136 -33114 -3968 -33092
rect -4136 -33175 -4122 -33114
rect -4054 -33153 -3968 -33114
rect -3900 -33153 -3864 -33092
rect -4054 -33175 -3864 -33153
rect -4136 -33200 -3864 -33175
rect -4198 -34382 -3878 -34379
rect -4198 -34404 -3874 -34382
rect -4198 -34415 -4001 -34404
rect -4198 -34513 -4166 -34415
rect -4075 -34502 -4001 -34415
rect -3910 -34502 -3874 -34404
rect -4075 -34513 -3874 -34502
rect -4198 -34540 -3874 -34513
rect -3976 -35596 -3874 -34540
rect -1245 -34691 -1188 -34461
rect -3674 -34909 -3609 -34735
rect -3694 -35541 -3588 -34909
rect -3701 -35567 -3399 -35541
rect -3701 -35569 -3515 -35567
rect -4005 -35693 -3852 -35596
rect -3701 -35637 -3675 -35569
rect -3605 -35635 -3515 -35569
rect -3445 -35635 -3399 -35567
rect -3605 -35637 -3399 -35635
rect -3701 -35667 -3399 -35637
rect -4005 -35770 -3975 -35693
rect -3883 -35770 -3852 -35693
rect -4005 -35838 -3852 -35770
rect -4005 -35935 -3985 -35838
rect -3866 -35935 -3852 -35838
rect -4005 -35959 -3852 -35935
rect 4068 -36216 4467 -32657
rect 4068 -36297 4082 -36216
rect 4138 -36297 4243 -36216
rect 4299 -36218 4467 -36216
rect 4299 -36297 4400 -36218
rect 4068 -36299 4400 -36297
rect 4456 -36299 4467 -36218
rect -7146 -37013 -6819 -37010
rect -7146 -37018 -6968 -37013
rect -7146 -37113 -7127 -37018
rect -7050 -37108 -6968 -37018
rect -6891 -37105 -6819 -37013
rect -6742 -37105 -6734 -37010
rect -6891 -37108 -6734 -37105
rect -7050 -37113 -6734 -37108
rect -7146 -37125 -6734 -37113
rect -4742 -37031 -4410 -36958
rect -4742 -37038 -4584 -37031
rect -4742 -37121 -4705 -37038
rect -4648 -37114 -4584 -37038
rect -4527 -37114 -4410 -37031
rect -4648 -37121 -4410 -37114
rect -7915 -37553 -7505 -37536
rect -7915 -37556 -7588 -37553
rect -7915 -37561 -7737 -37556
rect -7915 -37656 -7896 -37561
rect -7819 -37651 -7737 -37561
rect -7660 -37648 -7588 -37556
rect -7511 -37648 -7505 -37553
rect -7660 -37651 -7505 -37648
rect -7819 -37656 -7505 -37651
rect -7915 -37729 -7505 -37656
rect -7915 -37732 -7591 -37729
rect -7915 -37737 -7740 -37732
rect -7915 -37832 -7899 -37737
rect -7822 -37827 -7740 -37737
rect -7663 -37824 -7591 -37732
rect -7514 -37824 -7505 -37729
rect -7663 -37827 -7505 -37824
rect -7822 -37832 -7505 -37827
rect -7915 -37888 -7505 -37832
rect -7915 -37891 -7589 -37888
rect -7915 -37896 -7738 -37891
rect -7915 -37991 -7897 -37896
rect -7820 -37986 -7738 -37896
rect -7661 -37983 -7589 -37891
rect -7512 -37983 -7505 -37888
rect -7661 -37986 -7505 -37983
rect -7820 -37991 -7505 -37986
rect -7915 -38046 -7505 -37991
rect -7915 -38049 -7590 -38046
rect -7915 -38054 -7739 -38049
rect -7915 -38149 -7898 -38054
rect -7821 -38144 -7739 -38054
rect -7662 -38141 -7590 -38049
rect -7513 -38141 -7505 -38046
rect -7662 -38144 -7505 -38141
rect -7821 -38149 -7505 -38144
rect -7915 -38161 -7505 -38149
rect -7146 -37649 -6747 -37125
rect -4742 -37153 -4410 -37121
rect -7146 -37658 -6858 -37649
rect -7146 -37663 -6982 -37658
rect -7146 -37744 -7132 -37663
rect -7076 -37739 -6982 -37663
rect -6926 -37730 -6858 -37658
rect -6802 -37730 -6747 -37649
rect -6926 -37739 -6747 -37730
rect -7076 -37744 -6747 -37739
rect -7915 -38182 -7516 -38161
rect -7146 -38182 -6747 -37744
rect 4068 -37536 4467 -36299
rect 4832 51319 5231 55224
rect 14634 54809 15033 55873
rect 15320 55849 15719 55873
rect 15320 55832 15731 55849
rect 15320 55829 15648 55832
rect 15320 55824 15499 55829
rect 15320 55729 15340 55824
rect 15417 55734 15499 55824
rect 15576 55737 15648 55829
rect 15725 55737 15731 55832
rect 15576 55734 15731 55737
rect 15417 55729 15731 55734
rect 15320 55656 15731 55729
rect 15320 55653 15645 55656
rect 15320 55648 15496 55653
rect 15320 55553 15337 55648
rect 15414 55558 15496 55648
rect 15573 55561 15645 55653
rect 15722 55561 15731 55656
rect 15573 55558 15731 55561
rect 15414 55553 15731 55558
rect 15320 55497 15731 55553
rect 15320 55494 15647 55497
rect 15320 55489 15498 55494
rect 15320 55394 15339 55489
rect 15416 55399 15498 55489
rect 15575 55402 15647 55494
rect 15724 55402 15731 55497
rect 15575 55399 15731 55402
rect 15416 55394 15731 55399
rect 15320 55339 15731 55394
rect 15320 55336 15646 55339
rect 15320 55331 15497 55336
rect 15320 55236 15338 55331
rect 15415 55241 15497 55331
rect 15574 55244 15646 55336
rect 15723 55244 15731 55339
rect 15574 55241 15731 55244
rect 15415 55236 15731 55241
rect 15320 55224 15731 55236
rect 14633 54792 15043 54809
rect 14633 54789 14960 54792
rect 14633 54784 14811 54789
rect 14633 54689 14652 54784
rect 14729 54694 14811 54784
rect 14888 54697 14960 54789
rect 15037 54697 15043 54792
rect 14888 54694 15043 54697
rect 14729 54689 15043 54694
rect 14633 54616 15043 54689
rect 14633 54613 14957 54616
rect 14633 54608 14808 54613
rect 14633 54513 14649 54608
rect 14726 54518 14808 54608
rect 14885 54521 14957 54613
rect 15034 54521 15043 54616
rect 14885 54518 15043 54521
rect 14726 54513 15043 54518
rect 14633 54457 15043 54513
rect 14633 54454 14959 54457
rect 14633 54449 14810 54454
rect 14633 54354 14651 54449
rect 14728 54359 14810 54449
rect 14887 54362 14959 54454
rect 15036 54362 15043 54457
rect 14887 54359 15043 54362
rect 14728 54354 15043 54359
rect 14633 54299 15043 54354
rect 14633 54296 14958 54299
rect 14633 54291 14809 54296
rect 14633 54196 14650 54291
rect 14727 54201 14809 54291
rect 14886 54204 14958 54296
rect 15035 54204 15043 54299
rect 14886 54201 15043 54204
rect 14727 54196 15043 54201
rect 14633 54184 15043 54196
rect 6673 52463 6767 52472
rect 6502 52450 6774 52463
rect 6502 52372 6516 52450
rect 6594 52372 6681 52450
rect 6759 52372 6774 52450
rect 6502 52357 6774 52372
rect 6356 52196 6489 52215
rect 6356 52089 6370 52196
rect 6477 52089 6489 52196
rect 6356 51989 6489 52089
rect 6356 51884 6371 51989
rect 6476 51884 6489 51989
rect 6356 51868 6489 51884
rect 4832 51316 5158 51319
rect 4832 51240 4845 51316
rect 4907 51315 5158 51316
rect 4907 51240 4973 51315
rect 4832 51239 4973 51240
rect 5035 51243 5158 51315
rect 5220 51243 5231 51319
rect 5035 51239 5231 51243
rect 4832 47688 5231 51239
rect 6370 51144 6477 51868
rect 6673 51780 6767 52357
rect 6673 51770 6769 51780
rect 6672 51694 6681 51770
rect 6673 51692 6681 51694
rect 6759 51692 6769 51770
rect 6673 51606 6769 51692
rect 6673 51530 6682 51606
rect 6758 51530 6769 51606
rect 6673 51518 6769 51530
rect 6351 51129 6497 51144
rect 6351 51018 6368 51129
rect 6479 51018 6497 51129
rect 6351 50902 6497 51018
rect 6351 50793 6369 50902
rect 6478 50793 6497 50902
rect 6351 50772 6522 50793
rect 6353 50682 6522 50772
rect 4832 47685 4979 47688
rect 4832 47616 4844 47685
rect 4902 47619 4979 47685
rect 5037 47686 5231 47688
rect 5037 47619 5128 47686
rect 4902 47617 5128 47619
rect 5186 47617 5231 47686
rect 4902 47616 5231 47617
rect 4832 46294 5231 47616
rect 4832 46291 4981 46294
rect 4832 46228 4849 46291
rect 4909 46231 4981 46291
rect 5041 46291 5231 46294
rect 5041 46231 5115 46291
rect 4909 46228 5115 46231
rect 5175 46228 5231 46291
rect 4832 43020 5231 46228
rect 4832 43010 4980 43020
rect 4832 42920 4840 43010
rect 4920 42930 4980 43010
rect 5060 43010 5231 43020
rect 5060 42930 5120 43010
rect 4920 42920 5120 42930
rect 5200 42920 5231 43010
rect 4832 40595 5231 42920
rect 4832 40588 4972 40595
rect 4832 40532 4855 40588
rect 4907 40539 4972 40588
rect 5024 40592 5231 40595
rect 5024 40539 5089 40592
rect 4907 40536 5089 40539
rect 5141 40536 5231 40592
rect 4907 40532 5231 40536
rect 4832 39244 5231 40532
rect 4832 39237 4973 39244
rect 4832 39181 4856 39237
rect 4908 39188 4973 39237
rect 5025 39241 5231 39244
rect 5025 39188 5090 39241
rect 4908 39185 5090 39188
rect 5142 39185 5231 39241
rect 4908 39181 5231 39185
rect 4832 34494 5231 39181
rect 4832 34492 5137 34494
rect 4832 34423 4841 34492
rect 4906 34423 4991 34492
rect 5056 34425 5137 34492
rect 5202 34425 5231 34494
rect 5056 34423 5231 34425
rect 4832 30740 5231 34423
rect 6205 39694 6292 39734
rect 6205 39631 6222 39694
rect 6275 39631 6292 39694
rect 6205 39556 6292 39631
rect 6205 39493 6223 39556
rect 6276 39493 6292 39556
rect 6205 31131 6292 39493
rect 6415 38967 6522 50682
rect 6415 38892 6437 38967
rect 6512 38892 6522 38967
rect 6415 38796 6522 38892
rect 6415 38721 6435 38796
rect 6510 38721 6522 38796
rect 6415 38709 6522 38721
rect 6673 38541 6767 51518
rect 14634 50297 15033 54184
rect 14634 50294 14792 50297
rect 14634 50231 14660 50294
rect 14720 50234 14792 50294
rect 14852 50294 15033 50297
rect 14852 50234 14926 50294
rect 14720 50231 14926 50234
rect 14986 50231 15033 50294
rect 8105 49063 8161 49221
rect 7491 47824 7547 47971
rect 8555 46817 8611 46979
rect 6967 46663 7166 46678
rect 6967 46608 6977 46663
rect 7032 46608 7098 46663
rect 7153 46608 7166 46663
rect 6967 46597 7166 46608
rect 7052 44147 7131 46597
rect 7841 46018 7912 46096
rect 7012 44118 7225 44147
rect 7012 44117 7145 44118
rect 7012 44062 7031 44117
rect 7083 44063 7145 44117
rect 7197 44063 7225 44118
rect 7083 44062 7225 44063
rect 7012 44035 7225 44062
rect 7819 43964 7933 46018
rect 13950 45231 14058 45269
rect 13950 45136 13967 45231
rect 14044 45136 14058 45231
rect 13950 45055 14058 45136
rect 13950 44960 13964 45055
rect 14041 44960 14058 45055
rect 13950 44896 14058 44960
rect 13950 44801 13966 44896
rect 14043 44801 14058 44896
rect 13950 44738 14058 44801
rect 13950 44643 13965 44738
rect 14042 44643 14058 44738
rect 13747 44188 13852 44243
rect 13747 44093 13767 44188
rect 13844 44093 13852 44188
rect 13747 44012 13852 44093
rect 7807 43946 7945 43964
rect 7807 43868 7834 43946
rect 7910 43868 7945 43946
rect 7807 43762 7945 43868
rect 7807 43684 7842 43762
rect 7918 43684 7945 43762
rect 7807 43640 7945 43684
rect 13747 43917 13764 44012
rect 13841 43917 13852 44012
rect 13747 43853 13852 43917
rect 13747 43758 13766 43853
rect 13843 43758 13852 43853
rect 13747 43695 13852 43758
rect 7819 43637 7933 43640
rect 13747 43600 13765 43695
rect 13842 43600 13852 43695
rect 13747 42638 13852 43600
rect 13950 42707 14058 44643
rect 14634 41904 15033 50231
rect 14634 41900 14923 41904
rect 14634 41899 14802 41900
rect 14634 41843 14659 41899
rect 14711 41844 14802 41899
rect 14854 41848 14923 41900
rect 14975 41848 15033 41904
rect 14854 41844 15033 41848
rect 14711 41843 15033 41844
rect 7287 41554 7474 41555
rect 7109 41542 7474 41554
rect 7109 41541 7232 41542
rect 7109 41487 7119 41541
rect 7173 41487 7232 41541
rect 7109 41486 7232 41487
rect 7288 41486 7474 41542
rect 7109 41472 7474 41486
rect 7109 41471 7296 41472
rect 7368 38782 7451 41472
rect 9493 41260 9549 41583
rect 9496 40381 9552 40630
rect 7318 38699 7451 38782
rect 6666 38523 6775 38541
rect 6665 38431 6674 38523
rect 6766 38431 6775 38523
rect 6666 38345 6775 38431
rect 6666 38251 6673 38345
rect 6767 38251 6775 38345
rect 6666 38235 6775 38251
rect 6455 35767 6563 35813
rect 6455 35709 6484 35767
rect 6549 35709 6563 35767
rect 6455 35640 6563 35709
rect 6455 35582 6480 35640
rect 6545 35582 6563 35640
rect 6455 32201 6563 35582
rect 7002 33192 7125 33206
rect 7002 33113 7022 33192
rect 7113 33113 7125 33192
rect 7002 33098 7125 33113
rect 7318 33098 7401 38699
rect 9545 38029 9602 38281
rect 13790 37020 13898 37050
rect 13790 36925 13806 37020
rect 13883 36925 13898 37020
rect 13790 36844 13898 36925
rect 13790 36749 13803 36844
rect 13880 36749 13898 36844
rect 13790 36685 13898 36749
rect 13790 36590 13805 36685
rect 13882 36590 13898 36685
rect 13790 36527 13898 36590
rect 13790 36432 13804 36527
rect 13881 36432 13898 36527
rect 13587 35760 13692 35799
rect 13587 35665 13601 35760
rect 13678 35665 13692 35760
rect 13587 35584 13692 35665
rect 13587 35489 13598 35584
rect 13675 35489 13692 35584
rect 13587 35425 13692 35489
rect 13587 35330 13600 35425
rect 13677 35330 13692 35425
rect 13587 35267 13692 35330
rect 13587 35172 13599 35267
rect 13676 35172 13692 35267
rect 13587 34151 13692 35172
rect 13790 34160 13898 36432
rect 7002 33040 7401 33098
rect 7002 32961 7018 33040
rect 7109 33015 7401 33040
rect 14634 33437 15033 41843
rect 14634 33433 14768 33437
rect 14634 33377 14655 33433
rect 14707 33381 14768 33433
rect 14820 33433 15033 33437
rect 14820 33381 14881 33433
rect 14707 33377 14881 33381
rect 14933 33377 15033 33433
rect 7109 32961 7125 33015
rect 7002 32949 7125 32961
rect 9333 32531 9389 32718
rect 6455 32129 6477 32201
rect 6543 32129 6563 32201
rect 6455 32044 6563 32129
rect 6455 31972 6478 32044
rect 6544 31972 6563 32044
rect 6455 31951 6563 31972
rect 9336 31876 9392 32111
rect 6690 31174 6813 31188
rect 6690 31131 6710 31174
rect 6205 31095 6710 31131
rect 6801 31095 6813 31174
rect 6205 31044 6813 31095
rect 6690 31022 6813 31044
rect 6690 30943 6706 31022
rect 6797 30943 6813 31022
rect 6690 30931 6813 30943
rect 4832 30739 5127 30740
rect 4832 30736 4971 30739
rect 4832 30672 4839 30736
rect 4895 30675 4971 30736
rect 5027 30676 5127 30739
rect 5183 30676 5231 30740
rect 5027 30675 5231 30676
rect 4895 30672 5231 30675
rect 4832 26025 5231 30672
rect 6045 30367 6502 30406
rect 6045 30256 6064 30367
rect 6175 30366 6502 30367
rect 6175 30257 6367 30366
rect 6476 30257 6502 30366
rect 6175 30256 6502 30257
rect 6045 30244 6502 30256
rect 6064 28369 6175 30244
rect 6409 29838 6753 29857
rect 6409 29837 6631 29838
rect 6409 29735 6427 29837
rect 6529 29735 6631 29837
rect 6409 29734 6631 29735
rect 6735 29734 6753 29838
rect 6409 29713 6753 29734
rect 6426 28486 6530 29713
rect 9385 29521 9442 29772
rect 6411 28470 6782 28486
rect 6411 28469 6658 28470
rect 6049 28351 6188 28369
rect 6411 28367 6432 28469
rect 6534 28367 6658 28469
rect 6411 28366 6658 28367
rect 6762 28366 6782 28470
rect 6411 28351 6782 28366
rect 13826 28459 13934 28498
rect 13826 28364 13845 28459
rect 13922 28364 13934 28459
rect 6049 28240 6064 28351
rect 6175 28240 6188 28351
rect 6049 28099 6188 28240
rect 6049 27990 6065 28099
rect 6174 27990 6188 28099
rect 6049 27972 6188 27990
rect 4832 26021 5134 26025
rect 4832 25923 4846 26021
rect 4915 26020 5134 26021
rect 4915 25923 4986 26020
rect 4832 25922 4986 25923
rect 5055 25927 5134 26020
rect 5203 25927 5231 26025
rect 5055 25922 5231 25927
rect 4832 22739 5231 25922
rect 5556 24108 5745 24109
rect 5556 24101 5749 24108
rect 5556 24044 5684 24101
rect 5737 24044 5749 24101
rect 5556 24035 5749 24044
rect 5556 23978 5571 24035
rect 5624 23978 5749 24035
rect 5556 23948 5749 23978
rect 5556 23891 5678 23948
rect 5731 23891 5749 23948
rect 5556 23870 5749 23891
rect 5556 23813 5574 23870
rect 5627 23813 5749 23870
rect 5556 23799 5749 23813
rect 4832 22738 5132 22739
rect 4832 22737 4991 22738
rect 4832 22675 4847 22737
rect 4911 22676 4991 22737
rect 5055 22677 5132 22738
rect 5196 22677 5231 22739
rect 5055 22676 5231 22677
rect 4911 22675 5231 22676
rect 4832 17012 5231 22675
rect 5559 19200 5749 23799
rect 6064 22347 6175 27972
rect 6064 22281 6085 22347
rect 6151 22281 6175 22347
rect 6064 22192 6175 22281
rect 6064 22124 6084 22192
rect 6152 22124 6175 22192
rect 6064 21040 6175 22124
rect 6426 21850 6530 28351
rect 13826 28283 13934 28364
rect 13826 28188 13842 28283
rect 13919 28188 13934 28283
rect 13826 28124 13934 28188
rect 13826 28029 13844 28124
rect 13921 28029 13934 28124
rect 13826 27966 13934 28029
rect 13826 27871 13843 27966
rect 13920 27871 13934 27966
rect 13623 27348 13728 27390
rect 13623 27253 13645 27348
rect 13722 27253 13728 27348
rect 13623 27172 13728 27253
rect 13623 27077 13642 27172
rect 13719 27077 13728 27172
rect 13623 27013 13728 27077
rect 13623 26918 13644 27013
rect 13721 26918 13728 27013
rect 13623 26855 13728 26918
rect 13623 26760 13643 26855
rect 13720 26760 13728 26855
rect 13623 26248 13728 26760
rect 13826 26086 13934 27871
rect 7039 25142 7162 25156
rect 7039 25063 7059 25142
rect 7150 25063 7162 25142
rect 7039 24990 7162 25063
rect 7039 24911 7055 24990
rect 7146 24911 7162 24990
rect 7039 24899 7162 24911
rect 9369 24388 9425 24598
rect 9372 23884 9428 24127
rect 14634 23673 15033 33377
rect 14634 23617 14654 23673
rect 14706 23672 15033 23673
rect 14706 23617 14782 23672
rect 14634 23616 14782 23617
rect 14834 23671 15033 23672
rect 14834 23616 14921 23671
rect 14634 23615 14921 23616
rect 14973 23615 15033 23671
rect 6708 23211 6831 23225
rect 6708 23132 6728 23211
rect 6819 23132 6831 23211
rect 6708 23059 6831 23132
rect 6708 22980 6724 23059
rect 6815 22980 6831 23059
rect 6708 22968 6831 22980
rect 6418 21824 6751 21850
rect 6417 21720 6426 21824
rect 6530 21823 6751 21824
rect 6530 21721 6637 21823
rect 6739 21721 6751 21823
rect 6530 21720 6751 21721
rect 6418 21704 6751 21720
rect 6052 21019 6189 21040
rect 6052 20907 6064 21019
rect 6175 20907 6189 21019
rect 6052 20793 6189 20907
rect 6052 20679 6064 20793
rect 6175 20679 6189 20793
rect 6052 20668 6189 20679
rect 5559 19116 5587 19200
rect 5719 19116 5749 19200
rect 5559 19046 5749 19116
rect 5559 18962 5591 19046
rect 5723 18962 5749 19046
rect 5559 18930 5749 18962
rect 4832 17011 5081 17012
rect 4832 16940 4841 17011
rect 4898 16940 4961 17011
rect 5018 16941 5081 17011
rect 5138 16941 5231 17012
rect 5018 16940 5231 16941
rect 4832 13220 5231 16940
rect 4832 13215 4981 13220
rect 4832 13151 4848 13215
rect 4910 13156 4981 13215
rect 5043 13156 5121 13220
rect 5183 13156 5231 13220
rect 4910 13151 5231 13156
rect 4832 11694 5231 13151
rect 4832 11693 4983 11694
rect 4832 11605 4843 11693
rect 4904 11606 4983 11693
rect 5044 11688 5231 11694
rect 5044 11606 5124 11688
rect 4904 11605 5124 11606
rect 4832 11600 5124 11605
rect 5185 11600 5231 11688
rect 4832 4338 5231 11600
rect 4832 4332 5142 4338
rect 4832 4328 4990 4332
rect 4832 4259 4842 4328
rect 4897 4263 4990 4328
rect 5045 4269 5142 4332
rect 5197 4269 5231 4338
rect 5045 4263 5231 4269
rect 4897 4259 5231 4263
rect 4832 844 5231 4259
rect 4832 841 4977 844
rect 4832 781 4848 841
rect 4910 784 4977 841
rect 5039 784 5110 844
rect 5172 784 5231 844
rect 4910 781 5231 784
rect 4832 -1078 5231 781
rect 4832 -1083 5158 -1078
rect 4832 -1084 4997 -1083
rect 4832 -1153 4847 -1084
rect 4902 -1152 4997 -1084
rect 5052 -1147 5158 -1083
rect 5213 -1147 5231 -1078
rect 5052 -1152 5231 -1147
rect 4902 -1153 5231 -1152
rect 4832 -4899 5231 -1153
rect 4832 -5001 4843 -4899
rect 4922 -4900 5139 -4899
rect 4922 -5001 4993 -4900
rect 4832 -5002 4993 -5001
rect 5072 -5001 5139 -4900
rect 5218 -5001 5231 -4899
rect 5072 -5002 5231 -5001
rect 4832 -7379 5231 -5002
rect 4832 -7383 5123 -7379
rect 4832 -7384 4996 -7383
rect 4832 -7438 4869 -7384
rect 4926 -7437 4996 -7384
rect 5053 -7433 5123 -7383
rect 5180 -7433 5231 -7379
rect 5053 -7437 5231 -7433
rect 4926 -7438 5231 -7437
rect 4832 -8742 5231 -7438
rect 4832 -8746 5100 -8742
rect 4832 -8747 4973 -8746
rect 4832 -8801 4846 -8747
rect 4903 -8800 4973 -8747
rect 5030 -8796 5100 -8746
rect 5157 -8796 5231 -8742
rect 5030 -8800 5231 -8796
rect 4903 -8801 5231 -8800
rect 4832 -9856 5231 -8801
rect 4832 -9858 5133 -9856
rect 4832 -9932 4844 -9858
rect 4899 -9860 5133 -9858
rect 4899 -9932 4983 -9860
rect 4832 -9934 4983 -9932
rect 5038 -9930 5133 -9860
rect 5188 -9930 5231 -9856
rect 5038 -9934 5231 -9930
rect 4832 -13533 5231 -9934
rect 5719 17462 5911 17485
rect 5719 17386 5770 17462
rect 5852 17386 5911 17462
rect 5719 17296 5911 17386
rect 5719 17220 5773 17296
rect 5855 17220 5911 17296
rect 5719 17128 5911 17220
rect 5719 17052 5779 17128
rect 5861 17052 5911 17128
rect 5719 14497 5911 17052
rect 5719 14431 5833 14497
rect 5892 14431 5911 14497
rect 5719 14318 5911 14431
rect 5719 14252 5826 14318
rect 5885 14252 5911 14318
rect 5719 2335 5911 14252
rect 6064 12876 6175 20668
rect 6426 20595 6530 21704
rect 9421 21537 9478 21774
rect 6416 20584 6543 20595
rect 6416 20480 6426 20584
rect 6530 20480 6543 20584
rect 6416 20346 6543 20480
rect 6416 20244 6427 20346
rect 6529 20244 6543 20346
rect 6416 20231 6543 20244
rect 6043 12849 6195 12876
rect 6043 12721 6064 12849
rect 6175 12721 6195 12849
rect 6043 12652 6195 12721
rect 6043 12543 6065 12652
rect 6174 12543 6195 12652
rect 6043 12527 6195 12543
rect 6426 12317 6530 20231
rect 13640 19413 13748 19451
rect 13640 19318 13661 19413
rect 13738 19318 13748 19413
rect 13640 19237 13748 19318
rect 13640 19142 13658 19237
rect 13735 19142 13748 19237
rect 13640 19078 13748 19142
rect 13640 18983 13660 19078
rect 13737 18983 13748 19078
rect 13640 18920 13748 18983
rect 13640 18825 13659 18920
rect 13736 18825 13748 18920
rect 13437 18337 13542 18368
rect 13437 18242 13455 18337
rect 13532 18242 13542 18337
rect 13437 18161 13542 18242
rect 13437 18066 13452 18161
rect 13529 18066 13542 18161
rect 13437 18002 13542 18066
rect 13437 17907 13454 18002
rect 13531 17907 13542 18002
rect 13437 17844 13542 17907
rect 13437 17749 13453 17844
rect 13530 17749 13542 17844
rect 13437 16625 13542 17749
rect 13640 16580 13748 18825
rect 14634 15993 15033 23615
rect 14634 15990 14896 15993
rect 14634 15934 14661 15990
rect 14713 15934 14775 15990
rect 14827 15937 14896 15990
rect 14948 15937 15033 15993
rect 14827 15934 15033 15937
rect 6877 15582 6964 15603
rect 6877 15526 6890 15582
rect 6946 15526 6964 15582
rect 6877 15471 6964 15526
rect 6877 15415 6886 15471
rect 6942 15415 6964 15471
rect 6877 15400 6964 15415
rect 9183 14835 9239 15099
rect 9186 14346 9242 14579
rect 6631 13730 6718 13751
rect 6631 13674 6644 13730
rect 6700 13674 6718 13730
rect 6631 13619 6718 13674
rect 6631 13563 6640 13619
rect 6696 13563 6718 13619
rect 6631 13548 6718 13563
rect 6227 12302 6544 12317
rect 6227 12301 6426 12302
rect 6227 12199 6254 12301
rect 6356 12199 6426 12301
rect 6227 12198 6426 12199
rect 6530 12198 6544 12302
rect 6227 12184 6544 12198
rect 9235 12024 9292 12255
rect 13854 7396 13962 7429
rect 13854 7301 13878 7396
rect 13955 7301 13962 7396
rect 13854 7220 13962 7301
rect 13854 7125 13875 7220
rect 13952 7125 13962 7220
rect 13854 7061 13962 7125
rect 13854 6966 13877 7061
rect 13954 6966 13962 7061
rect 13854 6903 13962 6966
rect 13854 6808 13876 6903
rect 13953 6808 13962 6903
rect 13655 6185 13756 6188
rect 13651 6162 13756 6185
rect 13651 6067 13673 6162
rect 13750 6067 13756 6162
rect 13651 5986 13756 6067
rect 13651 5891 13670 5986
rect 13747 5891 13756 5986
rect 13651 5827 13756 5891
rect 13651 5732 13672 5827
rect 13749 5732 13756 5827
rect 13651 5669 13756 5732
rect 13651 5574 13671 5669
rect 13748 5574 13756 5669
rect 13651 4072 13756 5574
rect 13854 4238 13962 6808
rect 14634 3468 15033 15934
rect 14634 3463 14923 3468
rect 14634 3456 14798 3463
rect 14634 3400 14651 3456
rect 14703 3407 14798 3456
rect 14850 3412 14923 3463
rect 14975 3412 15033 3468
rect 14850 3407 15033 3412
rect 14703 3400 15033 3407
rect 7103 3168 7190 3189
rect 7103 3112 7116 3168
rect 7172 3112 7190 3168
rect 7103 3057 7190 3112
rect 7103 3001 7112 3057
rect 7168 3001 7190 3057
rect 7103 2986 7190 3001
rect 9397 2467 9453 2675
rect 5719 2266 5832 2335
rect 5896 2266 5911 2335
rect 5719 2169 5911 2266
rect 5719 2100 5831 2169
rect 5895 2100 5911 2169
rect 5719 -12009 5911 2100
rect 9400 1989 9456 2229
rect 6759 1266 6846 1287
rect 6759 1210 6772 1266
rect 6828 1210 6846 1266
rect 6759 1155 6846 1210
rect 6759 1099 6768 1155
rect 6824 1099 6846 1155
rect 6759 1084 6846 1099
rect 9449 -370 9506 -120
rect 13833 -2429 13941 -2404
rect 13833 -2455 13942 -2429
rect 13833 -2550 13859 -2455
rect 13936 -2550 13942 -2455
rect 13833 -2631 13942 -2550
rect 13833 -2726 13856 -2631
rect 13933 -2726 13942 -2631
rect 13833 -2790 13942 -2726
rect 13833 -2885 13858 -2790
rect 13935 -2885 13942 -2790
rect 13833 -2948 13942 -2885
rect 13833 -3043 13857 -2948
rect 13934 -3043 13942 -2948
rect 13833 -3066 13942 -3043
rect 13630 -3500 13735 -3492
rect 13630 -3526 13739 -3500
rect 13630 -3621 13656 -3526
rect 13733 -3621 13739 -3526
rect 13630 -3702 13739 -3621
rect 13630 -3797 13653 -3702
rect 13730 -3797 13739 -3702
rect 13630 -3861 13739 -3797
rect 13630 -3956 13655 -3861
rect 13732 -3956 13739 -3861
rect 13630 -4019 13739 -3956
rect 13630 -4114 13654 -4019
rect 13731 -4114 13739 -4019
rect 13630 -4137 13739 -4114
rect 13630 -5431 13735 -4137
rect 13833 -5480 13941 -3066
rect 7086 -6370 7173 -6349
rect 7086 -6426 7099 -6370
rect 7155 -6426 7173 -6370
rect 7086 -6481 7173 -6426
rect 7086 -6537 7095 -6481
rect 7151 -6537 7173 -6481
rect 7086 -6552 7173 -6537
rect 9376 -7140 9432 -6922
rect 14634 -7236 15033 3400
rect 14634 -7237 14900 -7236
rect 14634 -7238 14766 -7237
rect 14634 -7294 14647 -7238
rect 14699 -7293 14766 -7238
rect 14818 -7292 14900 -7237
rect 14952 -7292 15033 -7236
rect 14818 -7293 15033 -7292
rect 14699 -7294 15033 -7293
rect 9379 -7613 9435 -7367
rect 6460 -8328 6745 -8295
rect 6460 -8410 6473 -8328
rect 6555 -8410 6638 -8328
rect 6720 -8410 6745 -8328
rect 6460 -8448 6745 -8410
rect 9428 -9966 9485 -9708
rect 6176 -10177 6613 -10168
rect 6176 -10305 6184 -10177
rect 6312 -10305 6474 -10177
rect 6602 -10305 6613 -10177
rect 6176 -10319 6613 -10305
rect 6474 -10866 6586 -10319
rect 6459 -10880 6869 -10866
rect 6459 -10992 6474 -10880
rect 6586 -10881 6869 -10880
rect 6586 -10991 6747 -10881
rect 6857 -10991 6869 -10881
rect 6586 -10992 6869 -10991
rect 6459 -11004 6869 -10992
rect 13841 -11381 13949 -11321
rect 13841 -11476 13862 -11381
rect 13939 -11476 13949 -11381
rect 13841 -11557 13949 -11476
rect 13841 -11652 13859 -11557
rect 13936 -11652 13949 -11557
rect 13841 -11716 13949 -11652
rect 13841 -11811 13861 -11716
rect 13938 -11811 13949 -11716
rect 13841 -11874 13949 -11811
rect 13841 -11969 13860 -11874
rect 13937 -11969 13949 -11874
rect 6237 -12009 6395 -11995
rect 5719 -12060 6395 -12009
rect 5719 -12133 6271 -12060
rect 6370 -12133 6395 -12060
rect 5719 -12201 6395 -12133
rect 4832 -13536 5122 -13533
rect 4832 -13610 4844 -13536
rect 4907 -13539 5122 -13536
rect 4907 -13610 5001 -13539
rect 4832 -13613 5001 -13610
rect 5064 -13607 5122 -13539
rect 5185 -13607 5231 -13533
rect 5064 -13613 5231 -13607
rect 4832 -17196 5231 -13613
rect 6237 -12216 6395 -12201
rect 6237 -12289 6271 -12216
rect 6370 -12289 6395 -12216
rect 6237 -12372 6395 -12289
rect 6237 -12445 6266 -12372
rect 6365 -12445 6395 -12372
rect 13638 -12396 13743 -12381
rect 6237 -15840 6395 -12445
rect 13634 -12422 13743 -12396
rect 13634 -12517 13652 -12422
rect 13729 -12517 13743 -12422
rect 13634 -12598 13743 -12517
rect 13634 -12693 13649 -12598
rect 13726 -12693 13743 -12598
rect 13634 -12757 13743 -12693
rect 13634 -12852 13651 -12757
rect 13728 -12852 13743 -12757
rect 13634 -12915 13743 -12852
rect 13634 -13010 13650 -12915
rect 13727 -13010 13743 -12915
rect 13634 -13033 13743 -13010
rect 13638 -13885 13743 -13033
rect 13841 -13802 13949 -11969
rect 14634 -14527 15033 -7294
rect 14634 -14583 14645 -14527
rect 14697 -14583 14761 -14527
rect 14813 -14531 15033 -14527
rect 14813 -14583 14876 -14531
rect 14634 -14587 14876 -14583
rect 14928 -14587 15033 -14531
rect 7092 -14862 7179 -14841
rect 7092 -14918 7105 -14862
rect 7161 -14918 7179 -14862
rect 7092 -14973 7179 -14918
rect 7092 -15029 7101 -14973
rect 7157 -14975 7179 -14973
rect 7157 -15029 7309 -14975
rect 7092 -15044 7309 -15029
rect 7160 -15052 7309 -15044
rect 6237 -15919 6286 -15840
rect 6347 -15919 6395 -15840
rect 6237 -16023 6395 -15919
rect 6237 -16102 6285 -16023
rect 6346 -16102 6395 -16023
rect 6237 -16288 6395 -16102
rect 4832 -17199 4966 -17196
rect 4832 -17269 4843 -17199
rect 4901 -17266 4966 -17199
rect 5024 -17197 5231 -17196
rect 5024 -17266 5105 -17197
rect 4901 -17267 5105 -17266
rect 5163 -17267 5231 -17197
rect 4901 -17269 5231 -17267
rect 4832 -18959 5231 -17269
rect 4832 -18961 5148 -18959
rect 4832 -19035 4848 -18961
rect 4911 -19035 4986 -18961
rect 5049 -19033 5148 -18961
rect 5211 -19033 5231 -18959
rect 5049 -19035 5231 -19033
rect 4832 -21627 5231 -19035
rect 5825 -20218 5925 -20140
rect 5825 -20282 5842 -20218
rect 5908 -20282 5925 -20218
rect 5825 -20374 5925 -20282
rect 5408 -20448 5503 -20418
rect 5408 -20504 5431 -20448
rect 5486 -20504 5503 -20448
rect 5408 -20578 5503 -20504
rect 5408 -20634 5426 -20578
rect 5481 -20634 5503 -20578
rect 5408 -20655 5503 -20634
rect 5825 -20438 5842 -20374
rect 5908 -20438 5925 -20374
rect 6271 -20166 6362 -16288
rect 6633 -16765 6771 -16748
rect 6633 -16836 6667 -16765
rect 6738 -16836 6771 -16765
rect 6633 -16941 6771 -16836
rect 6633 -17012 6663 -16941
rect 6734 -17012 6771 -16941
rect 6633 -17022 6771 -17012
rect 6271 -20226 6286 -20166
rect 6343 -20226 6362 -20166
rect 6271 -20312 6362 -20226
rect 6271 -20372 6284 -20312
rect 6341 -20372 6362 -20312
rect 6271 -20388 6362 -20372
rect 6704 -18133 6798 -18118
rect 6704 -18194 6721 -18133
rect 6780 -18194 6798 -18133
rect 6704 -18261 6798 -18194
rect 6704 -18322 6724 -18261
rect 6783 -18322 6798 -18261
rect 4832 -21631 4996 -21627
rect 4832 -21726 4842 -21631
rect 4915 -21722 4996 -21631
rect 5069 -21629 5231 -21627
rect 5069 -21722 5143 -21629
rect 4915 -21724 5143 -21722
rect 5216 -21724 5231 -21629
rect 4915 -21726 5231 -21724
rect 4832 -25402 5231 -21726
rect 4832 -25406 5117 -25402
rect 4832 -25462 4859 -25406
rect 4911 -25407 5117 -25406
rect 4911 -25462 5002 -25407
rect 4832 -25463 5002 -25462
rect 5054 -25458 5117 -25407
rect 5169 -25458 5231 -25402
rect 5054 -25463 5231 -25458
rect 4832 -26564 5231 -25463
rect 4832 -26565 4985 -26564
rect 4832 -26658 4840 -26565
rect 4913 -26657 4985 -26565
rect 5058 -26567 5231 -26564
rect 5058 -26657 5131 -26567
rect 4913 -26658 5131 -26657
rect 4832 -26660 5131 -26658
rect 5204 -26660 5231 -26567
rect 4832 -29790 5231 -26660
rect 4832 -29793 4991 -29790
rect 4832 -29869 4844 -29793
rect 4918 -29866 4991 -29793
rect 5065 -29791 5231 -29790
rect 5065 -29866 5139 -29791
rect 4918 -29867 5139 -29866
rect 5213 -29867 5231 -29791
rect 4918 -29869 5231 -29867
rect 4832 -33417 5231 -29869
rect 4832 -33419 4998 -33417
rect 4832 -33486 4841 -33419
rect 4907 -33484 4998 -33419
rect 5064 -33418 5231 -33417
rect 5064 -33484 5135 -33418
rect 4907 -33485 5135 -33484
rect 5201 -33485 5231 -33418
rect 4907 -33486 5231 -33485
rect 4832 -35027 5231 -33486
rect 4832 -35030 4985 -35027
rect 4832 -35093 4853 -35030
rect 4913 -35090 4985 -35030
rect 5045 -35030 5231 -35027
rect 5045 -35090 5119 -35030
rect 4913 -35093 5119 -35090
rect 5179 -35093 5231 -35030
rect 4832 -36500 5231 -35093
rect 5409 -35236 5504 -20655
rect 5580 -20796 5675 -20764
rect 5580 -20851 5597 -20796
rect 5655 -20851 5675 -20796
rect 5580 -20939 5675 -20851
rect 5580 -20994 5597 -20939
rect 5655 -20994 5675 -20939
rect 5580 -34522 5675 -20994
rect 5825 -23779 5925 -20438
rect 6704 -20827 6798 -18322
rect 6986 -20452 7080 -18604
rect 6986 -20505 7005 -20452
rect 7063 -20505 7080 -20452
rect 6986 -20575 7080 -20505
rect 6986 -20628 7004 -20575
rect 7062 -20628 7080 -20575
rect 6986 -20646 7080 -20628
rect 6988 -20657 7077 -20646
rect 6527 -20855 6800 -20827
rect 6527 -20911 6573 -20855
rect 6637 -20862 6800 -20855
rect 6637 -20911 6714 -20862
rect 6527 -20918 6714 -20911
rect 6778 -20918 6800 -20862
rect 6527 -20965 6800 -20918
rect 7232 -23218 7309 -15052
rect 9384 -15588 9440 -15426
rect 9387 -16080 9443 -15816
rect 9436 -18395 9493 -18174
rect 13965 -19445 14073 -19428
rect 13962 -19471 14073 -19445
rect 13962 -19566 13980 -19471
rect 14057 -19566 14073 -19471
rect 13962 -19647 14073 -19566
rect 13962 -19742 13977 -19647
rect 14054 -19742 14073 -19647
rect 13962 -19806 14073 -19742
rect 13962 -19901 13979 -19806
rect 14056 -19901 14073 -19806
rect 13962 -19964 14073 -19901
rect 13962 -20059 13978 -19964
rect 14055 -20059 14073 -19964
rect 13962 -20082 14073 -20059
rect 13762 -20487 13867 -20471
rect 13760 -20513 13867 -20487
rect 13760 -20608 13778 -20513
rect 13855 -20608 13867 -20513
rect 13760 -20689 13867 -20608
rect 13760 -20784 13775 -20689
rect 13852 -20784 13867 -20689
rect 13760 -20848 13867 -20784
rect 13760 -20943 13777 -20848
rect 13854 -20943 13867 -20848
rect 13760 -21006 13867 -20943
rect 13760 -21101 13776 -21006
rect 13853 -21101 13867 -21006
rect 13760 -21124 13867 -21101
rect 13762 -21919 13867 -21124
rect 13965 -21963 14073 -20082
rect 14634 -22571 15033 -14587
rect 14634 -22578 14765 -22571
rect 14634 -22634 14652 -22578
rect 14704 -22627 14765 -22578
rect 14817 -22627 14888 -22571
rect 14940 -22627 15033 -22571
rect 14704 -22634 15033 -22627
rect 14634 -23006 15033 -22634
rect 14634 -23013 14771 -23006
rect 14634 -23069 14658 -23013
rect 14710 -23062 14771 -23013
rect 14823 -23062 14894 -23006
rect 14946 -23062 15033 -23006
rect 14710 -23069 15033 -23062
rect 7232 -23295 7352 -23218
rect 5825 -23869 5976 -23779
rect 5823 -23940 5976 -23869
rect 5823 -24003 5833 -23940
rect 5909 -24003 5976 -23940
rect 5823 -24097 5976 -24003
rect 5823 -24160 5834 -24097
rect 5910 -24160 5976 -24097
rect 5823 -24171 5976 -24160
rect 5580 -34579 5606 -34522
rect 5663 -34579 5675 -34522
rect 5580 -34668 5675 -34579
rect 5580 -34723 5607 -34668
rect 5662 -34723 5675 -34668
rect 5580 -34737 5675 -34723
rect 5409 -35299 5426 -35236
rect 5486 -35299 5504 -35236
rect 5409 -35369 5504 -35299
rect 5409 -35432 5426 -35369
rect 5486 -35432 5504 -35369
rect 5409 -35453 5504 -35432
rect 4832 -36517 5243 -36500
rect 4832 -36520 5160 -36517
rect 4832 -36525 5011 -36520
rect 4832 -36620 4852 -36525
rect 4929 -36615 5011 -36525
rect 5088 -36612 5160 -36520
rect 5237 -36612 5243 -36517
rect 5088 -36615 5243 -36612
rect 4929 -36620 5243 -36615
rect 4832 -36693 5243 -36620
rect 4832 -36696 5157 -36693
rect 4832 -36701 5008 -36696
rect 4832 -36796 4849 -36701
rect 4926 -36791 5008 -36701
rect 5085 -36788 5157 -36696
rect 5234 -36788 5243 -36693
rect 5085 -36791 5243 -36788
rect 4926 -36796 5243 -36791
rect 4832 -36852 5243 -36796
rect 4832 -36855 5159 -36852
rect 4832 -36860 5010 -36855
rect 4832 -36955 4851 -36860
rect 4928 -36950 5010 -36860
rect 5087 -36947 5159 -36855
rect 5236 -36947 5243 -36852
rect 5087 -36950 5243 -36947
rect 4928 -36955 5243 -36950
rect 4832 -37010 5243 -36955
rect 4832 -37013 5158 -37010
rect 4832 -37018 5009 -37013
rect 4832 -37113 4850 -37018
rect 4927 -37108 5009 -37018
rect 5086 -37105 5158 -37013
rect 5235 -37105 5243 -37010
rect 5825 -37027 5976 -24171
rect 7275 -24908 7352 -23295
rect 9508 -23729 9564 -23542
rect 9511 -24268 9567 -24048
rect 6656 -24974 6999 -24908
rect 6656 -24990 6880 -24974
rect 6656 -25067 6666 -24990
rect 6734 -25051 6880 -24990
rect 6948 -25051 6999 -24974
rect 6734 -25067 6999 -25051
rect 6656 -25121 6999 -25067
rect 7275 -24937 7532 -24908
rect 7275 -24987 7446 -24937
rect 7275 -25063 7285 -24987
rect 7353 -25013 7446 -24987
rect 7514 -25013 7532 -24937
rect 7353 -25063 7532 -25013
rect 7275 -25077 7532 -25063
rect 6406 -25762 6508 -25749
rect 6399 -25772 6515 -25762
rect 6399 -25848 6419 -25772
rect 6495 -25848 6515 -25772
rect 6399 -25854 6424 -25848
rect 6490 -25854 6515 -25848
rect 6399 -25962 6515 -25854
rect 6399 -26030 6423 -25962
rect 6491 -26030 6515 -25962
rect 6399 -27469 6515 -26030
rect 6696 -26315 6813 -26290
rect 6696 -26390 6710 -26315
rect 6785 -26390 6813 -26315
rect 6696 -26394 6813 -26390
rect 6687 -26481 6813 -26394
rect 6687 -26558 6709 -26481
rect 6786 -26558 6813 -26481
rect 6687 -26576 6813 -26558
rect 6687 -27136 6811 -26576
rect 9560 -26611 9617 -26365
rect 6687 -27221 6707 -27136
rect 6785 -27221 6811 -27136
rect 6687 -27296 6811 -27221
rect 6687 -27381 6709 -27296
rect 6787 -27381 6811 -27296
rect 6392 -27521 6516 -27469
rect 6392 -27601 6418 -27521
rect 6498 -27601 6516 -27521
rect 6392 -27678 6516 -27601
rect 6392 -27758 6415 -27678
rect 6495 -27758 6516 -27678
rect 6392 -27789 6516 -27758
rect 6399 -30446 6515 -27789
rect 6399 -30527 6412 -30446
rect 6492 -30527 6515 -30446
rect 6399 -30587 6515 -30527
rect 6399 -30668 6415 -30587
rect 6495 -30668 6515 -30587
rect 6399 -35533 6515 -30668
rect 6687 -29611 6811 -27381
rect 6687 -29667 6708 -29611
rect 6764 -29667 6811 -29611
rect 6687 -29724 6811 -29667
rect 6687 -29780 6708 -29724
rect 6764 -29780 6811 -29724
rect 6122 -35545 6536 -35533
rect 6122 -35558 6399 -35545
rect 6122 -35648 6128 -35558
rect 6218 -35648 6399 -35558
rect 6122 -35661 6399 -35648
rect 6495 -35661 6536 -35545
rect 6122 -35681 6536 -35661
rect 6687 -35815 6811 -29780
rect 14634 -30719 15033 -23069
rect 14634 -30722 14792 -30719
rect 14634 -30785 14660 -30722
rect 14720 -30782 14792 -30722
rect 14852 -30722 15033 -30719
rect 14852 -30782 14926 -30722
rect 14720 -30785 14926 -30782
rect 14986 -30785 15033 -30722
rect 14634 -31150 15033 -30785
rect 14634 -31153 14792 -31150
rect 14634 -31216 14660 -31153
rect 14720 -31213 14792 -31153
rect 14852 -31153 15033 -31150
rect 14852 -31213 14926 -31153
rect 14720 -31216 14926 -31213
rect 14986 -31216 15033 -31153
rect 8166 -32267 8222 -32120
rect 7552 -33487 7608 -33353
rect 8616 -34549 8672 -34355
rect 6366 -35839 6828 -35815
rect 6366 -35844 6687 -35839
rect 6366 -35931 6418 -35844
rect 6526 -35931 6687 -35844
rect 6366 -35936 6687 -35931
rect 6811 -35936 6828 -35839
rect 6366 -35982 6828 -35936
rect 14634 -36328 15033 -31216
rect 14634 -36332 14793 -36328
rect 14634 -36414 14656 -36332
rect 14723 -36410 14793 -36332
rect 14860 -36332 15033 -36328
rect 14860 -36410 14935 -36332
rect 14723 -36414 14935 -36410
rect 15002 -36414 15033 -36332
rect 5086 -37108 5243 -37105
rect 4927 -37113 5243 -37108
rect 4832 -37125 5243 -37113
rect 5764 -37071 6006 -37027
rect 5764 -37076 5919 -37071
rect 4068 -37553 4480 -37536
rect 4068 -37556 4397 -37553
rect 4068 -37561 4248 -37556
rect 4068 -37656 4089 -37561
rect 4166 -37651 4248 -37561
rect 4325 -37648 4397 -37556
rect 4474 -37648 4480 -37553
rect 4325 -37651 4480 -37648
rect 4166 -37656 4480 -37651
rect 4068 -37729 4480 -37656
rect 4068 -37732 4394 -37729
rect 4068 -37737 4245 -37732
rect 4068 -37832 4086 -37737
rect 4163 -37827 4245 -37737
rect 4322 -37824 4394 -37732
rect 4471 -37824 4480 -37729
rect 4322 -37827 4480 -37824
rect 4163 -37832 4480 -37827
rect 4068 -37888 4480 -37832
rect 4068 -37891 4396 -37888
rect 4068 -37896 4247 -37891
rect 4068 -37991 4088 -37896
rect 4165 -37986 4247 -37896
rect 4324 -37983 4396 -37891
rect 4473 -37983 4480 -37888
rect 4324 -37986 4480 -37983
rect 4165 -37991 4480 -37986
rect 4068 -38046 4480 -37991
rect 4068 -38049 4395 -38046
rect 4068 -38054 4246 -38049
rect 4068 -38149 4087 -38054
rect 4164 -38144 4246 -38054
rect 4323 -38141 4395 -38049
rect 4472 -38141 4480 -38046
rect 4323 -38144 4480 -38141
rect 4164 -38149 4480 -38144
rect 4068 -38161 4480 -38149
rect 4832 -37714 5231 -37125
rect 5764 -37158 5792 -37076
rect 5848 -37153 5919 -37076
rect 5975 -37153 6006 -37071
rect 5848 -37158 6006 -37153
rect 5764 -37188 6006 -37158
rect 14634 -37544 15033 -36414
rect 15320 51242 15719 55224
rect 25331 54811 25730 55873
rect 26017 55849 26416 55873
rect 26017 55832 26427 55849
rect 26017 55829 26344 55832
rect 26017 55824 26195 55829
rect 26017 55729 26036 55824
rect 26113 55734 26195 55824
rect 26272 55737 26344 55829
rect 26421 55737 26427 55832
rect 26272 55734 26427 55737
rect 26113 55729 26427 55734
rect 26017 55656 26427 55729
rect 26017 55653 26341 55656
rect 26017 55648 26192 55653
rect 26017 55553 26033 55648
rect 26110 55558 26192 55648
rect 26269 55561 26341 55653
rect 26418 55561 26427 55656
rect 26269 55558 26427 55561
rect 26110 55553 26427 55558
rect 26017 55497 26427 55553
rect 26017 55494 26343 55497
rect 26017 55489 26194 55494
rect 26017 55394 26035 55489
rect 26112 55399 26194 55489
rect 26271 55402 26343 55494
rect 26420 55402 26427 55497
rect 26271 55399 26427 55402
rect 26112 55394 26427 55399
rect 26017 55339 26427 55394
rect 26017 55336 26342 55339
rect 26017 55331 26193 55336
rect 26017 55236 26034 55331
rect 26111 55241 26193 55331
rect 26270 55244 26342 55336
rect 26419 55244 26427 55339
rect 26270 55241 26427 55244
rect 26111 55236 26427 55241
rect 26017 55224 26427 55236
rect 25328 54794 25738 54811
rect 25328 54791 25655 54794
rect 25328 54786 25506 54791
rect 25328 54691 25347 54786
rect 25424 54696 25506 54786
rect 25583 54699 25655 54791
rect 25732 54699 25738 54794
rect 25583 54696 25738 54699
rect 25424 54691 25738 54696
rect 25328 54618 25738 54691
rect 25328 54615 25652 54618
rect 25328 54610 25503 54615
rect 25328 54515 25344 54610
rect 25421 54520 25503 54610
rect 25580 54523 25652 54615
rect 25729 54523 25738 54618
rect 25580 54520 25738 54523
rect 25421 54515 25738 54520
rect 25328 54459 25738 54515
rect 25328 54456 25654 54459
rect 25328 54451 25505 54456
rect 25328 54356 25346 54451
rect 25423 54361 25505 54451
rect 25582 54364 25654 54456
rect 25731 54364 25738 54459
rect 25582 54361 25738 54364
rect 25423 54356 25738 54361
rect 25328 54301 25738 54356
rect 25328 54298 25653 54301
rect 25328 54293 25504 54298
rect 25328 54198 25345 54293
rect 25422 54203 25504 54293
rect 25581 54206 25653 54298
rect 25730 54206 25738 54301
rect 25581 54203 25738 54206
rect 25422 54198 25738 54203
rect 25328 54186 25738 54198
rect 24595 53602 24703 53634
rect 24595 53507 24616 53602
rect 24693 53507 24703 53602
rect 24595 53426 24703 53507
rect 24595 53331 24613 53426
rect 24690 53331 24703 53426
rect 24595 53267 24703 53331
rect 24595 53172 24615 53267
rect 24692 53172 24703 53267
rect 24595 53109 24703 53172
rect 24595 53014 24614 53109
rect 24691 53014 24703 53109
rect 24392 52557 24497 52596
rect 16644 52468 17105 52473
rect 16644 52461 17106 52468
rect 16644 52362 16664 52461
rect 16763 52460 17106 52461
rect 16763 52363 16857 52460
rect 16954 52363 17106 52460
rect 16763 52362 17106 52363
rect 16644 52348 17106 52362
rect 15320 51153 15334 51242
rect 15395 51241 15719 51242
rect 15395 51153 15482 51241
rect 15320 51152 15482 51153
rect 15543 51152 15644 51241
rect 15705 51152 15719 51241
rect 15320 48912 15719 51152
rect 15320 48909 15482 48912
rect 15320 48846 15350 48909
rect 15410 48849 15482 48909
rect 15542 48909 15719 48912
rect 15542 48849 15616 48909
rect 15410 48846 15616 48849
rect 15676 48846 15719 48909
rect 15320 47557 15719 48846
rect 15320 47554 15474 47557
rect 15320 47491 15342 47554
rect 15402 47494 15474 47554
rect 15534 47554 15719 47557
rect 15534 47494 15608 47554
rect 15402 47491 15608 47494
rect 15668 47491 15719 47554
rect 15320 42945 15719 47491
rect 16526 49916 16635 49968
rect 16526 49846 16552 49916
rect 16623 49846 16635 49916
rect 16526 49745 16635 49846
rect 16526 49675 16549 49745
rect 16620 49675 16635 49745
rect 15320 42943 15464 42945
rect 15320 42872 15330 42943
rect 15389 42874 15464 42943
rect 15523 42874 15601 42945
rect 15660 42874 15719 42945
rect 15389 42872 15719 42874
rect 15320 39172 15719 42872
rect 16254 45105 16393 45174
rect 16254 45017 16282 45105
rect 16382 45017 16393 45105
rect 16254 44907 16393 45017
rect 16254 44819 16272 44907
rect 16372 44819 16393 44907
rect 16254 40529 16393 44819
rect 16254 40463 16299 40529
rect 16363 40463 16393 40529
rect 16254 40391 16393 40463
rect 16254 40325 16301 40391
rect 16365 40325 16393 40391
rect 16254 40239 16393 40325
rect 16254 40173 16289 40239
rect 16353 40173 16393 40239
rect 16254 39880 16393 40173
rect 16526 41532 16635 49675
rect 16526 41459 16546 41532
rect 16617 41459 16635 41532
rect 16526 41362 16635 41459
rect 16526 41289 16541 41362
rect 16612 41289 16635 41362
rect 15320 39116 15353 39172
rect 15405 39166 15719 39172
rect 15405 39162 15594 39166
rect 15405 39116 15470 39162
rect 15320 39106 15470 39116
rect 15522 39110 15594 39162
rect 15646 39110 15719 39166
rect 15522 39106 15719 39110
rect 15320 34440 15719 39106
rect 15320 34439 15622 34440
rect 15320 34362 15327 34439
rect 15402 34362 15478 34439
rect 15553 34363 15622 34439
rect 15697 34363 15719 34440
rect 15553 34362 15719 34363
rect 15320 30696 15719 34362
rect 16259 35984 16388 39880
rect 16526 37256 16635 41289
rect 16752 48012 16861 48061
rect 16752 47952 16787 48012
rect 16840 47952 16861 48012
rect 16752 47869 16861 47952
rect 16752 47809 16781 47869
rect 16834 47809 16861 47869
rect 16752 39657 16861 47809
rect 17012 46852 17106 52348
rect 24392 52462 24412 52557
rect 24489 52462 24497 52557
rect 24392 52381 24497 52462
rect 24392 52286 24409 52381
rect 24486 52286 24497 52381
rect 24392 52222 24497 52286
rect 17262 52195 17412 52214
rect 17262 52090 17284 52195
rect 17389 52090 17412 52195
rect 17262 51993 17412 52090
rect 17262 51886 17283 51993
rect 17390 51886 17412 51993
rect 17262 51875 17412 51886
rect 24392 52127 24411 52222
rect 24488 52127 24497 52222
rect 24392 52064 24497 52127
rect 24392 51969 24410 52064
rect 24487 51969 24497 52064
rect 17283 47179 17390 51875
rect 24392 51581 24497 51969
rect 24392 51525 24420 51581
rect 24475 51525 24497 51581
rect 24392 50924 24497 51525
rect 24595 51442 24703 53014
rect 24595 51386 24626 51442
rect 24681 51386 24703 51442
rect 24595 50977 24703 51386
rect 20141 49940 20736 49942
rect 20138 49886 20736 49940
rect 20138 49776 20194 49886
rect 20141 48919 20197 48938
rect 20141 48865 20142 48919
rect 20196 48865 20197 48919
rect 20141 48758 20197 48865
rect 17283 47072 17838 47179
rect 16994 46829 17122 46852
rect 16994 46737 17013 46829
rect 17105 46737 17122 46829
rect 16994 46668 17122 46737
rect 16994 46574 17012 46668
rect 17106 46574 17122 46668
rect 16994 46560 17122 46574
rect 16745 39643 16868 39657
rect 16745 39564 16765 39643
rect 16856 39564 16868 39643
rect 16745 39491 16868 39564
rect 16745 39412 16761 39491
rect 16852 39412 16868 39491
rect 16745 39400 16868 39412
rect 16752 37600 16861 39400
rect 17012 38435 17106 46560
rect 17283 38792 17390 47072
rect 24601 45228 24709 45273
rect 24601 45133 24617 45228
rect 24694 45133 24709 45228
rect 24601 45052 24709 45133
rect 24601 44957 24614 45052
rect 24691 44957 24709 45052
rect 24601 44893 24709 44957
rect 24601 44798 24616 44893
rect 24693 44798 24709 44893
rect 24601 44735 24709 44798
rect 24601 44640 24615 44735
rect 24692 44640 24709 44735
rect 24398 44188 24503 44237
rect 24398 44093 24415 44188
rect 24492 44093 24503 44188
rect 24398 44012 24503 44093
rect 24398 43917 24412 44012
rect 24489 43917 24503 44012
rect 24398 43853 24503 43917
rect 24398 43758 24414 43853
rect 24491 43758 24503 43853
rect 24398 43695 24503 43758
rect 24398 43600 24413 43695
rect 24490 43600 24503 43695
rect 24398 42617 24503 43600
rect 24601 42578 24709 44640
rect 25331 42019 25730 54186
rect 25331 42016 25485 42019
rect 25331 41953 25353 42016
rect 25413 41956 25485 42016
rect 25545 42016 25730 42019
rect 25545 41956 25619 42016
rect 25413 41953 25619 41956
rect 25679 41953 25730 42016
rect 17838 41565 17961 41579
rect 17838 41486 17858 41565
rect 17949 41486 17961 41565
rect 17838 41413 17961 41486
rect 17838 41334 17854 41413
rect 17945 41334 17961 41413
rect 17838 41322 17961 41334
rect 20144 40930 20200 41268
rect 20147 40297 20203 40527
rect 17283 38685 17848 38792
rect 16996 38419 17117 38435
rect 16996 38327 17013 38419
rect 17105 38327 17117 38419
rect 16996 38260 17117 38327
rect 16996 38166 17012 38260
rect 17106 38166 17117 38260
rect 16996 38144 17117 38166
rect 20196 37974 20253 38198
rect 16752 37491 17241 37600
rect 16526 37147 16956 37256
rect 16259 35921 16285 35984
rect 16365 35921 16388 35984
rect 16259 35818 16388 35921
rect 16259 35755 16281 35818
rect 16361 35755 16388 35818
rect 16259 31739 16388 35755
rect 16561 34941 16677 35056
rect 16561 34867 16585 34941
rect 16649 34867 16677 34941
rect 16561 34797 16677 34867
rect 16561 34723 16589 34797
rect 16653 34786 16677 34797
rect 16653 34723 16682 34786
rect 16561 34703 16682 34723
rect 16563 32212 16682 34703
rect 16847 33071 16956 37147
rect 16847 33000 16873 33071
rect 16940 33000 16956 33071
rect 16847 32888 16956 33000
rect 16847 32817 16864 32888
rect 16931 32817 16956 32888
rect 16564 32171 16681 32212
rect 16564 32101 16584 32171
rect 16661 32101 16681 32171
rect 16564 32007 16681 32101
rect 16564 31937 16583 32007
rect 16660 31937 16681 32007
rect 16564 31913 16681 31937
rect 16259 31605 16601 31739
rect 15320 30690 15459 30696
rect 15320 30634 15339 30690
rect 15391 30640 15459 30690
rect 15511 30640 15595 30696
rect 15647 30640 15719 30696
rect 15391 30634 15719 30640
rect 15320 26441 15719 30634
rect 15320 26365 15331 26441
rect 15402 26365 15484 26441
rect 15555 26438 15719 26441
rect 15555 26365 15637 26438
rect 15320 26362 15637 26365
rect 15708 26362 15719 26438
rect 15320 21232 15719 26362
rect 16450 22620 16601 31605
rect 16847 25378 16956 32817
rect 17132 31133 17241 37491
rect 24685 37016 24793 37075
rect 24685 36921 24704 37016
rect 24781 36921 24793 37016
rect 24685 36840 24793 36921
rect 24685 36745 24701 36840
rect 24778 36745 24793 36840
rect 24685 36681 24793 36745
rect 24685 36586 24703 36681
rect 24780 36586 24793 36681
rect 24685 36523 24793 36586
rect 24685 36428 24702 36523
rect 24779 36428 24793 36523
rect 24482 35766 24587 35821
rect 24482 35671 24503 35766
rect 24580 35671 24587 35766
rect 24482 35590 24587 35671
rect 24482 35495 24500 35590
rect 24577 35495 24587 35590
rect 24482 35431 24587 35495
rect 24482 35336 24502 35431
rect 24579 35336 24587 35431
rect 24482 35273 24587 35336
rect 24482 35178 24501 35273
rect 24578 35178 24587 35273
rect 24482 34057 24587 35178
rect 24685 34137 24793 36428
rect 25331 33512 25730 41953
rect 25331 33509 25488 33512
rect 25331 33446 25356 33509
rect 25416 33449 25488 33509
rect 25548 33509 25730 33512
rect 25548 33449 25622 33509
rect 25416 33446 25622 33449
rect 25682 33446 25730 33509
rect 17889 33195 18012 33209
rect 17889 33116 17909 33195
rect 18000 33116 18012 33195
rect 17889 33043 18012 33116
rect 17889 32964 17905 33043
rect 17996 32964 18012 33043
rect 17889 32952 18012 32964
rect 20228 32255 20284 32577
rect 20231 31879 20287 32073
rect 17132 31119 17283 31133
rect 17132 31040 17180 31119
rect 17271 31040 17283 31119
rect 17132 30967 17283 31040
rect 17132 30888 17176 30967
rect 17267 30888 17283 30967
rect 17132 30876 17283 30888
rect 16780 25337 16973 25378
rect 16780 25231 16819 25337
rect 16940 25231 16973 25337
rect 16780 25117 16973 25231
rect 16780 25011 16814 25117
rect 16935 25011 16973 25117
rect 16780 24982 16973 25011
rect 17132 24723 17241 30876
rect 17440 30304 17538 30329
rect 17440 30238 17459 30304
rect 17525 30238 17538 30304
rect 17440 30138 17538 30238
rect 17440 30105 17458 30138
rect 17439 30070 17458 30105
rect 17526 30070 17538 30138
rect 17439 30055 17538 30070
rect 17439 28836 17522 30055
rect 17636 29778 17749 29810
rect 17636 29701 17655 29778
rect 17732 29701 17749 29778
rect 17636 29632 17749 29701
rect 17636 29593 17646 29632
rect 17630 29555 17646 29593
rect 17724 29555 17749 29632
rect 17630 29532 17749 29555
rect 17427 28824 17529 28836
rect 17427 28741 17439 28824
rect 17522 28741 17531 28824
rect 17427 28677 17529 28741
rect 17427 28590 17439 28677
rect 17522 28590 17529 28677
rect 17427 28578 17529 28590
rect 16949 24614 17241 24723
rect 16949 23299 17058 24614
rect 17439 24339 17522 28578
rect 17630 27152 17725 29532
rect 20280 29505 20337 29734
rect 18511 28460 18650 28480
rect 18511 28356 18531 28460
rect 18635 28356 18650 28460
rect 18511 28277 18650 28356
rect 18511 28175 18532 28277
rect 18634 28175 18650 28277
rect 18511 28158 18650 28175
rect 17881 28036 18025 28105
rect 17881 27925 17899 28036
rect 18010 27925 18025 28036
rect 17881 27787 18025 27925
rect 17881 27678 17900 27787
rect 18009 27678 18025 27787
rect 17881 27658 18025 27678
rect 17619 27140 17734 27152
rect 17619 27137 17631 27140
rect 17724 27137 17734 27140
rect 17619 27042 17630 27137
rect 17725 27042 17734 27137
rect 17619 26970 17734 27042
rect 17619 26875 17630 26970
rect 17725 26875 17734 26970
rect 17619 26867 17734 26875
rect 17195 24256 17522 24339
rect 16872 23252 17065 23299
rect 16872 23144 16922 23252
rect 17027 23144 17065 23252
rect 16872 23039 17065 23144
rect 16872 22931 16914 23039
rect 17019 22931 17065 23039
rect 16872 22899 17065 22931
rect 16853 22620 17070 22626
rect 16450 22415 17070 22620
rect 15320 21228 15443 21232
rect 15320 21172 15336 21228
rect 15388 21176 15443 21228
rect 15495 21228 15719 21232
rect 15495 21176 15568 21228
rect 15388 21172 15568 21176
rect 15620 21172 15719 21228
rect 15320 16920 15719 21172
rect 15320 16842 15334 16920
rect 15388 16917 15719 16920
rect 15388 16842 15475 16917
rect 15320 16839 15475 16842
rect 15529 16916 15719 16917
rect 15529 16839 15626 16916
rect 15320 16838 15626 16839
rect 15680 16838 15719 16916
rect 15320 13245 15719 16838
rect 15320 13238 15595 13245
rect 15320 13236 15459 13238
rect 15320 13180 15341 13236
rect 15393 13182 15459 13236
rect 15511 13189 15595 13238
rect 15647 13189 15719 13245
rect 15511 13182 15719 13189
rect 15393 13180 15719 13182
rect 15320 11531 15719 13180
rect 15320 11530 15493 11531
rect 15320 11452 15340 11530
rect 15394 11453 15493 11530
rect 15547 11522 15719 11531
rect 15547 11453 15626 11522
rect 15394 11452 15626 11453
rect 15320 11444 15626 11452
rect 15680 11444 15719 11522
rect 15320 4522 15719 11444
rect 15320 4519 15584 4522
rect 15320 4463 15344 4519
rect 15396 4463 15472 4519
rect 15524 4466 15584 4519
rect 15636 4466 15719 4522
rect 15524 4463 15719 4466
rect 15320 833 15719 4463
rect 16853 14566 17070 22415
rect 16853 14511 17004 14566
rect 17059 14511 17070 14566
rect 16853 14424 17070 14511
rect 16853 14369 17000 14424
rect 17055 14369 17070 14424
rect 16853 2229 17070 14369
rect 17195 11842 17278 24256
rect 17630 24042 17725 26867
rect 17896 26001 18007 27658
rect 18531 26610 18635 28158
rect 18530 26390 18635 26610
rect 18531 26381 18635 26390
rect 17881 25964 18020 26001
rect 17881 25855 17897 25964
rect 18006 25855 18020 25964
rect 17881 25750 18020 25855
rect 17881 25639 17896 25750
rect 18007 25639 18020 25750
rect 17881 25616 18020 25639
rect 17355 23947 17725 24042
rect 18814 23982 18870 24127
rect 17355 12350 17450 23947
rect 25331 23614 25730 33446
rect 25331 23611 25480 23614
rect 25331 23548 25348 23611
rect 25408 23551 25480 23611
rect 25540 23611 25730 23614
rect 25540 23551 25614 23611
rect 25408 23548 25614 23551
rect 25674 23548 25730 23611
rect 18200 22759 18256 22889
rect 19264 21719 19320 21916
rect 17638 21601 17856 21611
rect 17638 21600 17790 21601
rect 17638 21545 17650 21600
rect 17705 21545 17790 21600
rect 17638 21544 17790 21545
rect 17847 21544 17856 21601
rect 17638 21535 17856 21544
rect 17644 19579 17748 21535
rect 18550 20962 18621 21035
rect 18533 19877 18637 20962
rect 18270 19864 18676 19877
rect 18270 19863 18527 19864
rect 18270 19729 18278 19863
rect 18412 19729 18527 19863
rect 18270 19728 18527 19729
rect 18663 19728 18676 19864
rect 18270 19716 18676 19728
rect 17628 19539 17769 19579
rect 17628 19459 17656 19539
rect 17738 19459 17769 19539
rect 17628 19367 17769 19459
rect 17628 19287 17656 19367
rect 17738 19287 17769 19367
rect 17628 19256 17769 19287
rect 24697 19416 24805 19451
rect 24697 19321 24721 19416
rect 24798 19321 24805 19416
rect 24697 19240 24805 19321
rect 24697 19145 24718 19240
rect 24795 19145 24805 19240
rect 24697 19081 24805 19145
rect 24697 18986 24720 19081
rect 24797 18986 24805 19081
rect 24697 18923 24805 18986
rect 24697 18828 24719 18923
rect 24796 18828 24805 18923
rect 24494 18330 24599 18363
rect 24494 18235 24516 18330
rect 24593 18235 24599 18330
rect 24494 18154 24599 18235
rect 24494 18059 24513 18154
rect 24590 18059 24599 18154
rect 24494 17995 24599 18059
rect 24494 17900 24515 17995
rect 24592 17900 24599 17995
rect 24494 17837 24599 17900
rect 24494 17742 24514 17837
rect 24591 17742 24599 17837
rect 24494 16631 24599 17742
rect 24697 16624 24805 18828
rect 25331 15988 25730 23548
rect 25331 15985 25480 15988
rect 25331 15922 25348 15985
rect 25408 15925 25480 15985
rect 25540 15985 25730 15988
rect 25540 15925 25614 15985
rect 25408 15922 25614 15925
rect 25674 15922 25730 15985
rect 17940 15592 18027 15613
rect 17940 15536 17953 15592
rect 18009 15536 18027 15592
rect 17940 15481 18027 15536
rect 17940 15425 17949 15481
rect 18005 15425 18027 15481
rect 17940 15410 18027 15425
rect 20240 14887 20296 15086
rect 20243 14378 20299 14628
rect 17627 13700 17714 13721
rect 17627 13644 17640 13700
rect 17696 13644 17714 13700
rect 17627 13589 17714 13644
rect 17627 13533 17636 13589
rect 17692 13533 17714 13589
rect 17627 13518 17714 13533
rect 17355 12333 17605 12350
rect 17355 12332 17522 12333
rect 17355 12257 17365 12332
rect 17441 12257 17522 12332
rect 17355 12256 17522 12257
rect 17599 12256 17608 12333
rect 17355 12246 17605 12256
rect 17355 12244 17450 12246
rect 20292 12042 20349 12283
rect 17195 11759 17945 11842
rect 24697 7389 24805 7417
rect 24697 7294 24719 7389
rect 24796 7294 24805 7389
rect 24697 7213 24805 7294
rect 24697 7118 24716 7213
rect 24793 7118 24805 7213
rect 24697 7054 24805 7118
rect 24697 6959 24718 7054
rect 24795 6959 24805 7054
rect 24697 6896 24805 6959
rect 24697 6801 24717 6896
rect 24794 6801 24805 6896
rect 24494 6184 24599 6208
rect 24494 6158 24600 6184
rect 24494 6063 24517 6158
rect 24594 6063 24600 6158
rect 24494 5982 24600 6063
rect 24494 5887 24514 5982
rect 24591 5887 24600 5982
rect 24494 5823 24600 5887
rect 24494 5728 24516 5823
rect 24593 5728 24600 5823
rect 24494 5665 24600 5728
rect 24494 5570 24515 5665
rect 24592 5570 24600 5665
rect 24494 5547 24600 5570
rect 24494 4108 24599 5547
rect 24697 4143 24805 6801
rect 25331 3251 25730 15922
rect 25331 3248 25486 3251
rect 25331 3185 25354 3248
rect 25414 3188 25486 3248
rect 25546 3248 25730 3251
rect 25546 3188 25620 3248
rect 25414 3185 25620 3188
rect 25680 3185 25730 3248
rect 17949 3088 18036 3109
rect 17949 3032 17962 3088
rect 18018 3032 18036 3088
rect 17949 2977 18036 3032
rect 17949 2921 17958 2977
rect 18014 2921 18036 2977
rect 17949 2906 18036 2921
rect 20240 2344 20296 2555
rect 15320 830 15590 833
rect 15320 774 15350 830
rect 15402 774 15478 830
rect 15530 777 15590 830
rect 15642 777 15719 833
rect 15530 774 15719 777
rect 15320 722 15719 774
rect 15320 719 15591 722
rect 15320 663 15351 719
rect 15403 663 15479 719
rect 15531 666 15591 719
rect 15643 666 15719 722
rect 15531 663 15719 666
rect 15320 -656 15719 663
rect 15320 -658 15606 -656
rect 15320 -733 15332 -658
rect 15395 -662 15606 -658
rect 15395 -733 15474 -662
rect 15320 -737 15474 -733
rect 15537 -731 15606 -662
rect 15669 -731 15719 -656
rect 15537 -737 15719 -731
rect 15320 -5009 15719 -737
rect 15320 -5013 15462 -5009
rect 15320 -5084 15330 -5013
rect 15396 -5080 15462 -5013
rect 15528 -5012 15719 -5009
rect 15528 -5080 15623 -5012
rect 15396 -5083 15623 -5080
rect 15689 -5083 15719 -5012
rect 15396 -5084 15719 -5083
rect 15320 -5196 15719 -5084
rect 15320 -5198 15632 -5196
rect 15320 -5269 15328 -5198
rect 15394 -5200 15632 -5198
rect 15394 -5269 15478 -5200
rect 15320 -5271 15478 -5269
rect 15544 -5267 15632 -5200
rect 15698 -5267 15719 -5196
rect 15544 -5271 15719 -5267
rect 15320 -8676 15719 -5271
rect 15320 -8736 15330 -8676
rect 15384 -8736 15461 -8676
rect 15515 -8678 15719 -8676
rect 15515 -8736 15602 -8678
rect 15320 -8738 15602 -8736
rect 15656 -8738 15719 -8678
rect 15320 -9669 15719 -8738
rect 15320 -9672 15585 -9669
rect 15320 -9681 15463 -9672
rect 15320 -9737 15334 -9681
rect 15386 -9728 15463 -9681
rect 15515 -9725 15585 -9672
rect 15637 -9725 15719 -9669
rect 15515 -9728 15719 -9725
rect 15386 -9737 15719 -9728
rect 15320 -13652 15719 -9737
rect 15320 -13654 15467 -13652
rect 15320 -13727 15328 -13654
rect 15382 -13725 15467 -13654
rect 15521 -13654 15719 -13652
rect 15521 -13725 15611 -13654
rect 15382 -13727 15611 -13725
rect 15665 -13727 15719 -13654
rect 15320 -17266 15719 -13727
rect 16031 2211 17070 2229
rect 16031 2151 17002 2211
rect 17058 2151 17070 2211
rect 16031 2036 17070 2151
rect 16031 1976 16999 2036
rect 17055 1976 17070 2036
rect 16031 1959 17070 1976
rect 16031 -11530 16301 1959
rect 16908 1949 17070 1959
rect 20243 1851 20299 2101
rect 17564 1148 17651 1169
rect 17564 1092 17577 1148
rect 17633 1092 17651 1148
rect 17564 1037 17651 1092
rect 17564 981 17573 1037
rect 17629 981 17651 1037
rect 17564 966 17651 981
rect 16031 -11606 16091 -11530
rect 16172 -11606 16301 -11530
rect 16031 -11738 16301 -11606
rect 16675 -195 16810 -175
rect 16675 -270 16703 -195
rect 16778 -270 16810 -195
rect 16675 -409 16810 -270
rect 16675 -486 16702 -409
rect 16779 -486 16810 -409
rect 16675 -1246 16810 -486
rect 20292 -506 20349 -245
rect 16675 -1323 16700 -1246
rect 16778 -1323 16810 -1246
rect 16675 -1410 16810 -1323
rect 16675 -1487 16705 -1410
rect 16783 -1487 16810 -1410
rect 16675 -4365 16810 -1487
rect 16675 -4437 16703 -4365
rect 16775 -4437 16810 -4365
rect 16675 -4528 16810 -4437
rect 16675 -4602 16702 -4528
rect 16776 -4602 16810 -4528
rect 16675 -11607 16810 -4602
rect 16996 -688 17131 -654
rect 16996 -765 17013 -688
rect 17091 -765 17131 -688
rect 16996 -852 17131 -765
rect 16996 -929 17018 -852
rect 17096 -929 17131 -852
rect 16996 -5027 17131 -929
rect 16996 -5029 17282 -5027
rect 16996 -5076 17659 -5029
rect 16996 -5077 17541 -5076
rect 16996 -5135 17262 -5077
rect 17318 -5083 17541 -5077
rect 17318 -5135 17380 -5083
rect 16996 -5141 17380 -5135
rect 17436 -5134 17541 -5083
rect 17597 -5134 17659 -5076
rect 17436 -5141 17659 -5134
rect 16996 -5192 17659 -5141
rect 16996 -5204 17200 -5192
rect 16996 -11284 17131 -5204
rect 18846 -6908 18902 -6750
rect 25331 -7280 25730 3185
rect 25331 -7283 25486 -7280
rect 25331 -7346 25354 -7283
rect 25414 -7343 25486 -7283
rect 25546 -7283 25730 -7280
rect 25546 -7343 25620 -7283
rect 25414 -7346 25620 -7343
rect 25680 -7346 25730 -7283
rect 18232 -8013 18288 -7906
rect 19296 -9185 19352 -9000
rect 17304 -9304 17503 -9291
rect 17304 -9361 17316 -9304
rect 17373 -9359 17437 -9304
rect 17492 -9359 17503 -9304
rect 17373 -9361 17503 -9359
rect 17304 -9368 17503 -9361
rect 17311 -10855 17446 -9368
rect 17282 -10865 17758 -10855
rect 17282 -11004 17294 -10865
rect 17433 -10867 17758 -10865
rect 17433 -11004 17605 -10867
rect 17742 -11004 17758 -10867
rect 17282 -11018 17758 -11004
rect 16985 -11301 17147 -11284
rect 16985 -11437 16996 -11301
rect 17131 -11437 17147 -11301
rect 16031 -11814 16087 -11738
rect 16168 -11814 16301 -11738
rect 16031 -15889 16301 -11814
rect 16663 -11623 16822 -11607
rect 16663 -11759 16675 -11623
rect 16810 -11759 16822 -11623
rect 16663 -11977 16822 -11759
rect 16985 -11634 17147 -11437
rect 16985 -11770 16996 -11634
rect 17131 -11770 17147 -11634
rect 16985 -11785 17147 -11770
rect 24685 -11381 24793 -11333
rect 24685 -11476 24703 -11381
rect 24780 -11476 24793 -11381
rect 24685 -11557 24793 -11476
rect 24685 -11652 24700 -11557
rect 24777 -11652 24793 -11557
rect 24685 -11716 24793 -11652
rect 16663 -12113 16675 -11977
rect 16810 -12113 16822 -11977
rect 16663 -12125 16822 -12113
rect 16031 -15892 16448 -15889
rect 16031 -15950 16457 -15892
rect 16031 -16020 16378 -15950
rect 16441 -16020 16457 -15950
rect 16031 -16138 16457 -16020
rect 16031 -16208 16380 -16138
rect 16443 -16208 16457 -16138
rect 16031 -16346 16457 -16208
rect 15320 -17273 15588 -17266
rect 15320 -17280 15472 -17273
rect 15320 -17336 15331 -17280
rect 15383 -17329 15472 -17280
rect 15524 -17322 15588 -17273
rect 15640 -17322 15719 -17266
rect 15524 -17329 15719 -17322
rect 15383 -17336 15719 -17329
rect 15320 -18973 15719 -17336
rect 15320 -18974 15628 -18973
rect 15320 -19047 15336 -18974
rect 15390 -18975 15628 -18974
rect 15390 -19047 15472 -18975
rect 15320 -19048 15472 -19047
rect 15526 -19046 15628 -18975
rect 15682 -19046 15719 -18973
rect 15526 -19048 15719 -19046
rect 15320 -21704 15719 -19048
rect 15320 -21705 15612 -21704
rect 15320 -21777 15332 -21705
rect 15388 -21708 15612 -21705
rect 15388 -21777 15472 -21708
rect 15320 -21780 15472 -21777
rect 15528 -21776 15612 -21708
rect 15668 -21776 15719 -21704
rect 15528 -21780 15719 -21776
rect 15320 -25325 15719 -21780
rect 15320 -25336 15457 -25325
rect 15320 -25392 15341 -25336
rect 15393 -25381 15457 -25336
rect 15509 -25330 15719 -25325
rect 15509 -25381 15582 -25330
rect 15393 -25386 15582 -25381
rect 15634 -25386 15719 -25330
rect 15393 -25392 15719 -25386
rect 15320 -26949 15719 -25392
rect 15320 -26951 15480 -26949
rect 15320 -27044 15336 -26951
rect 15401 -27042 15480 -26951
rect 15545 -26951 15719 -26949
rect 15545 -27042 15622 -26951
rect 15401 -27044 15622 -27042
rect 15687 -27044 15719 -26951
rect 15320 -30094 15719 -27044
rect 15320 -30098 15636 -30094
rect 15320 -30101 15479 -30098
rect 15320 -30191 15334 -30101
rect 15405 -30188 15479 -30101
rect 15550 -30184 15636 -30098
rect 15707 -30184 15719 -30094
rect 15550 -30188 15719 -30184
rect 15405 -30191 15719 -30188
rect 15320 -33462 15719 -30191
rect 16367 -31652 16457 -16346
rect 16675 -18022 16810 -12125
rect 16996 -17509 17131 -11785
rect 24685 -11811 24702 -11716
rect 24779 -11811 24793 -11716
rect 24685 -11874 24793 -11811
rect 24685 -11969 24701 -11874
rect 24778 -11969 24793 -11874
rect 24482 -12418 24587 -12381
rect 24482 -12513 24502 -12418
rect 24579 -12513 24587 -12418
rect 24482 -12594 24587 -12513
rect 24482 -12689 24499 -12594
rect 24576 -12689 24587 -12594
rect 24482 -12753 24587 -12689
rect 24482 -12848 24501 -12753
rect 24578 -12848 24587 -12753
rect 24482 -12911 24587 -12848
rect 24482 -13006 24500 -12911
rect 24577 -13006 24587 -12911
rect 24482 -13885 24587 -13006
rect 24685 -13923 24793 -11969
rect 25331 -14490 25730 -7346
rect 25331 -14493 25492 -14490
rect 25331 -14556 25360 -14493
rect 25420 -14553 25492 -14493
rect 25552 -14493 25730 -14490
rect 25552 -14553 25626 -14493
rect 25420 -14556 25626 -14553
rect 25686 -14556 25730 -14493
rect 17933 -14910 18020 -14889
rect 17933 -14966 17946 -14910
rect 18002 -14966 18020 -14910
rect 17933 -15021 18020 -14966
rect 17933 -15077 17942 -15021
rect 17998 -15077 18020 -15021
rect 17933 -15092 18020 -15077
rect 20228 -15689 20284 -15418
rect 20231 -16145 20287 -15884
rect 17414 -16820 17552 -16803
rect 17414 -16891 17448 -16820
rect 17519 -16891 17552 -16820
rect 17414 -16996 17552 -16891
rect 17414 -17067 17444 -16996
rect 17515 -17067 17552 -16996
rect 17414 -17077 17552 -17067
rect 16996 -17575 17042 -17509
rect 17108 -17575 17131 -17509
rect 16996 -17698 17131 -17575
rect 16996 -17764 17042 -17698
rect 17108 -17764 17131 -17698
rect 16996 -17792 17131 -17764
rect 16675 -18099 16702 -18022
rect 16779 -18099 16810 -18022
rect 16675 -18191 16810 -18099
rect 16675 -18266 16703 -18191
rect 16778 -18266 16810 -18191
rect 16675 -18328 16810 -18266
rect 20280 -18484 20337 -18244
rect 24673 -19466 24781 -19440
rect 24673 -19561 24692 -19466
rect 24769 -19561 24781 -19466
rect 24673 -19642 24781 -19561
rect 24673 -19737 24689 -19642
rect 24766 -19737 24781 -19642
rect 24673 -19801 24781 -19737
rect 24673 -19896 24691 -19801
rect 24768 -19896 24781 -19801
rect 24673 -19959 24781 -19896
rect 24673 -20054 24690 -19959
rect 24767 -20054 24781 -19959
rect 17073 -20217 17173 -20171
rect 17073 -20325 17089 -20217
rect 17158 -20325 17173 -20217
rect 17073 -20463 17173 -20325
rect 17073 -20571 17089 -20463
rect 17158 -20571 17173 -20463
rect 24470 -20487 24575 -20471
rect 17073 -20592 17173 -20571
rect 24467 -20513 24575 -20487
rect 17073 -23643 17171 -20592
rect 24467 -20608 24485 -20513
rect 24562 -20608 24575 -20513
rect 24467 -20689 24575 -20608
rect 24467 -20784 24482 -20689
rect 24559 -20784 24575 -20689
rect 24467 -20848 24575 -20784
rect 24467 -20943 24484 -20848
rect 24561 -20943 24575 -20848
rect 24467 -21006 24575 -20943
rect 24467 -21101 24483 -21006
rect 24560 -21101 24575 -21006
rect 24467 -21124 24575 -21101
rect 24470 -21950 24575 -21124
rect 24673 -21926 24781 -20054
rect 25331 -22616 25730 -14556
rect 25331 -22619 25485 -22616
rect 25331 -22682 25353 -22619
rect 25413 -22679 25485 -22619
rect 25545 -22619 25730 -22616
rect 25545 -22679 25619 -22619
rect 25413 -22682 25619 -22679
rect 25679 -22682 25730 -22619
rect 25331 -23042 25730 -22682
rect 25331 -23045 25486 -23042
rect 25331 -23108 25354 -23045
rect 25414 -23105 25486 -23045
rect 25546 -23045 25730 -23042
rect 25546 -23105 25620 -23045
rect 25414 -23108 25620 -23105
rect 25680 -23108 25730 -23045
rect 17002 -23651 17171 -23643
rect 16972 -23765 17171 -23651
rect 20216 -23706 20272 -23507
rect 16972 -23782 17172 -23765
rect 16972 -23870 17087 -23782
rect 17153 -23870 17172 -23782
rect 16972 -23957 17172 -23870
rect 16972 -24045 17086 -23957
rect 17152 -24045 17172 -23957
rect 16972 -24061 17172 -24045
rect 16972 -24063 17171 -24061
rect 17002 -24068 17171 -24063
rect 15320 -33465 15480 -33462
rect 15320 -33528 15348 -33465
rect 15408 -33525 15480 -33465
rect 15540 -33465 15719 -33462
rect 15540 -33525 15614 -33465
rect 15408 -33528 15614 -33525
rect 15674 -33528 15719 -33465
rect 15320 -35017 15719 -33528
rect 15320 -35021 15601 -35017
rect 15320 -35111 15333 -35021
rect 15404 -35111 15470 -35021
rect 15541 -35107 15601 -35021
rect 15672 -35107 15719 -35017
rect 15541 -35111 15719 -35107
rect 15320 -36500 15719 -35111
rect 16340 -31906 16484 -31652
rect 16340 -31985 16383 -31906
rect 16454 -31985 16484 -31906
rect 16340 -32112 16484 -31985
rect 16340 -32191 16384 -32112
rect 16455 -32191 16484 -32112
rect 15316 -36517 15726 -36500
rect 15316 -36520 15643 -36517
rect 15316 -36525 15494 -36520
rect 15316 -36620 15335 -36525
rect 15412 -36615 15494 -36525
rect 15571 -36612 15643 -36520
rect 15720 -36612 15726 -36517
rect 15571 -36615 15726 -36612
rect 15412 -36620 15726 -36615
rect 15316 -36693 15726 -36620
rect 15316 -36696 15640 -36693
rect 15316 -36701 15491 -36696
rect 15316 -36796 15332 -36701
rect 15409 -36791 15491 -36701
rect 15568 -36788 15640 -36696
rect 15717 -36788 15726 -36693
rect 15568 -36791 15726 -36788
rect 15409 -36796 15726 -36791
rect 15316 -36852 15726 -36796
rect 15316 -36855 15642 -36852
rect 15316 -36860 15493 -36855
rect 15316 -36955 15334 -36860
rect 15411 -36950 15493 -36860
rect 15570 -36947 15642 -36855
rect 15719 -36947 15726 -36852
rect 15570 -36950 15726 -36947
rect 15411 -36955 15726 -36950
rect 15316 -37010 15726 -36955
rect 15316 -37013 15641 -37010
rect 15316 -37018 15492 -37013
rect 15316 -37113 15333 -37018
rect 15410 -37108 15492 -37018
rect 15569 -37105 15641 -37013
rect 15718 -37105 15726 -37010
rect 15569 -37108 15726 -37105
rect 15410 -37113 15726 -37108
rect 15316 -37125 15726 -37113
rect 4832 -37716 5125 -37714
rect 4832 -37804 4856 -37716
rect 4919 -37804 4998 -37716
rect 5061 -37802 5125 -37716
rect 5188 -37802 5231 -37714
rect 5061 -37804 5231 -37802
rect 4068 -38182 4467 -38161
rect 4832 -38182 5231 -37804
rect 14630 -37561 15040 -37544
rect 14630 -37564 14957 -37561
rect 14630 -37569 14808 -37564
rect 14630 -37664 14649 -37569
rect 14726 -37659 14808 -37569
rect 14885 -37656 14957 -37564
rect 15034 -37656 15040 -37561
rect 14885 -37659 15040 -37656
rect 14726 -37664 15040 -37659
rect 14630 -37737 15040 -37664
rect 14630 -37740 14954 -37737
rect 14630 -37745 14805 -37740
rect 14630 -37840 14646 -37745
rect 14723 -37835 14805 -37745
rect 14882 -37832 14954 -37740
rect 15031 -37832 15040 -37737
rect 14882 -37835 15040 -37832
rect 14723 -37840 15040 -37835
rect 14630 -37896 15040 -37840
rect 14630 -37899 14956 -37896
rect 14630 -37904 14807 -37899
rect 14630 -37999 14648 -37904
rect 14725 -37994 14807 -37904
rect 14884 -37991 14956 -37899
rect 15033 -37991 15040 -37896
rect 14884 -37994 15040 -37991
rect 14725 -37999 15040 -37994
rect 14630 -38054 15040 -37999
rect 14630 -38057 14955 -38054
rect 14630 -38062 14806 -38057
rect 14630 -38157 14647 -38062
rect 14724 -38152 14806 -38062
rect 14883 -38149 14955 -38057
rect 15032 -38149 15040 -38054
rect 14883 -38152 15040 -38149
rect 14724 -38157 15040 -38152
rect 14630 -38169 15040 -38157
rect 15320 -37840 15719 -37125
rect 16340 -37152 16484 -32191
rect 17002 -34971 17147 -24068
rect 20219 -24185 20275 -24019
rect 17320 -24952 17731 -24878
rect 17320 -24962 17593 -24952
rect 17320 -25055 17338 -24962
rect 17421 -25045 17593 -24962
rect 17676 -25045 17731 -24952
rect 17421 -25055 17731 -25045
rect 17320 -25100 17731 -25055
rect 17455 -33037 17563 -25100
rect 20268 -26533 20325 -26286
rect 24722 -27513 24830 -27472
rect 24722 -27608 24741 -27513
rect 24818 -27608 24830 -27513
rect 24722 -27689 24830 -27608
rect 24722 -27784 24738 -27689
rect 24815 -27784 24830 -27689
rect 24722 -27848 24830 -27784
rect 24722 -27943 24740 -27848
rect 24817 -27943 24830 -27848
rect 24722 -28006 24830 -27943
rect 24722 -28101 24739 -28006
rect 24816 -28101 24830 -28006
rect 24519 -28555 24624 -28515
rect 24519 -28650 24539 -28555
rect 24616 -28650 24624 -28555
rect 24519 -28731 24624 -28650
rect 24519 -28826 24536 -28731
rect 24613 -28826 24624 -28731
rect 24519 -28890 24624 -28826
rect 24519 -28985 24538 -28890
rect 24615 -28985 24624 -28890
rect 24519 -29048 24624 -28985
rect 24519 -29143 24537 -29048
rect 24614 -29143 24624 -29048
rect 24519 -30085 24624 -29143
rect 24722 -30130 24830 -28101
rect 20265 -31788 20321 -31609
rect 20268 -32341 20324 -32156
rect 17455 -33091 17772 -33037
rect 17455 -33093 17683 -33091
rect 17455 -33157 17525 -33093
rect 17583 -33155 17683 -33093
rect 17741 -33155 17772 -33091
rect 17583 -33157 17772 -33155
rect 17455 -33160 17772 -33157
rect 17512 -33184 17772 -33160
rect 17352 -34405 17660 -34373
rect 17352 -34469 17381 -34405
rect 17446 -34469 17499 -34405
rect 17564 -34469 17660 -34405
rect 17352 -34500 17660 -34469
rect 16198 -37199 16484 -37152
rect 16806 -35116 17147 -34971
rect 16806 -37162 16951 -35116
rect 17534 -35833 17659 -34500
rect 20317 -34659 20374 -34433
rect 17889 -34889 17952 -34750
rect 17870 -35340 17971 -34889
rect 17852 -35419 17989 -35340
rect 17852 -35499 17882 -35419
rect 17963 -35499 17989 -35419
rect 17852 -35559 17989 -35499
rect 17852 -35639 17881 -35559
rect 17962 -35639 17989 -35559
rect 17852 -35667 17989 -35639
rect 17870 -35669 17971 -35667
rect 17218 -35857 17659 -35833
rect 17218 -35861 17557 -35857
rect 17218 -35938 17255 -35861
rect 17337 -35862 17557 -35861
rect 17337 -35938 17403 -35862
rect 17218 -35939 17403 -35938
rect 17485 -35934 17557 -35862
rect 17639 -35934 17659 -35857
rect 17485 -35939 17659 -35934
rect 17218 -35958 17659 -35939
rect 16198 -37205 16357 -37199
rect 16198 -37266 16226 -37205
rect 16291 -37260 16357 -37205
rect 16422 -37260 16484 -37199
rect 16291 -37266 16484 -37260
rect 16198 -37296 16484 -37266
rect 16799 -37200 17156 -37162
rect 16799 -37202 17067 -37200
rect 16799 -37209 16950 -37202
rect 16799 -37283 16823 -37209
rect 16883 -37276 16950 -37209
rect 17010 -37274 17067 -37202
rect 17127 -37274 17156 -37200
rect 17010 -37276 17156 -37274
rect 16883 -37283 17156 -37276
rect 16799 -37301 17156 -37283
rect 15320 -37841 15617 -37840
rect 15320 -37923 15331 -37841
rect 15398 -37923 15466 -37841
rect 15533 -37922 15617 -37841
rect 15684 -37922 15719 -37840
rect 15533 -37923 15719 -37922
rect 14634 -38182 15033 -38169
rect 15320 -38182 15719 -37923
rect 25331 -37533 25730 -23108
rect 26017 51265 26416 55224
rect 26017 51262 26325 51265
rect 26017 51260 26161 51262
rect 26017 51178 26024 51260
rect 26083 51180 26161 51260
rect 26220 51183 26325 51262
rect 26384 51183 26416 51265
rect 26220 51180 26416 51183
rect 26083 51178 26416 51180
rect 26017 47642 26416 51178
rect 26017 47638 26306 47642
rect 26017 47556 26026 47638
rect 26085 47556 26164 47638
rect 26223 47560 26306 47638
rect 26365 47560 26416 47642
rect 26223 47556 26416 47560
rect 26017 46002 26416 47556
rect 26017 46000 26174 46002
rect 26017 45918 26034 46000
rect 26093 45920 26174 46000
rect 26233 46001 26416 46002
rect 26233 45920 26325 46001
rect 26093 45919 26325 45920
rect 26384 45919 26416 46001
rect 26093 45918 26416 45919
rect 26017 42866 26416 45918
rect 36836 52572 37235 55873
rect 37522 53623 37921 55873
rect 37522 53606 37932 53623
rect 37522 53603 37849 53606
rect 37522 53598 37700 53603
rect 37522 53503 37541 53598
rect 37618 53508 37700 53598
rect 37777 53511 37849 53603
rect 37926 53511 37932 53606
rect 37777 53508 37932 53511
rect 37618 53503 37932 53508
rect 37522 53430 37932 53503
rect 37522 53427 37846 53430
rect 37522 53422 37697 53427
rect 37522 53327 37538 53422
rect 37615 53332 37697 53422
rect 37774 53335 37846 53427
rect 37923 53335 37932 53430
rect 37774 53332 37932 53335
rect 37615 53327 37932 53332
rect 37522 53271 37932 53327
rect 37522 53268 37848 53271
rect 37522 53263 37699 53268
rect 37522 53168 37540 53263
rect 37617 53173 37699 53263
rect 37776 53176 37848 53268
rect 37925 53176 37932 53271
rect 37776 53173 37932 53176
rect 37617 53168 37932 53173
rect 37522 53113 37932 53168
rect 37522 53110 37847 53113
rect 37522 53105 37698 53110
rect 37522 53010 37539 53105
rect 37616 53015 37698 53105
rect 37775 53018 37847 53110
rect 37924 53018 37932 53113
rect 37775 53015 37932 53018
rect 37616 53010 37932 53015
rect 37522 53000 37932 53010
rect 36836 52555 37250 52572
rect 36836 52552 37167 52555
rect 36836 52547 37018 52552
rect 36836 52452 36859 52547
rect 36936 52457 37018 52547
rect 37095 52460 37167 52552
rect 37244 52460 37250 52555
rect 37095 52457 37250 52460
rect 36936 52452 37250 52457
rect 36836 52379 37250 52452
rect 36836 52376 37164 52379
rect 36836 52371 37015 52376
rect 36836 52276 36856 52371
rect 36933 52281 37015 52371
rect 37092 52284 37164 52376
rect 37241 52284 37250 52379
rect 37092 52281 37250 52284
rect 36933 52276 37250 52281
rect 36836 52220 37250 52276
rect 36836 52217 37166 52220
rect 36836 52212 37017 52217
rect 36836 52117 36858 52212
rect 36935 52122 37017 52212
rect 37094 52125 37166 52217
rect 37243 52125 37250 52220
rect 37094 52122 37250 52125
rect 36935 52117 37250 52122
rect 36836 52062 37250 52117
rect 36836 52059 37165 52062
rect 36836 52054 37016 52059
rect 36836 51959 36857 52054
rect 36934 51964 37016 52054
rect 37093 51967 37165 52059
rect 37242 51967 37250 52062
rect 37093 51964 37250 51967
rect 36934 51959 37250 51964
rect 36836 51949 37250 51959
rect 35573 45231 35681 45266
rect 35573 45136 35592 45231
rect 35669 45136 35681 45231
rect 35573 45055 35681 45136
rect 35573 44960 35589 45055
rect 35666 44960 35681 45055
rect 35573 44896 35681 44960
rect 35573 44801 35591 44896
rect 35668 44801 35681 44896
rect 35573 44738 35681 44801
rect 35573 44643 35590 44738
rect 35667 44643 35681 44738
rect 26017 42861 26169 42866
rect 26017 42786 26028 42861
rect 26087 42791 26169 42861
rect 26228 42865 26416 42866
rect 26228 42791 26323 42865
rect 26087 42790 26323 42791
rect 26382 42790 26416 42865
rect 26087 42786 26416 42790
rect 26017 39265 26416 42786
rect 35370 44191 35475 44248
rect 35370 44096 35389 44191
rect 35466 44096 35475 44191
rect 35370 44015 35475 44096
rect 35370 43920 35386 44015
rect 35463 43920 35475 44015
rect 35370 43856 35475 43920
rect 35370 43761 35388 43856
rect 35465 43761 35475 43856
rect 35370 43698 35475 43761
rect 35370 43603 35387 43698
rect 35464 43603 35475 43698
rect 35370 42687 35475 43603
rect 35573 42608 35681 44643
rect 36836 44203 37235 51949
rect 37522 45246 37921 53000
rect 37522 45229 37932 45246
rect 37522 45226 37849 45229
rect 37522 45221 37700 45226
rect 37522 45126 37541 45221
rect 37618 45131 37700 45221
rect 37777 45134 37849 45226
rect 37926 45134 37932 45229
rect 37777 45131 37932 45134
rect 37618 45126 37932 45131
rect 37522 45053 37932 45126
rect 37522 45050 37846 45053
rect 37522 45045 37697 45050
rect 37522 44950 37538 45045
rect 37615 44955 37697 45045
rect 37774 44958 37846 45050
rect 37923 44958 37932 45053
rect 37774 44955 37932 44958
rect 37615 44950 37932 44955
rect 37522 44894 37932 44950
rect 37522 44891 37848 44894
rect 37522 44886 37699 44891
rect 37522 44791 37540 44886
rect 37617 44796 37699 44886
rect 37776 44799 37848 44891
rect 37925 44799 37932 44894
rect 37776 44796 37932 44799
rect 37617 44791 37932 44796
rect 37522 44736 37932 44791
rect 37522 44733 37847 44736
rect 37522 44728 37698 44733
rect 37522 44633 37539 44728
rect 37616 44638 37698 44728
rect 37775 44641 37847 44733
rect 37924 44641 37932 44736
rect 37775 44638 37932 44641
rect 37616 44633 37932 44638
rect 37522 44623 37932 44633
rect 36836 44186 37246 44203
rect 36836 44183 37163 44186
rect 36836 44178 37014 44183
rect 36836 44083 36855 44178
rect 36932 44088 37014 44178
rect 37091 44091 37163 44183
rect 37240 44091 37246 44186
rect 37091 44088 37246 44091
rect 36932 44083 37246 44088
rect 36836 44010 37246 44083
rect 36836 44007 37160 44010
rect 36836 44002 37011 44007
rect 36836 43907 36852 44002
rect 36929 43912 37011 44002
rect 37088 43915 37160 44007
rect 37237 43915 37246 44010
rect 37088 43912 37246 43915
rect 36929 43907 37246 43912
rect 36836 43851 37246 43907
rect 36836 43848 37162 43851
rect 36836 43843 37013 43848
rect 36836 43748 36854 43843
rect 36931 43753 37013 43843
rect 37090 43756 37162 43848
rect 37239 43756 37246 43851
rect 37090 43753 37246 43756
rect 36931 43748 37246 43753
rect 36836 43693 37246 43748
rect 36836 43690 37161 43693
rect 36836 43685 37012 43690
rect 36836 43590 36853 43685
rect 36930 43595 37012 43685
rect 37089 43598 37161 43690
rect 37238 43598 37246 43693
rect 37089 43595 37246 43598
rect 36930 43590 37246 43595
rect 36836 43580 37246 43590
rect 28791 41689 28914 41703
rect 28791 41610 28811 41689
rect 28902 41610 28914 41689
rect 28791 41537 28914 41610
rect 28791 41458 28807 41537
rect 28898 41458 28914 41537
rect 28791 41446 28914 41458
rect 31116 41326 31172 41657
rect 27286 40613 27390 40627
rect 27286 40558 27306 40613
rect 27364 40558 27390 40613
rect 27286 40469 27390 40558
rect 27286 40414 27311 40469
rect 27369 40414 27390 40469
rect 31119 40418 31175 40639
rect 27286 40343 27390 40414
rect 27286 40294 27309 40343
rect 26017 39262 26181 39265
rect 26017 39199 26049 39262
rect 26109 39202 26181 39262
rect 26241 39262 26416 39265
rect 26241 39202 26315 39262
rect 26109 39199 26315 39202
rect 26375 39199 26416 39262
rect 26017 34406 26416 39199
rect 26017 34311 26028 34406
rect 26101 34311 26176 34406
rect 26249 34311 26330 34406
rect 26403 34311 26416 34406
rect 26017 30765 26416 34311
rect 26017 30762 26181 30765
rect 26017 30699 26049 30762
rect 26109 30702 26181 30762
rect 26241 30762 26416 30765
rect 26241 30702 26315 30762
rect 26109 30699 26315 30702
rect 26375 30699 26416 30762
rect 26017 26165 26416 30699
rect 26017 26162 26165 26165
rect 26017 26087 26025 26162
rect 26084 26090 26165 26162
rect 26224 26090 26312 26165
rect 26371 26090 26416 26165
rect 26084 26087 26416 26090
rect 26017 21180 26416 26087
rect 26017 21177 26174 21180
rect 26017 21114 26042 21177
rect 26102 21117 26174 21177
rect 26234 21177 26416 21180
rect 26234 21117 26308 21177
rect 26102 21114 26308 21117
rect 26368 21114 26416 21177
rect 26017 16954 26416 21114
rect 27284 40288 27309 40294
rect 27367 40294 27390 40343
rect 27367 40288 27402 40294
rect 27284 35598 27402 40288
rect 28461 39732 28584 39746
rect 28461 39653 28481 39732
rect 28572 39653 28584 39732
rect 28461 39580 28584 39653
rect 28461 39501 28477 39580
rect 28568 39501 28584 39580
rect 28461 39489 28584 39501
rect 27929 38873 28138 38892
rect 27929 38805 27946 38873
rect 28014 38872 28138 38873
rect 28014 38806 28070 38872
rect 28136 38806 28138 38872
rect 28014 38805 28138 38806
rect 27929 38783 28138 38805
rect 27284 35524 27309 35598
rect 27388 35524 27402 35598
rect 27284 35415 27402 35524
rect 27284 35341 27308 35415
rect 27387 35341 27402 35415
rect 27284 17813 27402 35341
rect 27537 32161 27700 32190
rect 27537 32083 27573 32161
rect 27664 32083 27700 32161
rect 27537 31954 27700 32083
rect 27537 31876 27582 31954
rect 27673 31876 27700 31954
rect 27537 27887 27700 31876
rect 27936 30569 28024 38783
rect 28286 38345 28404 38385
rect 28286 38270 28308 38345
rect 28383 38270 28404 38345
rect 28286 38197 28404 38270
rect 28286 38120 28307 38197
rect 28384 38120 28404 38197
rect 27918 30555 28036 30569
rect 27918 30469 27932 30555
rect 28018 30469 28036 30555
rect 27918 30393 28036 30469
rect 27918 30305 27936 30393
rect 28024 30305 28036 30393
rect 27918 30282 28036 30305
rect 28286 29890 28404 38120
rect 31168 38025 31225 38297
rect 35592 37016 35700 37045
rect 35592 36921 35612 37016
rect 35689 36921 35700 37016
rect 35592 36840 35700 36921
rect 35592 36745 35609 36840
rect 35686 36745 35700 36840
rect 35592 36681 35700 36745
rect 35592 36586 35611 36681
rect 35688 36586 35700 36681
rect 35592 36523 35700 36586
rect 35592 36428 35610 36523
rect 35687 36428 35700 36523
rect 35389 35760 35494 35799
rect 35389 35665 35407 35760
rect 35484 35665 35494 35760
rect 35389 35584 35494 35665
rect 35389 35489 35404 35584
rect 35481 35489 35494 35584
rect 35389 35425 35494 35489
rect 35389 35330 35406 35425
rect 35483 35330 35494 35425
rect 35389 35267 35494 35330
rect 35389 35172 35405 35267
rect 35482 35172 35494 35267
rect 35389 34188 35494 35172
rect 35592 34136 35700 36428
rect 36836 35776 37235 43580
rect 37522 37023 37921 44623
rect 37522 37006 37932 37023
rect 37522 37003 37849 37006
rect 37522 36998 37700 37003
rect 37522 36903 37541 36998
rect 37618 36908 37700 36998
rect 37777 36911 37849 37003
rect 37926 36911 37932 37006
rect 37777 36908 37932 36911
rect 37618 36903 37932 36908
rect 37522 36830 37932 36903
rect 37522 36827 37846 36830
rect 37522 36822 37697 36827
rect 37522 36727 37538 36822
rect 37615 36732 37697 36822
rect 37774 36735 37846 36827
rect 37923 36735 37932 36830
rect 37774 36732 37932 36735
rect 37615 36727 37932 36732
rect 37522 36671 37932 36727
rect 37522 36668 37848 36671
rect 37522 36663 37699 36668
rect 37522 36568 37540 36663
rect 37617 36573 37699 36663
rect 37776 36576 37848 36668
rect 37925 36576 37932 36671
rect 37776 36573 37932 36576
rect 37617 36568 37932 36573
rect 37522 36513 37932 36568
rect 37522 36510 37847 36513
rect 37522 36505 37698 36510
rect 37522 36410 37539 36505
rect 37616 36415 37698 36505
rect 37775 36418 37847 36510
rect 37924 36418 37932 36513
rect 37775 36415 37932 36418
rect 37616 36410 37932 36415
rect 37522 36400 37932 36410
rect 36832 35759 37242 35776
rect 36832 35756 37159 35759
rect 36832 35751 37010 35756
rect 36832 35656 36851 35751
rect 36928 35661 37010 35751
rect 37087 35664 37159 35756
rect 37236 35664 37242 35759
rect 37087 35661 37242 35664
rect 36928 35656 37242 35661
rect 36832 35583 37242 35656
rect 36832 35580 37156 35583
rect 36832 35575 37007 35580
rect 36832 35480 36848 35575
rect 36925 35485 37007 35575
rect 37084 35488 37156 35580
rect 37233 35488 37242 35583
rect 37084 35485 37242 35488
rect 36925 35480 37242 35485
rect 36832 35424 37242 35480
rect 36832 35421 37158 35424
rect 36832 35416 37009 35421
rect 36832 35321 36850 35416
rect 36927 35326 37009 35416
rect 37086 35329 37158 35421
rect 37235 35329 37242 35424
rect 37086 35326 37242 35329
rect 36927 35321 37242 35326
rect 36832 35266 37242 35321
rect 36832 35263 37157 35266
rect 36832 35258 37008 35263
rect 36832 35163 36849 35258
rect 36926 35168 37008 35258
rect 37085 35171 37157 35263
rect 37234 35171 37242 35266
rect 37085 35168 37242 35171
rect 36926 35163 37242 35168
rect 36832 35153 37242 35163
rect 28805 33195 28928 33209
rect 28805 33116 28825 33195
rect 28916 33116 28928 33195
rect 28805 33043 28928 33116
rect 28805 32964 28821 33043
rect 28912 32964 28928 33043
rect 28805 32952 28928 32964
rect 31135 32438 31191 32661
rect 31138 31923 31194 32141
rect 28530 31229 28653 31243
rect 28530 31150 28550 31229
rect 28641 31150 28653 31229
rect 28530 31077 28653 31150
rect 28530 30998 28546 31077
rect 28637 30998 28653 31077
rect 28530 30986 28653 30998
rect 28286 29848 28569 29890
rect 28286 29773 28460 29848
rect 28540 29773 28569 29848
rect 28286 29772 28569 29773
rect 28441 29684 28564 29772
rect 28441 29607 28462 29684
rect 28539 29607 28564 29684
rect 28441 29587 28564 29607
rect 27539 27809 27685 27887
rect 27539 27714 27567 27809
rect 27650 27714 27685 27809
rect 27539 27576 27685 27714
rect 27539 27481 27571 27576
rect 27654 27481 27685 27576
rect 27539 27425 27685 27481
rect 28441 27323 28560 29587
rect 31187 29573 31244 29799
rect 28761 29315 28819 29479
rect 28733 28856 28848 29315
rect 28731 28833 28849 28856
rect 28731 28749 28754 28833
rect 28820 28749 28849 28833
rect 28731 28696 28849 28749
rect 28731 28612 28756 28696
rect 28822 28612 28849 28696
rect 28731 28579 28849 28612
rect 28441 27292 28566 27323
rect 28441 27197 28462 27292
rect 28557 27197 28566 27292
rect 28441 27136 28566 27197
rect 28441 27043 28463 27136
rect 28556 27043 28566 27136
rect 28441 27009 28566 27043
rect 28441 26510 28560 27009
rect 28166 26494 28576 26510
rect 28166 26493 28441 26494
rect 28166 26376 28178 26493
rect 28295 26376 28441 26493
rect 28166 26375 28441 26376
rect 28560 26375 28576 26494
rect 28166 26361 28576 26375
rect 28733 25949 28848 28579
rect 36836 27368 37235 35153
rect 37522 28466 37921 36400
rect 37522 28449 37936 28466
rect 37522 28446 37853 28449
rect 37522 28441 37704 28446
rect 37522 28346 37545 28441
rect 37622 28351 37704 28441
rect 37781 28354 37853 28446
rect 37930 28354 37936 28449
rect 37781 28351 37936 28354
rect 37622 28346 37936 28351
rect 37522 28273 37936 28346
rect 37522 28270 37850 28273
rect 37522 28265 37701 28270
rect 37522 28170 37542 28265
rect 37619 28175 37701 28265
rect 37778 28178 37850 28270
rect 37927 28178 37936 28273
rect 37778 28175 37936 28178
rect 37619 28170 37936 28175
rect 37522 28114 37936 28170
rect 37522 28111 37852 28114
rect 37522 28106 37703 28111
rect 37522 28011 37544 28106
rect 37621 28016 37703 28106
rect 37780 28019 37852 28111
rect 37929 28019 37936 28114
rect 37780 28016 37936 28019
rect 37621 28011 37936 28016
rect 37522 27956 37936 28011
rect 37522 27953 37851 27956
rect 37522 27948 37702 27953
rect 37522 27853 37543 27948
rect 37620 27858 37702 27948
rect 37779 27861 37851 27953
rect 37928 27861 37936 27956
rect 37779 27858 37936 27861
rect 37620 27853 37936 27858
rect 37522 27843 37936 27853
rect 36832 27351 37242 27368
rect 36832 27348 37159 27351
rect 36832 27343 37010 27348
rect 36832 27248 36851 27343
rect 36928 27253 37010 27343
rect 37087 27256 37159 27348
rect 37236 27256 37242 27351
rect 37087 27253 37242 27256
rect 36928 27248 37242 27253
rect 36832 27175 37242 27248
rect 36832 27172 37156 27175
rect 36832 27167 37007 27172
rect 36832 27072 36848 27167
rect 36925 27077 37007 27167
rect 37084 27080 37156 27172
rect 37233 27080 37242 27175
rect 37084 27077 37242 27080
rect 36925 27072 37242 27077
rect 36832 27016 37242 27072
rect 36832 27013 37158 27016
rect 36832 27008 37009 27013
rect 36832 26913 36850 27008
rect 36927 26918 37009 27008
rect 37086 26921 37158 27013
rect 37235 26921 37242 27016
rect 37086 26918 37242 26921
rect 36927 26913 37242 26918
rect 36832 26858 37242 26913
rect 36832 26855 37157 26858
rect 36832 26850 37008 26855
rect 36832 26755 36849 26850
rect 36926 26760 37008 26850
rect 37085 26763 37157 26855
rect 37234 26763 37242 26858
rect 37085 26760 37242 26763
rect 36926 26755 37242 26760
rect 36832 26745 37242 26755
rect 28708 25948 28848 25949
rect 28572 25939 28848 25948
rect 28548 25924 28848 25939
rect 28548 25824 28588 25924
rect 28572 25815 28588 25824
rect 28697 25824 28848 25924
rect 28697 25815 28712 25824
rect 28572 25654 28712 25815
rect 28572 25543 28587 25654
rect 28698 25543 28712 25654
rect 28572 25536 28712 25543
rect 28587 25534 28698 25536
rect 29510 23944 29566 24073
rect 28896 22703 28952 22869
rect 29960 21655 30016 21846
rect 28463 21538 28574 21569
rect 28463 21483 28493 21538
rect 28548 21483 28574 21538
rect 28463 21419 28574 21483
rect 28463 21364 28493 21419
rect 28548 21364 28574 21419
rect 28463 20546 28574 21364
rect 28455 20531 28838 20546
rect 28455 20422 28464 20531
rect 28573 20422 28713 20531
rect 28822 20422 28838 20531
rect 28455 20408 28838 20422
rect 35605 19440 35706 19442
rect 35592 19416 35706 19440
rect 35592 19321 35623 19416
rect 35700 19321 35706 19416
rect 35592 19240 35706 19321
rect 35592 19145 35620 19240
rect 35697 19145 35706 19240
rect 35592 19081 35706 19145
rect 35592 18986 35622 19081
rect 35699 18986 35706 19081
rect 35592 18923 35706 18986
rect 35592 18828 35621 18923
rect 35698 18828 35706 18923
rect 35592 18805 35706 18828
rect 27205 17778 27402 17813
rect 27205 17660 27251 17778
rect 27369 17660 27402 17778
rect 27205 17543 27402 17660
rect 27205 17425 27246 17543
rect 27364 17425 27402 17543
rect 27205 17388 27402 17425
rect 35389 18352 35494 18368
rect 35389 18326 35500 18352
rect 35389 18231 35417 18326
rect 35494 18231 35500 18326
rect 35389 18150 35500 18231
rect 35389 18055 35414 18150
rect 35491 18055 35500 18150
rect 35389 17991 35500 18055
rect 35389 17896 35416 17991
rect 35493 17896 35500 17991
rect 35389 17833 35500 17896
rect 35389 17738 35415 17833
rect 35492 17738 35500 17833
rect 35389 17715 35500 17738
rect 26017 16951 26319 16954
rect 26017 16946 26180 16951
rect 26017 16873 26025 16946
rect 26082 16878 26180 16946
rect 26237 16881 26319 16951
rect 26376 16881 26416 16954
rect 26237 16878 26416 16881
rect 26082 16873 26416 16878
rect 26017 14600 26416 16873
rect 35389 16582 35494 17715
rect 35592 16597 35700 18805
rect 36836 18333 37235 26745
rect 37522 19415 37921 27843
rect 37522 19398 37932 19415
rect 37522 19395 37849 19398
rect 37522 19390 37700 19395
rect 37522 19295 37541 19390
rect 37618 19300 37700 19390
rect 37777 19303 37849 19395
rect 37926 19303 37932 19398
rect 37777 19300 37932 19303
rect 37618 19295 37932 19300
rect 37522 19222 37932 19295
rect 37522 19219 37846 19222
rect 37522 19214 37697 19219
rect 37522 19119 37538 19214
rect 37615 19124 37697 19214
rect 37774 19127 37846 19219
rect 37923 19127 37932 19222
rect 37774 19124 37932 19127
rect 37615 19119 37932 19124
rect 37522 19063 37932 19119
rect 37522 19060 37848 19063
rect 37522 19055 37699 19060
rect 37522 18960 37540 19055
rect 37617 18965 37699 19055
rect 37776 18968 37848 19060
rect 37925 18968 37932 19063
rect 37776 18965 37932 18968
rect 37617 18960 37932 18965
rect 37522 18905 37932 18960
rect 37522 18902 37847 18905
rect 37522 18897 37698 18902
rect 37522 18802 37539 18897
rect 37616 18807 37698 18897
rect 37775 18810 37847 18902
rect 37924 18810 37932 18905
rect 37775 18807 37932 18810
rect 37616 18802 37932 18807
rect 37522 18792 37932 18802
rect 36836 18316 37246 18333
rect 36836 18313 37163 18316
rect 36836 18308 37014 18313
rect 36836 18213 36855 18308
rect 36932 18218 37014 18308
rect 37091 18221 37163 18313
rect 37240 18221 37246 18316
rect 37091 18218 37246 18221
rect 36932 18213 37246 18218
rect 36836 18140 37246 18213
rect 36836 18137 37160 18140
rect 36836 18132 37011 18137
rect 36836 18037 36852 18132
rect 36929 18042 37011 18132
rect 37088 18045 37160 18137
rect 37237 18045 37246 18140
rect 37088 18042 37246 18045
rect 36929 18037 37246 18042
rect 36836 17981 37246 18037
rect 36836 17978 37162 17981
rect 36836 17973 37013 17978
rect 36836 17878 36854 17973
rect 36931 17883 37013 17973
rect 37090 17886 37162 17978
rect 37239 17886 37246 17981
rect 37090 17883 37246 17886
rect 36931 17878 37246 17883
rect 36836 17823 37246 17878
rect 36836 17820 37161 17823
rect 36836 17815 37012 17820
rect 36836 17720 36853 17815
rect 36930 17725 37012 17815
rect 37089 17728 37161 17820
rect 37238 17728 37246 17823
rect 37089 17725 37246 17728
rect 36930 17720 37246 17725
rect 36836 17710 37246 17720
rect 28851 15585 28938 15606
rect 28851 15529 28864 15585
rect 28920 15529 28938 15585
rect 28851 15474 28938 15529
rect 28851 15418 28860 15474
rect 28916 15418 28938 15474
rect 28851 15403 28938 15418
rect 31135 14882 31191 15089
rect 26017 14597 26195 14600
rect 26017 14534 26063 14597
rect 26123 14537 26195 14597
rect 26255 14597 26416 14600
rect 26255 14537 26329 14597
rect 26123 14534 26329 14537
rect 26389 14534 26416 14597
rect 26017 13245 26416 14534
rect 31138 14372 31194 14620
rect 28527 13723 28614 13744
rect 28527 13667 28540 13723
rect 28596 13667 28614 13723
rect 28527 13612 28614 13667
rect 28527 13556 28536 13612
rect 28592 13556 28614 13612
rect 28527 13541 28614 13556
rect 26017 13242 26187 13245
rect 26017 13179 26055 13242
rect 26115 13182 26187 13242
rect 26247 13242 26416 13245
rect 26247 13182 26321 13242
rect 26115 13179 26321 13182
rect 26381 13179 26416 13242
rect 26017 11526 26416 13179
rect 26017 11521 26173 11526
rect 26017 11448 26033 11521
rect 26090 11453 26173 11521
rect 26230 11525 26416 11526
rect 26230 11453 26325 11525
rect 26090 11452 26325 11453
rect 26382 11452 26416 11525
rect 26090 11448 26416 11452
rect 26017 4421 26416 11448
rect 26017 4411 26319 4421
rect 26017 4406 26174 4411
rect 26017 4336 26031 4406
rect 26099 4341 26174 4406
rect 26242 4351 26319 4411
rect 26387 4351 26416 4421
rect 26242 4341 26416 4351
rect 26099 4336 26416 4341
rect 26017 4266 26416 4336
rect 26017 4263 26327 4266
rect 26017 4193 26032 4263
rect 26100 4193 26176 4263
rect 26244 4196 26327 4263
rect 26395 4196 26416 4266
rect 26244 4193 26416 4196
rect 26017 1858 26416 4193
rect 26017 1855 26198 1858
rect 26017 1792 26066 1855
rect 26126 1795 26198 1855
rect 26258 1855 26416 1858
rect 26258 1795 26332 1855
rect 26126 1792 26332 1795
rect 26392 1792 26416 1855
rect 26017 508 26416 1792
rect 26017 505 26187 508
rect 26017 442 26055 505
rect 26115 445 26187 505
rect 26247 505 26416 508
rect 26247 445 26321 505
rect 26115 442 26321 445
rect 26381 442 26416 505
rect 26017 -793 26416 442
rect 26017 -795 26319 -793
rect 26017 -799 26183 -795
rect 26017 -898 26033 -799
rect 26100 -894 26183 -799
rect 26250 -892 26319 -795
rect 26386 -892 26416 -793
rect 26250 -894 26416 -892
rect 26100 -898 26416 -894
rect 26017 -4746 26416 -898
rect 26017 -4824 26022 -4746
rect 26093 -4747 26416 -4746
rect 26093 -4824 26177 -4747
rect 26017 -4825 26177 -4824
rect 26248 -4750 26416 -4747
rect 26248 -4825 26330 -4750
rect 26017 -4828 26330 -4825
rect 26401 -4828 26416 -4750
rect 26017 -9723 26416 -4828
rect 26017 -9726 26183 -9723
rect 26017 -9789 26051 -9726
rect 26111 -9786 26183 -9726
rect 26243 -9726 26416 -9723
rect 26243 -9786 26317 -9726
rect 26111 -9789 26317 -9786
rect 26377 -9789 26416 -9726
rect 26017 -13571 26416 -9789
rect 26017 -13579 26180 -13571
rect 26017 -13657 26027 -13579
rect 26088 -13649 26180 -13579
rect 26241 -13572 26416 -13571
rect 26241 -13649 26339 -13572
rect 26088 -13650 26339 -13649
rect 26400 -13650 26416 -13572
rect 26088 -13657 26416 -13650
rect 26017 -15897 26416 -13657
rect 26017 -15900 26173 -15897
rect 26017 -15963 26041 -15900
rect 26101 -15960 26173 -15900
rect 26233 -15900 26416 -15897
rect 26233 -15960 26307 -15900
rect 26101 -15963 26307 -15960
rect 26367 -15963 26416 -15900
rect 26017 -17246 26416 -15963
rect 26017 -17249 26173 -17246
rect 26017 -17312 26041 -17249
rect 26101 -17309 26173 -17249
rect 26233 -17249 26416 -17246
rect 26233 -17309 26307 -17249
rect 26101 -17312 26307 -17309
rect 26367 -17312 26416 -17249
rect 26017 -18951 26416 -17312
rect 27801 12849 27912 12878
rect 27801 12783 27828 12849
rect 27894 12783 27912 12849
rect 27801 12694 27912 12783
rect 27801 12628 27828 12694
rect 27894 12628 27912 12694
rect 27801 111 27912 12628
rect 28107 12348 28204 12349
rect 28107 12326 28205 12348
rect 28107 12251 28119 12326
rect 28194 12251 28205 12326
rect 28107 12152 28205 12251
rect 28107 12075 28118 12152
rect 28195 12075 28205 12152
rect 28107 12067 28205 12075
rect 27801 43 27820 111
rect 27888 43 27912 111
rect 27801 -75 27912 43
rect 27801 -141 27821 -75
rect 27887 -141 27912 -75
rect 27801 -4956 27912 -141
rect 28108 -399 28205 12067
rect 31187 12033 31244 12283
rect 35365 7418 35473 7429
rect 35365 7392 35474 7418
rect 35365 7297 35391 7392
rect 35468 7297 35474 7392
rect 35365 7216 35474 7297
rect 35365 7121 35388 7216
rect 35465 7121 35474 7216
rect 35365 7057 35474 7121
rect 35365 6962 35390 7057
rect 35467 6962 35474 7057
rect 35365 6899 35474 6962
rect 35365 6804 35389 6899
rect 35466 6804 35474 6899
rect 35365 6781 35474 6804
rect 35162 6181 35267 6208
rect 35162 6155 35273 6181
rect 35162 6060 35190 6155
rect 35267 6060 35273 6155
rect 35162 5979 35273 6060
rect 35162 5884 35187 5979
rect 35264 5884 35273 5979
rect 35162 5820 35273 5884
rect 35162 5725 35189 5820
rect 35266 5725 35273 5820
rect 35162 5662 35273 5725
rect 35162 5567 35188 5662
rect 35265 5567 35273 5662
rect 35162 5544 35273 5567
rect 35162 3821 35267 5544
rect 35365 3868 35473 6781
rect 36836 6176 37235 17710
rect 37522 7396 37921 18792
rect 37522 7379 37940 7396
rect 37522 7376 37857 7379
rect 37522 7371 37708 7376
rect 37522 7276 37549 7371
rect 37626 7281 37708 7371
rect 37785 7284 37857 7376
rect 37934 7284 37940 7379
rect 37785 7281 37940 7284
rect 37626 7276 37940 7281
rect 37522 7203 37940 7276
rect 37522 7200 37854 7203
rect 37522 7195 37705 7200
rect 37522 7100 37546 7195
rect 37623 7105 37705 7195
rect 37782 7108 37854 7200
rect 37931 7108 37940 7203
rect 37782 7105 37940 7108
rect 37623 7100 37940 7105
rect 37522 7044 37940 7100
rect 37522 7041 37856 7044
rect 37522 7036 37707 7041
rect 37522 6941 37548 7036
rect 37625 6946 37707 7036
rect 37784 6949 37856 7041
rect 37933 6949 37940 7044
rect 37784 6946 37940 6949
rect 37625 6941 37940 6946
rect 37522 6886 37940 6941
rect 37522 6883 37855 6886
rect 37522 6878 37706 6883
rect 37522 6783 37547 6878
rect 37624 6788 37706 6878
rect 37783 6791 37855 6883
rect 37932 6791 37940 6886
rect 37783 6788 37940 6791
rect 37624 6783 37940 6788
rect 37522 6773 37940 6783
rect 36836 6159 37250 6176
rect 36836 6156 37167 6159
rect 36836 6151 37018 6156
rect 36836 6056 36859 6151
rect 36936 6061 37018 6151
rect 37095 6064 37167 6156
rect 37244 6064 37250 6159
rect 37095 6061 37250 6064
rect 36936 6056 37250 6061
rect 36836 5983 37250 6056
rect 36836 5980 37164 5983
rect 36836 5975 37015 5980
rect 36836 5880 36856 5975
rect 36933 5885 37015 5975
rect 37092 5888 37164 5980
rect 37241 5888 37250 5983
rect 37092 5885 37250 5888
rect 36933 5880 37250 5885
rect 36836 5824 37250 5880
rect 36836 5821 37166 5824
rect 36836 5816 37017 5821
rect 36836 5721 36858 5816
rect 36935 5726 37017 5816
rect 37094 5729 37166 5821
rect 37243 5729 37250 5824
rect 37094 5726 37250 5729
rect 36935 5721 37250 5726
rect 36836 5666 37250 5721
rect 36836 5663 37165 5666
rect 36836 5658 37016 5663
rect 36836 5563 36857 5658
rect 36934 5568 37016 5658
rect 37093 5571 37165 5663
rect 37242 5571 37250 5666
rect 37093 5568 37250 5571
rect 36934 5563 37250 5568
rect 36836 5553 37250 5563
rect 28609 2863 28696 2884
rect 28609 2807 28622 2863
rect 28678 2807 28696 2863
rect 28609 2752 28696 2807
rect 28609 2696 28618 2752
rect 28674 2696 28696 2752
rect 28609 2681 28696 2696
rect 30908 2101 30964 2320
rect 30917 1628 30973 1882
rect 28335 951 28422 972
rect 28335 895 28348 951
rect 28404 895 28422 951
rect 28335 840 28422 895
rect 28335 784 28344 840
rect 28400 784 28422 840
rect 28335 769 28422 784
rect 28107 -418 28206 -399
rect 28107 -493 28121 -418
rect 28197 -493 28206 -418
rect 28107 -563 28206 -493
rect 28107 -640 28118 -563
rect 28195 -640 28206 -563
rect 28107 -659 28206 -640
rect 28108 -4397 28205 -659
rect 30960 -731 31017 -464
rect 36836 -3525 37235 5553
rect 37522 -2455 37921 6773
rect 37522 -2472 37932 -2455
rect 37522 -2475 37849 -2472
rect 37522 -2480 37700 -2475
rect 37522 -2575 37541 -2480
rect 37618 -2570 37700 -2480
rect 37777 -2567 37849 -2475
rect 37926 -2567 37932 -2472
rect 37777 -2570 37932 -2567
rect 37618 -2575 37932 -2570
rect 37522 -2648 37932 -2575
rect 37522 -2651 37846 -2648
rect 37522 -2656 37697 -2651
rect 37522 -2751 37538 -2656
rect 37615 -2746 37697 -2656
rect 37774 -2743 37846 -2651
rect 37923 -2743 37932 -2648
rect 37774 -2746 37932 -2743
rect 37615 -2751 37932 -2746
rect 37522 -2807 37932 -2751
rect 37522 -2810 37848 -2807
rect 37522 -2815 37699 -2810
rect 37522 -2910 37540 -2815
rect 37617 -2905 37699 -2815
rect 37776 -2902 37848 -2810
rect 37925 -2902 37932 -2807
rect 37776 -2905 37932 -2902
rect 37617 -2910 37932 -2905
rect 37522 -2965 37932 -2910
rect 37522 -2968 37847 -2965
rect 37522 -2973 37698 -2968
rect 37522 -3068 37539 -2973
rect 37616 -3063 37698 -2973
rect 37775 -3060 37847 -2968
rect 37924 -3060 37932 -2965
rect 37775 -3063 37932 -3060
rect 37616 -3068 37932 -3063
rect 37522 -3078 37932 -3068
rect 36832 -3542 37242 -3525
rect 36832 -3545 37159 -3542
rect 36832 -3550 37010 -3545
rect 36832 -3645 36851 -3550
rect 36928 -3640 37010 -3550
rect 37087 -3637 37159 -3545
rect 37236 -3637 37242 -3542
rect 37087 -3640 37242 -3637
rect 36928 -3645 37242 -3640
rect 36832 -3718 37242 -3645
rect 36832 -3721 37156 -3718
rect 36832 -3726 37007 -3721
rect 36832 -3821 36848 -3726
rect 36925 -3816 37007 -3726
rect 37084 -3813 37156 -3721
rect 37233 -3813 37242 -3718
rect 37084 -3816 37242 -3813
rect 36925 -3821 37242 -3816
rect 36832 -3877 37242 -3821
rect 36832 -3880 37158 -3877
rect 36832 -3885 37009 -3880
rect 36832 -3980 36850 -3885
rect 36927 -3975 37009 -3885
rect 37086 -3972 37158 -3880
rect 37235 -3972 37242 -3877
rect 37086 -3975 37242 -3972
rect 36927 -3980 37242 -3975
rect 36832 -4035 37242 -3980
rect 36832 -4038 37157 -4035
rect 36832 -4043 37008 -4038
rect 36832 -4138 36849 -4043
rect 36926 -4133 37008 -4043
rect 37085 -4130 37157 -4038
rect 37234 -4130 37242 -4035
rect 37085 -4133 37242 -4130
rect 36926 -4138 37242 -4133
rect 36832 -4148 37242 -4138
rect 28098 -4423 28444 -4397
rect 28098 -4488 28133 -4423
rect 28197 -4426 28444 -4423
rect 28197 -4488 28315 -4426
rect 28098 -4491 28315 -4488
rect 28379 -4491 28444 -4426
rect 28098 -4515 28444 -4491
rect 27801 -5031 27820 -4956
rect 27892 -5031 27912 -4956
rect 27801 -5133 27912 -5031
rect 27801 -5208 27815 -5133
rect 27887 -5208 27912 -5133
rect 27801 -17639 27912 -5208
rect 27801 -17705 27827 -17639
rect 27893 -17705 27912 -17639
rect 27801 -17804 27912 -17705
rect 27801 -17872 27826 -17804
rect 27894 -17872 27912 -17804
rect 27801 -17980 27912 -17872
rect 26017 -18961 26321 -18951
rect 26017 -18970 26187 -18961
rect 26017 -19048 26035 -18970
rect 26096 -19039 26187 -18970
rect 26248 -19029 26321 -18961
rect 26382 -19029 26416 -18951
rect 26248 -19039 26416 -19029
rect 26096 -19048 26416 -19039
rect 26017 -21624 26416 -19048
rect 26017 -21627 26307 -21624
rect 26017 -21708 26028 -21627
rect 26084 -21708 26172 -21627
rect 26228 -21705 26307 -21627
rect 26363 -21705 26416 -21624
rect 26228 -21708 26416 -21705
rect 26017 -24007 26416 -21708
rect 26017 -24010 26175 -24007
rect 26017 -24073 26043 -24010
rect 26103 -24070 26175 -24010
rect 26235 -24010 26416 -24007
rect 26235 -24070 26309 -24010
rect 26103 -24073 26309 -24070
rect 26369 -24073 26416 -24010
rect 26017 -25352 26416 -24073
rect 26017 -25355 26177 -25352
rect 26017 -25418 26045 -25355
rect 26105 -25415 26177 -25355
rect 26237 -25355 26416 -25352
rect 26237 -25415 26311 -25355
rect 26105 -25418 26311 -25415
rect 26371 -25418 26416 -25355
rect 26017 -26878 26416 -25418
rect 27804 -25702 27912 -17980
rect 27804 -25770 27825 -25702
rect 27893 -25770 27912 -25702
rect 27804 -25877 27912 -25770
rect 27804 -25943 27826 -25877
rect 27892 -25943 27912 -25877
rect 27804 -25965 27912 -25943
rect 28108 -18000 28205 -4515
rect 29530 -6954 29586 -6823
rect 28916 -8193 28972 -8041
rect 29980 -9241 30036 -9046
rect 28503 -9359 28587 -9341
rect 28503 -9416 28516 -9359
rect 28573 -9416 28587 -9359
rect 28503 -9484 28587 -9416
rect 28503 -9543 28518 -9484
rect 28577 -9543 28587 -9484
rect 28503 -11925 28587 -9543
rect 29266 -10004 29337 -9890
rect 29238 -11121 29364 -10004
rect 29218 -11130 29364 -11121
rect 29218 -11230 29254 -11130
rect 29339 -11230 29364 -11130
rect 29218 -11306 29364 -11230
rect 29218 -11406 29243 -11306
rect 29328 -11406 29364 -11306
rect 29218 -11421 29364 -11406
rect 35382 -11377 35490 -11345
rect 29218 -11426 29347 -11421
rect 35382 -11472 35400 -11377
rect 35477 -11472 35490 -11377
rect 35382 -11553 35490 -11472
rect 35382 -11648 35397 -11553
rect 35474 -11648 35490 -11553
rect 35382 -11712 35490 -11648
rect 35382 -11807 35399 -11712
rect 35476 -11807 35490 -11712
rect 35382 -11870 35490 -11807
rect 28489 -11974 28601 -11925
rect 28489 -12026 28521 -11974
rect 28576 -12026 28601 -11974
rect 28489 -12109 28601 -12026
rect 28489 -12161 28512 -12109
rect 28567 -12161 28601 -12109
rect 28489 -12182 28601 -12161
rect 35382 -11965 35398 -11870
rect 35475 -11965 35490 -11870
rect 35179 -12422 35284 -12357
rect 35179 -12517 35199 -12422
rect 35276 -12517 35284 -12422
rect 35179 -12598 35284 -12517
rect 35179 -12693 35196 -12598
rect 35273 -12693 35284 -12598
rect 35179 -12757 35284 -12693
rect 35179 -12852 35198 -12757
rect 35275 -12852 35284 -12757
rect 35179 -12915 35284 -12852
rect 35179 -13010 35197 -12915
rect 35274 -13010 35284 -12915
rect 35179 -13946 35284 -13010
rect 35382 -13887 35490 -11965
rect 36836 -12415 37235 -4148
rect 37522 -11376 37921 -3078
rect 37522 -11393 37932 -11376
rect 37522 -11396 37849 -11393
rect 37522 -11401 37700 -11396
rect 37522 -11496 37541 -11401
rect 37618 -11491 37700 -11401
rect 37777 -11488 37849 -11396
rect 37926 -11488 37932 -11393
rect 37777 -11491 37932 -11488
rect 37618 -11496 37932 -11491
rect 37522 -11569 37932 -11496
rect 37522 -11572 37846 -11569
rect 37522 -11577 37697 -11572
rect 37522 -11672 37538 -11577
rect 37615 -11667 37697 -11577
rect 37774 -11664 37846 -11572
rect 37923 -11664 37932 -11569
rect 37774 -11667 37932 -11664
rect 37615 -11672 37932 -11667
rect 37522 -11728 37932 -11672
rect 37522 -11731 37848 -11728
rect 37522 -11736 37699 -11731
rect 37522 -11831 37540 -11736
rect 37617 -11826 37699 -11736
rect 37776 -11823 37848 -11731
rect 37925 -11823 37932 -11728
rect 37776 -11826 37932 -11823
rect 37617 -11831 37932 -11826
rect 37522 -11886 37932 -11831
rect 37522 -11889 37847 -11886
rect 37522 -11894 37698 -11889
rect 37522 -11989 37539 -11894
rect 37616 -11984 37698 -11894
rect 37775 -11981 37847 -11889
rect 37924 -11981 37932 -11886
rect 37775 -11984 37932 -11981
rect 37616 -11989 37932 -11984
rect 37522 -11999 37932 -11989
rect 36836 -12432 37246 -12415
rect 36836 -12435 37163 -12432
rect 36836 -12440 37014 -12435
rect 36836 -12535 36855 -12440
rect 36932 -12530 37014 -12440
rect 37091 -12527 37163 -12435
rect 37240 -12527 37246 -12432
rect 37091 -12530 37246 -12527
rect 36932 -12535 37246 -12530
rect 36836 -12608 37246 -12535
rect 36836 -12611 37160 -12608
rect 36836 -12616 37011 -12611
rect 36836 -12711 36852 -12616
rect 36929 -12706 37011 -12616
rect 37088 -12703 37160 -12611
rect 37237 -12703 37246 -12608
rect 37088 -12706 37246 -12703
rect 36929 -12711 37246 -12706
rect 36836 -12767 37246 -12711
rect 36836 -12770 37162 -12767
rect 36836 -12775 37013 -12770
rect 36836 -12870 36854 -12775
rect 36931 -12865 37013 -12775
rect 37090 -12862 37162 -12770
rect 37239 -12862 37246 -12767
rect 37090 -12865 37246 -12862
rect 36931 -12870 37246 -12865
rect 36836 -12925 37246 -12870
rect 36836 -12928 37161 -12925
rect 36836 -12933 37012 -12928
rect 36836 -13028 36853 -12933
rect 36930 -13023 37012 -12933
rect 37089 -13020 37161 -12928
rect 37238 -13020 37246 -12925
rect 37089 -13023 37246 -13020
rect 36930 -13028 37246 -13023
rect 36836 -13038 37246 -13028
rect 28638 -14904 28725 -14883
rect 28638 -14960 28651 -14904
rect 28707 -14960 28725 -14904
rect 28638 -15015 28725 -14960
rect 28638 -15071 28647 -15015
rect 28703 -15071 28725 -15015
rect 28638 -15086 28725 -15071
rect 30925 -15625 30981 -15384
rect 30928 -16120 30984 -15918
rect 28305 -16761 28443 -16744
rect 28305 -16832 28339 -16761
rect 28410 -16832 28443 -16761
rect 28305 -16937 28443 -16832
rect 28305 -17008 28335 -16937
rect 28406 -17008 28443 -16937
rect 28305 -17018 28443 -17008
rect 28108 -18017 28214 -18000
rect 28108 -18094 28123 -18017
rect 28200 -18094 28214 -18017
rect 28108 -18166 28214 -18094
rect 28108 -18241 28124 -18166
rect 28199 -18241 28214 -18166
rect 28108 -18278 28214 -18241
rect 28108 -26099 28205 -18278
rect 30977 -18455 31034 -18214
rect 35402 -19445 35510 -19421
rect 35398 -19471 35510 -19445
rect 35398 -19566 35416 -19471
rect 35493 -19566 35510 -19471
rect 35398 -19647 35510 -19566
rect 35398 -19742 35413 -19647
rect 35490 -19742 35510 -19647
rect 35398 -19806 35510 -19742
rect 35398 -19901 35415 -19806
rect 35492 -19901 35510 -19806
rect 35398 -19964 35510 -19901
rect 35398 -20059 35414 -19964
rect 35491 -20059 35510 -19964
rect 35398 -20082 35510 -20059
rect 35199 -20487 35304 -20465
rect 35195 -20513 35304 -20487
rect 35195 -20608 35213 -20513
rect 35290 -20608 35304 -20513
rect 35195 -20689 35304 -20608
rect 35195 -20784 35210 -20689
rect 35287 -20784 35304 -20689
rect 35195 -20848 35304 -20784
rect 35195 -20943 35212 -20848
rect 35289 -20943 35304 -20848
rect 35195 -21006 35304 -20943
rect 35195 -21101 35211 -21006
rect 35288 -21101 35304 -21006
rect 35195 -21124 35304 -21101
rect 35199 -21894 35304 -21124
rect 35402 -21920 35510 -20082
rect 36836 -20498 37235 -13038
rect 37522 -19458 37921 -11999
rect 37522 -19475 37932 -19458
rect 37522 -19478 37849 -19475
rect 37522 -19483 37700 -19478
rect 37522 -19578 37541 -19483
rect 37618 -19573 37700 -19483
rect 37777 -19570 37849 -19478
rect 37926 -19570 37932 -19475
rect 37777 -19573 37932 -19570
rect 37618 -19578 37932 -19573
rect 37522 -19651 37932 -19578
rect 37522 -19654 37846 -19651
rect 37522 -19659 37697 -19654
rect 37522 -19754 37538 -19659
rect 37615 -19749 37697 -19659
rect 37774 -19746 37846 -19654
rect 37923 -19746 37932 -19651
rect 37774 -19749 37932 -19746
rect 37615 -19754 37932 -19749
rect 37522 -19810 37932 -19754
rect 37522 -19813 37848 -19810
rect 37522 -19818 37699 -19813
rect 37522 -19913 37540 -19818
rect 37617 -19908 37699 -19818
rect 37776 -19905 37848 -19813
rect 37925 -19905 37932 -19810
rect 37776 -19908 37932 -19905
rect 37617 -19913 37932 -19908
rect 37522 -19968 37932 -19913
rect 37522 -19971 37847 -19968
rect 37522 -19976 37698 -19971
rect 37522 -20071 37539 -19976
rect 37616 -20066 37698 -19976
rect 37775 -20063 37847 -19971
rect 37924 -20063 37932 -19968
rect 37775 -20066 37932 -20063
rect 37616 -20071 37932 -20066
rect 37522 -20081 37932 -20071
rect 36832 -20515 37242 -20498
rect 36832 -20518 37159 -20515
rect 36832 -20523 37010 -20518
rect 36832 -20618 36851 -20523
rect 36928 -20613 37010 -20523
rect 37087 -20610 37159 -20518
rect 37236 -20610 37242 -20515
rect 37087 -20613 37242 -20610
rect 36928 -20618 37242 -20613
rect 36832 -20691 37242 -20618
rect 36832 -20694 37156 -20691
rect 36832 -20699 37007 -20694
rect 36832 -20794 36848 -20699
rect 36925 -20789 37007 -20699
rect 37084 -20786 37156 -20694
rect 37233 -20786 37242 -20691
rect 37084 -20789 37242 -20786
rect 36925 -20794 37242 -20789
rect 36832 -20850 37242 -20794
rect 36832 -20853 37158 -20850
rect 36832 -20858 37009 -20853
rect 36832 -20953 36850 -20858
rect 36927 -20948 37009 -20858
rect 37086 -20945 37158 -20853
rect 37235 -20945 37242 -20850
rect 37086 -20948 37242 -20945
rect 36927 -20953 37242 -20948
rect 36832 -21008 37242 -20953
rect 36832 -21011 37157 -21008
rect 36832 -21016 37008 -21011
rect 36832 -21111 36849 -21016
rect 36926 -21106 37008 -21016
rect 37085 -21103 37157 -21011
rect 37234 -21103 37242 -21008
rect 37085 -21106 37242 -21103
rect 36926 -21111 37242 -21106
rect 36832 -21121 37242 -21111
rect 30945 -23767 31001 -23490
rect 30948 -24230 31004 -23989
rect 28308 -24912 28480 -24908
rect 28308 -24969 28407 -24912
rect 28463 -24969 28480 -24912
rect 28308 -25015 28480 -24969
rect 28308 -25072 28314 -25015
rect 28370 -25072 28480 -25015
rect 28308 -25084 28480 -25072
rect 28095 -26122 28222 -26099
rect 28095 -26197 28123 -26122
rect 28198 -26197 28222 -26122
rect 28095 -26277 28222 -26197
rect 28095 -26352 28119 -26277
rect 28195 -26352 28222 -26277
rect 28095 -26389 28222 -26352
rect 30997 -26553 31054 -26320
rect 26017 -26979 26027 -26878
rect 26103 -26880 26416 -26878
rect 26103 -26882 26333 -26880
rect 26103 -26979 26184 -26882
rect 26017 -26983 26184 -26979
rect 26260 -26981 26333 -26882
rect 26409 -26981 26416 -26880
rect 26260 -26983 26416 -26981
rect 26017 -29772 26416 -26983
rect 26017 -29775 26318 -29772
rect 26017 -29845 26023 -29775
rect 26089 -29776 26318 -29775
rect 26089 -29845 26175 -29776
rect 26017 -29846 26175 -29845
rect 26241 -29842 26318 -29776
rect 26384 -29842 26416 -29772
rect 26241 -29846 26416 -29842
rect 26017 -33395 26416 -29846
rect 26017 -33399 26311 -33395
rect 26017 -33469 26028 -33399
rect 26094 -33469 26162 -33399
rect 26228 -33465 26311 -33399
rect 26377 -33465 26416 -33395
rect 26228 -33469 26416 -33465
rect 26017 -35083 26416 -33469
rect 26017 -35085 26175 -35083
rect 26017 -35155 26033 -35085
rect 26099 -35153 26175 -35085
rect 26241 -35088 26416 -35083
rect 26241 -35153 26315 -35088
rect 26099 -35155 26315 -35153
rect 26017 -35158 26315 -35155
rect 26381 -35158 26416 -35088
rect 26017 -36500 26416 -35158
rect 36836 -28537 37235 -21121
rect 37522 -27501 37921 -20081
rect 37522 -27518 37932 -27501
rect 37522 -27521 37849 -27518
rect 37522 -27526 37700 -27521
rect 37522 -27621 37541 -27526
rect 37618 -27616 37700 -27526
rect 37777 -27613 37849 -27521
rect 37926 -27613 37932 -27518
rect 37777 -27616 37932 -27613
rect 37618 -27621 37932 -27616
rect 37522 -27694 37932 -27621
rect 37522 -27697 37846 -27694
rect 37522 -27702 37697 -27697
rect 37522 -27797 37538 -27702
rect 37615 -27792 37697 -27702
rect 37774 -27789 37846 -27697
rect 37923 -27789 37932 -27694
rect 37774 -27792 37932 -27789
rect 37615 -27797 37932 -27792
rect 37522 -27853 37932 -27797
rect 37522 -27856 37848 -27853
rect 37522 -27861 37699 -27856
rect 37522 -27956 37540 -27861
rect 37617 -27951 37699 -27861
rect 37776 -27948 37848 -27856
rect 37925 -27948 37932 -27853
rect 37776 -27951 37932 -27948
rect 37617 -27956 37932 -27951
rect 37522 -28011 37932 -27956
rect 37522 -28014 37847 -28011
rect 37522 -28019 37698 -28014
rect 37522 -28114 37539 -28019
rect 37616 -28109 37698 -28019
rect 37775 -28106 37847 -28014
rect 37924 -28106 37932 -28011
rect 37775 -28109 37932 -28106
rect 37616 -28114 37932 -28109
rect 37522 -28124 37932 -28114
rect 36836 -28554 37250 -28537
rect 36836 -28557 37167 -28554
rect 36836 -28562 37018 -28557
rect 36836 -28657 36859 -28562
rect 36936 -28652 37018 -28562
rect 37095 -28649 37167 -28557
rect 37244 -28649 37250 -28554
rect 37095 -28652 37250 -28649
rect 36936 -28657 37250 -28652
rect 36836 -28730 37250 -28657
rect 36836 -28733 37164 -28730
rect 36836 -28738 37015 -28733
rect 36836 -28833 36856 -28738
rect 36933 -28828 37015 -28738
rect 37092 -28825 37164 -28733
rect 37241 -28825 37250 -28730
rect 37092 -28828 37250 -28825
rect 36933 -28833 37250 -28828
rect 36836 -28889 37250 -28833
rect 36836 -28892 37166 -28889
rect 36836 -28897 37017 -28892
rect 36836 -28992 36858 -28897
rect 36935 -28987 37017 -28897
rect 37094 -28984 37166 -28892
rect 37243 -28984 37250 -28889
rect 37094 -28987 37250 -28984
rect 36935 -28992 37250 -28987
rect 36836 -29047 37250 -28992
rect 36836 -29050 37165 -29047
rect 36836 -29055 37016 -29050
rect 36836 -29150 36857 -29055
rect 36934 -29145 37016 -29055
rect 37093 -29142 37165 -29050
rect 37242 -29142 37250 -29047
rect 37093 -29145 37250 -29142
rect 36934 -29150 37250 -29145
rect 36836 -29160 37250 -29150
rect 26017 -36517 26431 -36500
rect 26017 -36520 26348 -36517
rect 26017 -36525 26199 -36520
rect 26017 -36620 26040 -36525
rect 26117 -36615 26199 -36525
rect 26276 -36612 26348 -36520
rect 26425 -36612 26431 -36517
rect 26276 -36615 26431 -36612
rect 26117 -36620 26431 -36615
rect 26017 -36693 26431 -36620
rect 26017 -36696 26345 -36693
rect 26017 -36701 26196 -36696
rect 26017 -36796 26037 -36701
rect 26114 -36791 26196 -36701
rect 26273 -36788 26345 -36696
rect 26422 -36788 26431 -36693
rect 26273 -36791 26431 -36788
rect 26114 -36796 26431 -36791
rect 26017 -36852 26431 -36796
rect 26017 -36855 26347 -36852
rect 26017 -36860 26198 -36855
rect 26017 -36955 26039 -36860
rect 26116 -36950 26198 -36860
rect 26275 -36947 26347 -36855
rect 26424 -36947 26431 -36852
rect 26275 -36950 26431 -36947
rect 26116 -36955 26431 -36950
rect 26017 -37010 26431 -36955
rect 26017 -37013 26346 -37010
rect 26017 -37018 26197 -37013
rect 26017 -37113 26038 -37018
rect 26115 -37108 26197 -37018
rect 26274 -37105 26346 -37013
rect 26423 -37105 26431 -37010
rect 26274 -37108 26431 -37105
rect 26115 -37113 26431 -37108
rect 26017 -37125 26431 -37113
rect 25331 -37550 25744 -37533
rect 25331 -37553 25661 -37550
rect 25331 -37558 25512 -37553
rect 25331 -37653 25353 -37558
rect 25430 -37648 25512 -37558
rect 25589 -37645 25661 -37553
rect 25738 -37645 25744 -37550
rect 25589 -37648 25744 -37645
rect 25430 -37653 25744 -37648
rect 25331 -37726 25744 -37653
rect 25331 -37729 25658 -37726
rect 25331 -37734 25509 -37729
rect 25331 -37829 25350 -37734
rect 25427 -37824 25509 -37734
rect 25586 -37821 25658 -37729
rect 25735 -37821 25744 -37726
rect 25586 -37824 25744 -37821
rect 25427 -37829 25744 -37824
rect 25331 -37885 25744 -37829
rect 25331 -37888 25660 -37885
rect 25331 -37893 25511 -37888
rect 25331 -37988 25352 -37893
rect 25429 -37983 25511 -37893
rect 25588 -37980 25660 -37888
rect 25737 -37980 25744 -37885
rect 25588 -37983 25744 -37980
rect 25429 -37988 25744 -37983
rect 25331 -38043 25744 -37988
rect 25331 -38046 25659 -38043
rect 25331 -38051 25510 -38046
rect 25331 -38146 25351 -38051
rect 25428 -38141 25510 -38051
rect 25587 -38138 25659 -38046
rect 25736 -38138 25744 -38043
rect 25587 -38141 25744 -38138
rect 25428 -38146 25744 -38141
rect 25331 -38158 25744 -38146
rect 25331 -38182 25730 -38158
rect 26017 -38182 26416 -37125
rect 36836 -38182 37235 -29160
rect 37522 -38182 37921 -28124
rect -56707 -38745 -56683 -38680
rect -56580 -38745 -56561 -38680
rect -56707 -38816 -56561 -38745
rect -56707 -38881 -56690 -38816
rect -56587 -38881 -56561 -38816
rect -56707 -38906 -56561 -38881
rect -57036 -39128 -57012 -39064
rect -56931 -39128 -56888 -39064
rect -57036 -39190 -56888 -39128
rect -57036 -39254 -57008 -39190
rect -56927 -39254 -56888 -39190
rect -57036 -39315 -56888 -39254
rect -57036 -39379 -57010 -39315
rect -56929 -39379 -56888 -39315
rect -57036 -39409 -56888 -39379
<< via2 >>
rect -65675 55729 -65598 55824
rect -65516 55734 -65439 55829
rect -65367 55737 -65290 55832
rect -65678 55553 -65601 55648
rect -65519 55558 -65442 55653
rect -65370 55561 -65293 55656
rect -65676 55394 -65599 55489
rect -65517 55399 -65440 55494
rect -65368 55402 -65291 55497
rect -65677 55236 -65600 55331
rect -65518 55241 -65441 55336
rect -65369 55244 -65292 55339
rect -66362 54691 -66285 54786
rect -66203 54696 -66126 54791
rect -66054 54699 -65977 54794
rect -66365 54515 -66288 54610
rect -66206 54520 -66129 54615
rect -66057 54523 -65980 54618
rect -66363 54356 -66286 54451
rect -66204 54361 -66127 54456
rect -66055 54364 -65978 54459
rect -66364 54198 -66287 54293
rect -66205 54203 -66128 54298
rect -66056 54206 -65979 54301
rect -70203 53504 -70126 53599
rect -70044 53509 -69967 53604
rect -69895 53512 -69818 53607
rect -70206 53328 -70129 53423
rect -70047 53333 -69970 53428
rect -69898 53336 -69821 53431
rect -70204 53169 -70127 53264
rect -70045 53174 -69968 53269
rect -69896 53177 -69819 53272
rect -70205 53011 -70128 53106
rect -70046 53016 -69969 53111
rect -69897 53019 -69820 53114
rect -70899 52456 -70822 52551
rect -70740 52461 -70663 52556
rect -70591 52464 -70514 52559
rect -70902 52280 -70825 52375
rect -70743 52285 -70666 52380
rect -70594 52288 -70517 52383
rect -70900 52121 -70823 52216
rect -70741 52126 -70664 52221
rect -70592 52129 -70515 52224
rect -70901 51963 -70824 52058
rect -70742 51968 -70665 52063
rect -70593 51971 -70516 52066
rect -70203 45129 -70126 45224
rect -70044 45134 -69967 45229
rect -69895 45137 -69818 45232
rect -70206 44953 -70129 45048
rect -70047 44958 -69970 45053
rect -69898 44961 -69821 45056
rect -70204 44794 -70127 44889
rect -70045 44799 -69968 44894
rect -69896 44802 -69819 44897
rect -70205 44636 -70128 44731
rect -70046 44641 -69969 44736
rect -69897 44644 -69820 44739
rect -70895 44086 -70818 44181
rect -70736 44091 -70659 44186
rect -70587 44094 -70510 44189
rect -70898 43910 -70821 44005
rect -70739 43915 -70662 44010
rect -70590 43918 -70513 44013
rect -70896 43751 -70819 43846
rect -70737 43756 -70660 43851
rect -70588 43759 -70511 43854
rect -70897 43593 -70820 43688
rect -70738 43598 -70661 43693
rect -70589 43601 -70512 43696
rect -69407 41042 -69346 41107
rect -69513 39225 -69434 39299
rect -70203 36912 -70126 37007
rect -70044 36917 -69967 37012
rect -69895 36920 -69818 37015
rect -70206 36736 -70129 36831
rect -70047 36741 -69970 36836
rect -69898 36744 -69821 36839
rect -70204 36577 -70127 36672
rect -70045 36582 -69968 36677
rect -69896 36585 -69819 36680
rect -70205 36419 -70128 36514
rect -70046 36424 -69969 36519
rect -69897 36427 -69820 36522
rect -70891 35661 -70814 35756
rect -70732 35666 -70655 35761
rect -70583 35669 -70506 35764
rect -70894 35485 -70817 35580
rect -70735 35490 -70658 35585
rect -70586 35493 -70509 35588
rect -70892 35326 -70815 35421
rect -70733 35331 -70656 35426
rect -70584 35334 -70507 35429
rect -70893 35168 -70816 35263
rect -70734 35173 -70657 35268
rect -70585 35176 -70508 35271
rect -70207 28355 -70130 28450
rect -70048 28360 -69971 28455
rect -69899 28363 -69822 28458
rect -70210 28179 -70133 28274
rect -70051 28184 -69974 28279
rect -69902 28187 -69825 28282
rect -70208 28020 -70131 28115
rect -70049 28025 -69972 28120
rect -69900 28028 -69823 28123
rect -70209 27862 -70132 27957
rect -70050 27867 -69973 27962
rect -69901 27870 -69824 27965
rect -70891 27245 -70814 27340
rect -70732 27250 -70655 27345
rect -70583 27253 -70506 27348
rect -70894 27069 -70817 27164
rect -70735 27074 -70658 27169
rect -70586 27077 -70509 27172
rect -70892 26910 -70815 27005
rect -70733 26915 -70656 27010
rect -70584 26918 -70507 27013
rect -70893 26752 -70816 26847
rect -70734 26757 -70657 26852
rect -70585 26760 -70508 26855
rect -70203 19297 -70126 19392
rect -70044 19302 -69967 19397
rect -69895 19305 -69818 19400
rect -70206 19121 -70129 19216
rect -70047 19126 -69970 19221
rect -69898 19129 -69821 19224
rect -70204 18962 -70127 19057
rect -70045 18967 -69968 19062
rect -69896 18970 -69819 19065
rect -70205 18804 -70128 18899
rect -70046 18809 -69969 18904
rect -69897 18812 -69820 18907
rect -70895 18216 -70818 18311
rect -70736 18221 -70659 18316
rect -70587 18224 -70510 18319
rect -70898 18040 -70821 18135
rect -70739 18045 -70662 18140
rect -70590 18048 -70513 18143
rect -70896 17881 -70819 17976
rect -70737 17886 -70660 17981
rect -70588 17889 -70511 17984
rect -70897 17723 -70820 17818
rect -70738 17728 -70661 17823
rect -70589 17731 -70512 17826
rect -71904 11197 -71787 11310
rect -71610 11194 -71493 11307
rect -71907 10899 -71790 11012
rect -71617 10899 -71500 11012
rect -70203 7277 -70126 7372
rect -70044 7282 -69967 7377
rect -69895 7285 -69818 7380
rect -70206 7101 -70129 7196
rect -70047 7106 -69970 7201
rect -69898 7109 -69821 7204
rect -70204 6942 -70127 7037
rect -70045 6947 -69968 7042
rect -69896 6950 -69819 7045
rect -70205 6784 -70128 6879
rect -70046 6789 -69969 6884
rect -69897 6792 -69820 6887
rect -70899 6047 -70822 6142
rect -70740 6052 -70663 6147
rect -70591 6055 -70514 6150
rect -70902 5871 -70825 5966
rect -70743 5876 -70666 5971
rect -70594 5879 -70517 5974
rect -70900 5712 -70823 5807
rect -70741 5717 -70664 5812
rect -70592 5720 -70515 5815
rect -70901 5554 -70824 5649
rect -70742 5559 -70665 5654
rect -70593 5562 -70516 5657
rect -70203 -2564 -70126 -2469
rect -70044 -2559 -69967 -2464
rect -69895 -2556 -69818 -2461
rect -70206 -2740 -70129 -2645
rect -70047 -2735 -69970 -2640
rect -69898 -2732 -69821 -2637
rect -70204 -2899 -70127 -2804
rect -70045 -2894 -69968 -2799
rect -69896 -2891 -69819 -2796
rect -70205 -3057 -70128 -2962
rect -70046 -3052 -69969 -2957
rect -69897 -3049 -69820 -2954
rect -70891 -3645 -70814 -3550
rect -70732 -3640 -70655 -3545
rect -70583 -3637 -70506 -3542
rect -70894 -3821 -70817 -3726
rect -70735 -3816 -70658 -3721
rect -70586 -3813 -70509 -3718
rect -70892 -3980 -70815 -3885
rect -70733 -3975 -70656 -3880
rect -70584 -3972 -70507 -3877
rect -70893 -4138 -70816 -4043
rect -70734 -4133 -70657 -4038
rect -70585 -4130 -70508 -4035
rect -70199 -11489 -70122 -11394
rect -70040 -11484 -69963 -11389
rect -69891 -11481 -69814 -11386
rect -70202 -11665 -70125 -11570
rect -70043 -11660 -69966 -11565
rect -69894 -11657 -69817 -11562
rect -70200 -11824 -70123 -11729
rect -70041 -11819 -69964 -11724
rect -69892 -11816 -69815 -11721
rect -70201 -11982 -70124 -11887
rect -70042 -11977 -69965 -11882
rect -69893 -11974 -69816 -11879
rect -70887 -12533 -70810 -12438
rect -70728 -12528 -70651 -12433
rect -70579 -12525 -70502 -12430
rect -70890 -12709 -70813 -12614
rect -70731 -12704 -70654 -12609
rect -70582 -12701 -70505 -12606
rect -70888 -12868 -70811 -12773
rect -70729 -12863 -70652 -12768
rect -70580 -12860 -70503 -12765
rect -70889 -13026 -70812 -12931
rect -70730 -13021 -70653 -12926
rect -70581 -13018 -70504 -12923
rect -70203 -19578 -70126 -19483
rect -70044 -19573 -69967 -19478
rect -69895 -19570 -69818 -19475
rect -70206 -19754 -70129 -19659
rect -70047 -19749 -69970 -19654
rect -69898 -19746 -69821 -19651
rect -70204 -19913 -70127 -19818
rect -70045 -19908 -69968 -19813
rect -69896 -19905 -69819 -19810
rect -70205 -20071 -70128 -19976
rect -70046 -20066 -69969 -19971
rect -69897 -20063 -69820 -19968
rect -70895 -20618 -70818 -20523
rect -70736 -20613 -70659 -20518
rect -70587 -20610 -70510 -20515
rect -70898 -20794 -70821 -20699
rect -70739 -20789 -70662 -20694
rect -70590 -20786 -70513 -20691
rect -70896 -20953 -70819 -20858
rect -70737 -20948 -70660 -20853
rect -70588 -20945 -70511 -20850
rect -70897 -21111 -70820 -21016
rect -70738 -21106 -70661 -21011
rect -70589 -21103 -70512 -21008
rect -68318 31130 -68237 31187
rect -68348 22714 -68263 22803
rect -68333 13646 -68258 13716
rect -68328 1064 -68246 1157
rect -68380 -7936 -68289 -7856
rect -68379 -8111 -68288 -8031
rect -68375 -16749 -68295 -16634
rect -68377 -17006 -68297 -16891
rect -66855 -23497 -66759 -23417
rect -70203 -27626 -70126 -27531
rect -70044 -27621 -69967 -27526
rect -69895 -27618 -69818 -27523
rect -70206 -27802 -70129 -27707
rect -70047 -27797 -69970 -27702
rect -69898 -27794 -69821 -27699
rect -70204 -27961 -70127 -27866
rect -70045 -27956 -69968 -27861
rect -69896 -27953 -69819 -27858
rect -70205 -28119 -70128 -28024
rect -70046 -28114 -69969 -28019
rect -69897 -28111 -69820 -28016
rect -70887 -28657 -70810 -28562
rect -70728 -28652 -70651 -28557
rect -70579 -28649 -70502 -28554
rect -70890 -28833 -70813 -28738
rect -70731 -28828 -70654 -28733
rect -70582 -28825 -70505 -28730
rect -70888 -28992 -70811 -28897
rect -70729 -28987 -70652 -28892
rect -70580 -28984 -70503 -28889
rect -70889 -29150 -70812 -29055
rect -70730 -29145 -70653 -29050
rect -70581 -29142 -70504 -29047
rect -55274 55728 -55197 55823
rect -55115 55733 -55038 55828
rect -54966 55736 -54889 55831
rect -55277 55552 -55200 55647
rect -55118 55557 -55041 55652
rect -54969 55560 -54892 55655
rect -55275 55393 -55198 55488
rect -55116 55398 -55039 55493
rect -54967 55401 -54890 55496
rect -55276 55235 -55199 55330
rect -55117 55240 -55040 55335
rect -54968 55243 -54891 55338
rect -55922 54693 -55845 54788
rect -55763 54698 -55686 54793
rect -55614 54701 -55537 54796
rect -55925 54517 -55848 54612
rect -55766 54522 -55689 54617
rect -55617 54525 -55540 54620
rect -55923 54358 -55846 54453
rect -55764 54363 -55687 54458
rect -55615 54366 -55538 54461
rect -55924 54200 -55847 54295
rect -55765 54205 -55688 54300
rect -55616 54208 -55539 54303
rect -63590 40847 -63479 40954
rect -63103 38910 -62992 39017
rect -56569 36925 -56492 37020
rect -56572 36749 -56495 36844
rect -56570 36590 -56493 36685
rect -56571 36432 -56494 36527
rect -56777 35668 -56700 35763
rect -56780 35492 -56703 35587
rect -56778 35333 -56701 35428
rect -56779 35175 -56702 35270
rect -63356 33209 -63265 33288
rect -63360 33057 -63269 33136
rect -63769 31271 -63678 31350
rect -63773 31119 -63682 31198
rect -56557 19314 -56480 19409
rect -56560 19138 -56483 19233
rect -56558 18979 -56481 19074
rect -56559 18821 -56482 18916
rect -56752 18231 -56675 18326
rect -56755 18055 -56678 18150
rect -56753 17896 -56676 17991
rect -56754 17738 -56677 17833
rect -63321 15647 -63265 15703
rect -63325 15536 -63269 15592
rect -63611 13707 -63555 13763
rect -63615 13596 -63559 13652
rect -56569 7301 -56492 7396
rect -56572 7125 -56495 7220
rect -56570 6966 -56493 7061
rect -56571 6808 -56494 6903
rect -56773 6062 -56696 6157
rect -56776 5886 -56699 5981
rect -56774 5727 -56697 5822
rect -56775 5569 -56698 5664
rect -63329 3324 -63273 3380
rect -63333 3213 -63277 3269
rect -63742 1354 -63686 1410
rect -63746 1243 -63690 1299
rect -56591 -2550 -56514 -2455
rect -56594 -2726 -56517 -2631
rect -56592 -2885 -56515 -2790
rect -56593 -3043 -56516 -2948
rect -56794 -3621 -56717 -3526
rect -56797 -3797 -56720 -3702
rect -56795 -3956 -56718 -3861
rect -56796 -4114 -56719 -4019
rect -63338 -6178 -63282 -6122
rect -63342 -6289 -63286 -6233
rect -64331 -8142 -64275 -8086
rect -64335 -8253 -64279 -8197
rect -56585 -11476 -56508 -11381
rect -56588 -11652 -56511 -11557
rect -56586 -11811 -56509 -11716
rect -56587 -11969 -56510 -11874
rect -56792 -12516 -56715 -12421
rect -56795 -12692 -56718 -12597
rect -56793 -12851 -56716 -12756
rect -56794 -13009 -56717 -12914
rect -63334 -14965 -63278 -14909
rect -63338 -15076 -63282 -15020
rect -63656 -16935 -63600 -16879
rect -63660 -17046 -63604 -16990
rect -56627 -19571 -56550 -19476
rect -56630 -19747 -56553 -19652
rect -56628 -19906 -56551 -19811
rect -56629 -20064 -56552 -19969
rect -56831 -20608 -56754 -20513
rect -56834 -20784 -56757 -20689
rect -56832 -20943 -56755 -20848
rect -56833 -21101 -56756 -21006
rect -63383 -23068 -63327 -23012
rect -63387 -23179 -63331 -23123
rect -63726 -25008 -63670 -24952
rect -63730 -25119 -63674 -25063
rect -65675 -36624 -65598 -36529
rect -65516 -36619 -65439 -36524
rect -65367 -36616 -65290 -36521
rect -65678 -36800 -65601 -36705
rect -65519 -36795 -65442 -36700
rect -65370 -36792 -65293 -36697
rect -65676 -36959 -65599 -36864
rect -65517 -36954 -65440 -36859
rect -65368 -36951 -65291 -36856
rect -65677 -37117 -65600 -37022
rect -65518 -37112 -65441 -37017
rect -65369 -37109 -65292 -37014
rect -66371 -37656 -66294 -37561
rect -66212 -37651 -66135 -37556
rect -66063 -37648 -65986 -37553
rect -66374 -37832 -66297 -37737
rect -66215 -37827 -66138 -37732
rect -66066 -37824 -65989 -37729
rect -66372 -37991 -66295 -37896
rect -66213 -37986 -66136 -37891
rect -66064 -37983 -65987 -37888
rect -66373 -38149 -66296 -38054
rect -66214 -38144 -66137 -38049
rect -66065 -38141 -65988 -38046
rect -56365 -32969 -56276 -32893
rect -56370 -33160 -56281 -33084
rect -44920 55731 -44843 55826
rect -44761 55736 -44684 55831
rect -44612 55739 -44535 55834
rect -44923 55555 -44846 55650
rect -44764 55560 -44687 55655
rect -44615 55563 -44538 55658
rect -44921 55396 -44844 55491
rect -44762 55401 -44685 55496
rect -44613 55404 -44536 55499
rect -44922 55238 -44845 55333
rect -44763 55243 -44686 55338
rect -44614 55246 -44537 55341
rect -45742 54706 -45665 54801
rect -45583 54711 -45506 54806
rect -45434 54714 -45357 54809
rect -45745 54530 -45668 54625
rect -45586 54535 -45509 54630
rect -45437 54538 -45360 54633
rect -45743 54371 -45666 54466
rect -45584 54376 -45507 54471
rect -45435 54379 -45358 54474
rect -45744 54213 -45667 54308
rect -45585 54218 -45508 54313
rect -45436 54221 -45359 54316
rect -46395 53507 -46318 53602
rect -46398 53331 -46321 53426
rect -46396 53172 -46319 53267
rect -46397 53014 -46320 53109
rect -46599 52477 -46522 52572
rect -46600 52274 -46523 52369
rect -46601 52072 -46524 52167
rect -53252 50012 -53161 50091
rect -53256 49860 -53165 49939
rect -46389 45133 -46312 45228
rect -46392 44957 -46315 45052
rect -46390 44798 -46313 44893
rect -46391 44640 -46314 44735
rect -46592 44096 -46515 44191
rect -46595 43920 -46518 44015
rect -46593 43761 -46516 43856
rect -46594 43603 -46517 43698
rect -53175 41678 -53084 41757
rect -53179 41526 -53088 41605
rect -46396 36925 -46319 37020
rect -46399 36749 -46322 36844
rect -46397 36590 -46320 36685
rect -46398 36432 -46321 36527
rect -46601 35668 -46524 35763
rect -46604 35492 -46527 35587
rect -46602 35333 -46525 35428
rect -46603 35175 -46526 35270
rect -53184 33214 -53093 33293
rect -53188 33062 -53097 33141
rect -53483 31271 -53392 31350
rect -53487 31119 -53396 31198
rect -46406 19314 -46329 19409
rect -46409 19138 -46332 19233
rect -46407 18979 -46330 19074
rect -46408 18821 -46331 18916
rect -46605 18227 -46528 18322
rect -46608 18051 -46531 18146
rect -46606 17892 -46529 17987
rect -46607 17734 -46530 17829
rect -53166 15877 -53110 15933
rect -53170 15766 -53114 15822
rect -53461 13979 -53405 14035
rect -53465 13868 -53409 13924
rect -46419 7301 -46342 7396
rect -46422 7125 -46345 7220
rect -46420 6966 -46343 7061
rect -46421 6808 -46344 6903
rect -46623 6066 -46546 6161
rect -46626 5890 -46549 5985
rect -46624 5731 -46547 5826
rect -46625 5573 -46548 5668
rect -53194 2993 -53138 3049
rect -53198 2882 -53142 2938
rect -53627 1038 -53571 1094
rect -53631 927 -53575 983
rect -53009 984 -52949 1062
rect -52878 995 -52818 1073
rect -46430 -19566 -46353 -19471
rect -46433 -19742 -46356 -19647
rect -46431 -19901 -46354 -19806
rect -46432 -20059 -46355 -19964
rect -46636 -20604 -46559 -20509
rect -46639 -20780 -46562 -20685
rect -46637 -20939 -46560 -20844
rect -46638 -21097 -46561 -21002
rect -53191 -23036 -53135 -22980
rect -53195 -23147 -53139 -23091
rect -53526 -24971 -53467 -24909
rect -53543 -25109 -53484 -25047
rect -46396 -27608 -46319 -27513
rect -46399 -27784 -46322 -27689
rect -46397 -27943 -46320 -27848
rect -46398 -28101 -46321 -28006
rect -46607 -28650 -46530 -28555
rect -46610 -28826 -46533 -28731
rect -46608 -28985 -46531 -28890
rect -46609 -29143 -46532 -29048
rect -53633 -33086 -53555 -33085
rect -53633 -33162 -53632 -33086
rect -53632 -33162 -53556 -33086
rect -53556 -33162 -53555 -33086
rect -53633 -33163 -53555 -33162
rect -53468 -33163 -53390 -33085
rect -55277 -36613 -55200 -36518
rect -55118 -36608 -55041 -36513
rect -54969 -36605 -54892 -36510
rect -55280 -36789 -55203 -36694
rect -55121 -36784 -55044 -36689
rect -54972 -36781 -54895 -36686
rect -55278 -36948 -55201 -36853
rect -55119 -36943 -55042 -36848
rect -54970 -36940 -54893 -36845
rect -55279 -37106 -55202 -37011
rect -55120 -37101 -55043 -37006
rect -54971 -37098 -54894 -37003
rect -55919 -37659 -55842 -37564
rect -55760 -37654 -55683 -37559
rect -55611 -37651 -55534 -37556
rect -55922 -37835 -55845 -37740
rect -55763 -37830 -55686 -37735
rect -55614 -37827 -55537 -37732
rect -55920 -37994 -55843 -37899
rect -55761 -37989 -55684 -37894
rect -55612 -37986 -55535 -37891
rect -55921 -38152 -55844 -38057
rect -55762 -38147 -55685 -38052
rect -55613 -38144 -55536 -38049
rect -34684 55728 -34607 55823
rect -34525 55733 -34448 55828
rect -34376 55736 -34299 55831
rect -34687 55552 -34610 55647
rect -34528 55557 -34451 55652
rect -34379 55560 -34302 55655
rect -34685 55393 -34608 55488
rect -34526 55398 -34449 55493
rect -34377 55401 -34300 55496
rect -34686 55235 -34609 55330
rect -34527 55240 -34450 55335
rect -34378 55243 -34301 55338
rect -35374 54693 -35297 54788
rect -35215 54698 -35138 54793
rect -35066 54701 -34989 54796
rect -35377 54517 -35300 54612
rect -35218 54522 -35141 54617
rect -35069 54525 -34992 54620
rect -35375 54358 -35298 54453
rect -35216 54363 -35139 54458
rect -35067 54366 -34990 54461
rect -35376 54200 -35299 54295
rect -35217 54205 -35140 54300
rect -35068 54208 -34991 54303
rect -36016 53520 -35939 53615
rect -36019 53344 -35942 53439
rect -36017 53185 -35940 53280
rect -36018 53027 -35941 53122
rect -36236 52468 -36159 52563
rect -36239 52292 -36162 52387
rect -36237 52133 -36160 52228
rect -36238 51975 -36161 52070
rect -42873 49905 -42782 49984
rect -42877 49753 -42786 49832
rect -36083 45136 -36006 45231
rect -36086 44960 -36009 45055
rect -36084 44801 -36007 44896
rect -36085 44643 -36008 44738
rect -36289 44093 -36212 44188
rect -36292 43917 -36215 44012
rect -36290 43758 -36213 43853
rect -36291 43600 -36214 43695
rect -42854 41708 -42763 41787
rect -42858 41556 -42767 41635
rect -36023 36925 -35946 37020
rect -36026 36749 -35949 36844
rect -36024 36590 -35947 36685
rect -36025 36432 -35948 36527
rect -36221 35671 -36144 35766
rect -36224 35495 -36147 35590
rect -36222 35336 -36145 35431
rect -36223 35178 -36146 35273
rect -42790 33185 -42699 33264
rect -42794 33033 -42703 33112
rect -43109 31240 -43018 31319
rect -43113 31088 -43022 31167
rect -36223 28364 -36146 28459
rect -36226 28188 -36149 28283
rect -36224 28029 -36147 28124
rect -36225 27871 -36148 27966
rect -36430 27249 -36353 27344
rect -36433 27073 -36356 27168
rect -36431 26914 -36354 27009
rect -36432 26756 -36355 26851
rect -43004 24774 -42913 24853
rect -43008 24622 -42917 24701
rect -43303 22834 -43212 22913
rect -43307 22682 -43216 22761
rect -42963 15566 -42907 15622
rect -42967 15455 -42911 15511
rect -36194 19321 -36117 19416
rect -36197 19145 -36120 19240
rect -36195 18986 -36118 19081
rect -36196 18828 -36119 18923
rect -36400 18231 -36323 18326
rect -36403 18055 -36326 18150
rect -36401 17896 -36324 17991
rect -36402 17738 -36325 17833
rect -43268 13608 -43212 13664
rect -42693 13635 -42628 13718
rect -42561 13639 -42496 13722
rect -43272 13497 -43216 13553
rect -36009 7298 -35932 7393
rect -36012 7122 -35935 7217
rect -36010 6963 -35933 7058
rect -36011 6805 -35934 6900
rect -36217 6059 -36140 6154
rect -36220 5883 -36143 5978
rect -36218 5724 -36141 5819
rect -36219 5566 -36142 5661
rect -42778 2760 -42722 2816
rect -42782 2649 -42726 2705
rect -43134 851 -43078 907
rect -43138 740 -43082 796
rect -36040 -2550 -35963 -2455
rect -36043 -2726 -35966 -2631
rect -36041 -2885 -35964 -2790
rect -36042 -3043 -35965 -2948
rect -36247 -3624 -36170 -3529
rect -36250 -3800 -36173 -3705
rect -36248 -3959 -36171 -3864
rect -36249 -4117 -36172 -4022
rect -42799 -6203 -42743 -6147
rect -42803 -6314 -42747 -6258
rect -43097 -8116 -43015 -8034
rect -43097 -8281 -43015 -8199
rect -42673 -8223 -42605 -8137
rect -42509 -8219 -42441 -8133
rect -36198 -11472 -36121 -11377
rect -36201 -11648 -36124 -11553
rect -36199 -11807 -36122 -11712
rect -36200 -11965 -36123 -11870
rect -36403 -12517 -36326 -12422
rect -36406 -12693 -36329 -12598
rect -36404 -12852 -36327 -12757
rect -36405 -13010 -36328 -12915
rect -42972 -15155 -42916 -15099
rect -42976 -15266 -42920 -15210
rect -43324 -17028 -43268 -16972
rect -43328 -17139 -43272 -17083
rect -36053 -19561 -35976 -19466
rect -36056 -19737 -35979 -19642
rect -36054 -19896 -35977 -19801
rect -36055 -20054 -35978 -19959
rect -36260 -20608 -36183 -20513
rect -36263 -20784 -36186 -20689
rect -36261 -20943 -36184 -20848
rect -36262 -21101 -36185 -21006
rect -42800 -23045 -42744 -22989
rect -42804 -23156 -42748 -23100
rect -43341 -25117 -43267 -25050
rect -43186 -25104 -43112 -25037
rect -42676 -25098 -42616 -25027
rect -42538 -25094 -42478 -25023
rect -44920 -36620 -44843 -36525
rect -44761 -36615 -44684 -36520
rect -44612 -36612 -44535 -36517
rect -44923 -36796 -44846 -36701
rect -44764 -36791 -44687 -36696
rect -44615 -36788 -44538 -36693
rect -44921 -36955 -44844 -36860
rect -44762 -36950 -44685 -36855
rect -44613 -36947 -44536 -36852
rect -44922 -37113 -44845 -37018
rect -44763 -37108 -44686 -37013
rect -44614 -37105 -44537 -37010
rect -45742 -37659 -45665 -37564
rect -45583 -37654 -45506 -37559
rect -45434 -37651 -45357 -37556
rect -45745 -37835 -45668 -37740
rect -45586 -37830 -45509 -37735
rect -45437 -37827 -45360 -37732
rect -45743 -37994 -45666 -37899
rect -45584 -37989 -45507 -37894
rect -45435 -37986 -45358 -37891
rect -45744 -38152 -45667 -38057
rect -45585 -38147 -45508 -38052
rect -45436 -38144 -45359 -38049
rect -36007 -27604 -35930 -27509
rect -36010 -27780 -35933 -27685
rect -36008 -27939 -35931 -27844
rect -36009 -28097 -35932 -28002
rect -36214 -28646 -36137 -28551
rect -36217 -28822 -36140 -28727
rect -36215 -28981 -36138 -28886
rect -36216 -29139 -36139 -29044
rect -43133 -33147 -43077 -33088
rect -43020 -33144 -42964 -33085
rect -23375 55728 -23298 55823
rect -23216 55733 -23139 55828
rect -23067 55736 -22990 55831
rect -23378 55552 -23301 55647
rect -23219 55557 -23142 55652
rect -23070 55560 -22993 55655
rect -23376 55393 -23299 55488
rect -23217 55398 -23140 55493
rect -23068 55401 -22991 55496
rect -23377 55235 -23300 55330
rect -23218 55240 -23141 55335
rect -23069 55243 -22992 55338
rect -24170 54689 -24093 54784
rect -24011 54694 -23934 54789
rect -23862 54697 -23785 54792
rect -24173 54513 -24096 54608
rect -24014 54518 -23937 54613
rect -23865 54521 -23788 54616
rect -24171 54354 -24094 54449
rect -24012 54359 -23935 54454
rect -23863 54362 -23786 54457
rect -24172 54196 -24095 54291
rect -24013 54201 -23936 54296
rect -23864 54204 -23787 54299
rect -32478 49929 -32359 50028
rect -32484 49707 -32365 49806
rect -32467 41675 -32362 41759
rect -32472 41484 -32367 41568
rect -24963 36925 -24886 37020
rect -24966 36749 -24889 36844
rect -24964 36590 -24887 36685
rect -24965 36432 -24888 36527
rect -25161 35665 -25084 35760
rect -25164 35489 -25087 35584
rect -25162 35330 -25085 35425
rect -25163 35172 -25086 35267
rect -31731 33029 -31640 33108
rect -31735 32877 -31644 32956
rect -32035 31055 -31944 31134
rect -32039 30903 -31948 30982
rect -11204 53507 -11127 53602
rect -11207 53331 -11130 53426
rect -11205 53172 -11128 53267
rect -11206 53014 -11129 53109
rect -11417 52461 -11340 52556
rect -11420 52285 -11343 52380
rect -11418 52126 -11341 52221
rect -11419 51968 -11342 52063
rect -17978 49888 -17887 49967
rect -17982 49736 -17891 49815
rect -7126 55729 -7049 55824
rect -6967 55734 -6890 55829
rect -6818 55737 -6741 55832
rect -7129 55553 -7052 55648
rect -6970 55558 -6893 55653
rect -6821 55561 -6744 55656
rect -7127 55394 -7050 55489
rect -6968 55399 -6891 55494
rect -6819 55402 -6742 55497
rect -7128 55236 -7051 55331
rect -6969 55241 -6892 55336
rect -6820 55244 -6743 55339
rect -7899 54693 -7822 54788
rect -7740 54698 -7663 54793
rect -7591 54701 -7514 54796
rect -7902 54517 -7825 54612
rect -7743 54522 -7666 54617
rect -7594 54525 -7517 54620
rect -7900 54358 -7823 54453
rect -7741 54363 -7664 54458
rect -7592 54366 -7515 54461
rect -7901 54200 -7824 54295
rect -7742 54205 -7665 54300
rect -7593 54208 -7516 54303
rect -11035 45136 -10958 45231
rect -11038 44960 -10961 45055
rect -11036 44801 -10959 44896
rect -11037 44643 -10960 44738
rect -11241 44093 -11164 44188
rect -11244 43917 -11167 44012
rect -25823 19318 -25746 19413
rect -25826 19142 -25749 19237
rect -25824 18983 -25747 19078
rect -25825 18825 -25748 18920
rect -26029 18231 -25952 18326
rect -26032 18055 -25955 18150
rect -26030 17896 -25953 17991
rect -26031 17738 -25954 17833
rect -32593 15704 -32537 15760
rect -32597 15593 -32541 15649
rect -24175 14008 -24069 14094
rect -23950 14010 -23844 14096
rect -32931 13796 -32875 13852
rect -32935 13685 -32879 13741
rect -27090 7294 -27013 7389
rect -27093 7118 -27016 7213
rect -27091 6959 -27014 7054
rect -27092 6801 -27015 6896
rect -27916 6066 -27839 6161
rect -27919 5890 -27842 5985
rect -27917 5731 -27840 5826
rect -27918 5573 -27841 5668
rect -32474 2762 -32418 2818
rect -32478 2651 -32422 2707
rect -32833 911 -32777 967
rect -32837 800 -32781 856
rect -25102 -11472 -25025 -11377
rect -25105 -11648 -25028 -11553
rect -25103 -11807 -25026 -11712
rect -25104 -11965 -25027 -11870
rect -25303 -12517 -25226 -12422
rect -25306 -12693 -25229 -12598
rect -25304 -12852 -25227 -12757
rect -25305 -13010 -25228 -12915
rect -31855 -15052 -31799 -14996
rect -31859 -15163 -31803 -15107
rect -32183 -16887 -32114 -16809
rect -32183 -17069 -32114 -16991
rect -34681 -36616 -34604 -36521
rect -34522 -36611 -34445 -36516
rect -34373 -36608 -34296 -36513
rect -34684 -36792 -34607 -36697
rect -34525 -36787 -34448 -36692
rect -34376 -36784 -34299 -36689
rect -34682 -36951 -34605 -36856
rect -34523 -36946 -34446 -36851
rect -34374 -36943 -34297 -36848
rect -34683 -37109 -34606 -37014
rect -34524 -37104 -34447 -37009
rect -34375 -37101 -34298 -37006
rect -35371 -37663 -35294 -37568
rect -35212 -37658 -35135 -37563
rect -35063 -37655 -34986 -37560
rect -35374 -37839 -35297 -37744
rect -35215 -37834 -35138 -37739
rect -35066 -37831 -34989 -37736
rect -35372 -37998 -35295 -37903
rect -35213 -37993 -35136 -37898
rect -35064 -37990 -34987 -37895
rect -35373 -38156 -35296 -38061
rect -35214 -38151 -35137 -38056
rect -35065 -38148 -34988 -38053
rect -11242 43758 -11165 43853
rect -11243 43600 -11166 43695
rect -17805 41576 -17714 41655
rect -17809 41424 -17718 41503
rect -19287 33156 -19196 33244
rect -19284 32949 -19193 33037
rect -21211 19320 -21134 19415
rect -11137 36925 -11060 37020
rect -11140 36749 -11063 36844
rect -11138 36590 -11061 36685
rect -11139 36432 -11062 36527
rect -11338 35675 -11261 35770
rect -11341 35499 -11264 35594
rect -11339 35340 -11262 35435
rect -11340 35182 -11263 35277
rect -17916 33071 -17825 33150
rect -17920 32919 -17829 32998
rect -18207 31095 -18116 31174
rect -18211 30943 -18120 31022
rect -11847 28361 -11770 28456
rect -11850 28185 -11773 28280
rect -11848 28026 -11771 28121
rect -11849 27868 -11772 27963
rect -12047 27263 -11970 27358
rect -12050 27087 -11973 27182
rect -12048 26928 -11971 27023
rect -12049 26770 -11972 26865
rect -18615 24812 -18524 24891
rect -18619 24660 -18528 24739
rect -19029 22886 -18938 22965
rect -19033 22734 -18942 22813
rect -21214 19144 -21137 19239
rect -21212 18985 -21135 19080
rect -21213 18827 -21136 18922
rect -20728 18251 -20651 18346
rect -20731 18075 -20654 18170
rect -20729 17916 -20652 18011
rect -20730 17758 -20653 17853
rect -8395 24801 -8259 24913
rect -8407 24531 -8271 24643
rect -20225 15320 -20135 15406
rect -20229 15115 -20139 15201
rect -9885 15037 -9818 15113
rect -9726 15038 -9659 15114
rect -20237 13625 -20151 13726
rect -20022 13628 -19936 13729
rect -8891 13624 -8801 13727
rect -8685 13627 -8595 13730
rect -18798 9756 -18733 9831
rect -18798 8635 -18733 8703
rect -18798 8504 -18733 8569
rect -12562 -2550 -12485 -2455
rect -12565 -2726 -12488 -2631
rect -12563 -2885 -12486 -2790
rect -12564 -3043 -12487 -2948
rect -12768 -3628 -12691 -3533
rect -12771 -3804 -12694 -3709
rect -12769 -3963 -12692 -3868
rect -12770 -4121 -12693 -4026
rect -19334 -6239 -19278 -6183
rect -19338 -6350 -19282 -6294
rect -19850 -8314 -19768 -8232
rect -19685 -8314 -19603 -8232
rect -11090 -11472 -11013 -11377
rect -11093 -11648 -11016 -11553
rect -11091 -11807 -11014 -11712
rect -11092 -11965 -11015 -11870
rect -11291 -12517 -11214 -12422
rect -11294 -12693 -11217 -12598
rect -11292 -12852 -11215 -12757
rect -11293 -13010 -11216 -12915
rect -17851 -15128 -17795 -15072
rect -17855 -15239 -17799 -15183
rect -18441 -17051 -18359 -16969
rect -18276 -17051 -18194 -16969
rect -11142 -19566 -11065 -19471
rect -11145 -19742 -11068 -19647
rect -11143 -19901 -11066 -19806
rect -11144 -20059 -11067 -19964
rect -11345 -20608 -11268 -20513
rect -11348 -20784 -11271 -20689
rect -11346 -20943 -11269 -20848
rect -11347 -21101 -11270 -21006
rect -17892 -23057 -17836 -23001
rect -17896 -23168 -17840 -23112
rect -18255 -24936 -18173 -24854
rect -18255 -25101 -18173 -25019
rect -11180 -27608 -11103 -27513
rect -11183 -27784 -11106 -27689
rect -11181 -27943 -11104 -27848
rect -11182 -28101 -11105 -28006
rect -11386 -28646 -11309 -28551
rect -23381 -36620 -23304 -36525
rect -23222 -36615 -23145 -36520
rect -23073 -36612 -22996 -36517
rect -23384 -36796 -23307 -36701
rect -23225 -36791 -23148 -36696
rect -23076 -36788 -22999 -36693
rect -11389 -28822 -11312 -28727
rect -11387 -28981 -11310 -28886
rect -11388 -29139 -11311 -29044
rect -18438 -33149 -18377 -33081
rect -18259 -33147 -18198 -33079
rect -23382 -36955 -23305 -36860
rect -23223 -36950 -23146 -36855
rect -23074 -36947 -22997 -36852
rect -23383 -37113 -23306 -37018
rect -23224 -37108 -23147 -37013
rect -23075 -37105 -22998 -37010
rect -24170 -37652 -24093 -37557
rect -24011 -37647 -23934 -37552
rect -23862 -37644 -23785 -37549
rect -24173 -37828 -24096 -37733
rect -24014 -37823 -23937 -37728
rect -23865 -37820 -23788 -37725
rect -24171 -37987 -24094 -37892
rect -24012 -37982 -23935 -37887
rect -23863 -37979 -23786 -37884
rect -24172 -38145 -24095 -38050
rect -24013 -38140 -23936 -38045
rect -23864 -38137 -23787 -38042
rect 4854 55729 4931 55824
rect 5013 55734 5090 55829
rect 5162 55737 5239 55832
rect 4851 55553 4928 55648
rect 5010 55558 5087 55653
rect 5159 55561 5236 55656
rect 4853 55394 4930 55489
rect 5012 55399 5089 55494
rect 5161 55402 5238 55497
rect 4852 55236 4929 55331
rect 5011 55241 5088 55336
rect 5160 55244 5237 55339
rect 4089 54691 4166 54786
rect 4248 54696 4325 54791
rect 4397 54699 4474 54794
rect 4086 54515 4163 54610
rect 4245 54520 4322 54615
rect 4394 54523 4471 54618
rect 4088 54356 4165 54451
rect 4247 54361 4324 54456
rect 4396 54364 4473 54459
rect 4087 54198 4164 54293
rect 4246 54203 4323 54298
rect 4395 54206 4472 54301
rect 2900 53500 2977 53595
rect 2897 53324 2974 53419
rect 2899 53165 2976 53260
rect 2898 53007 2975 53102
rect 2693 52461 2770 52556
rect 2690 52285 2767 52380
rect 2692 52126 2769 52221
rect 2691 51968 2768 52063
rect -3887 49925 -3796 50004
rect -3891 49773 -3800 49852
rect 2839 36925 2916 37020
rect 2836 36749 2913 36844
rect 2838 36590 2915 36685
rect 2837 36432 2914 36527
rect 2631 35665 2708 35760
rect 2628 35489 2705 35584
rect 2630 35330 2707 35425
rect 2629 35172 2706 35267
rect -3954 33116 -3863 33195
rect -3958 32964 -3867 33043
rect -4250 31146 -4159 31225
rect -4254 30994 -4163 31073
rect 3012 19321 3089 19416
rect 3009 19145 3086 19240
rect 3011 18986 3088 19081
rect 3010 18828 3087 18923
rect 2810 18238 2887 18333
rect 2807 18062 2884 18157
rect 2809 17903 2886 17998
rect 2808 17745 2885 17840
rect -3755 15612 -3699 15668
rect -3759 15501 -3703 15557
rect -4098 13685 -4042 13741
rect -4102 13574 -4046 13630
rect 3048 7297 3125 7392
rect 3045 7121 3122 7216
rect 3047 6962 3124 7057
rect 3046 6804 3123 6899
rect 2843 6060 2920 6155
rect 2840 5884 2917 5979
rect 2842 5725 2919 5820
rect 2841 5567 2918 5662
rect -3707 2919 -3651 2975
rect -3711 2808 -3655 2864
rect -4071 984 -4015 1040
rect -4075 873 -4019 929
rect -5294 -22926 -5194 -22845
rect -5295 -23127 -5195 -23046
rect -4927 -24811 -4830 -24701
rect -4929 -25097 -4832 -24987
rect 3091 -11476 3168 -11381
rect 3088 -11652 3165 -11557
rect 3090 -11811 3167 -11716
rect 3089 -11969 3166 -11874
rect 2889 -12517 2966 -12422
rect 2886 -12693 2963 -12598
rect 2888 -12852 2965 -12757
rect 2887 -13010 2964 -12915
rect -3669 -14935 -3613 -14879
rect -3673 -15046 -3617 -14990
rect -4002 -16819 -3932 -16754
rect -4008 -16978 -3938 -16913
rect 3174 -27608 3251 -27513
rect 3171 -27784 3248 -27689
rect 3173 -27943 3250 -27848
rect 3172 -28101 3249 -28006
rect 2980 -28650 3057 -28555
rect 2977 -28826 3054 -28731
rect 2979 -28985 3056 -28890
rect 2978 -29143 3055 -29048
rect -7125 -36620 -7048 -36525
rect -6966 -36615 -6889 -36520
rect -6817 -36612 -6740 -36517
rect -7128 -36796 -7051 -36701
rect -6969 -36791 -6892 -36696
rect -6820 -36788 -6743 -36693
rect -7126 -36955 -7049 -36860
rect -6967 -36950 -6890 -36855
rect -6818 -36947 -6741 -36852
rect -4122 -33175 -4054 -33114
rect -3968 -33153 -3900 -33092
rect -7127 -37113 -7050 -37018
rect -6968 -37108 -6891 -37013
rect -6819 -37105 -6742 -37010
rect -7896 -37656 -7819 -37561
rect -7737 -37651 -7660 -37556
rect -7588 -37648 -7511 -37553
rect -7899 -37832 -7822 -37737
rect -7740 -37827 -7663 -37732
rect -7591 -37824 -7514 -37729
rect -7897 -37991 -7820 -37896
rect -7738 -37986 -7661 -37891
rect -7589 -37983 -7512 -37888
rect -7898 -38149 -7821 -38054
rect -7739 -38144 -7662 -38049
rect -7590 -38141 -7513 -38046
rect 15340 55729 15417 55824
rect 15499 55734 15576 55829
rect 15648 55737 15725 55832
rect 15337 55553 15414 55648
rect 15496 55558 15573 55653
rect 15645 55561 15722 55656
rect 15339 55394 15416 55489
rect 15498 55399 15575 55494
rect 15647 55402 15724 55497
rect 15338 55236 15415 55331
rect 15497 55241 15574 55336
rect 15646 55244 15723 55339
rect 14652 54689 14729 54784
rect 14811 54694 14888 54789
rect 14960 54697 15037 54792
rect 14649 54513 14726 54608
rect 14808 54518 14885 54613
rect 14957 54521 15034 54616
rect 14651 54354 14728 54449
rect 14810 54359 14887 54454
rect 14959 54362 15036 54457
rect 14650 54196 14727 54291
rect 14809 54201 14886 54296
rect 14958 54204 15035 54299
rect 13967 45136 14044 45231
rect 13964 44960 14041 45055
rect 13966 44801 14043 44896
rect 13965 44643 14042 44738
rect 13767 44093 13844 44188
rect 13764 43917 13841 44012
rect 13766 43758 13843 43853
rect 13765 43600 13842 43695
rect 7022 33113 7113 33192
rect 13806 36925 13883 37020
rect 13803 36749 13880 36844
rect 13805 36590 13882 36685
rect 13804 36432 13881 36527
rect 13601 35665 13678 35760
rect 13598 35489 13675 35584
rect 13600 35330 13677 35425
rect 13599 35172 13676 35267
rect 7018 32961 7109 33040
rect 6710 31095 6801 31174
rect 6706 30943 6797 31022
rect 13845 28364 13922 28459
rect 13842 28188 13919 28283
rect 13844 28029 13921 28124
rect 13843 27871 13920 27966
rect 13645 27253 13722 27348
rect 13642 27077 13719 27172
rect 13644 26918 13721 27013
rect 13643 26760 13720 26855
rect 7059 25063 7150 25142
rect 7055 24911 7146 24990
rect 6728 23132 6819 23211
rect 6724 22980 6815 23059
rect 13661 19318 13738 19413
rect 13658 19142 13735 19237
rect 13660 18983 13737 19078
rect 13659 18825 13736 18920
rect 13455 18242 13532 18337
rect 13452 18066 13529 18161
rect 13454 17907 13531 18002
rect 13453 17749 13530 17844
rect 6890 15526 6946 15582
rect 6886 15415 6942 15471
rect 6644 13674 6700 13730
rect 6640 13563 6696 13619
rect 13878 7301 13955 7396
rect 13875 7125 13952 7220
rect 13877 6966 13954 7061
rect 13876 6808 13953 6903
rect 13673 6067 13750 6162
rect 13670 5891 13747 5986
rect 13672 5732 13749 5827
rect 13671 5574 13748 5669
rect 7116 3112 7172 3168
rect 7112 3001 7168 3057
rect 6772 1210 6828 1266
rect 6768 1099 6824 1155
rect 13859 -2550 13936 -2455
rect 13856 -2726 13933 -2631
rect 13858 -2885 13935 -2790
rect 13857 -3043 13934 -2948
rect 13656 -3621 13733 -3526
rect 13653 -3797 13730 -3702
rect 13655 -3956 13732 -3861
rect 13654 -4114 13731 -4019
rect 7099 -6426 7155 -6370
rect 7095 -6537 7151 -6481
rect 6473 -8410 6555 -8328
rect 6638 -8410 6720 -8328
rect 13862 -11476 13939 -11381
rect 13859 -11652 13936 -11557
rect 13861 -11811 13938 -11716
rect 13860 -11969 13937 -11874
rect 13652 -12517 13729 -12422
rect 13649 -12693 13726 -12598
rect 13651 -12852 13728 -12757
rect 13650 -13010 13727 -12915
rect 7105 -14918 7161 -14862
rect 7101 -15029 7157 -14973
rect 6667 -16836 6738 -16765
rect 6663 -17012 6734 -16941
rect 13980 -19566 14057 -19471
rect 13977 -19742 14054 -19647
rect 13979 -19901 14056 -19806
rect 13978 -20059 14055 -19964
rect 13778 -20608 13855 -20513
rect 13775 -20784 13852 -20689
rect 13777 -20943 13854 -20848
rect 13776 -21101 13853 -21006
rect 4852 -36620 4929 -36525
rect 5011 -36615 5088 -36520
rect 5160 -36612 5237 -36517
rect 4849 -36796 4926 -36701
rect 5008 -36791 5085 -36696
rect 5157 -36788 5234 -36693
rect 4851 -36955 4928 -36860
rect 5010 -36950 5087 -36855
rect 5159 -36947 5236 -36852
rect 4850 -37113 4927 -37018
rect 5009 -37108 5086 -37013
rect 5158 -37105 5235 -37010
rect 6666 -25067 6734 -24990
rect 6880 -25051 6948 -24974
rect 7285 -25063 7353 -24987
rect 7446 -25013 7514 -24937
rect 4089 -37656 4166 -37561
rect 4248 -37651 4325 -37556
rect 4397 -37648 4474 -37553
rect 4086 -37832 4163 -37737
rect 4245 -37827 4322 -37732
rect 4394 -37824 4471 -37729
rect 4088 -37991 4165 -37896
rect 4247 -37986 4324 -37891
rect 4396 -37983 4473 -37888
rect 4087 -38149 4164 -38054
rect 4246 -38144 4323 -38049
rect 4395 -38141 4472 -38046
rect 26036 55729 26113 55824
rect 26195 55734 26272 55829
rect 26344 55737 26421 55832
rect 26033 55553 26110 55648
rect 26192 55558 26269 55653
rect 26341 55561 26418 55656
rect 26035 55394 26112 55489
rect 26194 55399 26271 55494
rect 26343 55402 26420 55497
rect 26034 55236 26111 55331
rect 26193 55241 26270 55336
rect 26342 55244 26419 55339
rect 25347 54691 25424 54786
rect 25506 54696 25583 54791
rect 25655 54699 25732 54794
rect 25344 54515 25421 54610
rect 25503 54520 25580 54615
rect 25652 54523 25729 54618
rect 25346 54356 25423 54451
rect 25505 54361 25582 54456
rect 25654 54364 25731 54459
rect 25345 54198 25422 54293
rect 25504 54203 25581 54298
rect 25653 54206 25730 54301
rect 24616 53507 24693 53602
rect 24613 53331 24690 53426
rect 24615 53172 24692 53267
rect 24614 53014 24691 53109
rect 24412 52462 24489 52557
rect 24409 52286 24486 52381
rect 24411 52127 24488 52222
rect 24410 51969 24487 52064
rect 16765 39564 16856 39643
rect 16761 39412 16852 39491
rect 24617 45133 24694 45228
rect 24614 44957 24691 45052
rect 24616 44798 24693 44893
rect 24615 44640 24692 44735
rect 24415 44093 24492 44188
rect 24412 43917 24489 44012
rect 24414 43758 24491 43853
rect 24413 43600 24490 43695
rect 17858 41486 17949 41565
rect 17854 41334 17945 41413
rect 24704 36921 24781 37016
rect 24701 36745 24778 36840
rect 24703 36586 24780 36681
rect 24702 36428 24779 36523
rect 24503 35671 24580 35766
rect 24500 35495 24577 35590
rect 24502 35336 24579 35431
rect 24501 35178 24578 35273
rect 17909 33116 18000 33195
rect 17905 32964 17996 33043
rect 17180 31040 17271 31119
rect 17176 30888 17267 30967
rect 16819 25231 16940 25337
rect 16814 25011 16935 25117
rect 16922 23144 17027 23252
rect 16914 22931 17019 23039
rect 24721 19321 24798 19416
rect 24718 19145 24795 19240
rect 24720 18986 24797 19081
rect 24719 18828 24796 18923
rect 24516 18235 24593 18330
rect 24513 18059 24590 18154
rect 24515 17900 24592 17995
rect 24514 17742 24591 17837
rect 17953 15536 18009 15592
rect 17949 15425 18005 15481
rect 17640 13644 17696 13700
rect 17636 13533 17692 13589
rect 24719 7294 24796 7389
rect 24716 7118 24793 7213
rect 24718 6959 24795 7054
rect 24717 6801 24794 6896
rect 24517 6063 24594 6158
rect 24514 5887 24591 5982
rect 24516 5728 24593 5823
rect 24515 5570 24592 5665
rect 17962 3032 18018 3088
rect 17958 2921 18014 2977
rect 17577 1092 17633 1148
rect 17573 981 17629 1037
rect 24703 -11476 24780 -11381
rect 24700 -11652 24777 -11557
rect 24702 -11811 24779 -11716
rect 24701 -11969 24778 -11874
rect 24502 -12513 24579 -12418
rect 24499 -12689 24576 -12594
rect 24501 -12848 24578 -12753
rect 24500 -13006 24577 -12911
rect 17946 -14966 18002 -14910
rect 17942 -15077 17998 -15021
rect 17448 -16891 17519 -16820
rect 17444 -17067 17515 -16996
rect 24692 -19561 24769 -19466
rect 24689 -19737 24766 -19642
rect 24691 -19896 24768 -19801
rect 24690 -20054 24767 -19959
rect 24485 -20608 24562 -20513
rect 24482 -20784 24559 -20689
rect 24484 -20943 24561 -20848
rect 24483 -21101 24560 -21006
rect 15335 -36620 15412 -36525
rect 15494 -36615 15571 -36520
rect 15643 -36612 15720 -36517
rect 15332 -36796 15409 -36701
rect 15491 -36791 15568 -36696
rect 15640 -36788 15717 -36693
rect 15334 -36955 15411 -36860
rect 15493 -36950 15570 -36855
rect 15642 -36947 15719 -36852
rect 15333 -37113 15410 -37018
rect 15492 -37108 15569 -37013
rect 15641 -37105 15718 -37010
rect 14649 -37664 14726 -37569
rect 14808 -37659 14885 -37564
rect 14957 -37656 15034 -37561
rect 14646 -37840 14723 -37745
rect 14805 -37835 14882 -37740
rect 14954 -37832 15031 -37737
rect 14648 -37999 14725 -37904
rect 14807 -37994 14884 -37899
rect 14956 -37991 15033 -37896
rect 14647 -38157 14724 -38062
rect 14806 -38152 14883 -38057
rect 14955 -38149 15032 -38054
rect 17338 -25055 17421 -24962
rect 17593 -25045 17676 -24952
rect 24741 -27608 24818 -27513
rect 24738 -27784 24815 -27689
rect 24740 -27943 24817 -27848
rect 24739 -28101 24816 -28006
rect 24539 -28650 24616 -28555
rect 24536 -28826 24613 -28731
rect 24538 -28985 24615 -28890
rect 24537 -29143 24614 -29048
rect 17525 -33157 17583 -33093
rect 17683 -33155 17741 -33091
rect 37541 53503 37618 53598
rect 37700 53508 37777 53603
rect 37849 53511 37926 53606
rect 37538 53327 37615 53422
rect 37697 53332 37774 53427
rect 37846 53335 37923 53430
rect 37540 53168 37617 53263
rect 37699 53173 37776 53268
rect 37848 53176 37925 53271
rect 37539 53010 37616 53105
rect 37698 53015 37775 53110
rect 37847 53018 37924 53113
rect 36859 52452 36936 52547
rect 37018 52457 37095 52552
rect 37167 52460 37244 52555
rect 36856 52276 36933 52371
rect 37015 52281 37092 52376
rect 37164 52284 37241 52379
rect 36858 52117 36935 52212
rect 37017 52122 37094 52217
rect 37166 52125 37243 52220
rect 36857 51959 36934 52054
rect 37016 51964 37093 52059
rect 37165 51967 37242 52062
rect 35592 45136 35669 45231
rect 35589 44960 35666 45055
rect 35591 44801 35668 44896
rect 35590 44643 35667 44738
rect 35389 44096 35466 44191
rect 35386 43920 35463 44015
rect 35388 43761 35465 43856
rect 35387 43603 35464 43698
rect 37541 45126 37618 45221
rect 37700 45131 37777 45226
rect 37849 45134 37926 45229
rect 37538 44950 37615 45045
rect 37697 44955 37774 45050
rect 37846 44958 37923 45053
rect 37540 44791 37617 44886
rect 37699 44796 37776 44891
rect 37848 44799 37925 44894
rect 37539 44633 37616 44728
rect 37698 44638 37775 44733
rect 37847 44641 37924 44736
rect 36855 44083 36932 44178
rect 37014 44088 37091 44183
rect 37163 44091 37240 44186
rect 36852 43907 36929 44002
rect 37011 43912 37088 44007
rect 37160 43915 37237 44010
rect 36854 43748 36931 43843
rect 37013 43753 37090 43848
rect 37162 43756 37239 43851
rect 36853 43590 36930 43685
rect 37012 43595 37089 43690
rect 37161 43598 37238 43693
rect 28811 41610 28902 41689
rect 28807 41458 28898 41537
rect 28481 39653 28572 39732
rect 28477 39501 28568 39580
rect 35612 36921 35689 37016
rect 35609 36745 35686 36840
rect 35611 36586 35688 36681
rect 35610 36428 35687 36523
rect 35407 35665 35484 35760
rect 35404 35489 35481 35584
rect 35406 35330 35483 35425
rect 35405 35172 35482 35267
rect 37541 36903 37618 36998
rect 37700 36908 37777 37003
rect 37849 36911 37926 37006
rect 37538 36727 37615 36822
rect 37697 36732 37774 36827
rect 37846 36735 37923 36830
rect 37540 36568 37617 36663
rect 37699 36573 37776 36668
rect 37848 36576 37925 36671
rect 37539 36410 37616 36505
rect 37698 36415 37775 36510
rect 37847 36418 37924 36513
rect 36851 35656 36928 35751
rect 37010 35661 37087 35756
rect 37159 35664 37236 35759
rect 36848 35480 36925 35575
rect 37007 35485 37084 35580
rect 37156 35488 37233 35583
rect 36850 35321 36927 35416
rect 37009 35326 37086 35421
rect 37158 35329 37235 35424
rect 36849 35163 36926 35258
rect 37008 35168 37085 35263
rect 37157 35171 37234 35266
rect 28825 33116 28916 33195
rect 28821 32964 28912 33043
rect 28550 31150 28641 31229
rect 28546 30998 28637 31077
rect 37545 28346 37622 28441
rect 37704 28351 37781 28446
rect 37853 28354 37930 28449
rect 37542 28170 37619 28265
rect 37701 28175 37778 28270
rect 37850 28178 37927 28273
rect 37544 28011 37621 28106
rect 37703 28016 37780 28111
rect 37852 28019 37929 28114
rect 37543 27853 37620 27948
rect 37702 27858 37779 27953
rect 37851 27861 37928 27956
rect 36851 27248 36928 27343
rect 37010 27253 37087 27348
rect 37159 27256 37236 27351
rect 36848 27072 36925 27167
rect 37007 27077 37084 27172
rect 37156 27080 37233 27175
rect 36850 26913 36927 27008
rect 37009 26918 37086 27013
rect 37158 26921 37235 27016
rect 36849 26755 36926 26850
rect 37008 26760 37085 26855
rect 37157 26763 37234 26858
rect 35623 19321 35700 19416
rect 35620 19145 35697 19240
rect 35622 18986 35699 19081
rect 35621 18828 35698 18923
rect 35417 18231 35494 18326
rect 35414 18055 35491 18150
rect 35416 17896 35493 17991
rect 35415 17738 35492 17833
rect 37541 19295 37618 19390
rect 37700 19300 37777 19395
rect 37849 19303 37926 19398
rect 37538 19119 37615 19214
rect 37697 19124 37774 19219
rect 37846 19127 37923 19222
rect 37540 18960 37617 19055
rect 37699 18965 37776 19060
rect 37848 18968 37925 19063
rect 37539 18802 37616 18897
rect 37698 18807 37775 18902
rect 37847 18810 37924 18905
rect 36855 18213 36932 18308
rect 37014 18218 37091 18313
rect 37163 18221 37240 18316
rect 36852 18037 36929 18132
rect 37011 18042 37088 18137
rect 37160 18045 37237 18140
rect 36854 17878 36931 17973
rect 37013 17883 37090 17978
rect 37162 17886 37239 17981
rect 36853 17720 36930 17815
rect 37012 17725 37089 17820
rect 37161 17728 37238 17823
rect 28864 15529 28920 15585
rect 28860 15418 28916 15474
rect 28540 13667 28596 13723
rect 28536 13556 28592 13612
rect 35391 7297 35468 7392
rect 35388 7121 35465 7216
rect 35390 6962 35467 7057
rect 35389 6804 35466 6899
rect 35190 6060 35267 6155
rect 35187 5884 35264 5979
rect 35189 5725 35266 5820
rect 35188 5567 35265 5662
rect 37549 7276 37626 7371
rect 37708 7281 37785 7376
rect 37857 7284 37934 7379
rect 37546 7100 37623 7195
rect 37705 7105 37782 7200
rect 37854 7108 37931 7203
rect 37548 6941 37625 7036
rect 37707 6946 37784 7041
rect 37856 6949 37933 7044
rect 37547 6783 37624 6878
rect 37706 6788 37783 6883
rect 37855 6791 37932 6886
rect 36859 6056 36936 6151
rect 37018 6061 37095 6156
rect 37167 6064 37244 6159
rect 36856 5880 36933 5975
rect 37015 5885 37092 5980
rect 37164 5888 37241 5983
rect 36858 5721 36935 5816
rect 37017 5726 37094 5821
rect 37166 5729 37243 5824
rect 36857 5563 36934 5658
rect 37016 5568 37093 5663
rect 37165 5571 37242 5666
rect 28622 2807 28678 2863
rect 28618 2696 28674 2752
rect 28348 895 28404 951
rect 28344 784 28400 840
rect 37541 -2575 37618 -2480
rect 37700 -2570 37777 -2475
rect 37849 -2567 37926 -2472
rect 37538 -2751 37615 -2656
rect 37697 -2746 37774 -2651
rect 37846 -2743 37923 -2648
rect 37540 -2910 37617 -2815
rect 37699 -2905 37776 -2810
rect 37848 -2902 37925 -2807
rect 37539 -3068 37616 -2973
rect 37698 -3063 37775 -2968
rect 37847 -3060 37924 -2965
rect 36851 -3645 36928 -3550
rect 37010 -3640 37087 -3545
rect 37159 -3637 37236 -3542
rect 36848 -3821 36925 -3726
rect 37007 -3816 37084 -3721
rect 37156 -3813 37233 -3718
rect 36850 -3980 36927 -3885
rect 37009 -3975 37086 -3880
rect 37158 -3972 37235 -3877
rect 36849 -4138 36926 -4043
rect 37008 -4133 37085 -4038
rect 37157 -4130 37234 -4035
rect 35400 -11472 35477 -11377
rect 35397 -11648 35474 -11553
rect 35399 -11807 35476 -11712
rect 35398 -11965 35475 -11870
rect 35199 -12517 35276 -12422
rect 35196 -12693 35273 -12598
rect 35198 -12852 35275 -12757
rect 35197 -13010 35274 -12915
rect 37541 -11496 37618 -11401
rect 37700 -11491 37777 -11396
rect 37849 -11488 37926 -11393
rect 37538 -11672 37615 -11577
rect 37697 -11667 37774 -11572
rect 37846 -11664 37923 -11569
rect 37540 -11831 37617 -11736
rect 37699 -11826 37776 -11731
rect 37848 -11823 37925 -11728
rect 37539 -11989 37616 -11894
rect 37698 -11984 37775 -11889
rect 37847 -11981 37924 -11886
rect 36855 -12535 36932 -12440
rect 37014 -12530 37091 -12435
rect 37163 -12527 37240 -12432
rect 36852 -12711 36929 -12616
rect 37011 -12706 37088 -12611
rect 37160 -12703 37237 -12608
rect 36854 -12870 36931 -12775
rect 37013 -12865 37090 -12770
rect 37162 -12862 37239 -12767
rect 36853 -13028 36930 -12933
rect 37012 -13023 37089 -12928
rect 37161 -13020 37238 -12925
rect 28651 -14960 28707 -14904
rect 28647 -15071 28703 -15015
rect 28339 -16832 28410 -16761
rect 28335 -17008 28406 -16937
rect 35416 -19566 35493 -19471
rect 35413 -19742 35490 -19647
rect 35415 -19901 35492 -19806
rect 35414 -20059 35491 -19964
rect 35213 -20608 35290 -20513
rect 35210 -20784 35287 -20689
rect 35212 -20943 35289 -20848
rect 35211 -21101 35288 -21006
rect 37541 -19578 37618 -19483
rect 37700 -19573 37777 -19478
rect 37849 -19570 37926 -19475
rect 37538 -19754 37615 -19659
rect 37697 -19749 37774 -19654
rect 37846 -19746 37923 -19651
rect 37540 -19913 37617 -19818
rect 37699 -19908 37776 -19813
rect 37848 -19905 37925 -19810
rect 37539 -20071 37616 -19976
rect 37698 -20066 37775 -19971
rect 37847 -20063 37924 -19968
rect 36851 -20618 36928 -20523
rect 37010 -20613 37087 -20518
rect 37159 -20610 37236 -20515
rect 36848 -20794 36925 -20699
rect 37007 -20789 37084 -20694
rect 37156 -20786 37233 -20691
rect 36850 -20953 36927 -20858
rect 37009 -20948 37086 -20853
rect 37158 -20945 37235 -20850
rect 36849 -21111 36926 -21016
rect 37008 -21106 37085 -21011
rect 37157 -21103 37234 -21008
rect 28407 -24969 28463 -24912
rect 28314 -25072 28370 -25015
rect 37541 -27621 37618 -27526
rect 37700 -27616 37777 -27521
rect 37849 -27613 37926 -27518
rect 37538 -27797 37615 -27702
rect 37697 -27792 37774 -27697
rect 37846 -27789 37923 -27694
rect 37540 -27956 37617 -27861
rect 37699 -27951 37776 -27856
rect 37848 -27948 37925 -27853
rect 37539 -28114 37616 -28019
rect 37698 -28109 37775 -28014
rect 37847 -28106 37924 -28011
rect 36859 -28657 36936 -28562
rect 37018 -28652 37095 -28557
rect 37167 -28649 37244 -28554
rect 36856 -28833 36933 -28738
rect 37015 -28828 37092 -28733
rect 37164 -28825 37241 -28730
rect 36858 -28992 36935 -28897
rect 37017 -28987 37094 -28892
rect 37166 -28984 37243 -28889
rect 36857 -29150 36934 -29055
rect 37016 -29145 37093 -29050
rect 37165 -29142 37242 -29047
rect 26040 -36620 26117 -36525
rect 26199 -36615 26276 -36520
rect 26348 -36612 26425 -36517
rect 26037 -36796 26114 -36701
rect 26196 -36791 26273 -36696
rect 26345 -36788 26422 -36693
rect 26039 -36955 26116 -36860
rect 26198 -36950 26275 -36855
rect 26347 -36947 26424 -36852
rect 26038 -37113 26115 -37018
rect 26197 -37108 26274 -37013
rect 26346 -37105 26423 -37010
rect 25353 -37653 25430 -37558
rect 25512 -37648 25589 -37553
rect 25661 -37645 25738 -37550
rect 25350 -37829 25427 -37734
rect 25509 -37824 25586 -37729
rect 25658 -37821 25735 -37726
rect 25352 -37988 25429 -37893
rect 25511 -37983 25588 -37888
rect 25660 -37980 25737 -37885
rect 25351 -38146 25428 -38051
rect 25510 -38141 25587 -38046
rect 25659 -38138 25736 -38043
<< metal3 >>
rect -70936 55834 37954 55868
rect -70936 55832 -44612 55834
rect -70936 55829 -65367 55832
rect -70936 55824 -65516 55829
rect -70936 55729 -65675 55824
rect -65598 55734 -65516 55824
rect -65439 55737 -65367 55829
rect -65290 55831 -44612 55832
rect -65290 55828 -54966 55831
rect -65290 55823 -55115 55828
rect -65290 55737 -55274 55823
rect -65439 55734 -55274 55737
rect -65598 55729 -55274 55734
rect -70936 55728 -55274 55729
rect -55197 55733 -55115 55823
rect -55038 55736 -54966 55828
rect -54889 55826 -44761 55831
rect -54889 55736 -44920 55826
rect -55038 55733 -44920 55736
rect -55197 55731 -44920 55733
rect -44843 55736 -44761 55826
rect -44684 55739 -44612 55831
rect -44535 55832 37954 55834
rect -44535 55831 -6818 55832
rect -44535 55828 -34376 55831
rect -44535 55823 -34525 55828
rect -44535 55739 -34684 55823
rect -44684 55736 -34684 55739
rect -44843 55731 -34684 55736
rect -55197 55728 -34684 55731
rect -34607 55733 -34525 55823
rect -34448 55736 -34376 55828
rect -34299 55828 -23067 55831
rect -34299 55823 -23216 55828
rect -34299 55736 -23375 55823
rect -34448 55733 -23375 55736
rect -34607 55728 -23375 55733
rect -23298 55733 -23216 55823
rect -23139 55736 -23067 55828
rect -22990 55829 -6818 55831
rect -22990 55824 -6967 55829
rect -22990 55736 -7126 55824
rect -23139 55733 -7126 55736
rect -23298 55729 -7126 55733
rect -7049 55734 -6967 55824
rect -6890 55737 -6818 55829
rect -6741 55829 5162 55832
rect -6741 55824 5013 55829
rect -6741 55737 4854 55824
rect -6890 55734 4854 55737
rect -7049 55729 4854 55734
rect 4931 55734 5013 55824
rect 5090 55737 5162 55829
rect 5239 55829 15648 55832
rect 5239 55824 15499 55829
rect 5239 55737 15340 55824
rect 5090 55734 15340 55737
rect 4931 55729 15340 55734
rect 15417 55734 15499 55824
rect 15576 55737 15648 55829
rect 15725 55829 26344 55832
rect 15725 55824 26195 55829
rect 15725 55737 26036 55824
rect 15576 55734 26036 55737
rect 15417 55729 26036 55734
rect 26113 55734 26195 55824
rect 26272 55737 26344 55829
rect 26421 55737 37954 55832
rect 26272 55734 37954 55737
rect 26113 55729 37954 55734
rect -23298 55728 37954 55729
rect -70936 55658 37954 55728
rect -70936 55656 -44615 55658
rect -70936 55653 -65370 55656
rect -70936 55648 -65519 55653
rect -70936 55553 -65678 55648
rect -65601 55558 -65519 55648
rect -65442 55561 -65370 55653
rect -65293 55655 -44615 55656
rect -65293 55652 -54969 55655
rect -65293 55647 -55118 55652
rect -65293 55561 -55277 55647
rect -65442 55558 -55277 55561
rect -65601 55553 -55277 55558
rect -70936 55552 -55277 55553
rect -55200 55557 -55118 55647
rect -55041 55560 -54969 55652
rect -54892 55650 -44764 55655
rect -54892 55560 -44923 55650
rect -55041 55557 -44923 55560
rect -55200 55555 -44923 55557
rect -44846 55560 -44764 55650
rect -44687 55563 -44615 55655
rect -44538 55656 37954 55658
rect -44538 55655 -6821 55656
rect -44538 55652 -34379 55655
rect -44538 55647 -34528 55652
rect -44538 55563 -34687 55647
rect -44687 55560 -34687 55563
rect -44846 55555 -34687 55560
rect -55200 55552 -34687 55555
rect -34610 55557 -34528 55647
rect -34451 55560 -34379 55652
rect -34302 55652 -23070 55655
rect -34302 55647 -23219 55652
rect -34302 55560 -23378 55647
rect -34451 55557 -23378 55560
rect -34610 55552 -23378 55557
rect -23301 55557 -23219 55647
rect -23142 55560 -23070 55652
rect -22993 55653 -6821 55655
rect -22993 55648 -6970 55653
rect -22993 55560 -7129 55648
rect -23142 55557 -7129 55560
rect -23301 55553 -7129 55557
rect -7052 55558 -6970 55648
rect -6893 55561 -6821 55653
rect -6744 55653 5159 55656
rect -6744 55648 5010 55653
rect -6744 55561 4851 55648
rect -6893 55558 4851 55561
rect -7052 55553 4851 55558
rect 4928 55558 5010 55648
rect 5087 55561 5159 55653
rect 5236 55653 15645 55656
rect 5236 55648 15496 55653
rect 5236 55561 15337 55648
rect 5087 55558 15337 55561
rect 4928 55553 15337 55558
rect 15414 55558 15496 55648
rect 15573 55561 15645 55653
rect 15722 55653 26341 55656
rect 15722 55648 26192 55653
rect 15722 55561 26033 55648
rect 15573 55558 26033 55561
rect 15414 55553 26033 55558
rect 26110 55558 26192 55648
rect 26269 55561 26341 55653
rect 26418 55561 37954 55656
rect 26269 55558 37954 55561
rect 26110 55553 37954 55558
rect -23301 55552 37954 55553
rect -70936 55499 37954 55552
rect -70936 55497 -44613 55499
rect -70936 55494 -65368 55497
rect -70936 55489 -65517 55494
rect -70936 55394 -65676 55489
rect -65599 55399 -65517 55489
rect -65440 55402 -65368 55494
rect -65291 55496 -44613 55497
rect -65291 55493 -54967 55496
rect -65291 55488 -55116 55493
rect -65291 55402 -55275 55488
rect -65440 55399 -55275 55402
rect -65599 55394 -55275 55399
rect -70936 55393 -55275 55394
rect -55198 55398 -55116 55488
rect -55039 55401 -54967 55493
rect -54890 55491 -44762 55496
rect -54890 55401 -44921 55491
rect -55039 55398 -44921 55401
rect -55198 55396 -44921 55398
rect -44844 55401 -44762 55491
rect -44685 55404 -44613 55496
rect -44536 55497 37954 55499
rect -44536 55496 -6819 55497
rect -44536 55493 -34377 55496
rect -44536 55488 -34526 55493
rect -44536 55404 -34685 55488
rect -44685 55401 -34685 55404
rect -44844 55396 -34685 55401
rect -55198 55393 -34685 55396
rect -34608 55398 -34526 55488
rect -34449 55401 -34377 55493
rect -34300 55493 -23068 55496
rect -34300 55488 -23217 55493
rect -34300 55401 -23376 55488
rect -34449 55398 -23376 55401
rect -34608 55393 -23376 55398
rect -23299 55398 -23217 55488
rect -23140 55401 -23068 55493
rect -22991 55494 -6819 55496
rect -22991 55489 -6968 55494
rect -22991 55401 -7127 55489
rect -23140 55398 -7127 55401
rect -23299 55394 -7127 55398
rect -7050 55399 -6968 55489
rect -6891 55402 -6819 55494
rect -6742 55494 5161 55497
rect -6742 55489 5012 55494
rect -6742 55402 4853 55489
rect -6891 55399 4853 55402
rect -7050 55394 4853 55399
rect 4930 55399 5012 55489
rect 5089 55402 5161 55494
rect 5238 55494 15647 55497
rect 5238 55489 15498 55494
rect 5238 55402 15339 55489
rect 5089 55399 15339 55402
rect 4930 55394 15339 55399
rect 15416 55399 15498 55489
rect 15575 55402 15647 55494
rect 15724 55494 26343 55497
rect 15724 55489 26194 55494
rect 15724 55402 26035 55489
rect 15575 55399 26035 55402
rect 15416 55394 26035 55399
rect 26112 55399 26194 55489
rect 26271 55402 26343 55494
rect 26420 55402 37954 55497
rect 26271 55399 37954 55402
rect 26112 55394 37954 55399
rect -23299 55393 37954 55394
rect -70936 55341 37954 55393
rect -70936 55339 -44614 55341
rect -70936 55336 -65369 55339
rect -70936 55331 -65518 55336
rect -70936 55236 -65677 55331
rect -65600 55241 -65518 55331
rect -65441 55244 -65369 55336
rect -65292 55338 -44614 55339
rect -65292 55335 -54968 55338
rect -65292 55330 -55117 55335
rect -65292 55244 -55276 55330
rect -65441 55241 -55276 55244
rect -65600 55236 -55276 55241
rect -70936 55235 -55276 55236
rect -55199 55240 -55117 55330
rect -55040 55243 -54968 55335
rect -54891 55333 -44763 55338
rect -54891 55243 -44922 55333
rect -55040 55240 -44922 55243
rect -55199 55238 -44922 55240
rect -44845 55243 -44763 55333
rect -44686 55246 -44614 55338
rect -44537 55339 37954 55341
rect -44537 55338 -6820 55339
rect -44537 55335 -34378 55338
rect -44537 55330 -34527 55335
rect -44537 55246 -34686 55330
rect -44686 55243 -34686 55246
rect -44845 55238 -34686 55243
rect -55199 55235 -34686 55238
rect -34609 55240 -34527 55330
rect -34450 55243 -34378 55335
rect -34301 55335 -23069 55338
rect -34301 55330 -23218 55335
rect -34301 55243 -23377 55330
rect -34450 55240 -23377 55243
rect -34609 55235 -23377 55240
rect -23300 55240 -23218 55330
rect -23141 55243 -23069 55335
rect -22992 55336 -6820 55338
rect -22992 55331 -6969 55336
rect -22992 55243 -7128 55331
rect -23141 55240 -7128 55243
rect -23300 55236 -7128 55240
rect -7051 55241 -6969 55331
rect -6892 55244 -6820 55336
rect -6743 55336 5160 55339
rect -6743 55331 5011 55336
rect -6743 55244 4852 55331
rect -6892 55241 4852 55244
rect -7051 55236 4852 55241
rect 4929 55241 5011 55331
rect 5088 55244 5160 55336
rect 5237 55336 15646 55339
rect 5237 55331 15497 55336
rect 5237 55244 15338 55331
rect 5088 55241 15338 55244
rect 4929 55236 15338 55241
rect 15415 55241 15497 55331
rect 15574 55244 15646 55336
rect 15723 55336 26342 55339
rect 15723 55331 26193 55336
rect 15723 55244 26034 55331
rect 15574 55241 26034 55244
rect 15415 55236 26034 55241
rect 26111 55241 26193 55331
rect 26270 55244 26342 55336
rect 26419 55244 37954 55339
rect 26270 55241 37954 55244
rect 26111 55236 37954 55241
rect -23300 55235 37954 55236
rect -70936 55222 37954 55235
rect -45498 54834 -45349 54837
rect -45599 54831 -45349 54834
rect -70936 54809 37954 54831
rect -70936 54806 -45434 54809
rect -70936 54801 -45583 54806
rect -70936 54796 -45742 54801
rect -70936 54794 -55614 54796
rect -70936 54791 -66054 54794
rect -70936 54786 -66203 54791
rect -70936 54691 -66362 54786
rect -66285 54696 -66203 54786
rect -66126 54699 -66054 54791
rect -65977 54793 -55614 54794
rect -65977 54788 -55763 54793
rect -65977 54699 -55922 54788
rect -66126 54696 -55922 54699
rect -66285 54693 -55922 54696
rect -55845 54698 -55763 54788
rect -55686 54701 -55614 54793
rect -55537 54706 -45742 54796
rect -45665 54711 -45583 54801
rect -45506 54714 -45434 54806
rect -45357 54796 37954 54809
rect -45357 54793 -35066 54796
rect -45357 54788 -35215 54793
rect -45357 54714 -35374 54788
rect -45506 54711 -35374 54714
rect -45665 54706 -35374 54711
rect -55537 54701 -35374 54706
rect -55686 54698 -35374 54701
rect -55845 54693 -35374 54698
rect -35297 54698 -35215 54788
rect -35138 54701 -35066 54793
rect -34989 54793 -7591 54796
rect -34989 54792 -7740 54793
rect -34989 54789 -23862 54792
rect -34989 54784 -24011 54789
rect -34989 54701 -24170 54784
rect -35138 54698 -24170 54701
rect -35297 54693 -24170 54698
rect -66285 54691 -24170 54693
rect -70936 54689 -24170 54691
rect -24093 54694 -24011 54784
rect -23934 54697 -23862 54789
rect -23785 54788 -7740 54792
rect -23785 54697 -7899 54788
rect -23934 54694 -7899 54697
rect -24093 54693 -7899 54694
rect -7822 54698 -7740 54788
rect -7663 54701 -7591 54793
rect -7514 54794 37954 54796
rect -7514 54791 4397 54794
rect -7514 54786 4248 54791
rect -7514 54701 4089 54786
rect -7663 54698 4089 54701
rect -7822 54693 4089 54698
rect -24093 54691 4089 54693
rect 4166 54696 4248 54786
rect 4325 54699 4397 54791
rect 4474 54792 25655 54794
rect 4474 54789 14960 54792
rect 4474 54784 14811 54789
rect 4474 54699 14652 54784
rect 4325 54696 14652 54699
rect 4166 54691 14652 54696
rect -24093 54689 14652 54691
rect 14729 54694 14811 54784
rect 14888 54697 14960 54789
rect 15037 54791 25655 54792
rect 15037 54786 25506 54791
rect 15037 54697 25347 54786
rect 14888 54694 25347 54697
rect 14729 54691 25347 54694
rect 25424 54696 25506 54786
rect 25583 54699 25655 54791
rect 25732 54699 37954 54794
rect 25583 54696 37954 54699
rect 25424 54691 37954 54696
rect 14729 54689 37954 54691
rect -70936 54633 37954 54689
rect -70936 54630 -45437 54633
rect -70936 54625 -45586 54630
rect -70936 54620 -45745 54625
rect -70936 54618 -55617 54620
rect -70936 54615 -66057 54618
rect -70936 54610 -66206 54615
rect -70936 54515 -66365 54610
rect -66288 54520 -66206 54610
rect -66129 54523 -66057 54615
rect -65980 54617 -55617 54618
rect -65980 54612 -55766 54617
rect -65980 54523 -55925 54612
rect -66129 54520 -55925 54523
rect -66288 54517 -55925 54520
rect -55848 54522 -55766 54612
rect -55689 54525 -55617 54617
rect -55540 54530 -45745 54620
rect -45668 54535 -45586 54625
rect -45509 54538 -45437 54630
rect -45360 54620 37954 54633
rect -45360 54617 -35069 54620
rect -45360 54612 -35218 54617
rect -45360 54538 -35377 54612
rect -45509 54535 -35377 54538
rect -45668 54530 -35377 54535
rect -55540 54525 -35377 54530
rect -55689 54522 -35377 54525
rect -55848 54517 -35377 54522
rect -35300 54522 -35218 54612
rect -35141 54525 -35069 54617
rect -34992 54617 -7594 54620
rect -34992 54616 -7743 54617
rect -34992 54613 -23865 54616
rect -34992 54608 -24014 54613
rect -34992 54525 -24173 54608
rect -35141 54522 -24173 54525
rect -35300 54517 -24173 54522
rect -66288 54515 -24173 54517
rect -70936 54513 -24173 54515
rect -24096 54518 -24014 54608
rect -23937 54521 -23865 54613
rect -23788 54612 -7743 54616
rect -23788 54521 -7902 54612
rect -23937 54518 -7902 54521
rect -24096 54517 -7902 54518
rect -7825 54522 -7743 54612
rect -7666 54525 -7594 54617
rect -7517 54618 37954 54620
rect -7517 54615 4394 54618
rect -7517 54610 4245 54615
rect -7517 54525 4086 54610
rect -7666 54522 4086 54525
rect -7825 54517 4086 54522
rect -24096 54515 4086 54517
rect 4163 54520 4245 54610
rect 4322 54523 4394 54615
rect 4471 54616 25652 54618
rect 4471 54613 14957 54616
rect 4471 54608 14808 54613
rect 4471 54523 14649 54608
rect 4322 54520 14649 54523
rect 4163 54515 14649 54520
rect -24096 54513 14649 54515
rect 14726 54518 14808 54608
rect 14885 54521 14957 54613
rect 15034 54615 25652 54616
rect 15034 54610 25503 54615
rect 15034 54521 25344 54610
rect 14885 54518 25344 54521
rect 14726 54515 25344 54518
rect 25421 54520 25503 54610
rect 25580 54523 25652 54615
rect 25729 54523 37954 54618
rect 25580 54520 37954 54523
rect 25421 54515 37954 54520
rect 14726 54513 37954 54515
rect -70936 54474 37954 54513
rect -70936 54471 -45435 54474
rect -70936 54466 -45584 54471
rect -70936 54461 -45743 54466
rect -70936 54459 -55615 54461
rect -70936 54456 -66055 54459
rect -70936 54451 -66204 54456
rect -70936 54356 -66363 54451
rect -66286 54361 -66204 54451
rect -66127 54364 -66055 54456
rect -65978 54458 -55615 54459
rect -65978 54453 -55764 54458
rect -65978 54364 -55923 54453
rect -66127 54361 -55923 54364
rect -66286 54358 -55923 54361
rect -55846 54363 -55764 54453
rect -55687 54366 -55615 54458
rect -55538 54371 -45743 54461
rect -45666 54376 -45584 54466
rect -45507 54379 -45435 54471
rect -45358 54461 37954 54474
rect -45358 54458 -35067 54461
rect -45358 54453 -35216 54458
rect -45358 54379 -35375 54453
rect -45507 54376 -35375 54379
rect -45666 54371 -35375 54376
rect -55538 54366 -35375 54371
rect -55687 54363 -35375 54366
rect -55846 54358 -35375 54363
rect -35298 54363 -35216 54453
rect -35139 54366 -35067 54458
rect -34990 54458 -7592 54461
rect -34990 54457 -7741 54458
rect -34990 54454 -23863 54457
rect -34990 54449 -24012 54454
rect -34990 54366 -24171 54449
rect -35139 54363 -24171 54366
rect -35298 54358 -24171 54363
rect -66286 54356 -24171 54358
rect -70936 54354 -24171 54356
rect -24094 54359 -24012 54449
rect -23935 54362 -23863 54454
rect -23786 54453 -7741 54457
rect -23786 54362 -7900 54453
rect -23935 54359 -7900 54362
rect -24094 54358 -7900 54359
rect -7823 54363 -7741 54453
rect -7664 54366 -7592 54458
rect -7515 54459 37954 54461
rect -7515 54456 4396 54459
rect -7515 54451 4247 54456
rect -7515 54366 4088 54451
rect -7664 54363 4088 54366
rect -7823 54358 4088 54363
rect -24094 54356 4088 54358
rect 4165 54361 4247 54451
rect 4324 54364 4396 54456
rect 4473 54457 25654 54459
rect 4473 54454 14959 54457
rect 4473 54449 14810 54454
rect 4473 54364 14651 54449
rect 4324 54361 14651 54364
rect 4165 54356 14651 54361
rect -24094 54354 14651 54356
rect 14728 54359 14810 54449
rect 14887 54362 14959 54454
rect 15036 54456 25654 54457
rect 15036 54451 25505 54456
rect 15036 54362 25346 54451
rect 14887 54359 25346 54362
rect 14728 54356 25346 54359
rect 25423 54361 25505 54451
rect 25582 54364 25654 54456
rect 25731 54364 37954 54459
rect 25582 54361 37954 54364
rect 25423 54356 37954 54361
rect 14728 54354 37954 54356
rect -70936 54316 37954 54354
rect -70936 54313 -45436 54316
rect -70936 54308 -45585 54313
rect -70936 54303 -45744 54308
rect -70936 54301 -55616 54303
rect -70936 54298 -66056 54301
rect -70936 54293 -66205 54298
rect -70936 54198 -66364 54293
rect -66287 54203 -66205 54293
rect -66128 54206 -66056 54298
rect -65979 54300 -55616 54301
rect -65979 54295 -55765 54300
rect -65979 54206 -55924 54295
rect -66128 54203 -55924 54206
rect -66287 54200 -55924 54203
rect -55847 54205 -55765 54295
rect -55688 54208 -55616 54300
rect -55539 54213 -45744 54303
rect -45667 54218 -45585 54308
rect -45508 54221 -45436 54313
rect -45359 54303 37954 54316
rect -45359 54300 -35068 54303
rect -45359 54295 -35217 54300
rect -45359 54221 -35376 54295
rect -45508 54218 -35376 54221
rect -45667 54213 -35376 54218
rect -55539 54208 -35376 54213
rect -55688 54205 -35376 54208
rect -55847 54200 -35376 54205
rect -35299 54205 -35217 54295
rect -35140 54208 -35068 54300
rect -34991 54300 -7593 54303
rect -34991 54299 -7742 54300
rect -34991 54296 -23864 54299
rect -34991 54291 -24013 54296
rect -34991 54208 -24172 54291
rect -35140 54205 -24172 54208
rect -35299 54200 -24172 54205
rect -66287 54198 -24172 54200
rect -70936 54196 -24172 54198
rect -24095 54201 -24013 54291
rect -23936 54204 -23864 54296
rect -23787 54295 -7742 54299
rect -23787 54204 -7901 54295
rect -23936 54201 -7901 54204
rect -24095 54200 -7901 54201
rect -7824 54205 -7742 54295
rect -7665 54208 -7593 54300
rect -7516 54301 37954 54303
rect -7516 54298 4395 54301
rect -7516 54293 4246 54298
rect -7516 54208 4087 54293
rect -7665 54205 4087 54208
rect -7824 54200 4087 54205
rect -24095 54198 4087 54200
rect 4164 54203 4246 54293
rect 4323 54206 4395 54298
rect 4472 54299 25653 54301
rect 4472 54296 14958 54299
rect 4472 54291 14809 54296
rect 4472 54206 14650 54291
rect 4323 54203 14650 54206
rect 4164 54198 14650 54203
rect -24095 54196 14650 54198
rect 14727 54201 14809 54291
rect 14886 54204 14958 54296
rect 15035 54298 25653 54299
rect 15035 54293 25504 54298
rect 15035 54204 25345 54293
rect 14886 54201 25345 54204
rect 14727 54198 25345 54201
rect 25422 54203 25504 54293
rect 25581 54206 25653 54298
rect 25730 54206 37954 54301
rect 25581 54203 37954 54206
rect 25422 54198 37954 54203
rect 14727 54196 37954 54198
rect -70936 54185 37954 54196
rect -24189 54184 -23779 54185
rect 14633 54184 15043 54185
rect -44767 53634 -44666 53638
rect -36027 53634 -35933 53639
rect -70936 53615 37954 53634
rect -70936 53607 -36016 53615
rect -70936 53604 -69895 53607
rect -70936 53599 -70044 53604
rect -70936 53504 -70203 53599
rect -70126 53509 -70044 53599
rect -69967 53512 -69895 53604
rect -69818 53602 -36016 53607
rect -69818 53512 -46395 53602
rect -69967 53509 -46395 53512
rect -70126 53507 -46395 53509
rect -46318 53520 -36016 53602
rect -35939 53606 37954 53615
rect -35939 53603 37849 53606
rect -35939 53602 37700 53603
rect -35939 53520 -11204 53602
rect -46318 53507 -11204 53520
rect -11127 53595 24616 53602
rect -11127 53507 2900 53595
rect -70126 53504 2900 53507
rect -70936 53500 2900 53504
rect 2977 53507 24616 53595
rect 24693 53598 37700 53602
rect 24693 53507 37541 53598
rect 2977 53503 37541 53507
rect 37618 53508 37700 53598
rect 37777 53511 37849 53603
rect 37926 53511 37954 53606
rect 37777 53508 37954 53511
rect 37618 53503 37954 53508
rect 2977 53500 37954 53503
rect -70936 53439 37954 53500
rect -70936 53431 -36019 53439
rect -70936 53428 -69898 53431
rect -70936 53423 -70047 53428
rect -70936 53328 -70206 53423
rect -70129 53333 -70047 53423
rect -69970 53336 -69898 53428
rect -69821 53426 -36019 53431
rect -69821 53336 -46398 53426
rect -69970 53333 -46398 53336
rect -70129 53331 -46398 53333
rect -46321 53344 -36019 53426
rect -35942 53430 37954 53439
rect -35942 53427 37846 53430
rect -35942 53426 37697 53427
rect -35942 53344 -11207 53426
rect -46321 53331 -11207 53344
rect -11130 53419 24613 53426
rect -11130 53331 2897 53419
rect -70129 53328 2897 53331
rect -70936 53324 2897 53328
rect 2974 53331 24613 53419
rect 24690 53422 37697 53426
rect 24690 53331 37538 53422
rect 2974 53327 37538 53331
rect 37615 53332 37697 53422
rect 37774 53335 37846 53427
rect 37923 53335 37954 53430
rect 37774 53332 37954 53335
rect 37615 53327 37954 53332
rect 2974 53324 37954 53327
rect -70936 53280 37954 53324
rect -70936 53272 -36017 53280
rect -70936 53269 -69896 53272
rect -70936 53264 -70045 53269
rect -70936 53169 -70204 53264
rect -70127 53174 -70045 53264
rect -69968 53177 -69896 53269
rect -69819 53267 -36017 53272
rect -69819 53177 -46396 53267
rect -69968 53174 -46396 53177
rect -70127 53172 -46396 53174
rect -46319 53185 -36017 53267
rect -35940 53271 37954 53280
rect -35940 53268 37848 53271
rect -35940 53267 37699 53268
rect -35940 53185 -11205 53267
rect -46319 53172 -11205 53185
rect -11128 53260 24615 53267
rect -11128 53172 2899 53260
rect -70127 53169 2899 53172
rect -70936 53165 2899 53169
rect 2976 53172 24615 53260
rect 24692 53263 37699 53267
rect 24692 53172 37540 53263
rect 2976 53168 37540 53172
rect 37617 53173 37699 53263
rect 37776 53176 37848 53268
rect 37925 53176 37954 53271
rect 37776 53173 37954 53176
rect 37617 53168 37954 53173
rect 2976 53165 37954 53168
rect -70936 53122 37954 53165
rect -70936 53114 -36018 53122
rect -70936 53111 -69897 53114
rect -70936 53106 -70046 53111
rect -70936 53011 -70205 53106
rect -70128 53016 -70046 53106
rect -69969 53019 -69897 53111
rect -69820 53109 -36018 53114
rect -69820 53019 -46397 53109
rect -69969 53016 -46397 53019
rect -70128 53014 -46397 53016
rect -46320 53027 -36018 53109
rect -35941 53113 37954 53122
rect -35941 53110 37847 53113
rect -35941 53109 37698 53110
rect -35941 53027 -11206 53109
rect -46320 53014 -11206 53027
rect -11129 53102 24614 53109
rect -11129 53014 2898 53102
rect -70128 53011 2898 53014
rect -70936 53007 2898 53011
rect 2975 53014 24614 53102
rect 24691 53105 37698 53109
rect 24691 53014 37539 53105
rect 2975 53010 37539 53014
rect 37616 53015 37698 53105
rect 37775 53018 37847 53110
rect 37924 53018 37954 53113
rect 37775 53015 37954 53018
rect 37616 53010 37954 53015
rect 2975 53007 37954 53010
rect -70936 52988 37954 53007
rect -70936 52572 37954 52597
rect -70936 52559 -46599 52572
rect -70936 52556 -70591 52559
rect -70936 52551 -70740 52556
rect -70936 52456 -70899 52551
rect -70822 52461 -70740 52551
rect -70663 52464 -70591 52556
rect -70514 52477 -46599 52559
rect -46522 52563 37954 52572
rect -46522 52477 -36236 52563
rect -70514 52468 -36236 52477
rect -36159 52557 37954 52563
rect -36159 52556 24412 52557
rect -36159 52468 -11417 52556
rect -70514 52464 -11417 52468
rect -70663 52461 -11417 52464
rect -11340 52461 2693 52556
rect 2770 52462 24412 52556
rect 24489 52555 37954 52557
rect 24489 52552 37167 52555
rect 24489 52547 37018 52552
rect 24489 52462 36859 52547
rect 2770 52461 36859 52462
rect -70822 52456 36859 52461
rect -70936 52452 36859 52456
rect 36936 52457 37018 52547
rect 37095 52460 37167 52552
rect 37244 52460 37954 52555
rect 37095 52457 37954 52460
rect 36936 52452 37954 52457
rect -70936 52387 37954 52452
rect -70936 52383 -36239 52387
rect -70936 52380 -70594 52383
rect -70936 52375 -70743 52380
rect -70936 52280 -70902 52375
rect -70825 52285 -70743 52375
rect -70666 52288 -70594 52380
rect -70517 52369 -36239 52383
rect -70517 52288 -46600 52369
rect -70666 52285 -46600 52288
rect -70825 52280 -46600 52285
rect -70936 52274 -46600 52280
rect -46523 52292 -36239 52369
rect -36162 52381 37954 52387
rect -36162 52380 24409 52381
rect -36162 52292 -11420 52380
rect -46523 52285 -11420 52292
rect -11343 52285 2690 52380
rect 2767 52286 24409 52380
rect 24486 52379 37954 52381
rect 24486 52376 37164 52379
rect 24486 52371 37015 52376
rect 24486 52286 36856 52371
rect 2767 52285 36856 52286
rect -46523 52276 36856 52285
rect 36933 52281 37015 52371
rect 37092 52284 37164 52376
rect 37241 52284 37954 52379
rect 37092 52281 37954 52284
rect 36933 52276 37954 52281
rect -46523 52274 37954 52276
rect -70936 52228 37954 52274
rect -70936 52224 -36237 52228
rect -70936 52221 -70592 52224
rect -70936 52216 -70741 52221
rect -70936 52121 -70900 52216
rect -70823 52126 -70741 52216
rect -70664 52129 -70592 52221
rect -70515 52167 -36237 52224
rect -70515 52129 -46601 52167
rect -70664 52126 -46601 52129
rect -70823 52121 -46601 52126
rect -70936 52072 -46601 52121
rect -46524 52133 -36237 52167
rect -36160 52222 37954 52228
rect -36160 52221 24411 52222
rect -36160 52133 -11418 52221
rect -46524 52126 -11418 52133
rect -11341 52126 2692 52221
rect 2769 52127 24411 52221
rect 24488 52220 37954 52222
rect 24488 52217 37166 52220
rect 24488 52212 37017 52217
rect 24488 52127 36858 52212
rect 2769 52126 36858 52127
rect -46524 52117 36858 52126
rect 36935 52122 37017 52212
rect 37094 52125 37166 52217
rect 37243 52125 37954 52220
rect 37094 52122 37954 52125
rect 36935 52117 37954 52122
rect -46524 52072 37954 52117
rect -70936 52070 37954 52072
rect -70936 52066 -36238 52070
rect -70936 52063 -70593 52066
rect -70936 52058 -70742 52063
rect -70936 51963 -70901 52058
rect -70824 51968 -70742 52058
rect -70665 51971 -70593 52063
rect -70516 51975 -36238 52066
rect -36161 52064 37954 52070
rect -36161 52063 24410 52064
rect -36161 51975 -11419 52063
rect -70516 51971 -11419 51975
rect -70665 51968 -11419 51971
rect -11342 51968 2691 52063
rect 2768 51969 24410 52063
rect 24487 52062 37954 52064
rect 24487 52059 37165 52062
rect 24487 52054 37016 52059
rect 24487 51969 36857 52054
rect 2768 51968 36857 51969
rect -70824 51963 36857 51968
rect -70936 51959 36857 51963
rect 36934 51964 37016 52054
rect 37093 51967 37165 52059
rect 37242 51967 37954 52062
rect 37093 51964 37954 51967
rect 36934 51959 37954 51964
rect -70936 51951 37954 51959
rect -70915 51950 -70508 51951
rect 36839 51949 37251 51951
rect -53272 50091 -53149 50105
rect -53272 50012 -53252 50091
rect -53161 50062 -53149 50091
rect -53161 50012 -52841 50062
rect -53272 49970 -52841 50012
rect -32518 50028 -32331 50077
rect -42893 49984 -42770 49998
rect -42893 49970 -42873 49984
rect -53272 49939 -42873 49970
rect -53272 49860 -53256 49939
rect -53165 49905 -42873 49939
rect -42782 49970 -42770 49984
rect -32518 49970 -32478 50028
rect -42782 49929 -32478 49970
rect -32359 49970 -32331 50028
rect -3907 50004 -3784 50018
rect -17998 49970 -17875 49981
rect -3907 49970 -3887 50004
rect -32359 49967 -3887 49970
rect -32359 49929 -17978 49967
rect -42782 49905 -17978 49929
rect -53165 49888 -17978 49905
rect -17887 49925 -3887 49967
rect -3796 49925 -3784 50004
rect -17887 49888 -3784 49925
rect -53165 49860 -3784 49888
rect -53272 49852 -3784 49860
rect -53272 49848 -3891 49852
rect -53116 49832 -3891 49848
rect -53116 49784 -42877 49832
rect -42893 49753 -42877 49784
rect -42786 49815 -3891 49832
rect -42786 49806 -17982 49815
rect -42786 49784 -32484 49806
rect -42786 49753 -42770 49784
rect -42893 49741 -42770 49753
rect -32518 49707 -32484 49784
rect -32365 49784 -17982 49806
rect -32365 49707 -32331 49784
rect -17998 49736 -17982 49784
rect -17891 49784 -3891 49815
rect -17891 49736 -17875 49784
rect -3907 49773 -3891 49784
rect -3800 49773 -3784 49852
rect -3907 49761 -3784 49773
rect -17998 49724 -17875 49736
rect -32518 49685 -32331 49707
rect -70936 45232 37954 45266
rect -70936 45229 -69895 45232
rect -70936 45224 -70044 45229
rect -70936 45129 -70203 45224
rect -70126 45134 -70044 45224
rect -69967 45137 -69895 45229
rect -69818 45231 37954 45232
rect -69818 45228 -36083 45231
rect -69818 45137 -46389 45228
rect -69967 45134 -46389 45137
rect -70126 45133 -46389 45134
rect -46312 45136 -36083 45228
rect -36006 45136 -11035 45231
rect -10958 45136 13967 45231
rect 14044 45228 35592 45231
rect 14044 45136 24617 45228
rect -46312 45133 24617 45136
rect 24694 45136 35592 45228
rect 35669 45229 37954 45231
rect 35669 45226 37849 45229
rect 35669 45221 37700 45226
rect 35669 45136 37541 45221
rect 24694 45133 37541 45136
rect -70126 45129 37541 45133
rect -70936 45126 37541 45129
rect 37618 45131 37700 45221
rect 37777 45134 37849 45226
rect 37926 45134 37954 45229
rect 37777 45131 37954 45134
rect 37618 45126 37954 45131
rect -70936 45056 37954 45126
rect -70936 45053 -69898 45056
rect -70936 45048 -70047 45053
rect -70936 44953 -70206 45048
rect -70129 44958 -70047 45048
rect -69970 44961 -69898 45053
rect -69821 45055 37954 45056
rect -69821 45052 -36086 45055
rect -69821 44961 -46392 45052
rect -69970 44958 -46392 44961
rect -70129 44957 -46392 44958
rect -46315 44960 -36086 45052
rect -36009 44960 -11038 45055
rect -10961 44960 13964 45055
rect 14041 45052 35589 45055
rect 14041 44960 24614 45052
rect -46315 44957 24614 44960
rect 24691 44960 35589 45052
rect 35666 45053 37954 45055
rect 35666 45050 37846 45053
rect 35666 45045 37697 45050
rect 35666 44960 37538 45045
rect 24691 44957 37538 44960
rect -70129 44953 37538 44957
rect -70936 44950 37538 44953
rect 37615 44955 37697 45045
rect 37774 44958 37846 45050
rect 37923 44958 37954 45053
rect 37774 44955 37954 44958
rect 37615 44950 37954 44955
rect -70936 44897 37954 44950
rect -70936 44894 -69896 44897
rect -70936 44889 -70045 44894
rect -70936 44794 -70204 44889
rect -70127 44799 -70045 44889
rect -69968 44802 -69896 44894
rect -69819 44896 37954 44897
rect -69819 44893 -36084 44896
rect -69819 44802 -46390 44893
rect -69968 44799 -46390 44802
rect -70127 44798 -46390 44799
rect -46313 44801 -36084 44893
rect -36007 44801 -11036 44896
rect -10959 44801 13966 44896
rect 14043 44893 35591 44896
rect 14043 44801 24616 44893
rect -46313 44798 24616 44801
rect 24693 44801 35591 44893
rect 35668 44894 37954 44896
rect 35668 44891 37848 44894
rect 35668 44886 37699 44891
rect 35668 44801 37540 44886
rect 24693 44798 37540 44801
rect -70127 44794 37540 44798
rect -70936 44791 37540 44794
rect 37617 44796 37699 44886
rect 37776 44799 37848 44891
rect 37925 44799 37954 44894
rect 37776 44796 37954 44799
rect 37617 44791 37954 44796
rect -70936 44739 37954 44791
rect -70936 44736 -69897 44739
rect -70936 44731 -70046 44736
rect -70936 44636 -70205 44731
rect -70128 44641 -70046 44731
rect -69969 44644 -69897 44736
rect -69820 44738 37954 44739
rect -69820 44735 -36085 44738
rect -69820 44644 -46391 44735
rect -69969 44641 -46391 44644
rect -70128 44640 -46391 44641
rect -46314 44643 -36085 44735
rect -36008 44643 -11037 44738
rect -10960 44643 13965 44738
rect 14042 44735 35590 44738
rect 14042 44643 24615 44735
rect -46314 44640 24615 44643
rect 24692 44643 35590 44735
rect 35667 44736 37954 44738
rect 35667 44733 37847 44736
rect 35667 44728 37698 44733
rect 35667 44643 37539 44728
rect 24692 44640 37539 44643
rect -70128 44636 37539 44640
rect -70936 44633 37539 44636
rect 37616 44638 37698 44728
rect 37775 44641 37847 44733
rect 37924 44641 37954 44736
rect 37775 44638 37954 44641
rect 37616 44633 37954 44638
rect -70936 44620 37954 44633
rect -70936 44191 37954 44229
rect -70936 44189 -46592 44191
rect -70936 44186 -70587 44189
rect -70936 44181 -70736 44186
rect -70936 44086 -70895 44181
rect -70818 44091 -70736 44181
rect -70659 44094 -70587 44186
rect -70510 44096 -46592 44189
rect -46515 44188 35389 44191
rect -46515 44096 -36289 44188
rect -70510 44094 -36289 44096
rect -70659 44093 -36289 44094
rect -36212 44093 -11241 44188
rect -11164 44093 13767 44188
rect 13844 44093 24415 44188
rect 24492 44096 35389 44188
rect 35466 44186 37954 44191
rect 35466 44183 37163 44186
rect 35466 44178 37014 44183
rect 35466 44096 36855 44178
rect 24492 44093 36855 44096
rect -70659 44091 36855 44093
rect -70818 44086 36855 44091
rect -70936 44083 36855 44086
rect 36932 44088 37014 44178
rect 37091 44091 37163 44183
rect 37240 44091 37954 44186
rect 37091 44088 37954 44091
rect 36932 44083 37954 44088
rect -70936 44015 37954 44083
rect -70936 44013 -46595 44015
rect -70936 44010 -70590 44013
rect -70936 44005 -70739 44010
rect -70936 43910 -70898 44005
rect -70821 43915 -70739 44005
rect -70662 43918 -70590 44010
rect -70513 43920 -46595 44013
rect -46518 44012 35386 44015
rect -46518 43920 -36292 44012
rect -70513 43918 -36292 43920
rect -70662 43917 -36292 43918
rect -36215 43917 -11244 44012
rect -11167 43917 13764 44012
rect 13841 43917 24412 44012
rect 24489 43920 35386 44012
rect 35463 44010 37954 44015
rect 35463 44007 37160 44010
rect 35463 44002 37011 44007
rect 35463 43920 36852 44002
rect 24489 43917 36852 43920
rect -70662 43915 36852 43917
rect -70821 43910 36852 43915
rect -70936 43907 36852 43910
rect 36929 43912 37011 44002
rect 37088 43915 37160 44007
rect 37237 43915 37954 44010
rect 37088 43912 37954 43915
rect 36929 43907 37954 43912
rect -70936 43856 37954 43907
rect -70936 43854 -46593 43856
rect -70936 43851 -70588 43854
rect -70936 43846 -70737 43851
rect -70936 43751 -70896 43846
rect -70819 43756 -70737 43846
rect -70660 43759 -70588 43851
rect -70511 43761 -46593 43854
rect -46516 43853 35388 43856
rect -46516 43761 -36290 43853
rect -70511 43759 -36290 43761
rect -70660 43758 -36290 43759
rect -36213 43758 -11242 43853
rect -11165 43758 13766 43853
rect 13843 43758 24414 43853
rect 24491 43761 35388 43853
rect 35465 43851 37954 43856
rect 35465 43848 37162 43851
rect 35465 43843 37013 43848
rect 35465 43761 36854 43843
rect 24491 43758 36854 43761
rect -70660 43756 36854 43758
rect -70819 43751 36854 43756
rect -70936 43748 36854 43751
rect 36931 43753 37013 43843
rect 37090 43756 37162 43848
rect 37239 43756 37954 43851
rect 37090 43753 37954 43756
rect 36931 43748 37954 43753
rect -70936 43698 37954 43748
rect -70936 43696 -46594 43698
rect -70936 43693 -70589 43696
rect -70936 43688 -70738 43693
rect -70936 43593 -70897 43688
rect -70820 43598 -70738 43688
rect -70661 43601 -70589 43693
rect -70512 43603 -46594 43696
rect -46517 43695 35387 43698
rect -46517 43603 -36291 43695
rect -70512 43601 -36291 43603
rect -70661 43600 -36291 43601
rect -36214 43600 -11243 43695
rect -11166 43600 13765 43695
rect 13842 43600 24413 43695
rect 24490 43603 35387 43695
rect 35464 43693 37954 43698
rect 35464 43690 37161 43693
rect 35464 43685 37012 43690
rect 35464 43603 36853 43685
rect 24490 43600 36853 43603
rect -70661 43598 36853 43600
rect -70820 43593 36853 43598
rect -70936 43590 36853 43593
rect 36930 43595 37012 43685
rect 37089 43598 37161 43690
rect 37238 43598 37954 43693
rect 37089 43595 37954 43598
rect 36930 43590 37954 43595
rect -70936 43583 37954 43590
rect -70911 43580 -70504 43583
rect 36835 43580 37247 43583
rect -42874 41787 -42751 41801
rect -53195 41757 -53072 41771
rect -53195 41678 -53175 41757
rect -53084 41707 -53072 41757
rect -42874 41708 -42854 41787
rect -42763 41708 -42751 41787
rect -42874 41707 -42751 41708
rect -32499 41759 -32337 41790
rect -32499 41707 -32467 41759
rect -53084 41678 -32467 41707
rect -53195 41675 -32467 41678
rect -32362 41707 -32337 41759
rect -32362 41675 -17726 41707
rect -53195 41669 -17726 41675
rect 28791 41689 28914 41703
rect -53195 41655 -17702 41669
rect -53195 41635 -17805 41655
rect -53195 41605 -42858 41635
rect -53195 41526 -53179 41605
rect -53088 41556 -42858 41605
rect -42767 41576 -17805 41635
rect -17714 41576 -17702 41655
rect 28791 41610 28811 41689
rect 28902 41610 28914 41689
rect -42767 41568 -17702 41576
rect -42767 41556 -32472 41568
rect -53088 41547 -32472 41556
rect -53088 41526 -53072 41547
rect -42874 41544 -42751 41547
rect -53195 41514 -53072 41526
rect -32499 41484 -32472 41547
rect -32367 41547 -17702 41568
rect -32367 41484 -32337 41547
rect -32499 41461 -32337 41484
rect -17825 41503 -17702 41547
rect -17825 41424 -17809 41503
rect -17718 41424 -17702 41503
rect -17825 41412 -17702 41424
rect 17838 41565 17961 41579
rect 17838 41486 17858 41565
rect 17949 41545 17961 41565
rect 28791 41545 28914 41610
rect 17949 41537 28914 41545
rect 17949 41486 28807 41537
rect 17838 41458 28807 41486
rect 28898 41458 28914 41537
rect 17838 41413 28914 41458
rect 17838 41334 17854 41413
rect 17945 41364 28914 41413
rect 17945 41334 17961 41364
rect 17838 41322 17961 41334
rect -69427 41107 -69286 41132
rect -69427 41042 -69407 41107
rect -69346 41042 -69286 41107
rect -69427 40978 -69286 41042
rect -63615 40978 -63448 40988
rect -69427 40954 -63448 40978
rect -69427 40847 -63590 40954
rect -63479 40847 -63448 40954
rect -69427 40837 -63448 40847
rect -63615 40821 -63448 40837
rect 28461 39732 28584 39746
rect 16745 39643 16868 39657
rect 16745 39564 16765 39643
rect 16856 39609 16868 39643
rect 28461 39653 28481 39732
rect 28572 39653 28584 39732
rect 28461 39609 28584 39653
rect 16856 39580 28588 39609
rect 16856 39564 28477 39580
rect 16745 39501 28477 39564
rect 28568 39501 28588 39580
rect 16745 39491 28588 39501
rect 16745 39412 16761 39491
rect 16852 39418 28588 39491
rect 16852 39412 16868 39418
rect 16745 39400 16868 39412
rect -69535 39299 -69394 39328
rect -69535 39225 -69513 39299
rect -69434 39225 -69394 39299
rect -69535 39041 -69394 39225
rect -63128 39041 -62961 39051
rect -69535 39017 -62961 39041
rect -69535 38910 -63103 39017
rect -62992 38910 -62961 39017
rect -69535 38900 -62961 38910
rect -63128 38884 -62961 38900
rect -70936 37020 37954 37052
rect -70936 37015 -56569 37020
rect -70936 37012 -69895 37015
rect -70936 37007 -70044 37012
rect -70936 36912 -70203 37007
rect -70126 36917 -70044 37007
rect -69967 36920 -69895 37012
rect -69818 36925 -56569 37015
rect -56492 36925 -46396 37020
rect -46319 36925 -36023 37020
rect -35946 36925 -24963 37020
rect -24886 36925 -11137 37020
rect -11060 36925 2839 37020
rect 2916 36925 13806 37020
rect 13883 37016 37954 37020
rect 13883 36925 24704 37016
rect -69818 36921 24704 36925
rect 24781 36921 35612 37016
rect 35689 37006 37954 37016
rect 35689 37003 37849 37006
rect 35689 36998 37700 37003
rect 35689 36921 37541 36998
rect -69818 36920 37541 36921
rect -69967 36917 37541 36920
rect -70126 36912 37541 36917
rect -70936 36903 37541 36912
rect 37618 36908 37700 36998
rect 37777 36911 37849 37003
rect 37926 36911 37954 37006
rect 37777 36908 37954 36911
rect 37618 36903 37954 36908
rect -70936 36844 37954 36903
rect -70936 36839 -56572 36844
rect -70936 36836 -69898 36839
rect -70936 36831 -70047 36836
rect -70936 36736 -70206 36831
rect -70129 36741 -70047 36831
rect -69970 36744 -69898 36836
rect -69821 36749 -56572 36839
rect -56495 36749 -46399 36844
rect -46322 36749 -36026 36844
rect -35949 36749 -24966 36844
rect -24889 36749 -11140 36844
rect -11063 36749 2836 36844
rect 2913 36749 13803 36844
rect 13880 36840 37954 36844
rect 13880 36749 24701 36840
rect -69821 36745 24701 36749
rect 24778 36745 35609 36840
rect 35686 36830 37954 36840
rect 35686 36827 37846 36830
rect 35686 36822 37697 36827
rect 35686 36745 37538 36822
rect -69821 36744 37538 36745
rect -69970 36741 37538 36744
rect -70129 36736 37538 36741
rect -70936 36727 37538 36736
rect 37615 36732 37697 36822
rect 37774 36735 37846 36827
rect 37923 36735 37954 36830
rect 37774 36732 37954 36735
rect 37615 36727 37954 36732
rect -70936 36685 37954 36727
rect -70936 36680 -56570 36685
rect -70936 36677 -69896 36680
rect -70936 36672 -70045 36677
rect -70936 36577 -70204 36672
rect -70127 36582 -70045 36672
rect -69968 36585 -69896 36677
rect -69819 36590 -56570 36680
rect -56493 36590 -46397 36685
rect -46320 36590 -36024 36685
rect -35947 36590 -24964 36685
rect -24887 36590 -11138 36685
rect -11061 36590 2838 36685
rect 2915 36590 13805 36685
rect 13882 36681 37954 36685
rect 13882 36590 24703 36681
rect -69819 36586 24703 36590
rect 24780 36586 35611 36681
rect 35688 36671 37954 36681
rect 35688 36668 37848 36671
rect 35688 36663 37699 36668
rect 35688 36586 37540 36663
rect -69819 36585 37540 36586
rect -69968 36582 37540 36585
rect -70127 36577 37540 36582
rect -70936 36568 37540 36577
rect 37617 36573 37699 36663
rect 37776 36576 37848 36668
rect 37925 36576 37954 36671
rect 37776 36573 37954 36576
rect 37617 36568 37954 36573
rect -70936 36527 37954 36568
rect -70936 36522 -56571 36527
rect -70936 36519 -69897 36522
rect -70936 36514 -70046 36519
rect -70936 36419 -70205 36514
rect -70128 36424 -70046 36514
rect -69969 36427 -69897 36519
rect -69820 36432 -56571 36522
rect -56494 36432 -46398 36527
rect -46321 36432 -36025 36527
rect -35948 36432 -24965 36527
rect -24888 36432 -11139 36527
rect -11062 36432 2837 36527
rect 2914 36432 13804 36527
rect 13881 36523 37954 36527
rect 13881 36432 24702 36523
rect -69820 36428 24702 36432
rect 24779 36428 35610 36523
rect 35687 36513 37954 36523
rect 35687 36510 37847 36513
rect 35687 36505 37698 36510
rect 35687 36428 37539 36505
rect -69820 36427 37539 36428
rect -69969 36424 37539 36427
rect -70128 36419 37539 36424
rect -70936 36410 37539 36419
rect 37616 36415 37698 36505
rect 37775 36418 37847 36510
rect 37924 36418 37954 36513
rect 37775 36415 37954 36418
rect 37616 36410 37954 36415
rect -70936 36406 37954 36410
rect 37521 36400 37933 36406
rect -70936 35770 37954 35800
rect -70936 35766 -11338 35770
rect -70936 35764 -36221 35766
rect -70936 35761 -70583 35764
rect -70936 35756 -70732 35761
rect -70936 35661 -70891 35756
rect -70814 35666 -70732 35756
rect -70655 35669 -70583 35761
rect -70506 35763 -36221 35764
rect -70506 35669 -56777 35763
rect -70655 35668 -56777 35669
rect -56700 35668 -46601 35763
rect -46524 35671 -36221 35763
rect -36144 35760 -11338 35766
rect -36144 35671 -25161 35760
rect -46524 35668 -25161 35671
rect -70655 35666 -25161 35668
rect -70814 35665 -25161 35666
rect -25084 35675 -11338 35760
rect -11261 35766 37954 35770
rect -11261 35760 24503 35766
rect -11261 35675 2631 35760
rect -25084 35665 2631 35675
rect 2708 35665 13601 35760
rect 13678 35671 24503 35760
rect 24580 35760 37954 35766
rect 24580 35671 35407 35760
rect 13678 35665 35407 35671
rect 35484 35759 37954 35760
rect 35484 35756 37159 35759
rect 35484 35751 37010 35756
rect 35484 35665 36851 35751
rect -70814 35661 36851 35665
rect -70936 35656 36851 35661
rect 36928 35661 37010 35751
rect 37087 35664 37159 35756
rect 37236 35664 37954 35759
rect 37087 35661 37954 35664
rect 36928 35656 37954 35661
rect -70936 35594 37954 35656
rect -70936 35590 -11341 35594
rect -70936 35588 -36224 35590
rect -70936 35585 -70586 35588
rect -70936 35580 -70735 35585
rect -70936 35485 -70894 35580
rect -70817 35490 -70735 35580
rect -70658 35493 -70586 35585
rect -70509 35587 -36224 35588
rect -70509 35493 -56780 35587
rect -70658 35492 -56780 35493
rect -56703 35492 -46604 35587
rect -46527 35495 -36224 35587
rect -36147 35584 -11341 35590
rect -36147 35495 -25164 35584
rect -46527 35492 -25164 35495
rect -70658 35490 -25164 35492
rect -70817 35489 -25164 35490
rect -25087 35499 -11341 35584
rect -11264 35590 37954 35594
rect -11264 35584 24500 35590
rect -11264 35499 2628 35584
rect -25087 35489 2628 35499
rect 2705 35489 13598 35584
rect 13675 35495 24500 35584
rect 24577 35584 37954 35590
rect 24577 35495 35404 35584
rect 13675 35489 35404 35495
rect 35481 35583 37954 35584
rect 35481 35580 37156 35583
rect 35481 35575 37007 35580
rect 35481 35489 36848 35575
rect -70817 35485 36848 35489
rect -70936 35480 36848 35485
rect 36925 35485 37007 35575
rect 37084 35488 37156 35580
rect 37233 35488 37954 35583
rect 37084 35485 37954 35488
rect 36925 35480 37954 35485
rect -70936 35435 37954 35480
rect -70936 35431 -11339 35435
rect -70936 35429 -36222 35431
rect -70936 35426 -70584 35429
rect -70936 35421 -70733 35426
rect -70936 35326 -70892 35421
rect -70815 35331 -70733 35421
rect -70656 35334 -70584 35426
rect -70507 35428 -36222 35429
rect -70507 35334 -56778 35428
rect -70656 35333 -56778 35334
rect -56701 35333 -46602 35428
rect -46525 35336 -36222 35428
rect -36145 35425 -11339 35431
rect -36145 35336 -25162 35425
rect -46525 35333 -25162 35336
rect -70656 35331 -25162 35333
rect -70815 35330 -25162 35331
rect -25085 35340 -11339 35425
rect -11262 35431 37954 35435
rect -11262 35425 24502 35431
rect -11262 35340 2630 35425
rect -25085 35330 2630 35340
rect 2707 35330 13600 35425
rect 13677 35336 24502 35425
rect 24579 35425 37954 35431
rect 24579 35336 35406 35425
rect 13677 35330 35406 35336
rect 35483 35424 37954 35425
rect 35483 35421 37158 35424
rect 35483 35416 37009 35421
rect 35483 35330 36850 35416
rect -70815 35326 36850 35330
rect -70936 35321 36850 35326
rect 36927 35326 37009 35416
rect 37086 35329 37158 35421
rect 37235 35329 37954 35424
rect 37086 35326 37954 35329
rect 36927 35321 37954 35326
rect -70936 35277 37954 35321
rect -70936 35273 -11340 35277
rect -70936 35271 -36223 35273
rect -70936 35268 -70585 35271
rect -70936 35263 -70734 35268
rect -70936 35168 -70893 35263
rect -70816 35173 -70734 35263
rect -70657 35176 -70585 35268
rect -70508 35270 -36223 35271
rect -70508 35176 -56779 35270
rect -70657 35175 -56779 35176
rect -56702 35175 -46603 35270
rect -46526 35178 -36223 35270
rect -36146 35267 -11340 35273
rect -36146 35178 -25163 35267
rect -46526 35175 -25163 35178
rect -70657 35173 -25163 35175
rect -70816 35172 -25163 35173
rect -25086 35182 -11340 35267
rect -11263 35273 37954 35277
rect -11263 35267 24501 35273
rect -11263 35182 2629 35267
rect -25086 35172 2629 35182
rect 2706 35172 13599 35267
rect 13676 35178 24501 35267
rect 24578 35267 37954 35273
rect 24578 35178 35405 35267
rect 13676 35172 35405 35178
rect 35482 35266 37954 35267
rect 35482 35263 37157 35266
rect 35482 35258 37008 35263
rect 35482 35172 36849 35258
rect -70816 35168 36849 35172
rect -70936 35163 36849 35168
rect 36926 35168 37008 35258
rect 37085 35171 37157 35263
rect 37234 35171 37954 35266
rect 37085 35168 37954 35171
rect 36926 35163 37954 35168
rect -70936 35154 37954 35163
rect 36831 35153 37243 35154
rect -63376 33288 -63253 33302
rect -63376 33209 -63356 33288
rect -63265 33269 -63253 33288
rect -53204 33293 -53081 33307
rect -53204 33269 -53184 33293
rect -63265 33214 -53184 33269
rect -53093 33269 -53081 33293
rect -42810 33269 -42687 33278
rect -19314 33269 -19162 33285
rect -53093 33264 7121 33269
rect -53093 33214 -42790 33264
rect -63265 33209 -42790 33214
rect -63376 33185 -42790 33209
rect -42699 33244 7121 33264
rect -42699 33185 -19287 33244
rect -63376 33156 -19287 33185
rect -19196 33206 7121 33244
rect -19196 33195 7125 33206
rect -19196 33156 -3954 33195
rect -63376 33150 -3954 33156
rect -63376 33141 -17916 33150
rect -63376 33136 -53188 33141
rect -63376 33057 -63360 33136
rect -63269 33080 -53188 33136
rect -63269 33057 -63253 33080
rect -63376 33045 -63253 33057
rect -53204 33062 -53188 33080
rect -53097 33112 -17916 33141
rect -53097 33080 -42794 33112
rect -53097 33062 -53081 33080
rect -53204 33050 -53081 33062
rect -42810 33033 -42794 33080
rect -42703 33108 -17916 33112
rect -42703 33080 -31731 33108
rect -42703 33033 -42687 33080
rect -42810 33021 -42687 33033
rect -31751 33029 -31731 33080
rect -31640 33080 -17916 33108
rect -31640 33029 -31628 33080
rect -31751 32956 -31628 33029
rect -31751 32877 -31735 32956
rect -31644 32877 -31628 32956
rect -19314 33037 -19162 33080
rect -19314 32949 -19284 33037
rect -19193 32949 -19162 33037
rect -19314 32922 -19162 32949
rect -17936 33071 -17916 33080
rect -17825 33116 -3954 33150
rect -3863 33192 7125 33195
rect -3863 33116 7022 33192
rect -17825 33113 7022 33116
rect 7113 33113 7125 33192
rect -17825 33080 7125 33113
rect -17825 33071 -17813 33080
rect -17936 32998 -17813 33071
rect -17936 32919 -17920 32998
rect -17829 32919 -17813 32998
rect -3974 33043 -3851 33080
rect -3974 32964 -3958 33043
rect -3867 32964 -3851 33043
rect -3974 32952 -3851 32964
rect 7002 33040 7125 33080
rect 7002 32961 7018 33040
rect 7109 32961 7125 33040
rect 7002 32949 7125 32961
rect 17889 33195 18012 33209
rect 17889 33116 17909 33195
rect 18000 33152 18012 33195
rect 28805 33195 28928 33209
rect 28805 33152 28825 33195
rect 18000 33116 28825 33152
rect 28916 33116 28928 33195
rect 17889 33043 28928 33116
rect 17889 32964 17905 33043
rect 17996 32982 28821 33043
rect 17996 32964 18012 32982
rect 17889 32952 18012 32964
rect 28805 32964 28821 32982
rect 28912 32964 28928 33043
rect 28805 32952 28928 32964
rect -17936 32907 -17813 32919
rect -31751 32865 -31628 32877
rect -63789 31350 -63666 31364
rect -63789 31323 -63769 31350
rect -68364 31271 -63769 31323
rect -63678 31323 -63666 31350
rect -53503 31350 -53380 31364
rect -53503 31323 -53483 31350
rect -63678 31271 -53483 31323
rect -53392 31323 -53380 31350
rect -43129 31323 -43006 31333
rect -53392 31319 6848 31323
rect -53392 31271 -43109 31319
rect -68364 31240 -43109 31271
rect -43018 31240 6848 31319
rect -68364 31225 6848 31240
rect -68364 31198 -4250 31225
rect -68364 31187 -63773 31198
rect -68364 31130 -68318 31187
rect -68237 31131 -63773 31187
rect -68237 31130 -68172 31131
rect -68364 31016 -68172 31130
rect -63789 31119 -63773 31131
rect -63682 31131 -53487 31198
rect -63682 31119 -63666 31131
rect -63789 31107 -63666 31119
rect -53503 31119 -53487 31131
rect -53396 31174 -4250 31198
rect -53396 31167 -18207 31174
rect -53396 31131 -43113 31167
rect -53396 31119 -53380 31131
rect -53503 31107 -53380 31119
rect -43129 31088 -43113 31131
rect -43022 31134 -18207 31167
rect -43022 31131 -32035 31134
rect -43022 31088 -43006 31131
rect -43129 31076 -43006 31088
rect -32055 31055 -32035 31131
rect -31944 31131 -18207 31134
rect -31944 31055 -31932 31131
rect -32055 30982 -31932 31055
rect -32055 30903 -32039 30982
rect -31948 30903 -31932 30982
rect -18227 31095 -18207 31131
rect -18116 31146 -4250 31174
rect -4159 31174 6848 31225
rect -4159 31146 6710 31174
rect -18116 31131 6710 31146
rect -18116 31095 -18104 31131
rect -18227 31022 -18104 31095
rect -18227 30943 -18211 31022
rect -18120 30943 -18104 31022
rect -4270 31073 -4147 31131
rect -4270 30994 -4254 31073
rect -4163 30994 -4147 31073
rect -4270 30982 -4147 30994
rect 6656 31095 6710 31131
rect 6801 31095 6848 31174
rect 28530 31229 28653 31243
rect 28530 31150 28550 31229
rect 28641 31150 28653 31229
rect 6656 31022 6848 31095
rect -18227 30931 -18104 30943
rect 6656 30943 6706 31022
rect 6797 30943 6848 31022
rect 6656 30929 6848 30943
rect 17160 31119 17283 31133
rect 17160 31040 17180 31119
rect 17271 31083 17283 31119
rect 28530 31083 28653 31150
rect 17271 31077 28658 31083
rect 17271 31040 28546 31077
rect 17160 30998 28546 31040
rect 28637 30998 28658 31077
rect 17160 30967 28658 30998
rect -32055 30891 -31932 30903
rect 17160 30888 17176 30967
rect 17267 30900 28658 30967
rect 17267 30888 17283 30900
rect 17160 30876 17283 30888
rect -70936 28459 37954 28492
rect -70936 28458 -36223 28459
rect -70936 28455 -69899 28458
rect -70936 28450 -70048 28455
rect -70936 28355 -70207 28450
rect -70130 28360 -70048 28450
rect -69971 28363 -69899 28455
rect -69822 28364 -36223 28458
rect -36146 28456 13845 28459
rect -36146 28364 -11847 28456
rect -69822 28363 -11847 28364
rect -69971 28361 -11847 28363
rect -11770 28364 13845 28456
rect 13922 28449 37954 28459
rect 13922 28446 37853 28449
rect 13922 28441 37704 28446
rect 13922 28364 37545 28441
rect -11770 28361 37545 28364
rect -69971 28360 37545 28361
rect -70130 28355 37545 28360
rect -70936 28346 37545 28355
rect 37622 28351 37704 28441
rect 37781 28354 37853 28446
rect 37930 28354 37954 28449
rect 37781 28351 37954 28354
rect 37622 28346 37954 28351
rect -70936 28283 37954 28346
rect -70936 28282 -36226 28283
rect -70936 28279 -69902 28282
rect -70936 28274 -70051 28279
rect -70936 28179 -70210 28274
rect -70133 28184 -70051 28274
rect -69974 28187 -69902 28279
rect -69825 28188 -36226 28282
rect -36149 28280 13842 28283
rect -36149 28188 -11850 28280
rect -69825 28187 -11850 28188
rect -69974 28185 -11850 28187
rect -11773 28188 13842 28280
rect 13919 28273 37954 28283
rect 13919 28270 37850 28273
rect 13919 28265 37701 28270
rect 13919 28188 37542 28265
rect -11773 28185 37542 28188
rect -69974 28184 37542 28185
rect -70133 28179 37542 28184
rect -70936 28170 37542 28179
rect 37619 28175 37701 28265
rect 37778 28178 37850 28270
rect 37927 28178 37954 28273
rect 37778 28175 37954 28178
rect 37619 28170 37954 28175
rect -70936 28124 37954 28170
rect -70936 28123 -36224 28124
rect -70936 28120 -69900 28123
rect -70936 28115 -70049 28120
rect -70936 28020 -70208 28115
rect -70131 28025 -70049 28115
rect -69972 28028 -69900 28120
rect -69823 28029 -36224 28123
rect -36147 28121 13844 28124
rect -36147 28029 -11848 28121
rect -69823 28028 -11848 28029
rect -69972 28026 -11848 28028
rect -11771 28029 13844 28121
rect 13921 28114 37954 28124
rect 13921 28111 37852 28114
rect 13921 28106 37703 28111
rect 13921 28029 37544 28106
rect -11771 28026 37544 28029
rect -69972 28025 37544 28026
rect -70131 28020 37544 28025
rect -70936 28011 37544 28020
rect 37621 28016 37703 28106
rect 37780 28019 37852 28111
rect 37929 28019 37954 28114
rect 37780 28016 37954 28019
rect 37621 28011 37954 28016
rect -70936 27966 37954 28011
rect -70936 27965 -36225 27966
rect -70936 27962 -69901 27965
rect -70936 27957 -70050 27962
rect -70936 27862 -70209 27957
rect -70132 27867 -70050 27957
rect -69973 27870 -69901 27962
rect -69824 27871 -36225 27965
rect -36148 27963 13843 27966
rect -36148 27871 -11849 27963
rect -69824 27870 -11849 27871
rect -69973 27868 -11849 27870
rect -11772 27871 13843 27963
rect 13920 27956 37954 27966
rect 13920 27953 37851 27956
rect 13920 27948 37702 27953
rect 13920 27871 37543 27948
rect -11772 27868 37543 27871
rect -69973 27867 37543 27868
rect -70132 27862 37543 27867
rect -70936 27853 37543 27862
rect 37620 27858 37702 27948
rect 37779 27861 37851 27953
rect 37928 27861 37954 27956
rect 37779 27858 37954 27861
rect 37620 27853 37954 27858
rect -70936 27846 37954 27853
rect 37525 27843 37937 27846
rect -70936 27358 37954 27388
rect -70936 27348 -12047 27358
rect -70936 27345 -70583 27348
rect -70936 27340 -70732 27345
rect -70936 27245 -70891 27340
rect -70814 27250 -70732 27340
rect -70655 27253 -70583 27345
rect -70506 27344 -12047 27348
rect -70506 27253 -36430 27344
rect -70655 27250 -36430 27253
rect -70814 27249 -36430 27250
rect -36353 27263 -12047 27344
rect -11970 27351 37954 27358
rect -11970 27348 37159 27351
rect -11970 27263 13645 27348
rect -36353 27253 13645 27263
rect 13722 27343 37010 27348
rect 13722 27253 36851 27343
rect -36353 27249 36851 27253
rect -70814 27248 36851 27249
rect 36928 27253 37010 27343
rect 37087 27256 37159 27348
rect 37236 27256 37954 27351
rect 37087 27253 37954 27256
rect 36928 27248 37954 27253
rect -70814 27245 37954 27248
rect -70936 27182 37954 27245
rect -70936 27172 -12050 27182
rect -70936 27169 -70586 27172
rect -70936 27164 -70735 27169
rect -70936 27069 -70894 27164
rect -70817 27074 -70735 27164
rect -70658 27077 -70586 27169
rect -70509 27168 -12050 27172
rect -70509 27077 -36433 27168
rect -70658 27074 -36433 27077
rect -70817 27073 -36433 27074
rect -36356 27087 -12050 27168
rect -11973 27175 37954 27182
rect -11973 27172 37156 27175
rect -11973 27087 13642 27172
rect -36356 27077 13642 27087
rect 13719 27167 37007 27172
rect 13719 27077 36848 27167
rect -36356 27073 36848 27077
rect -70817 27072 36848 27073
rect 36925 27077 37007 27167
rect 37084 27080 37156 27172
rect 37233 27080 37954 27175
rect 37084 27077 37954 27080
rect 36925 27072 37954 27077
rect -70817 27069 37954 27072
rect -70936 27023 37954 27069
rect -70936 27013 -12048 27023
rect -70936 27010 -70584 27013
rect -70936 27005 -70733 27010
rect -70936 26910 -70892 27005
rect -70815 26915 -70733 27005
rect -70656 26918 -70584 27010
rect -70507 27009 -12048 27013
rect -70507 26918 -36431 27009
rect -70656 26915 -36431 26918
rect -70815 26914 -36431 26915
rect -36354 26928 -12048 27009
rect -11971 27016 37954 27023
rect -11971 27013 37158 27016
rect -11971 26928 13644 27013
rect -36354 26918 13644 26928
rect 13721 27008 37009 27013
rect 13721 26918 36850 27008
rect -36354 26914 36850 26918
rect -70815 26913 36850 26914
rect 36927 26918 37009 27008
rect 37086 26921 37158 27013
rect 37235 26921 37954 27016
rect 37086 26918 37954 26921
rect 36927 26913 37954 26918
rect -70815 26910 37954 26913
rect -70936 26865 37954 26910
rect -70936 26855 -12049 26865
rect -70936 26852 -70585 26855
rect -70936 26847 -70734 26852
rect -70936 26752 -70893 26847
rect -70816 26757 -70734 26847
rect -70657 26760 -70585 26852
rect -70508 26851 -12049 26855
rect -70508 26760 -36432 26851
rect -70657 26757 -36432 26760
rect -70816 26756 -36432 26757
rect -36355 26770 -12049 26851
rect -11972 26858 37954 26865
rect -11972 26855 37157 26858
rect -11972 26770 13643 26855
rect -36355 26760 13643 26770
rect 13720 26850 37008 26855
rect 13720 26760 36849 26850
rect -36355 26756 36849 26760
rect -70816 26755 36849 26756
rect 36926 26760 37008 26850
rect 37085 26763 37157 26855
rect 37234 26763 37954 26858
rect 37085 26760 37954 26763
rect 36926 26755 37954 26760
rect -70816 26752 37954 26755
rect -70936 26742 37954 26752
rect -70907 26739 -70500 26742
rect 16780 25377 16973 25378
rect 16780 25337 16974 25377
rect 16780 25231 16819 25337
rect 16940 25231 16974 25337
rect 16780 25176 16974 25231
rect 6986 25142 16974 25176
rect 6986 25063 7059 25142
rect 7150 25117 16974 25142
rect 7150 25063 16814 25117
rect 6986 25011 16814 25063
rect 16935 25011 16974 25117
rect -8429 24913 -8229 25001
rect -18635 24891 -18512 24905
rect -43024 24853 -42901 24867
rect -43024 24774 -43004 24853
rect -42913 24824 -42901 24853
rect -18635 24824 -18615 24891
rect -42913 24812 -18615 24824
rect -18524 24824 -18512 24891
rect -8429 24824 -8395 24913
rect -18524 24812 -8395 24824
rect -42913 24801 -8395 24812
rect -8259 24824 -8229 24913
rect 6986 24990 16974 25011
rect 6986 24911 7055 24990
rect 7146 24983 16974 24990
rect 7146 24911 7179 24983
rect 16780 24982 16973 24983
rect 6986 24824 7179 24911
rect -8259 24801 7179 24824
rect -42913 24774 7179 24801
rect -43024 24739 7179 24774
rect -43024 24701 -18619 24739
rect -43024 24622 -43008 24701
rect -42917 24660 -18619 24701
rect -18528 24660 7179 24739
rect -42917 24643 7179 24660
rect -42917 24631 -8407 24643
rect -42917 24622 -42901 24631
rect -43024 24610 -42901 24622
rect -8429 24531 -8407 24631
rect -8271 24631 7179 24643
rect -8271 24531 -8229 24631
rect -8429 24503 -8229 24531
rect 16872 23252 17065 23299
rect 6708 23211 6831 23225
rect 6708 23139 6728 23211
rect 6135 23132 6728 23139
rect 6819 23139 6831 23211
rect 16872 23144 16922 23252
rect 17027 23144 17065 23252
rect 16872 23139 17065 23144
rect 6819 23132 17065 23139
rect 6135 23059 17065 23132
rect 6135 22980 6724 23059
rect 6815 23039 17065 23059
rect 6815 22980 16914 23039
rect -19049 22965 -18926 22979
rect -43323 22913 -43200 22927
rect -43323 22878 -43303 22913
rect -68369 22834 -43303 22878
rect -43212 22878 -43200 22913
rect -19049 22886 -19029 22965
rect -18938 22886 -18926 22965
rect -19049 22878 -18926 22886
rect 6135 22948 16914 22980
rect 6135 22878 6326 22948
rect 16872 22931 16914 22948
rect 17019 22931 17065 23039
rect 16872 22899 17065 22931
rect -43212 22834 6326 22878
rect -68369 22813 6326 22834
rect -68369 22803 -19033 22813
rect -68369 22714 -68348 22803
rect -68263 22761 -19033 22803
rect -68263 22714 -43307 22761
rect -68369 22687 -43307 22714
rect -43323 22682 -43307 22687
rect -43216 22734 -19033 22761
rect -18942 22734 6326 22813
rect -43216 22687 6326 22734
rect -43216 22682 -43200 22687
rect -43323 22670 -43200 22682
rect -36212 19435 -36111 19442
rect -25841 19435 -25740 19439
rect -21233 19435 -21128 19437
rect 2994 19435 3095 19442
rect 13643 19435 13744 19439
rect 24703 19435 24804 19442
rect 35605 19435 35706 19442
rect -70936 19416 37954 19435
rect -70936 19409 -36194 19416
rect -70936 19400 -56557 19409
rect -70936 19397 -69895 19400
rect -70936 19392 -70044 19397
rect -70936 19297 -70203 19392
rect -70126 19302 -70044 19392
rect -69967 19305 -69895 19397
rect -69818 19314 -56557 19400
rect -56480 19314 -46406 19409
rect -46329 19321 -36194 19409
rect -36117 19415 3012 19416
rect -36117 19413 -21211 19415
rect -36117 19321 -25823 19413
rect -46329 19318 -25823 19321
rect -25746 19320 -21211 19413
rect -21134 19321 3012 19415
rect 3089 19413 24721 19416
rect 3089 19321 13661 19413
rect -21134 19320 13661 19321
rect -25746 19318 13661 19320
rect 13738 19321 24721 19413
rect 24798 19321 35623 19416
rect 35700 19398 37954 19416
rect 35700 19395 37849 19398
rect 35700 19390 37700 19395
rect 35700 19321 37541 19390
rect 13738 19318 37541 19321
rect -46329 19314 37541 19318
rect -69818 19305 37541 19314
rect -69967 19302 37541 19305
rect -70126 19297 37541 19302
rect -70936 19295 37541 19297
rect 37618 19300 37700 19390
rect 37777 19303 37849 19395
rect 37926 19303 37954 19398
rect 37777 19300 37954 19303
rect 37618 19295 37954 19300
rect -70936 19240 37954 19295
rect -70936 19233 -36197 19240
rect -70936 19224 -56560 19233
rect -70936 19221 -69898 19224
rect -70936 19216 -70047 19221
rect -70936 19121 -70206 19216
rect -70129 19126 -70047 19216
rect -69970 19129 -69898 19221
rect -69821 19138 -56560 19224
rect -56483 19138 -46409 19233
rect -46332 19145 -36197 19233
rect -36120 19239 3009 19240
rect -36120 19237 -21214 19239
rect -36120 19145 -25826 19237
rect -46332 19142 -25826 19145
rect -25749 19144 -21214 19237
rect -21137 19145 3009 19239
rect 3086 19237 24718 19240
rect 3086 19145 13658 19237
rect -21137 19144 13658 19145
rect -25749 19142 13658 19144
rect 13735 19145 24718 19237
rect 24795 19145 35620 19240
rect 35697 19222 37954 19240
rect 35697 19219 37846 19222
rect 35697 19214 37697 19219
rect 35697 19145 37538 19214
rect 13735 19142 37538 19145
rect -46332 19138 37538 19142
rect -69821 19129 37538 19138
rect -69970 19126 37538 19129
rect -70129 19121 37538 19126
rect -70936 19119 37538 19121
rect 37615 19124 37697 19214
rect 37774 19127 37846 19219
rect 37923 19127 37954 19222
rect 37774 19124 37954 19127
rect 37615 19119 37954 19124
rect -70936 19081 37954 19119
rect -70936 19074 -36195 19081
rect -70936 19065 -56558 19074
rect -70936 19062 -69896 19065
rect -70936 19057 -70045 19062
rect -70936 18962 -70204 19057
rect -70127 18967 -70045 19057
rect -69968 18970 -69896 19062
rect -69819 18979 -56558 19065
rect -56481 18979 -46407 19074
rect -46330 18986 -36195 19074
rect -36118 19080 3011 19081
rect -36118 19078 -21212 19080
rect -36118 18986 -25824 19078
rect -46330 18983 -25824 18986
rect -25747 18985 -21212 19078
rect -21135 18986 3011 19080
rect 3088 19078 24720 19081
rect 3088 18986 13660 19078
rect -21135 18985 13660 18986
rect -25747 18983 13660 18985
rect 13737 18986 24720 19078
rect 24797 18986 35622 19081
rect 35699 19063 37954 19081
rect 35699 19060 37848 19063
rect 35699 19055 37699 19060
rect 35699 18986 37540 19055
rect 13737 18983 37540 18986
rect -46330 18979 37540 18983
rect -69819 18970 37540 18979
rect -69968 18967 37540 18970
rect -70127 18962 37540 18967
rect -70936 18960 37540 18962
rect 37617 18965 37699 19055
rect 37776 18968 37848 19060
rect 37925 18968 37954 19063
rect 37776 18965 37954 18968
rect 37617 18960 37954 18965
rect -70936 18923 37954 18960
rect -70936 18916 -36196 18923
rect -70936 18907 -56559 18916
rect -70936 18904 -69897 18907
rect -70936 18899 -70046 18904
rect -70936 18804 -70205 18899
rect -70128 18809 -70046 18899
rect -69969 18812 -69897 18904
rect -69820 18821 -56559 18907
rect -56482 18821 -46408 18916
rect -46331 18828 -36196 18916
rect -36119 18922 3010 18923
rect -36119 18920 -21213 18922
rect -36119 18828 -25825 18920
rect -46331 18825 -25825 18828
rect -25748 18827 -21213 18920
rect -21136 18828 3010 18922
rect 3087 18920 24719 18923
rect 3087 18828 13659 18920
rect -21136 18827 13659 18828
rect -25748 18825 13659 18827
rect 13736 18828 24719 18920
rect 24796 18828 35621 18923
rect 35698 18905 37954 18923
rect 35698 18902 37847 18905
rect 35698 18897 37698 18902
rect 35698 18828 37539 18897
rect 13736 18825 37539 18828
rect -46331 18821 37539 18825
rect -69820 18812 37539 18821
rect -69969 18809 37539 18812
rect -70128 18804 37539 18809
rect -70936 18802 37539 18804
rect 37616 18807 37698 18897
rect 37775 18810 37847 18902
rect 37924 18810 37954 18905
rect 37775 18807 37954 18810
rect 37616 18802 37954 18807
rect -70936 18789 37954 18802
rect -20750 18354 -20645 18368
rect 2792 18354 2893 18359
rect 13437 18354 13538 18363
rect 24498 18354 24599 18356
rect -70936 18346 37954 18354
rect -70936 18326 -20728 18346
rect -70936 18319 -56752 18326
rect -70936 18316 -70587 18319
rect -70936 18311 -70736 18316
rect -70936 18216 -70895 18311
rect -70818 18221 -70736 18311
rect -70659 18224 -70587 18316
rect -70510 18231 -56752 18319
rect -56675 18322 -36400 18326
rect -56675 18231 -46605 18322
rect -70510 18227 -46605 18231
rect -46528 18231 -36400 18322
rect -36323 18231 -26029 18326
rect -25952 18251 -20728 18326
rect -20651 18337 37954 18346
rect -20651 18333 13455 18337
rect -20651 18251 2810 18333
rect -25952 18238 2810 18251
rect 2887 18242 13455 18333
rect 13532 18330 37954 18337
rect 13532 18242 24516 18330
rect 2887 18238 24516 18242
rect -25952 18235 24516 18238
rect 24593 18326 37954 18330
rect 24593 18235 35417 18326
rect -25952 18231 35417 18235
rect 35494 18316 37954 18326
rect 35494 18313 37163 18316
rect 35494 18308 37014 18313
rect 35494 18231 36855 18308
rect -46528 18227 36855 18231
rect -70510 18224 36855 18227
rect -70659 18221 36855 18224
rect -70818 18216 36855 18221
rect -70936 18213 36855 18216
rect 36932 18218 37014 18308
rect 37091 18221 37163 18313
rect 37240 18221 37954 18316
rect 37091 18218 37954 18221
rect 36932 18213 37954 18218
rect -70936 18170 37954 18213
rect -70936 18150 -20731 18170
rect -70936 18143 -56755 18150
rect -70936 18140 -70590 18143
rect -70936 18135 -70739 18140
rect -70936 18040 -70898 18135
rect -70821 18045 -70739 18135
rect -70662 18048 -70590 18140
rect -70513 18055 -56755 18143
rect -56678 18146 -36403 18150
rect -56678 18055 -46608 18146
rect -70513 18051 -46608 18055
rect -46531 18055 -36403 18146
rect -36326 18055 -26032 18150
rect -25955 18075 -20731 18150
rect -20654 18161 37954 18170
rect -20654 18157 13452 18161
rect -20654 18075 2807 18157
rect -25955 18062 2807 18075
rect 2884 18066 13452 18157
rect 13529 18154 37954 18161
rect 13529 18066 24513 18154
rect 2884 18062 24513 18066
rect -25955 18059 24513 18062
rect 24590 18150 37954 18154
rect 24590 18059 35414 18150
rect -25955 18055 35414 18059
rect 35491 18140 37954 18150
rect 35491 18137 37160 18140
rect 35491 18132 37011 18137
rect 35491 18055 36852 18132
rect -46531 18051 36852 18055
rect -70513 18048 36852 18051
rect -70662 18045 36852 18048
rect -70821 18040 36852 18045
rect -70936 18037 36852 18040
rect 36929 18042 37011 18132
rect 37088 18045 37160 18137
rect 37237 18045 37954 18140
rect 37088 18042 37954 18045
rect 36929 18037 37954 18042
rect -70936 18011 37954 18037
rect -70936 17991 -20729 18011
rect -70936 17984 -56753 17991
rect -70936 17981 -70588 17984
rect -70936 17976 -70737 17981
rect -70936 17881 -70896 17976
rect -70819 17886 -70737 17976
rect -70660 17889 -70588 17981
rect -70511 17896 -56753 17984
rect -56676 17987 -36401 17991
rect -56676 17896 -46606 17987
rect -70511 17892 -46606 17896
rect -46529 17896 -36401 17987
rect -36324 17896 -26030 17991
rect -25953 17916 -20729 17991
rect -20652 18002 37954 18011
rect -20652 17998 13454 18002
rect -20652 17916 2809 17998
rect -25953 17903 2809 17916
rect 2886 17907 13454 17998
rect 13531 17995 37954 18002
rect 13531 17907 24515 17995
rect 2886 17903 24515 17907
rect -25953 17900 24515 17903
rect 24592 17991 37954 17995
rect 24592 17900 35416 17991
rect -25953 17896 35416 17900
rect 35493 17981 37954 17991
rect 35493 17978 37162 17981
rect 35493 17973 37013 17978
rect 35493 17896 36854 17973
rect -46529 17892 36854 17896
rect -70511 17889 36854 17892
rect -70660 17886 36854 17889
rect -70819 17881 36854 17886
rect -70936 17878 36854 17881
rect 36931 17883 37013 17973
rect 37090 17886 37162 17978
rect 37239 17886 37954 17981
rect 37090 17883 37954 17886
rect 36931 17878 37954 17883
rect -70936 17853 37954 17878
rect -70936 17833 -20730 17853
rect -70936 17826 -56754 17833
rect -70936 17823 -70589 17826
rect -70936 17818 -70738 17823
rect -70936 17723 -70897 17818
rect -70820 17728 -70738 17818
rect -70661 17731 -70589 17823
rect -70512 17738 -56754 17826
rect -56677 17829 -36402 17833
rect -56677 17738 -46607 17829
rect -70512 17734 -46607 17738
rect -46530 17738 -36402 17829
rect -36325 17738 -26031 17833
rect -25954 17758 -20730 17833
rect -20653 17844 37954 17853
rect -20653 17840 13453 17844
rect -20653 17758 2808 17840
rect -25954 17745 2808 17758
rect 2885 17749 13453 17840
rect 13530 17837 37954 17844
rect 13530 17749 24514 17837
rect 2885 17745 24514 17749
rect -25954 17742 24514 17745
rect 24591 17833 37954 17837
rect 24591 17742 35415 17833
rect -25954 17738 35415 17742
rect 35492 17823 37954 17833
rect 35492 17820 37161 17823
rect 35492 17815 37012 17820
rect 35492 17738 36853 17815
rect -46530 17734 36853 17738
rect -70512 17731 36853 17734
rect -70661 17728 36853 17731
rect -70820 17723 36853 17728
rect -70936 17720 36853 17723
rect 36930 17725 37012 17815
rect 37089 17728 37161 17820
rect 37238 17728 37954 17823
rect 37089 17725 37954 17728
rect 36930 17720 37954 17725
rect -70936 17708 37954 17720
rect -53208 15933 -53063 15965
rect -53208 15877 -53166 15933
rect -53110 15877 -53063 15933
rect -53208 15822 -53063 15877
rect -53208 15766 -53170 15822
rect -53114 15766 -53063 15822
rect -63334 15703 -63247 15724
rect -63334 15647 -63321 15703
rect -63265 15690 -63247 15703
rect -53208 15690 -53063 15766
rect -32606 15760 -32519 15781
rect -32606 15704 -32593 15760
rect -32537 15704 -32519 15760
rect -32606 15690 -32519 15704
rect -63265 15649 -20108 15690
rect -3768 15673 -3681 15689
rect -63265 15647 -32597 15649
rect -63334 15622 -32597 15647
rect -63334 15592 -42963 15622
rect -63334 15536 -63325 15592
rect -63269 15566 -42963 15592
rect -42907 15593 -32597 15622
rect -32541 15593 -20108 15649
rect -42907 15566 -20108 15593
rect -63269 15545 -20108 15566
rect -63269 15536 -63247 15545
rect -63334 15521 -63247 15536
rect -42976 15511 -42889 15545
rect -42976 15455 -42967 15511
rect -42911 15455 -42889 15511
rect -42976 15440 -42889 15455
rect -20253 15406 -20108 15545
rect -20253 15320 -20225 15406
rect -20135 15320 -20108 15406
rect -20253 15201 -20108 15320
rect -20253 15115 -20229 15201
rect -20139 15115 -20108 15201
rect -9008 15668 28925 15673
rect -9008 15612 -3755 15668
rect -3699 15612 28925 15668
rect -9008 15606 28925 15612
rect -9008 15592 28938 15606
rect -9008 15582 17953 15592
rect -9008 15557 6890 15582
rect -9008 15541 -3759 15557
rect -9008 15153 -8876 15541
rect -3768 15501 -3759 15541
rect -3703 15541 6890 15557
rect -3703 15501 -3681 15541
rect -3768 15486 -3681 15501
rect 6877 15526 6890 15541
rect 6946 15541 17953 15582
rect 6946 15526 6964 15541
rect 6877 15471 6964 15526
rect 6877 15415 6886 15471
rect 6942 15415 6964 15471
rect 6877 15400 6964 15415
rect 17940 15536 17953 15541
rect 18009 15585 28938 15592
rect 18009 15541 28864 15585
rect 18009 15536 18027 15541
rect 17940 15481 18027 15536
rect 17940 15425 17949 15481
rect 18005 15425 18027 15481
rect 17940 15410 18027 15425
rect 28851 15529 28864 15541
rect 28920 15529 28938 15585
rect 28851 15474 28938 15529
rect 28851 15418 28860 15474
rect 28916 15418 28938 15474
rect 28851 15403 28938 15418
rect -20253 15090 -20108 15115
rect -9905 15114 -8876 15153
rect -9905 15113 -9726 15114
rect -9905 15037 -9885 15113
rect -9818 15038 -9726 15113
rect -9659 15038 -8876 15114
rect -9818 15037 -8876 15038
rect -9905 15021 -8876 15037
rect -24194 14096 -19559 14117
rect -24194 14094 -23950 14096
rect -53486 14035 -53359 14069
rect -53486 13979 -53461 14035
rect -53405 13979 -53359 14035
rect -24194 14008 -24175 14094
rect -24069 14010 -23950 14094
rect -23844 14010 -19559 14096
rect -24069 14008 -19559 14010
rect -24194 13988 -19559 14008
rect -53486 13924 -53359 13979
rect -53486 13868 -53465 13924
rect -53409 13868 -53359 13924
rect -63624 13763 -63537 13785
rect -63624 13749 -63611 13763
rect -68360 13716 -63611 13749
rect -68360 13646 -68333 13716
rect -68258 13707 -63611 13716
rect -63555 13749 -63537 13763
rect -53486 13749 -53359 13868
rect -32944 13852 -32857 13873
rect -32944 13796 -32931 13852
rect -32875 13796 -32857 13852
rect -32944 13749 -32857 13796
rect -8912 13768 -8567 13774
rect -20257 13749 -19895 13763
rect -63555 13741 -19895 13749
rect -63555 13722 -32935 13741
rect -63555 13718 -42561 13722
rect -63555 13707 -42693 13718
rect -68258 13664 -42693 13707
rect -68258 13652 -43268 13664
rect -68258 13646 -63615 13652
rect -68360 13622 -63615 13646
rect -63624 13596 -63615 13622
rect -63559 13622 -43268 13652
rect -63559 13596 -63537 13622
rect -63624 13581 -63537 13596
rect -43281 13608 -43268 13622
rect -43212 13635 -42693 13664
rect -42628 13639 -42561 13718
rect -42496 13685 -32935 13722
rect -32879 13729 -19895 13741
rect -32879 13726 -20022 13729
rect -32879 13685 -20237 13726
rect -42496 13639 -20237 13685
rect -42628 13635 -20237 13639
rect -43212 13625 -20237 13635
rect -20151 13628 -20022 13726
rect -19936 13628 -19895 13729
rect -20151 13625 -19895 13628
rect -43212 13622 -19895 13625
rect -43212 13608 -43194 13622
rect -20257 13609 -19895 13622
rect -8912 13741 28701 13768
rect -8912 13730 -4098 13741
rect -8912 13727 -8685 13730
rect -8912 13624 -8891 13727
rect -8801 13627 -8685 13727
rect -8595 13685 -4098 13730
rect -4042 13730 28701 13741
rect -4042 13685 6644 13730
rect -8595 13674 6644 13685
rect 6700 13723 28701 13730
rect 6700 13700 28540 13723
rect 6700 13674 17640 13700
rect -8595 13644 17640 13674
rect 17696 13667 28540 13700
rect 28596 13667 28701 13723
rect 17696 13644 28701 13667
rect -8595 13630 28701 13644
rect -8595 13627 -4102 13630
rect -8801 13624 -4102 13627
rect -43281 13553 -43194 13608
rect -8912 13607 -4102 13624
rect -8912 13590 -8567 13607
rect -4111 13574 -4102 13607
rect -4046 13619 28701 13630
rect -4046 13607 6640 13619
rect -4046 13574 -4024 13607
rect -4111 13559 -4024 13574
rect 6631 13563 6640 13607
rect 6696 13612 28701 13619
rect 6696 13607 28536 13612
rect 6696 13563 6718 13607
rect -43281 13497 -43272 13553
rect -43216 13497 -43194 13553
rect 6631 13548 6718 13563
rect 17627 13589 17714 13607
rect 17627 13533 17636 13589
rect 17692 13533 17714 13589
rect 28527 13556 28536 13607
rect 28592 13607 28701 13612
rect 28592 13556 28614 13607
rect 28527 13541 28614 13556
rect 17627 13518 17714 13533
rect -43281 13482 -43194 13497
rect -71933 11310 -70484 11335
rect -71933 11197 -71904 11310
rect -71787 11307 -70484 11310
rect -71787 11197 -71610 11307
rect -71933 11194 -71610 11197
rect -71493 11194 -70484 11307
rect -71933 11012 -70484 11194
rect -71933 10899 -71907 11012
rect -71790 10899 -71617 11012
rect -71500 10899 -70484 11012
rect -71933 10868 -70484 10899
rect -70951 9624 -70484 10868
rect -18808 9846 -18709 9847
rect -18815 9831 -18709 9846
rect -18815 9756 -18798 9831
rect -18733 9756 -18709 9831
rect -18815 9744 -18709 9756
rect -18815 9743 -18716 9744
rect -70951 9517 -21319 9624
rect -70951 9264 -21250 9517
rect -70951 9157 -21319 9264
rect -18798 8715 -18733 9743
rect -16592 9493 -16536 9590
rect -18818 8703 -18712 8715
rect -18818 8635 -18798 8703
rect -18733 8635 -18712 8703
rect -18818 8569 -18712 8635
rect -18818 8504 -18798 8569
rect -18733 8504 -18712 8569
rect -18818 8483 -18712 8504
rect -15955 7636 -15780 7723
rect -15867 7632 -15782 7636
rect -56587 7419 -56486 7422
rect -46437 7419 -46336 7422
rect 13860 7419 13961 7422
rect -70936 7396 -27005 7419
rect -70936 7380 -56569 7396
rect -70936 7377 -69895 7380
rect -70936 7372 -70044 7377
rect -70936 7277 -70203 7372
rect -70126 7282 -70044 7372
rect -69967 7285 -69895 7377
rect -69818 7301 -56569 7380
rect -56492 7301 -46419 7396
rect -46342 7393 -27005 7396
rect -46342 7301 -36009 7393
rect -69818 7298 -36009 7301
rect -35932 7389 -27005 7393
rect -35932 7298 -27090 7389
rect -69818 7294 -27090 7298
rect -27013 7294 -27005 7389
rect -69818 7285 -27005 7294
rect -69967 7282 -27005 7285
rect -70126 7277 -27005 7282
rect -70936 7220 -27005 7277
rect -70936 7204 -56572 7220
rect -70936 7201 -69898 7204
rect -70936 7196 -70047 7201
rect -70936 7101 -70206 7196
rect -70129 7106 -70047 7196
rect -69970 7109 -69898 7201
rect -69821 7125 -56572 7204
rect -56495 7125 -46422 7220
rect -46345 7217 -27005 7220
rect -46345 7125 -36012 7217
rect -69821 7122 -36012 7125
rect -35935 7213 -27005 7217
rect -35935 7122 -27093 7213
rect -69821 7118 -27093 7122
rect -27016 7118 -27005 7213
rect -69821 7109 -27005 7118
rect -69970 7106 -27005 7109
rect -70129 7101 -27005 7106
rect -70936 7061 -27005 7101
rect -70936 7045 -56570 7061
rect -70936 7042 -69896 7045
rect -70936 7037 -70045 7042
rect -70936 6942 -70204 7037
rect -70127 6947 -70045 7037
rect -69968 6950 -69896 7042
rect -69819 6966 -56570 7045
rect -56493 6966 -46420 7061
rect -46343 7058 -27005 7061
rect -46343 6966 -36010 7058
rect -69819 6963 -36010 6966
rect -35933 7054 -27005 7058
rect -35933 6963 -27091 7054
rect -69819 6959 -27091 6963
rect -27014 6959 -27005 7054
rect -69819 6950 -27005 6959
rect -69968 6947 -27005 6950
rect -70127 6942 -27005 6947
rect -70936 6903 -27005 6942
rect -70936 6887 -56571 6903
rect -70936 6884 -69897 6887
rect -70936 6879 -70046 6884
rect -70936 6784 -70205 6879
rect -70128 6789 -70046 6879
rect -69969 6792 -69897 6884
rect -69820 6808 -56571 6887
rect -56494 6808 -46421 6903
rect -46344 6900 -27005 6903
rect -46344 6808 -36011 6900
rect -69820 6805 -36011 6808
rect -35934 6896 -27005 6900
rect -35934 6805 -27092 6896
rect -69820 6801 -27092 6805
rect -27015 6801 -27005 6896
rect -69820 6792 -27005 6801
rect -69969 6789 -27005 6792
rect -70128 6784 -27005 6789
rect -70936 6773 -27005 6784
rect 3014 7396 37954 7419
rect 3014 7392 13878 7396
rect 3014 7297 3048 7392
rect 3125 7301 13878 7392
rect 13955 7392 37954 7396
rect 13955 7389 35391 7392
rect 13955 7301 24719 7389
rect 3125 7297 24719 7301
rect 3014 7294 24719 7297
rect 24796 7297 35391 7389
rect 35468 7379 37954 7392
rect 35468 7376 37857 7379
rect 35468 7371 37708 7376
rect 35468 7297 37549 7371
rect 24796 7294 37549 7297
rect 3014 7276 37549 7294
rect 37626 7281 37708 7371
rect 37785 7284 37857 7376
rect 37934 7284 37954 7379
rect 37785 7281 37954 7284
rect 37626 7276 37954 7281
rect 3014 7220 37954 7276
rect 3014 7216 13875 7220
rect 3014 7121 3045 7216
rect 3122 7125 13875 7216
rect 13952 7216 37954 7220
rect 13952 7213 35388 7216
rect 13952 7125 24716 7213
rect 3122 7121 24716 7125
rect 3014 7118 24716 7121
rect 24793 7121 35388 7213
rect 35465 7203 37954 7216
rect 35465 7200 37854 7203
rect 35465 7195 37705 7200
rect 35465 7121 37546 7195
rect 24793 7118 37546 7121
rect 3014 7100 37546 7118
rect 37623 7105 37705 7195
rect 37782 7108 37854 7200
rect 37931 7108 37954 7203
rect 37782 7105 37954 7108
rect 37623 7100 37954 7105
rect 3014 7061 37954 7100
rect 3014 7057 13877 7061
rect 3014 6962 3047 7057
rect 3124 6966 13877 7057
rect 13954 7057 37954 7061
rect 13954 7054 35390 7057
rect 13954 6966 24718 7054
rect 3124 6962 24718 6966
rect 3014 6959 24718 6962
rect 24795 6962 35390 7054
rect 35467 7044 37954 7057
rect 35467 7041 37856 7044
rect 35467 7036 37707 7041
rect 35467 6962 37548 7036
rect 24795 6959 37548 6962
rect 3014 6941 37548 6959
rect 37625 6946 37707 7036
rect 37784 6949 37856 7041
rect 37933 6949 37954 7044
rect 37784 6946 37954 6949
rect 37625 6941 37954 6946
rect 3014 6903 37954 6941
rect 3014 6899 13876 6903
rect 3014 6804 3046 6899
rect 3123 6808 13876 6899
rect 13953 6899 37954 6903
rect 13953 6896 35389 6899
rect 13953 6808 24717 6896
rect 3123 6804 24717 6808
rect 3014 6801 24717 6804
rect 24794 6804 35389 6896
rect 35466 6886 37954 6899
rect 35466 6883 37855 6886
rect 35466 6878 37706 6883
rect 35466 6804 37547 6878
rect 24794 6801 37547 6804
rect 3014 6783 37547 6801
rect 37624 6788 37706 6878
rect 37783 6791 37855 6883
rect 37932 6791 37954 6886
rect 37783 6788 37954 6791
rect 37624 6783 37954 6788
rect 3014 6773 37954 6783
rect -70219 6771 -69812 6773
rect -70936 6161 -27810 6188
rect -70936 6157 -46623 6161
rect -70936 6150 -56773 6157
rect -70936 6147 -70591 6150
rect -70936 6142 -70740 6147
rect -70936 6047 -70899 6142
rect -70822 6052 -70740 6142
rect -70663 6055 -70591 6147
rect -70514 6062 -56773 6150
rect -56696 6066 -46623 6157
rect -46546 6154 -27916 6161
rect -46546 6066 -36217 6154
rect -56696 6062 -36217 6066
rect -70514 6059 -36217 6062
rect -36140 6066 -27916 6154
rect -27839 6066 -27810 6161
rect -36140 6059 -27810 6066
rect -70514 6055 -27810 6059
rect -70663 6052 -27810 6055
rect -70822 6047 -27810 6052
rect -70936 5985 -27810 6047
rect -70936 5981 -46626 5985
rect -70936 5974 -56776 5981
rect -70936 5971 -70594 5974
rect -70936 5966 -70743 5971
rect -70936 5871 -70902 5966
rect -70825 5876 -70743 5966
rect -70666 5879 -70594 5971
rect -70517 5886 -56776 5974
rect -56699 5890 -46626 5981
rect -46549 5978 -27919 5985
rect -46549 5890 -36220 5978
rect -56699 5886 -36220 5890
rect -70517 5883 -36220 5886
rect -36143 5890 -27919 5978
rect -27842 5890 -27810 5985
rect 2814 6162 37954 6188
rect 2814 6155 13673 6162
rect 2814 6060 2843 6155
rect 2920 6067 13673 6155
rect 13750 6159 37954 6162
rect 13750 6158 37167 6159
rect 13750 6067 24517 6158
rect 2920 6063 24517 6067
rect 24594 6156 37167 6158
rect 24594 6155 37018 6156
rect 24594 6063 35190 6155
rect 2920 6060 35190 6063
rect 35267 6151 37018 6155
rect 35267 6060 36859 6151
rect 2814 6056 36859 6060
rect 36936 6061 37018 6151
rect 37095 6064 37167 6156
rect 37244 6064 37954 6159
rect 37095 6061 37954 6064
rect 36936 6056 37954 6061
rect 2814 5986 37954 6056
rect 2814 5979 13670 5986
rect -15885 5917 -15765 5978
rect -36143 5883 -27810 5890
rect -70517 5879 -27810 5883
rect -70666 5876 -27810 5879
rect -70825 5871 -27810 5876
rect -70936 5826 -27810 5871
rect -70936 5822 -46624 5826
rect -70936 5815 -56774 5822
rect -70936 5812 -70592 5815
rect -70936 5807 -70741 5812
rect -70936 5712 -70900 5807
rect -70823 5717 -70741 5807
rect -70664 5720 -70592 5812
rect -70515 5727 -56774 5815
rect -56697 5731 -46624 5822
rect -46547 5819 -27917 5826
rect -46547 5731 -36218 5819
rect -56697 5727 -36218 5731
rect -70515 5724 -36218 5727
rect -36141 5731 -27917 5819
rect -27840 5731 -27810 5826
rect -36141 5724 -27810 5731
rect -70515 5720 -27810 5724
rect -70664 5717 -27810 5720
rect -70823 5712 -27810 5717
rect -70936 5668 -27810 5712
rect -70936 5664 -46625 5668
rect -70936 5657 -56775 5664
rect -70936 5654 -70593 5657
rect -70936 5649 -70742 5654
rect -70936 5554 -70901 5649
rect -70824 5559 -70742 5649
rect -70665 5562 -70593 5654
rect -70516 5569 -56775 5657
rect -56698 5573 -46625 5664
rect -46548 5661 -27918 5668
rect -46548 5573 -36219 5661
rect -56698 5569 -36219 5573
rect -70516 5566 -36219 5569
rect -36142 5573 -27918 5661
rect -27841 5573 -27810 5668
rect -36142 5566 -27810 5573
rect -70516 5562 -27810 5566
rect -70665 5559 -27810 5562
rect -70824 5554 -27810 5559
rect -70936 5542 -27810 5554
rect 2814 5884 2840 5979
rect 2917 5891 13670 5979
rect 13747 5983 37954 5986
rect 13747 5982 37164 5983
rect 13747 5891 24514 5982
rect 2917 5887 24514 5891
rect 24591 5980 37164 5982
rect 24591 5979 37015 5980
rect 24591 5887 35187 5979
rect 2917 5884 35187 5887
rect 35264 5975 37015 5979
rect 35264 5884 36856 5975
rect 2814 5880 36856 5884
rect 36933 5885 37015 5975
rect 37092 5888 37164 5980
rect 37241 5888 37954 5983
rect 37092 5885 37954 5888
rect 36933 5880 37954 5885
rect 2814 5827 37954 5880
rect 2814 5820 13672 5827
rect 2814 5725 2842 5820
rect 2919 5732 13672 5820
rect 13749 5824 37954 5827
rect 13749 5823 37166 5824
rect 13749 5732 24516 5823
rect 2919 5728 24516 5732
rect 24593 5821 37166 5823
rect 24593 5820 37017 5821
rect 24593 5728 35189 5820
rect 2919 5725 35189 5728
rect 35266 5816 37017 5820
rect 35266 5725 36858 5816
rect 2814 5721 36858 5725
rect 36935 5726 37017 5816
rect 37094 5729 37166 5821
rect 37243 5729 37954 5824
rect 37094 5726 37954 5729
rect 36935 5721 37954 5726
rect 2814 5669 37954 5721
rect 2814 5662 13671 5669
rect 2814 5567 2841 5662
rect 2918 5574 13671 5662
rect 13748 5666 37954 5669
rect 13748 5665 37165 5666
rect 13748 5574 24515 5665
rect 2918 5570 24515 5574
rect 24592 5663 37165 5665
rect 24592 5662 37016 5663
rect 24592 5570 35188 5662
rect 2918 5567 35188 5570
rect 35265 5658 37016 5662
rect 35265 5567 36857 5658
rect 2814 5563 36857 5567
rect 36934 5568 37016 5658
rect 37093 5571 37165 5663
rect 37242 5571 37954 5666
rect 37093 5568 37954 5571
rect 36934 5563 37954 5568
rect 2814 5542 37954 5563
rect -70915 5541 -70508 5542
rect -12824 5052 -12600 5117
rect -63342 3380 -63255 3401
rect -63342 3324 -63329 3380
rect -63273 3357 -63255 3380
rect -63273 3324 28723 3357
rect -63342 3269 28723 3324
rect -63342 3213 -63333 3269
rect -63277 3230 28723 3269
rect -63277 3213 -63255 3230
rect -63342 3198 -63255 3213
rect -53222 3049 -53095 3230
rect -53222 2993 -53194 3049
rect -53138 2993 -53095 3049
rect -53222 2938 -53095 2993
rect -53222 2882 -53198 2938
rect -53142 2882 -53095 2938
rect -53222 2854 -53095 2882
rect -42830 2816 -42703 3230
rect -42830 2760 -42778 2816
rect -42722 2760 -42703 2816
rect -42830 2705 -42703 2760
rect -42830 2649 -42782 2705
rect -42726 2649 -42703 2705
rect -32546 2839 -32419 3230
rect -3803 2996 -3676 3230
rect 7061 3168 7250 3230
rect 7061 3112 7116 3168
rect 7172 3151 7250 3168
rect 7172 3112 7190 3151
rect 7061 3069 7190 3112
rect 7103 3057 7190 3069
rect 7103 3001 7112 3057
rect 7168 3001 7190 3057
rect -3803 2975 -3633 2996
rect 7103 2986 7190 3001
rect 17915 3088 18042 3230
rect 17915 3032 17962 3088
rect 18018 3032 18042 3088
rect 17915 2987 18042 3032
rect -3803 2919 -3707 2975
rect -3651 2919 -3633 2975
rect -3803 2864 -3633 2919
rect 17949 2977 18036 2987
rect 17949 2921 17958 2977
rect 18014 2921 18036 2977
rect 17949 2906 18036 2921
rect -3803 2843 -3711 2864
rect -32546 2818 -32400 2839
rect -32546 2762 -32474 2818
rect -32418 2762 -32400 2818
rect -3720 2808 -3711 2843
rect -3655 2808 -3633 2864
rect -3720 2793 -3633 2808
rect 28596 2863 28723 3230
rect 28596 2807 28622 2863
rect 28678 2807 28723 2863
rect -32546 2707 -32400 2762
rect 28596 2752 28723 2807
rect 28596 2743 28618 2752
rect -32546 2656 -32478 2707
rect -42830 2631 -42703 2649
rect -32487 2651 -32478 2656
rect -32422 2651 -32400 2707
rect 28609 2696 28618 2743
rect 28674 2743 28723 2752
rect 28674 2696 28696 2743
rect 28609 2681 28696 2696
rect -32487 2636 -32400 2651
rect -63781 1410 -63644 1453
rect -63781 1354 -63742 1410
rect -63686 1354 -63644 1410
rect -63781 1299 -63644 1354
rect -63781 1243 -63746 1299
rect -63690 1243 -63644 1299
rect -68362 1157 -68225 1175
rect -68362 1064 -68328 1157
rect -68246 1106 -68225 1157
rect -63781 1106 -63644 1243
rect 6759 1266 6846 1287
rect 6759 1210 6772 1266
rect 6828 1210 6846 1266
rect 6759 1155 6846 1210
rect 6759 1129 6768 1155
rect -53640 1106 -53553 1115
rect -68246 1094 -43366 1106
rect -68246 1064 -53627 1094
rect -68362 1038 -53627 1064
rect -53571 1073 -43366 1094
rect -53571 1062 -52878 1073
rect -53571 1038 -53009 1062
rect -68362 984 -53009 1038
rect -52949 995 -52878 1062
rect -52818 995 -43366 1073
rect 6403 1099 6768 1129
rect 6824 1129 6846 1155
rect 17564 1148 17651 1169
rect 17564 1129 17577 1148
rect 6824 1099 17577 1129
rect 6403 1092 17577 1099
rect 17633 1129 17651 1148
rect 17633 1092 28175 1129
rect -52949 984 -43366 995
rect -4084 1040 -3997 1061
rect -68362 983 -43366 984
rect -68362 969 -53631 983
rect -53640 927 -53631 969
rect -53575 969 -43366 983
rect -53575 927 -53553 969
rect -53640 912 -53553 927
rect -43503 941 -43366 969
rect -32846 967 -32759 988
rect -32846 941 -32833 967
rect -43503 911 -32833 941
rect -32777 941 -32759 967
rect -4084 984 -4071 1040
rect -4015 984 -3997 1040
rect -4084 941 -3997 984
rect 6403 1037 28175 1092
rect 6403 992 17573 1037
rect 6403 941 6540 992
rect 17564 981 17573 992
rect 17629 992 28175 1037
rect 17629 981 17651 992
rect 17564 966 17651 981
rect -32777 929 6540 941
rect -32777 911 -4075 929
rect -43503 907 -4075 911
rect -43503 851 -43134 907
rect -43078 873 -4075 907
rect -4019 873 6540 929
rect -43078 856 6540 873
rect -43078 851 -32837 856
rect -43503 804 -32837 851
rect -43147 796 -43060 804
rect -43147 740 -43138 796
rect -43082 740 -43060 796
rect -32846 800 -32837 804
rect -32781 804 6540 856
rect 28038 917 28175 992
rect 28335 951 28422 972
rect 28335 917 28348 951
rect 28038 895 28348 917
rect 28404 917 28422 951
rect 28404 895 28611 917
rect 28038 840 28611 895
rect -32781 800 -32759 804
rect -32846 785 -32759 800
rect 28038 784 28344 840
rect 28400 784 28611 840
rect 28038 780 28611 784
rect 28335 769 28422 780
rect -43147 725 -43060 740
rect -70936 -2455 37954 -2429
rect -70936 -2461 -56591 -2455
rect -70936 -2464 -69895 -2461
rect -70936 -2469 -70044 -2464
rect -70936 -2564 -70203 -2469
rect -70126 -2559 -70044 -2469
rect -69967 -2556 -69895 -2464
rect -69818 -2550 -56591 -2461
rect -56514 -2550 -36040 -2455
rect -35963 -2550 -12562 -2455
rect -12485 -2550 13859 -2455
rect 13936 -2472 37954 -2455
rect 13936 -2475 37849 -2472
rect 13936 -2480 37700 -2475
rect 13936 -2550 37541 -2480
rect -69818 -2556 37541 -2550
rect -69967 -2559 37541 -2556
rect -70126 -2564 37541 -2559
rect -70936 -2575 37541 -2564
rect 37618 -2570 37700 -2480
rect 37777 -2567 37849 -2475
rect 37926 -2567 37954 -2472
rect 37777 -2570 37954 -2567
rect 37618 -2575 37954 -2570
rect -70936 -2631 37954 -2575
rect -70936 -2637 -56594 -2631
rect -70936 -2640 -69898 -2637
rect -70936 -2645 -70047 -2640
rect -70936 -2740 -70206 -2645
rect -70129 -2735 -70047 -2645
rect -69970 -2732 -69898 -2640
rect -69821 -2726 -56594 -2637
rect -56517 -2726 -36043 -2631
rect -35966 -2726 -12565 -2631
rect -12488 -2726 13856 -2631
rect 13933 -2648 37954 -2631
rect 13933 -2651 37846 -2648
rect 13933 -2656 37697 -2651
rect 13933 -2726 37538 -2656
rect -69821 -2732 37538 -2726
rect -69970 -2735 37538 -2732
rect -70129 -2740 37538 -2735
rect -70936 -2751 37538 -2740
rect 37615 -2746 37697 -2656
rect 37774 -2743 37846 -2651
rect 37923 -2743 37954 -2648
rect 37774 -2746 37954 -2743
rect 37615 -2751 37954 -2746
rect -70936 -2790 37954 -2751
rect -70936 -2796 -56592 -2790
rect -70936 -2799 -69896 -2796
rect -70936 -2804 -70045 -2799
rect -70936 -2899 -70204 -2804
rect -70127 -2894 -70045 -2804
rect -69968 -2891 -69896 -2799
rect -69819 -2885 -56592 -2796
rect -56515 -2885 -36041 -2790
rect -35964 -2885 -12563 -2790
rect -12486 -2885 13858 -2790
rect 13935 -2807 37954 -2790
rect 13935 -2810 37848 -2807
rect 13935 -2815 37699 -2810
rect 13935 -2885 37540 -2815
rect -69819 -2891 37540 -2885
rect -69968 -2894 37540 -2891
rect -70127 -2899 37540 -2894
rect -70936 -2910 37540 -2899
rect 37617 -2905 37699 -2815
rect 37776 -2902 37848 -2810
rect 37925 -2902 37954 -2807
rect 37776 -2905 37954 -2902
rect 37617 -2910 37954 -2905
rect -70936 -2948 37954 -2910
rect -70936 -2954 -56593 -2948
rect -70936 -2957 -69897 -2954
rect -70936 -2962 -70046 -2957
rect -70936 -3057 -70205 -2962
rect -70128 -3052 -70046 -2962
rect -69969 -3049 -69897 -2957
rect -69820 -3043 -56593 -2954
rect -56516 -3043 -36042 -2948
rect -35965 -3043 -12564 -2948
rect -12487 -3043 13857 -2948
rect 13934 -2965 37954 -2948
rect 13934 -2968 37847 -2965
rect 13934 -2973 37698 -2968
rect 13934 -3043 37539 -2973
rect -69820 -3049 37539 -3043
rect -69969 -3052 37539 -3049
rect -70128 -3057 37539 -3052
rect -70936 -3068 37539 -3057
rect 37616 -3063 37698 -2973
rect 37775 -3060 37847 -2968
rect 37924 -3060 37954 -2965
rect 37775 -3063 37954 -3060
rect 37616 -3068 37954 -3063
rect -70936 -3075 37954 -3068
rect 37521 -3078 37933 -3075
rect -56812 -3501 -56711 -3500
rect 13638 -3501 13739 -3500
rect -70936 -3526 37954 -3501
rect -70936 -3542 -56794 -3526
rect -70936 -3545 -70583 -3542
rect -70936 -3550 -70732 -3545
rect -70936 -3645 -70891 -3550
rect -70814 -3640 -70732 -3550
rect -70655 -3637 -70583 -3545
rect -70506 -3621 -56794 -3542
rect -56717 -3529 13656 -3526
rect -56717 -3621 -36247 -3529
rect -70506 -3624 -36247 -3621
rect -36170 -3533 13656 -3529
rect -36170 -3624 -12768 -3533
rect -70506 -3628 -12768 -3624
rect -12691 -3621 13656 -3533
rect 13733 -3542 37954 -3526
rect 13733 -3545 37159 -3542
rect 13733 -3550 37010 -3545
rect 13733 -3621 36851 -3550
rect -12691 -3628 36851 -3621
rect -70506 -3637 36851 -3628
rect -70655 -3640 36851 -3637
rect -70814 -3645 36851 -3640
rect 36928 -3640 37010 -3550
rect 37087 -3637 37159 -3545
rect 37236 -3637 37954 -3542
rect 37087 -3640 37954 -3637
rect 36928 -3645 37954 -3640
rect -70936 -3702 37954 -3645
rect -70936 -3718 -56797 -3702
rect -70936 -3721 -70586 -3718
rect -70936 -3726 -70735 -3721
rect -70936 -3821 -70894 -3726
rect -70817 -3816 -70735 -3726
rect -70658 -3813 -70586 -3721
rect -70509 -3797 -56797 -3718
rect -56720 -3705 13653 -3702
rect -56720 -3797 -36250 -3705
rect -70509 -3800 -36250 -3797
rect -36173 -3709 13653 -3705
rect -36173 -3800 -12771 -3709
rect -70509 -3804 -12771 -3800
rect -12694 -3797 13653 -3709
rect 13730 -3718 37954 -3702
rect 13730 -3721 37156 -3718
rect 13730 -3726 37007 -3721
rect 13730 -3797 36848 -3726
rect -12694 -3804 36848 -3797
rect -70509 -3813 36848 -3804
rect -70658 -3816 36848 -3813
rect -70817 -3821 36848 -3816
rect 36925 -3816 37007 -3726
rect 37084 -3813 37156 -3721
rect 37233 -3813 37954 -3718
rect 37084 -3816 37954 -3813
rect 36925 -3821 37954 -3816
rect -70936 -3861 37954 -3821
rect -70936 -3877 -56795 -3861
rect -70936 -3880 -70584 -3877
rect -70936 -3885 -70733 -3880
rect -70936 -3980 -70892 -3885
rect -70815 -3975 -70733 -3885
rect -70656 -3972 -70584 -3880
rect -70507 -3956 -56795 -3877
rect -56718 -3864 13655 -3861
rect -56718 -3956 -36248 -3864
rect -70507 -3959 -36248 -3956
rect -36171 -3868 13655 -3864
rect -36171 -3959 -12769 -3868
rect -70507 -3963 -12769 -3959
rect -12692 -3956 13655 -3868
rect 13732 -3877 37954 -3861
rect 13732 -3880 37158 -3877
rect 13732 -3885 37009 -3880
rect 13732 -3956 36850 -3885
rect -12692 -3963 36850 -3956
rect -70507 -3972 36850 -3963
rect -70656 -3975 36850 -3972
rect -70815 -3980 36850 -3975
rect 36927 -3975 37009 -3885
rect 37086 -3972 37158 -3880
rect 37235 -3972 37954 -3877
rect 37086 -3975 37954 -3972
rect 36927 -3980 37954 -3975
rect -70936 -4019 37954 -3980
rect -70936 -4035 -56796 -4019
rect -70936 -4038 -70585 -4035
rect -70936 -4043 -70734 -4038
rect -70936 -4138 -70893 -4043
rect -70816 -4133 -70734 -4043
rect -70657 -4130 -70585 -4038
rect -70508 -4114 -56796 -4035
rect -56719 -4022 13654 -4019
rect -56719 -4114 -36249 -4022
rect -70508 -4117 -36249 -4114
rect -36172 -4026 13654 -4022
rect -36172 -4117 -12770 -4026
rect -70508 -4121 -12770 -4117
rect -12693 -4114 13654 -4026
rect 13731 -4035 37954 -4019
rect 13731 -4038 37157 -4035
rect 13731 -4043 37008 -4038
rect 13731 -4114 36849 -4043
rect -12693 -4121 36849 -4114
rect -70508 -4130 36849 -4121
rect -70657 -4133 36849 -4130
rect -70816 -4138 36849 -4133
rect 36926 -4133 37008 -4043
rect 37085 -4130 37157 -4038
rect 37234 -4130 37954 -4035
rect 37085 -4133 37954 -4130
rect 36926 -4138 37954 -4133
rect -70936 -4147 37954 -4138
rect -70907 -4151 -70500 -4147
rect 36831 -4148 37243 -4147
rect -63401 -6101 -63270 -6038
rect -63401 -6122 -63264 -6101
rect -63401 -6178 -63338 -6122
rect -63282 -6178 -63264 -6122
rect -63401 -6233 -63264 -6178
rect -63401 -6289 -63342 -6233
rect -63286 -6289 -63264 -6233
rect -63401 -6304 -63264 -6289
rect -42817 -6147 -42686 -6122
rect -42817 -6203 -42799 -6147
rect -42743 -6203 -42686 -6147
rect -42817 -6258 -42686 -6203
rect -63401 -6374 -63270 -6304
rect -42817 -6314 -42803 -6258
rect -42747 -6314 -42686 -6258
rect -42817 -6374 -42686 -6314
rect -19355 -6183 -19224 -6156
rect -19355 -6239 -19334 -6183
rect -19278 -6239 -19224 -6183
rect -19355 -6294 -19224 -6239
rect -19355 -6350 -19338 -6294
rect -19282 -6350 -19224 -6294
rect -19355 -6374 -19224 -6350
rect 7086 -6370 7173 -6349
rect 7086 -6374 7099 -6370
rect -63401 -6426 7099 -6374
rect 7155 -6426 7173 -6370
rect -63401 -6481 7173 -6426
rect -63401 -6505 7095 -6481
rect 7086 -6537 7095 -6505
rect 7151 -6537 7173 -6481
rect 7086 -6552 7173 -6537
rect -68404 -7856 -68270 -7804
rect -68404 -7936 -68380 -7856
rect -68289 -7936 -68270 -7856
rect -68404 -8031 -68270 -7936
rect -68404 -8111 -68379 -8031
rect -68288 -8103 -68270 -8031
rect -43130 -8034 -42977 -8009
rect -64344 -8086 -64257 -8065
rect -64344 -8103 -64331 -8086
rect -68288 -8111 -64331 -8103
rect -68404 -8142 -64331 -8111
rect -64275 -8103 -64257 -8086
rect -43130 -8103 -43097 -8034
rect -64275 -8116 -43097 -8103
rect -43015 -8103 -42977 -8034
rect -42686 -8103 -42426 -8102
rect -43015 -8116 6589 -8103
rect -64275 -8133 6589 -8116
rect -64275 -8137 -42509 -8133
rect -64275 -8142 -42673 -8137
rect -68404 -8197 -42673 -8142
rect -68404 -8237 -64335 -8197
rect -64344 -8253 -64335 -8237
rect -64279 -8199 -42673 -8197
rect -64279 -8237 -43097 -8199
rect -64279 -8253 -64257 -8237
rect -64344 -8268 -64257 -8253
rect -43130 -8281 -43097 -8237
rect -43015 -8223 -42673 -8199
rect -42605 -8219 -42509 -8137
rect -42441 -8219 6589 -8133
rect -42605 -8223 6589 -8219
rect -43015 -8232 6589 -8223
rect -43015 -8237 -19850 -8232
rect -43015 -8281 -42977 -8237
rect -43130 -8294 -42977 -8281
rect -19867 -8314 -19850 -8237
rect -19768 -8314 -19685 -8232
rect -19603 -8237 6589 -8232
rect -19603 -8314 -19572 -8237
rect -19867 -8361 -19572 -8314
rect 6455 -8295 6589 -8237
rect 6455 -8328 6745 -8295
rect 6455 -8410 6473 -8328
rect 6555 -8410 6638 -8328
rect 6720 -8410 6745 -8328
rect 6455 -8448 6745 -8410
rect 6455 -8450 6589 -8448
rect -36216 -11353 -36115 -11351
rect -25120 -11353 -25019 -11351
rect -11108 -11353 -11007 -11351
rect 35382 -11353 35483 -11351
rect -70936 -11377 37954 -11353
rect -70936 -11381 -36198 -11377
rect -70936 -11386 -56585 -11381
rect -70936 -11389 -69891 -11386
rect -70936 -11394 -70040 -11389
rect -70936 -11489 -70199 -11394
rect -70122 -11484 -70040 -11394
rect -69963 -11481 -69891 -11389
rect -69814 -11476 -56585 -11386
rect -56508 -11472 -36198 -11381
rect -36121 -11472 -25102 -11377
rect -25025 -11472 -11090 -11377
rect -11013 -11381 35400 -11377
rect -11013 -11472 3091 -11381
rect -56508 -11476 3091 -11472
rect 3168 -11476 13862 -11381
rect 13939 -11476 24703 -11381
rect 24780 -11472 35400 -11381
rect 35477 -11393 37954 -11377
rect 35477 -11396 37849 -11393
rect 35477 -11401 37700 -11396
rect 35477 -11472 37541 -11401
rect 24780 -11476 37541 -11472
rect -69814 -11481 37541 -11476
rect -69963 -11484 37541 -11481
rect -70122 -11489 37541 -11484
rect -70936 -11496 37541 -11489
rect 37618 -11491 37700 -11401
rect 37777 -11488 37849 -11396
rect 37926 -11488 37954 -11393
rect 37777 -11491 37954 -11488
rect 37618 -11496 37954 -11491
rect -70936 -11553 37954 -11496
rect -70936 -11557 -36201 -11553
rect -70936 -11562 -56588 -11557
rect -70936 -11565 -69894 -11562
rect -70936 -11570 -70043 -11565
rect -70936 -11665 -70202 -11570
rect -70125 -11660 -70043 -11570
rect -69966 -11657 -69894 -11565
rect -69817 -11652 -56588 -11562
rect -56511 -11648 -36201 -11557
rect -36124 -11648 -25105 -11553
rect -25028 -11648 -11093 -11553
rect -11016 -11557 35397 -11553
rect -11016 -11648 3088 -11557
rect -56511 -11652 3088 -11648
rect 3165 -11652 13859 -11557
rect 13936 -11652 24700 -11557
rect 24777 -11648 35397 -11557
rect 35474 -11569 37954 -11553
rect 35474 -11572 37846 -11569
rect 35474 -11577 37697 -11572
rect 35474 -11648 37538 -11577
rect 24777 -11652 37538 -11648
rect -69817 -11657 37538 -11652
rect -69966 -11660 37538 -11657
rect -70125 -11665 37538 -11660
rect -70936 -11672 37538 -11665
rect 37615 -11667 37697 -11577
rect 37774 -11664 37846 -11572
rect 37923 -11664 37954 -11569
rect 37774 -11667 37954 -11664
rect 37615 -11672 37954 -11667
rect -70936 -11712 37954 -11672
rect -70936 -11716 -36199 -11712
rect -70936 -11721 -56586 -11716
rect -70936 -11724 -69892 -11721
rect -70936 -11729 -70041 -11724
rect -70936 -11824 -70200 -11729
rect -70123 -11819 -70041 -11729
rect -69964 -11816 -69892 -11724
rect -69815 -11811 -56586 -11721
rect -56509 -11807 -36199 -11716
rect -36122 -11807 -25103 -11712
rect -25026 -11807 -11091 -11712
rect -11014 -11716 35399 -11712
rect -11014 -11807 3090 -11716
rect -56509 -11811 3090 -11807
rect 3167 -11811 13861 -11716
rect 13938 -11811 24702 -11716
rect 24779 -11807 35399 -11716
rect 35476 -11728 37954 -11712
rect 35476 -11731 37848 -11728
rect 35476 -11736 37699 -11731
rect 35476 -11807 37540 -11736
rect 24779 -11811 37540 -11807
rect -69815 -11816 37540 -11811
rect -69964 -11819 37540 -11816
rect -70123 -11824 37540 -11819
rect -70936 -11831 37540 -11824
rect 37617 -11826 37699 -11736
rect 37776 -11823 37848 -11731
rect 37925 -11823 37954 -11728
rect 37776 -11826 37954 -11823
rect 37617 -11831 37954 -11826
rect -70936 -11870 37954 -11831
rect -70936 -11874 -36200 -11870
rect -70936 -11879 -56587 -11874
rect -70936 -11882 -69893 -11879
rect -70936 -11887 -70042 -11882
rect -70936 -11982 -70201 -11887
rect -70124 -11977 -70042 -11887
rect -69965 -11974 -69893 -11882
rect -69816 -11969 -56587 -11879
rect -56510 -11965 -36200 -11874
rect -36123 -11965 -25104 -11870
rect -25027 -11965 -11092 -11870
rect -11015 -11874 35398 -11870
rect -11015 -11965 3089 -11874
rect -56510 -11969 3089 -11965
rect 3166 -11969 13860 -11874
rect 13937 -11969 24701 -11874
rect 24778 -11965 35398 -11874
rect 35475 -11886 37954 -11870
rect 35475 -11889 37847 -11886
rect 35475 -11894 37698 -11889
rect 35475 -11965 37539 -11894
rect 24778 -11969 37539 -11965
rect -69816 -11974 37539 -11969
rect -69965 -11977 37539 -11974
rect -70124 -11982 37539 -11977
rect -70936 -11989 37539 -11982
rect 37616 -11984 37698 -11894
rect 37775 -11981 37847 -11889
rect 37924 -11981 37954 -11886
rect 37775 -11984 37954 -11981
rect 37616 -11989 37954 -11984
rect -70936 -11999 37954 -11989
rect -70936 -12418 37954 -12390
rect -70936 -12421 24502 -12418
rect -70936 -12430 -56792 -12421
rect -70936 -12433 -70579 -12430
rect -70936 -12438 -70728 -12433
rect -70936 -12533 -70887 -12438
rect -70810 -12528 -70728 -12438
rect -70651 -12525 -70579 -12433
rect -70502 -12516 -56792 -12430
rect -56715 -12422 24502 -12421
rect -56715 -12516 -36403 -12422
rect -70502 -12517 -36403 -12516
rect -36326 -12517 -25303 -12422
rect -25226 -12517 -11291 -12422
rect -11214 -12517 2889 -12422
rect 2966 -12517 13652 -12422
rect 13729 -12513 24502 -12422
rect 24579 -12422 37954 -12418
rect 24579 -12513 35199 -12422
rect 13729 -12517 35199 -12513
rect 35276 -12432 37954 -12422
rect 35276 -12435 37163 -12432
rect 35276 -12440 37014 -12435
rect 35276 -12517 36855 -12440
rect -70502 -12525 36855 -12517
rect -70651 -12528 36855 -12525
rect -70810 -12533 36855 -12528
rect -70936 -12535 36855 -12533
rect 36932 -12530 37014 -12440
rect 37091 -12527 37163 -12435
rect 37240 -12527 37954 -12432
rect 37091 -12530 37954 -12527
rect 36932 -12535 37954 -12530
rect -70936 -12594 37954 -12535
rect -70936 -12597 24499 -12594
rect -70936 -12606 -56795 -12597
rect -70936 -12609 -70582 -12606
rect -70936 -12614 -70731 -12609
rect -70936 -12709 -70890 -12614
rect -70813 -12704 -70731 -12614
rect -70654 -12701 -70582 -12609
rect -70505 -12692 -56795 -12606
rect -56718 -12598 24499 -12597
rect -56718 -12692 -36406 -12598
rect -70505 -12693 -36406 -12692
rect -36329 -12693 -25306 -12598
rect -25229 -12693 -11294 -12598
rect -11217 -12693 2886 -12598
rect 2963 -12693 13649 -12598
rect 13726 -12689 24499 -12598
rect 24576 -12598 37954 -12594
rect 24576 -12689 35196 -12598
rect 13726 -12693 35196 -12689
rect 35273 -12608 37954 -12598
rect 35273 -12611 37160 -12608
rect 35273 -12616 37011 -12611
rect 35273 -12693 36852 -12616
rect -70505 -12701 36852 -12693
rect -70654 -12704 36852 -12701
rect -70813 -12709 36852 -12704
rect -70936 -12711 36852 -12709
rect 36929 -12706 37011 -12616
rect 37088 -12703 37160 -12611
rect 37237 -12703 37954 -12608
rect 37088 -12706 37954 -12703
rect 36929 -12711 37954 -12706
rect -70936 -12753 37954 -12711
rect -70936 -12756 24501 -12753
rect -70936 -12765 -56793 -12756
rect -70936 -12768 -70580 -12765
rect -70936 -12773 -70729 -12768
rect -70936 -12868 -70888 -12773
rect -70811 -12863 -70729 -12773
rect -70652 -12860 -70580 -12768
rect -70503 -12851 -56793 -12765
rect -56716 -12757 24501 -12756
rect -56716 -12851 -36404 -12757
rect -70503 -12852 -36404 -12851
rect -36327 -12852 -25304 -12757
rect -25227 -12852 -11292 -12757
rect -11215 -12852 2888 -12757
rect 2965 -12852 13651 -12757
rect 13728 -12848 24501 -12757
rect 24578 -12757 37954 -12753
rect 24578 -12848 35198 -12757
rect 13728 -12852 35198 -12848
rect 35275 -12767 37954 -12757
rect 35275 -12770 37162 -12767
rect 35275 -12775 37013 -12770
rect 35275 -12852 36854 -12775
rect -70503 -12860 36854 -12852
rect -70652 -12863 36854 -12860
rect -70811 -12868 36854 -12863
rect -70936 -12870 36854 -12868
rect 36931 -12865 37013 -12775
rect 37090 -12862 37162 -12770
rect 37239 -12862 37954 -12767
rect 37090 -12865 37954 -12862
rect 36931 -12870 37954 -12865
rect -70936 -12911 37954 -12870
rect -70936 -12914 24500 -12911
rect -70936 -12923 -56794 -12914
rect -70936 -12926 -70581 -12923
rect -70936 -12931 -70730 -12926
rect -70936 -13026 -70889 -12931
rect -70812 -13021 -70730 -12931
rect -70653 -13018 -70581 -12926
rect -70504 -13009 -56794 -12923
rect -56717 -12915 24500 -12914
rect -56717 -13009 -36405 -12915
rect -70504 -13010 -36405 -13009
rect -36328 -13010 -25305 -12915
rect -25228 -13010 -11293 -12915
rect -11216 -13010 2887 -12915
rect 2964 -13010 13650 -12915
rect 13727 -13006 24500 -12915
rect 24577 -12915 37954 -12911
rect 24577 -13006 35197 -12915
rect 13727 -13010 35197 -13006
rect 35274 -12925 37954 -12915
rect 35274 -12928 37161 -12925
rect 35274 -12933 37012 -12928
rect 35274 -13010 36853 -12933
rect -70504 -13018 36853 -13010
rect -70653 -13021 36853 -13018
rect -70812 -13026 36853 -13021
rect -70936 -13028 36853 -13026
rect 36930 -13023 37012 -12933
rect 37089 -13020 37161 -12928
rect 37238 -13020 37954 -12925
rect 37089 -13023 37954 -13020
rect 36930 -13028 37954 -13023
rect -70936 -13036 37954 -13028
rect -70903 -13039 -70496 -13036
rect 36835 -13038 37247 -13036
rect -3682 -14879 -3595 -14858
rect -63347 -14909 -63260 -14888
rect -63347 -14965 -63334 -14909
rect -63278 -14923 -63260 -14909
rect -63278 -14965 -17744 -14923
rect -63347 -14996 -17744 -14965
rect -63347 -15020 -31855 -14996
rect -63347 -15076 -63338 -15020
rect -63282 -15052 -31855 -15020
rect -31799 -15052 -17744 -14996
rect -63282 -15057 -17744 -15052
rect -3682 -14935 -3669 -14879
rect -3613 -14903 -3595 -14879
rect 7092 -14862 7179 -14841
rect 7092 -14903 7105 -14862
rect -3613 -14918 7105 -14903
rect 7161 -14903 7179 -14862
rect 17933 -14903 18020 -14889
rect 28638 -14903 28725 -14883
rect 7161 -14904 28725 -14903
rect 7161 -14910 28651 -14904
rect 7161 -14918 17946 -14910
rect -3613 -14935 17946 -14918
rect -3682 -14966 17946 -14935
rect 18002 -14960 28651 -14910
rect 28707 -14960 28725 -14904
rect 18002 -14966 28725 -14960
rect -3682 -14973 28725 -14966
rect -3682 -14990 7101 -14973
rect -3682 -15046 -3673 -14990
rect -3617 -15029 7101 -14990
rect 7157 -15015 28725 -14973
rect 7157 -15021 28647 -15015
rect 7157 -15029 17942 -15021
rect -3617 -15039 17942 -15029
rect -3617 -15046 -3595 -15039
rect 7092 -15044 7179 -15039
rect -63282 -15076 -63260 -15057
rect -63347 -15091 -63260 -15076
rect -43012 -15099 -42878 -15057
rect -43012 -15155 -42972 -15099
rect -42916 -15155 -42878 -15099
rect -43012 -15210 -42878 -15155
rect -31868 -15107 -31781 -15057
rect -31868 -15163 -31859 -15107
rect -31803 -15163 -31781 -15107
rect -31868 -15178 -31781 -15163
rect -17864 -15072 -17777 -15057
rect -3682 -15061 -3595 -15046
rect -17864 -15128 -17851 -15072
rect -17795 -15128 -17777 -15072
rect 17933 -15077 17942 -15039
rect 17998 -15039 28647 -15021
rect 17998 -15077 18020 -15039
rect 17933 -15092 18020 -15077
rect 28638 -15071 28647 -15039
rect 28703 -15071 28725 -15015
rect 28638 -15086 28725 -15071
rect -43012 -15266 -42976 -15210
rect -42920 -15266 -42878 -15210
rect -17864 -15183 -17777 -15128
rect -17864 -15239 -17855 -15183
rect -17799 -15239 -17777 -15183
rect -17864 -15254 -17777 -15239
rect -43012 -15303 -42878 -15266
rect -68398 -16634 -68278 -16601
rect -68398 -16749 -68375 -16634
rect -68295 -16749 -68278 -16634
rect -68398 -16891 -68278 -16749
rect -4046 -16754 -3896 -16730
rect -32218 -16809 -32087 -16789
rect -68398 -17006 -68377 -16891
rect -68297 -16901 -68278 -16891
rect -63669 -16879 -63582 -16858
rect -63669 -16901 -63656 -16879
rect -68297 -16935 -63656 -16901
rect -63600 -16901 -63582 -16879
rect -32218 -16887 -32183 -16809
rect -32114 -16887 -32087 -16809
rect -32218 -16901 -32087 -16887
rect -4046 -16819 -4002 -16754
rect -3932 -16819 -3896 -16754
rect -4046 -16829 -3896 -16819
rect 6633 -16765 6771 -16748
rect 6633 -16829 6667 -16765
rect -4046 -16836 6667 -16829
rect 6738 -16829 6771 -16765
rect 28305 -16761 28443 -16744
rect 17414 -16820 17552 -16803
rect 17414 -16829 17448 -16820
rect 6738 -16836 17448 -16829
rect -4046 -16891 17448 -16836
rect 17519 -16829 17552 -16820
rect 28305 -16829 28339 -16761
rect 17519 -16832 28339 -16829
rect 28410 -16829 28443 -16761
rect 28410 -16832 28501 -16829
rect 17519 -16891 28501 -16832
rect -63600 -16935 -18122 -16901
rect -68297 -16969 -18122 -16935
rect -68297 -16972 -18441 -16969
rect -68297 -16990 -43324 -16972
rect -68297 -17006 -63660 -16990
rect -68398 -17021 -63660 -17006
rect -63669 -17046 -63660 -17021
rect -63604 -17021 -43324 -16990
rect -63604 -17046 -63582 -17021
rect -63669 -17061 -63582 -17046
rect -43337 -17028 -43324 -17021
rect -43268 -16991 -18441 -16972
rect -43268 -17021 -32183 -16991
rect -43268 -17028 -43250 -17021
rect -43337 -17083 -43250 -17028
rect -32218 -17069 -32183 -17021
rect -32114 -17021 -18441 -16991
rect -32114 -17069 -32087 -17021
rect -32218 -17083 -32087 -17069
rect -18454 -17051 -18441 -17021
rect -18359 -17051 -18276 -16969
rect -18194 -17021 -18122 -16969
rect -4046 -16913 28501 -16891
rect -4046 -16978 -4008 -16913
rect -3938 -16937 28501 -16913
rect -3938 -16941 28335 -16937
rect -3938 -16964 6663 -16941
rect -3938 -16978 -3896 -16964
rect -4046 -16995 -3896 -16978
rect 6633 -17012 6663 -16964
rect 6734 -16964 28335 -16941
rect 6734 -17012 6771 -16964
rect -18194 -17051 -18169 -17021
rect 6633 -17022 6771 -17012
rect 17414 -16996 17552 -16964
rect -43337 -17139 -43328 -17083
rect -43272 -17139 -43250 -17083
rect -18454 -17089 -18169 -17051
rect 17414 -17067 17444 -16996
rect 17515 -17067 17552 -16996
rect 28305 -17008 28335 -16964
rect 28406 -16964 28501 -16937
rect 28406 -17008 28443 -16964
rect 28305 -17018 28443 -17008
rect 17414 -17077 17552 -17067
rect -43337 -17154 -43250 -17139
rect -36071 -19442 -35970 -19440
rect 24674 -19442 24775 -19440
rect -70936 -19466 37954 -19442
rect -70936 -19471 -36053 -19466
rect -70936 -19475 -46430 -19471
rect -70936 -19478 -69895 -19475
rect -70936 -19483 -70044 -19478
rect -70936 -19578 -70203 -19483
rect -70126 -19573 -70044 -19483
rect -69967 -19570 -69895 -19478
rect -69818 -19476 -46430 -19475
rect -69818 -19570 -56627 -19476
rect -69967 -19571 -56627 -19570
rect -56550 -19566 -46430 -19476
rect -46353 -19561 -36053 -19471
rect -35976 -19471 24692 -19466
rect -35976 -19561 -11142 -19471
rect -46353 -19566 -11142 -19561
rect -11065 -19566 13980 -19471
rect 14057 -19561 24692 -19471
rect 24769 -19471 37954 -19466
rect 24769 -19561 35416 -19471
rect 14057 -19566 35416 -19561
rect 35493 -19475 37954 -19471
rect 35493 -19478 37849 -19475
rect 35493 -19483 37700 -19478
rect 35493 -19566 37541 -19483
rect -56550 -19571 37541 -19566
rect -69967 -19573 37541 -19571
rect -70126 -19578 37541 -19573
rect 37618 -19573 37700 -19483
rect 37777 -19570 37849 -19478
rect 37926 -19570 37954 -19475
rect 37777 -19573 37954 -19570
rect 37618 -19578 37954 -19573
rect -70936 -19642 37954 -19578
rect -70936 -19647 -36056 -19642
rect -70936 -19651 -46433 -19647
rect -70936 -19654 -69898 -19651
rect -70936 -19659 -70047 -19654
rect -70936 -19754 -70206 -19659
rect -70129 -19749 -70047 -19659
rect -69970 -19746 -69898 -19654
rect -69821 -19652 -46433 -19651
rect -69821 -19746 -56630 -19652
rect -69970 -19747 -56630 -19746
rect -56553 -19742 -46433 -19652
rect -46356 -19737 -36056 -19647
rect -35979 -19647 24689 -19642
rect -35979 -19737 -11145 -19647
rect -46356 -19742 -11145 -19737
rect -11068 -19742 13977 -19647
rect 14054 -19737 24689 -19647
rect 24766 -19647 37954 -19642
rect 24766 -19737 35413 -19647
rect 14054 -19742 35413 -19737
rect 35490 -19651 37954 -19647
rect 35490 -19654 37846 -19651
rect 35490 -19659 37697 -19654
rect 35490 -19742 37538 -19659
rect -56553 -19747 37538 -19742
rect -69970 -19749 37538 -19747
rect -70129 -19754 37538 -19749
rect 37615 -19749 37697 -19659
rect 37774 -19746 37846 -19654
rect 37923 -19746 37954 -19651
rect 37774 -19749 37954 -19746
rect 37615 -19754 37954 -19749
rect -70936 -19801 37954 -19754
rect -70936 -19806 -36054 -19801
rect -70936 -19810 -46431 -19806
rect -70936 -19813 -69896 -19810
rect -70936 -19818 -70045 -19813
rect -70936 -19913 -70204 -19818
rect -70127 -19908 -70045 -19818
rect -69968 -19905 -69896 -19813
rect -69819 -19811 -46431 -19810
rect -69819 -19905 -56628 -19811
rect -69968 -19906 -56628 -19905
rect -56551 -19901 -46431 -19811
rect -46354 -19896 -36054 -19806
rect -35977 -19806 24691 -19801
rect -35977 -19896 -11143 -19806
rect -46354 -19901 -11143 -19896
rect -11066 -19901 13979 -19806
rect 14056 -19896 24691 -19806
rect 24768 -19806 37954 -19801
rect 24768 -19896 35415 -19806
rect 14056 -19901 35415 -19896
rect 35492 -19810 37954 -19806
rect 35492 -19813 37848 -19810
rect 35492 -19818 37699 -19813
rect 35492 -19901 37540 -19818
rect -56551 -19906 37540 -19901
rect -69968 -19908 37540 -19906
rect -70127 -19913 37540 -19908
rect 37617 -19908 37699 -19818
rect 37776 -19905 37848 -19813
rect 37925 -19905 37954 -19810
rect 37776 -19908 37954 -19905
rect 37617 -19913 37954 -19908
rect -70936 -19959 37954 -19913
rect -70936 -19964 -36055 -19959
rect -70936 -19968 -46432 -19964
rect -70936 -19971 -69897 -19968
rect -70936 -19976 -70046 -19971
rect -70936 -20071 -70205 -19976
rect -70128 -20066 -70046 -19976
rect -69969 -20063 -69897 -19971
rect -69820 -19969 -46432 -19968
rect -69820 -20063 -56629 -19969
rect -69969 -20064 -56629 -20063
rect -56552 -20059 -46432 -19969
rect -46355 -20054 -36055 -19964
rect -35978 -19964 24690 -19959
rect -35978 -20054 -11144 -19964
rect -46355 -20059 -11144 -20054
rect -11067 -20059 13978 -19964
rect 14055 -20054 24690 -19964
rect 24767 -19964 37954 -19959
rect 24767 -20054 35414 -19964
rect 14055 -20059 35414 -20054
rect 35491 -19968 37954 -19964
rect 35491 -19971 37847 -19968
rect 35491 -19976 37698 -19971
rect 35491 -20059 37539 -19976
rect -56552 -20064 37539 -20059
rect -69969 -20066 37539 -20064
rect -70128 -20071 37539 -20066
rect 37616 -20066 37698 -19976
rect 37775 -20063 37847 -19971
rect 37924 -20063 37954 -19968
rect 37775 -20066 37954 -20063
rect 37616 -20071 37954 -20066
rect -70936 -20088 37954 -20071
rect -70936 -20509 37954 -20479
rect -70936 -20513 -46636 -20509
rect -70936 -20515 -56831 -20513
rect -70936 -20518 -70587 -20515
rect -70936 -20523 -70736 -20518
rect -70936 -20618 -70895 -20523
rect -70818 -20613 -70736 -20523
rect -70659 -20610 -70587 -20518
rect -70510 -20608 -56831 -20515
rect -56754 -20604 -46636 -20513
rect -46559 -20513 37954 -20509
rect -46559 -20604 -36260 -20513
rect -56754 -20608 -36260 -20604
rect -36183 -20608 -11345 -20513
rect -11268 -20608 13778 -20513
rect 13855 -20608 24485 -20513
rect 24562 -20608 35213 -20513
rect 35290 -20515 37954 -20513
rect 35290 -20518 37159 -20515
rect 35290 -20523 37010 -20518
rect 35290 -20608 36851 -20523
rect -70510 -20610 36851 -20608
rect -70659 -20613 36851 -20610
rect -70818 -20618 36851 -20613
rect 36928 -20613 37010 -20523
rect 37087 -20610 37159 -20518
rect 37236 -20610 37954 -20515
rect 37087 -20613 37954 -20610
rect 36928 -20618 37954 -20613
rect -70936 -20685 37954 -20618
rect -70936 -20689 -46639 -20685
rect -70936 -20691 -56834 -20689
rect -70936 -20694 -70590 -20691
rect -70936 -20699 -70739 -20694
rect -70936 -20794 -70898 -20699
rect -70821 -20789 -70739 -20699
rect -70662 -20786 -70590 -20694
rect -70513 -20784 -56834 -20691
rect -56757 -20780 -46639 -20689
rect -46562 -20689 37954 -20685
rect -46562 -20780 -36263 -20689
rect -56757 -20784 -36263 -20780
rect -36186 -20784 -11348 -20689
rect -11271 -20784 13775 -20689
rect 13852 -20784 24482 -20689
rect 24559 -20784 35210 -20689
rect 35287 -20691 37954 -20689
rect 35287 -20694 37156 -20691
rect 35287 -20699 37007 -20694
rect 35287 -20784 36848 -20699
rect -70513 -20786 36848 -20784
rect -70662 -20789 36848 -20786
rect -70821 -20794 36848 -20789
rect 36925 -20789 37007 -20699
rect 37084 -20786 37156 -20694
rect 37233 -20786 37954 -20691
rect 37084 -20789 37954 -20786
rect 36925 -20794 37954 -20789
rect -70936 -20844 37954 -20794
rect -70936 -20848 -46637 -20844
rect -70936 -20850 -56832 -20848
rect -70936 -20853 -70588 -20850
rect -70936 -20858 -70737 -20853
rect -70936 -20953 -70896 -20858
rect -70819 -20948 -70737 -20858
rect -70660 -20945 -70588 -20853
rect -70511 -20943 -56832 -20850
rect -56755 -20939 -46637 -20848
rect -46560 -20848 37954 -20844
rect -46560 -20939 -36261 -20848
rect -56755 -20943 -36261 -20939
rect -36184 -20943 -11346 -20848
rect -11269 -20943 13777 -20848
rect 13854 -20943 24484 -20848
rect 24561 -20943 35212 -20848
rect 35289 -20850 37954 -20848
rect 35289 -20853 37158 -20850
rect 35289 -20858 37009 -20853
rect 35289 -20943 36850 -20858
rect -70511 -20945 36850 -20943
rect -70660 -20948 36850 -20945
rect -70819 -20953 36850 -20948
rect 36927 -20948 37009 -20858
rect 37086 -20945 37158 -20853
rect 37235 -20945 37954 -20850
rect 37086 -20948 37954 -20945
rect 36927 -20953 37954 -20948
rect -70936 -21002 37954 -20953
rect -70936 -21006 -46638 -21002
rect -70936 -21008 -56833 -21006
rect -70936 -21011 -70589 -21008
rect -70936 -21016 -70738 -21011
rect -70936 -21111 -70897 -21016
rect -70820 -21106 -70738 -21016
rect -70661 -21103 -70589 -21011
rect -70512 -21101 -56833 -21008
rect -56756 -21097 -46638 -21006
rect -46561 -21006 37954 -21002
rect -46561 -21097 -36262 -21006
rect -56756 -21101 -36262 -21097
rect -36185 -21101 -11347 -21006
rect -11270 -21101 13776 -21006
rect 13853 -21101 24483 -21006
rect 24560 -21101 35211 -21006
rect 35288 -21008 37954 -21006
rect 35288 -21011 37157 -21008
rect 35288 -21016 37008 -21011
rect 35288 -21101 36849 -21016
rect -70512 -21103 36849 -21101
rect -70661 -21106 36849 -21103
rect -70820 -21111 36849 -21106
rect 36926 -21106 37008 -21016
rect 37085 -21103 37157 -21011
rect 37234 -21103 37954 -21008
rect 37085 -21106 37954 -21103
rect 36926 -21111 37954 -21106
rect -70936 -21125 37954 -21111
rect -5312 -22845 -5178 -22802
rect -5312 -22926 -5294 -22845
rect -5194 -22926 -5178 -22845
rect -53204 -22980 -53117 -22959
rect -63396 -23010 -63309 -22991
rect -53204 -23010 -53191 -22980
rect -63396 -23012 -53191 -23010
rect -63396 -23068 -63383 -23012
rect -63327 -23036 -53191 -23012
rect -53135 -23010 -53117 -22980
rect -42813 -22989 -42726 -22968
rect -42813 -23010 -42800 -22989
rect -53135 -23036 -42800 -23010
rect -63327 -23045 -42800 -23036
rect -42744 -23010 -42726 -22989
rect -17905 -23001 -17818 -22980
rect -17905 -23010 -17892 -23001
rect -42744 -23045 -17892 -23010
rect -63327 -23057 -17892 -23045
rect -17836 -23010 -17818 -23001
rect -5312 -23010 -5178 -22926
rect -17836 -23046 -5178 -23010
rect -17836 -23057 -5295 -23046
rect -63327 -23068 -5295 -23057
rect -63396 -23091 -5295 -23068
rect -63396 -23123 -53195 -23091
rect -63396 -23179 -63387 -23123
rect -63331 -23144 -53195 -23123
rect -63331 -23179 -63309 -23144
rect -53204 -23147 -53195 -23144
rect -53139 -23100 -5295 -23091
rect -53139 -23144 -42804 -23100
rect -53139 -23147 -53117 -23144
rect -53204 -23162 -53117 -23147
rect -42813 -23156 -42804 -23144
rect -42748 -23112 -5295 -23100
rect -42748 -23144 -17896 -23112
rect -42748 -23156 -42726 -23144
rect -42813 -23171 -42726 -23156
rect -17905 -23168 -17896 -23144
rect -17840 -23127 -5295 -23112
rect -5195 -23127 -5178 -23046
rect -17840 -23144 -5178 -23127
rect -17840 -23168 -17818 -23144
rect -63396 -23194 -63309 -23179
rect -17905 -23183 -17818 -23168
rect -66896 -23417 -66488 -23396
rect -66896 -23497 -66855 -23417
rect -66759 -23497 -66488 -23417
rect -66896 -23547 -66488 -23497
rect -66639 -24975 -66488 -23547
rect -4953 -24701 -4802 -24665
rect -4953 -24811 -4927 -24701
rect -4830 -24811 -4802 -24701
rect -18293 -24854 -18140 -24841
rect -53561 -24909 -53410 -24883
rect -63739 -24952 -63652 -24931
rect -63739 -24975 -63726 -24952
rect -66639 -25008 -63726 -24975
rect -63670 -24975 -63652 -24952
rect -53561 -24971 -53526 -24909
rect -53467 -24971 -53410 -24909
rect -53561 -24975 -53410 -24971
rect -18293 -24936 -18255 -24854
rect -18173 -24936 -18140 -24854
rect -43355 -24975 -43028 -24974
rect -42701 -24975 -42445 -24973
rect -18293 -24975 -18140 -24936
rect -4953 -24975 -4802 -24811
rect 17320 -24908 17731 -24878
rect -63670 -24987 -4802 -24975
rect -63670 -25008 -4929 -24987
rect -66639 -25019 -4929 -25008
rect -66639 -25023 -18255 -25019
rect -66639 -25027 -42538 -25023
rect -66639 -25037 -42676 -25027
rect -66639 -25047 -43186 -25037
rect -66639 -25063 -53543 -25047
rect -66639 -25119 -63730 -25063
rect -63674 -25109 -53543 -25063
rect -53484 -25050 -43186 -25047
rect -53484 -25109 -43341 -25050
rect -63674 -25117 -43341 -25109
rect -43267 -25104 -43186 -25050
rect -43112 -25098 -42676 -25037
rect -42616 -25094 -42538 -25027
rect -42478 -25094 -18255 -25023
rect -42616 -25098 -18255 -25094
rect -43112 -25101 -18255 -25098
rect -18173 -25097 -4929 -25019
rect -4832 -25097 -4802 -24987
rect 6654 -24912 28480 -24908
rect 6654 -24937 28407 -24912
rect 6654 -24974 7446 -24937
rect 6654 -24990 6880 -24974
rect 6654 -25067 6666 -24990
rect 6734 -25051 6880 -24990
rect 6948 -24987 7446 -24974
rect 6948 -25051 7285 -24987
rect 6734 -25063 7285 -25051
rect 7353 -25013 7446 -24987
rect 7514 -24952 28407 -24937
rect 7514 -24962 17593 -24952
rect 7514 -25013 17338 -24962
rect 7353 -25055 17338 -25013
rect 17421 -25045 17593 -24962
rect 17676 -24969 28407 -24952
rect 28463 -24969 28480 -24912
rect 17676 -25015 28480 -24969
rect 17676 -25045 28314 -25015
rect 17421 -25055 28314 -25045
rect 7353 -25063 28314 -25055
rect 6734 -25067 28314 -25063
rect 6654 -25072 28314 -25067
rect 28370 -25072 28480 -25015
rect 6654 -25080 28480 -25072
rect -18173 -25101 -4802 -25097
rect -43112 -25104 -4802 -25101
rect -43267 -25117 -4802 -25104
rect -63674 -25119 -4802 -25117
rect -66639 -25126 -4802 -25119
rect 6656 -25121 6999 -25080
rect 17320 -25100 17731 -25080
rect 28308 -25084 28480 -25080
rect -70936 -27509 37954 -27482
rect -70936 -27513 -36007 -27509
rect -70936 -27523 -46396 -27513
rect -70936 -27526 -69895 -27523
rect -70936 -27531 -70044 -27526
rect -70936 -27626 -70203 -27531
rect -70126 -27621 -70044 -27531
rect -69967 -27618 -69895 -27526
rect -69818 -27608 -46396 -27523
rect -46319 -27604 -36007 -27513
rect -35930 -27513 37954 -27509
rect -35930 -27604 -11180 -27513
rect -46319 -27608 -11180 -27604
rect -11103 -27608 3174 -27513
rect 3251 -27608 24741 -27513
rect 24818 -27518 37954 -27513
rect 24818 -27521 37849 -27518
rect 24818 -27526 37700 -27521
rect 24818 -27608 37541 -27526
rect -69818 -27618 37541 -27608
rect -69967 -27621 37541 -27618
rect 37618 -27616 37700 -27526
rect 37777 -27613 37849 -27521
rect 37926 -27613 37954 -27518
rect 37777 -27616 37954 -27613
rect 37618 -27621 37954 -27616
rect -70126 -27626 37954 -27621
rect -70936 -27685 37954 -27626
rect -70936 -27689 -36010 -27685
rect -70936 -27699 -46399 -27689
rect -70936 -27702 -69898 -27699
rect -70936 -27707 -70047 -27702
rect -70936 -27802 -70206 -27707
rect -70129 -27797 -70047 -27707
rect -69970 -27794 -69898 -27702
rect -69821 -27784 -46399 -27699
rect -46322 -27780 -36010 -27689
rect -35933 -27689 37954 -27685
rect -35933 -27780 -11183 -27689
rect -46322 -27784 -11183 -27780
rect -11106 -27784 3171 -27689
rect 3248 -27784 24738 -27689
rect 24815 -27694 37954 -27689
rect 24815 -27697 37846 -27694
rect 24815 -27702 37697 -27697
rect 24815 -27784 37538 -27702
rect -69821 -27794 37538 -27784
rect -69970 -27797 37538 -27794
rect 37615 -27792 37697 -27702
rect 37774 -27789 37846 -27697
rect 37923 -27789 37954 -27694
rect 37774 -27792 37954 -27789
rect 37615 -27797 37954 -27792
rect -70129 -27802 37954 -27797
rect -70936 -27844 37954 -27802
rect -70936 -27848 -36008 -27844
rect -70936 -27858 -46397 -27848
rect -70936 -27861 -69896 -27858
rect -70936 -27866 -70045 -27861
rect -70936 -27961 -70204 -27866
rect -70127 -27956 -70045 -27866
rect -69968 -27953 -69896 -27861
rect -69819 -27943 -46397 -27858
rect -46320 -27939 -36008 -27848
rect -35931 -27848 37954 -27844
rect -35931 -27939 -11181 -27848
rect -46320 -27943 -11181 -27939
rect -11104 -27943 3173 -27848
rect 3250 -27943 24740 -27848
rect 24817 -27853 37954 -27848
rect 24817 -27856 37848 -27853
rect 24817 -27861 37699 -27856
rect 24817 -27943 37540 -27861
rect -69819 -27953 37540 -27943
rect -69968 -27956 37540 -27953
rect 37617 -27951 37699 -27861
rect 37776 -27948 37848 -27856
rect 37925 -27948 37954 -27853
rect 37776 -27951 37954 -27948
rect 37617 -27956 37954 -27951
rect -70127 -27961 37954 -27956
rect -70936 -28002 37954 -27961
rect -70936 -28006 -36009 -28002
rect -70936 -28016 -46398 -28006
rect -70936 -28019 -69897 -28016
rect -70936 -28024 -70046 -28019
rect -70936 -28119 -70205 -28024
rect -70128 -28114 -70046 -28024
rect -69969 -28111 -69897 -28019
rect -69820 -28101 -46398 -28016
rect -46321 -28097 -36009 -28006
rect -35932 -28006 37954 -28002
rect -35932 -28097 -11182 -28006
rect -46321 -28101 -11182 -28097
rect -11105 -28101 3172 -28006
rect 3249 -28101 24739 -28006
rect 24816 -28011 37954 -28006
rect 24816 -28014 37847 -28011
rect 24816 -28019 37698 -28014
rect 24816 -28101 37539 -28019
rect -69820 -28111 37539 -28101
rect -69969 -28114 37539 -28111
rect 37616 -28109 37698 -28019
rect 37775 -28106 37847 -28014
rect 37924 -28106 37954 -28011
rect 37775 -28109 37954 -28106
rect 37616 -28114 37954 -28109
rect -70128 -28119 37954 -28114
rect -70936 -28128 37954 -28119
rect -70219 -28132 -69812 -28128
rect -70936 -28551 37954 -28519
rect -70936 -28554 -36214 -28551
rect -70936 -28557 -70579 -28554
rect -70936 -28562 -70728 -28557
rect -70936 -28657 -70887 -28562
rect -70810 -28652 -70728 -28562
rect -70651 -28649 -70579 -28557
rect -70502 -28555 -36214 -28554
rect -70502 -28649 -46607 -28555
rect -70651 -28650 -46607 -28649
rect -46530 -28646 -36214 -28555
rect -36137 -28646 -11386 -28551
rect -11309 -28554 37954 -28551
rect -11309 -28555 37167 -28554
rect -11309 -28646 2980 -28555
rect -46530 -28650 2980 -28646
rect 3057 -28650 24539 -28555
rect 24616 -28557 37167 -28555
rect 24616 -28562 37018 -28557
rect 24616 -28650 36859 -28562
rect -70651 -28652 36859 -28650
rect -70810 -28657 36859 -28652
rect 36936 -28652 37018 -28562
rect 37095 -28649 37167 -28557
rect 37244 -28649 37954 -28554
rect 37095 -28652 37954 -28649
rect 36936 -28657 37954 -28652
rect -70936 -28727 37954 -28657
rect -70936 -28730 -36217 -28727
rect -70936 -28733 -70582 -28730
rect -70936 -28738 -70731 -28733
rect -70936 -28833 -70890 -28738
rect -70813 -28828 -70731 -28738
rect -70654 -28825 -70582 -28733
rect -70505 -28731 -36217 -28730
rect -70505 -28825 -46610 -28731
rect -70654 -28826 -46610 -28825
rect -46533 -28822 -36217 -28731
rect -36140 -28822 -11389 -28727
rect -11312 -28730 37954 -28727
rect -11312 -28731 37164 -28730
rect -11312 -28822 2977 -28731
rect -46533 -28826 2977 -28822
rect 3054 -28826 24536 -28731
rect 24613 -28733 37164 -28731
rect 24613 -28738 37015 -28733
rect 24613 -28826 36856 -28738
rect -70654 -28828 36856 -28826
rect -70813 -28833 36856 -28828
rect 36933 -28828 37015 -28738
rect 37092 -28825 37164 -28733
rect 37241 -28825 37954 -28730
rect 37092 -28828 37954 -28825
rect 36933 -28833 37954 -28828
rect -70936 -28886 37954 -28833
rect -70936 -28889 -36215 -28886
rect -70936 -28892 -70580 -28889
rect -70936 -28897 -70729 -28892
rect -70936 -28992 -70888 -28897
rect -70811 -28987 -70729 -28897
rect -70652 -28984 -70580 -28892
rect -70503 -28890 -36215 -28889
rect -70503 -28984 -46608 -28890
rect -70652 -28985 -46608 -28984
rect -46531 -28981 -36215 -28890
rect -36138 -28981 -11387 -28886
rect -11310 -28889 37954 -28886
rect -11310 -28890 37166 -28889
rect -11310 -28981 2979 -28890
rect -46531 -28985 2979 -28981
rect 3056 -28985 24538 -28890
rect 24615 -28892 37166 -28890
rect 24615 -28897 37017 -28892
rect 24615 -28985 36858 -28897
rect -70652 -28987 36858 -28985
rect -70811 -28992 36858 -28987
rect 36935 -28987 37017 -28897
rect 37094 -28984 37166 -28892
rect 37243 -28984 37954 -28889
rect 37094 -28987 37954 -28984
rect 36935 -28992 37954 -28987
rect -70936 -29044 37954 -28992
rect -70936 -29047 -36216 -29044
rect -70936 -29050 -70581 -29047
rect -70936 -29055 -70730 -29050
rect -70936 -29150 -70889 -29055
rect -70812 -29145 -70730 -29055
rect -70653 -29142 -70581 -29050
rect -70504 -29048 -36216 -29047
rect -70504 -29142 -46609 -29048
rect -70653 -29143 -46609 -29142
rect -46532 -29139 -36216 -29048
rect -36139 -29139 -11388 -29044
rect -11311 -29047 37954 -29044
rect -11311 -29048 37165 -29047
rect -11311 -29139 2978 -29048
rect -46532 -29143 2978 -29139
rect 3055 -29143 24537 -29048
rect 24614 -29050 37165 -29048
rect 24614 -29055 37016 -29050
rect 24614 -29143 36857 -29055
rect -70653 -29145 36857 -29143
rect -70812 -29150 36857 -29145
rect 36934 -29145 37016 -29055
rect 37093 -29142 37165 -29050
rect 37242 -29142 37954 -29047
rect 37093 -29145 37954 -29142
rect 36934 -29150 37954 -29145
rect -70936 -29165 37954 -29150
rect -46625 -29166 -46524 -29165
rect 2962 -29166 3063 -29165
rect 24521 -29166 24622 -29165
rect -56388 -32893 -56253 -32836
rect -56388 -32969 -56365 -32893
rect -56276 -32969 -56253 -32893
rect -56388 -33046 -56253 -32969
rect -53649 -33046 -53369 -33030
rect -53224 -33046 -53089 -33045
rect -18454 -33046 -18146 -33026
rect 17512 -33046 17772 -33037
rect -56388 -33079 17772 -33046
rect -56388 -33081 -18259 -33079
rect -56388 -33084 -18438 -33081
rect -56388 -33160 -56370 -33084
rect -56281 -33085 -18438 -33084
rect -56281 -33160 -53633 -33085
rect -56388 -33163 -53633 -33160
rect -53555 -33163 -53468 -33085
rect -53390 -33088 -43020 -33085
rect -53390 -33147 -43133 -33088
rect -43077 -33144 -43020 -33088
rect -42964 -33144 -18438 -33085
rect -43077 -33147 -18438 -33144
rect -53390 -33149 -18438 -33147
rect -18377 -33147 -18259 -33081
rect -18198 -33091 17772 -33079
rect -18198 -33092 17683 -33091
rect -18198 -33114 -3968 -33092
rect -18198 -33147 -4122 -33114
rect -18377 -33149 -4122 -33147
rect -53390 -33163 -4122 -33149
rect -56388 -33175 -4122 -33163
rect -4054 -33153 -3968 -33114
rect -3900 -33093 17683 -33092
rect -3900 -33153 17525 -33093
rect -4054 -33157 17525 -33153
rect 17583 -33155 17683 -33093
rect 17741 -33155 17772 -33091
rect 17583 -33157 17772 -33155
rect -4054 -33175 17772 -33157
rect -56388 -33181 17772 -33175
rect -53649 -33213 -53369 -33181
rect -4136 -33200 -3864 -33181
rect 17512 -33184 17772 -33181
rect -70936 -36510 37954 -36480
rect -70936 -36513 -54969 -36510
rect -70936 -36518 -55118 -36513
rect -70936 -36521 -55277 -36518
rect -70936 -36524 -65367 -36521
rect -70936 -36529 -65516 -36524
rect -70936 -36624 -65675 -36529
rect -65598 -36619 -65516 -36529
rect -65439 -36616 -65367 -36524
rect -65290 -36613 -55277 -36521
rect -55200 -36608 -55118 -36518
rect -55041 -36605 -54969 -36513
rect -54892 -36513 37954 -36510
rect -54892 -36516 -34373 -36513
rect -54892 -36517 -34522 -36516
rect -54892 -36520 -44612 -36517
rect -54892 -36525 -44761 -36520
rect -54892 -36605 -44920 -36525
rect -55041 -36608 -44920 -36605
rect -55200 -36613 -44920 -36608
rect -65290 -36616 -44920 -36613
rect -65439 -36619 -44920 -36616
rect -65598 -36620 -44920 -36619
rect -44843 -36615 -44761 -36525
rect -44684 -36612 -44612 -36520
rect -44535 -36521 -34522 -36517
rect -44535 -36612 -34681 -36521
rect -44684 -36615 -34681 -36612
rect -44843 -36616 -34681 -36615
rect -34604 -36611 -34522 -36521
rect -34445 -36608 -34373 -36516
rect -34296 -36517 37954 -36513
rect -34296 -36520 -23073 -36517
rect -34296 -36525 -23222 -36520
rect -34296 -36608 -23381 -36525
rect -34445 -36611 -23381 -36608
rect -34604 -36616 -23381 -36611
rect -44843 -36620 -23381 -36616
rect -23304 -36615 -23222 -36525
rect -23145 -36612 -23073 -36520
rect -22996 -36520 -6817 -36517
rect -22996 -36525 -6966 -36520
rect -22996 -36612 -7125 -36525
rect -23145 -36615 -7125 -36612
rect -23304 -36620 -7125 -36615
rect -7048 -36615 -6966 -36525
rect -6889 -36612 -6817 -36520
rect -6740 -36520 5160 -36517
rect -6740 -36525 5011 -36520
rect -6740 -36612 4852 -36525
rect -6889 -36615 4852 -36612
rect -7048 -36620 4852 -36615
rect 4929 -36615 5011 -36525
rect 5088 -36612 5160 -36520
rect 5237 -36520 15643 -36517
rect 5237 -36525 15494 -36520
rect 5237 -36612 15335 -36525
rect 5088 -36615 15335 -36612
rect 4929 -36620 15335 -36615
rect 15412 -36615 15494 -36525
rect 15571 -36612 15643 -36520
rect 15720 -36520 26348 -36517
rect 15720 -36525 26199 -36520
rect 15720 -36612 26040 -36525
rect 15571 -36615 26040 -36612
rect 15412 -36620 26040 -36615
rect 26117 -36615 26199 -36525
rect 26276 -36612 26348 -36520
rect 26425 -36612 37954 -36517
rect 26276 -36615 37954 -36612
rect 26117 -36620 37954 -36615
rect -65598 -36624 37954 -36620
rect -70936 -36686 37954 -36624
rect -70936 -36689 -54972 -36686
rect -70936 -36694 -55121 -36689
rect -70936 -36697 -55280 -36694
rect -70936 -36700 -65370 -36697
rect -70936 -36705 -65519 -36700
rect -70936 -36800 -65678 -36705
rect -65601 -36795 -65519 -36705
rect -65442 -36792 -65370 -36700
rect -65293 -36789 -55280 -36697
rect -55203 -36784 -55121 -36694
rect -55044 -36781 -54972 -36689
rect -54895 -36689 37954 -36686
rect -54895 -36692 -34376 -36689
rect -54895 -36693 -34525 -36692
rect -54895 -36696 -44615 -36693
rect -54895 -36701 -44764 -36696
rect -54895 -36781 -44923 -36701
rect -55044 -36784 -44923 -36781
rect -55203 -36789 -44923 -36784
rect -65293 -36792 -44923 -36789
rect -65442 -36795 -44923 -36792
rect -65601 -36796 -44923 -36795
rect -44846 -36791 -44764 -36701
rect -44687 -36788 -44615 -36696
rect -44538 -36697 -34525 -36693
rect -44538 -36788 -34684 -36697
rect -44687 -36791 -34684 -36788
rect -44846 -36792 -34684 -36791
rect -34607 -36787 -34525 -36697
rect -34448 -36784 -34376 -36692
rect -34299 -36693 37954 -36689
rect -34299 -36696 -23076 -36693
rect -34299 -36701 -23225 -36696
rect -34299 -36784 -23384 -36701
rect -34448 -36787 -23384 -36784
rect -34607 -36792 -23384 -36787
rect -44846 -36796 -23384 -36792
rect -23307 -36791 -23225 -36701
rect -23148 -36788 -23076 -36696
rect -22999 -36696 -6820 -36693
rect -22999 -36701 -6969 -36696
rect -22999 -36788 -7128 -36701
rect -23148 -36791 -7128 -36788
rect -23307 -36796 -7128 -36791
rect -7051 -36791 -6969 -36701
rect -6892 -36788 -6820 -36696
rect -6743 -36696 5157 -36693
rect -6743 -36701 5008 -36696
rect -6743 -36788 4849 -36701
rect -6892 -36791 4849 -36788
rect -7051 -36796 4849 -36791
rect 4926 -36791 5008 -36701
rect 5085 -36788 5157 -36696
rect 5234 -36696 15640 -36693
rect 5234 -36701 15491 -36696
rect 5234 -36788 15332 -36701
rect 5085 -36791 15332 -36788
rect 4926 -36796 15332 -36791
rect 15409 -36791 15491 -36701
rect 15568 -36788 15640 -36696
rect 15717 -36696 26345 -36693
rect 15717 -36701 26196 -36696
rect 15717 -36788 26037 -36701
rect 15568 -36791 26037 -36788
rect 15409 -36796 26037 -36791
rect 26114 -36791 26196 -36701
rect 26273 -36788 26345 -36696
rect 26422 -36788 37954 -36693
rect 26273 -36791 37954 -36788
rect 26114 -36796 37954 -36791
rect -65601 -36800 37954 -36796
rect -70936 -36845 37954 -36800
rect -70936 -36848 -54970 -36845
rect -70936 -36853 -55119 -36848
rect -70936 -36856 -55278 -36853
rect -70936 -36859 -65368 -36856
rect -70936 -36864 -65517 -36859
rect -70936 -36959 -65676 -36864
rect -65599 -36954 -65517 -36864
rect -65440 -36951 -65368 -36859
rect -65291 -36948 -55278 -36856
rect -55201 -36943 -55119 -36853
rect -55042 -36940 -54970 -36848
rect -54893 -36848 37954 -36845
rect -54893 -36851 -34374 -36848
rect -54893 -36852 -34523 -36851
rect -54893 -36855 -44613 -36852
rect -54893 -36860 -44762 -36855
rect -54893 -36940 -44921 -36860
rect -55042 -36943 -44921 -36940
rect -55201 -36948 -44921 -36943
rect -65291 -36951 -44921 -36948
rect -65440 -36954 -44921 -36951
rect -65599 -36955 -44921 -36954
rect -44844 -36950 -44762 -36860
rect -44685 -36947 -44613 -36855
rect -44536 -36856 -34523 -36852
rect -44536 -36947 -34682 -36856
rect -44685 -36950 -34682 -36947
rect -44844 -36951 -34682 -36950
rect -34605 -36946 -34523 -36856
rect -34446 -36943 -34374 -36851
rect -34297 -36852 37954 -36848
rect -34297 -36855 -23074 -36852
rect -34297 -36860 -23223 -36855
rect -34297 -36943 -23382 -36860
rect -34446 -36946 -23382 -36943
rect -34605 -36951 -23382 -36946
rect -44844 -36955 -23382 -36951
rect -23305 -36950 -23223 -36860
rect -23146 -36947 -23074 -36855
rect -22997 -36855 -6818 -36852
rect -22997 -36860 -6967 -36855
rect -22997 -36947 -7126 -36860
rect -23146 -36950 -7126 -36947
rect -23305 -36955 -7126 -36950
rect -7049 -36950 -6967 -36860
rect -6890 -36947 -6818 -36855
rect -6741 -36855 5159 -36852
rect -6741 -36860 5010 -36855
rect -6741 -36947 4851 -36860
rect -6890 -36950 4851 -36947
rect -7049 -36955 4851 -36950
rect 4928 -36950 5010 -36860
rect 5087 -36947 5159 -36855
rect 5236 -36855 15642 -36852
rect 5236 -36860 15493 -36855
rect 5236 -36947 15334 -36860
rect 5087 -36950 15334 -36947
rect 4928 -36955 15334 -36950
rect 15411 -36950 15493 -36860
rect 15570 -36947 15642 -36855
rect 15719 -36855 26347 -36852
rect 15719 -36860 26198 -36855
rect 15719 -36947 26039 -36860
rect 15570 -36950 26039 -36947
rect 15411 -36955 26039 -36950
rect 26116 -36950 26198 -36860
rect 26275 -36947 26347 -36855
rect 26424 -36947 37954 -36852
rect 26275 -36950 37954 -36947
rect 26116 -36955 37954 -36950
rect -65599 -36959 37954 -36955
rect -70936 -37003 37954 -36959
rect -70936 -37006 -54971 -37003
rect -70936 -37011 -55120 -37006
rect -70936 -37014 -55279 -37011
rect -70936 -37017 -65369 -37014
rect -70936 -37022 -65518 -37017
rect -70936 -37117 -65677 -37022
rect -65600 -37112 -65518 -37022
rect -65441 -37109 -65369 -37017
rect -65292 -37106 -55279 -37014
rect -55202 -37101 -55120 -37011
rect -55043 -37098 -54971 -37006
rect -54894 -37006 37954 -37003
rect -54894 -37009 -34375 -37006
rect -54894 -37010 -34524 -37009
rect -54894 -37013 -44614 -37010
rect -54894 -37018 -44763 -37013
rect -54894 -37098 -44922 -37018
rect -55043 -37101 -44922 -37098
rect -55202 -37106 -44922 -37101
rect -65292 -37109 -44922 -37106
rect -65441 -37112 -44922 -37109
rect -65600 -37113 -44922 -37112
rect -44845 -37108 -44763 -37018
rect -44686 -37105 -44614 -37013
rect -44537 -37014 -34524 -37010
rect -44537 -37105 -34683 -37014
rect -44686 -37108 -34683 -37105
rect -44845 -37109 -34683 -37108
rect -34606 -37104 -34524 -37014
rect -34447 -37101 -34375 -37009
rect -34298 -37010 37954 -37006
rect -34298 -37013 -23075 -37010
rect -34298 -37018 -23224 -37013
rect -34298 -37101 -23383 -37018
rect -34447 -37104 -23383 -37101
rect -34606 -37109 -23383 -37104
rect -44845 -37113 -23383 -37109
rect -23306 -37108 -23224 -37018
rect -23147 -37105 -23075 -37013
rect -22998 -37013 -6819 -37010
rect -22998 -37018 -6968 -37013
rect -22998 -37105 -7127 -37018
rect -23147 -37108 -7127 -37105
rect -23306 -37113 -7127 -37108
rect -7050 -37108 -6968 -37018
rect -6891 -37105 -6819 -37013
rect -6742 -37013 5158 -37010
rect -6742 -37018 5009 -37013
rect -6742 -37105 4850 -37018
rect -6891 -37108 4850 -37105
rect -7050 -37113 4850 -37108
rect 4927 -37108 5009 -37018
rect 5086 -37105 5158 -37013
rect 5235 -37013 15641 -37010
rect 5235 -37018 15492 -37013
rect 5235 -37105 15333 -37018
rect 5086 -37108 15333 -37105
rect 4927 -37113 15333 -37108
rect 15410 -37108 15492 -37018
rect 15569 -37105 15641 -37013
rect 15718 -37013 26346 -37010
rect 15718 -37018 26197 -37013
rect 15718 -37105 26038 -37018
rect 15569 -37108 26038 -37105
rect 15410 -37113 26038 -37108
rect 26115 -37108 26197 -37018
rect 26274 -37105 26346 -37013
rect 26423 -37105 37954 -37010
rect 26274 -37108 37954 -37105
rect 26115 -37113 37954 -37108
rect -65600 -37117 37954 -37113
rect -70936 -37126 37954 -37117
rect -65694 -37129 -65284 -37126
rect -70936 -37549 37954 -37517
rect -70936 -37552 -23862 -37549
rect -70936 -37553 -24011 -37552
rect -70936 -37556 -66063 -37553
rect -70936 -37561 -66212 -37556
rect -70936 -37656 -66371 -37561
rect -66294 -37651 -66212 -37561
rect -66135 -37648 -66063 -37556
rect -65986 -37556 -24011 -37553
rect -65986 -37559 -55611 -37556
rect -65986 -37564 -55760 -37559
rect -65986 -37648 -55919 -37564
rect -66135 -37651 -55919 -37648
rect -66294 -37656 -55919 -37651
rect -70936 -37659 -55919 -37656
rect -55842 -37654 -55760 -37564
rect -55683 -37651 -55611 -37559
rect -55534 -37559 -45434 -37556
rect -55534 -37564 -45583 -37559
rect -55534 -37651 -45742 -37564
rect -55683 -37654 -45742 -37651
rect -55842 -37659 -45742 -37654
rect -45665 -37654 -45583 -37564
rect -45506 -37651 -45434 -37559
rect -45357 -37557 -24011 -37556
rect -45357 -37560 -24170 -37557
rect -45357 -37563 -35063 -37560
rect -45357 -37568 -35212 -37563
rect -45357 -37651 -35371 -37568
rect -45506 -37654 -35371 -37651
rect -45665 -37659 -35371 -37654
rect -70936 -37663 -35371 -37659
rect -35294 -37658 -35212 -37568
rect -35135 -37655 -35063 -37563
rect -34986 -37652 -24170 -37560
rect -24093 -37647 -24011 -37557
rect -23934 -37644 -23862 -37552
rect -23785 -37550 37954 -37549
rect -23785 -37553 25661 -37550
rect -23785 -37556 -7588 -37553
rect -23785 -37561 -7737 -37556
rect -23785 -37644 -7896 -37561
rect -23934 -37647 -7896 -37644
rect -24093 -37652 -7896 -37647
rect -34986 -37655 -7896 -37652
rect -35135 -37656 -7896 -37655
rect -7819 -37651 -7737 -37561
rect -7660 -37648 -7588 -37556
rect -7511 -37556 4397 -37553
rect -7511 -37561 4248 -37556
rect -7511 -37648 4089 -37561
rect -7660 -37651 4089 -37648
rect -7819 -37656 4089 -37651
rect 4166 -37651 4248 -37561
rect 4325 -37648 4397 -37556
rect 4474 -37558 25512 -37553
rect 4474 -37561 25353 -37558
rect 4474 -37564 14957 -37561
rect 4474 -37569 14808 -37564
rect 4474 -37648 14649 -37569
rect 4325 -37651 14649 -37648
rect 4166 -37656 14649 -37651
rect -35135 -37658 14649 -37656
rect -35294 -37663 14649 -37658
rect -70936 -37664 14649 -37663
rect 14726 -37659 14808 -37569
rect 14885 -37656 14957 -37564
rect 15034 -37653 25353 -37561
rect 25430 -37648 25512 -37558
rect 25589 -37645 25661 -37553
rect 25738 -37645 37954 -37550
rect 25589 -37648 37954 -37645
rect 25430 -37653 37954 -37648
rect 15034 -37656 37954 -37653
rect 14885 -37659 37954 -37656
rect 14726 -37664 37954 -37659
rect -70936 -37725 37954 -37664
rect -70936 -37728 -23865 -37725
rect -70936 -37729 -24014 -37728
rect -70936 -37732 -66066 -37729
rect -70936 -37737 -66215 -37732
rect -70936 -37832 -66374 -37737
rect -66297 -37827 -66215 -37737
rect -66138 -37824 -66066 -37732
rect -65989 -37732 -24014 -37729
rect -65989 -37735 -55614 -37732
rect -65989 -37740 -55763 -37735
rect -65989 -37824 -55922 -37740
rect -66138 -37827 -55922 -37824
rect -66297 -37832 -55922 -37827
rect -70936 -37835 -55922 -37832
rect -55845 -37830 -55763 -37740
rect -55686 -37827 -55614 -37735
rect -55537 -37735 -45437 -37732
rect -55537 -37740 -45586 -37735
rect -55537 -37827 -45745 -37740
rect -55686 -37830 -45745 -37827
rect -55845 -37835 -45745 -37830
rect -45668 -37830 -45586 -37740
rect -45509 -37827 -45437 -37735
rect -45360 -37733 -24014 -37732
rect -45360 -37736 -24173 -37733
rect -45360 -37739 -35066 -37736
rect -45360 -37744 -35215 -37739
rect -45360 -37827 -35374 -37744
rect -45509 -37830 -35374 -37827
rect -45668 -37835 -35374 -37830
rect -70936 -37839 -35374 -37835
rect -35297 -37834 -35215 -37744
rect -35138 -37831 -35066 -37739
rect -34989 -37828 -24173 -37736
rect -24096 -37823 -24014 -37733
rect -23937 -37820 -23865 -37728
rect -23788 -37726 37954 -37725
rect -23788 -37729 25658 -37726
rect -23788 -37732 -7591 -37729
rect -23788 -37737 -7740 -37732
rect -23788 -37820 -7899 -37737
rect -23937 -37823 -7899 -37820
rect -24096 -37828 -7899 -37823
rect -34989 -37831 -7899 -37828
rect -35138 -37832 -7899 -37831
rect -7822 -37827 -7740 -37737
rect -7663 -37824 -7591 -37732
rect -7514 -37732 4394 -37729
rect -7514 -37737 4245 -37732
rect -7514 -37824 4086 -37737
rect -7663 -37827 4086 -37824
rect -7822 -37832 4086 -37827
rect 4163 -37827 4245 -37737
rect 4322 -37824 4394 -37732
rect 4471 -37734 25509 -37729
rect 4471 -37737 25350 -37734
rect 4471 -37740 14954 -37737
rect 4471 -37745 14805 -37740
rect 4471 -37824 14646 -37745
rect 4322 -37827 14646 -37824
rect 4163 -37832 14646 -37827
rect -35138 -37834 14646 -37832
rect -35297 -37839 14646 -37834
rect -70936 -37840 14646 -37839
rect 14723 -37835 14805 -37745
rect 14882 -37832 14954 -37740
rect 15031 -37829 25350 -37737
rect 25427 -37824 25509 -37734
rect 25586 -37821 25658 -37729
rect 25735 -37821 37954 -37726
rect 25586 -37824 37954 -37821
rect 25427 -37829 37954 -37824
rect 15031 -37832 37954 -37829
rect 14882 -37835 37954 -37832
rect 14723 -37840 37954 -37835
rect -70936 -37884 37954 -37840
rect -70936 -37887 -23863 -37884
rect -70936 -37888 -24012 -37887
rect -70936 -37891 -66064 -37888
rect -70936 -37896 -66213 -37891
rect -70936 -37991 -66372 -37896
rect -66295 -37986 -66213 -37896
rect -66136 -37983 -66064 -37891
rect -65987 -37891 -24012 -37888
rect -65987 -37894 -55612 -37891
rect -65987 -37899 -55761 -37894
rect -65987 -37983 -55920 -37899
rect -66136 -37986 -55920 -37983
rect -66295 -37991 -55920 -37986
rect -70936 -37994 -55920 -37991
rect -55843 -37989 -55761 -37899
rect -55684 -37986 -55612 -37894
rect -55535 -37894 -45435 -37891
rect -55535 -37899 -45584 -37894
rect -55535 -37986 -45743 -37899
rect -55684 -37989 -45743 -37986
rect -55843 -37994 -45743 -37989
rect -45666 -37989 -45584 -37899
rect -45507 -37986 -45435 -37894
rect -45358 -37892 -24012 -37891
rect -45358 -37895 -24171 -37892
rect -45358 -37898 -35064 -37895
rect -45358 -37903 -35213 -37898
rect -45358 -37986 -35372 -37903
rect -45507 -37989 -35372 -37986
rect -45666 -37994 -35372 -37989
rect -70936 -37998 -35372 -37994
rect -35295 -37993 -35213 -37903
rect -35136 -37990 -35064 -37898
rect -34987 -37987 -24171 -37895
rect -24094 -37982 -24012 -37892
rect -23935 -37979 -23863 -37887
rect -23786 -37885 37954 -37884
rect -23786 -37888 25660 -37885
rect -23786 -37891 -7589 -37888
rect -23786 -37896 -7738 -37891
rect -23786 -37979 -7897 -37896
rect -23935 -37982 -7897 -37979
rect -24094 -37987 -7897 -37982
rect -34987 -37990 -7897 -37987
rect -35136 -37991 -7897 -37990
rect -7820 -37986 -7738 -37896
rect -7661 -37983 -7589 -37891
rect -7512 -37891 4396 -37888
rect -7512 -37896 4247 -37891
rect -7512 -37983 4088 -37896
rect -7661 -37986 4088 -37983
rect -7820 -37991 4088 -37986
rect 4165 -37986 4247 -37896
rect 4324 -37983 4396 -37891
rect 4473 -37893 25511 -37888
rect 4473 -37896 25352 -37893
rect 4473 -37899 14956 -37896
rect 4473 -37904 14807 -37899
rect 4473 -37983 14648 -37904
rect 4324 -37986 14648 -37983
rect 4165 -37991 14648 -37986
rect -35136 -37993 14648 -37991
rect -35295 -37998 14648 -37993
rect -70936 -37999 14648 -37998
rect 14725 -37994 14807 -37904
rect 14884 -37991 14956 -37899
rect 15033 -37988 25352 -37896
rect 25429 -37983 25511 -37893
rect 25588 -37980 25660 -37888
rect 25737 -37980 37954 -37885
rect 25588 -37983 37954 -37980
rect 25429 -37988 37954 -37983
rect 15033 -37991 37954 -37988
rect 14884 -37994 37954 -37991
rect 14725 -37999 37954 -37994
rect -70936 -38042 37954 -37999
rect -70936 -38045 -23864 -38042
rect -70936 -38046 -24013 -38045
rect -70936 -38049 -66065 -38046
rect -70936 -38054 -66214 -38049
rect -70936 -38149 -66373 -38054
rect -66296 -38144 -66214 -38054
rect -66137 -38141 -66065 -38049
rect -65988 -38049 -24013 -38046
rect -65988 -38052 -55613 -38049
rect -65988 -38057 -55762 -38052
rect -65988 -38141 -55921 -38057
rect -66137 -38144 -55921 -38141
rect -66296 -38149 -55921 -38144
rect -70936 -38152 -55921 -38149
rect -55844 -38147 -55762 -38057
rect -55685 -38144 -55613 -38052
rect -55536 -38052 -45436 -38049
rect -55536 -38057 -45585 -38052
rect -55536 -38144 -45744 -38057
rect -55685 -38147 -45744 -38144
rect -55844 -38152 -45744 -38147
rect -45667 -38147 -45585 -38057
rect -45508 -38144 -45436 -38052
rect -45359 -38050 -24013 -38049
rect -45359 -38053 -24172 -38050
rect -45359 -38056 -35065 -38053
rect -45359 -38061 -35214 -38056
rect -45359 -38144 -35373 -38061
rect -45508 -38147 -35373 -38144
rect -45667 -38152 -35373 -38147
rect -70936 -38156 -35373 -38152
rect -35296 -38151 -35214 -38061
rect -35137 -38148 -35065 -38056
rect -34988 -38145 -24172 -38053
rect -24095 -38140 -24013 -38050
rect -23936 -38137 -23864 -38045
rect -23787 -38043 37954 -38042
rect -23787 -38046 25659 -38043
rect -23787 -38049 -7590 -38046
rect -23787 -38054 -7739 -38049
rect -23787 -38137 -7898 -38054
rect -23936 -38140 -7898 -38137
rect -24095 -38145 -7898 -38140
rect -34988 -38148 -7898 -38145
rect -35137 -38149 -7898 -38148
rect -7821 -38144 -7739 -38054
rect -7662 -38141 -7590 -38049
rect -7513 -38049 4395 -38046
rect -7513 -38054 4246 -38049
rect -7513 -38141 4087 -38054
rect -7662 -38144 4087 -38141
rect -7821 -38149 4087 -38144
rect 4164 -38144 4246 -38054
rect 4323 -38141 4395 -38049
rect 4472 -38051 25510 -38046
rect 4472 -38054 25351 -38051
rect 4472 -38057 14955 -38054
rect 4472 -38062 14806 -38057
rect 4472 -38141 14647 -38062
rect 4323 -38144 14647 -38141
rect 4164 -38149 14647 -38144
rect -35137 -38151 14647 -38149
rect -35296 -38156 14647 -38151
rect -70936 -38157 14647 -38156
rect 14724 -38152 14806 -38062
rect 14883 -38149 14955 -38057
rect 15032 -38146 25351 -38054
rect 25428 -38141 25510 -38051
rect 25587 -38138 25659 -38046
rect 25736 -38138 37954 -38043
rect 25587 -38141 37954 -38138
rect 25428 -38146 37954 -38141
rect 15032 -38149 37954 -38146
rect 14883 -38152 37954 -38149
rect 14724 -38157 37954 -38152
rect -70936 -38163 37954 -38157
rect -55938 -38164 -55528 -38163
rect -45761 -38164 -45351 -38163
rect -35390 -38168 -34980 -38163
rect 14630 -38169 15040 -38163
use Buff_4x  Buff_4x_0
timestamp 1694601504
transform -1 0 -67571 0 1 37319
box -175 -237 958 1180
use Buff_4x  Buff_4x_1
timestamp 1694601504
transform 1 0 -69311 0 1 38859
box -175 -237 958 1180
use Buff_4x  Buff_4x_2
timestamp 1694601504
transform -1 0 -66792 0 1 42497
box -175 -237 958 1180
use Buff_4x  Buff_4x_3
timestamp 1694601504
transform 1 0 -69232 0 1 42509
box -175 -237 958 1180
use Buff_4x  Buff_4x_4
timestamp 1694601504
transform -1 0 -66849 0 1 40662
box -175 -237 958 1180
use Buff_4x  Buff_4x_5
timestamp 1694601504
transform 1 0 -69218 0 1 40669
box -175 -237 958 1180
use Buff_4x  Buff_4x_6
timestamp 1694601504
transform -1 0 -66844 0 1 38883
box -175 -237 958 1180
use Buff_4x  Buff_4x_7
timestamp 1694601504
transform 1 0 -57987 0 1 -36016
box -175 -237 958 1180
use Buff_4x  Buff_4x_8
timestamp 1694601504
transform 1 0 -49413 0 1 -37824
box -175 -237 958 1180
use Buff_4x  Buff_4x_9
timestamp 1694601504
transform 1 0 -27725 0 1 -37413
box -175 -237 958 1180
use Buff_4x  Buff_4x_10
timestamp 1694601504
transform 1 0 -12109 0 1 -37523
box -175 -237 958 1180
use Buff_4x  Buff_4x_11
timestamp 1694601504
transform 1 0 11940 0 1 -37706
box -175 -237 958 1180
use Buff_4x  Buff_4x_12
timestamp 1694601504
transform 1 0 708 0 1 -37587
box -175 -237 958 1180
use Buff_4x  Buff_4x_13
timestamp 1694601504
transform -1 0 21328 0 1 -37708
box -175 -237 958 1180
use Buff_16x  Buff_16x_0
timestamp 1694601232
transform -1 0 -66728 0 1 30655
box -160 -230 1608 1426
use Buff_16x  Buff_16x_1
timestamp 1694601232
transform 1 0 -68519 0 1 -26996
box -160 -230 1608 1426
use Buff_16x  Buff_16x_2
timestamp 1694601232
transform -1 0 -66735 0 1 22276
box -160 -230 1608 1426
use Buff_16x  Buff_16x_3
timestamp 1694601232
transform -1 0 -66751 0 1 13199
box -160 -230 1608 1426
use Buff_16x  Buff_16x_4
timestamp 1694601232
transform -1 0 -66752 0 1 631
box -160 -230 1608 1426
use Buff_16x  Buff_16x_5
timestamp 1694601232
transform -1 0 -66746 0 1 -8480
box -160 -230 1608 1426
use Buff_16x  Buff_16x_6
timestamp 1694601232
transform 1 0 -68426 0 1 -23943
box -160 -230 1608 1426
use Buff_16x  Buff_16x_7
timestamp 1694601232
transform 1 0 -56874 0 1 -36023
box -160 -230 1608 1426
use Buff_16x  Buff_16x_8
timestamp 1694601232
transform 1 0 -48300 0 1 -37831
box -160 -230 1608 1426
use Buff_16x  Buff_16x_9
timestamp 1694601232
transform 1 0 -26612 0 1 -37420
box -160 -230 1608 1426
use Buff_16x  Buff_16x_10
timestamp 1694601232
transform 1 0 -10996 0 1 -37530
box -160 -230 1608 1426
use Buff_16x  Buff_16x_11
timestamp 1694601232
transform 1 0 1821 0 1 -37594
box -160 -230 1608 1426
use Buff_16x  Buff_16x_12
timestamp 1694601232
transform -1 0 20215 0 1 -37715
box -160 -230 1608 1426
use Buff_16x  Buff_16x_13
timestamp 1694601232
transform 1 0 13053 0 1 -37713
box -160 -230 1608 1426
use CM_32_C  CM_32_C_0
timestamp 1693898149
transform 1 0 -32639 0 -1 -5340
box -789 -525 6929 5146
use CM_32_C  CM_32_C_1
timestamp 1693898149
transform 1 0 -32088 0 1 20988
box -789 -525 6929 5146
use CM_32_C  CM_32_C_2
timestamp 1693898149
transform 1 0 -4160 0 1 21215
box -789 -525 6929 5146
use CM_32_C  CM_32_C_3
timestamp 1693898149
transform 1 0 -3153 0 -1 -5132
box -789 -525 6929 5146
use CM_32_C  CM_32_C_4
timestamp 1693898149
transform 1 0 -31252 0 1 38293
box -789 -525 6929 5146
use CM_32_C  CM_32_C_5
timestamp 1693898149
transform 1 0 -52850 0 -1 -13710
box -789 -525 6929 5146
use CM_32_C  CM_32_C_6
timestamp 1693898149
transform 1 0 -3065 0 1 38218
box -789 -525 6929 5146
use CM_32_C  CM_32_C_7
timestamp 1693898149
transform 1 0 18219 0 1 21395
box -789 -525 6929 5146
use CM_32_C  CM_32_C_8
timestamp 1693898149
transform 1 0 18251 0 1 -9510
box -789 -525 6929 5146
use CM_32_C  CM_32_C_9
timestamp 1693898149
transform 1 0 -3109 0 1 -26408
box -789 -525 6929 5146
use CM_32_C  CM_32_C_10
timestamp 1693898149
transform 1 0 -31275 0 1 -26453
box -789 -525 6929 5146
use CM_32_C  CM_32_C_11
timestamp 1693898149
transform 1 0 -52897 0 1 -9549
box -789 -525 6929 5146
use CM_32_C  CM_32_C_12
timestamp 1693898149
transform 1 0 -52865 0 1 21357
box -789 -525 6929 5146
use CM_32_C  CM_32_C_13
timestamp 1693898149
transform 1 0 -31336 0 1 46498
box -789 -525 6929 5146
use CM_32_C  CM_32_C_14
timestamp 1693898149
transform 1 0 -31240 0 1 -34751
box -789 -525 6929 5146
use CM_32_C  CM_32_C_15
timestamp 1693898149
transform 1 0 7510 0 1 46458
box -789 -525 6929 5146
use CM_32_C  CM_32_C_16
timestamp 1693898149
transform 1 0 28915 0 1 21333
box -789 -525 6929 5146
use CM_32_C  CM_32_C_17
timestamp 1693898149
transform 1 0 28935 0 1 -9565
box -789 -525 6929 5146
use CM_32_C  CM_32_C_18
timestamp 1693898149
transform 1 0 7571 0 1 -34873
box -789 -525 6929 5146
use CM_32_C  CM_32_C_19
timestamp 1693898149
transform 1 0 -63250 0 1 21435
box -789 -525 6929 5146
use Current_Mirror_Top  Current_Mirror_Top_0
timestamp 1697714711
transform -1 0 -72254 0 -1 18354
box -186 -209 4486 6364
use INV_BUFF  INV_BUFF_0
timestamp 1694585882
transform 1 0 -33565 0 1 5082
box -90 0 858 813
use INV_BUFF  INV_BUFF_1
timestamp 1694585882
transform 1 0 -63023 0 1 5081
box -90 0 858 813
use INV_BUFF  INV_BUFF_2
timestamp 1694585882
transform 1 0 -33547 0 1 9621
box -90 0 858 813
use INV_BUFF  INV_BUFF_3
timestamp 1694585882
transform 1 0 -63015 0 1 6010
box -90 0 858 813
use INV_BUFF  INV_BUFF_4
timestamp 1694585882
transform 1 0 -63008 0 1 6924
box -90 0 858 813
use INV_BUFF  INV_BUFF_5
timestamp 1694585882
transform 1 0 -63008 0 1 7831
box -90 0 858 813
use INV_BUFF  INV_BUFF_6
timestamp 1694585882
transform 1 0 -63015 0 1 8745
box -90 0 858 813
use INV_BUFF  INV_BUFF_7
timestamp 1694585882
transform 1 0 -9864 0 1 46912
box -90 0 858 813
use INV_BUFF  INV_BUFF_8
timestamp 1694585882
transform 1 0 -63015 0 1 9659
box -90 0 858 813
use INV_BUFF  INV_BUFF_9
timestamp 1694585882
transform 1 0 -33557 0 1 5988
box -90 0 858 813
use INV_BUFF  INV_BUFF_10
timestamp 1694585882
transform 1 0 -33557 0 1 6902
box -90 0 858 813
use INV_BUFF  INV_BUFF_11
timestamp 1694585882
transform 1 0 -33549 0 1 7783
box -90 0 858 813
use INV_BUFF  INV_BUFF_12
timestamp 1694585882
transform 1 0 -33557 0 1 8721
box -90 0 858 813
use INV_BUFF  INV_BUFF_13
timestamp 1694585882
transform 1 0 -10468 0 1 25432
box -90 0 858 813
use INV_BUFF  INV_BUFF_14
timestamp 1694585882
transform 1 0 -59423 0 1 48813
box -90 0 858 813
use INV_BUFF  INV_BUFF_15
timestamp 1694585882
transform 1 0 -59404 0 1 45847
box -90 0 858 813
use INV_BUFF  INV_BUFF_16
timestamp 1694585882
transform 1 0 -59404 0 1 47320
box -90 0 858 813
use INV_BUFF  INV_BUFF_17
timestamp 1694585882
transform 1 0 -67689 0 1 -33292
box -90 0 858 813
use INV_BUFF  INV_BUFF_18
timestamp 1694585882
transform 1 0 -68533 0 1 45925
box -90 0 858 813
use INV_BUFF  INV_BUFF_19
timestamp 1694585882
transform 1 0 -68591 0 1 47370
box -90 0 858 813
use INV_BUFF  INV_BUFF_20
timestamp 1694585882
transform 1 0 -68590 0 1 48798
box -90 0 858 813
use INV_BUFF  INV_BUFF_21
timestamp 1694585882
transform 1 0 -67686 0 1 -31806
box -90 0 858 813
use INV_BUFF  INV_BUFF_22
timestamp 1694585882
transform 1 0 -69407 0 1 -31806
box -90 0 858 813
use INV_BUFF  INV_BUFF_23
timestamp 1694585882
transform 1 0 -67674 0 1 -34458
box -90 0 858 813
use INV_BUFF  INV_BUFF_24
timestamp 1694585882
transform 1 0 -69454 0 1 -34458
box -90 0 858 813
use INV_BUFF  INV_BUFF_25
timestamp 1694585882
transform 1 0 -69431 0 1 -33291
box -90 0 858 813
use LSBs_magic_TG  LSBs_magic_TG_0
timestamp 1694400330
transform 1 0 -15298 0 1 10723
box -6506 -12515 6485 6731
use MSB_Unit_Cell  MSB_Unit_Cell_0
timestamp 1695284343
transform 1 0 -29575 0 1 -3123
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_1
timestamp 1695284343
transform 1 0 -40058 0 1 -21095
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_2
timestamp 1695284343
transform 1 0 -813 0 1 -3021
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_3
timestamp 1695284343
transform 1 0 -39896 0 1 -12172
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_4
timestamp 1695284343
transform 1 0 -846 0 1 9661
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_5
timestamp 1695284343
transform 1 0 -14992 0 1 27080
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_6
timestamp 1695284343
transform 1 0 -1020 0 1 27144
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_7
timestamp 1695284343
transform 1 0 9954 0 1 27083
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_8
timestamp 1695284343
transform 1 0 9990 0 1 19084
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_9
timestamp 1695284343
transform 1 0 9804 0 1 9564
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_10
timestamp 1695284343
transform 1 0 10018 0 1 -2808
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_11
timestamp 1695284343
transform 1 0 9997 0 1 -12395
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_12
timestamp 1695284343
transform 1 0 10005 0 1 -20862
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_13
timestamp 1695284343
transform 1 0 -761 0 1 -20888
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_14
timestamp 1695284343
transform 1 0 -14949 0 1 -21038
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_15
timestamp 1695284343
transform 1 0 -28962 0 1 -20963
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_16
timestamp 1695284343
transform 1 0 -28814 0 1 27025
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_17
timestamp 1695284343
transform 1 0 -39878 0 1 27210
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_18
timestamp 1695284343
transform 1 0 -40078 0 1 18787
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_19
timestamp 1695284343
transform 1 0 -40053 0 1 9613
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_20
timestamp 1695284343
transform 1 0 -39873 0 1 -3205
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_21
timestamp 1695284343
transform 1 0 -14995 0 1 -29026
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_22
timestamp 1695284343
transform 1 0 -39907 0 1 -28997
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_23
timestamp 1695284343
transform 1 0 -14888 0 1 35592
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_24
timestamp 1695284343
transform 1 0 10114 0 1 35592
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_25
timestamp 1695284343
transform 1 0 -39935 0 1 35733
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_26
timestamp 1695284343
transform 1 0 -50241 0 1 35685
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_27
timestamp 1695284343
transform 1 0 -50252 0 1 27237
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_28
timestamp 1695284343
transform 1 0 -29683 0 1 9797
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_29
timestamp 1695284343
transform 1 0 -50260 0 1 9951
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_30
timestamp 1695284343
transform 1 0 -50283 0 1 -2977
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_31
timestamp 1695284343
transform 1 0 -50289 0 1 -28963
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_32
timestamp 1695284343
transform 1 0 20765 0 1 35508
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_33
timestamp 1695284343
transform 1 0 20849 0 1 -20927
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_34
timestamp 1695284343
transform 1 0 10129 0 1 -29051
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_35
timestamp 1695284343
transform 1 0 20837 0 1 -28978
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_36
timestamp 1695284343
transform 1 0 20861 0 1 -2931
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_37
timestamp 1695284343
transform 1 0 20849 0 1 27041
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_38
timestamp 1695284343
transform 1 0 20861 0 1 9596
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_39
timestamp 1695284343
transform 1 0 31566 0 1 -29013
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_40
timestamp 1695284343
transform 1 0 -50249 0 1 44017
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_41
timestamp 1695284343
transform 1 0 -39888 0 1 43904
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_42
timestamp 1695284343
transform 1 0 -16425 0 1 -12286
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_43
timestamp 1695284343
transform 1 0 -15065 0 1 43904
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_44
timestamp 1695284343
transform 1 0 -961 0 1 43960
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_45
timestamp 1695284343
transform 1 0 20759 0 1 43904
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_46
timestamp 1695284343
transform 1 0 31737 0 1 35609
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_47
timestamp 1695284343
transform 1 0 31756 0 1 27112
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_48
timestamp 1695284343
transform 1 0 31756 0 1 9590
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_49
timestamp 1695284343
transform 1 0 31529 0 1 -3154
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_50
timestamp 1695284343
transform 1 0 31546 0 1 -20902
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_51
timestamp 1695284343
transform 1 0 -60478 0 1 -29024
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_52
timestamp 1695284343
transform 1 0 -60428 0 1 27244
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_53
timestamp 1695284343
transform 1 0 -60409 0 1 9674
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_54
timestamp 1695284343
transform 1 0 -60427 0 1 -2638
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_55
timestamp 1695284343
transform 1 0 -60446 0 1 -12150
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_56
timestamp 1695284343
transform 1 0 -60446 0 1 -20926
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_57
timestamp 1695284343
transform 1 0 -39868 0 1 -37104
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_58
timestamp 1695284343
transform 1 0 -15702 0 1 18848
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_59
timestamp 1695284343
transform 1 0 -50256 0 1 -37104
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_60
timestamp 1695284343
transform 1 0 -15038 0 1 -37045
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_61
timestamp 1695284343
transform 1 0 -676 0 1 -37144
box -3642 1970 4332 7695
use MSB_Unit_Cell  MSB_Unit_Cell_62
timestamp 1695284343
transform 1 0 20886 0 1 -37123
box -3642 1970 4332 7695
use pmos_3p3_KG2TLM  pmos_3p3_KG2TLM_0
timestamp 1697714711
transform 1 0 -71407 0 1 12006
box -326 -190 326 190
use ppolyf_u_JWZPDU  ppolyf_u_JWZPDU_0
timestamp 1699423221
transform 1 0 -68761 0 1 59317
box -2844 -1287 2844 1287
use ppolyf_u_JWZPDU  ppolyf_u_JWZPDU_1
timestamp 1699423221
transform 1 0 -62944 0 1 59317
box -2844 -1287 2844 1287
use therm_Dec  therm_Dec_0
timestamp 1694585882
transform -1 0 -59160 0 1 42410
box -842 -4784 4258 891
use therm_Dec  therm_Dec_1
timestamp 1694585882
transform 1 0 -63356 0 1 -30910
box -842 -4784 4258 891
<< labels >>
flabel metal1 -62922 42795 -62922 42795 0 FreeSans 1600 180 0 0 R6
port 0 nsew
flabel metal1 -62697 42033 -62697 42033 0 FreeSans 1600 180 0 0 R5
port 1 nsew
flabel metal1 -62686 41842 -62686 41842 0 FreeSans 1600 180 0 0 R3
port 2 nsew
flabel metal1 -63016 39941 -63016 39941 0 FreeSans 1600 180 0 0 R2
port 4 nsew
flabel metal1 -61745 38976 -61745 38976 0 FreeSans 1600 180 0 0 R1
port 5 nsew
flabel metal1 -59622 -30510 -59622 -30510 0 FreeSans 1600 180 0 0 C6
port 7 nsew
flabel metal1 -59751 -31268 -59751 -31268 0 FreeSans 1600 180 0 0 C5
port 8 nsew
flabel metal1 -59767 -31480 -59767 -31480 0 FreeSans 1600 180 0 0 C3
port 9 nsew
flabel metal1 -59471 -32414 -59471 -32414 0 FreeSans 1600 180 0 0 C4
port 10 nsew
flabel metal1 -59496 -33364 -59495 -33363 0 FreeSans 1600 180 0 0 C2
port 11 nsew
flabel metal1 -60799 -34342 -60799 -34342 0 FreeSans 1600 180 0 0 C1
port 12 nsew
flabel metal1 -59069 -35292 -59069 -35292 0 FreeSans 1600 180 0 0 C0
port 13 nsew
flabel metal2 -66205 56961 -66205 56961 0 FreeSans 1600 0 0 0 VDD
port 14 nsew
flabel metal2 -65500 56961 -65500 56961 0 FreeSans 1600 0 0 0 VSS
port 15 nsew
flabel metal2 -70055 56960 -70055 56960 0 FreeSans 1600 0 0 0 OUT+
port 16 nsew
flabel metal2 -70725 56960 -70725 56960 0 FreeSans 1600 0 0 0 OUT-
port 17 nsew
flabel metal1 -71054 46329 -71054 46329 0 FreeSans 1600 0 0 0 B12
port 18 nsew
flabel metal1 -71158 47757 -71158 47757 0 FreeSans 1600 0 0 0 B11
port 19 nsew
flabel metal1 -71158 49217 -71158 49217 0 FreeSans 1600 0 0 0 B10
port 20 nsew
flabel metal1 -58264 46244 -58264 46244 0 FreeSans 1600 0 0 0 B12D
port 21 nsew
flabel metal1 -58248 47725 -58248 47725 0 FreeSans 1600 0 0 0 B11D
port 22 nsew
flabel metal1 -58312 49206 -58312 49206 0 FreeSans 1600 0 0 0 B10D
port 23 nsew
flabel metal1 -70997 -31385 -70997 -31385 0 FreeSans 1600 0 0 0 B9
port 24 nsew
flabel metal1 -70997 -32886 -70997 -32886 0 FreeSans 1600 0 0 0 B8
port 25 nsew
flabel metal1 -70995 -34041 -70995 -34041 0 FreeSans 1600 0 0 0 B7
port 26 nsew
flabel metal1 -64949 -31394 -64949 -31394 0 FreeSans 1600 0 0 0 B9D
port 27 nsew
flabel metal1 -64965 -32894 -64965 -32894 0 FreeSans 1600 0 0 0 B8D
port 28 nsew
flabel metal1 -64614 -33411 -64614 -33411 0 FreeSans 1600 0 0 0 B7D
port 29 nsew
flabel metal2 -8462 56671 -8462 56671 0 FreeSans 1600 0 0 0 SEL_L
port 30 nsew
flabel metal2 -9262 17224 -9262 17224 0 FreeSans 1600 0 0 0 SEL
port 31 nsew
flabel metal1 -71287 9158 -71287 9158 0 FreeSans 1600 0 0 0 B2
port 33 nsew
flabel metal1 -71238 8231 -71238 8231 0 FreeSans 1600 0 0 0 B3
port 34 nsew
flabel metal1 -71247 7330 -71247 7330 0 FreeSans 1600 0 0 0 B4
port 35 nsew
flabel metal1 -71260 6425 -71260 6425 0 FreeSans 1600 0 0 0 B5
port 36 nsew
flabel metal1 -71260 5476 -71260 5476 0 FreeSans 1600 0 0 0 B6
port 37 nsew
flabel metal1 -21771 6563 -21771 6563 0 FreeSans 1600 0 0 0 B2D
port 39 nsew
flabel metal1 -21838 5726 -21838 5726 0 FreeSans 1600 0 0 0 B3D
port 40 nsew
flabel metal1 -21869 4349 -21869 4349 0 FreeSans 1600 0 0 0 B5D
port 42 nsew
flabel metal1 -21749 4144 -21749 4144 0 FreeSans 1600 0 0 0 B6D
port 43 nsew
flabel metal3 -71716 11087 -71716 11087 0 FreeSans 1600 0 0 0 ITAIL
port 44 nsew
flabel metal1 -61942 49189 -61942 49189 0 FreeSans 1600 0 0 0 B10M
port 45 nsew
flabel metal1 -61889 47752 -61889 47752 0 FreeSans 1600 0 0 0 B11M
port 46 nsew
flabel metal1 -61880 46317 -61880 46317 0 FreeSans 1600 0 0 0 B12M
port 47 nsew
flabel metal1 -61926 10074 -61926 10074 0 FreeSans 1600 0 0 0 B1M
port 48 nsew
flabel metal1 -61926 9131 -61926 9131 0 FreeSans 1600 0 0 0 B2M
port 49 nsew
flabel metal1 -61840 8246 -61840 8246 0 FreeSans 1600 0 0 0 B3M
port 50 nsew
flabel metal1 -61859 6418 -61859 6418 0 FreeSans 1600 0 0 0 B5M
port 52 nsew
flabel metal1 -61859 5447 -61859 5447 0 FreeSans 1600 0 0 0 B6M
port 53 nsew
flabel metal1 -68193 -31413 -68193 -31413 0 FreeSans 1600 0 0 0 B9M
port 54 nsew
flabel metal1 -68241 -32892 -68241 -32892 0 FreeSans 1600 0 0 0 B8M
port 55 nsew
flabel metal1 -68246 -34064 -68246 -34064 0 FreeSans 1600 0 0 0 B7M
port 56 nsew
flabel metal2 -18625 -1475 -18625 -1475 0 FreeSans 1600 0 0 0 cur_1_d
port 57 nsew
flabel metal2 -18615 -1717 -18615 -1717 0 FreeSans 1600 0 0 0 cur_1_u
port 58 nsew
flabel metal2 -3712 -9514 -3712 -9514 0 FreeSans 1600 0 0 0 cur_2_u
port 59 nsew
flabel metal2 -3891 -10256 -3891 -10256 0 FreeSans 1600 0 0 0 cur_2_d
port 60 nsew
flabel metal2 -33153 -9733 -33153 -9733 0 FreeSans 1600 0 0 0 cur_3_u
port 61 nsew
flabel metal2 -33326 -10496 -33326 -10496 0 FreeSans 1600 0 0 0 cur_3_d
port 62 nsew
flabel via1 17434 -5121 17434 -5121 0 FreeSans 1600 0 0 0 cur_6_u
port 67 nsew
flabel via1 16728 -4415 16728 -4415 0 FreeSans 1600 0 0 0 cur_6_d
port 68 nsew
flabel via1 28346 -4449 28346 -4449 0 FreeSans 1600 0 0 0 cur_7_d
port 69 nsew
flabel via1 27847 -5178 27847 -5178 0 FreeSans 1600 0 0 0 cur_7_u
port 70 nsew
flabel metal2 6740 -29695 6740 -29695 0 FreeSans 1600 0 0 0 cur_8_d
port 71 nsew
flabel metal2 6444 -30543 6444 -30543 0 FreeSans 1600 0 0 0 cur_8_u
port 72 nsew
flabel via1 -3741 -22006 -3741 -22006 0 FreeSans 1600 0 0 0 cur_9_u
port 73 nsew
flabel via1 -3988 -21299 -3988 -21299 0 FreeSans 1600 0 0 0 cur_9_d
port 74 nsew
flabel metal2 -32268 -21425 -32268 -21425 0 FreeSans 1600 0 0 0 cur_10_d
port 75 nsew
flabel via1 -31914 -22050 -31914 -22050 0 FreeSans 1600 0 0 0 cur_10_u
port 76 nsew
flabel metal2 -32937 -30261 -32937 -30261 0 FreeSans 1600 0 0 0 cur_11_u
port 77 nsew
flabel metal2 -32633 -29584 -32633 -29584 0 FreeSans 1600 0 0 0 cur_11_d
port 78 nsew
flabel via1 -53963 -18822 -53963 -18822 0 FreeSans 1600 0 0 0 cur_12_d
port 79 nsew
flabel via1 -53385 -18108 -53385 -18108 0 FreeSans 1600 0 0 0 cur_12_u
port 80 nsew
flabel via1 -53526 -5156 -53526 -5156 0 FreeSans 1600 0 0 0 cur_13_u
port 81 nsew
flabel metal2 -53981 -4478 -53981 -4478 0 FreeSans 1600 0 0 0 cur_13_d
port 82 nsew
flabel metal2 -53480 25727 -53480 25727 0 FreeSans 1600 0 0 0 cur_14_u
port 83 nsew
flabel via1 -53847 26452 -53847 26452 0 FreeSans 1600 0 0 0 cur_14_d
port 84 nsew
flabel metal2 -64350 26491 -64350 26491 0 FreeSans 1600 0 0 0 cur_15_d
port 85 nsew
flabel via1 -64061 25827 -64061 25827 0 FreeSans 1600 0 0 0 cur_15_u
port 86 nsew
flabel metal2 -3887 43403 -3887 43403 0 FreeSans 1600 0 0 0 cur_18_d
port 91 nsew
flabel metal2 -4424 42632 -4424 42632 0 FreeSans 1600 0 0 0 cur_18_u
port 92 nsew
flabel via1 6457 50857 6457 50857 0 FreeSans 1600 0 0 0 cur_19_u
port 93 nsew
flabel via1 6716 51570 6716 51570 0 FreeSans 1600 0 0 0 cur_19_d
port 94 nsew
flabel metal2 17943 25792 17943 25792 0 FreeSans 1600 0 0 0 cur_20_u
port 95 nsew
flabel metal2 18577 26426 18577 26426 0 FreeSans 1600 0 0 0 cur_20_d
port 96 nsew
flabel via1 28291 26430 28291 26430 0 FreeSans 1600 0 0 0 cur_21_d
port 97 nsew
flabel metal2 28628 25710 28628 25710 0 FreeSans 1600 0 0 0 cur_21_u
port 98 nsew
flabel via1 -9289 38682 -9289 38682 0 FreeSans 1600 0 0 0 SEL_M
port 99 nsew
flabel via1 -33670 26100 -33670 26100 0 FreeSans 1600 0 0 0 cur_4_d
port 100 nsew
flabel metal1 -32670 25370 -32670 25370 0 FreeSans 1600 0 0 0 cur_4_u
port 101 nsew
flabel metal1 -4650 25590 -4650 25590 0 FreeSans 1600 0 0 0 cur_5_u
port 104 nsew
flabel via1 -5310 26320 -5310 26320 0 FreeSans 1600 0 0 0 cur_5_d
port 105 nsew
flabel metal1 -61670 7460 -61670 7460 0 FreeSans 1600 0 0 0 B4M
port 106 nsew
flabel via1 -67754 42934 -67754 42934 0 FreeSans 1600 0 0 0 R6m
port 107 nsew
flabel via1 -68313 42929 -68313 42929 0 FreeSans 1600 0 0 0 R5m
port 108 nsew
flabel via1 -67759 41087 -67759 41087 0 FreeSans 1600 0 0 0 R3m
port 109 nsew
flabel via1 -68323 41082 -68323 41082 0 FreeSans 1600 0 0 0 R4m
port 110 nsew
flabel via1 -67859 39291 -67859 39291 0 FreeSans 1600 0 0 0 R2m
port 111 nsew
flabel via1 -68403 39276 -68403 39276 0 FreeSans 1600 0 0 0 R1m
port 112 nsew
flabel via1 -68462 37729 -68462 37729 0 FreeSans 1600 0 0 0 R0m
port 113 nsew
flabel via2 -68271 31142 -68271 31142 0 FreeSans 1600 0 0 0 R6D
port 114 nsew
flabel via2 -68296 22772 -68296 22772 0 FreeSans 1600 0 0 0 R5D
port 115 nsew
flabel via2 -68296 13683 -68296 13683 0 FreeSans 1600 0 0 0 R4D
port 116 nsew
flabel via2 -68286 1107 -68286 1107 0 FreeSans 1600 0 0 0 R3D
port 117 nsew
flabel metal3 -68326 -8002 -68326 -8002 0 FreeSans 1600 0 0 0 R2D
port 118 nsew
flabel via2 -66806 -23468 -66806 -23468 0 FreeSans 1600 0 0 0 R1D
port 119 nsew
flabel via1 -66911 -26510 -66911 -26510 0 FreeSans 1600 0 0 0 R0D
port 120 nsew
flabel via1 -54378 -35576 -54378 -35576 0 FreeSans 1600 0 0 0 C0D
port 121 nsew
flabel metal2 -43846 -37370 -43846 -37370 0 FreeSans 1600 0 0 0 C1D
port 122 nsew
flabel metal2 -19358 -32063 -19358 -32063 0 FreeSans 1600 0 0 0 C2D
port 123 nsew
flabel metal2 -4539 -32103 -4539 -32103 0 FreeSans 1600 0 0 0 C3D
port 124 nsew
flabel metal2 5900 -37155 5900 -37155 0 FreeSans 1600 0 0 0 C4D
port 125 nsew
flabel metal2 16347 -37236 16347 -37236 0 FreeSans 1600 0 0 0 C6D
port 126 nsew
flabel metal2 16932 -37236 16932 -37236 0 FreeSans 1600 0 0 0 C5D
port 127 nsew
flabel metal1 20378 -37270 20378 -37270 0 FreeSans 1600 0 0 0 C5M
port 128 nsew
flabel metal1 12961 -37286 12961 -37286 0 FreeSans 1600 0 0 0 C6M
port 129 nsew
flabel metal1 1657 -37174 1657 -37174 0 FreeSans 1600 0 0 0 C4M
port 130 nsew
flabel metal1 -11174 -37146 -11174 -37146 0 FreeSans 1600 0 0 0 C3M
port 131 nsew
flabel metal1 -26775 -37147 -26775 -37147 0 FreeSans 1600 0 0 0 C2M
port 132 nsew
flabel metal1 -48442 -37356 -48442 -37356 0 FreeSans 1600 0 0 0 C1M
port 133 nsew
flabel metal1 -57065 -35603 -57065 -35603 0 FreeSans 1600 0 0 0 C0M
port 134 nsew
flabel metal1 -10820 16440 -10820 16440 0 FreeSans 1600 0 0 0 GT1
port 135 nsew
flabel metal1 -10815 14571 -10815 14571 0 FreeSans 1600 0 0 0 GT2
port 136 nsew
flabel metal1 -9121 16161 -9119 16165 0 FreeSans 1600 0 0 0 O-
port 137 nsew
flabel metal1 -9504 14319 -9504 14319 0 FreeSans 1600 0 0 0 O+
port 138 nsew
flabel metal1 -31821 43405 -31821 43405 0 FreeSans 1600 0 0 0 cur_16_d
port 87 nsew
flabel metal1 -31863 42688 -31863 42688 0 FreeSans 1600 0 0 0 cur_16_u
port 88 nsew
flabel via1 -32368 50912 -32368 50912 0 FreeSans 1600 0 0 0 cur_17_u
port 90 nsew
flabel via1 -32141 51608 -32141 51608 0 FreeSans 1600 0 0 0 cur_17_d
port 89 nsew
flabel metal1 -13396 12789 -13396 12789 0 FreeSans 1600 0 0 0 OUT6
port 139 nsew
flabel metal1 -13911 11641 -13911 11641 0 FreeSans 1600 0 0 0 OUT5
port 140 nsew
flabel metal1 -18100 9177 -18100 9177 0 FreeSans 1600 0 0 0 OUT4
port 141 nsew
flabel metal1 -15828 9182 -15828 9182 0 FreeSans 1600 0 0 0 OUT3
port 142 nsew
flabel metal3 -16568 9556 -16568 9556 0 FreeSans 1600 0 0 0 OUT2
port 143 nsew
flabel metal1 -17113 9757 -17113 9757 0 FreeSans 1600 0 0 0 OUT1
port 144 nsew
flabel metal2 -19472 12956 -19472 12956 0 FreeSans 1600 0 0 0 SD3_1
port 145 nsew
flabel metal1 -19341 11991 -19341 11991 0 FreeSans 1600 0 0 0 IT
port 146 nsew
flabel metal1 -17366 11810 -17366 11810 0 FreeSans 1600 0 0 0 SD0_2
port 147 nsew
flabel metal1 -14374 11345 -14374 11345 0 FreeSans 1600 0 0 0 SD0_1
port 148 nsew
flabel metal1 -18127 10606 -18127 10606 0 FreeSans 1600 0 0 0 G1_1
port 149 nsew
flabel metal1 -18040 10323 -18040 10323 0 FreeSans 1600 0 0 0 G1_2
port 150 nsew
flabel metal1 -18884 10428 -18884 10428 0 FreeSans 1600 0 0 0 SD1_1
port 151 nsew
flabel metal1 -19255 9535 -19255 9535 0 FreeSans 1600 0 0 0 SD2_1
port 152 nsew
flabel metal1 -18302 9532 -18302 9532 0 FreeSans 1600 0 0 0 SD2_5
port 153 nsew
flabel metal1 -17772 9520 -17772 9520 0 FreeSans 1600 0 0 0 SD2_4
port 154 nsew
flabel metal1 -17439 9580 -17439 9580 0 FreeSans 1600 0 0 0 SD2_3
port 155 nsew
flabel metal1 -16887 9403 -16887 9403 0 FreeSans 1600 0 0 0 G2_1
port 156 nsew
flabel metal1 -16899 9653 -16899 9653 0 FreeSans 1600 0 0 0 SD2_2
port 157 nsew
flabel metal3 -15823 7676 -15823 7676 0 FreeSans 1600 0 0 0 b1
port 158 nsew
flabel metal1 -15900 7456 -15900 7456 0 FreeSans 1600 0 0 0 b1b
port 159 nsew
flabel metal1 -15864 6804 -15864 6804 0 FreeSans 1600 0 0 0 b2
port 160 nsew
flabel metal1 -15891 6592 -15891 6592 0 FreeSans 1600 0 0 0 b2b
port 161 nsew
flabel metal3 -15828 5944 -15828 5944 0 FreeSans 1600 0 0 0 b3
port 162 nsew
flabel metal1 -15958 5733 -15958 5733 0 FreeSans 1600 0 0 0 b3b
port 163 nsew
flabel metal2 -15925 5083 -15925 5083 0 FreeSans 1600 0 0 0 b4
port 164 nsew
flabel metal1 -16035 4865 -16035 4865 0 FreeSans 1600 0 0 0 b4b
port 165 nsew
flabel metal1 -14409 6086 -14409 6086 0 FreeSans 1600 0 0 0 b5b
port 166 nsew
flabel metal2 -14381 5080 -14381 5080 0 FreeSans 1600 0 0 0 b5
port 167 nsew
flabel metal3 -12757 5084 -12757 5084 0 FreeSans 1600 0 0 0 b6
port 168 nsew
flabel metal1 -12919 4832 -12919 4832 0 FreeSans 1600 0 0 0 b6b
port 169 nsew
flabel metal2 -17015 3011 -17015 3011 0 FreeSans 1600 0 0 0 SDc1_1
port 170 nsew
flabel metal1 -18271 2108 -18271 2108 0 FreeSans 1600 0 0 0 Gc1_1
port 171 nsew
flabel metal1 -17285 1764 -17285 1764 0 FreeSans 1600 0 0 0 Gc1_2
port 172 nsew
flabel metal2 -17878 766 -17878 766 0 FreeSans 1600 0 0 0 SDc1_2
port 173 nsew
flabel metal2 -50839 50027 -50839 50027 0 FreeSans 1600 0 0 0 QB1
port 174 nsew
flabel via1 -50844 49004 -50844 49004 0 FreeSans 1600 0 0 0 Q1
port 175 nsew
flabel via1 -50788 46498 -50788 46498 0 FreeSans 1600 0 0 0 SDM_1
port 176 nsew
flabel metal1 -53012 46760 -53012 46760 0 FreeSans 1600 0 0 0 OUTM_1
port 177 nsew
flabel metal1 -42654 46649 -42654 46649 0 FreeSans 1600 0 0 0 OUTM_2
port 178 nsew
flabel via1 -40430 46382 -40430 46382 0 FreeSans 1600 0 0 0 SDM_2
port 179 nsew
flabel metal2 -40482 49696 -40482 49696 0 FreeSans 1600 0 0 0 QB2
port 180 nsew
flabel via1 -40471 48890 -40471 48890 0 FreeSans 1600 0 0 0 Q2
port 181 nsew
flabel metal2 -15653 49679 -15653 49679 0 FreeSans 1600 0 0 0 QB3
port 182 nsew
flabel via1 -15659 48891 -15659 48891 0 FreeSans 1600 0 0 0 Q3
port 183 nsew
flabel via1 -15609 46387 -15609 46387 0 FreeSans 1600 0 0 0 SDM_3
port 184 nsew
flabel metal1 -16195 46647 -16195 46647 0 FreeSans 1600 0 0 0 OUTM_3
port 185 nsew
flabel metal1 -1537 49974 -1537 49974 0 FreeSans 1600 0 0 0 QB4
port 186 nsew
flabel via1 -1558 48945 -1558 48945 0 FreeSans 1600 0 0 0 Q4
port 187 nsew
flabel via1 -1503 46452 -1503 46452 0 FreeSans 1600 0 0 0 SDM_4
port 188 nsew
flabel metal1 -2081 46712 -2081 46712 0 FreeSans 1600 0 0 0 OUTM_4
port 189 nsew
flabel metal1 19194 46651 19194 46651 0 FreeSans 1600 0 0 0 OUTM_5
port 190 nsew
flabel via1 20222 46389 20222 46389 0 FreeSans 1600 0 0 0 SDM_5
port 191 nsew
flabel via1 20169 48898 20169 48898 0 FreeSans 1600 0 0 0 Q5
port 192 nsew
flabel metal2 20204 49916 20204 49916 0 FreeSans 1600 0 0 0 QB5
port 193 nsew
flabel metal2 -50836 41318 -50836 41318 0 FreeSans 1600 0 0 0 QB6
port 194 nsew
flabel via1 -50842 40674 -50842 40674 0 FreeSans 1600 0 0 0 Q6
port 195 nsew
flabel via1 -50785 38172 -50785 38172 0 FreeSans 1600 0 0 0 SDM_6
port 196 nsew
flabel metal1 -51838 38425 -51838 38425 0 FreeSans 1600 0 0 0 OUTM_6
port 197 nsew
flabel metal1 -41498 38478 -41498 38478 0 FreeSans 1600 0 0 0 OUTM_7
port 198 nsew
flabel via1 -40476 38221 -40476 38221 0 FreeSans 1600 0 0 0 SDM_7
port 199 nsew
flabel via1 -40526 40716 -40526 40716 0 FreeSans 1600 0 0 0 Q7
port 200 nsew
flabel metal2 -40522 41755 -40522 41755 0 FreeSans 1600 0 0 0 QB7
port 201 nsew
flabel metal2 -15483 41601 -15483 41601 0 FreeSans 1600 0 0 0 QB8
port 202 nsew
flabel via1 -15483 40584 -15483 40584 0 FreeSans 1600 0 0 0 Q8
port 203 nsew
flabel via1 -15422 38081 -15422 38081 0 FreeSans 1600 0 0 0 SDM_8
port 204 nsew
flabel metal1 -16435 38337 -16435 38337 0 FreeSans 1600 0 0 0 OUTM_8
port 205 nsew
flabel metal1 8099 38339 8099 38339 0 FreeSans 1600 0 0 0 OUTM_9
port 206 nsew
flabel metal2 9569 38074 9569 38074 0 FreeSans 1600 0 0 0 SDM_9
port 207 nsew
flabel metal2 9524 40594 9524 40594 0 FreeSans 1600 0 0 0 Q9
port 208 nsew
flabel metal2 20167 41210 20167 41210 0 FreeSans 1600 0 0 0 QB10
port 210 nsew
flabel metal2 20171 40498 20171 40498 0 FreeSans 1600 0 0 0 Q10
port 211 nsew
flabel metal2 20209 37998 20209 37998 0 FreeSans 1600 0 0 0 SDM_10
port 212 nsew
flabel metal1 18843 38251 18843 38251 0 FreeSans 1600 0 0 0 OUTM_10
port 213 nsew
flabel metal1 30172 38353 30172 38353 0 FreeSans 1600 0 0 0 OUTM_11
port 214 nsew
flabel metal2 31193 38093 31193 38093 0 FreeSans 1600 0 0 0 SDM_11
port 215 nsew
flabel metal2 31151 40617 31151 40617 0 FreeSans 1600 0 0 0 Q11
port 216 nsew
flabel metal2 31138 41621 31138 41621 0 FreeSans 1600 0 0 0 QB11
port 217 nsew
flabel metal2 -61018 32872 -61018 32872 0 FreeSans 1600 0 0 0 QB12
port 218 nsew
flabel metal2 -61018 32226 -61018 32226 0 FreeSans 1600 0 0 0 Q12
port 219 nsew
flabel metal1 -61636 29988 -61636 29988 0 FreeSans 1600 0 0 0 OUTM_12
port 220 nsew
flabel metal2 -60973 29735 -60973 29735 0 FreeSans 1600 0 0 0 SDM_12
port 221 nsew
flabel metal2 -50791 29724 -50791 29724 0 FreeSans 1600 0 0 0 SDM_13
port 222 nsew
flabel metal1 -51530 29988 -51530 29988 0 FreeSans 1600 0 0 0 OUTM_13
port 223 nsew
flabel metal2 -50837 32233 -50837 32233 0 FreeSans 1600 0 0 0 Q13
port 224 nsew
flabel metal2 -50845 32929 -50845 32929 0 FreeSans 1600 0 0 0 QB13
port 225 nsew
flabel metal2 -40475 32810 -40475 32810 0 FreeSans 1600 0 0 0 QB14
port 226 nsew
flabel metal2 -40469 32192 -40469 32192 0 FreeSans 1600 0 0 0 Q14
port 227 nsew
flabel metal1 -41091 29960 -41091 29960 0 FreeSans 1600 0 0 0 OUTM_14
port 228 nsew
flabel metal2 -40421 29696 -40421 29696 0 FreeSans 1600 0 0 0 SDM_14
port 229 nsew
flabel metal2 -29358 29512 -29358 29512 0 FreeSans 1600 0 0 0 SDM_15
port 230 nsew
flabel metal1 -29973 29774 -29973 29774 0 FreeSans 1600 0 0 0 OUTM_15
port 231 nsew
flabel metal2 -29411 32006 -29411 32006 0 FreeSans 1600 0 0 0 Q15
port 232 nsew
flabel metal2 -29407 32614 -29407 32614 0 FreeSans 1600 0 0 0 QB15
port 233 nsew
flabel metal2 -15590 32619 -15590 32619 0 FreeSans 1600 0 0 0 QB16
port 234 nsew
flabel metal2 -15577 32056 -15577 32056 0 FreeSans 1600 0 0 0 Q16
port 235 nsew
flabel metal1 -14556 29833 -14556 29833 0 FreeSans 1600 0 0 0 OUTM_16
port 236 nsew
flabel metal2 -15537 29568 -15537 29568 0 FreeSans 1600 0 0 0 SDM_16
port 237 nsew
flabel metal2 -1567 29628 -1567 29628 0 FreeSans 1600 0 0 0 SDM_17
port 238 nsew
flabel metal1 -2165 29900 -2165 29900 0 FreeSans 1600 0 0 0 OUTM_17
port 239 nsew
flabel metal2 -1608 32119 -1608 32119 0 FreeSans 1600 0 0 0 Q17
port 240 nsew
flabel metal2 -1617 32509 -1617 32509 0 FreeSans 1600 0 0 0 QB17
port 241 nsew
flabel metal2 9370 32624 9370 32624 0 FreeSans 1600 0 0 0 QB18
port 242 nsew
flabel metal2 9366 32067 9366 32067 0 FreeSans 1600 0 0 0 Q18
port 243 nsew
flabel metal1 8705 29832 8705 29832 0 FreeSans 1600 0 0 0 OUTM_18
port 244 nsew
flabel metal2 9418 29576 9418 29576 0 FreeSans 1600 0 0 0 SDM_18
port 245 nsew
flabel metal2 20311 29529 20311 29529 0 FreeSans 1600 0 0 0 SDM_19
port 246 nsew
flabel metal1 19686 29794 19686 29794 0 FreeSans 1600 0 0 0 OUTM_19
port 247 nsew
flabel metal2 20252 32480 20252 32480 0 FreeSans 1600 0 0 0 QB19
port 248 nsew
flabel metal2 20252 32020 20252 32020 0 FreeSans 1600 0 0 0 Q19
port 249 nsew
flabel metal2 31159 32534 31159 32534 0 FreeSans 1600 0 0 0 QB20
port 250 nsew
flabel metal2 31166 32077 31166 32077 0 FreeSans 1600 0 0 0 Q20
port 251 nsew
flabel metal2 31214 29606 31214 29606 0 FreeSans 1600 0 0 0 SDM_20
port 252 nsew
flabel metal1 30693 29867 30693 29867 0 FreeSans 1600 0 0 0 OUTM_20
port 253 nsew
flabel metal1 -41219 21542 -41219 21542 0 FreeSans 1600 0 0 0 OUTM_21
port 254 nsew
flabel metal2 -40619 21271 -40619 21271 0 FreeSans 1600 0 0 0 SDM_21
port 255 nsew
flabel metal2 -40670 24142 -40670 24142 0 FreeSans 1600 0 0 0 QB21
port 256 nsew
flabel metal2 -40666 23756 -40666 23756 0 FreeSans 1600 0 0 0 Q21
port 257 nsew
flabel metal2 -16295 23835 -16295 23835 0 FreeSans 1600 0 0 0 Q22
port 258 nsew
flabel metal2 -16286 24146 -16286 24146 0 FreeSans 1600 0 0 0 QB22
port 259 nsew
flabel metal2 -16243 21324 -16243 21324 0 FreeSans 1600 0 0 0 SDM_22
port 260 nsew
flabel metal1 -16436 21594 -16436 21594 0 FreeSans 1600 0 0 0 OUTM_22
port 261 nsew
flabel metal1 9249 21828 9249 21828 0 FreeSans 1600 0 0 0 OUTM_23
port 262 nsew
flabel metal2 9443 21568 9443 21568 0 FreeSans 1600 0 0 0 SDM_23
port 263 nsew
flabel metal2 9398 24499 9398 24499 0 FreeSans 1600 0 0 0 QB23
port 264 nsew
flabel metal2 9398 24063 9398 24063 0 FreeSans 1600 0 0 0 Q23
port 265 nsew
flabel metal2 -61005 14640 -61005 14640 0 FreeSans 1600 0 0 0 Q24
port 266 nsew
flabel metal2 -61010 15069 -61010 15069 0 FreeSans 1600 0 0 0 QB24
port 267 nsew
flabel metal2 -60957 12145 -60957 12145 0 FreeSans 1600 0 0 0 SDM_24
port 268 nsew
flabel metal1 -61475 12424 -61475 12424 0 FreeSans 1600 0 0 0 OUTM_24
port 269 nsew
flabel metal1 -51413 12703 -51413 12703 0 FreeSans 1600 0 0 0 OUTM_25
port 270 nsew
flabel metal2 -50795 12429 -50795 12429 0 FreeSans 1600 0 0 0 SDM_25
port 271 nsew
flabel metal2 -50856 15325 -50856 15325 0 FreeSans 1600 0 0 0 QB25
port 272 nsew
flabel metal2 -50853 14943 -50853 14943 0 FreeSans 1600 0 0 0 Q25
port 273 nsew
flabel metal2 -40642 14598 -40642 14598 0 FreeSans 1600 0 0 0 Q26
port 274 nsew
flabel metal2 -40640 14940 -40640 14940 0 FreeSans 1600 0 0 0 QB26
port 275 nsew
flabel metal1 -41203 12361 -41203 12361 0 FreeSans 1600 0 0 0 OUTM_26
port 276 nsew
flabel metal2 -40590 12100 -40590 12100 0 FreeSans 1600 0 0 0 SDM_26
port 277 nsew
flabel metal2 -30225 12279 -30225 12279 0 FreeSans 1600 0 0 0 SDM_27
port 279 nsew
flabel metal1 -30858 12548 -30858 12548 0 FreeSans 1600 0 0 0 OUTM_27
port 280 nsew
flabel metal2 -30273 14779 -30273 14779 0 FreeSans 1600 0 0 0 Q27
port 281 nsew
flabel metal2 -30283 15196 -30283 15196 0 FreeSans 1600 0 0 0 QB27
port 282 nsew
flabel metal2 -1444 15033 -1444 15033 0 FreeSans 1600 0 0 0 QB28
port 283 nsew
flabel metal2 -1436 14645 -1436 14645 0 FreeSans 1600 0 0 0 Q28
port 284 nsew
flabel metal2 -1385 12143 -1385 12143 0 FreeSans 1600 0 0 0 SDM_28
port 285 nsew
flabel metal1 -1995 12420 -1995 12420 0 FreeSans 1600 0 0 0 OUTM_28
port 286 nsew
flabel metal1 8734 12316 8734 12316 0 FreeSans 1600 0 0 0 OUTM_29
port 287 nsew
flabel metal2 9262 12052 9262 12052 0 FreeSans 1600 0 0 0 SDM_29
port 288 nsew
flabel metal2 9216 14920 9216 14920 0 FreeSans 1600 0 0 0 QB29
port 289 nsew
flabel metal2 9210 14495 9210 14495 0 FreeSans 1600 0 0 0 Q29
port 290 nsew
flabel metal2 20265 14595 20265 14595 0 FreeSans 1600 0 0 0 Q30
port 291 nsew
flabel metal2 20277 14973 20277 14973 0 FreeSans 1600 0 0 0 QB30
port 292 nsew
flabel metal2 20323 12083 20323 12083 0 FreeSans 1600 0 0 0 SDM_30
port 293 nsew
flabel metal1 19701 12344 19701 12344 0 FreeSans 1600 0 0 0 OUTM_30
port 294 nsew
flabel metal1 30613 12343 30613 12343 0 FreeSans 1600 0 0 0 OUTM_31
port 295 nsew
flabel metal2 31218 12069 31218 12069 0 FreeSans 1600 0 0 0 SDM_31
port 296 nsew
flabel metal2 31165 14566 31165 14566 0 FreeSans 1600 0 0 0 Q31
port 297 nsew
flabel metal2 31160 14967 31160 14967 0 FreeSans 1600 0 0 0 QB31
port 298 nsew
flabel metal2 -61030 2737 -61030 2737 0 FreeSans 1600 0 0 0 QB32
port 299 nsew
flabel metal2 -61020 2298 -61020 2298 0 FreeSans 1600 0 0 0 Q32
port 300 nsew
flabel metal2 -60965 -145 -60965 -145 0 FreeSans 1600 0 0 0 SDM_32
port 301 nsew
flabel metal1 -61422 112 -61422 112 0 FreeSans 1600 0 0 0 OUTM_32
port 302 nsew
flabel metal1 -51436 -225 -51436 -225 0 FreeSans 1600 0 0 0 OUTM_33
port 303 nsew
flabel metal2 -50831 -496 -50831 -496 0 FreeSans 1600 0 0 0 SDM_33
port 304 nsew
flabel metal2 -50879 2001 -50879 2001 0 FreeSans 1600 0 0 0 Q33
port 305 nsew
flabel metal2 -50871 2373 -50871 2373 0 FreeSans 1600 0 0 0 QB33
port 306 nsew
flabel metal2 -40464 2145 -40464 2145 0 FreeSans 1600 0 0 0 QB34
port 307 nsew
flabel metal2 -40466 1633 -40466 1633 0 FreeSans 1600 0 0 0 Q34
port 308 nsew
flabel metal2 -40421 -721 -40421 -721 0 FreeSans 1600 0 0 0 SDM_34
port 309 nsew
flabel metal1 -41024 -453 -41024 -453 0 FreeSans 1600 0 0 0 OUTM_34
port 310 nsew
flabel metal1 -30696 -374 -30696 -374 0 FreeSans 1600 0 0 0 OUTM_35
port 311 nsew
flabel metal2 -30123 -636 -30123 -636 0 FreeSans 1600 0 0 0 SDM_35
port 312 nsew
flabel metal2 -30173 1853 -30173 1853 0 FreeSans 1600 0 0 0 Q35
port 313 nsew
flabel metal2 -30160 2230 -30160 2230 0 FreeSans 1600 0 0 0 QB35
port 314 nsew
flabel metal2 -1409 2359 -1409 2359 0 FreeSans 1600 0 0 0 QB36
port 315 nsew
flabel metal2 -1401 1886 -1401 1886 0 FreeSans 1600 0 0 0 Q36
port 316 nsew
flabel metal2 -1353 -558 -1353 -558 0 FreeSans 1600 0 0 0 SDM_36
port 317 nsew
flabel metal1 -1962 -270 -1962 -270 0 FreeSans 1600 0 0 0 OUTM_36
port 318 nsew
flabel metal1 8872 -59 8872 -59 0 FreeSans 1600 0 0 0 OUTM_37
port 319 nsew
flabel metal2 9473 -324 9473 -324 0 FreeSans 1600 0 0 0 SDM_37
port 320 nsew
flabel metal2 9417 2538 9417 2538 0 FreeSans 1600 0 0 0 QB37
port 321 nsew
flabel metal2 9433 2092 9433 2092 0 FreeSans 1600 0 0 0 Q37
port 322 nsew
flabel metal2 20264 1967 20264 1967 0 FreeSans 1600 0 0 0 Q38
port 323 nsew
flabel metal2 20272 2436 20272 2436 0 FreeSans 1600 0 0 0 QB38
port 324 nsew
flabel metal2 20322 -441 20322 -441 0 FreeSans 1600 0 0 0 SDM_38
port 325 nsew
flabel metal1 19706 -182 19706 -182 0 FreeSans 1600 0 0 0 OUTM_38
port 326 nsew
flabel metal1 30393 -406 30393 -406 0 FreeSans 1600 0 0 0 OUTM_39
port 327 nsew
flabel metal2 30983 -671 30983 -671 0 FreeSans 1600 0 0 0 SDM_39
port 328 nsew
flabel metal2 30932 2196 30932 2196 0 FreeSans 1600 0 0 0 QB39
port 329 nsew
flabel metal2 30940 1777 30940 1777 0 FreeSans 1600 0 0 0 Q39
port 330 nsew
flabel metal2 -61046 -7221 -61043 -7221 0 FreeSans 1600 0 0 0 Q40
port 331 nsew
flabel metal2 -61035 -6786 -61032 -6786 0 FreeSans 1600 0 0 0 QB40
port 332 nsew
flabel metal2 -60984 -9670 -60984 -9670 0 FreeSans 1600 0 0 0 SDM_40
port 333 nsew
flabel metal1 -61591 -9397 -61591 -9397 0 FreeSans 1600 0 0 0 OUTM_40
port 334 nsew
flabel metal1 -41042 -9419 -41042 -9419 0 FreeSans 1600 0 0 0 OUTM_41
port 335 nsew
flabel metal2 -40440 -9681 -40440 -9681 0 FreeSans 1600 0 0 0 SDM_41
port 336 nsew
flabel metal2 -40492 -6848 -40492 -6848 0 FreeSans 1600 0 0 0 QB41
port 337 nsew
flabel metal2 -40484 -7218 -40484 -7218 0 FreeSans 1600 0 0 0 Q41
port 338 nsew
flabel metal2 -17018 -7285 -17018 -7285 0 FreeSans 1600 0 0 0 Q42
port 339 nsew
flabel metal2 -17018 -6934 -17018 -6934 0 FreeSans 1600 0 0 0 QB42
port 340 nsew
flabel metal2 -16964 -9790 -16964 -9790 0 FreeSans 1600 0 0 0 SDM_42
port 341 nsew
flabel metal1 -17591 -9536 -17591 -9536 0 FreeSans 1600 0 0 0 OUTM_42
port 342 nsew
flabel metal1 8856 -9647 8856 -9647 0 FreeSans 1600 0 0 0 OUTM_43
port 343 nsew
flabel metal2 9448 -9908 9448 -9908 0 FreeSans 1600 0 0 0 SDM_43
port 344 nsew
flabel metal2 9399 -7406 9399 -7406 0 FreeSans 1600 0 0 0 Q43
port 345 nsew
flabel metal2 9399 -7041 9399 -7041 0 FreeSans 1600 0 0 0 QB43
port 346 nsew
flabel metal2 -61051 -15610 -61051 -15610 0 FreeSans 1600 0 0 0 QB44
port 347 nsew
flabel metal2 -61042 -16000 -61042 -16000 0 FreeSans 1600 0 0 0 Q44
port 348 nsew
flabel metal1 -61594 -18177 -61594 -18177 0 FreeSans 1600 0 0 0 OUTM_44
port 349 nsew
flabel metal2 -60992 -18444 -60992 -18444 0 FreeSans 1600 0 0 0 SDM_44
port 350 nsew
flabel metal2 -40607 -18603 -40607 -18603 0 FreeSans 1600 0 0 0 SDM_45
port 351 nsew
flabel metal1 -41211 -18344 -41211 -18344 0 FreeSans 1600 0 0 0 OUTM_45
port 352 nsew
flabel metal2 -40649 -16156 -40649 -16156 0 FreeSans 1600 0 0 0 Q45
port 353 nsew
flabel metal2 -40655 -15727 -40655 -15727 0 FreeSans 1600 0 0 0 QB45
port 354 nsew
flabel metal2 -29562 -15641 -29562 -15641 0 FreeSans 1600 0 0 0 QB46
port 355 nsew
flabel metal2 -29553 -16035 -29553 -16035 0 FreeSans 1600 0 0 0 Q46
port 356 nsew
flabel metal2 -29505 -18460 -29505 -18460 0 FreeSans 1600 0 0 0 SDM_46
port 357 nsew
flabel metal1 -30120 -18212 -30120 -18212 0 FreeSans 1600 0 0 0 OUTM_46
port 358 nsew
flabel metal1 -16109 -18286 -16109 -18286 0 FreeSans 1600 0 0 0 OUTM_47
port 359 nsew
flabel metal2 -15496 -18552 -15496 -18552 0 FreeSans 1600 0 0 0 SDM_47
port 360 nsew
flabel metal2 -15542 -16145 -15542 -16145 0 FreeSans 1600 0 0 0 Q47
port 361 nsew
flabel metal2 -15548 -15706 -15548 -15706 0 FreeSans 1600 0 0 0 QB47
port 362 nsew
flabel metal2 -1367 -15513 -1367 -15513 0 FreeSans 1600 0 0 0 QB48
port 363 nsew
flabel metal2 -1352 -15971 -1352 -15971 0 FreeSans 1600 0 0 0 Q48
port 364 nsew
flabel metal2 -1302 -18395 -1302 -18395 0 FreeSans 1600 0 0 0 SDM_48
port 365 nsew
flabel metal1 -1909 -18140 -1909 -18140 0 FreeSans 1600 0 0 0 OUTM_48
port 366 nsew
flabel metal1 8849 -18110 8849 -18110 0 FreeSans 1600 0 0 0 OUTM_49
port 367 nsew
flabel metal2 9458 -18364 9458 -18364 0 FreeSans 1600 0 0 0 SDM_49
port 368 nsew
flabel metal2 9413 -15936 9413 -15936 0 FreeSans 1600 0 0 0 Q49
port 369 nsew
flabel metal2 9416 -15469 9416 -15469 0 FreeSans 1600 0 0 0 QB49
port 370 nsew
flabel metal2 20253 -15585 20253 -15585 0 FreeSans 1600 0 0 0 QB50
port 371 nsew
flabel metal2 20256 -15955 20256 -15955 0 FreeSans 1600 0 0 0 Q50
port 372 nsew
flabel metal2 20305 -18438 20305 -18438 0 FreeSans 1600 0 0 0 SDM_50
port 373 nsew
flabel metal1 19704 -18176 19704 -18176 0 FreeSans 1600 0 0 0 OUTM_50
port 374 nsew
flabel metal1 30390 -18153 30390 -18153 0 FreeSans 1600 0 0 0 OUTM_51
port 375 nsew
flabel metal2 31000 -18397 31000 -18397 0 FreeSans 1600 0 0 0 SDM_51
port 376 nsew
flabel metal2 30949 -16022 30949 -16022 0 FreeSans 1600 0 0 0 Q51
port 377 nsew
flabel metal2 30957 -15529 30957 -15529 0 FreeSans 1600 0 0 0 QB51
port 378 nsew
flabel metal2 -61078 -23697 -61078 -23697 0 FreeSans 1600 0 0 0 QB52
port 379 nsew
flabel metal2 -61058 -24102 -61058 -24102 0 FreeSans 1600 0 0 0 Q52
port 380 nsew
flabel metal2 -61022 -26529 -61022 -26529 0 FreeSans 1600 0 0 0 SDM_52
port 381 nsew
flabel metal1 -61625 -26273 -61625 -26273 0 FreeSans 1600 0 0 0 OUTM_52
port 382 nsew
flabel metal1 -51427 -26213 -51427 -26213 0 FreeSans 1600 0 0 0 OUTM_53
port 383 nsew
flabel metal2 -50832 -26455 -50832 -26455 0 FreeSans 1600 0 0 0 SDM_53
port 384 nsew
flabel metal2 -50890 -24067 -50890 -24067 0 FreeSans 1600 0 0 0 Q53
port 385 nsew
flabel metal2 -50885 -23656 -50885 -23656 0 FreeSans 1600 0 0 0 QB53
port 386 nsew
flabel metal2 -40501 -23608 -40501 -23608 0 FreeSans 1600 0 0 0 QB54
port 387 nsew
flabel metal2 -40504 -24077 -40504 -24077 0 FreeSans 1600 0 0 0 Q54
port 388 nsew
flabel metal2 -40449 -26494 -40449 -26494 0 FreeSans 1600 0 0 0 SDM_54
port 389 nsew
flabel metal1 -41065 -26246 -41065 -26246 0 FreeSans 1600 0 0 0 OUTM_54
port 390 nsew
flabel metal1 -16159 -26281 -16159 -26281 0 FreeSans 1600 0 0 0 OUTM_55
port 391 nsew
flabel metal2 -15536 -26528 -15536 -26528 0 FreeSans 1600 0 0 0 SDM_55
port 392 nsew
flabel metal2 -15597 -23669 -15597 -23669 0 FreeSans 1600 0 0 0 QB55
port 393 nsew
flabel metal2 -15583 -24107 -15583 -24107 0 FreeSans 1600 0 0 0 Q55
port 394 nsew
flabel metal2 9527 -24138 9527 -24138 0 FreeSans 1600 0 0 0 Q56
port 395 nsew
flabel metal2 9527 -23640 9527 -23640 0 FreeSans 1600 0 0 0 QB56
port 396 nsew
flabel metal2 9586 -26564 9586 -26564 0 FreeSans 1600 0 0 0 SDM_56
port 397 nsew
flabel metal1 8981 -26302 8981 -26302 0 FreeSans 1600 0 0 0 OUTM_56
port 398 nsew
flabel metal1 19679 -26233 19679 -26233 0 FreeSans 1600 0 0 0 OUTM_57
port 399 nsew
flabel metal2 20288 -26481 20290 -26481 0 FreeSans 1600 0 0 0 SDM_57
port 400 nsew
flabel metal2 20239 -24082 20239 -24082 0 FreeSans 1600 0 0 0 Q57
port 401 nsew
flabel metal2 20239 -23616 20239 -23616 0 FreeSans 1600 0 0 0 QB57
port 402 nsew
flabel metal2 30970 -23643 30970 -23643 0 FreeSans 1600 0 0 0 QB58
port 403 nsew
flabel metal2 30978 -24069 30978 -24069 0 FreeSans 1600 0 0 0 Q58
port 404 nsew
flabel metal2 31027 -26509 31027 -26509 0 FreeSans 1600 0 0 0 SDM_58
port 405 nsew
flabel metal1 30417 -26269 30417 -26269 0 FreeSans 1600 0 0 0 OUTM_58
port 406 nsew
flabel metal1 -51425 -34357 -51425 -34357 0 FreeSans 1600 0 0 0 OUTM_59
port 407 nsew
flabel metal2 -50796 -34600 -50796 -34600 0 FreeSans 1600 0 0 0 SDM_59
port 408 nsew
flabel metal2 -50849 -32190 -50849 -32190 0 FreeSans 1600 0 0 0 Q59
port 409 nsew
flabel metal2 -50849 -31667 -50849 -31667 0 FreeSans 1600 0 0 0 QB59
port 410 nsew
flabel metal2 -40471 -31620 -40471 -31620 0 FreeSans 1600 0 0 0 QB60
port 411 nsew
flabel metal2 -40454 -32193 -40454 -32193 0 FreeSans 1600 0 0 0 Q60
port 412 nsew
flabel metal2 -40400 -34611 -40400 -34611 0 FreeSans 1600 0 0 0 SDM_60
port 413 nsew
flabel metal1 -41013 -34355 -41013 -34355 0 FreeSans 1600 0 0 0 OUTM_60
port 414 nsew
flabel metal1 -16192 -34296 -16192 -34296 0 FreeSans 1600 0 0 0 OUTM_61
port 415 nsew
flabel metal2 -15583 -34540 -15583 -34540 0 FreeSans 1600 0 0 0 SDM_61
port 416 nsew
flabel metal2 -15637 -32076 -15637 -32076 0 FreeSans 1600 0 0 0 Q61
port 417 nsew
flabel metal2 -15628 -31648 -15628 -31648 0 FreeSans 1600 0 0 0 QB61
port 418 nsew
flabel metal2 -1280 -31747 -1280 -31747 0 FreeSans 1600 0 0 0 QB62
port 419 nsew
flabel metal2 -1269 -32280 -1269 -32280 0 FreeSans 1600 0 0 0 Q62
port 420 nsew
flabel metal1 -1819 -34398 -1819 -34398 0 FreeSans 1600 0 0 0 OUTM_62
port 421 nsew
flabel metal2 -1221 -34628 -1221 -34628 0 FreeSans 1600 0 0 0 SDM_62
port 422 nsew
flabel metal2 20342 -34616 20342 -34616 0 FreeSans 1600 0 0 0 SDM_63
port 423 nsew
flabel metal1 19737 -34377 19737 -34377 0 FreeSans 1600 0 0 0 OUTM_63
port 424 nsew
flabel metal2 20284 -32259 20284 -32259 0 FreeSans 1600 0 0 0 Q63
port 425 nsew
flabel metal2 20282 -31711 20282 -31711 0 FreeSans 1600 0 0 0 QB63
port 426 nsew
flabel metal2 -30266 46983 -30266 46983 0 FreeSans 1600 0 0 0 C1_0
port 427 nsew
flabel metal1 -30719 47750 -30719 47750 0 FreeSans 1600 0 0 0 C1_1
port 428 nsew
flabel metal2 -31323 47896 -31323 47896 0 FreeSans 1600 0 0 0 C1_2
port 429 nsew
flabel metal2 -30715 49131 -30714 49131 0 FreeSans 1600 0 0 0 C1_3
port 430 nsew
flabel metal2 8581 46944 8581 46944 0 FreeSans 1600 0 0 0 C2_0
port 431 nsew
flabel metal1 8124 47715 8124 47715 0 FreeSans 1600 0 0 0 C2_1
port 432 nsew
flabel metal2 7513 47904 7513 47904 0 FreeSans 1600 0 0 0 C2_2
port 433 nsew
flabel metal2 8131 49091 8131 49091 0 FreeSans 1600 0 0 0 C2_3
port 434 nsew
flabel metal2 -30178 38770 -30178 38770 0 FreeSans 1600 0 0 0 C3_0
port 435 nsew
flabel metal1 -30641 39556 -30641 39556 0 FreeSans 1600 0 0 0 C3_1
port 436 nsew
flabel metal2 -31256 39766 -31256 39766 0 FreeSans 1600 0 0 0 C3_2
port 437 nsew
flabel metal2 -30630 40925 -30630 40925 0 FreeSans 1600 0 0 0 C3_3
port 438 nsew
flabel metal2 -1993 38700 -1993 38700 0 FreeSans 1600 0 0 0 C4_0
port 439 nsew
flabel metal1 -2437 39500 -2437 39500 0 FreeSans 1600 0 0 0 C4_1
port 440 nsew
flabel metal2 -3066 39694 -3066 39694 0 FreeSans 1600 0 0 0 C4_2
port 441 nsew
flabel metal2 -2443 40853 -2443 40853 0 FreeSans 1600 0 0 0 C4_3
port 442 nsew
flabel metal2 -62178 21920 -62178 21920 0 FreeSans 1600 0 0 0 C5_0
port 443 nsew
flabel metal1 -62630 22915 -62630 22915 0 FreeSans 1600 0 0 0 C5_1
port 444 nsew
flabel metal2 -63242 22948 -63242 22948 0 FreeSans 1600 0 0 0 C5_2
port 445 nsew
flabel metal2 -62633 24076 -62633 24076 0 FreeSans 1600 0 0 0 C5_3
port 446 nsew
flabel metal2 -51790 21843 -51790 21843 0 FreeSans 1600 0 0 0 C6_0
port 447 nsew
flabel metal1 -52246 22619 -52246 22619 0 FreeSans 1600 0 0 0 C6_1
port 448 nsew
flabel metal2 -52857 22932 -52857 22932 0 FreeSans 1600 0 0 0 C6_2
port 449 nsew
flabel metal2 -52248 23999 -52248 23999 0 FreeSans 1600 0 0 0 C6_3
port 450 nsew
flabel metal2 -31020 21469 -31020 21469 0 FreeSans 1600 0 0 0 C7_0
port 451 nsew
flabel metal1 -31475 22256 -31475 22256 0 FreeSans 1600 0 0 0 C7_1
port 452 nsew
flabel metal2 -32087 22472 -32087 22472 0 FreeSans 1600 0 0 0 C7_2
port 453 nsew
flabel metal2 -31469 23625 -31469 23625 0 FreeSans 1600 0 0 0 C7_3
port 454 nsew
flabel metal2 -3096 21704 -3094 21704 0 FreeSans 1600 0 0 0 C8_0
port 455 nsew
flabel metal1 -3540 22485 -3540 22485 0 FreeSans 1600 0 0 0 C8_1
port 456 nsew
flabel metal2 -4145 22610 -4145 22610 0 FreeSans 1600 0 0 0 C8_2
port 457 nsew
flabel metal2 -3537 23849 -3537 23849 0 FreeSans 1600 0 0 0 C8_3
port 458 nsew
flabel metal2 19287 21883 19287 21883 0 FreeSans 1600 0 0 0 C9_0
port 459 nsew
flabel metal1 18839 22672 18839 22672 0 FreeSans 1600 0 0 0 C9_1
port 460 nsew
flabel metal2 18227 22862 18227 22862 0 FreeSans 1600 0 0 0 C9_2
port 461 nsew
flabel metal2 18840 24025 18840 24025 0 FreeSans 1600 0 0 0 C9_3
port 462 nsew
flabel metal2 29980 21775 29980 21775 0 FreeSans 1600 0 0 0 C10_0
port 463 nsew
flabel metal1 29538 22600 29538 22600 0 FreeSans 1600 0 0 0 C10_1
port 464 nsew
flabel metal2 28935 22794 28935 22794 0 FreeSans 1600 0 0 0 C10_2
port 465 nsew
flabel metal2 29530 23984 29530 23984 0 FreeSans 1600 0 0 0 C10_3
port 466 nsew
flabel metal2 -51826 -9071 -51826 -9071 0 FreeSans 1600 0 0 0 C11_0
port 467 nsew
flabel metal1 -52275 -8285 -52275 -8285 0 FreeSans 1600 0 0 0 C11_1
port 468 nsew
flabel metal2 -52895 -8076 -52895 -8076 0 FreeSans 1600 0 0 0 C11_2
port 469 nsew
flabel metal2 -52273 -6853 -52273 -6853 0 FreeSans 1600 0 0 0 C11_3
port 470 nsew
flabel metal2 -31568 -5827 -31567 -5826 0 FreeSans 1600 0 0 0 C12_0
port 471 nsew
flabel metal1 -32011 -6604 -32011 -6604 0 FreeSans 1600 0 0 0 C12_1
port 472 nsew
flabel metal2 -32630 -6727 -32630 -6727 0 FreeSans 1600 0 0 0 C12_2
port 473 nsew
flabel metal2 -32018 -7976 -32018 -7976 0 FreeSans 1600 0 0 0 C12_3
port 474 nsew
flabel metal2 -2080 -5606 -2080 -5606 0 FreeSans 1600 0 0 0 C13_0
port 475 nsew
flabel metal1 -2535 -6605 -2535 -6605 0 FreeSans 1600 0 0 0 C13_1
port 476 nsew
flabel metal2 -3149 -6616 -3149 -6616 0 FreeSans 1600 0 0 0 C13_2
port 477 nsew
flabel metal2 -2529 -7765 -2529 -7765 0 FreeSans 1600 0 0 0 C13_3
port 478 nsew
flabel metal2 19316 -9034 19316 -9034 0 FreeSans 1600 0 0 0 C14_0
port 479 nsew
flabel metal1 18866 -8225 18866 -8225 0 FreeSans 1600 0 0 0 C14_1
port 480 nsew
flabel metal2 18259 -7966 18259 -7966 0 FreeSans 1600 0 0 0 C14_2
port 481 nsew
flabel metal2 18866 -6880 18866 -6880 0 FreeSans 1600 0 0 0 C14_3
port 482 nsew
flabel metal2 30008 -9084 30008 -9084 0 FreeSans 1600 0 0 0 C15_0
port 483 nsew
flabel metal1 29555 -8290 29555 -8290 0 FreeSans 1600 0 0 0 C15_1
port 484 nsew
flabel metal2 28940 -8093 28940 -8093 0 FreeSans 1600 0 0 0 C15_2
port 485 nsew
flabel metal2 29550 -6929 29550 -6929 0 FreeSans 1600 0 0 0 C15_3
port 486 nsew
flabel metal2 -51783 -14187 -51783 -14187 0 FreeSans 1600 0 0 0 C16_0
port 487 nsew
flabel metal1 -52226 -15204 -52226 -15204 0 FreeSans 1600 0 0 0 C16_1
port 488 nsew
flabel metal2 -52826 -15181 -52826 -15181 0 FreeSans 1600 0 0 0 C16_2
port 489 nsew
flabel metal2 -52236 -16349 -52236 -16349 0 FreeSans 1600 0 0 0 C16_3
port 490 nsew
flabel metal2 -30208 -25963 -30208 -25963 0 FreeSans 1600 0 0 0 C17_0
port 491 nsew
flabel metal1 -30655 -25166 -30655 -25166 0 FreeSans 1600 0 0 0 C17_1
port 492 nsew
flabel metal2 -31270 -24898 -31270 -24898 0 FreeSans 1600 0 0 0 C17_2
port 493 nsew
flabel metal2 -30656 -23822 -30656 -23822 0 FreeSans 1600 0 0 0 C17_3
port 494 nsew
flabel metal2 -2052 -25929 -2052 -25929 0 FreeSans 1600 0 0 0 C18_0
port 495 nsew
flabel metal1 -2488 -25136 -2488 -25136 0 FreeSans 1600 0 0 0 C18_1
port 496 nsew
flabel metal2 -3096 -24959 -3096 -24959 0 FreeSans 1600 0 0 0 C18_2
port 497 nsew
flabel metal2 -2491 -23783 -2491 -23783 0 FreeSans 1600 0 0 0 C18_3
port 498 nsew
flabel metal2 -30167 -34271 -30167 -34271 0 FreeSans 1600 0 0 0 C19_0
port 499 nsew
flabel metal1 -30615 -33463 -30615 -33463 0 FreeSans 1600 0 0 0 C19_1
port 500 nsew
flabel metal2 -31237 -33264 -31237 -33264 0 FreeSans 1600 0 0 0 C19_2
port 501 nsew
flabel metal2 -30614 -32122 -30614 -32122 0 FreeSans 1600 0 0 0 C19_3
port 502 nsew
flabel metal2 8641 -34386 8641 -34386 0 FreeSans 1600 0 0 0 C20_0
port 503 nsew
flabel metal1 8187 -33590 8187 -33590 0 FreeSans 1600 0 0 0 C20_1
port 504 nsew
flabel metal2 7573 -33459 7573 -33459 0 FreeSans 1600 0 0 0 C20_2
port 505 nsew
flabel metal2 8196 -32239 8196 -32239 0 FreeSans 1600 0 0 0 C20_3
port 506 nsew
flabel metal1 -71862 12311 -71862 12311 0 FreeSans 1600 0 0 0 G_source_dn
port 508 nsew
flabel metal1 -72117 18325 -72117 18325 0 FreeSans 1600 0 0 0 ITAIL_TOP
port 509 nsew
flabel metal1 9471 41606 9471 41606 0 FreeSans 1600 0 0 0 QB9
port 510 nsew
flabel metal1 -21802 7446 -21802 7446 0 FreeSans 1600 0 0 0 B1D
port 512 nsew
flabel metal1 -21827 4862 -21827 4862 0 FreeSans 1600 0 0 0 B4D
port 513 nsew
flabel metal1 -63456 38012 -63456 38012 0 FreeSans 1600 0 0 0 R0
port 514 nsew
flabel metal1 -63073 40896 -63073 40896 0 FreeSans 1600 0 0 0 R4
port 515 nsew
flabel metal1 -71884 12519 -71884 12519 0 FreeSans 1600 0 0 0 G_source_up
port 507 nsew
flabel metal1 -71339 10064 -71339 10064 0 FreeSans 1600 0 0 0 B1
port 517 nsew
<< end >>
