magic
tech gf180mcuC
magscale 1 10
timestamp 1699960019
<< nwell >>
rect -10910 -1423 -10506 -672
rect 2718 -8715 9137 -3142
rect 20948 -10345 27414 -1631
<< psubdiff >>
rect -10866 -4411 -10577 -4388
rect -10866 -4457 -10837 -4411
rect -10791 -4457 -10743 -4411
rect -10697 -4457 -10649 -4411
rect -10603 -4457 -10577 -4411
rect -10866 -4490 -10577 -4457
<< nsubdiff >>
rect -10827 -764 -10620 -733
rect -10827 -810 -10783 -764
rect -10737 -810 -10689 -764
rect -10643 -810 -10620 -764
rect -10827 -882 -10620 -810
rect -10827 -928 -10784 -882
rect -10738 -928 -10690 -882
rect -10644 -928 -10620 -882
rect -10827 -952 -10620 -928
rect 20984 -1697 27354 -1684
rect 20984 -1743 20997 -1697
rect 21043 -1743 21091 -1697
rect 21137 -1743 21185 -1697
rect 21231 -1743 21279 -1697
rect 21325 -1743 21373 -1697
rect 21419 -1743 21467 -1697
rect 21513 -1743 21561 -1697
rect 21607 -1743 21655 -1697
rect 21701 -1743 21749 -1697
rect 21795 -1743 21843 -1697
rect 21889 -1743 21937 -1697
rect 21983 -1743 22031 -1697
rect 22077 -1743 22125 -1697
rect 22171 -1743 22219 -1697
rect 22265 -1743 22313 -1697
rect 22359 -1743 22407 -1697
rect 22453 -1743 22501 -1697
rect 22547 -1743 22595 -1697
rect 22641 -1743 22689 -1697
rect 22735 -1743 22783 -1697
rect 22829 -1743 22877 -1697
rect 22923 -1743 22971 -1697
rect 23017 -1743 23065 -1697
rect 23111 -1743 23159 -1697
rect 23205 -1743 23253 -1697
rect 23299 -1743 23347 -1697
rect 23393 -1743 23441 -1697
rect 23487 -1743 23535 -1697
rect 23581 -1743 23629 -1697
rect 23675 -1743 23723 -1697
rect 23769 -1743 23817 -1697
rect 23863 -1743 23911 -1697
rect 23957 -1743 24005 -1697
rect 24051 -1743 24099 -1697
rect 24145 -1743 24193 -1697
rect 24239 -1743 24287 -1697
rect 24333 -1743 24381 -1697
rect 24427 -1743 24475 -1697
rect 24521 -1743 24569 -1697
rect 24615 -1743 24663 -1697
rect 24709 -1743 24757 -1697
rect 24803 -1743 24851 -1697
rect 24897 -1743 24945 -1697
rect 24991 -1743 25039 -1697
rect 25085 -1743 25133 -1697
rect 25179 -1743 25227 -1697
rect 25273 -1743 25321 -1697
rect 25367 -1743 25415 -1697
rect 25461 -1743 25509 -1697
rect 25555 -1743 25603 -1697
rect 25649 -1743 25697 -1697
rect 25743 -1743 25791 -1697
rect 25837 -1743 25885 -1697
rect 25931 -1743 25979 -1697
rect 26025 -1743 26073 -1697
rect 26119 -1743 26167 -1697
rect 26213 -1743 26261 -1697
rect 26307 -1743 26355 -1697
rect 26401 -1743 26449 -1697
rect 26495 -1743 26543 -1697
rect 26589 -1743 26637 -1697
rect 26683 -1743 26731 -1697
rect 26777 -1743 26825 -1697
rect 26871 -1743 26919 -1697
rect 26965 -1743 27013 -1697
rect 27059 -1743 27107 -1697
rect 27153 -1743 27201 -1697
rect 27247 -1743 27295 -1697
rect 27341 -1743 27354 -1697
rect 20984 -1756 27354 -1743
rect 20984 -1791 21056 -1756
rect 20984 -1837 20997 -1791
rect 21043 -1837 21056 -1791
rect 20984 -1885 21056 -1837
rect 20984 -1931 20997 -1885
rect 21043 -1931 21056 -1885
rect 20984 -1979 21056 -1931
rect 20984 -2025 20997 -1979
rect 21043 -2025 21056 -1979
rect 20984 -2073 21056 -2025
rect 20984 -2119 20997 -2073
rect 21043 -2119 21056 -2073
rect 20984 -2167 21056 -2119
rect 20984 -2213 20997 -2167
rect 21043 -2213 21056 -2167
rect 20984 -2261 21056 -2213
rect 20984 -2307 20997 -2261
rect 21043 -2307 21056 -2261
rect 20984 -2355 21056 -2307
rect 20984 -2401 20997 -2355
rect 21043 -2401 21056 -2355
rect 20984 -2449 21056 -2401
rect 20984 -2495 20997 -2449
rect 21043 -2495 21056 -2449
rect 20984 -2543 21056 -2495
rect 20984 -2589 20997 -2543
rect 21043 -2589 21056 -2543
rect 20984 -2637 21056 -2589
rect 20984 -2683 20997 -2637
rect 21043 -2683 21056 -2637
rect 20984 -2731 21056 -2683
rect 20984 -2777 20997 -2731
rect 21043 -2777 21056 -2731
rect 20984 -2825 21056 -2777
rect 20984 -2871 20997 -2825
rect 21043 -2871 21056 -2825
rect 20984 -2919 21056 -2871
rect 20984 -2965 20997 -2919
rect 21043 -2965 21056 -2919
rect 20984 -3013 21056 -2965
rect 20984 -3059 20997 -3013
rect 21043 -3059 21056 -3013
rect 20984 -3107 21056 -3059
rect 20984 -3153 20997 -3107
rect 21043 -3153 21056 -3107
rect 2743 -3180 9113 -3167
rect 2743 -3226 2756 -3180
rect 2802 -3226 2850 -3180
rect 2896 -3226 2944 -3180
rect 2990 -3226 3038 -3180
rect 3084 -3226 3132 -3180
rect 3178 -3226 3226 -3180
rect 3272 -3226 3320 -3180
rect 3366 -3226 3414 -3180
rect 3460 -3226 3508 -3180
rect 3554 -3226 3602 -3180
rect 3648 -3226 3696 -3180
rect 3742 -3226 3790 -3180
rect 3836 -3226 3884 -3180
rect 3930 -3226 3978 -3180
rect 4024 -3226 4072 -3180
rect 4118 -3226 4166 -3180
rect 4212 -3226 4260 -3180
rect 4306 -3226 4354 -3180
rect 4400 -3226 4448 -3180
rect 4494 -3226 4542 -3180
rect 4588 -3226 4636 -3180
rect 4682 -3226 4730 -3180
rect 4776 -3226 4824 -3180
rect 4870 -3226 4918 -3180
rect 4964 -3226 5012 -3180
rect 5058 -3226 5106 -3180
rect 5152 -3226 5200 -3180
rect 5246 -3226 5294 -3180
rect 5340 -3226 5388 -3180
rect 5434 -3226 5482 -3180
rect 5528 -3226 5576 -3180
rect 5622 -3226 5670 -3180
rect 5716 -3226 5764 -3180
rect 5810 -3226 5858 -3180
rect 5904 -3226 5952 -3180
rect 5998 -3226 6046 -3180
rect 6092 -3226 6140 -3180
rect 6186 -3226 6234 -3180
rect 6280 -3226 6328 -3180
rect 6374 -3226 6422 -3180
rect 6468 -3226 6516 -3180
rect 6562 -3226 6610 -3180
rect 6656 -3226 6704 -3180
rect 6750 -3226 6798 -3180
rect 6844 -3226 6892 -3180
rect 6938 -3226 6986 -3180
rect 7032 -3226 7080 -3180
rect 7126 -3226 7174 -3180
rect 7220 -3226 7268 -3180
rect 7314 -3226 7362 -3180
rect 7408 -3226 7456 -3180
rect 7502 -3226 7550 -3180
rect 7596 -3226 7644 -3180
rect 7690 -3226 7738 -3180
rect 7784 -3226 7832 -3180
rect 7878 -3226 7926 -3180
rect 7972 -3226 8020 -3180
rect 8066 -3226 8114 -3180
rect 8160 -3226 8208 -3180
rect 8254 -3226 8302 -3180
rect 8348 -3226 8396 -3180
rect 8442 -3226 8490 -3180
rect 8536 -3226 8584 -3180
rect 8630 -3226 8678 -3180
rect 8724 -3226 8772 -3180
rect 8818 -3226 8866 -3180
rect 8912 -3226 8960 -3180
rect 9006 -3226 9054 -3180
rect 9100 -3226 9113 -3180
rect 2743 -3239 9113 -3226
rect 2743 -3274 2815 -3239
rect 2743 -3320 2756 -3274
rect 2802 -3320 2815 -3274
rect 2743 -3368 2815 -3320
rect 2743 -3414 2756 -3368
rect 2802 -3414 2815 -3368
rect 2743 -3462 2815 -3414
rect 2743 -3508 2756 -3462
rect 2802 -3508 2815 -3462
rect 2743 -3556 2815 -3508
rect 2743 -3602 2756 -3556
rect 2802 -3602 2815 -3556
rect 2743 -3650 2815 -3602
rect 2743 -3696 2756 -3650
rect 2802 -3696 2815 -3650
rect 2743 -3744 2815 -3696
rect 2743 -3790 2756 -3744
rect 2802 -3790 2815 -3744
rect 2743 -3838 2815 -3790
rect 2743 -3884 2756 -3838
rect 2802 -3884 2815 -3838
rect 2743 -3932 2815 -3884
rect 2743 -3978 2756 -3932
rect 2802 -3978 2815 -3932
rect 2743 -4026 2815 -3978
rect 2743 -4072 2756 -4026
rect 2802 -4072 2815 -4026
rect 2743 -4120 2815 -4072
rect 2743 -4166 2756 -4120
rect 2802 -4166 2815 -4120
rect 2743 -4214 2815 -4166
rect 2743 -4260 2756 -4214
rect 2802 -4260 2815 -4214
rect 2743 -4308 2815 -4260
rect 2743 -4354 2756 -4308
rect 2802 -4354 2815 -4308
rect 2743 -4402 2815 -4354
rect 2743 -4448 2756 -4402
rect 2802 -4448 2815 -4402
rect 2743 -4496 2815 -4448
rect 2743 -4542 2756 -4496
rect 2802 -4542 2815 -4496
rect 2743 -4590 2815 -4542
rect 2743 -4636 2756 -4590
rect 2802 -4636 2815 -4590
rect 2743 -4684 2815 -4636
rect 2743 -4730 2756 -4684
rect 2802 -4730 2815 -4684
rect 2743 -4778 2815 -4730
rect 2743 -4824 2756 -4778
rect 2802 -4824 2815 -4778
rect 2743 -4872 2815 -4824
rect 2743 -4918 2756 -4872
rect 2802 -4918 2815 -4872
rect 2743 -4966 2815 -4918
rect 2743 -5012 2756 -4966
rect 2802 -5012 2815 -4966
rect 2743 -5060 2815 -5012
rect 2743 -5106 2756 -5060
rect 2802 -5106 2815 -5060
rect 2743 -5154 2815 -5106
rect 2743 -5200 2756 -5154
rect 2802 -5200 2815 -5154
rect 2743 -5248 2815 -5200
rect 2743 -5294 2756 -5248
rect 2802 -5294 2815 -5248
rect 2743 -5342 2815 -5294
rect 2743 -5388 2756 -5342
rect 2802 -5388 2815 -5342
rect 2743 -5436 2815 -5388
rect 2743 -5482 2756 -5436
rect 2802 -5482 2815 -5436
rect 2743 -5530 2815 -5482
rect 2743 -5576 2756 -5530
rect 2802 -5576 2815 -5530
rect 2743 -5624 2815 -5576
rect 2743 -5670 2756 -5624
rect 2802 -5670 2815 -5624
rect 2743 -5718 2815 -5670
rect 2743 -5764 2756 -5718
rect 2802 -5764 2815 -5718
rect 2743 -5812 2815 -5764
rect 2743 -5858 2756 -5812
rect 2802 -5858 2815 -5812
rect 2743 -5906 2815 -5858
rect 2743 -5952 2756 -5906
rect 2802 -5952 2815 -5906
rect 2743 -6000 2815 -5952
rect 2743 -6046 2756 -6000
rect 2802 -6046 2815 -6000
rect 2743 -6094 2815 -6046
rect 2743 -6140 2756 -6094
rect 2802 -6140 2815 -6094
rect 2743 -6188 2815 -6140
rect 2743 -6234 2756 -6188
rect 2802 -6234 2815 -6188
rect 2743 -6282 2815 -6234
rect 2743 -6328 2756 -6282
rect 2802 -6328 2815 -6282
rect 2743 -6376 2815 -6328
rect 2743 -6422 2756 -6376
rect 2802 -6422 2815 -6376
rect 2743 -6470 2815 -6422
rect 2743 -6516 2756 -6470
rect 2802 -6516 2815 -6470
rect 2743 -6564 2815 -6516
rect 2743 -6610 2756 -6564
rect 2802 -6610 2815 -6564
rect 2743 -6658 2815 -6610
rect 2743 -6704 2756 -6658
rect 2802 -6704 2815 -6658
rect 2743 -6752 2815 -6704
rect 2743 -6798 2756 -6752
rect 2802 -6798 2815 -6752
rect 2743 -6846 2815 -6798
rect 2743 -6892 2756 -6846
rect 2802 -6892 2815 -6846
rect 2743 -6940 2815 -6892
rect 2743 -6986 2756 -6940
rect 2802 -6986 2815 -6940
rect 2743 -7034 2815 -6986
rect 2743 -7080 2756 -7034
rect 2802 -7080 2815 -7034
rect 2743 -7128 2815 -7080
rect 2743 -7174 2756 -7128
rect 2802 -7174 2815 -7128
rect 2743 -7222 2815 -7174
rect 2743 -7268 2756 -7222
rect 2802 -7268 2815 -7222
rect 2743 -7316 2815 -7268
rect 2743 -7362 2756 -7316
rect 2802 -7362 2815 -7316
rect 2743 -7410 2815 -7362
rect 2743 -7456 2756 -7410
rect 2802 -7456 2815 -7410
rect 2743 -7504 2815 -7456
rect 2743 -7550 2756 -7504
rect 2802 -7550 2815 -7504
rect 2743 -7598 2815 -7550
rect 2743 -7644 2756 -7598
rect 2802 -7644 2815 -7598
rect 2743 -7692 2815 -7644
rect 2743 -7738 2756 -7692
rect 2802 -7738 2815 -7692
rect 2743 -7786 2815 -7738
rect 2743 -7832 2756 -7786
rect 2802 -7832 2815 -7786
rect 2743 -7880 2815 -7832
rect 2743 -7926 2756 -7880
rect 2802 -7926 2815 -7880
rect 2743 -7974 2815 -7926
rect 2743 -8020 2756 -7974
rect 2802 -8020 2815 -7974
rect 2743 -8068 2815 -8020
rect 2743 -8114 2756 -8068
rect 2802 -8114 2815 -8068
rect 2743 -8162 2815 -8114
rect 2743 -8208 2756 -8162
rect 2802 -8208 2815 -8162
rect 2743 -8256 2815 -8208
rect 2743 -8302 2756 -8256
rect 2802 -8302 2815 -8256
rect 2743 -8350 2815 -8302
rect 2743 -8396 2756 -8350
rect 2802 -8396 2815 -8350
rect 2743 -8444 2815 -8396
rect 2743 -8490 2756 -8444
rect 2802 -8490 2815 -8444
rect 2743 -8538 2815 -8490
rect 2743 -8584 2756 -8538
rect 2802 -8584 2815 -8538
rect 2743 -8619 2815 -8584
rect 9041 -3274 9113 -3239
rect 9041 -3320 9054 -3274
rect 9100 -3320 9113 -3274
rect 9041 -3368 9113 -3320
rect 9041 -3414 9054 -3368
rect 9100 -3414 9113 -3368
rect 9041 -3462 9113 -3414
rect 9041 -3508 9054 -3462
rect 9100 -3508 9113 -3462
rect 9041 -3556 9113 -3508
rect 9041 -3602 9054 -3556
rect 9100 -3602 9113 -3556
rect 9041 -3650 9113 -3602
rect 9041 -3696 9054 -3650
rect 9100 -3696 9113 -3650
rect 9041 -3744 9113 -3696
rect 9041 -3790 9054 -3744
rect 9100 -3790 9113 -3744
rect 9041 -3838 9113 -3790
rect 9041 -3884 9054 -3838
rect 9100 -3884 9113 -3838
rect 9041 -3932 9113 -3884
rect 9041 -3978 9054 -3932
rect 9100 -3978 9113 -3932
rect 9041 -4026 9113 -3978
rect 9041 -4072 9054 -4026
rect 9100 -4072 9113 -4026
rect 9041 -4120 9113 -4072
rect 9041 -4166 9054 -4120
rect 9100 -4166 9113 -4120
rect 9041 -4214 9113 -4166
rect 9041 -4260 9054 -4214
rect 9100 -4260 9113 -4214
rect 9041 -4308 9113 -4260
rect 9041 -4354 9054 -4308
rect 9100 -4354 9113 -4308
rect 9041 -4402 9113 -4354
rect 9041 -4448 9054 -4402
rect 9100 -4448 9113 -4402
rect 9041 -4496 9113 -4448
rect 9041 -4542 9054 -4496
rect 9100 -4542 9113 -4496
rect 9041 -4590 9113 -4542
rect 9041 -4636 9054 -4590
rect 9100 -4636 9113 -4590
rect 9041 -4684 9113 -4636
rect 9041 -4730 9054 -4684
rect 9100 -4730 9113 -4684
rect 9041 -4778 9113 -4730
rect 9041 -4824 9054 -4778
rect 9100 -4824 9113 -4778
rect 9041 -4872 9113 -4824
rect 9041 -4918 9054 -4872
rect 9100 -4918 9113 -4872
rect 9041 -4966 9113 -4918
rect 9041 -5012 9054 -4966
rect 9100 -5012 9113 -4966
rect 9041 -5060 9113 -5012
rect 9041 -5106 9054 -5060
rect 9100 -5106 9113 -5060
rect 9041 -5154 9113 -5106
rect 9041 -5200 9054 -5154
rect 9100 -5200 9113 -5154
rect 9041 -5248 9113 -5200
rect 9041 -5294 9054 -5248
rect 9100 -5294 9113 -5248
rect 9041 -5342 9113 -5294
rect 9041 -5388 9054 -5342
rect 9100 -5388 9113 -5342
rect 9041 -5436 9113 -5388
rect 9041 -5482 9054 -5436
rect 9100 -5482 9113 -5436
rect 9041 -5530 9113 -5482
rect 9041 -5576 9054 -5530
rect 9100 -5576 9113 -5530
rect 9041 -5624 9113 -5576
rect 9041 -5670 9054 -5624
rect 9100 -5670 9113 -5624
rect 9041 -5718 9113 -5670
rect 9041 -5764 9054 -5718
rect 9100 -5764 9113 -5718
rect 9041 -5812 9113 -5764
rect 9041 -5858 9054 -5812
rect 9100 -5858 9113 -5812
rect 9041 -5906 9113 -5858
rect 9041 -5952 9054 -5906
rect 9100 -5952 9113 -5906
rect 9041 -6000 9113 -5952
rect 9041 -6046 9054 -6000
rect 9100 -6046 9113 -6000
rect 9041 -6094 9113 -6046
rect 9041 -6140 9054 -6094
rect 9100 -6140 9113 -6094
rect 9041 -6188 9113 -6140
rect 9041 -6234 9054 -6188
rect 9100 -6234 9113 -6188
rect 9041 -6282 9113 -6234
rect 9041 -6328 9054 -6282
rect 9100 -6328 9113 -6282
rect 9041 -6376 9113 -6328
rect 9041 -6422 9054 -6376
rect 9100 -6422 9113 -6376
rect 9041 -6470 9113 -6422
rect 9041 -6516 9054 -6470
rect 9100 -6516 9113 -6470
rect 9041 -6564 9113 -6516
rect 9041 -6610 9054 -6564
rect 9100 -6610 9113 -6564
rect 9041 -6658 9113 -6610
rect 9041 -6704 9054 -6658
rect 9100 -6704 9113 -6658
rect 9041 -6752 9113 -6704
rect 9041 -6798 9054 -6752
rect 9100 -6798 9113 -6752
rect 9041 -6846 9113 -6798
rect 9041 -6892 9054 -6846
rect 9100 -6892 9113 -6846
rect 9041 -6940 9113 -6892
rect 9041 -6986 9054 -6940
rect 9100 -6986 9113 -6940
rect 9041 -7034 9113 -6986
rect 9041 -7080 9054 -7034
rect 9100 -7080 9113 -7034
rect 9041 -7128 9113 -7080
rect 9041 -7174 9054 -7128
rect 9100 -7174 9113 -7128
rect 9041 -7222 9113 -7174
rect 9041 -7268 9054 -7222
rect 9100 -7268 9113 -7222
rect 9041 -7316 9113 -7268
rect 9041 -7362 9054 -7316
rect 9100 -7362 9113 -7316
rect 9041 -7410 9113 -7362
rect 9041 -7456 9054 -7410
rect 9100 -7456 9113 -7410
rect 9041 -7504 9113 -7456
rect 9041 -7550 9054 -7504
rect 9100 -7550 9113 -7504
rect 9041 -7598 9113 -7550
rect 9041 -7644 9054 -7598
rect 9100 -7644 9113 -7598
rect 9041 -7692 9113 -7644
rect 9041 -7738 9054 -7692
rect 9100 -7738 9113 -7692
rect 9041 -7786 9113 -7738
rect 9041 -7832 9054 -7786
rect 9100 -7832 9113 -7786
rect 9041 -7880 9113 -7832
rect 9041 -7926 9054 -7880
rect 9100 -7926 9113 -7880
rect 9041 -7974 9113 -7926
rect 9041 -8020 9054 -7974
rect 9100 -8020 9113 -7974
rect 9041 -8068 9113 -8020
rect 9041 -8114 9054 -8068
rect 9100 -8114 9113 -8068
rect 9041 -8162 9113 -8114
rect 9041 -8208 9054 -8162
rect 9100 -8208 9113 -8162
rect 9041 -8256 9113 -8208
rect 9041 -8302 9054 -8256
rect 9100 -8302 9113 -8256
rect 9041 -8350 9113 -8302
rect 9041 -8396 9054 -8350
rect 9100 -8396 9113 -8350
rect 9041 -8444 9113 -8396
rect 9041 -8490 9054 -8444
rect 9100 -8490 9113 -8444
rect 9041 -8538 9113 -8490
rect 9041 -8584 9054 -8538
rect 9100 -8584 9113 -8538
rect 9041 -8619 9113 -8584
rect 2743 -8632 9113 -8619
rect 2743 -8678 2756 -8632
rect 2802 -8678 2850 -8632
rect 2896 -8678 2944 -8632
rect 2990 -8678 3038 -8632
rect 3084 -8678 3132 -8632
rect 3178 -8678 3226 -8632
rect 3272 -8678 3320 -8632
rect 3366 -8678 3414 -8632
rect 3460 -8678 3508 -8632
rect 3554 -8678 3602 -8632
rect 3648 -8678 3696 -8632
rect 3742 -8678 3790 -8632
rect 3836 -8678 3884 -8632
rect 3930 -8678 3978 -8632
rect 4024 -8678 4072 -8632
rect 4118 -8678 4166 -8632
rect 4212 -8678 4260 -8632
rect 4306 -8678 4354 -8632
rect 4400 -8678 4448 -8632
rect 4494 -8678 4542 -8632
rect 4588 -8678 4636 -8632
rect 4682 -8678 4730 -8632
rect 4776 -8678 4824 -8632
rect 4870 -8678 4918 -8632
rect 4964 -8678 5012 -8632
rect 5058 -8678 5106 -8632
rect 5152 -8678 5200 -8632
rect 5246 -8678 5294 -8632
rect 5340 -8678 5388 -8632
rect 5434 -8678 5482 -8632
rect 5528 -8678 5576 -8632
rect 5622 -8678 5670 -8632
rect 5716 -8678 5764 -8632
rect 5810 -8678 5858 -8632
rect 5904 -8678 5952 -8632
rect 5998 -8678 6046 -8632
rect 6092 -8678 6140 -8632
rect 6186 -8678 6234 -8632
rect 6280 -8678 6328 -8632
rect 6374 -8678 6422 -8632
rect 6468 -8678 6516 -8632
rect 6562 -8678 6610 -8632
rect 6656 -8678 6704 -8632
rect 6750 -8678 6798 -8632
rect 6844 -8678 6892 -8632
rect 6938 -8678 6986 -8632
rect 7032 -8678 7080 -8632
rect 7126 -8678 7174 -8632
rect 7220 -8678 7268 -8632
rect 7314 -8678 7362 -8632
rect 7408 -8678 7456 -8632
rect 7502 -8678 7550 -8632
rect 7596 -8678 7644 -8632
rect 7690 -8678 7738 -8632
rect 7784 -8678 7832 -8632
rect 7878 -8678 7926 -8632
rect 7972 -8678 8020 -8632
rect 8066 -8678 8114 -8632
rect 8160 -8678 8208 -8632
rect 8254 -8678 8302 -8632
rect 8348 -8678 8396 -8632
rect 8442 -8678 8490 -8632
rect 8536 -8678 8584 -8632
rect 8630 -8678 8678 -8632
rect 8724 -8678 8772 -8632
rect 8818 -8678 8866 -8632
rect 8912 -8678 8960 -8632
rect 9006 -8678 9054 -8632
rect 9100 -8678 9113 -8632
rect 2743 -8691 9113 -8678
rect 20984 -3201 21056 -3153
rect 20984 -3247 20997 -3201
rect 21043 -3247 21056 -3201
rect 20984 -3295 21056 -3247
rect 20984 -3341 20997 -3295
rect 21043 -3341 21056 -3295
rect 20984 -3389 21056 -3341
rect 20984 -3435 20997 -3389
rect 21043 -3435 21056 -3389
rect 20984 -3483 21056 -3435
rect 20984 -3529 20997 -3483
rect 21043 -3529 21056 -3483
rect 20984 -3577 21056 -3529
rect 20984 -3623 20997 -3577
rect 21043 -3623 21056 -3577
rect 20984 -3671 21056 -3623
rect 20984 -3717 20997 -3671
rect 21043 -3717 21056 -3671
rect 20984 -3765 21056 -3717
rect 20984 -3811 20997 -3765
rect 21043 -3811 21056 -3765
rect 20984 -3859 21056 -3811
rect 20984 -3905 20997 -3859
rect 21043 -3905 21056 -3859
rect 20984 -3953 21056 -3905
rect 20984 -3999 20997 -3953
rect 21043 -3999 21056 -3953
rect 20984 -4047 21056 -3999
rect 20984 -4093 20997 -4047
rect 21043 -4093 21056 -4047
rect 20984 -4141 21056 -4093
rect 20984 -4187 20997 -4141
rect 21043 -4187 21056 -4141
rect 20984 -4235 21056 -4187
rect 20984 -4281 20997 -4235
rect 21043 -4281 21056 -4235
rect 20984 -4329 21056 -4281
rect 20984 -4375 20997 -4329
rect 21043 -4375 21056 -4329
rect 20984 -4423 21056 -4375
rect 20984 -4469 20997 -4423
rect 21043 -4469 21056 -4423
rect 20984 -4517 21056 -4469
rect 20984 -4563 20997 -4517
rect 21043 -4563 21056 -4517
rect 20984 -4611 21056 -4563
rect 20984 -4657 20997 -4611
rect 21043 -4657 21056 -4611
rect 20984 -4705 21056 -4657
rect 20984 -4751 20997 -4705
rect 21043 -4751 21056 -4705
rect 20984 -4799 21056 -4751
rect 20984 -4845 20997 -4799
rect 21043 -4845 21056 -4799
rect 20984 -4893 21056 -4845
rect 20984 -4939 20997 -4893
rect 21043 -4939 21056 -4893
rect 20984 -4987 21056 -4939
rect 20984 -5033 20997 -4987
rect 21043 -5033 21056 -4987
rect 20984 -5081 21056 -5033
rect 20984 -5127 20997 -5081
rect 21043 -5127 21056 -5081
rect 20984 -5175 21056 -5127
rect 20984 -5221 20997 -5175
rect 21043 -5221 21056 -5175
rect 20984 -5269 21056 -5221
rect 20984 -5315 20997 -5269
rect 21043 -5315 21056 -5269
rect 20984 -5363 21056 -5315
rect 20984 -5409 20997 -5363
rect 21043 -5409 21056 -5363
rect 20984 -5457 21056 -5409
rect 20984 -5503 20997 -5457
rect 21043 -5503 21056 -5457
rect 20984 -5551 21056 -5503
rect 20984 -5597 20997 -5551
rect 21043 -5597 21056 -5551
rect 20984 -5645 21056 -5597
rect 20984 -5691 20997 -5645
rect 21043 -5691 21056 -5645
rect 20984 -5739 21056 -5691
rect 20984 -5785 20997 -5739
rect 21043 -5785 21056 -5739
rect 20984 -5833 21056 -5785
rect 20984 -5879 20997 -5833
rect 21043 -5879 21056 -5833
rect 20984 -5927 21056 -5879
rect 20984 -5973 20997 -5927
rect 21043 -5973 21056 -5927
rect 20984 -6021 21056 -5973
rect 20984 -6067 20997 -6021
rect 21043 -6067 21056 -6021
rect 20984 -6115 21056 -6067
rect 20984 -6161 20997 -6115
rect 21043 -6161 21056 -6115
rect 20984 -6209 21056 -6161
rect 20984 -6255 20997 -6209
rect 21043 -6255 21056 -6209
rect 20984 -6303 21056 -6255
rect 20984 -6349 20997 -6303
rect 21043 -6349 21056 -6303
rect 20984 -6397 21056 -6349
rect 20984 -6443 20997 -6397
rect 21043 -6443 21056 -6397
rect 20984 -6491 21056 -6443
rect 20984 -6537 20997 -6491
rect 21043 -6537 21056 -6491
rect 20984 -6585 21056 -6537
rect 20984 -6631 20997 -6585
rect 21043 -6631 21056 -6585
rect 20984 -6679 21056 -6631
rect 20984 -6725 20997 -6679
rect 21043 -6725 21056 -6679
rect 20984 -6773 21056 -6725
rect 20984 -6819 20997 -6773
rect 21043 -6819 21056 -6773
rect 20984 -6867 21056 -6819
rect 20984 -6913 20997 -6867
rect 21043 -6913 21056 -6867
rect 20984 -6961 21056 -6913
rect 20984 -7007 20997 -6961
rect 21043 -7007 21056 -6961
rect 20984 -7055 21056 -7007
rect 20984 -7101 20997 -7055
rect 21043 -7101 21056 -7055
rect 20984 -7149 21056 -7101
rect 20984 -7195 20997 -7149
rect 21043 -7195 21056 -7149
rect 20984 -7243 21056 -7195
rect 20984 -7289 20997 -7243
rect 21043 -7289 21056 -7243
rect 20984 -7337 21056 -7289
rect 20984 -7383 20997 -7337
rect 21043 -7383 21056 -7337
rect 20984 -7431 21056 -7383
rect 20984 -7477 20997 -7431
rect 21043 -7477 21056 -7431
rect 20984 -7525 21056 -7477
rect 20984 -7571 20997 -7525
rect 21043 -7571 21056 -7525
rect 20984 -7619 21056 -7571
rect 20984 -7665 20997 -7619
rect 21043 -7665 21056 -7619
rect 20984 -7713 21056 -7665
rect 20984 -7759 20997 -7713
rect 21043 -7759 21056 -7713
rect 20984 -7807 21056 -7759
rect 20984 -7853 20997 -7807
rect 21043 -7853 21056 -7807
rect 20984 -7901 21056 -7853
rect 20984 -7947 20997 -7901
rect 21043 -7947 21056 -7901
rect 20984 -7995 21056 -7947
rect 20984 -8041 20997 -7995
rect 21043 -8041 21056 -7995
rect 20984 -8089 21056 -8041
rect 20984 -8135 20997 -8089
rect 21043 -8135 21056 -8089
rect 20984 -8183 21056 -8135
rect 20984 -8229 20997 -8183
rect 21043 -8229 21056 -8183
rect 20984 -8277 21056 -8229
rect 20984 -8323 20997 -8277
rect 21043 -8323 21056 -8277
rect 20984 -8371 21056 -8323
rect 20984 -8417 20997 -8371
rect 21043 -8417 21056 -8371
rect 20984 -8465 21056 -8417
rect 20984 -8511 20997 -8465
rect 21043 -8511 21056 -8465
rect 20984 -8559 21056 -8511
rect 20984 -8605 20997 -8559
rect 21043 -8605 21056 -8559
rect 20984 -8653 21056 -8605
rect 20984 -8699 20997 -8653
rect 21043 -8699 21056 -8653
rect 20984 -8747 21056 -8699
rect 20984 -8793 20997 -8747
rect 21043 -8793 21056 -8747
rect 20984 -8841 21056 -8793
rect 20984 -8887 20997 -8841
rect 21043 -8887 21056 -8841
rect 20984 -8935 21056 -8887
rect 20984 -8981 20997 -8935
rect 21043 -8981 21056 -8935
rect 20984 -9029 21056 -8981
rect 20984 -9075 20997 -9029
rect 21043 -9075 21056 -9029
rect 20984 -9123 21056 -9075
rect 20984 -9169 20997 -9123
rect 21043 -9169 21056 -9123
rect 20984 -9217 21056 -9169
rect 20984 -9263 20997 -9217
rect 21043 -9263 21056 -9217
rect 20984 -9311 21056 -9263
rect 20984 -9357 20997 -9311
rect 21043 -9357 21056 -9311
rect 20984 -9405 21056 -9357
rect 20984 -9451 20997 -9405
rect 21043 -9451 21056 -9405
rect 20984 -9499 21056 -9451
rect 20984 -9545 20997 -9499
rect 21043 -9545 21056 -9499
rect 20984 -9593 21056 -9545
rect 20984 -9639 20997 -9593
rect 21043 -9639 21056 -9593
rect 20984 -9687 21056 -9639
rect 20984 -9733 20997 -9687
rect 21043 -9733 21056 -9687
rect 20984 -9781 21056 -9733
rect 20984 -9827 20997 -9781
rect 21043 -9827 21056 -9781
rect 20984 -9875 21056 -9827
rect 20984 -9921 20997 -9875
rect 21043 -9921 21056 -9875
rect 20984 -9969 21056 -9921
rect 20984 -10015 20997 -9969
rect 21043 -10015 21056 -9969
rect 20984 -10063 21056 -10015
rect 20984 -10109 20997 -10063
rect 21043 -10109 21056 -10063
rect 20984 -10157 21056 -10109
rect 20984 -10203 20997 -10157
rect 21043 -10203 21056 -10157
rect 20984 -10238 21056 -10203
rect 27282 -1791 27354 -1756
rect 27282 -1837 27295 -1791
rect 27341 -1837 27354 -1791
rect 27282 -1885 27354 -1837
rect 27282 -1931 27295 -1885
rect 27341 -1931 27354 -1885
rect 27282 -1979 27354 -1931
rect 27282 -2025 27295 -1979
rect 27341 -2025 27354 -1979
rect 27282 -2073 27354 -2025
rect 27282 -2119 27295 -2073
rect 27341 -2119 27354 -2073
rect 27282 -2167 27354 -2119
rect 27282 -2213 27295 -2167
rect 27341 -2213 27354 -2167
rect 27282 -2261 27354 -2213
rect 27282 -2307 27295 -2261
rect 27341 -2307 27354 -2261
rect 27282 -2355 27354 -2307
rect 27282 -2401 27295 -2355
rect 27341 -2401 27354 -2355
rect 27282 -2449 27354 -2401
rect 27282 -2495 27295 -2449
rect 27341 -2495 27354 -2449
rect 27282 -2543 27354 -2495
rect 27282 -2589 27295 -2543
rect 27341 -2589 27354 -2543
rect 27282 -2637 27354 -2589
rect 27282 -2683 27295 -2637
rect 27341 -2683 27354 -2637
rect 27282 -2731 27354 -2683
rect 27282 -2777 27295 -2731
rect 27341 -2777 27354 -2731
rect 27282 -2825 27354 -2777
rect 27282 -2871 27295 -2825
rect 27341 -2871 27354 -2825
rect 27282 -2919 27354 -2871
rect 27282 -2965 27295 -2919
rect 27341 -2965 27354 -2919
rect 27282 -3013 27354 -2965
rect 27282 -3059 27295 -3013
rect 27341 -3059 27354 -3013
rect 27282 -3107 27354 -3059
rect 27282 -3153 27295 -3107
rect 27341 -3153 27354 -3107
rect 27282 -3201 27354 -3153
rect 27282 -3247 27295 -3201
rect 27341 -3247 27354 -3201
rect 27282 -3295 27354 -3247
rect 27282 -3341 27295 -3295
rect 27341 -3341 27354 -3295
rect 27282 -3389 27354 -3341
rect 27282 -3435 27295 -3389
rect 27341 -3435 27354 -3389
rect 27282 -3483 27354 -3435
rect 27282 -3529 27295 -3483
rect 27341 -3529 27354 -3483
rect 27282 -3577 27354 -3529
rect 27282 -3623 27295 -3577
rect 27341 -3623 27354 -3577
rect 27282 -3671 27354 -3623
rect 27282 -3717 27295 -3671
rect 27341 -3717 27354 -3671
rect 27282 -3765 27354 -3717
rect 27282 -3811 27295 -3765
rect 27341 -3811 27354 -3765
rect 27282 -3859 27354 -3811
rect 27282 -3905 27295 -3859
rect 27341 -3905 27354 -3859
rect 27282 -3953 27354 -3905
rect 27282 -3999 27295 -3953
rect 27341 -3999 27354 -3953
rect 27282 -4047 27354 -3999
rect 27282 -4093 27295 -4047
rect 27341 -4093 27354 -4047
rect 27282 -4141 27354 -4093
rect 27282 -4187 27295 -4141
rect 27341 -4187 27354 -4141
rect 27282 -4235 27354 -4187
rect 27282 -4281 27295 -4235
rect 27341 -4281 27354 -4235
rect 27282 -4329 27354 -4281
rect 27282 -4375 27295 -4329
rect 27341 -4375 27354 -4329
rect 27282 -4423 27354 -4375
rect 27282 -4469 27295 -4423
rect 27341 -4469 27354 -4423
rect 27282 -4517 27354 -4469
rect 27282 -4563 27295 -4517
rect 27341 -4563 27354 -4517
rect 27282 -4611 27354 -4563
rect 27282 -4657 27295 -4611
rect 27341 -4657 27354 -4611
rect 27282 -4705 27354 -4657
rect 27282 -4751 27295 -4705
rect 27341 -4751 27354 -4705
rect 27282 -4799 27354 -4751
rect 27282 -4845 27295 -4799
rect 27341 -4845 27354 -4799
rect 27282 -4893 27354 -4845
rect 27282 -4939 27295 -4893
rect 27341 -4939 27354 -4893
rect 27282 -4987 27354 -4939
rect 27282 -5033 27295 -4987
rect 27341 -5033 27354 -4987
rect 27282 -5081 27354 -5033
rect 27282 -5127 27295 -5081
rect 27341 -5127 27354 -5081
rect 27282 -5175 27354 -5127
rect 27282 -5221 27295 -5175
rect 27341 -5221 27354 -5175
rect 27282 -5269 27354 -5221
rect 27282 -5315 27295 -5269
rect 27341 -5315 27354 -5269
rect 27282 -5363 27354 -5315
rect 27282 -5409 27295 -5363
rect 27341 -5409 27354 -5363
rect 27282 -5457 27354 -5409
rect 27282 -5503 27295 -5457
rect 27341 -5503 27354 -5457
rect 27282 -5551 27354 -5503
rect 27282 -5597 27295 -5551
rect 27341 -5597 27354 -5551
rect 27282 -5645 27354 -5597
rect 27282 -5691 27295 -5645
rect 27341 -5691 27354 -5645
rect 27282 -5739 27354 -5691
rect 27282 -5785 27295 -5739
rect 27341 -5785 27354 -5739
rect 27282 -5833 27354 -5785
rect 27282 -5879 27295 -5833
rect 27341 -5879 27354 -5833
rect 27282 -5927 27354 -5879
rect 27282 -5973 27295 -5927
rect 27341 -5973 27354 -5927
rect 27282 -6021 27354 -5973
rect 27282 -6067 27295 -6021
rect 27341 -6067 27354 -6021
rect 27282 -6115 27354 -6067
rect 27282 -6161 27295 -6115
rect 27341 -6161 27354 -6115
rect 27282 -6209 27354 -6161
rect 27282 -6255 27295 -6209
rect 27341 -6255 27354 -6209
rect 27282 -6303 27354 -6255
rect 27282 -6349 27295 -6303
rect 27341 -6349 27354 -6303
rect 27282 -6397 27354 -6349
rect 27282 -6443 27295 -6397
rect 27341 -6443 27354 -6397
rect 27282 -6491 27354 -6443
rect 27282 -6537 27295 -6491
rect 27341 -6537 27354 -6491
rect 27282 -6585 27354 -6537
rect 27282 -6631 27295 -6585
rect 27341 -6631 27354 -6585
rect 27282 -6679 27354 -6631
rect 27282 -6725 27295 -6679
rect 27341 -6725 27354 -6679
rect 27282 -6773 27354 -6725
rect 27282 -6819 27295 -6773
rect 27341 -6819 27354 -6773
rect 27282 -6867 27354 -6819
rect 27282 -6913 27295 -6867
rect 27341 -6913 27354 -6867
rect 27282 -6961 27354 -6913
rect 27282 -7007 27295 -6961
rect 27341 -7007 27354 -6961
rect 27282 -7055 27354 -7007
rect 27282 -7101 27295 -7055
rect 27341 -7101 27354 -7055
rect 27282 -7149 27354 -7101
rect 27282 -7195 27295 -7149
rect 27341 -7195 27354 -7149
rect 27282 -7243 27354 -7195
rect 27282 -7289 27295 -7243
rect 27341 -7289 27354 -7243
rect 27282 -7337 27354 -7289
rect 27282 -7383 27295 -7337
rect 27341 -7383 27354 -7337
rect 27282 -7431 27354 -7383
rect 27282 -7477 27295 -7431
rect 27341 -7477 27354 -7431
rect 27282 -7525 27354 -7477
rect 27282 -7571 27295 -7525
rect 27341 -7571 27354 -7525
rect 27282 -7619 27354 -7571
rect 27282 -7665 27295 -7619
rect 27341 -7665 27354 -7619
rect 27282 -7713 27354 -7665
rect 27282 -7759 27295 -7713
rect 27341 -7759 27354 -7713
rect 27282 -7807 27354 -7759
rect 27282 -7853 27295 -7807
rect 27341 -7853 27354 -7807
rect 27282 -7901 27354 -7853
rect 27282 -7947 27295 -7901
rect 27341 -7947 27354 -7901
rect 27282 -7995 27354 -7947
rect 27282 -8041 27295 -7995
rect 27341 -8041 27354 -7995
rect 27282 -8089 27354 -8041
rect 27282 -8135 27295 -8089
rect 27341 -8135 27354 -8089
rect 27282 -8183 27354 -8135
rect 27282 -8229 27295 -8183
rect 27341 -8229 27354 -8183
rect 27282 -8277 27354 -8229
rect 27282 -8323 27295 -8277
rect 27341 -8323 27354 -8277
rect 27282 -8371 27354 -8323
rect 27282 -8417 27295 -8371
rect 27341 -8417 27354 -8371
rect 27282 -8465 27354 -8417
rect 27282 -8511 27295 -8465
rect 27341 -8511 27354 -8465
rect 27282 -8559 27354 -8511
rect 27282 -8605 27295 -8559
rect 27341 -8605 27354 -8559
rect 27282 -8653 27354 -8605
rect 27282 -8699 27295 -8653
rect 27341 -8699 27354 -8653
rect 27282 -8747 27354 -8699
rect 27282 -8793 27295 -8747
rect 27341 -8793 27354 -8747
rect 27282 -8841 27354 -8793
rect 27282 -8887 27295 -8841
rect 27341 -8887 27354 -8841
rect 27282 -8935 27354 -8887
rect 27282 -8981 27295 -8935
rect 27341 -8981 27354 -8935
rect 27282 -9029 27354 -8981
rect 27282 -9075 27295 -9029
rect 27341 -9075 27354 -9029
rect 27282 -9123 27354 -9075
rect 27282 -9169 27295 -9123
rect 27341 -9169 27354 -9123
rect 27282 -9217 27354 -9169
rect 27282 -9263 27295 -9217
rect 27341 -9263 27354 -9217
rect 27282 -9311 27354 -9263
rect 27282 -9357 27295 -9311
rect 27341 -9357 27354 -9311
rect 27282 -9405 27354 -9357
rect 27282 -9451 27295 -9405
rect 27341 -9451 27354 -9405
rect 27282 -9499 27354 -9451
rect 27282 -9545 27295 -9499
rect 27341 -9545 27354 -9499
rect 27282 -9593 27354 -9545
rect 27282 -9639 27295 -9593
rect 27341 -9639 27354 -9593
rect 27282 -9687 27354 -9639
rect 27282 -9733 27295 -9687
rect 27341 -9733 27354 -9687
rect 27282 -9781 27354 -9733
rect 27282 -9827 27295 -9781
rect 27341 -9827 27354 -9781
rect 27282 -9875 27354 -9827
rect 27282 -9921 27295 -9875
rect 27341 -9921 27354 -9875
rect 27282 -9969 27354 -9921
rect 27282 -10015 27295 -9969
rect 27341 -10015 27354 -9969
rect 27282 -10063 27354 -10015
rect 27282 -10109 27295 -10063
rect 27341 -10109 27354 -10063
rect 27282 -10157 27354 -10109
rect 27282 -10203 27295 -10157
rect 27341 -10203 27354 -10157
rect 27282 -10238 27354 -10203
rect 20984 -10251 27354 -10238
rect 20984 -10297 20997 -10251
rect 21043 -10297 21091 -10251
rect 21137 -10297 21185 -10251
rect 21231 -10297 21279 -10251
rect 21325 -10297 21373 -10251
rect 21419 -10297 21467 -10251
rect 21513 -10297 21561 -10251
rect 21607 -10297 21655 -10251
rect 21701 -10297 21749 -10251
rect 21795 -10297 21843 -10251
rect 21889 -10297 21937 -10251
rect 21983 -10297 22031 -10251
rect 22077 -10297 22125 -10251
rect 22171 -10297 22219 -10251
rect 22265 -10297 22313 -10251
rect 22359 -10297 22407 -10251
rect 22453 -10297 22501 -10251
rect 22547 -10297 22595 -10251
rect 22641 -10297 22689 -10251
rect 22735 -10297 22783 -10251
rect 22829 -10297 22877 -10251
rect 22923 -10297 22971 -10251
rect 23017 -10297 23065 -10251
rect 23111 -10297 23159 -10251
rect 23205 -10297 23253 -10251
rect 23299 -10297 23347 -10251
rect 23393 -10297 23441 -10251
rect 23487 -10297 23535 -10251
rect 23581 -10297 23629 -10251
rect 23675 -10297 23723 -10251
rect 23769 -10297 23817 -10251
rect 23863 -10297 23911 -10251
rect 23957 -10297 24005 -10251
rect 24051 -10297 24099 -10251
rect 24145 -10297 24193 -10251
rect 24239 -10297 24287 -10251
rect 24333 -10297 24381 -10251
rect 24427 -10297 24475 -10251
rect 24521 -10297 24569 -10251
rect 24615 -10297 24663 -10251
rect 24709 -10297 24757 -10251
rect 24803 -10297 24851 -10251
rect 24897 -10297 24945 -10251
rect 24991 -10297 25039 -10251
rect 25085 -10297 25133 -10251
rect 25179 -10297 25227 -10251
rect 25273 -10297 25321 -10251
rect 25367 -10297 25415 -10251
rect 25461 -10297 25509 -10251
rect 25555 -10297 25603 -10251
rect 25649 -10297 25697 -10251
rect 25743 -10297 25791 -10251
rect 25837 -10297 25885 -10251
rect 25931 -10297 25979 -10251
rect 26025 -10297 26073 -10251
rect 26119 -10297 26167 -10251
rect 26213 -10297 26261 -10251
rect 26307 -10297 26355 -10251
rect 26401 -10297 26449 -10251
rect 26495 -10297 26543 -10251
rect 26589 -10297 26637 -10251
rect 26683 -10297 26731 -10251
rect 26777 -10297 26825 -10251
rect 26871 -10297 26919 -10251
rect 26965 -10297 27013 -10251
rect 27059 -10297 27107 -10251
rect 27153 -10297 27201 -10251
rect 27247 -10297 27295 -10251
rect 27341 -10297 27354 -10251
rect 20984 -10310 27354 -10297
<< psubdiffcont >>
rect -10837 -4457 -10791 -4411
rect -10743 -4457 -10697 -4411
rect -10649 -4457 -10603 -4411
<< nsubdiffcont >>
rect -10783 -810 -10737 -764
rect -10689 -810 -10643 -764
rect -10784 -928 -10738 -882
rect -10690 -928 -10644 -882
rect 20997 -1743 21043 -1697
rect 21091 -1743 21137 -1697
rect 21185 -1743 21231 -1697
rect 21279 -1743 21325 -1697
rect 21373 -1743 21419 -1697
rect 21467 -1743 21513 -1697
rect 21561 -1743 21607 -1697
rect 21655 -1743 21701 -1697
rect 21749 -1743 21795 -1697
rect 21843 -1743 21889 -1697
rect 21937 -1743 21983 -1697
rect 22031 -1743 22077 -1697
rect 22125 -1743 22171 -1697
rect 22219 -1743 22265 -1697
rect 22313 -1743 22359 -1697
rect 22407 -1743 22453 -1697
rect 22501 -1743 22547 -1697
rect 22595 -1743 22641 -1697
rect 22689 -1743 22735 -1697
rect 22783 -1743 22829 -1697
rect 22877 -1743 22923 -1697
rect 22971 -1743 23017 -1697
rect 23065 -1743 23111 -1697
rect 23159 -1743 23205 -1697
rect 23253 -1743 23299 -1697
rect 23347 -1743 23393 -1697
rect 23441 -1743 23487 -1697
rect 23535 -1743 23581 -1697
rect 23629 -1743 23675 -1697
rect 23723 -1743 23769 -1697
rect 23817 -1743 23863 -1697
rect 23911 -1743 23957 -1697
rect 24005 -1743 24051 -1697
rect 24099 -1743 24145 -1697
rect 24193 -1743 24239 -1697
rect 24287 -1743 24333 -1697
rect 24381 -1743 24427 -1697
rect 24475 -1743 24521 -1697
rect 24569 -1743 24615 -1697
rect 24663 -1743 24709 -1697
rect 24757 -1743 24803 -1697
rect 24851 -1743 24897 -1697
rect 24945 -1743 24991 -1697
rect 25039 -1743 25085 -1697
rect 25133 -1743 25179 -1697
rect 25227 -1743 25273 -1697
rect 25321 -1743 25367 -1697
rect 25415 -1743 25461 -1697
rect 25509 -1743 25555 -1697
rect 25603 -1743 25649 -1697
rect 25697 -1743 25743 -1697
rect 25791 -1743 25837 -1697
rect 25885 -1743 25931 -1697
rect 25979 -1743 26025 -1697
rect 26073 -1743 26119 -1697
rect 26167 -1743 26213 -1697
rect 26261 -1743 26307 -1697
rect 26355 -1743 26401 -1697
rect 26449 -1743 26495 -1697
rect 26543 -1743 26589 -1697
rect 26637 -1743 26683 -1697
rect 26731 -1743 26777 -1697
rect 26825 -1743 26871 -1697
rect 26919 -1743 26965 -1697
rect 27013 -1743 27059 -1697
rect 27107 -1743 27153 -1697
rect 27201 -1743 27247 -1697
rect 27295 -1743 27341 -1697
rect 20997 -1837 21043 -1791
rect 20997 -1931 21043 -1885
rect 20997 -2025 21043 -1979
rect 20997 -2119 21043 -2073
rect 20997 -2213 21043 -2167
rect 20997 -2307 21043 -2261
rect 20997 -2401 21043 -2355
rect 20997 -2495 21043 -2449
rect 20997 -2589 21043 -2543
rect 20997 -2683 21043 -2637
rect 20997 -2777 21043 -2731
rect 20997 -2871 21043 -2825
rect 20997 -2965 21043 -2919
rect 20997 -3059 21043 -3013
rect 20997 -3153 21043 -3107
rect 2756 -3226 2802 -3180
rect 2850 -3226 2896 -3180
rect 2944 -3226 2990 -3180
rect 3038 -3226 3084 -3180
rect 3132 -3226 3178 -3180
rect 3226 -3226 3272 -3180
rect 3320 -3226 3366 -3180
rect 3414 -3226 3460 -3180
rect 3508 -3226 3554 -3180
rect 3602 -3226 3648 -3180
rect 3696 -3226 3742 -3180
rect 3790 -3226 3836 -3180
rect 3884 -3226 3930 -3180
rect 3978 -3226 4024 -3180
rect 4072 -3226 4118 -3180
rect 4166 -3226 4212 -3180
rect 4260 -3226 4306 -3180
rect 4354 -3226 4400 -3180
rect 4448 -3226 4494 -3180
rect 4542 -3226 4588 -3180
rect 4636 -3226 4682 -3180
rect 4730 -3226 4776 -3180
rect 4824 -3226 4870 -3180
rect 4918 -3226 4964 -3180
rect 5012 -3226 5058 -3180
rect 5106 -3226 5152 -3180
rect 5200 -3226 5246 -3180
rect 5294 -3226 5340 -3180
rect 5388 -3226 5434 -3180
rect 5482 -3226 5528 -3180
rect 5576 -3226 5622 -3180
rect 5670 -3226 5716 -3180
rect 5764 -3226 5810 -3180
rect 5858 -3226 5904 -3180
rect 5952 -3226 5998 -3180
rect 6046 -3226 6092 -3180
rect 6140 -3226 6186 -3180
rect 6234 -3226 6280 -3180
rect 6328 -3226 6374 -3180
rect 6422 -3226 6468 -3180
rect 6516 -3226 6562 -3180
rect 6610 -3226 6656 -3180
rect 6704 -3226 6750 -3180
rect 6798 -3226 6844 -3180
rect 6892 -3226 6938 -3180
rect 6986 -3226 7032 -3180
rect 7080 -3226 7126 -3180
rect 7174 -3226 7220 -3180
rect 7268 -3226 7314 -3180
rect 7362 -3226 7408 -3180
rect 7456 -3226 7502 -3180
rect 7550 -3226 7596 -3180
rect 7644 -3226 7690 -3180
rect 7738 -3226 7784 -3180
rect 7832 -3226 7878 -3180
rect 7926 -3226 7972 -3180
rect 8020 -3226 8066 -3180
rect 8114 -3226 8160 -3180
rect 8208 -3226 8254 -3180
rect 8302 -3226 8348 -3180
rect 8396 -3226 8442 -3180
rect 8490 -3226 8536 -3180
rect 8584 -3226 8630 -3180
rect 8678 -3226 8724 -3180
rect 8772 -3226 8818 -3180
rect 8866 -3226 8912 -3180
rect 8960 -3226 9006 -3180
rect 9054 -3226 9100 -3180
rect 2756 -3320 2802 -3274
rect 2756 -3414 2802 -3368
rect 2756 -3508 2802 -3462
rect 2756 -3602 2802 -3556
rect 2756 -3696 2802 -3650
rect 2756 -3790 2802 -3744
rect 2756 -3884 2802 -3838
rect 2756 -3978 2802 -3932
rect 2756 -4072 2802 -4026
rect 2756 -4166 2802 -4120
rect 2756 -4260 2802 -4214
rect 2756 -4354 2802 -4308
rect 2756 -4448 2802 -4402
rect 2756 -4542 2802 -4496
rect 2756 -4636 2802 -4590
rect 2756 -4730 2802 -4684
rect 2756 -4824 2802 -4778
rect 2756 -4918 2802 -4872
rect 2756 -5012 2802 -4966
rect 2756 -5106 2802 -5060
rect 2756 -5200 2802 -5154
rect 2756 -5294 2802 -5248
rect 2756 -5388 2802 -5342
rect 2756 -5482 2802 -5436
rect 2756 -5576 2802 -5530
rect 2756 -5670 2802 -5624
rect 2756 -5764 2802 -5718
rect 2756 -5858 2802 -5812
rect 2756 -5952 2802 -5906
rect 2756 -6046 2802 -6000
rect 2756 -6140 2802 -6094
rect 2756 -6234 2802 -6188
rect 2756 -6328 2802 -6282
rect 2756 -6422 2802 -6376
rect 2756 -6516 2802 -6470
rect 2756 -6610 2802 -6564
rect 2756 -6704 2802 -6658
rect 2756 -6798 2802 -6752
rect 2756 -6892 2802 -6846
rect 2756 -6986 2802 -6940
rect 2756 -7080 2802 -7034
rect 2756 -7174 2802 -7128
rect 2756 -7268 2802 -7222
rect 2756 -7362 2802 -7316
rect 2756 -7456 2802 -7410
rect 2756 -7550 2802 -7504
rect 2756 -7644 2802 -7598
rect 2756 -7738 2802 -7692
rect 2756 -7832 2802 -7786
rect 2756 -7926 2802 -7880
rect 2756 -8020 2802 -7974
rect 2756 -8114 2802 -8068
rect 2756 -8208 2802 -8162
rect 2756 -8302 2802 -8256
rect 2756 -8396 2802 -8350
rect 2756 -8490 2802 -8444
rect 2756 -8584 2802 -8538
rect 9054 -3320 9100 -3274
rect 9054 -3414 9100 -3368
rect 9054 -3508 9100 -3462
rect 9054 -3602 9100 -3556
rect 9054 -3696 9100 -3650
rect 9054 -3790 9100 -3744
rect 9054 -3884 9100 -3838
rect 9054 -3978 9100 -3932
rect 9054 -4072 9100 -4026
rect 9054 -4166 9100 -4120
rect 9054 -4260 9100 -4214
rect 9054 -4354 9100 -4308
rect 9054 -4448 9100 -4402
rect 9054 -4542 9100 -4496
rect 9054 -4636 9100 -4590
rect 9054 -4730 9100 -4684
rect 9054 -4824 9100 -4778
rect 9054 -4918 9100 -4872
rect 9054 -5012 9100 -4966
rect 9054 -5106 9100 -5060
rect 9054 -5200 9100 -5154
rect 9054 -5294 9100 -5248
rect 9054 -5388 9100 -5342
rect 9054 -5482 9100 -5436
rect 9054 -5576 9100 -5530
rect 9054 -5670 9100 -5624
rect 9054 -5764 9100 -5718
rect 9054 -5858 9100 -5812
rect 9054 -5952 9100 -5906
rect 9054 -6046 9100 -6000
rect 9054 -6140 9100 -6094
rect 9054 -6234 9100 -6188
rect 9054 -6328 9100 -6282
rect 9054 -6422 9100 -6376
rect 9054 -6516 9100 -6470
rect 9054 -6610 9100 -6564
rect 9054 -6704 9100 -6658
rect 9054 -6798 9100 -6752
rect 9054 -6892 9100 -6846
rect 9054 -6986 9100 -6940
rect 9054 -7080 9100 -7034
rect 9054 -7174 9100 -7128
rect 9054 -7268 9100 -7222
rect 9054 -7362 9100 -7316
rect 9054 -7456 9100 -7410
rect 9054 -7550 9100 -7504
rect 9054 -7644 9100 -7598
rect 9054 -7738 9100 -7692
rect 9054 -7832 9100 -7786
rect 9054 -7926 9100 -7880
rect 9054 -8020 9100 -7974
rect 9054 -8114 9100 -8068
rect 9054 -8208 9100 -8162
rect 9054 -8302 9100 -8256
rect 9054 -8396 9100 -8350
rect 9054 -8490 9100 -8444
rect 9054 -8584 9100 -8538
rect 2756 -8678 2802 -8632
rect 2850 -8678 2896 -8632
rect 2944 -8678 2990 -8632
rect 3038 -8678 3084 -8632
rect 3132 -8678 3178 -8632
rect 3226 -8678 3272 -8632
rect 3320 -8678 3366 -8632
rect 3414 -8678 3460 -8632
rect 3508 -8678 3554 -8632
rect 3602 -8678 3648 -8632
rect 3696 -8678 3742 -8632
rect 3790 -8678 3836 -8632
rect 3884 -8678 3930 -8632
rect 3978 -8678 4024 -8632
rect 4072 -8678 4118 -8632
rect 4166 -8678 4212 -8632
rect 4260 -8678 4306 -8632
rect 4354 -8678 4400 -8632
rect 4448 -8678 4494 -8632
rect 4542 -8678 4588 -8632
rect 4636 -8678 4682 -8632
rect 4730 -8678 4776 -8632
rect 4824 -8678 4870 -8632
rect 4918 -8678 4964 -8632
rect 5012 -8678 5058 -8632
rect 5106 -8678 5152 -8632
rect 5200 -8678 5246 -8632
rect 5294 -8678 5340 -8632
rect 5388 -8678 5434 -8632
rect 5482 -8678 5528 -8632
rect 5576 -8678 5622 -8632
rect 5670 -8678 5716 -8632
rect 5764 -8678 5810 -8632
rect 5858 -8678 5904 -8632
rect 5952 -8678 5998 -8632
rect 6046 -8678 6092 -8632
rect 6140 -8678 6186 -8632
rect 6234 -8678 6280 -8632
rect 6328 -8678 6374 -8632
rect 6422 -8678 6468 -8632
rect 6516 -8678 6562 -8632
rect 6610 -8678 6656 -8632
rect 6704 -8678 6750 -8632
rect 6798 -8678 6844 -8632
rect 6892 -8678 6938 -8632
rect 6986 -8678 7032 -8632
rect 7080 -8678 7126 -8632
rect 7174 -8678 7220 -8632
rect 7268 -8678 7314 -8632
rect 7362 -8678 7408 -8632
rect 7456 -8678 7502 -8632
rect 7550 -8678 7596 -8632
rect 7644 -8678 7690 -8632
rect 7738 -8678 7784 -8632
rect 7832 -8678 7878 -8632
rect 7926 -8678 7972 -8632
rect 8020 -8678 8066 -8632
rect 8114 -8678 8160 -8632
rect 8208 -8678 8254 -8632
rect 8302 -8678 8348 -8632
rect 8396 -8678 8442 -8632
rect 8490 -8678 8536 -8632
rect 8584 -8678 8630 -8632
rect 8678 -8678 8724 -8632
rect 8772 -8678 8818 -8632
rect 8866 -8678 8912 -8632
rect 8960 -8678 9006 -8632
rect 9054 -8678 9100 -8632
rect 20997 -3247 21043 -3201
rect 20997 -3341 21043 -3295
rect 20997 -3435 21043 -3389
rect 20997 -3529 21043 -3483
rect 20997 -3623 21043 -3577
rect 20997 -3717 21043 -3671
rect 20997 -3811 21043 -3765
rect 20997 -3905 21043 -3859
rect 20997 -3999 21043 -3953
rect 20997 -4093 21043 -4047
rect 20997 -4187 21043 -4141
rect 20997 -4281 21043 -4235
rect 20997 -4375 21043 -4329
rect 20997 -4469 21043 -4423
rect 20997 -4563 21043 -4517
rect 20997 -4657 21043 -4611
rect 20997 -4751 21043 -4705
rect 20997 -4845 21043 -4799
rect 20997 -4939 21043 -4893
rect 20997 -5033 21043 -4987
rect 20997 -5127 21043 -5081
rect 20997 -5221 21043 -5175
rect 20997 -5315 21043 -5269
rect 20997 -5409 21043 -5363
rect 20997 -5503 21043 -5457
rect 20997 -5597 21043 -5551
rect 20997 -5691 21043 -5645
rect 20997 -5785 21043 -5739
rect 20997 -5879 21043 -5833
rect 20997 -5973 21043 -5927
rect 20997 -6067 21043 -6021
rect 20997 -6161 21043 -6115
rect 20997 -6255 21043 -6209
rect 20997 -6349 21043 -6303
rect 20997 -6443 21043 -6397
rect 20997 -6537 21043 -6491
rect 20997 -6631 21043 -6585
rect 20997 -6725 21043 -6679
rect 20997 -6819 21043 -6773
rect 20997 -6913 21043 -6867
rect 20997 -7007 21043 -6961
rect 20997 -7101 21043 -7055
rect 20997 -7195 21043 -7149
rect 20997 -7289 21043 -7243
rect 20997 -7383 21043 -7337
rect 20997 -7477 21043 -7431
rect 20997 -7571 21043 -7525
rect 20997 -7665 21043 -7619
rect 20997 -7759 21043 -7713
rect 20997 -7853 21043 -7807
rect 20997 -7947 21043 -7901
rect 20997 -8041 21043 -7995
rect 20997 -8135 21043 -8089
rect 20997 -8229 21043 -8183
rect 20997 -8323 21043 -8277
rect 20997 -8417 21043 -8371
rect 20997 -8511 21043 -8465
rect 20997 -8605 21043 -8559
rect 20997 -8699 21043 -8653
rect 20997 -8793 21043 -8747
rect 20997 -8887 21043 -8841
rect 20997 -8981 21043 -8935
rect 20997 -9075 21043 -9029
rect 20997 -9169 21043 -9123
rect 20997 -9263 21043 -9217
rect 20997 -9357 21043 -9311
rect 20997 -9451 21043 -9405
rect 20997 -9545 21043 -9499
rect 20997 -9639 21043 -9593
rect 20997 -9733 21043 -9687
rect 20997 -9827 21043 -9781
rect 20997 -9921 21043 -9875
rect 20997 -10015 21043 -9969
rect 20997 -10109 21043 -10063
rect 20997 -10203 21043 -10157
rect 27295 -1837 27341 -1791
rect 27295 -1931 27341 -1885
rect 27295 -2025 27341 -1979
rect 27295 -2119 27341 -2073
rect 27295 -2213 27341 -2167
rect 27295 -2307 27341 -2261
rect 27295 -2401 27341 -2355
rect 27295 -2495 27341 -2449
rect 27295 -2589 27341 -2543
rect 27295 -2683 27341 -2637
rect 27295 -2777 27341 -2731
rect 27295 -2871 27341 -2825
rect 27295 -2965 27341 -2919
rect 27295 -3059 27341 -3013
rect 27295 -3153 27341 -3107
rect 27295 -3247 27341 -3201
rect 27295 -3341 27341 -3295
rect 27295 -3435 27341 -3389
rect 27295 -3529 27341 -3483
rect 27295 -3623 27341 -3577
rect 27295 -3717 27341 -3671
rect 27295 -3811 27341 -3765
rect 27295 -3905 27341 -3859
rect 27295 -3999 27341 -3953
rect 27295 -4093 27341 -4047
rect 27295 -4187 27341 -4141
rect 27295 -4281 27341 -4235
rect 27295 -4375 27341 -4329
rect 27295 -4469 27341 -4423
rect 27295 -4563 27341 -4517
rect 27295 -4657 27341 -4611
rect 27295 -4751 27341 -4705
rect 27295 -4845 27341 -4799
rect 27295 -4939 27341 -4893
rect 27295 -5033 27341 -4987
rect 27295 -5127 27341 -5081
rect 27295 -5221 27341 -5175
rect 27295 -5315 27341 -5269
rect 27295 -5409 27341 -5363
rect 27295 -5503 27341 -5457
rect 27295 -5597 27341 -5551
rect 27295 -5691 27341 -5645
rect 27295 -5785 27341 -5739
rect 27295 -5879 27341 -5833
rect 27295 -5973 27341 -5927
rect 27295 -6067 27341 -6021
rect 27295 -6161 27341 -6115
rect 27295 -6255 27341 -6209
rect 27295 -6349 27341 -6303
rect 27295 -6443 27341 -6397
rect 27295 -6537 27341 -6491
rect 27295 -6631 27341 -6585
rect 27295 -6725 27341 -6679
rect 27295 -6819 27341 -6773
rect 27295 -6913 27341 -6867
rect 27295 -7007 27341 -6961
rect 27295 -7101 27341 -7055
rect 27295 -7195 27341 -7149
rect 27295 -7289 27341 -7243
rect 27295 -7383 27341 -7337
rect 27295 -7477 27341 -7431
rect 27295 -7571 27341 -7525
rect 27295 -7665 27341 -7619
rect 27295 -7759 27341 -7713
rect 27295 -7853 27341 -7807
rect 27295 -7947 27341 -7901
rect 27295 -8041 27341 -7995
rect 27295 -8135 27341 -8089
rect 27295 -8229 27341 -8183
rect 27295 -8323 27341 -8277
rect 27295 -8417 27341 -8371
rect 27295 -8511 27341 -8465
rect 27295 -8605 27341 -8559
rect 27295 -8699 27341 -8653
rect 27295 -8793 27341 -8747
rect 27295 -8887 27341 -8841
rect 27295 -8981 27341 -8935
rect 27295 -9075 27341 -9029
rect 27295 -9169 27341 -9123
rect 27295 -9263 27341 -9217
rect 27295 -9357 27341 -9311
rect 27295 -9451 27341 -9405
rect 27295 -9545 27341 -9499
rect 27295 -9639 27341 -9593
rect 27295 -9733 27341 -9687
rect 27295 -9827 27341 -9781
rect 27295 -9921 27341 -9875
rect 27295 -10015 27341 -9969
rect 27295 -10109 27341 -10063
rect 27295 -10203 27341 -10157
rect 20997 -10297 21043 -10251
rect 21091 -10297 21137 -10251
rect 21185 -10297 21231 -10251
rect 21279 -10297 21325 -10251
rect 21373 -10297 21419 -10251
rect 21467 -10297 21513 -10251
rect 21561 -10297 21607 -10251
rect 21655 -10297 21701 -10251
rect 21749 -10297 21795 -10251
rect 21843 -10297 21889 -10251
rect 21937 -10297 21983 -10251
rect 22031 -10297 22077 -10251
rect 22125 -10297 22171 -10251
rect 22219 -10297 22265 -10251
rect 22313 -10297 22359 -10251
rect 22407 -10297 22453 -10251
rect 22501 -10297 22547 -10251
rect 22595 -10297 22641 -10251
rect 22689 -10297 22735 -10251
rect 22783 -10297 22829 -10251
rect 22877 -10297 22923 -10251
rect 22971 -10297 23017 -10251
rect 23065 -10297 23111 -10251
rect 23159 -10297 23205 -10251
rect 23253 -10297 23299 -10251
rect 23347 -10297 23393 -10251
rect 23441 -10297 23487 -10251
rect 23535 -10297 23581 -10251
rect 23629 -10297 23675 -10251
rect 23723 -10297 23769 -10251
rect 23817 -10297 23863 -10251
rect 23911 -10297 23957 -10251
rect 24005 -10297 24051 -10251
rect 24099 -10297 24145 -10251
rect 24193 -10297 24239 -10251
rect 24287 -10297 24333 -10251
rect 24381 -10297 24427 -10251
rect 24475 -10297 24521 -10251
rect 24569 -10297 24615 -10251
rect 24663 -10297 24709 -10251
rect 24757 -10297 24803 -10251
rect 24851 -10297 24897 -10251
rect 24945 -10297 24991 -10251
rect 25039 -10297 25085 -10251
rect 25133 -10297 25179 -10251
rect 25227 -10297 25273 -10251
rect 25321 -10297 25367 -10251
rect 25415 -10297 25461 -10251
rect 25509 -10297 25555 -10251
rect 25603 -10297 25649 -10251
rect 25697 -10297 25743 -10251
rect 25791 -10297 25837 -10251
rect 25885 -10297 25931 -10251
rect 25979 -10297 26025 -10251
rect 26073 -10297 26119 -10251
rect 26167 -10297 26213 -10251
rect 26261 -10297 26307 -10251
rect 26355 -10297 26401 -10251
rect 26449 -10297 26495 -10251
rect 26543 -10297 26589 -10251
rect 26637 -10297 26683 -10251
rect 26731 -10297 26777 -10251
rect 26825 -10297 26871 -10251
rect 26919 -10297 26965 -10251
rect 27013 -10297 27059 -10251
rect 27107 -10297 27153 -10251
rect 27201 -10297 27247 -10251
rect 27295 -10297 27341 -10251
<< polysilicon >>
rect -10736 -3030 -10680 -1336
rect -10909 -3045 -10680 -3030
rect -10909 -3093 -10894 -3045
rect -10830 -3093 -10680 -3045
rect -10909 -3106 -10680 -3093
rect -10736 -4194 -10680 -3106
<< polycontact >>
rect -10894 -3093 -10830 -3045
<< metal1 >>
rect 1270 14910 3980 15300
rect 1270 14800 5640 14910
rect 1270 14730 1770 14800
rect -16811 14442 1770 14730
rect -19056 14230 1770 14442
rect 3480 14410 5640 14800
rect -19056 14016 -16348 14230
rect -13843 14222 -12031 14230
rect -13872 11981 -13718 11998
rect -13872 11916 -13829 11981
rect -13765 11916 -13718 11981
rect -13872 11903 -13718 11916
rect -9952 11997 -9728 12025
rect -9952 11937 -9917 11997
rect -9857 11996 -9728 11997
rect -9857 11937 -9804 11996
rect -9952 11936 -9804 11937
rect -9744 11936 -9728 11996
rect -9952 11908 -9728 11936
rect -7207 12023 -7082 12024
rect -7207 12001 -6972 12023
rect -7207 11941 -7165 12001
rect -7105 11941 -7051 12001
rect -6991 11941 -6972 12001
rect -7207 11918 -6972 11941
rect 1270 10850 1770 14230
rect -13342 10002 -5484 10495
rect -13342 6759 -12849 10002
rect -13342 6678 -12501 6759
rect -13342 6625 -12170 6678
rect -13342 6623 -12850 6625
rect -13342 6571 -13264 6623
rect -13212 6571 -13160 6623
rect -13108 6571 -13056 6623
rect -13004 6573 -12850 6623
rect -12798 6573 -12746 6625
rect -12694 6573 -12642 6625
rect -12590 6618 -12170 6625
rect -12590 6573 -12487 6618
rect -13004 6571 -12487 6573
rect -13342 6566 -12487 6571
rect -12435 6566 -12383 6618
rect -12331 6566 -12279 6618
rect -12227 6566 -12170 6618
rect -13342 6521 -12170 6566
rect -13342 6519 -12850 6521
rect -13342 6467 -13264 6519
rect -13212 6467 -13160 6519
rect -13108 6467 -13056 6519
rect -13004 6469 -12850 6519
rect -12798 6469 -12746 6521
rect -12694 6469 -12642 6521
rect -12590 6514 -12170 6521
rect -12590 6469 -12487 6514
rect -13004 6467 -12487 6469
rect -13342 6462 -12487 6467
rect -12435 6462 -12383 6514
rect -12331 6462 -12279 6514
rect -12227 6462 -12170 6514
rect -13342 6417 -12170 6462
rect -13342 6415 -12850 6417
rect -13342 6363 -13264 6415
rect -13212 6363 -13160 6415
rect -13108 6363 -13056 6415
rect -13004 6365 -12850 6415
rect -12798 6365 -12746 6417
rect -12694 6365 -12642 6417
rect -12590 6410 -12170 6417
rect -12590 6365 -12487 6410
rect -13004 6363 -12487 6365
rect -13342 6358 -12487 6363
rect -12435 6358 -12383 6410
rect -12331 6358 -12279 6410
rect -12227 6358 -12170 6410
rect -13342 6207 -12170 6358
rect -13342 6155 -13262 6207
rect -13210 6155 -13158 6207
rect -13106 6155 -13054 6207
rect -13002 6190 -12170 6207
rect -13002 6155 -12820 6190
rect -13342 6138 -12820 6155
rect -12768 6138 -12716 6190
rect -12664 6138 -12612 6190
rect -12560 6183 -12170 6190
rect -12560 6138 -12457 6183
rect -13342 6131 -12457 6138
rect -12405 6131 -12353 6183
rect -12301 6131 -12249 6183
rect -12197 6131 -12170 6183
rect -13342 6103 -12170 6131
rect -13342 6051 -13262 6103
rect -13210 6051 -13158 6103
rect -13106 6051 -13054 6103
rect -13002 6086 -12170 6103
rect -13002 6051 -12820 6086
rect -13342 6034 -12820 6051
rect -12768 6034 -12716 6086
rect -12664 6034 -12612 6086
rect -12560 6079 -12170 6086
rect -12560 6034 -12457 6079
rect -13342 6027 -12457 6034
rect -12405 6027 -12353 6079
rect -12301 6027 -12249 6079
rect -12197 6027 -12170 6079
rect -13342 5999 -12170 6027
rect -13342 5947 -13262 5999
rect -13210 5947 -13158 5999
rect -13106 5947 -13054 5999
rect -13002 5982 -12170 5999
rect -13002 5947 -12820 5982
rect -13342 5930 -12820 5947
rect -12768 5930 -12716 5982
rect -12664 5930 -12612 5982
rect -12560 5975 -12170 5982
rect -12560 5930 -12457 5975
rect -13342 5923 -12457 5930
rect -12405 5923 -12353 5975
rect -12301 5923 -12249 5975
rect -12197 5923 -12170 5975
rect -13342 5855 -12170 5923
rect -13342 5800 -12501 5855
rect -13342 5766 -12849 5800
rect -13342 5714 -13262 5766
rect -13210 5714 -13158 5766
rect -13106 5714 -13054 5766
rect -13002 5714 -12849 5766
rect -13342 5662 -12849 5714
rect -13342 5610 -13262 5662
rect -13210 5610 -13158 5662
rect -13106 5610 -13054 5662
rect -13002 5610 -12849 5662
rect -13342 5558 -12849 5610
rect -13342 5506 -13262 5558
rect -13210 5506 -13158 5558
rect -13106 5506 -13054 5558
rect -13002 5506 -12849 5558
rect -13342 2376 -12849 5506
rect -18329 2337 -12849 2376
rect -21120 1921 -12849 2337
rect -18329 1883 -12849 1921
rect 361 -245 879 4609
rect 1981 -245 2499 1479
rect 3753 -245 4174 1477
rect 14007 216 14672 1303
rect 13977 215 14672 216
rect 13977 204 14387 215
rect 13977 152 13989 204
rect 14041 152 14093 204
rect 14145 152 14197 204
rect 14249 163 14387 204
rect 14439 163 14491 215
rect 14543 163 14595 215
rect 14647 163 14672 215
rect 14249 152 14672 163
rect 13977 111 14672 152
rect 13977 100 14387 111
rect 13977 48 13989 100
rect 14041 48 14093 100
rect 14145 48 14197 100
rect 14249 59 14387 100
rect 14439 59 14491 111
rect 14543 59 14595 111
rect 14647 59 14672 111
rect 14249 48 14672 59
rect 13977 7 14672 48
rect 13977 -4 14387 7
rect 13977 -56 13989 -4
rect 14041 -56 14093 -4
rect 14145 -56 14197 -4
rect 14249 -45 14387 -4
rect 14439 -45 14491 7
rect 14543 -45 14595 7
rect 14647 -45 14672 7
rect 14249 -56 14672 -45
rect 13977 -68 14672 -56
rect 14007 -106 14672 -68
rect -17089 -533 4174 -245
rect -19334 -745 4174 -533
rect -19334 -959 -16626 -745
rect -14121 -753 -12309 -745
rect -10873 -764 -10531 -745
rect -6309 -763 4174 -745
rect -10873 -810 -10783 -764
rect -10737 -810 -10689 -764
rect -10643 -810 -10531 -764
rect -10873 -852 -10531 -810
rect -10955 -882 -10445 -852
rect -10955 -928 -10784 -882
rect -10738 -928 -10690 -882
rect -10644 -928 -10445 -882
rect -10955 -965 -10445 -928
rect -10819 -2934 -10757 -965
rect -14173 -2993 -13989 -2968
rect -14173 -3049 -14136 -2993
rect -14072 -3049 -13989 -2993
rect -14173 -3070 -13989 -3049
rect -10971 -3043 -10816 -3027
rect -10971 -3099 -10942 -3043
rect -10878 -3045 -10816 -3043
rect -10830 -3093 -10816 -3045
rect -10878 -3099 -10816 -3093
rect -10971 -3111 -10816 -3099
rect -10661 -3032 -10591 -1131
rect 3753 -1723 4174 -763
rect 20566 -1298 20987 1018
rect 23003 -1298 23424 1054
rect 20566 -1670 23424 -1298
rect 20566 -1697 27368 -1670
rect 20566 -1723 20997 -1697
rect 3753 -1743 20997 -1723
rect 21043 -1743 21091 -1697
rect 21137 -1743 21185 -1697
rect 21231 -1743 21279 -1697
rect 21325 -1743 21373 -1697
rect 21419 -1743 21467 -1697
rect 21513 -1743 21561 -1697
rect 21607 -1743 21655 -1697
rect 21701 -1743 21749 -1697
rect 21795 -1743 21843 -1697
rect 21889 -1743 21937 -1697
rect 21983 -1743 22031 -1697
rect 22077 -1743 22125 -1697
rect 22171 -1743 22219 -1697
rect 22265 -1743 22313 -1697
rect 22359 -1743 22407 -1697
rect 22453 -1743 22501 -1697
rect 22547 -1743 22595 -1697
rect 22641 -1743 22689 -1697
rect 22735 -1743 22783 -1697
rect 22829 -1743 22877 -1697
rect 22923 -1743 22971 -1697
rect 23017 -1743 23065 -1697
rect 23111 -1743 23159 -1697
rect 23205 -1743 23253 -1697
rect 23299 -1743 23347 -1697
rect 23393 -1743 23441 -1697
rect 23487 -1743 23535 -1697
rect 23581 -1743 23629 -1697
rect 23675 -1743 23723 -1697
rect 23769 -1743 23817 -1697
rect 23863 -1743 23911 -1697
rect 23957 -1743 24005 -1697
rect 24051 -1743 24099 -1697
rect 24145 -1743 24193 -1697
rect 24239 -1743 24287 -1697
rect 24333 -1743 24381 -1697
rect 24427 -1743 24475 -1697
rect 24521 -1743 24569 -1697
rect 24615 -1743 24663 -1697
rect 24709 -1743 24757 -1697
rect 24803 -1743 24851 -1697
rect 24897 -1743 24945 -1697
rect 24991 -1743 25039 -1697
rect 25085 -1743 25133 -1697
rect 25179 -1743 25227 -1697
rect 25273 -1743 25321 -1697
rect 25367 -1743 25415 -1697
rect 25461 -1743 25509 -1697
rect 25555 -1743 25603 -1697
rect 25649 -1743 25697 -1697
rect 25743 -1743 25791 -1697
rect 25837 -1743 25885 -1697
rect 25931 -1743 25979 -1697
rect 26025 -1743 26073 -1697
rect 26119 -1743 26167 -1697
rect 26213 -1743 26261 -1697
rect 26307 -1743 26355 -1697
rect 26401 -1743 26449 -1697
rect 26495 -1743 26543 -1697
rect 26589 -1743 26637 -1697
rect 26683 -1743 26731 -1697
rect 26777 -1743 26825 -1697
rect 26871 -1743 26919 -1697
rect 26965 -1743 27013 -1697
rect 27059 -1743 27107 -1697
rect 27153 -1743 27201 -1697
rect 27247 -1743 27295 -1697
rect 27341 -1743 27368 -1697
rect 3753 -1770 27368 -1743
rect 3753 -1791 21070 -1770
rect 3753 -1837 20997 -1791
rect 21043 -1837 21070 -1791
rect 3753 -1885 21070 -1837
rect 27268 -1791 27368 -1770
rect 27268 -1837 27295 -1791
rect 27341 -1837 27368 -1791
rect 3753 -1931 20997 -1885
rect 21043 -1931 21070 -1885
rect 3753 -1979 21070 -1931
rect 25788 -1869 25968 -1857
rect 25788 -1921 25800 -1869
rect 25852 -1921 25904 -1869
rect 25956 -1921 25968 -1869
rect 25788 -1949 25968 -1921
rect 26277 -1870 26457 -1858
rect 26277 -1922 26289 -1870
rect 26341 -1922 26393 -1870
rect 26445 -1922 26457 -1870
rect 26277 -1946 26457 -1922
rect 27268 -1885 27368 -1837
rect 27268 -1931 27295 -1885
rect 27341 -1931 27368 -1885
rect 3753 -2025 20997 -1979
rect 21043 -2025 21070 -1979
rect 3753 -2073 21070 -2025
rect 3753 -2119 20997 -2073
rect 21043 -2119 21070 -2073
rect 3753 -2144 21070 -2119
rect 3753 -2724 4174 -2144
rect 20566 -2167 21070 -2144
rect 20566 -2213 20997 -2167
rect 21043 -2213 21070 -2167
rect 20566 -2244 21070 -2213
rect 21926 -2173 23106 -1962
rect 20566 -2261 21504 -2244
rect 20566 -2307 20997 -2261
rect 21043 -2307 21504 -2261
rect 20566 -2355 21504 -2307
rect 21926 -2349 22137 -2173
rect 20566 -2401 20997 -2355
rect 21043 -2367 21504 -2355
rect 21043 -2401 21070 -2367
rect 20566 -2449 21070 -2401
rect 20566 -2495 20997 -2449
rect 21043 -2495 21070 -2449
rect 20566 -2543 21070 -2495
rect 20566 -2589 20997 -2543
rect 21043 -2589 21070 -2543
rect 20566 -2637 21070 -2589
rect 20566 -2683 20997 -2637
rect 21043 -2683 21070 -2637
rect 22407 -2451 22618 -2275
rect 22895 -2349 23106 -2173
rect 23862 -2173 25042 -1962
rect 23376 -2451 23587 -2275
rect 23862 -2349 24073 -2173
rect 22407 -2662 23587 -2451
rect 24319 -2455 24530 -2275
rect 24831 -2349 25042 -2173
rect 25779 -1973 25990 -1949
rect 25779 -2025 25800 -1973
rect 25852 -2025 25904 -1973
rect 25956 -2025 25990 -1973
rect 25779 -2077 25990 -2025
rect 25779 -2129 25800 -2077
rect 25852 -2129 25904 -2077
rect 25956 -2129 25990 -2077
rect 25288 -2455 25499 -2275
rect 25779 -2336 25990 -2129
rect 26261 -1974 26472 -1946
rect 26261 -2026 26289 -1974
rect 26341 -2026 26393 -1974
rect 26445 -2026 26472 -1974
rect 26261 -2078 26472 -2026
rect 26261 -2130 26289 -2078
rect 26341 -2130 26393 -2078
rect 26445 -2130 26472 -2078
rect 26261 -2333 26472 -2130
rect 27268 -1979 27368 -1931
rect 27268 -2025 27295 -1979
rect 27341 -2025 27368 -1979
rect 27268 -2073 27368 -2025
rect 27268 -2119 27295 -2073
rect 27341 -2119 27368 -2073
rect 27268 -2167 27368 -2119
rect 27268 -2213 27295 -2167
rect 27341 -2213 27368 -2167
rect 27268 -2244 27368 -2213
rect 26820 -2261 27368 -2244
rect 26820 -2307 27295 -2261
rect 27341 -2307 27368 -2261
rect 26820 -2355 27368 -2307
rect 26820 -2367 27295 -2355
rect 24319 -2666 25499 -2455
rect 27268 -2401 27295 -2367
rect 27341 -2401 27368 -2355
rect 27268 -2449 27368 -2401
rect 27268 -2495 27295 -2449
rect 27341 -2495 27368 -2449
rect 27268 -2543 27368 -2495
rect 27268 -2589 27295 -2543
rect 27341 -2589 27368 -2543
rect 27268 -2637 27368 -2589
rect 20566 -2724 21070 -2683
rect 3753 -2731 21070 -2724
rect 3753 -2777 20997 -2731
rect 21043 -2777 21070 -2731
rect 3753 -2825 21070 -2777
rect 3753 -2871 20997 -2825
rect 21043 -2871 21070 -2825
rect 3753 -2919 21070 -2871
rect -10149 -2975 -9974 -2954
rect -10149 -2981 -10128 -2975
rect -10305 -3032 -10128 -2981
rect -10661 -3045 -10128 -3032
rect -10050 -3045 -9974 -2975
rect -10661 -3051 -9974 -3045
rect -10661 -3102 -10235 -3051
rect -10149 -3065 -9974 -3051
rect -7416 -2976 -7241 -2951
rect -7416 -3046 -7377 -2976
rect -7299 -3046 -7241 -2976
rect -7416 -3062 -7241 -3046
rect 3753 -2965 20997 -2919
rect 21043 -2965 21070 -2919
rect 3753 -3013 21070 -2965
rect 3753 -3059 20997 -3013
rect 21043 -3059 21070 -3013
rect -10821 -4345 -10759 -3162
rect -10661 -4198 -10591 -3102
rect 3753 -3107 21070 -3059
rect 3753 -3145 20997 -3107
rect 3753 -3153 9127 -3145
rect 2729 -3180 9127 -3153
rect 2729 -3226 2756 -3180
rect 2802 -3226 2850 -3180
rect 2896 -3226 2944 -3180
rect 2990 -3226 3038 -3180
rect 3084 -3226 3132 -3180
rect 3178 -3226 3226 -3180
rect 3272 -3226 3320 -3180
rect 3366 -3226 3414 -3180
rect 3460 -3226 3508 -3180
rect 3554 -3226 3602 -3180
rect 3648 -3226 3696 -3180
rect 3742 -3226 3790 -3180
rect 3836 -3226 3884 -3180
rect 3930 -3226 3978 -3180
rect 4024 -3226 4072 -3180
rect 4118 -3226 4166 -3180
rect 4212 -3226 4260 -3180
rect 4306 -3226 4354 -3180
rect 4400 -3226 4448 -3180
rect 4494 -3226 4542 -3180
rect 4588 -3226 4636 -3180
rect 4682 -3226 4730 -3180
rect 4776 -3226 4824 -3180
rect 4870 -3226 4918 -3180
rect 4964 -3226 5012 -3180
rect 5058 -3226 5106 -3180
rect 5152 -3226 5200 -3180
rect 5246 -3226 5294 -3180
rect 5340 -3226 5388 -3180
rect 5434 -3226 5482 -3180
rect 5528 -3226 5576 -3180
rect 5622 -3226 5670 -3180
rect 5716 -3226 5764 -3180
rect 5810 -3226 5858 -3180
rect 5904 -3226 5952 -3180
rect 5998 -3226 6046 -3180
rect 6092 -3226 6140 -3180
rect 6186 -3226 6234 -3180
rect 6280 -3226 6328 -3180
rect 6374 -3226 6422 -3180
rect 6468 -3226 6516 -3180
rect 6562 -3226 6610 -3180
rect 6656 -3226 6704 -3180
rect 6750 -3226 6798 -3180
rect 6844 -3226 6892 -3180
rect 6938 -3226 6986 -3180
rect 7032 -3226 7080 -3180
rect 7126 -3226 7174 -3180
rect 7220 -3226 7268 -3180
rect 7314 -3226 7362 -3180
rect 7408 -3226 7456 -3180
rect 7502 -3226 7550 -3180
rect 7596 -3226 7644 -3180
rect 7690 -3226 7738 -3180
rect 7784 -3226 7832 -3180
rect 7878 -3226 7926 -3180
rect 7972 -3226 8020 -3180
rect 8066 -3226 8114 -3180
rect 8160 -3226 8208 -3180
rect 8254 -3226 8302 -3180
rect 8348 -3226 8396 -3180
rect 8442 -3226 8490 -3180
rect 8536 -3226 8584 -3180
rect 8630 -3226 8678 -3180
rect 8724 -3226 8772 -3180
rect 8818 -3226 8866 -3180
rect 8912 -3226 8960 -3180
rect 9006 -3226 9054 -3180
rect 9100 -3226 9127 -3180
rect 2729 -3253 9127 -3226
rect 2729 -3274 2829 -3253
rect 2729 -3320 2756 -3274
rect 2802 -3320 2829 -3274
rect 2729 -3368 2829 -3320
rect 9027 -3274 9127 -3253
rect 9027 -3320 9054 -3274
rect 9100 -3320 9127 -3274
rect 2729 -3414 2756 -3368
rect 2802 -3414 2829 -3368
rect 7519 -3363 7699 -3351
rect 2729 -3462 2829 -3414
rect 2729 -3508 2756 -3462
rect 2802 -3508 2829 -3462
rect 2729 -3556 2829 -3508
rect 2729 -3602 2756 -3556
rect 2802 -3602 2829 -3556
rect 2729 -3650 2829 -3602
rect 2729 -3696 2756 -3650
rect 2802 -3669 2829 -3650
rect 3656 -3603 4836 -3392
rect 2802 -3696 3229 -3669
rect 2729 -3744 3229 -3696
rect 2729 -3790 2756 -3744
rect 2802 -3790 3229 -3744
rect 3656 -3779 3867 -3603
rect 2729 -3792 3229 -3790
rect 2729 -3838 2829 -3792
rect 2729 -3884 2756 -3838
rect 2802 -3884 2829 -3838
rect 2729 -3932 2829 -3884
rect 2729 -3978 2756 -3932
rect 2802 -3978 2829 -3932
rect 2729 -4026 2829 -3978
rect 2729 -4072 2756 -4026
rect 2802 -4072 2829 -4026
rect 2729 -4120 2829 -4072
rect 4137 -3881 4348 -3705
rect 4625 -3779 4836 -3603
rect 5592 -3603 6772 -3392
rect 7519 -3415 7531 -3363
rect 7583 -3415 7635 -3363
rect 7687 -3415 7699 -3363
rect 7519 -3467 7699 -3415
rect 7519 -3519 7531 -3467
rect 7583 -3519 7635 -3467
rect 7687 -3519 7699 -3467
rect 7519 -3554 7699 -3519
rect 8006 -3359 8186 -3347
rect 8006 -3411 8018 -3359
rect 8070 -3411 8122 -3359
rect 8174 -3411 8186 -3359
rect 8006 -3463 8186 -3411
rect 8006 -3515 8018 -3463
rect 8070 -3515 8122 -3463
rect 8174 -3515 8186 -3463
rect 8006 -3554 8186 -3515
rect 9027 -3368 9127 -3320
rect 9027 -3414 9054 -3368
rect 9100 -3414 9127 -3368
rect 9027 -3462 9127 -3414
rect 9027 -3508 9054 -3462
rect 9100 -3508 9127 -3462
rect 5106 -3881 5317 -3705
rect 5592 -3779 5803 -3603
rect 4137 -4092 5317 -3881
rect 6049 -3885 6260 -3705
rect 6561 -3779 6772 -3603
rect 7509 -3571 7720 -3554
rect 7509 -3623 7531 -3571
rect 7583 -3623 7635 -3571
rect 7687 -3623 7720 -3571
rect 7018 -3885 7229 -3705
rect 7509 -3766 7720 -3623
rect 7991 -3567 8202 -3554
rect 7991 -3619 8018 -3567
rect 8070 -3619 8122 -3567
rect 8174 -3619 8202 -3567
rect 7991 -3763 8202 -3619
rect 9027 -3556 9127 -3508
rect 9027 -3602 9054 -3556
rect 9100 -3602 9127 -3556
rect 9027 -3650 9127 -3602
rect 9027 -3675 9054 -3650
rect 8596 -3696 9054 -3675
rect 9100 -3696 9127 -3650
rect 8596 -3744 9127 -3696
rect 8596 -3790 9054 -3744
rect 9100 -3790 9127 -3744
rect 8596 -3798 9127 -3790
rect 6049 -4096 7229 -3885
rect 9027 -3838 9127 -3798
rect 9027 -3884 9054 -3838
rect 9100 -3884 9127 -3838
rect 9027 -3932 9127 -3884
rect 9027 -3978 9054 -3932
rect 9100 -3978 9127 -3932
rect 9027 -4026 9127 -3978
rect 9027 -4072 9054 -4026
rect 9100 -4072 9127 -4026
rect 2729 -4166 2756 -4120
rect 2802 -4166 2829 -4120
rect 2729 -4214 2829 -4166
rect 2729 -4260 2756 -4214
rect 2802 -4260 2829 -4214
rect 2729 -4308 2829 -4260
rect -10940 -4411 -10462 -4345
rect -10940 -4457 -10837 -4411
rect -10791 -4457 -10743 -4411
rect -10697 -4457 -10649 -4411
rect -10603 -4457 -10462 -4411
rect -10940 -4480 -10462 -4457
rect 2729 -4354 2756 -4308
rect 2802 -4354 2829 -4308
rect 2729 -4402 2829 -4354
rect 2729 -4448 2756 -4402
rect 2802 -4448 2829 -4402
rect -13620 -4973 -5762 -4480
rect 2729 -4496 2829 -4448
rect 2729 -4542 2756 -4496
rect 2802 -4542 2829 -4496
rect 2729 -4590 2829 -4542
rect 2729 -4636 2756 -4590
rect 2802 -4636 2829 -4590
rect 2729 -4684 2829 -4636
rect 2729 -4730 2756 -4684
rect 2802 -4730 2829 -4684
rect 2729 -4778 2829 -4730
rect 2729 -4824 2756 -4778
rect 2802 -4824 2829 -4778
rect 2729 -4872 2829 -4824
rect 2729 -4918 2756 -4872
rect 2802 -4918 2829 -4872
rect 2729 -4966 2829 -4918
rect -13620 -9409 -13127 -4973
rect 2729 -5012 2756 -4966
rect 2802 -5012 2829 -4966
rect 2729 -5060 2829 -5012
rect 2729 -5106 2756 -5060
rect 2802 -5106 2829 -5060
rect 2729 -5154 2829 -5106
rect 9027 -4120 9127 -4072
rect 9027 -4166 9054 -4120
rect 9100 -4166 9127 -4120
rect 9027 -4214 9127 -4166
rect 9027 -4260 9054 -4214
rect 9100 -4260 9127 -4214
rect 9027 -4308 9127 -4260
rect 10543 -4293 10964 -3145
rect 13154 -4277 13575 -3145
rect 14555 -3476 14977 -3467
rect 14073 -3517 14977 -3476
rect 14073 -3522 14462 -3517
rect 14073 -3574 14130 -3522
rect 14182 -3574 14234 -3522
rect 14286 -3574 14338 -3522
rect 14390 -3569 14462 -3522
rect 14514 -3569 14566 -3517
rect 14618 -3569 14670 -3517
rect 14722 -3569 14977 -3517
rect 14390 -3574 14977 -3569
rect 14073 -3621 14977 -3574
rect 14073 -3626 14462 -3621
rect 14073 -3678 14130 -3626
rect 14182 -3678 14234 -3626
rect 14286 -3678 14338 -3626
rect 14390 -3673 14462 -3626
rect 14514 -3673 14566 -3621
rect 14618 -3673 14670 -3621
rect 14722 -3673 14977 -3621
rect 14390 -3678 14977 -3673
rect 14073 -3725 14977 -3678
rect 14073 -3730 14462 -3725
rect 14073 -3782 14130 -3730
rect 14182 -3782 14234 -3730
rect 14286 -3782 14338 -3730
rect 14390 -3777 14462 -3730
rect 14514 -3777 14566 -3725
rect 14618 -3777 14670 -3725
rect 14722 -3777 14977 -3725
rect 14390 -3782 14977 -3777
rect 14073 -3857 14977 -3782
rect 14372 -3866 14977 -3857
rect 14372 -3918 14464 -3866
rect 14516 -3918 14568 -3866
rect 14620 -3918 14672 -3866
rect 14724 -3918 14977 -3866
rect 14372 -3970 14977 -3918
rect 14372 -4022 14464 -3970
rect 14516 -4022 14568 -3970
rect 14620 -4022 14672 -3970
rect 14724 -4022 14977 -3970
rect 14372 -4074 14977 -4022
rect 14372 -4126 14464 -4074
rect 14516 -4126 14568 -4074
rect 14620 -4126 14672 -4074
rect 14724 -4126 14977 -4074
rect 9027 -4354 9054 -4308
rect 9100 -4354 9127 -4308
rect 9027 -4402 9127 -4354
rect 9027 -4448 9054 -4402
rect 9100 -4448 9127 -4402
rect 9027 -4496 9127 -4448
rect 9027 -4542 9054 -4496
rect 9100 -4542 9127 -4496
rect 9027 -4590 9127 -4542
rect 9027 -4636 9054 -4590
rect 9100 -4636 9127 -4590
rect 9027 -4684 9127 -4636
rect 9027 -4730 9054 -4684
rect 9100 -4730 9127 -4684
rect 9027 -4778 9127 -4730
rect 9027 -4824 9054 -4778
rect 9100 -4824 9127 -4778
rect 9027 -4872 9127 -4824
rect 9027 -4918 9054 -4872
rect 9100 -4918 9127 -4872
rect 9027 -4966 9127 -4918
rect 9027 -5012 9054 -4966
rect 9100 -5012 9127 -4966
rect 9027 -5060 9127 -5012
rect 9027 -5106 9054 -5060
rect 9100 -5106 9127 -5060
rect 2729 -5200 2756 -5154
rect 2802 -5200 2829 -5154
rect 2729 -5248 2829 -5200
rect 2729 -5294 2756 -5248
rect 2802 -5294 2829 -5248
rect 2729 -5342 2829 -5294
rect 2729 -5388 2756 -5342
rect 2802 -5388 2829 -5342
rect 2729 -5421 2829 -5388
rect 4622 -5325 5802 -5114
rect 2729 -5436 3248 -5421
rect 2729 -5482 2756 -5436
rect 2802 -5482 3248 -5436
rect 2729 -5530 3248 -5482
rect 2729 -5576 2756 -5530
rect 2802 -5544 3248 -5530
rect 2802 -5576 2829 -5544
rect 2729 -5624 2829 -5576
rect 2729 -5670 2756 -5624
rect 2802 -5670 2829 -5624
rect 2729 -5718 2829 -5670
rect 2729 -5764 2756 -5718
rect 2802 -5764 2829 -5718
rect 2729 -5812 2829 -5764
rect 2729 -5858 2756 -5812
rect 2802 -5858 2829 -5812
rect 2729 -5906 2829 -5858
rect 2729 -5952 2756 -5906
rect 2802 -5952 2829 -5906
rect 2729 -6000 2829 -5952
rect 2729 -6046 2756 -6000
rect 2802 -6046 2829 -6000
rect 2729 -6094 2829 -6046
rect 2729 -6140 2756 -6094
rect 2802 -6140 2829 -6094
rect 2729 -6188 2829 -6140
rect 2729 -6234 2756 -6188
rect 2802 -6220 2829 -6188
rect 2802 -6234 3229 -6220
rect 2729 -6282 3229 -6234
rect 2729 -6328 2756 -6282
rect 2802 -6328 3229 -6282
rect 3655 -6317 3866 -5441
rect 4148 -6317 4359 -5441
rect 4622 -5501 4833 -5325
rect 5103 -5603 5314 -5427
rect 5591 -5501 5802 -5325
rect 6542 -5334 7722 -5123
rect 6072 -5603 6283 -5427
rect 6542 -5510 6753 -5334
rect 5103 -5814 6283 -5603
rect 7015 -5607 7226 -5427
rect 7511 -5510 7722 -5334
rect 9027 -5154 9127 -5106
rect 9027 -5200 9054 -5154
rect 9100 -5200 9127 -5154
rect 9027 -5248 9127 -5200
rect 9027 -5294 9054 -5248
rect 9100 -5294 9127 -5248
rect 9027 -5342 9127 -5294
rect 9027 -5388 9054 -5342
rect 9100 -5388 9127 -5342
rect 9027 -5421 9127 -5388
rect 7984 -5607 8195 -5427
rect 8586 -5436 9127 -5421
rect 8586 -5482 9054 -5436
rect 9100 -5482 9127 -5436
rect 8586 -5530 9127 -5482
rect 8586 -5544 9054 -5530
rect 7015 -5818 8195 -5607
rect 9027 -5576 9054 -5544
rect 9100 -5576 9127 -5530
rect 9027 -5624 9127 -5576
rect 9027 -5670 9054 -5624
rect 9100 -5670 9127 -5624
rect 9027 -5718 9127 -5670
rect 9027 -5764 9054 -5718
rect 9100 -5764 9127 -5718
rect 9027 -5812 9127 -5764
rect 9027 -5858 9054 -5812
rect 9100 -5858 9127 -5812
rect 9027 -5906 9127 -5858
rect 5103 -6155 6283 -5944
rect 2729 -6343 3229 -6328
rect 2729 -6376 2829 -6343
rect 2729 -6422 2756 -6376
rect 2802 -6422 2829 -6376
rect 2729 -6470 2829 -6422
rect 2729 -6516 2756 -6470
rect 2802 -6516 2829 -6470
rect 2729 -6564 2829 -6516
rect 2729 -6610 2756 -6564
rect 2802 -6610 2829 -6564
rect 2729 -6658 2829 -6610
rect 4622 -6433 4833 -6257
rect 5103 -6331 5314 -6155
rect 5591 -6433 5802 -6257
rect 6072 -6331 6283 -6155
rect 7015 -6151 8195 -5940
rect 4622 -6644 5802 -6433
rect 6542 -6424 6753 -6248
rect 7015 -6331 7226 -6151
rect 7511 -6424 7722 -6248
rect 7984 -6331 8195 -6151
rect 9027 -5952 9054 -5906
rect 9100 -5952 9127 -5906
rect 9027 -6000 9127 -5952
rect 9027 -6046 9054 -6000
rect 9100 -6046 9127 -6000
rect 9027 -6094 9127 -6046
rect 9027 -6140 9054 -6094
rect 9100 -6140 9127 -6094
rect 9027 -6188 9127 -6140
rect 9027 -6234 9054 -6188
rect 9100 -6234 9127 -6188
rect 9027 -6235 9127 -6234
rect 8562 -6282 9127 -6235
rect 8562 -6328 9054 -6282
rect 9100 -6328 9127 -6282
rect 8562 -6358 9127 -6328
rect 6542 -6635 7722 -6424
rect 9027 -6376 9127 -6358
rect 9027 -6422 9054 -6376
rect 9100 -6422 9127 -6376
rect 9027 -6470 9127 -6422
rect 9027 -6516 9054 -6470
rect 9100 -6516 9127 -6470
rect 9027 -6564 9127 -6516
rect 9027 -6610 9054 -6564
rect 9100 -6610 9127 -6564
rect 2729 -6704 2756 -6658
rect 2802 -6704 2829 -6658
rect 2729 -6752 2829 -6704
rect 2729 -6798 2756 -6752
rect 2802 -6798 2829 -6752
rect 2729 -6846 2829 -6798
rect 2729 -6892 2756 -6846
rect 2802 -6892 2829 -6846
rect 2729 -6940 2829 -6892
rect 2729 -6986 2756 -6940
rect 2802 -6986 2829 -6940
rect 2729 -7034 2829 -6986
rect 2729 -7080 2756 -7034
rect 2802 -7080 2829 -7034
rect 2729 -7128 2829 -7080
rect 2729 -7174 2756 -7128
rect 2802 -7174 2829 -7128
rect 2729 -7222 2829 -7174
rect 2729 -7268 2756 -7222
rect 2802 -7268 2829 -7222
rect 2729 -7316 2829 -7268
rect 2729 -7362 2756 -7316
rect 2802 -7362 2829 -7316
rect 2729 -7410 2829 -7362
rect 2729 -7456 2756 -7410
rect 2802 -7456 2829 -7410
rect 2729 -7504 2829 -7456
rect 2729 -7550 2756 -7504
rect 2802 -7550 2829 -7504
rect 2729 -7598 2829 -7550
rect 2729 -7644 2756 -7598
rect 2802 -7644 2829 -7598
rect 2729 -7692 2829 -7644
rect 9027 -6658 9127 -6610
rect 9027 -6704 9054 -6658
rect 9100 -6704 9127 -6658
rect 9027 -6752 9127 -6704
rect 9027 -6798 9054 -6752
rect 9100 -6798 9127 -6752
rect 9027 -6846 9127 -6798
rect 9027 -6892 9054 -6846
rect 9100 -6892 9127 -6846
rect 9027 -6940 9127 -6892
rect 9027 -6986 9054 -6940
rect 9100 -6986 9127 -6940
rect 9027 -7034 9127 -6986
rect 9027 -7080 9054 -7034
rect 9100 -7080 9127 -7034
rect 9027 -7128 9127 -7080
rect 9027 -7174 9054 -7128
rect 9100 -7174 9127 -7128
rect 9027 -7222 9127 -7174
rect 9027 -7268 9054 -7222
rect 9100 -7268 9127 -7222
rect 9027 -7316 9127 -7268
rect 9027 -7362 9054 -7316
rect 9100 -7362 9127 -7316
rect 9027 -7410 9127 -7362
rect 9027 -7456 9054 -7410
rect 9100 -7456 9127 -7410
rect 9027 -7504 9127 -7456
rect 9027 -7550 9054 -7504
rect 9100 -7550 9127 -7504
rect 9027 -7598 9127 -7550
rect 9027 -7644 9054 -7598
rect 9100 -7644 9127 -7598
rect 2729 -7738 2756 -7692
rect 2802 -7738 2829 -7692
rect 2729 -7786 2829 -7738
rect 2729 -7832 2756 -7786
rect 2802 -7832 2829 -7786
rect 2729 -7880 2829 -7832
rect 2729 -7926 2756 -7880
rect 2802 -7926 2829 -7880
rect 2729 -7962 2829 -7926
rect 4137 -7877 5317 -7666
rect 2729 -7974 3245 -7962
rect 2729 -8020 2756 -7974
rect 2802 -8020 3245 -7974
rect 2729 -8068 3245 -8020
rect 2729 -8114 2756 -8068
rect 2802 -8085 3245 -8068
rect 2802 -8114 2829 -8085
rect 2729 -8162 2829 -8114
rect 2729 -8208 2756 -8162
rect 2802 -8208 2829 -8162
rect 2729 -8256 2829 -8208
rect 2729 -8302 2756 -8256
rect 2802 -8302 2829 -8256
rect 2729 -8350 2829 -8302
rect 2729 -8396 2756 -8350
rect 2802 -8396 2829 -8350
rect 3656 -8155 3867 -7979
rect 4137 -8053 4348 -7877
rect 4625 -8155 4836 -7979
rect 5106 -8053 5317 -7877
rect 6049 -7873 7229 -7662
rect 3656 -8366 4836 -8155
rect 5592 -8155 5803 -7979
rect 6049 -8053 6260 -7873
rect 6561 -8155 6772 -7979
rect 7018 -8053 7229 -7873
rect 9027 -7692 9127 -7644
rect 9027 -7738 9054 -7692
rect 9100 -7738 9127 -7692
rect 9027 -7786 9127 -7738
rect 9027 -7832 9054 -7786
rect 9100 -7832 9127 -7786
rect 9027 -7880 9127 -7832
rect 9027 -7926 9054 -7880
rect 9100 -7926 9127 -7880
rect 9027 -7962 9127 -7926
rect 8571 -7974 9127 -7962
rect 5592 -8366 6772 -8155
rect 7509 -8191 7720 -7992
rect 7509 -8243 7540 -8191
rect 7592 -8243 7644 -8191
rect 7696 -8243 7720 -8191
rect 7509 -8295 7720 -8243
rect 7509 -8304 7540 -8295
rect 7528 -8347 7540 -8304
rect 7592 -8347 7644 -8295
rect 7696 -8304 7720 -8295
rect 7991 -8179 8202 -7995
rect 8571 -8020 9054 -7974
rect 9100 -8020 9127 -7974
rect 8571 -8068 9127 -8020
rect 8571 -8085 9054 -8068
rect 7991 -8231 8020 -8179
rect 8072 -8231 8124 -8179
rect 8176 -8231 8202 -8179
rect 7991 -8283 8202 -8231
rect 7991 -8304 8020 -8283
rect 7696 -8347 7708 -8304
rect 2729 -8444 2829 -8396
rect 2729 -8490 2756 -8444
rect 2802 -8490 2829 -8444
rect 7528 -8399 7708 -8347
rect 7528 -8451 7540 -8399
rect 7592 -8451 7644 -8399
rect 7696 -8451 7708 -8399
rect 8008 -8335 8020 -8304
rect 8072 -8335 8124 -8283
rect 8176 -8304 8202 -8283
rect 9027 -8114 9054 -8085
rect 9100 -8114 9127 -8068
rect 9027 -8162 9127 -8114
rect 9027 -8208 9054 -8162
rect 9100 -8208 9127 -8162
rect 9027 -8256 9127 -8208
rect 9027 -8302 9054 -8256
rect 9100 -8302 9127 -8256
rect 8176 -8335 8188 -8304
rect 8008 -8387 8188 -8335
rect 8008 -8439 8020 -8387
rect 8072 -8439 8124 -8387
rect 8176 -8439 8188 -8387
rect 8008 -8451 8188 -8439
rect 9027 -8350 9127 -8302
rect 9027 -8396 9054 -8350
rect 9100 -8396 9127 -8350
rect 9027 -8444 9127 -8396
rect 7528 -8463 7708 -8451
rect 2729 -8538 2829 -8490
rect 2729 -8584 2756 -8538
rect 2802 -8584 2829 -8538
rect 2729 -8605 2829 -8584
rect 9027 -8490 9054 -8444
rect 9100 -8490 9127 -8444
rect 9027 -8538 9127 -8490
rect 9027 -8584 9054 -8538
rect 9100 -8584 9127 -8538
rect 9027 -8605 9127 -8584
rect 2729 -8632 9127 -8605
rect 2729 -8678 2756 -8632
rect 2802 -8678 2850 -8632
rect 2896 -8678 2944 -8632
rect 2990 -8678 3038 -8632
rect 3084 -8678 3132 -8632
rect 3178 -8678 3226 -8632
rect 3272 -8678 3320 -8632
rect 3366 -8678 3414 -8632
rect 3460 -8678 3508 -8632
rect 3554 -8678 3602 -8632
rect 3648 -8678 3696 -8632
rect 3742 -8678 3790 -8632
rect 3836 -8678 3884 -8632
rect 3930 -8678 3978 -8632
rect 4024 -8678 4072 -8632
rect 4118 -8678 4166 -8632
rect 4212 -8678 4260 -8632
rect 4306 -8678 4354 -8632
rect 4400 -8678 4448 -8632
rect 4494 -8678 4542 -8632
rect 4588 -8678 4636 -8632
rect 4682 -8678 4730 -8632
rect 4776 -8678 4824 -8632
rect 4870 -8678 4918 -8632
rect 4964 -8678 5012 -8632
rect 5058 -8678 5106 -8632
rect 5152 -8678 5200 -8632
rect 5246 -8678 5294 -8632
rect 5340 -8678 5388 -8632
rect 5434 -8678 5482 -8632
rect 5528 -8678 5576 -8632
rect 5622 -8678 5670 -8632
rect 5716 -8678 5764 -8632
rect 5810 -8678 5858 -8632
rect 5904 -8678 5952 -8632
rect 5998 -8678 6046 -8632
rect 6092 -8678 6140 -8632
rect 6186 -8678 6234 -8632
rect 6280 -8678 6328 -8632
rect 6374 -8678 6422 -8632
rect 6468 -8678 6516 -8632
rect 6562 -8678 6610 -8632
rect 6656 -8678 6704 -8632
rect 6750 -8678 6798 -8632
rect 6844 -8678 6892 -8632
rect 6938 -8678 6986 -8632
rect 7032 -8678 7080 -8632
rect 7126 -8678 7174 -8632
rect 7220 -8678 7268 -8632
rect 7314 -8678 7362 -8632
rect 7408 -8678 7456 -8632
rect 7502 -8678 7550 -8632
rect 7596 -8678 7644 -8632
rect 7690 -8678 7738 -8632
rect 7784 -8678 7832 -8632
rect 7878 -8678 7926 -8632
rect 7972 -8678 8020 -8632
rect 8066 -8678 8114 -8632
rect 8160 -8678 8208 -8632
rect 8254 -8678 8302 -8632
rect 8348 -8678 8396 -8632
rect 8442 -8678 8490 -8632
rect 8536 -8678 8584 -8632
rect 8630 -8678 8678 -8632
rect 8724 -8678 8772 -8632
rect 8818 -8678 8866 -8632
rect 8912 -8678 8960 -8632
rect 9006 -8678 9054 -8632
rect 9100 -8678 9127 -8632
rect 2729 -8705 9127 -8678
rect 9589 -6561 9968 -6442
rect 12203 -6470 12572 -6443
rect 12203 -6540 12226 -6470
rect 12295 -6540 12347 -6470
rect 12416 -6540 12572 -6470
rect -13620 -9800 -3265 -9409
rect 9589 -9466 9708 -6561
rect 12203 -6562 12572 -6540
rect 10527 -8333 10949 -7945
rect 13078 -8333 13500 -7950
rect 14372 -8333 14977 -4126
rect 16144 -4277 16565 -3145
rect 18985 -4260 19406 -3145
rect 20566 -3153 20997 -3145
rect 21043 -3153 21070 -3107
rect 20566 -3201 21070 -3153
rect 20566 -3247 20997 -3201
rect 21043 -3247 21070 -3201
rect 20566 -3295 21070 -3247
rect 20566 -3341 20997 -3295
rect 21043 -3341 21070 -3295
rect 20566 -3389 21070 -3341
rect 20566 -3435 20997 -3389
rect 21043 -3435 21070 -3389
rect 20566 -3483 21070 -3435
rect 20566 -3529 20997 -3483
rect 21043 -3529 21070 -3483
rect 20566 -3577 21070 -3529
rect 20566 -3623 20997 -3577
rect 21043 -3623 21070 -3577
rect 20566 -3671 21070 -3623
rect 20566 -3717 20997 -3671
rect 21043 -3717 21070 -3671
rect 27268 -2683 27295 -2637
rect 27341 -2683 27368 -2637
rect 27268 -2731 27368 -2683
rect 27268 -2777 27295 -2731
rect 27341 -2777 27368 -2731
rect 27268 -2825 27368 -2777
rect 27268 -2871 27295 -2825
rect 27341 -2871 27368 -2825
rect 27268 -2919 27368 -2871
rect 27268 -2965 27295 -2919
rect 27341 -2965 27368 -2919
rect 27268 -3013 27368 -2965
rect 27268 -3059 27295 -3013
rect 27341 -3059 27368 -3013
rect 27268 -3107 27368 -3059
rect 27268 -3153 27295 -3107
rect 27341 -3153 27368 -3107
rect 27268 -3201 27368 -3153
rect 27268 -3247 27295 -3201
rect 27341 -3247 27368 -3201
rect 27268 -3295 27368 -3247
rect 27268 -3341 27295 -3295
rect 27341 -3341 27368 -3295
rect 27268 -3389 27368 -3341
rect 27268 -3435 27295 -3389
rect 27341 -3435 27368 -3389
rect 27268 -3483 27368 -3435
rect 27268 -3529 27295 -3483
rect 27341 -3529 27368 -3483
rect 27268 -3577 27368 -3529
rect 27268 -3623 27295 -3577
rect 27341 -3623 27368 -3577
rect 27268 -3671 27368 -3623
rect 20566 -3765 21070 -3717
rect 20566 -3811 20997 -3765
rect 21043 -3811 21070 -3765
rect 20566 -3859 21070 -3811
rect 20566 -3905 20997 -3859
rect 21043 -3905 21070 -3859
rect 20566 -3953 21070 -3905
rect 20566 -3999 20997 -3953
rect 21043 -3987 21070 -3953
rect 22892 -3895 24072 -3684
rect 21043 -3999 21509 -3987
rect 20566 -4047 21509 -3999
rect 20566 -4093 20997 -4047
rect 21043 -4093 21509 -4047
rect 20566 -4110 21509 -4093
rect 20566 -4141 21070 -4110
rect 20566 -4187 20997 -4141
rect 21043 -4187 21070 -4141
rect 20566 -4235 21070 -4187
rect 20566 -4281 20997 -4235
rect 21043 -4281 21070 -4235
rect 20566 -4329 21070 -4281
rect 20566 -4375 20997 -4329
rect 21043 -4375 21070 -4329
rect 20566 -4423 21070 -4375
rect 20566 -4469 20997 -4423
rect 21043 -4469 21070 -4423
rect 20566 -4517 21070 -4469
rect 20566 -4563 20997 -4517
rect 21043 -4563 21070 -4517
rect 20566 -4611 21070 -4563
rect 20566 -4657 20997 -4611
rect 21043 -4657 21070 -4611
rect 20566 -4705 21070 -4657
rect 20566 -4751 20997 -4705
rect 21043 -4751 21070 -4705
rect 20566 -4793 21070 -4751
rect 20566 -4799 21514 -4793
rect 20566 -4845 20997 -4799
rect 21043 -4845 21514 -4799
rect 20566 -4893 21514 -4845
rect 21925 -4887 22136 -4011
rect 22418 -4887 22629 -4011
rect 22892 -4071 23103 -3895
rect 23373 -4173 23584 -3997
rect 23861 -4071 24072 -3895
rect 24812 -3904 25992 -3693
rect 24342 -4173 24553 -3997
rect 24812 -4080 25023 -3904
rect 23373 -4384 24553 -4173
rect 25285 -4177 25496 -3997
rect 25781 -4080 25992 -3904
rect 27268 -3717 27295 -3671
rect 27341 -3717 27368 -3671
rect 27268 -3765 27368 -3717
rect 27268 -3811 27295 -3765
rect 27341 -3811 27368 -3765
rect 27268 -3859 27368 -3811
rect 27268 -3905 27295 -3859
rect 27341 -3905 27368 -3859
rect 27268 -3953 27368 -3905
rect 27268 -3979 27295 -3953
rect 26254 -4177 26465 -3997
rect 26854 -3999 27295 -3979
rect 27341 -3999 27368 -3953
rect 26854 -4047 27368 -3999
rect 26854 -4093 27295 -4047
rect 27341 -4093 27368 -4047
rect 26854 -4102 27368 -4093
rect 25285 -4388 26465 -4177
rect 27268 -4141 27368 -4102
rect 27268 -4187 27295 -4141
rect 27341 -4187 27368 -4141
rect 27268 -4235 27368 -4187
rect 27268 -4281 27295 -4235
rect 27341 -4281 27368 -4235
rect 27268 -4329 27368 -4281
rect 27268 -4375 27295 -4329
rect 27341 -4375 27368 -4329
rect 27268 -4423 27368 -4375
rect 27268 -4469 27295 -4423
rect 27341 -4469 27368 -4423
rect 23373 -4725 24553 -4514
rect 20566 -4939 20997 -4893
rect 21043 -4916 21514 -4893
rect 21043 -4939 21070 -4916
rect 20566 -4987 21070 -4939
rect 20566 -5033 20997 -4987
rect 21043 -5033 21070 -4987
rect 20566 -5081 21070 -5033
rect 20566 -5127 20997 -5081
rect 21043 -5127 21070 -5081
rect 20566 -5175 21070 -5127
rect 20566 -5221 20997 -5175
rect 21043 -5221 21070 -5175
rect 22892 -5003 23103 -4827
rect 23373 -4901 23584 -4725
rect 23861 -5003 24072 -4827
rect 24342 -4901 24553 -4725
rect 25285 -4721 26465 -4510
rect 22892 -5214 24072 -5003
rect 24812 -4994 25023 -4818
rect 25285 -4901 25496 -4721
rect 25781 -4994 25992 -4818
rect 26254 -4901 26465 -4721
rect 27268 -4517 27368 -4469
rect 27268 -4563 27295 -4517
rect 27341 -4563 27368 -4517
rect 27268 -4611 27368 -4563
rect 27268 -4657 27295 -4611
rect 27341 -4657 27368 -4611
rect 27268 -4705 27368 -4657
rect 27268 -4751 27295 -4705
rect 27341 -4751 27368 -4705
rect 27268 -4790 27368 -4751
rect 26827 -4799 27368 -4790
rect 26827 -4845 27295 -4799
rect 27341 -4845 27368 -4799
rect 26827 -4893 27368 -4845
rect 26827 -4913 27295 -4893
rect 24812 -5205 25992 -4994
rect 27268 -4939 27295 -4913
rect 27341 -4939 27368 -4893
rect 27268 -4987 27368 -4939
rect 27268 -5033 27295 -4987
rect 27341 -5033 27368 -4987
rect 27268 -5081 27368 -5033
rect 27268 -5127 27295 -5081
rect 27341 -5127 27368 -5081
rect 27268 -5175 27368 -5127
rect 20566 -5269 21070 -5221
rect 20566 -5315 20997 -5269
rect 21043 -5315 21070 -5269
rect 20566 -5363 21070 -5315
rect 20566 -5409 20997 -5363
rect 21043 -5409 21070 -5363
rect 20566 -5457 21070 -5409
rect 20566 -5503 20997 -5457
rect 21043 -5503 21070 -5457
rect 20566 -5551 21070 -5503
rect 20566 -5597 20997 -5551
rect 21043 -5597 21070 -5551
rect 20566 -5645 21070 -5597
rect 20566 -5691 20997 -5645
rect 21043 -5691 21070 -5645
rect 20566 -5739 21070 -5691
rect 20566 -5785 20997 -5739
rect 21043 -5785 21070 -5739
rect 20566 -5833 21070 -5785
rect 20566 -5879 20997 -5833
rect 21043 -5879 21070 -5833
rect 20566 -5927 21070 -5879
rect 20566 -5973 20997 -5927
rect 21043 -5973 21070 -5927
rect 20566 -6021 21070 -5973
rect 20566 -6067 20997 -6021
rect 21043 -6067 21070 -6021
rect 20566 -6115 21070 -6067
rect 20566 -6161 20997 -6115
rect 21043 -6161 21070 -6115
rect 20566 -6209 21070 -6161
rect 20566 -6255 20997 -6209
rect 21043 -6255 21070 -6209
rect 27268 -5221 27295 -5175
rect 27341 -5221 27368 -5175
rect 27268 -5269 27368 -5221
rect 27268 -5315 27295 -5269
rect 27341 -5315 27368 -5269
rect 27268 -5363 27368 -5315
rect 27268 -5409 27295 -5363
rect 27341 -5409 27368 -5363
rect 27268 -5457 27368 -5409
rect 27268 -5503 27295 -5457
rect 27341 -5503 27368 -5457
rect 27268 -5551 27368 -5503
rect 27268 -5597 27295 -5551
rect 27341 -5597 27368 -5551
rect 27268 -5645 27368 -5597
rect 27268 -5691 27295 -5645
rect 27341 -5691 27368 -5645
rect 27268 -5739 27368 -5691
rect 27268 -5785 27295 -5739
rect 27341 -5785 27368 -5739
rect 27268 -5833 27368 -5785
rect 27268 -5879 27295 -5833
rect 27341 -5879 27368 -5833
rect 27268 -5927 27368 -5879
rect 27268 -5973 27295 -5927
rect 27341 -5973 27368 -5927
rect 27268 -6021 27368 -5973
rect 27268 -6067 27295 -6021
rect 27341 -6067 27368 -6021
rect 27268 -6115 27368 -6067
rect 27268 -6161 27295 -6115
rect 27341 -6161 27368 -6115
rect 27268 -6209 27368 -6161
rect 20566 -6303 21070 -6255
rect 20566 -6349 20997 -6303
rect 21043 -6349 21070 -6303
rect 20566 -6397 21070 -6349
rect 20566 -6443 20997 -6397
rect 21043 -6443 21070 -6397
rect 15195 -6465 15564 -6445
rect 15195 -6535 15223 -6465
rect 15292 -6535 15344 -6465
rect 15413 -6535 15564 -6465
rect 15195 -6564 15564 -6535
rect 17977 -6473 18368 -6451
rect 17977 -6543 18001 -6473
rect 18070 -6543 18122 -6473
rect 18191 -6543 18368 -6473
rect 17977 -6572 18368 -6543
rect 20566 -6491 21070 -6443
rect 20566 -6537 20997 -6491
rect 21043 -6525 21070 -6491
rect 22407 -6447 23587 -6236
rect 21043 -6537 21515 -6525
rect 20566 -6585 21515 -6537
rect 20566 -6631 20997 -6585
rect 21043 -6631 21515 -6585
rect 20566 -6648 21515 -6631
rect 20566 -6679 21070 -6648
rect 20566 -6725 20997 -6679
rect 21043 -6725 21070 -6679
rect 20566 -6773 21070 -6725
rect 20566 -6819 20997 -6773
rect 21043 -6819 21070 -6773
rect 20566 -6867 21070 -6819
rect 20566 -6913 20997 -6867
rect 21043 -6913 21070 -6867
rect 20566 -6961 21070 -6913
rect 21926 -6725 22137 -6549
rect 22407 -6623 22618 -6447
rect 22895 -6725 23106 -6549
rect 23376 -6623 23587 -6447
rect 24319 -6443 25499 -6232
rect 21926 -6936 23106 -6725
rect 23862 -6725 24073 -6549
rect 24319 -6623 24530 -6443
rect 24831 -6725 25042 -6549
rect 25288 -6623 25499 -6443
rect 27268 -6255 27295 -6209
rect 27341 -6255 27368 -6209
rect 27268 -6303 27368 -6255
rect 27268 -6349 27295 -6303
rect 27341 -6349 27368 -6303
rect 27268 -6397 27368 -6349
rect 27268 -6443 27295 -6397
rect 27341 -6443 27368 -6397
rect 27268 -6491 27368 -6443
rect 27268 -6524 27295 -6491
rect 26835 -6537 27295 -6524
rect 27341 -6537 27368 -6491
rect 23862 -6936 25042 -6725
rect 25779 -6833 25990 -6562
rect 25729 -6845 26013 -6833
rect 25729 -6897 25741 -6845
rect 25793 -6897 25845 -6845
rect 25897 -6897 25949 -6845
rect 26001 -6897 26013 -6845
rect 20566 -7007 20997 -6961
rect 21043 -7007 21070 -6961
rect 20566 -7055 21070 -7007
rect 20566 -7101 20997 -7055
rect 21043 -7101 21070 -7055
rect 20566 -7149 21070 -7101
rect 25729 -6949 26013 -6897
rect 25729 -7001 25741 -6949
rect 25793 -7001 25845 -6949
rect 25897 -7001 25949 -6949
rect 26001 -7001 26013 -6949
rect 25729 -7053 26013 -7001
rect 25729 -7105 25741 -7053
rect 25793 -7105 25845 -7053
rect 25897 -7105 25949 -7053
rect 26001 -7105 26013 -7053
rect 25729 -7117 26013 -7105
rect 20566 -7195 20997 -7149
rect 21043 -7195 21070 -7149
rect 20566 -7243 21070 -7195
rect 20566 -7289 20997 -7243
rect 21043 -7289 21070 -7243
rect 20566 -7337 21070 -7289
rect 20566 -7383 20997 -7337
rect 21043 -7383 21070 -7337
rect 20566 -7431 21070 -7383
rect 20566 -7477 20997 -7431
rect 21043 -7477 21070 -7431
rect 20566 -7525 21070 -7477
rect 20566 -7571 20997 -7525
rect 21043 -7571 21070 -7525
rect 20566 -7619 21070 -7571
rect 20566 -7665 20997 -7619
rect 21043 -7665 21070 -7619
rect 20566 -7713 21070 -7665
rect 20566 -7759 20997 -7713
rect 21043 -7759 21070 -7713
rect 20566 -7807 21070 -7759
rect 20566 -7853 20997 -7807
rect 21043 -7840 21070 -7807
rect 21926 -7767 23106 -7556
rect 21043 -7853 21507 -7840
rect 20566 -7901 21507 -7853
rect 16204 -8333 16626 -7923
rect 19109 -8333 19531 -7941
rect 10527 -8755 19531 -8333
rect 20566 -7947 20997 -7901
rect 21043 -7947 21507 -7901
rect 21926 -7943 22137 -7767
rect 20566 -7963 21507 -7947
rect 20566 -7995 21070 -7963
rect 20566 -8041 20997 -7995
rect 21043 -8041 21070 -7995
rect 20566 -8089 21070 -8041
rect 20566 -8135 20997 -8089
rect 21043 -8135 21070 -8089
rect 20566 -8183 21070 -8135
rect 20566 -8229 20997 -8183
rect 21043 -8229 21070 -8183
rect 20566 -8277 21070 -8229
rect 22407 -8045 22618 -7869
rect 22895 -7943 23106 -7767
rect 23862 -7767 25042 -7556
rect 23376 -8045 23587 -7869
rect 23862 -7943 24073 -7767
rect 22407 -8256 23587 -8045
rect 24319 -8049 24530 -7869
rect 24831 -7943 25042 -7767
rect 25288 -8049 25499 -7869
rect 25779 -7930 25990 -7117
rect 26261 -7443 26472 -6565
rect 26835 -6585 27368 -6537
rect 26835 -6631 27295 -6585
rect 27341 -6631 27368 -6585
rect 26835 -6647 27368 -6631
rect 27268 -6679 27368 -6647
rect 27268 -6725 27295 -6679
rect 27341 -6725 27368 -6679
rect 27268 -6773 27368 -6725
rect 27268 -6819 27295 -6773
rect 27341 -6819 27368 -6773
rect 27268 -6867 27368 -6819
rect 27268 -6913 27295 -6867
rect 27341 -6913 27368 -6867
rect 27268 -6961 27368 -6913
rect 27268 -7007 27295 -6961
rect 27341 -7007 27368 -6961
rect 27268 -7055 27368 -7007
rect 27268 -7101 27295 -7055
rect 27341 -7101 27368 -7055
rect 27268 -7149 27368 -7101
rect 27268 -7195 27295 -7149
rect 27341 -7195 27368 -7149
rect 27268 -7243 27368 -7195
rect 27268 -7289 27295 -7243
rect 27341 -7289 27368 -7243
rect 27268 -7337 27368 -7289
rect 27268 -7383 27295 -7337
rect 27341 -7383 27368 -7337
rect 27268 -7431 27368 -7383
rect 26230 -7455 26514 -7443
rect 26230 -7507 26242 -7455
rect 26294 -7507 26346 -7455
rect 26398 -7507 26450 -7455
rect 26502 -7507 26514 -7455
rect 26230 -7559 26514 -7507
rect 26230 -7611 26242 -7559
rect 26294 -7611 26346 -7559
rect 26398 -7611 26450 -7559
rect 26502 -7611 26514 -7559
rect 26230 -7663 26514 -7611
rect 26230 -7715 26242 -7663
rect 26294 -7715 26346 -7663
rect 26398 -7715 26450 -7663
rect 26502 -7715 26514 -7663
rect 26230 -7727 26514 -7715
rect 27268 -7477 27295 -7431
rect 27341 -7477 27368 -7431
rect 27268 -7525 27368 -7477
rect 27268 -7571 27295 -7525
rect 27341 -7571 27368 -7525
rect 27268 -7619 27368 -7571
rect 27268 -7665 27295 -7619
rect 27341 -7665 27368 -7619
rect 27268 -7713 27368 -7665
rect 26261 -7927 26472 -7727
rect 27268 -7759 27295 -7713
rect 27341 -7759 27368 -7713
rect 27268 -7807 27368 -7759
rect 27268 -7835 27295 -7807
rect 26846 -7853 27295 -7835
rect 27341 -7853 27368 -7807
rect 26846 -7901 27368 -7853
rect 26846 -7947 27295 -7901
rect 27341 -7947 27368 -7901
rect 26846 -7958 27368 -7947
rect 24319 -8260 25499 -8049
rect 27268 -7995 27368 -7958
rect 27268 -8041 27295 -7995
rect 27341 -8041 27368 -7995
rect 27268 -8089 27368 -8041
rect 27268 -8135 27295 -8089
rect 27341 -8135 27368 -8089
rect 27268 -8183 27368 -8135
rect 27268 -8229 27295 -8183
rect 27341 -8229 27368 -8183
rect 20566 -8323 20997 -8277
rect 21043 -8323 21070 -8277
rect 20566 -8371 21070 -8323
rect 20566 -8417 20997 -8371
rect 21043 -8417 21070 -8371
rect 20566 -8465 21070 -8417
rect 20566 -8511 20997 -8465
rect 21043 -8511 21070 -8465
rect 20566 -8559 21070 -8511
rect 20566 -8605 20997 -8559
rect 21043 -8605 21070 -8559
rect 20566 -8653 21070 -8605
rect 20566 -8699 20997 -8653
rect 21043 -8699 21070 -8653
rect 20566 -8747 21070 -8699
rect 10755 -9432 10992 -9399
rect 10755 -9466 10787 -9432
rect 9589 -9501 10787 -9466
rect 10857 -9433 10992 -9432
rect 10857 -9501 10912 -9433
rect 9589 -9502 10912 -9501
rect 10982 -9502 10992 -9433
rect 9589 -9553 10992 -9502
rect 9589 -9585 10787 -9553
rect 10755 -9622 10787 -9585
rect 10857 -9554 10992 -9553
rect 10857 -9622 10912 -9554
rect 10755 -9623 10912 -9622
rect 10982 -9623 10992 -9554
rect 10755 -9651 10992 -9623
rect -13620 -9852 -3983 -9800
rect -3931 -9852 -3879 -9800
rect -3827 -9852 -3775 -9800
rect -3723 -9805 -3265 -9800
rect -3723 -9852 -3617 -9805
rect -13620 -9857 -3617 -9852
rect -3565 -9857 -3513 -9805
rect -3461 -9857 -3409 -9805
rect -3357 -9857 -3265 -9805
rect -13620 -9902 -3265 -9857
rect -13620 -11061 -13127 -9902
rect -4048 -9904 -3265 -9902
rect -4048 -9956 -3983 -9904
rect -3931 -9956 -3879 -9904
rect -3827 -9956 -3775 -9904
rect -3723 -9909 -3265 -9904
rect -3723 -9956 -3617 -9909
rect -4048 -9961 -3617 -9956
rect -3565 -9961 -3513 -9909
rect -3461 -9961 -3409 -9909
rect -3357 -9961 -3265 -9909
rect -4048 -10008 -3265 -9961
rect -4048 -10060 -3983 -10008
rect -3931 -10060 -3879 -10008
rect -3827 -10060 -3775 -10008
rect -3723 -10013 -3265 -10008
rect -3723 -10060 -3617 -10013
rect -4048 -10065 -3617 -10060
rect -3565 -10065 -3513 -10013
rect -3461 -10065 -3409 -10013
rect -3357 -10065 -3265 -10013
rect -4048 -10197 -3265 -10065
rect -4048 -10249 -3977 -10197
rect -3925 -10249 -3873 -10197
rect -3821 -10249 -3769 -10197
rect -3717 -10202 -3265 -10197
rect -3717 -10249 -3611 -10202
rect -4048 -10254 -3611 -10249
rect -3559 -10254 -3507 -10202
rect -3455 -10254 -3403 -10202
rect -3351 -10254 -3265 -10202
rect -4048 -10301 -3265 -10254
rect -4048 -10353 -3977 -10301
rect -3925 -10353 -3873 -10301
rect -3821 -10353 -3769 -10301
rect -3717 -10306 -3265 -10301
rect -3717 -10353 -3611 -10306
rect -4048 -10358 -3611 -10353
rect -3559 -10358 -3507 -10306
rect -3455 -10358 -3403 -10306
rect -3351 -10358 -3265 -10306
rect -4048 -10405 -3265 -10358
rect -4048 -10457 -3977 -10405
rect -3925 -10457 -3873 -10405
rect -3821 -10457 -3769 -10405
rect -3717 -10410 -3265 -10405
rect -3717 -10457 -3611 -10410
rect -4048 -10462 -3611 -10457
rect -3559 -10462 -3507 -10410
rect -3455 -10462 -3403 -10410
rect -3351 -10462 -3265 -10410
rect -4048 -10574 -3265 -10462
rect -4048 -10626 -3985 -10574
rect -3933 -10626 -3881 -10574
rect -3829 -10626 -3777 -10574
rect -3725 -10579 -3265 -10574
rect -3725 -10626 -3619 -10579
rect -4048 -10631 -3619 -10626
rect -3567 -10631 -3515 -10579
rect -3463 -10631 -3411 -10579
rect -3359 -10631 -3265 -10579
rect -4048 -10678 -3265 -10631
rect -4048 -10730 -3985 -10678
rect -3933 -10730 -3881 -10678
rect -3829 -10730 -3777 -10678
rect -3725 -10683 -3265 -10678
rect -3725 -10730 -3619 -10683
rect -4048 -10735 -3619 -10730
rect -3567 -10735 -3515 -10683
rect -3463 -10735 -3411 -10683
rect -3359 -10735 -3265 -10683
rect -4048 -10782 -3265 -10735
rect -4048 -10834 -3985 -10782
rect -3933 -10834 -3881 -10782
rect -3829 -10834 -3777 -10782
rect -3725 -10787 -3265 -10782
rect -3725 -10834 -3619 -10787
rect -4048 -10839 -3619 -10834
rect -3567 -10839 -3515 -10787
rect -3463 -10839 -3411 -10787
rect -3359 -10839 -3265 -10787
rect -4048 -10974 -3265 -10839
rect -4048 -11026 -3961 -10974
rect -3909 -11026 -3857 -10974
rect -3805 -11026 -3753 -10974
rect -3701 -10979 -3265 -10974
rect -3701 -11026 -3595 -10979
rect -4048 -11031 -3595 -11026
rect -3543 -11031 -3491 -10979
rect -3439 -11031 -3387 -10979
rect -3335 -11031 -3265 -10979
rect -4048 -11060 -3265 -11031
rect -7872 -11061 -7379 -11060
rect -4081 -11061 -3265 -11060
rect 1034 -11061 1527 -11060
rect 7292 -11061 7785 -11060
rect 11481 -11061 11974 -8755
rect 14933 -11061 15426 -8755
rect 18593 -11061 19086 -8755
rect 20566 -8793 20997 -8747
rect 21043 -8793 21070 -8747
rect 20566 -8841 21070 -8793
rect 20566 -8887 20997 -8841
rect 21043 -8887 21070 -8841
rect 20566 -8935 21070 -8887
rect 20566 -8981 20997 -8935
rect 21043 -8981 21070 -8935
rect 20566 -9029 21070 -8981
rect 20566 -9075 20997 -9029
rect 21043 -9075 21070 -9029
rect 20566 -9123 21070 -9075
rect 20566 -9169 20997 -9123
rect 21043 -9169 21070 -9123
rect 20566 -9217 21070 -9169
rect 20566 -9263 20997 -9217
rect 21043 -9263 21070 -9217
rect 20566 -9311 21070 -9263
rect 27268 -8277 27368 -8229
rect 27268 -8323 27295 -8277
rect 27341 -8323 27368 -8277
rect 27268 -8371 27368 -8323
rect 27268 -8417 27295 -8371
rect 27341 -8417 27368 -8371
rect 27268 -8465 27368 -8417
rect 27268 -8511 27295 -8465
rect 27341 -8511 27368 -8465
rect 27268 -8559 27368 -8511
rect 27268 -8605 27295 -8559
rect 27341 -8605 27368 -8559
rect 27268 -8653 27368 -8605
rect 27268 -8699 27295 -8653
rect 27341 -8699 27368 -8653
rect 27268 -8747 27368 -8699
rect 27268 -8793 27295 -8747
rect 27341 -8793 27368 -8747
rect 27268 -8841 27368 -8793
rect 27268 -8887 27295 -8841
rect 27341 -8887 27368 -8841
rect 27268 -8935 27368 -8887
rect 27268 -8981 27295 -8935
rect 27341 -8981 27368 -8935
rect 27268 -9029 27368 -8981
rect 27268 -9075 27295 -9029
rect 27341 -9075 27368 -9029
rect 27268 -9123 27368 -9075
rect 27268 -9169 27295 -9123
rect 27341 -9169 27368 -9123
rect 27268 -9217 27368 -9169
rect 27268 -9263 27295 -9217
rect 27341 -9263 27368 -9217
rect 20566 -9357 20997 -9311
rect 21043 -9357 21070 -9311
rect 20566 -9405 21070 -9357
rect 20566 -9451 20997 -9405
rect 21043 -9451 21070 -9405
rect 20566 -9499 21070 -9451
rect 20566 -9545 20997 -9499
rect 21043 -9545 21070 -9499
rect 20566 -9577 21070 -9545
rect 22892 -9489 24072 -9278
rect 20566 -9593 21510 -9577
rect 20566 -9639 20997 -9593
rect 21043 -9639 21510 -9593
rect 20566 -9687 21510 -9639
rect 20566 -9733 20997 -9687
rect 21043 -9700 21510 -9687
rect 21043 -9733 21070 -9700
rect 20566 -9781 21070 -9733
rect 20566 -9827 20997 -9781
rect 21043 -9827 21070 -9781
rect 20566 -9875 21070 -9827
rect 20566 -9921 20997 -9875
rect 21043 -9921 21070 -9875
rect 20566 -9969 21070 -9921
rect 20566 -10015 20997 -9969
rect 21043 -10015 21070 -9969
rect 21925 -9803 22136 -9605
rect 21925 -9855 21949 -9803
rect 22001 -9855 22053 -9803
rect 22105 -9855 22136 -9803
rect 21925 -9907 22136 -9855
rect 21925 -9959 21949 -9907
rect 22001 -9959 22053 -9907
rect 22105 -9959 22136 -9907
rect 21925 -9991 22136 -9959
rect 22418 -9789 22629 -9605
rect 22892 -9665 23103 -9489
rect 22418 -9841 22446 -9789
rect 22498 -9841 22550 -9789
rect 22602 -9841 22629 -9789
rect 22418 -9893 22629 -9841
rect 22418 -9945 22446 -9893
rect 22498 -9945 22550 -9893
rect 22602 -9945 22629 -9893
rect 22418 -9991 22629 -9945
rect 23373 -9767 23584 -9591
rect 23861 -9665 24072 -9489
rect 24812 -9498 25992 -9287
rect 24342 -9767 24553 -9591
rect 24812 -9674 25023 -9498
rect 23373 -9978 24553 -9767
rect 25285 -9771 25496 -9591
rect 25781 -9674 25992 -9498
rect 27268 -9311 27368 -9263
rect 27268 -9357 27295 -9311
rect 27341 -9357 27368 -9311
rect 27268 -9405 27368 -9357
rect 27268 -9451 27295 -9405
rect 27341 -9451 27368 -9405
rect 27268 -9499 27368 -9451
rect 27268 -9545 27295 -9499
rect 27341 -9545 27368 -9499
rect 27268 -9557 27368 -9545
rect 26254 -9771 26465 -9591
rect 26840 -9593 27368 -9557
rect 26840 -9639 27295 -9593
rect 27341 -9639 27368 -9593
rect 26840 -9680 27368 -9639
rect 25285 -9982 26465 -9771
rect 27268 -9687 27368 -9680
rect 27268 -9733 27295 -9687
rect 27341 -9733 27368 -9687
rect 27268 -9781 27368 -9733
rect 27268 -9827 27295 -9781
rect 27341 -9827 27368 -9781
rect 27268 -9875 27368 -9827
rect 27268 -9921 27295 -9875
rect 27341 -9921 27368 -9875
rect 27268 -9969 27368 -9921
rect 20566 -10063 21070 -10015
rect 20566 -10109 20997 -10063
rect 21043 -10109 21070 -10063
rect 21937 -10011 22117 -9991
rect 21937 -10063 21949 -10011
rect 22001 -10063 22053 -10011
rect 22105 -10063 22117 -10011
rect 22434 -9997 22614 -9991
rect 22434 -10049 22446 -9997
rect 22498 -10049 22550 -9997
rect 22602 -10049 22614 -9997
rect 22434 -10061 22614 -10049
rect 27268 -10015 27295 -9969
rect 27341 -10015 27368 -9969
rect 21937 -10075 22117 -10063
rect 27268 -10063 27368 -10015
rect 20566 -10144 21070 -10109
rect 20970 -10157 21070 -10144
rect 20970 -10203 20997 -10157
rect 21043 -10203 21070 -10157
rect 20970 -10224 21070 -10203
rect 27268 -10109 27295 -10063
rect 27341 -10109 27368 -10063
rect 27268 -10157 27368 -10109
rect 27268 -10203 27295 -10157
rect 27341 -10203 27368 -10157
rect 27268 -10224 27368 -10203
rect 20970 -10251 27368 -10224
rect 20970 -10297 20997 -10251
rect 21043 -10297 21091 -10251
rect 21137 -10297 21185 -10251
rect 21231 -10297 21279 -10251
rect 21325 -10297 21373 -10251
rect 21419 -10297 21467 -10251
rect 21513 -10297 21561 -10251
rect 21607 -10297 21655 -10251
rect 21701 -10297 21749 -10251
rect 21795 -10297 21843 -10251
rect 21889 -10297 21937 -10251
rect 21983 -10297 22031 -10251
rect 22077 -10297 22125 -10251
rect 22171 -10297 22219 -10251
rect 22265 -10297 22313 -10251
rect 22359 -10297 22407 -10251
rect 22453 -10297 22501 -10251
rect 22547 -10297 22595 -10251
rect 22641 -10297 22689 -10251
rect 22735 -10297 22783 -10251
rect 22829 -10297 22877 -10251
rect 22923 -10297 22971 -10251
rect 23017 -10297 23065 -10251
rect 23111 -10297 23159 -10251
rect 23205 -10297 23253 -10251
rect 23299 -10297 23347 -10251
rect 23393 -10297 23441 -10251
rect 23487 -10297 23535 -10251
rect 23581 -10297 23629 -10251
rect 23675 -10297 23723 -10251
rect 23769 -10297 23817 -10251
rect 23863 -10297 23911 -10251
rect 23957 -10297 24005 -10251
rect 24051 -10297 24099 -10251
rect 24145 -10297 24193 -10251
rect 24239 -10297 24287 -10251
rect 24333 -10297 24381 -10251
rect 24427 -10297 24475 -10251
rect 24521 -10297 24569 -10251
rect 24615 -10297 24663 -10251
rect 24709 -10297 24757 -10251
rect 24803 -10297 24851 -10251
rect 24897 -10297 24945 -10251
rect 24991 -10297 25039 -10251
rect 25085 -10297 25133 -10251
rect 25179 -10297 25227 -10251
rect 25273 -10297 25321 -10251
rect 25367 -10297 25415 -10251
rect 25461 -10297 25509 -10251
rect 25555 -10297 25603 -10251
rect 25649 -10297 25697 -10251
rect 25743 -10297 25791 -10251
rect 25837 -10297 25885 -10251
rect 25931 -10297 25979 -10251
rect 26025 -10297 26073 -10251
rect 26119 -10297 26167 -10251
rect 26213 -10297 26261 -10251
rect 26307 -10297 26355 -10251
rect 26401 -10297 26449 -10251
rect 26495 -10297 26543 -10251
rect 26589 -10297 26637 -10251
rect 26683 -10297 26731 -10251
rect 26777 -10297 26825 -10251
rect 26871 -10297 26919 -10251
rect 26965 -10297 27013 -10251
rect 27059 -10297 27107 -10251
rect 27153 -10297 27201 -10251
rect 27247 -10297 27295 -10251
rect 27341 -10297 27368 -10251
rect 20970 -10324 27368 -10297
rect -13620 -11078 19086 -11061
rect -13620 -11130 -3961 -11078
rect -3909 -11130 -3857 -11078
rect -3805 -11130 -3753 -11078
rect -3701 -11083 19086 -11078
rect -3701 -11130 -3595 -11083
rect -13620 -11135 -3595 -11130
rect -3543 -11135 -3491 -11083
rect -3439 -11135 -3387 -11083
rect -3335 -11135 19086 -11083
rect -13620 -11182 19086 -11135
rect -13620 -11234 -3961 -11182
rect -3909 -11234 -3857 -11182
rect -3805 -11234 -3753 -11182
rect -3701 -11187 19086 -11182
rect -3701 -11234 -3595 -11187
rect -13620 -11239 -3595 -11234
rect -3543 -11239 -3491 -11187
rect -3439 -11239 -3387 -11187
rect -3335 -11239 19086 -11187
rect -13620 -11554 19086 -11239
rect -13620 -12599 -13127 -11554
rect -7872 -12599 -7379 -11554
rect -4081 -12599 -3588 -11554
rect 1034 -12599 1527 -11554
rect 7292 -12599 7785 -11554
rect 11481 -12599 11974 -11554
rect 14933 -12599 15426 -11554
rect 18593 -12599 19086 -11554
rect -18607 -12638 19086 -12599
rect -21398 -13054 19086 -12638
rect -18607 -13092 19086 -13054
<< via1 >>
rect -13829 11916 -13765 11981
rect -9917 11937 -9857 11997
rect -9804 11936 -9744 11996
rect -7165 11941 -7105 12001
rect -7051 11941 -6991 12001
rect -13264 6571 -13212 6623
rect -13160 6571 -13108 6623
rect -13056 6571 -13004 6623
rect -12850 6573 -12798 6625
rect -12746 6573 -12694 6625
rect -12642 6573 -12590 6625
rect -12487 6566 -12435 6618
rect -12383 6566 -12331 6618
rect -12279 6566 -12227 6618
rect -13264 6467 -13212 6519
rect -13160 6467 -13108 6519
rect -13056 6467 -13004 6519
rect -12850 6469 -12798 6521
rect -12746 6469 -12694 6521
rect -12642 6469 -12590 6521
rect -12487 6462 -12435 6514
rect -12383 6462 -12331 6514
rect -12279 6462 -12227 6514
rect -13264 6363 -13212 6415
rect -13160 6363 -13108 6415
rect -13056 6363 -13004 6415
rect -12850 6365 -12798 6417
rect -12746 6365 -12694 6417
rect -12642 6365 -12590 6417
rect -12487 6358 -12435 6410
rect -12383 6358 -12331 6410
rect -12279 6358 -12227 6410
rect -13262 6155 -13210 6207
rect -13158 6155 -13106 6207
rect -13054 6155 -13002 6207
rect -12820 6138 -12768 6190
rect -12716 6138 -12664 6190
rect -12612 6138 -12560 6190
rect -12457 6131 -12405 6183
rect -12353 6131 -12301 6183
rect -12249 6131 -12197 6183
rect -13262 6051 -13210 6103
rect -13158 6051 -13106 6103
rect -13054 6051 -13002 6103
rect -12820 6034 -12768 6086
rect -12716 6034 -12664 6086
rect -12612 6034 -12560 6086
rect -12457 6027 -12405 6079
rect -12353 6027 -12301 6079
rect -12249 6027 -12197 6079
rect -13262 5947 -13210 5999
rect -13158 5947 -13106 5999
rect -13054 5947 -13002 5999
rect -12820 5930 -12768 5982
rect -12716 5930 -12664 5982
rect -12612 5930 -12560 5982
rect -12457 5923 -12405 5975
rect -12353 5923 -12301 5975
rect -12249 5923 -12197 5975
rect -13262 5714 -13210 5766
rect -13158 5714 -13106 5766
rect -13054 5714 -13002 5766
rect -13262 5610 -13210 5662
rect -13158 5610 -13106 5662
rect -13054 5610 -13002 5662
rect -13262 5506 -13210 5558
rect -13158 5506 -13106 5558
rect -13054 5506 -13002 5558
rect 13989 152 14041 204
rect 14093 152 14145 204
rect 14197 152 14249 204
rect 14387 163 14439 215
rect 14491 163 14543 215
rect 14595 163 14647 215
rect 13989 48 14041 100
rect 14093 48 14145 100
rect 14197 48 14249 100
rect 14387 59 14439 111
rect 14491 59 14543 111
rect 14595 59 14647 111
rect 13989 -56 14041 -4
rect 14093 -56 14145 -4
rect 14197 -56 14249 -4
rect 14387 -45 14439 7
rect 14491 -45 14543 7
rect 14595 -45 14647 7
rect -14136 -3049 -14072 -2993
rect -10942 -3045 -10878 -3043
rect -10942 -3093 -10894 -3045
rect -10894 -3093 -10878 -3045
rect -10942 -3099 -10878 -3093
rect 25800 -1921 25852 -1869
rect 25904 -1921 25956 -1869
rect 26289 -1922 26341 -1870
rect 26393 -1922 26445 -1870
rect 25800 -2025 25852 -1973
rect 25904 -2025 25956 -1973
rect 25800 -2129 25852 -2077
rect 25904 -2129 25956 -2077
rect 26289 -2026 26341 -1974
rect 26393 -2026 26445 -1974
rect 26289 -2130 26341 -2078
rect 26393 -2130 26445 -2078
rect -10128 -3045 -10050 -2975
rect -7377 -3046 -7299 -2976
rect 7531 -3415 7583 -3363
rect 7635 -3415 7687 -3363
rect 7531 -3519 7583 -3467
rect 7635 -3519 7687 -3467
rect 8018 -3411 8070 -3359
rect 8122 -3411 8174 -3359
rect 8018 -3515 8070 -3463
rect 8122 -3515 8174 -3463
rect 7531 -3623 7583 -3571
rect 7635 -3623 7687 -3571
rect 8018 -3619 8070 -3567
rect 8122 -3619 8174 -3567
rect 14130 -3574 14182 -3522
rect 14234 -3574 14286 -3522
rect 14338 -3574 14390 -3522
rect 14462 -3569 14514 -3517
rect 14566 -3569 14618 -3517
rect 14670 -3569 14722 -3517
rect 14130 -3678 14182 -3626
rect 14234 -3678 14286 -3626
rect 14338 -3678 14390 -3626
rect 14462 -3673 14514 -3621
rect 14566 -3673 14618 -3621
rect 14670 -3673 14722 -3621
rect 14130 -3782 14182 -3730
rect 14234 -3782 14286 -3730
rect 14338 -3782 14390 -3730
rect 14462 -3777 14514 -3725
rect 14566 -3777 14618 -3725
rect 14670 -3777 14722 -3725
rect 14464 -3918 14516 -3866
rect 14568 -3918 14620 -3866
rect 14672 -3918 14724 -3866
rect 14464 -4022 14516 -3970
rect 14568 -4022 14620 -3970
rect 14672 -4022 14724 -3970
rect 14464 -4126 14516 -4074
rect 14568 -4126 14620 -4074
rect 14672 -4126 14724 -4074
rect 7540 -8243 7592 -8191
rect 7644 -8243 7696 -8191
rect 7540 -8347 7592 -8295
rect 7644 -8347 7696 -8295
rect 8020 -8231 8072 -8179
rect 8124 -8231 8176 -8179
rect 7540 -8451 7592 -8399
rect 7644 -8451 7696 -8399
rect 8020 -8335 8072 -8283
rect 8124 -8335 8176 -8283
rect 8020 -8439 8072 -8387
rect 8124 -8439 8176 -8387
rect 12226 -6540 12295 -6470
rect 12347 -6540 12416 -6470
rect 15223 -6535 15292 -6465
rect 15344 -6535 15413 -6465
rect 18001 -6543 18070 -6473
rect 18122 -6543 18191 -6473
rect 25741 -6897 25793 -6845
rect 25845 -6897 25897 -6845
rect 25949 -6897 26001 -6845
rect 25741 -7001 25793 -6949
rect 25845 -7001 25897 -6949
rect 25949 -7001 26001 -6949
rect 25741 -7105 25793 -7053
rect 25845 -7105 25897 -7053
rect 25949 -7105 26001 -7053
rect 26242 -7507 26294 -7455
rect 26346 -7507 26398 -7455
rect 26450 -7507 26502 -7455
rect 26242 -7611 26294 -7559
rect 26346 -7611 26398 -7559
rect 26450 -7611 26502 -7559
rect 26242 -7715 26294 -7663
rect 26346 -7715 26398 -7663
rect 26450 -7715 26502 -7663
rect 10787 -9501 10857 -9432
rect 10912 -9502 10982 -9433
rect 10787 -9622 10857 -9553
rect 10912 -9623 10982 -9554
rect -3983 -9852 -3931 -9800
rect -3879 -9852 -3827 -9800
rect -3775 -9852 -3723 -9800
rect -3617 -9857 -3565 -9805
rect -3513 -9857 -3461 -9805
rect -3409 -9857 -3357 -9805
rect -3983 -9956 -3931 -9904
rect -3879 -9956 -3827 -9904
rect -3775 -9956 -3723 -9904
rect -3617 -9961 -3565 -9909
rect -3513 -9961 -3461 -9909
rect -3409 -9961 -3357 -9909
rect -3983 -10060 -3931 -10008
rect -3879 -10060 -3827 -10008
rect -3775 -10060 -3723 -10008
rect -3617 -10065 -3565 -10013
rect -3513 -10065 -3461 -10013
rect -3409 -10065 -3357 -10013
rect -3977 -10249 -3925 -10197
rect -3873 -10249 -3821 -10197
rect -3769 -10249 -3717 -10197
rect -3611 -10254 -3559 -10202
rect -3507 -10254 -3455 -10202
rect -3403 -10254 -3351 -10202
rect -3977 -10353 -3925 -10301
rect -3873 -10353 -3821 -10301
rect -3769 -10353 -3717 -10301
rect -3611 -10358 -3559 -10306
rect -3507 -10358 -3455 -10306
rect -3403 -10358 -3351 -10306
rect -3977 -10457 -3925 -10405
rect -3873 -10457 -3821 -10405
rect -3769 -10457 -3717 -10405
rect -3611 -10462 -3559 -10410
rect -3507 -10462 -3455 -10410
rect -3403 -10462 -3351 -10410
rect -3985 -10626 -3933 -10574
rect -3881 -10626 -3829 -10574
rect -3777 -10626 -3725 -10574
rect -3619 -10631 -3567 -10579
rect -3515 -10631 -3463 -10579
rect -3411 -10631 -3359 -10579
rect -3985 -10730 -3933 -10678
rect -3881 -10730 -3829 -10678
rect -3777 -10730 -3725 -10678
rect -3619 -10735 -3567 -10683
rect -3515 -10735 -3463 -10683
rect -3411 -10735 -3359 -10683
rect -3985 -10834 -3933 -10782
rect -3881 -10834 -3829 -10782
rect -3777 -10834 -3725 -10782
rect -3619 -10839 -3567 -10787
rect -3515 -10839 -3463 -10787
rect -3411 -10839 -3359 -10787
rect -3961 -11026 -3909 -10974
rect -3857 -11026 -3805 -10974
rect -3753 -11026 -3701 -10974
rect -3595 -11031 -3543 -10979
rect -3491 -11031 -3439 -10979
rect -3387 -11031 -3335 -10979
rect 21949 -9855 22001 -9803
rect 22053 -9855 22105 -9803
rect 21949 -9959 22001 -9907
rect 22053 -9959 22105 -9907
rect 22446 -9841 22498 -9789
rect 22550 -9841 22602 -9789
rect 22446 -9945 22498 -9893
rect 22550 -9945 22602 -9893
rect 21949 -10063 22001 -10011
rect 22053 -10063 22105 -10011
rect 22446 -10049 22498 -9997
rect 22550 -10049 22602 -9997
rect -3961 -11130 -3909 -11078
rect -3857 -11130 -3805 -11078
rect -3753 -11130 -3701 -11078
rect -3595 -11135 -3543 -11083
rect -3491 -11135 -3439 -11083
rect -3387 -11135 -3335 -11083
rect -3961 -11234 -3909 -11182
rect -3857 -11234 -3805 -11182
rect -3753 -11234 -3701 -11182
rect -3595 -11239 -3543 -11187
rect -3491 -11239 -3439 -11187
rect -3387 -11239 -3335 -11187
<< metal2 >>
rect 31218 14648 31502 15282
rect -1780 14386 -1349 14435
rect -1780 14330 -1762 14386
rect -1706 14330 -1658 14386
rect -1602 14330 -1554 14386
rect -1498 14330 -1349 14386
rect -1780 14282 -1349 14330
rect -1780 14226 -1762 14282
rect -1706 14226 -1658 14282
rect -1602 14226 -1554 14282
rect -1498 14226 -1349 14282
rect -1780 14178 -1349 14226
rect -1780 14122 -1762 14178
rect -1706 14122 -1658 14178
rect -1602 14122 -1554 14178
rect -1498 14122 -1349 14178
rect -13537 12937 -5324 13128
rect -14618 12525 -14334 12535
rect -14618 12469 -14608 12525
rect -14552 12469 -14504 12525
rect -14448 12469 -14400 12525
rect -14344 12469 -14334 12525
rect -14618 12431 -14334 12469
rect -14618 12421 -12768 12431
rect -14618 12365 -14608 12421
rect -14552 12365 -14504 12421
rect -14448 12365 -14400 12421
rect -14344 12365 -12768 12421
rect -14618 12317 -12768 12365
rect -14618 12261 -14608 12317
rect -14552 12261 -14504 12317
rect -14448 12261 -14400 12317
rect -14344 12306 -12768 12317
rect -14344 12261 -14334 12306
rect -14618 12251 -14334 12261
rect -15663 11981 -13711 12006
rect -15663 11916 -13829 11981
rect -13765 11916 -13711 11981
rect -15663 11892 -13711 11916
rect -15663 -2962 -15351 11892
rect -11238 7764 -10820 12937
rect -9337 12295 -5487 12470
rect -9952 11997 -9728 12025
rect -9952 11937 -9917 11997
rect -9857 11996 -9728 11997
rect -9857 11937 -9804 11996
rect -9952 11936 -9804 11937
rect -9744 11936 -9728 11996
rect -9952 11908 -9728 11936
rect -8927 12004 -8648 12037
rect -8927 11926 -8890 12004
rect -8824 11926 -8755 12004
rect -8689 11926 -8648 12004
rect -8927 8735 -8648 11926
rect -7735 9435 -7367 12295
rect -7207 12023 -7082 12024
rect -7207 12001 -6972 12023
rect -7207 11941 -7165 12001
rect -7105 11941 -7051 12001
rect -6991 11941 -6972 12001
rect -7207 11918 -6972 11941
rect -8082 9375 -7354 9435
rect -8082 9319 -8056 9375
rect -8000 9319 -7952 9375
rect -7896 9319 -7848 9375
rect -7792 9374 -7354 9375
rect -7792 9319 -7720 9374
rect -8082 9318 -7720 9319
rect -7664 9318 -7616 9374
rect -7560 9318 -7512 9374
rect -7456 9318 -7354 9374
rect -8082 9271 -7354 9318
rect -8082 9215 -8056 9271
rect -8000 9215 -7952 9271
rect -7896 9215 -7848 9271
rect -7792 9270 -7354 9271
rect -7792 9215 -7720 9270
rect -8082 9214 -7720 9215
rect -7664 9214 -7616 9270
rect -7560 9214 -7512 9270
rect -7456 9214 -7354 9270
rect -8082 9167 -7354 9214
rect -8082 9111 -8056 9167
rect -8000 9111 -7952 9167
rect -7896 9111 -7848 9167
rect -7792 9166 -7354 9167
rect -7792 9111 -7720 9166
rect -8082 9110 -7720 9111
rect -7664 9110 -7616 9166
rect -7560 9110 -7512 9166
rect -7456 9110 -7354 9166
rect -8082 9081 -7354 9110
rect -8927 8657 -8884 8735
rect -8818 8657 -8764 8735
rect -8698 8657 -8648 8735
rect -8927 8605 -8648 8657
rect -8927 8527 -8884 8605
rect -8818 8527 -8764 8605
rect -8698 8527 -8648 8605
rect -8927 8475 -8648 8527
rect -8927 8397 -8884 8475
rect -8818 8397 -8764 8475
rect -8698 8397 -8648 8475
rect -8927 8158 -8648 8397
rect -11238 7278 -2265 7764
rect -13337 6808 -3232 6828
rect -13338 6755 -3232 6808
rect -13338 6699 -4321 6755
rect -4265 6699 -4217 6755
rect -4161 6699 -4113 6755
rect -4057 6741 -3232 6755
rect -4057 6699 -3968 6741
rect -13338 6685 -3968 6699
rect -3912 6685 -3864 6741
rect -3808 6685 -3760 6741
rect -3704 6739 -3232 6741
rect -3704 6685 -3552 6739
rect -13338 6683 -3552 6685
rect -3496 6683 -3448 6739
rect -3392 6683 -3344 6739
rect -3288 6683 -3232 6739
rect -13338 6651 -3232 6683
rect -13338 6625 -4321 6651
rect -13338 6623 -12850 6625
rect -13338 6571 -13264 6623
rect -13212 6571 -13160 6623
rect -13108 6571 -13056 6623
rect -13004 6573 -12850 6623
rect -12798 6573 -12746 6625
rect -12694 6573 -12642 6625
rect -12590 6618 -4321 6625
rect -12590 6573 -12487 6618
rect -13004 6571 -12487 6573
rect -13338 6566 -12487 6571
rect -12435 6566 -12383 6618
rect -12331 6566 -12279 6618
rect -12227 6595 -4321 6618
rect -4265 6595 -4217 6651
rect -4161 6595 -4113 6651
rect -4057 6637 -3232 6651
rect -4057 6595 -3968 6637
rect -12227 6581 -3968 6595
rect -3912 6581 -3864 6637
rect -3808 6581 -3760 6637
rect -3704 6635 -3232 6637
rect -3704 6581 -3552 6635
rect -12227 6579 -3552 6581
rect -3496 6579 -3448 6635
rect -3392 6579 -3344 6635
rect -3288 6579 -3232 6635
rect -12227 6566 -3232 6579
rect -13338 6547 -3232 6566
rect -13338 6521 -4321 6547
rect -13338 6519 -12850 6521
rect -13338 6467 -13264 6519
rect -13212 6467 -13160 6519
rect -13108 6467 -13056 6519
rect -13004 6469 -12850 6519
rect -12798 6469 -12746 6521
rect -12694 6469 -12642 6521
rect -12590 6514 -4321 6521
rect -12590 6469 -12487 6514
rect -13004 6467 -12487 6469
rect -13338 6462 -12487 6467
rect -12435 6462 -12383 6514
rect -12331 6462 -12279 6514
rect -12227 6491 -4321 6514
rect -4265 6491 -4217 6547
rect -4161 6491 -4113 6547
rect -4057 6533 -3232 6547
rect -4057 6491 -3968 6533
rect -12227 6477 -3968 6491
rect -3912 6477 -3864 6533
rect -3808 6477 -3760 6533
rect -3704 6531 -3232 6533
rect -3704 6477 -3552 6531
rect -12227 6475 -3552 6477
rect -3496 6475 -3448 6531
rect -3392 6475 -3344 6531
rect -3288 6475 -3232 6531
rect -12227 6462 -3232 6475
rect -13338 6417 -3232 6462
rect -13338 6415 -12850 6417
rect -13338 6363 -13264 6415
rect -13212 6363 -13160 6415
rect -13108 6363 -13056 6415
rect -13004 6365 -12850 6415
rect -12798 6365 -12746 6417
rect -12694 6365 -12642 6417
rect -12590 6410 -3232 6417
rect -12590 6365 -12487 6410
rect -13004 6363 -12487 6365
rect -13338 6358 -12487 6363
rect -12435 6358 -12383 6410
rect -12331 6358 -12279 6410
rect -12227 6376 -3232 6410
rect -12227 6358 -4289 6376
rect -13338 6320 -4289 6358
rect -4233 6320 -4185 6376
rect -4129 6374 -3232 6376
rect -4129 6320 -4048 6374
rect -13338 6318 -4048 6320
rect -3992 6318 -3944 6374
rect -3888 6318 -3840 6374
rect -3784 6318 -3645 6374
rect -3589 6318 -3541 6374
rect -3485 6318 -3437 6374
rect -3381 6318 -3232 6374
rect -13338 6272 -3232 6318
rect -13338 6216 -4289 6272
rect -4233 6216 -4185 6272
rect -4129 6270 -3232 6272
rect -4129 6216 -4048 6270
rect -13338 6214 -4048 6216
rect -3992 6214 -3944 6270
rect -3888 6214 -3840 6270
rect -3784 6214 -3645 6270
rect -3589 6214 -3541 6270
rect -3485 6214 -3437 6270
rect -3381 6214 -3232 6270
rect -13338 6207 -3232 6214
rect -13338 6155 -13262 6207
rect -13210 6155 -13158 6207
rect -13106 6155 -13054 6207
rect -13002 6190 -3232 6207
rect -13002 6155 -12820 6190
rect -13338 6138 -12820 6155
rect -12768 6138 -12716 6190
rect -12664 6138 -12612 6190
rect -12560 6183 -3232 6190
rect -12560 6138 -12457 6183
rect -13338 6131 -12457 6138
rect -12405 6131 -12353 6183
rect -12301 6131 -12249 6183
rect -12197 6168 -3232 6183
rect -12197 6131 -4289 6168
rect -13338 6112 -4289 6131
rect -4233 6112 -4185 6168
rect -4129 6166 -3232 6168
rect -4129 6112 -4048 6166
rect -13338 6110 -4048 6112
rect -3992 6110 -3944 6166
rect -3888 6110 -3840 6166
rect -3784 6110 -3645 6166
rect -3589 6110 -3541 6166
rect -3485 6110 -3437 6166
rect -3381 6110 -3232 6166
rect -13338 6103 -3232 6110
rect -13338 6051 -13262 6103
rect -13210 6051 -13158 6103
rect -13106 6051 -13054 6103
rect -13002 6086 -3232 6103
rect -13002 6051 -12820 6086
rect -13338 6034 -12820 6051
rect -12768 6034 -12716 6086
rect -12664 6034 -12612 6086
rect -12560 6079 -3232 6086
rect -12560 6034 -12457 6079
rect -13338 6027 -12457 6034
rect -12405 6027 -12353 6079
rect -12301 6027 -12249 6079
rect -12197 6033 -3232 6079
rect -12197 6027 -4282 6033
rect -13338 5999 -4282 6027
rect -13338 5947 -13262 5999
rect -13210 5947 -13158 5999
rect -13106 5947 -13054 5999
rect -13002 5982 -4282 5999
rect -13002 5947 -12820 5982
rect -13338 5930 -12820 5947
rect -12768 5930 -12716 5982
rect -12664 5930 -12612 5982
rect -12560 5977 -4282 5982
rect -4226 5977 -4178 6033
rect -4122 6031 -3232 6033
rect -4122 5977 -4041 6031
rect -12560 5975 -4041 5977
rect -3985 5975 -3937 6031
rect -3881 5975 -3833 6031
rect -3777 5975 -3638 6031
rect -3582 5975 -3534 6031
rect -3478 5975 -3430 6031
rect -3374 5975 -3232 6031
rect -12560 5930 -12457 5975
rect -13338 5923 -12457 5930
rect -12405 5923 -12353 5975
rect -12301 5923 -12249 5975
rect -12197 5923 -3232 5975
rect -13338 5898 -3232 5923
rect -13338 5842 -4289 5898
rect -4233 5842 -4185 5898
rect -4129 5896 -3232 5898
rect -4129 5842 -4048 5896
rect -13338 5840 -4048 5842
rect -3992 5840 -3944 5896
rect -3888 5840 -3840 5896
rect -3784 5840 -3645 5896
rect -3589 5840 -3541 5896
rect -3485 5840 -3437 5896
rect -3381 5840 -3232 5896
rect -13338 5766 -3232 5840
rect -13338 5714 -13262 5766
rect -13210 5714 -13158 5766
rect -13106 5714 -13054 5766
rect -13002 5760 -3232 5766
rect -13002 5714 -12463 5760
rect -13338 5662 -12463 5714
rect -13338 5610 -13262 5662
rect -13210 5610 -13158 5662
rect -13106 5610 -13054 5662
rect -13002 5610 -12463 5662
rect -13338 5558 -12463 5610
rect -13338 5506 -13262 5558
rect -13210 5506 -13158 5558
rect -13106 5506 -13054 5558
rect -13002 5506 -12463 5558
rect -13338 5433 -12463 5506
rect -13338 5432 -12889 5433
rect -11415 -1803 -11131 -1793
rect -11415 -1847 -11405 -1803
rect -13815 -1859 -11405 -1847
rect -11349 -1859 -11301 -1803
rect -11245 -1859 -11197 -1803
rect -11141 -1847 -11131 -1803
rect -11141 -1859 -5602 -1847
rect -13815 -1907 -5602 -1859
rect -13815 -1963 -11405 -1907
rect -11349 -1963 -11301 -1907
rect -11245 -1963 -11197 -1907
rect -11141 -1963 -5602 -1907
rect -13815 -2011 -5602 -1963
rect -13815 -2038 -11405 -2011
rect -11415 -2067 -11405 -2038
rect -11349 -2067 -11301 -2011
rect -11245 -2067 -11197 -2011
rect -11141 -2038 -5602 -2011
rect -11141 -2067 -11131 -2038
rect -11415 -2077 -11131 -2067
rect -14896 -2450 -14612 -2440
rect -14896 -2506 -14886 -2450
rect -14830 -2506 -14782 -2450
rect -14726 -2506 -14678 -2450
rect -14622 -2506 -14612 -2450
rect -7968 -2453 -7643 -2432
rect -7968 -2505 -7953 -2453
rect -14896 -2544 -14612 -2506
rect -9615 -2509 -7953 -2505
rect -7897 -2509 -7849 -2453
rect -7793 -2509 -7745 -2453
rect -7689 -2505 -7643 -2453
rect -7689 -2509 -5765 -2505
rect -14896 -2554 -13046 -2544
rect -14896 -2610 -14886 -2554
rect -14830 -2610 -14782 -2554
rect -14726 -2610 -14678 -2554
rect -14622 -2610 -13046 -2554
rect -14896 -2658 -13046 -2610
rect -14896 -2714 -14886 -2658
rect -14830 -2714 -14782 -2658
rect -14726 -2714 -14678 -2658
rect -14622 -2669 -13046 -2658
rect -9615 -2557 -5765 -2509
rect -9615 -2613 -7953 -2557
rect -7897 -2613 -7849 -2557
rect -7793 -2613 -7745 -2557
rect -7689 -2613 -5765 -2557
rect -9615 -2661 -5765 -2613
rect -14622 -2714 -14612 -2669
rect -9615 -2680 -7953 -2661
rect -14896 -2724 -14612 -2714
rect -7968 -2717 -7953 -2680
rect -7897 -2717 -7849 -2661
rect -7793 -2717 -7745 -2661
rect -7689 -2680 -5765 -2661
rect -7689 -2717 -7643 -2680
rect -7967 -2737 -7643 -2717
rect -15663 -2993 -11534 -2962
rect -15663 -3049 -14136 -2993
rect -14072 -3023 -11534 -2993
rect -10170 -2975 -7231 -2953
rect -14072 -3043 -10810 -3023
rect -14072 -3049 -10942 -3043
rect -15663 -3073 -10942 -3049
rect -15663 -11960 -15351 -3073
rect -11645 -3099 -10942 -3073
rect -10878 -3099 -10810 -3043
rect -10170 -3045 -10128 -2975
rect -10050 -2976 -7231 -2975
rect -10050 -2978 -8744 -2976
rect -10050 -3045 -8905 -2978
rect -10170 -3056 -8905 -3045
rect -8839 -3054 -8744 -2978
rect -8678 -3046 -7377 -2976
rect -7299 -3046 -7231 -2976
rect -8678 -3054 -7231 -3046
rect -8839 -3056 -7231 -3054
rect -10170 -3070 -7231 -3056
rect -11645 -3134 -10810 -3099
rect -14956 -5588 -7648 -5557
rect -14956 -5590 -14531 -5588
rect -14956 -5646 -14913 -5590
rect -14857 -5646 -14809 -5590
rect -14753 -5646 -14705 -5590
rect -14649 -5644 -14531 -5590
rect -14475 -5644 -14427 -5588
rect -14371 -5644 -14323 -5588
rect -14267 -5596 -7648 -5588
rect -14267 -5644 -8354 -5596
rect -14649 -5646 -8354 -5644
rect -14956 -5652 -8354 -5646
rect -8298 -5652 -8250 -5596
rect -8194 -5652 -8146 -5596
rect -8090 -5601 -7648 -5596
rect -8090 -5652 -7998 -5601
rect -14956 -5657 -7998 -5652
rect -7942 -5657 -7894 -5601
rect -7838 -5657 -7790 -5601
rect -7734 -5657 -7648 -5601
rect -14956 -5692 -7648 -5657
rect -14956 -5694 -14531 -5692
rect -14956 -5750 -14913 -5694
rect -14857 -5750 -14809 -5694
rect -14753 -5750 -14705 -5694
rect -14649 -5748 -14531 -5694
rect -14475 -5748 -14427 -5692
rect -14371 -5748 -14323 -5692
rect -14267 -5700 -7648 -5692
rect -14267 -5748 -8354 -5700
rect -14649 -5750 -8354 -5748
rect -14956 -5756 -8354 -5750
rect -8298 -5756 -8250 -5700
rect -8194 -5756 -8146 -5700
rect -8090 -5705 -7648 -5700
rect -8090 -5756 -7998 -5705
rect -14956 -5761 -7998 -5756
rect -7942 -5761 -7894 -5705
rect -7838 -5761 -7790 -5705
rect -7734 -5761 -7648 -5705
rect -14956 -5796 -7648 -5761
rect -14956 -5798 -14531 -5796
rect -14956 -5854 -14913 -5798
rect -14857 -5854 -14809 -5798
rect -14753 -5854 -14705 -5798
rect -14649 -5852 -14531 -5798
rect -14475 -5852 -14427 -5796
rect -14371 -5852 -14323 -5796
rect -14267 -5804 -7648 -5796
rect -14267 -5852 -8354 -5804
rect -14649 -5854 -8354 -5852
rect -14956 -5860 -8354 -5854
rect -8298 -5860 -8250 -5804
rect -8194 -5860 -8146 -5804
rect -8090 -5809 -7648 -5804
rect -8090 -5860 -7998 -5809
rect -14956 -5865 -7998 -5860
rect -7942 -5865 -7894 -5809
rect -7838 -5865 -7790 -5809
rect -7734 -5865 -7648 -5809
rect -14956 -5882 -7648 -5865
rect -4283 -9800 -3269 5760
rect -2751 -6364 -2265 7278
rect -1780 -1034 -1349 14122
rect 32132 14045 32410 14744
rect -1048 13250 -617 13287
rect -1048 13194 -982 13250
rect -926 13194 -878 13250
rect -822 13194 -774 13250
rect -718 13194 -617 13250
rect -1048 13146 -617 13194
rect -1048 13090 -982 13146
rect -926 13090 -878 13146
rect -822 13090 -774 13146
rect -718 13090 -617 13146
rect -1048 13042 -617 13090
rect -1048 12986 -982 13042
rect -926 12986 -878 13042
rect -822 12986 -774 13042
rect -718 12986 -617 13042
rect -1048 -427 -617 12986
rect 6683 7072 6989 7091
rect 6683 7016 6707 7072
rect 6763 7016 6811 7072
rect 6867 7016 6915 7072
rect 6971 7016 6989 7072
rect 6683 6968 6989 7016
rect 6683 6912 6707 6968
rect 6763 6912 6811 6968
rect 6867 6912 6915 6968
rect 6971 6912 6989 6968
rect 6683 6864 6989 6912
rect 6683 6830 6707 6864
rect 6028 6808 6707 6830
rect 6763 6808 6811 6864
rect 6867 6808 6915 6864
rect 6971 6830 6989 6864
rect 9808 6977 10114 6996
rect 9808 6921 9832 6977
rect 9888 6921 9936 6977
rect 9992 6921 10040 6977
rect 10096 6921 10114 6977
rect 9808 6873 10114 6921
rect 16371 6960 16677 6979
rect 16371 6904 16395 6960
rect 16451 6904 16499 6960
rect 16555 6904 16603 6960
rect 16659 6904 16677 6960
rect 6971 6808 7022 6830
rect 6028 6745 7022 6808
rect 6028 6689 6149 6745
rect 6205 6737 7022 6745
rect 6205 6689 6255 6737
rect 6028 6681 6255 6689
rect 6311 6681 6359 6737
rect 6415 6681 6463 6737
rect 6519 6734 7022 6737
rect 6519 6681 6654 6734
rect 6028 6678 6654 6681
rect 6710 6678 6758 6734
rect 6814 6678 6862 6734
rect 6918 6678 7022 6734
rect 9808 6817 9832 6873
rect 9888 6817 9936 6873
rect 9992 6817 10040 6873
rect 10096 6817 10114 6873
rect 9808 6769 10114 6817
rect 9808 6713 9832 6769
rect 9888 6713 9936 6769
rect 9992 6713 10040 6769
rect 10096 6713 10114 6769
rect 9808 6684 10114 6713
rect 15954 6868 16260 6887
rect 15954 6812 15978 6868
rect 16034 6812 16082 6868
rect 16138 6812 16186 6868
rect 16242 6812 16260 6868
rect 15954 6764 16260 6812
rect 15954 6708 15978 6764
rect 16034 6708 16082 6764
rect 16138 6708 16186 6764
rect 16242 6708 16260 6764
rect 6028 6641 7022 6678
rect 6028 6585 6149 6641
rect 6205 6633 7022 6641
rect 6205 6585 6255 6633
rect 6028 6577 6255 6585
rect 6311 6577 6359 6633
rect 6415 6577 6463 6633
rect 6519 6630 7022 6633
rect 6519 6577 6654 6630
rect 6028 6574 6654 6577
rect 6710 6574 6758 6630
rect 6814 6574 6862 6630
rect 6918 6574 7022 6630
rect 15954 6660 16260 6708
rect 16371 6856 16677 6904
rect 16371 6800 16395 6856
rect 16451 6800 16499 6856
rect 16555 6800 16603 6856
rect 16659 6800 16677 6856
rect 16371 6752 16677 6800
rect 16371 6696 16395 6752
rect 16451 6696 16499 6752
rect 16555 6696 16603 6752
rect 16659 6696 16677 6752
rect 16371 6667 16677 6696
rect 15954 6604 15978 6660
rect 16034 6604 16082 6660
rect 16138 6604 16186 6660
rect 16242 6604 16260 6660
rect 15954 6575 16260 6604
rect 6028 6537 7022 6574
rect 6028 6481 6149 6537
rect 6205 6529 7022 6537
rect 6205 6481 6255 6529
rect 6028 6473 6255 6481
rect 6311 6473 6359 6529
rect 6415 6473 6463 6529
rect 6519 6526 7022 6529
rect 6519 6473 6654 6526
rect 6028 6470 6654 6473
rect 6710 6470 6758 6526
rect 6814 6470 6862 6526
rect 6918 6470 7022 6526
rect 6028 6412 7022 6470
rect 6028 6394 6167 6412
rect 6143 6356 6167 6394
rect 6223 6356 6271 6412
rect 6327 6356 6375 6412
rect 6431 6394 7022 6412
rect 15951 6522 16257 6541
rect 15951 6466 15975 6522
rect 16031 6466 16079 6522
rect 16135 6466 16183 6522
rect 16239 6466 16257 6522
rect 15951 6418 16257 6466
rect 6431 6356 6449 6394
rect 6143 6308 6449 6356
rect 6143 6252 6167 6308
rect 6223 6252 6271 6308
rect 6327 6252 6375 6308
rect 6431 6252 6449 6308
rect 6143 6204 6449 6252
rect 15951 6362 15975 6418
rect 16031 6362 16079 6418
rect 16135 6362 16183 6418
rect 16239 6362 16257 6418
rect 15951 6314 16257 6362
rect 15951 6258 15975 6314
rect 16031 6258 16079 6314
rect 16135 6258 16183 6314
rect 16239 6258 16257 6314
rect 15951 6229 16257 6258
rect 6143 6148 6167 6204
rect 6223 6148 6271 6204
rect 6327 6148 6375 6204
rect 6431 6148 6449 6204
rect 6143 6119 6449 6148
rect 28110 795 28394 798
rect 28070 787 28440 795
rect 28070 731 28120 787
rect 28176 731 28224 787
rect 28280 731 28328 787
rect 28384 731 28440 787
rect 28070 683 28440 731
rect 28070 627 28120 683
rect 28176 627 28224 683
rect 28280 627 28328 683
rect 28384 627 28440 683
rect 28070 579 28440 627
rect 28070 523 28120 579
rect 28176 523 28224 579
rect 28280 523 28328 579
rect 28384 523 28440 579
rect 14375 217 14659 227
rect 13977 206 14261 216
rect 13977 150 13987 206
rect 14043 150 14091 206
rect 14147 150 14195 206
rect 14251 150 14261 206
rect 13977 102 14261 150
rect 13977 46 13987 102
rect 14043 46 14091 102
rect 14147 46 14195 102
rect 14251 46 14261 102
rect 13977 -2 14261 46
rect 13977 -58 13987 -2
rect 14043 -58 14091 -2
rect 14147 -58 14195 -2
rect 14251 -58 14261 -2
rect 14375 161 14385 217
rect 14441 161 14489 217
rect 14545 161 14593 217
rect 14649 161 14659 217
rect 14375 113 14659 161
rect 14375 57 14385 113
rect 14441 57 14489 113
rect 14545 57 14593 113
rect 14649 57 14659 113
rect 14375 9 14659 57
rect 14375 -47 14385 9
rect 14441 -47 14489 9
rect 14545 -47 14593 9
rect 14649 -47 14659 9
rect 14375 -57 14659 -47
rect 13977 -68 14261 -58
rect -1048 -500 15407 -427
rect -1048 -556 12133 -500
rect 12189 -556 12237 -500
rect 12293 -556 12341 -500
rect 12397 -528 15407 -500
rect 12397 -547 26491 -528
rect 12397 -556 15098 -547
rect -1048 -603 15098 -556
rect 15154 -603 15202 -547
rect 15258 -603 15306 -547
rect 15362 -603 26491 -547
rect -1048 -604 26491 -603
rect -1048 -660 12133 -604
rect 12189 -660 12237 -604
rect 12293 -660 12341 -604
rect 12397 -651 26491 -604
rect 12397 -660 15098 -651
rect -1048 -707 15098 -660
rect 15154 -707 15202 -651
rect 15258 -707 15306 -651
rect 15362 -707 26491 -651
rect -1048 -708 26491 -707
rect -1048 -764 12133 -708
rect 12189 -764 12237 -708
rect 12293 -764 12341 -708
rect 12397 -755 26491 -708
rect 12397 -764 15098 -755
rect -1048 -811 15098 -764
rect 15154 -811 15202 -755
rect 15258 -811 15306 -755
rect 15362 -811 26491 -755
rect -1048 -833 26491 -811
rect -1048 -858 15407 -833
rect -1780 -1060 18191 -1034
rect -1780 -1079 26012 -1060
rect -1780 -1109 17896 -1079
rect -1780 -1165 9517 -1109
rect 9573 -1165 9621 -1109
rect 9677 -1165 9725 -1109
rect 9781 -1135 17896 -1109
rect 17952 -1135 18000 -1079
rect 18056 -1135 18104 -1079
rect 18160 -1135 26012 -1079
rect 9781 -1165 26012 -1135
rect -1780 -1183 26012 -1165
rect -1780 -1213 17896 -1183
rect -1780 -1269 9517 -1213
rect 9573 -1269 9621 -1213
rect 9677 -1269 9725 -1213
rect 9781 -1239 17896 -1213
rect 17952 -1239 18000 -1183
rect 18056 -1239 18104 -1183
rect 18160 -1239 26012 -1183
rect 9781 -1269 26012 -1239
rect -1780 -1287 26012 -1269
rect -1780 -1317 17896 -1287
rect -1780 -1373 9517 -1317
rect 9573 -1373 9621 -1317
rect 9677 -1373 9725 -1317
rect 9781 -1343 17896 -1317
rect 17952 -1343 18000 -1287
rect 18056 -1343 18104 -1287
rect 18160 -1343 26012 -1287
rect 9781 -1365 26012 -1343
rect 9781 -1373 18191 -1365
rect -1780 -1465 18191 -1373
rect 25767 -1869 26012 -1365
rect 25767 -1921 25800 -1869
rect 25852 -1921 25904 -1869
rect 25956 -1921 26012 -1869
rect 25767 -1973 26012 -1921
rect 25767 -2025 25800 -1973
rect 25852 -2025 25904 -1973
rect 25956 -2025 26012 -1973
rect 25767 -2077 26012 -2025
rect 25767 -2129 25800 -2077
rect 25852 -2129 25904 -2077
rect 25956 -2129 26012 -2077
rect 25767 -2151 26012 -2129
rect 26246 -1870 26491 -833
rect 26246 -1922 26289 -1870
rect 26341 -1922 26393 -1870
rect 26445 -1922 26491 -1870
rect 26246 -1974 26491 -1922
rect 26246 -2026 26289 -1974
rect 26341 -2026 26393 -1974
rect 26445 -2026 26491 -1974
rect 26246 -2078 26491 -2026
rect 26246 -2130 26289 -2078
rect 26341 -2130 26393 -2078
rect 26445 -2130 26491 -2078
rect 26246 -2149 26491 -2130
rect 12111 -2550 12416 -2531
rect 12111 -2561 12133 -2550
rect 7490 -2606 12133 -2561
rect 12189 -2606 12237 -2550
rect 12293 -2606 12341 -2550
rect 12397 -2606 12416 -2550
rect 7490 -2654 12416 -2606
rect 7490 -2710 12133 -2654
rect 12189 -2710 12237 -2654
rect 12293 -2710 12341 -2654
rect 12397 -2710 12416 -2654
rect 7490 -2758 12416 -2710
rect 7490 -2797 12133 -2758
rect 7490 -3363 7726 -2797
rect 12111 -2814 12133 -2797
rect 12189 -2814 12237 -2758
rect 12293 -2814 12341 -2758
rect 12397 -2814 12416 -2758
rect 12111 -2832 12416 -2814
rect 9497 -3008 9802 -2990
rect 7490 -3415 7531 -3363
rect 7583 -3415 7635 -3363
rect 7687 -3415 7726 -3363
rect 7490 -3467 7726 -3415
rect 7490 -3519 7531 -3467
rect 7583 -3519 7635 -3467
rect 7687 -3519 7726 -3467
rect 7490 -3571 7726 -3519
rect 7490 -3623 7531 -3571
rect 7583 -3623 7635 -3571
rect 7687 -3623 7726 -3571
rect 7490 -3657 7726 -3623
rect 7973 -3009 9802 -3008
rect 7973 -3065 9519 -3009
rect 9575 -3065 9623 -3009
rect 9679 -3065 9727 -3009
rect 9783 -3065 9802 -3009
rect 7973 -3113 9802 -3065
rect 7973 -3169 9519 -3113
rect 9575 -3169 9623 -3113
rect 9679 -3169 9727 -3113
rect 9783 -3169 9802 -3113
rect 7973 -3217 9802 -3169
rect 7973 -3244 9519 -3217
rect 7973 -3359 8209 -3244
rect 9497 -3273 9519 -3244
rect 9575 -3273 9623 -3217
rect 9679 -3273 9727 -3217
rect 9783 -3273 9802 -3217
rect 9497 -3291 9802 -3273
rect 7973 -3411 8018 -3359
rect 8070 -3411 8122 -3359
rect 8174 -3411 8209 -3359
rect 7973 -3463 8209 -3411
rect 7973 -3515 8018 -3463
rect 8070 -3515 8122 -3463
rect 8174 -3515 8209 -3463
rect 7973 -3567 8209 -3515
rect 7973 -3619 8018 -3567
rect 8070 -3619 8122 -3567
rect 8174 -3619 8209 -3567
rect 7973 -3676 8209 -3619
rect 9538 -6028 9774 -3291
rect 11694 -5389 11929 -5343
rect 11236 -5503 11929 -5389
rect 9538 -6153 10882 -6028
rect 9538 -6215 9774 -6153
rect -2774 -6395 -2035 -6364
rect -2774 -6451 -2742 -6395
rect -2686 -6451 -2638 -6395
rect -2582 -6451 -2534 -6395
rect -2478 -6398 -2035 -6395
rect -2478 -6451 -2343 -6398
rect -2774 -6454 -2343 -6451
rect -2287 -6454 -2239 -6398
rect -2183 -6454 -2135 -6398
rect -2079 -6454 -2035 -6398
rect -2774 -6499 -2035 -6454
rect -2774 -6555 -2742 -6499
rect -2686 -6555 -2638 -6499
rect -2582 -6555 -2534 -6499
rect -2478 -6502 -2035 -6499
rect -2478 -6555 -2343 -6502
rect -2774 -6558 -2343 -6555
rect -2287 -6558 -2239 -6502
rect -2183 -6558 -2135 -6502
rect -2079 -6558 -2035 -6502
rect -2774 -6603 -2035 -6558
rect -2774 -6659 -2742 -6603
rect -2686 -6659 -2638 -6603
rect -2582 -6659 -2534 -6603
rect -2478 -6606 -2035 -6603
rect -2478 -6659 -2343 -6606
rect -2774 -6662 -2343 -6659
rect -2287 -6662 -2239 -6606
rect -2183 -6662 -2135 -6606
rect -2079 -6662 -2035 -6606
rect -2774 -6697 -2035 -6662
rect 7493 -8191 7729 -8164
rect 7493 -8243 7540 -8191
rect 7592 -8243 7644 -8191
rect 7696 -8243 7729 -8191
rect 7493 -8295 7729 -8243
rect 7493 -8347 7540 -8295
rect 7592 -8347 7644 -8295
rect 7696 -8347 7729 -8295
rect 7493 -8399 7729 -8347
rect 7493 -8451 7540 -8399
rect 7592 -8451 7644 -8399
rect 7696 -8451 7729 -8399
rect 7493 -8857 7729 -8451
rect 7975 -8179 8210 -8159
rect 7975 -8231 8020 -8179
rect 8072 -8231 8124 -8179
rect 8176 -8231 8210 -8179
rect 7975 -8283 8210 -8231
rect 7975 -8335 8020 -8283
rect 8072 -8335 8124 -8283
rect 8176 -8335 8210 -8283
rect 7975 -8387 8210 -8335
rect 7975 -8439 8020 -8387
rect 8072 -8439 8124 -8387
rect 8176 -8439 8210 -8387
rect 7975 -8471 8210 -8439
rect 9944 -8409 10249 -8385
rect 9944 -8465 9967 -8409
rect 10023 -8465 10071 -8409
rect 10127 -8465 10175 -8409
rect 10231 -8465 10249 -8409
rect 9944 -8471 10249 -8465
rect 11694 -8471 11929 -5503
rect 12142 -6028 12378 -2832
rect 14073 -3515 14758 -3476
rect 14073 -3520 14460 -3515
rect 14073 -3576 14128 -3520
rect 14184 -3576 14232 -3520
rect 14288 -3576 14336 -3520
rect 14392 -3571 14460 -3520
rect 14516 -3571 14564 -3515
rect 14620 -3571 14668 -3515
rect 14724 -3571 14758 -3515
rect 14392 -3576 14758 -3571
rect 14073 -3619 14758 -3576
rect 14073 -3624 14460 -3619
rect 14073 -3680 14128 -3624
rect 14184 -3680 14232 -3624
rect 14288 -3680 14336 -3624
rect 14392 -3675 14460 -3624
rect 14516 -3675 14564 -3619
rect 14620 -3675 14668 -3619
rect 14724 -3675 14758 -3619
rect 14392 -3680 14758 -3675
rect 14073 -3723 14758 -3680
rect 14073 -3728 14460 -3723
rect 14073 -3784 14128 -3728
rect 14184 -3784 14232 -3728
rect 14288 -3784 14336 -3728
rect 14392 -3779 14460 -3728
rect 14516 -3779 14564 -3723
rect 14620 -3779 14668 -3723
rect 14724 -3779 14758 -3723
rect 14392 -3784 14758 -3779
rect 14073 -3857 14758 -3784
rect 14425 -3864 14741 -3857
rect 14425 -3920 14462 -3864
rect 14518 -3920 14566 -3864
rect 14622 -3920 14670 -3864
rect 14726 -3920 14741 -3864
rect 14425 -3968 14741 -3920
rect 14425 -4024 14462 -3968
rect 14518 -4024 14566 -3968
rect 14622 -4024 14670 -3968
rect 14726 -4024 14741 -3968
rect 14425 -4072 14741 -4024
rect 14425 -4128 14462 -4072
rect 14518 -4128 14566 -4072
rect 14622 -4128 14670 -4072
rect 14726 -4128 14741 -4072
rect 14425 -4160 14741 -4128
rect 14283 -5389 14519 -5345
rect 17222 -5389 17467 -5372
rect 20085 -5389 20719 -5342
rect 13951 -5503 14519 -5389
rect 16858 -5503 17467 -5389
rect 19765 -5503 20719 -5389
rect 12142 -6153 13273 -6028
rect 12142 -6208 12378 -6153
rect 12213 -6470 12429 -6458
rect 12213 -6540 12226 -6470
rect 12295 -6540 12347 -6470
rect 12416 -6540 12429 -6470
rect 12213 -6552 12429 -6540
rect 7975 -8513 11929 -8471
rect 7975 -8569 9967 -8513
rect 10023 -8569 10071 -8513
rect 10127 -8569 10175 -8513
rect 10231 -8569 11929 -8513
rect 7975 -8617 11929 -8569
rect 7975 -8673 9967 -8617
rect 10023 -8673 10071 -8617
rect 10127 -8673 10175 -8617
rect 10231 -8673 11929 -8617
rect 7975 -8706 11929 -8673
rect 14283 -8857 14519 -5503
rect 15091 -6008 15375 -5995
rect 15091 -6064 15101 -6008
rect 15157 -6064 15205 -6008
rect 15261 -6064 15309 -6008
rect 15365 -6028 15375 -6008
rect 15365 -6064 16199 -6028
rect 15091 -6112 16199 -6064
rect 15091 -6168 15101 -6112
rect 15157 -6168 15205 -6112
rect 15261 -6168 15309 -6112
rect 15365 -6153 16199 -6112
rect 15365 -6168 15375 -6153
rect 15091 -6178 15375 -6168
rect 15210 -6465 15426 -6453
rect 15210 -6535 15223 -6465
rect 15292 -6535 15344 -6465
rect 15413 -6535 15426 -6465
rect 15210 -6547 15426 -6535
rect 7493 -8909 14519 -8857
rect 7493 -8965 9293 -8909
rect 9349 -8965 9397 -8909
rect 9453 -8965 9501 -8909
rect 9557 -8965 14519 -8909
rect 7493 -9013 14519 -8965
rect 7493 -9069 9293 -9013
rect 9349 -9069 9397 -9013
rect 9453 -9069 9501 -9013
rect 9557 -9069 14519 -9013
rect 7493 -9093 14519 -9069
rect 9270 -9117 9575 -9093
rect 9270 -9173 9293 -9117
rect 9349 -9173 9397 -9117
rect 9453 -9173 9501 -9117
rect 9557 -9173 9575 -9117
rect 9270 -9189 9575 -9173
rect 10755 -9432 10992 -9399
rect 10755 -9501 10787 -9432
rect 10857 -9433 10992 -9432
rect 10857 -9501 10912 -9433
rect 10755 -9502 10912 -9501
rect 10982 -9502 10992 -9433
rect 10755 -9553 10992 -9502
rect 10755 -9622 10787 -9553
rect 10857 -9554 10992 -9553
rect 10857 -9622 10912 -9554
rect 10755 -9623 10912 -9622
rect 10982 -9623 10992 -9554
rect 10755 -9651 10992 -9623
rect -4283 -9852 -3983 -9800
rect -3931 -9852 -3879 -9800
rect -3827 -9852 -3775 -9800
rect -3723 -9805 -3269 -9800
rect -3723 -9852 -3617 -9805
rect -4283 -9857 -3617 -9852
rect -3565 -9857 -3513 -9805
rect -3461 -9857 -3409 -9805
rect -3357 -9857 -3269 -9805
rect -4283 -9904 -3269 -9857
rect -4283 -9956 -3983 -9904
rect -3931 -9956 -3879 -9904
rect -3827 -9956 -3775 -9904
rect -3723 -9909 -3269 -9904
rect -3723 -9956 -3617 -9909
rect -4283 -9961 -3617 -9956
rect -3565 -9961 -3513 -9909
rect -3461 -9961 -3409 -9909
rect -3357 -9961 -3269 -9909
rect -4283 -10008 -3269 -9961
rect -4283 -10060 -3983 -10008
rect -3931 -10060 -3879 -10008
rect -3827 -10060 -3775 -10008
rect -3723 -10013 -3269 -10008
rect -3723 -10060 -3617 -10013
rect -4283 -10065 -3617 -10060
rect -3565 -10065 -3513 -10013
rect -3461 -10065 -3409 -10013
rect -3357 -10065 -3269 -10013
rect -4283 -10197 -3269 -10065
rect -4283 -10249 -3977 -10197
rect -3925 -10249 -3873 -10197
rect -3821 -10249 -3769 -10197
rect -3717 -10202 -3269 -10197
rect -3717 -10249 -3611 -10202
rect -4283 -10254 -3611 -10249
rect -3559 -10254 -3507 -10202
rect -3455 -10254 -3403 -10202
rect -3351 -10254 -3269 -10202
rect -4283 -10301 -3269 -10254
rect -4283 -10353 -3977 -10301
rect -3925 -10353 -3873 -10301
rect -3821 -10353 -3769 -10301
rect -3717 -10306 -3269 -10301
rect -3717 -10353 -3611 -10306
rect -4283 -10358 -3611 -10353
rect -3559 -10358 -3507 -10306
rect -3455 -10358 -3403 -10306
rect -3351 -10358 -3269 -10306
rect -4283 -10405 -3269 -10358
rect -4283 -10457 -3977 -10405
rect -3925 -10457 -3873 -10405
rect -3821 -10457 -3769 -10405
rect -3717 -10410 -3269 -10405
rect -3717 -10457 -3611 -10410
rect -4283 -10462 -3611 -10457
rect -3559 -10462 -3507 -10410
rect -3455 -10462 -3403 -10410
rect -3351 -10462 -3269 -10410
rect -4283 -10574 -3269 -10462
rect -4283 -10626 -3985 -10574
rect -3933 -10626 -3881 -10574
rect -3829 -10626 -3777 -10574
rect -3725 -10579 -3269 -10574
rect -3725 -10626 -3619 -10579
rect -4283 -10631 -3619 -10626
rect -3567 -10631 -3515 -10579
rect -3463 -10631 -3411 -10579
rect -3359 -10631 -3269 -10579
rect -4283 -10678 -3269 -10631
rect -4283 -10730 -3985 -10678
rect -3933 -10730 -3881 -10678
rect -3829 -10730 -3777 -10678
rect -3725 -10683 -3269 -10678
rect -3725 -10730 -3619 -10683
rect -4283 -10735 -3619 -10730
rect -3567 -10735 -3515 -10683
rect -3463 -10735 -3411 -10683
rect -3359 -10735 -3269 -10683
rect -4283 -10782 -3269 -10735
rect -4283 -10834 -3985 -10782
rect -3933 -10834 -3881 -10782
rect -3829 -10834 -3777 -10782
rect -3725 -10787 -3269 -10782
rect -3725 -10834 -3619 -10787
rect -4283 -10839 -3619 -10834
rect -3567 -10839 -3515 -10787
rect -3463 -10839 -3411 -10787
rect -3359 -10839 -3269 -10787
rect -4283 -10974 -3269 -10839
rect -4283 -11026 -3961 -10974
rect -3909 -11026 -3857 -10974
rect -3805 -11026 -3753 -10974
rect -3701 -10979 -3269 -10974
rect -3701 -11026 -3595 -10979
rect -4283 -11031 -3595 -11026
rect -3543 -11031 -3491 -10979
rect -3439 -11031 -3387 -10979
rect -3335 -11031 -3269 -10979
rect -4283 -11078 -3269 -11031
rect -4283 -11130 -3961 -11078
rect -3909 -11130 -3857 -11078
rect -3805 -11130 -3753 -11078
rect -3701 -11083 -3269 -11078
rect -3701 -11130 -3595 -11083
rect -4283 -11135 -3595 -11130
rect -3543 -11135 -3491 -11083
rect -3439 -11135 -3387 -11083
rect -3335 -11135 -3269 -11083
rect 17222 -10865 17467 -5503
rect 20085 -5587 20719 -5503
rect 17881 -6007 18165 -5994
rect 17881 -6063 17891 -6007
rect 17947 -6063 17995 -6007
rect 18051 -6063 18099 -6007
rect 18155 -6028 18165 -6007
rect 18155 -6063 18994 -6028
rect 17881 -6111 18994 -6063
rect 17881 -6167 17891 -6111
rect 17947 -6167 17995 -6111
rect 18051 -6167 18099 -6111
rect 18155 -6153 18994 -6111
rect 18155 -6167 18165 -6153
rect 17881 -6177 18165 -6167
rect 17988 -6473 18204 -6461
rect 17988 -6543 18001 -6473
rect 18070 -6543 18122 -6473
rect 18191 -6543 18204 -6473
rect 17988 -6555 18204 -6543
rect 20474 -10470 20719 -5587
rect 28070 -6780 28440 523
rect 28868 387 29152 398
rect 28868 384 28878 387
rect 25630 -6845 28440 -6780
rect 25630 -6897 25741 -6845
rect 25793 -6897 25845 -6845
rect 25897 -6897 25949 -6845
rect 26001 -6897 28440 -6845
rect 25630 -6949 28440 -6897
rect 25630 -7001 25741 -6949
rect 25793 -7001 25845 -6949
rect 25897 -7001 25949 -6949
rect 26001 -7001 28440 -6949
rect 25630 -7053 28440 -7001
rect 25630 -7105 25741 -7053
rect 25793 -7105 25845 -7053
rect 25897 -7105 25949 -7053
rect 26001 -7105 28440 -7053
rect 25630 -7150 28440 -7105
rect 28838 331 28878 384
rect 28934 331 28982 387
rect 29038 331 29086 387
rect 29142 384 29152 387
rect 29142 331 29208 384
rect 28838 283 29208 331
rect 28838 227 28878 283
rect 28934 227 28982 283
rect 29038 227 29086 283
rect 29142 227 29208 283
rect 28838 179 29208 227
rect 28838 123 28878 179
rect 28934 123 28982 179
rect 29038 123 29086 179
rect 29142 123 29208 179
rect 28838 -7390 29208 123
rect 26180 -7455 29208 -7390
rect 26180 -7507 26242 -7455
rect 26294 -7507 26346 -7455
rect 26398 -7507 26450 -7455
rect 26502 -7507 29208 -7455
rect 26180 -7559 29208 -7507
rect 26180 -7611 26242 -7559
rect 26294 -7611 26346 -7559
rect 26398 -7611 26450 -7559
rect 26502 -7611 29208 -7559
rect 26180 -7663 29208 -7611
rect 26180 -7715 26242 -7663
rect 26294 -7715 26346 -7663
rect 26398 -7715 26450 -7663
rect 26502 -7715 29208 -7663
rect 26180 -7760 29208 -7715
rect 21908 -9803 22153 -9773
rect 21908 -9855 21949 -9803
rect 22001 -9855 22053 -9803
rect 22105 -9855 22153 -9803
rect 21908 -9907 22153 -9855
rect 21908 -9959 21949 -9907
rect 22001 -9959 22053 -9907
rect 22105 -9959 22153 -9907
rect 21908 -10011 22153 -9959
rect 21908 -10063 21949 -10011
rect 22001 -10063 22053 -10011
rect 22105 -10063 22153 -10011
rect 21908 -10470 22153 -10063
rect 20474 -10715 22153 -10470
rect 22394 -9789 22639 -9760
rect 22394 -9841 22446 -9789
rect 22498 -9841 22550 -9789
rect 22602 -9841 22639 -9789
rect 22394 -9893 22639 -9841
rect 22394 -9945 22446 -9893
rect 22498 -9945 22550 -9893
rect 22602 -9945 22639 -9893
rect 22394 -9997 22639 -9945
rect 22394 -10049 22446 -9997
rect 22498 -10049 22550 -9997
rect 22602 -10049 22639 -9997
rect 22394 -10865 22639 -10049
rect 17222 -11110 22639 -10865
rect -4283 -11182 -3269 -11135
rect -4283 -11234 -3961 -11182
rect -3909 -11234 -3857 -11182
rect -3805 -11234 -3753 -11182
rect -3701 -11187 -3269 -11182
rect -3701 -11234 -3595 -11187
rect -4283 -11239 -3595 -11234
rect -3543 -11239 -3491 -11187
rect -3439 -11239 -3387 -11187
rect -3335 -11239 -3269 -11187
rect -4283 -11403 -3269 -11239
rect -4283 -11411 -3596 -11403
rect -15663 -11984 11009 -11960
rect -15663 -12040 10799 -11984
rect 10855 -12040 10903 -11984
rect 10959 -12040 11009 -11984
rect -15663 -12088 11009 -12040
rect -15663 -12144 10799 -12088
rect 10855 -12144 10903 -12088
rect 10959 -12144 11009 -12088
rect -15663 -12192 11009 -12144
rect -15663 -12248 10799 -12192
rect 10855 -12248 10903 -12192
rect 10959 -12248 11009 -12192
rect -15663 -12272 11009 -12248
<< via2 >>
rect -1762 14330 -1706 14386
rect -1658 14330 -1602 14386
rect -1554 14330 -1498 14386
rect -1762 14226 -1706 14282
rect -1658 14226 -1602 14282
rect -1554 14226 -1498 14282
rect -1762 14122 -1706 14178
rect -1658 14122 -1602 14178
rect -1554 14122 -1498 14178
rect -14608 12469 -14552 12525
rect -14504 12469 -14448 12525
rect -14400 12469 -14344 12525
rect -14608 12365 -14552 12421
rect -14504 12365 -14448 12421
rect -14400 12365 -14344 12421
rect -14608 12261 -14552 12317
rect -14504 12261 -14448 12317
rect -14400 12261 -14344 12317
rect -9917 11937 -9857 11997
rect -9804 11936 -9744 11996
rect -8890 11926 -8824 12004
rect -8755 11926 -8689 12004
rect -7165 11941 -7105 12001
rect -7051 11941 -6991 12001
rect -8056 9319 -8000 9375
rect -7952 9319 -7896 9375
rect -7848 9319 -7792 9375
rect -7720 9318 -7664 9374
rect -7616 9318 -7560 9374
rect -7512 9318 -7456 9374
rect -8056 9215 -8000 9271
rect -7952 9215 -7896 9271
rect -7848 9215 -7792 9271
rect -7720 9214 -7664 9270
rect -7616 9214 -7560 9270
rect -7512 9214 -7456 9270
rect -8056 9111 -8000 9167
rect -7952 9111 -7896 9167
rect -7848 9111 -7792 9167
rect -7720 9110 -7664 9166
rect -7616 9110 -7560 9166
rect -7512 9110 -7456 9166
rect -8884 8657 -8818 8735
rect -8764 8657 -8698 8735
rect -8884 8527 -8818 8605
rect -8764 8527 -8698 8605
rect -8884 8397 -8818 8475
rect -8764 8397 -8698 8475
rect -4321 6699 -4265 6755
rect -4217 6699 -4161 6755
rect -4113 6699 -4057 6755
rect -3968 6685 -3912 6741
rect -3864 6685 -3808 6741
rect -3760 6685 -3704 6741
rect -3552 6683 -3496 6739
rect -3448 6683 -3392 6739
rect -3344 6683 -3288 6739
rect -4321 6595 -4265 6651
rect -4217 6595 -4161 6651
rect -4113 6595 -4057 6651
rect -3968 6581 -3912 6637
rect -3864 6581 -3808 6637
rect -3760 6581 -3704 6637
rect -3552 6579 -3496 6635
rect -3448 6579 -3392 6635
rect -3344 6579 -3288 6635
rect -4321 6491 -4265 6547
rect -4217 6491 -4161 6547
rect -4113 6491 -4057 6547
rect -3968 6477 -3912 6533
rect -3864 6477 -3808 6533
rect -3760 6477 -3704 6533
rect -3552 6475 -3496 6531
rect -3448 6475 -3392 6531
rect -3344 6475 -3288 6531
rect -4289 6320 -4233 6376
rect -4185 6320 -4129 6376
rect -4048 6318 -3992 6374
rect -3944 6318 -3888 6374
rect -3840 6318 -3784 6374
rect -3645 6318 -3589 6374
rect -3541 6318 -3485 6374
rect -3437 6318 -3381 6374
rect -4289 6216 -4233 6272
rect -4185 6216 -4129 6272
rect -4048 6214 -3992 6270
rect -3944 6214 -3888 6270
rect -3840 6214 -3784 6270
rect -3645 6214 -3589 6270
rect -3541 6214 -3485 6270
rect -3437 6214 -3381 6270
rect -4289 6112 -4233 6168
rect -4185 6112 -4129 6168
rect -4048 6110 -3992 6166
rect -3944 6110 -3888 6166
rect -3840 6110 -3784 6166
rect -3645 6110 -3589 6166
rect -3541 6110 -3485 6166
rect -3437 6110 -3381 6166
rect -4282 5977 -4226 6033
rect -4178 5977 -4122 6033
rect -4041 5975 -3985 6031
rect -3937 5975 -3881 6031
rect -3833 5975 -3777 6031
rect -3638 5975 -3582 6031
rect -3534 5975 -3478 6031
rect -3430 5975 -3374 6031
rect -4289 5842 -4233 5898
rect -4185 5842 -4129 5898
rect -4048 5840 -3992 5896
rect -3944 5840 -3888 5896
rect -3840 5840 -3784 5896
rect -3645 5840 -3589 5896
rect -3541 5840 -3485 5896
rect -3437 5840 -3381 5896
rect -11405 -1859 -11349 -1803
rect -11301 -1859 -11245 -1803
rect -11197 -1859 -11141 -1803
rect -11405 -1963 -11349 -1907
rect -11301 -1963 -11245 -1907
rect -11197 -1963 -11141 -1907
rect -11405 -2067 -11349 -2011
rect -11301 -2067 -11245 -2011
rect -11197 -2067 -11141 -2011
rect -14886 -2506 -14830 -2450
rect -14782 -2506 -14726 -2450
rect -14678 -2506 -14622 -2450
rect -7953 -2509 -7897 -2453
rect -7849 -2509 -7793 -2453
rect -7745 -2509 -7689 -2453
rect -14886 -2610 -14830 -2554
rect -14782 -2610 -14726 -2554
rect -14678 -2610 -14622 -2554
rect -14886 -2714 -14830 -2658
rect -14782 -2714 -14726 -2658
rect -14678 -2714 -14622 -2658
rect -7953 -2613 -7897 -2557
rect -7849 -2613 -7793 -2557
rect -7745 -2613 -7689 -2557
rect -7953 -2717 -7897 -2661
rect -7849 -2717 -7793 -2661
rect -7745 -2717 -7689 -2661
rect -8905 -3056 -8839 -2978
rect -8744 -3054 -8678 -2976
rect -14913 -5646 -14857 -5590
rect -14809 -5646 -14753 -5590
rect -14705 -5646 -14649 -5590
rect -14531 -5644 -14475 -5588
rect -14427 -5644 -14371 -5588
rect -14323 -5644 -14267 -5588
rect -8354 -5652 -8298 -5596
rect -8250 -5652 -8194 -5596
rect -8146 -5652 -8090 -5596
rect -7998 -5657 -7942 -5601
rect -7894 -5657 -7838 -5601
rect -7790 -5657 -7734 -5601
rect -14913 -5750 -14857 -5694
rect -14809 -5750 -14753 -5694
rect -14705 -5750 -14649 -5694
rect -14531 -5748 -14475 -5692
rect -14427 -5748 -14371 -5692
rect -14323 -5748 -14267 -5692
rect -8354 -5756 -8298 -5700
rect -8250 -5756 -8194 -5700
rect -8146 -5756 -8090 -5700
rect -7998 -5761 -7942 -5705
rect -7894 -5761 -7838 -5705
rect -7790 -5761 -7734 -5705
rect -14913 -5854 -14857 -5798
rect -14809 -5854 -14753 -5798
rect -14705 -5854 -14649 -5798
rect -14531 -5852 -14475 -5796
rect -14427 -5852 -14371 -5796
rect -14323 -5852 -14267 -5796
rect -8354 -5860 -8298 -5804
rect -8250 -5860 -8194 -5804
rect -8146 -5860 -8090 -5804
rect -7998 -5865 -7942 -5809
rect -7894 -5865 -7838 -5809
rect -7790 -5865 -7734 -5809
rect -982 13194 -926 13250
rect -878 13194 -822 13250
rect -774 13194 -718 13250
rect -982 13090 -926 13146
rect -878 13090 -822 13146
rect -774 13090 -718 13146
rect -982 12986 -926 13042
rect -878 12986 -822 13042
rect -774 12986 -718 13042
rect 6707 7016 6763 7072
rect 6811 7016 6867 7072
rect 6915 7016 6971 7072
rect 6707 6912 6763 6968
rect 6811 6912 6867 6968
rect 6915 6912 6971 6968
rect 6707 6808 6763 6864
rect 6811 6808 6867 6864
rect 6915 6808 6971 6864
rect 9832 6921 9888 6977
rect 9936 6921 9992 6977
rect 10040 6921 10096 6977
rect 16395 6904 16451 6960
rect 16499 6904 16555 6960
rect 16603 6904 16659 6960
rect 6149 6689 6205 6745
rect 6255 6681 6311 6737
rect 6359 6681 6415 6737
rect 6463 6681 6519 6737
rect 6654 6678 6710 6734
rect 6758 6678 6814 6734
rect 6862 6678 6918 6734
rect 9832 6817 9888 6873
rect 9936 6817 9992 6873
rect 10040 6817 10096 6873
rect 9832 6713 9888 6769
rect 9936 6713 9992 6769
rect 10040 6713 10096 6769
rect 15978 6812 16034 6868
rect 16082 6812 16138 6868
rect 16186 6812 16242 6868
rect 15978 6708 16034 6764
rect 16082 6708 16138 6764
rect 16186 6708 16242 6764
rect 6149 6585 6205 6641
rect 6255 6577 6311 6633
rect 6359 6577 6415 6633
rect 6463 6577 6519 6633
rect 6654 6574 6710 6630
rect 6758 6574 6814 6630
rect 6862 6574 6918 6630
rect 16395 6800 16451 6856
rect 16499 6800 16555 6856
rect 16603 6800 16659 6856
rect 16395 6696 16451 6752
rect 16499 6696 16555 6752
rect 16603 6696 16659 6752
rect 15978 6604 16034 6660
rect 16082 6604 16138 6660
rect 16186 6604 16242 6660
rect 6149 6481 6205 6537
rect 6255 6473 6311 6529
rect 6359 6473 6415 6529
rect 6463 6473 6519 6529
rect 6654 6470 6710 6526
rect 6758 6470 6814 6526
rect 6862 6470 6918 6526
rect 6167 6356 6223 6412
rect 6271 6356 6327 6412
rect 6375 6356 6431 6412
rect 15975 6466 16031 6522
rect 16079 6466 16135 6522
rect 16183 6466 16239 6522
rect 6167 6252 6223 6308
rect 6271 6252 6327 6308
rect 6375 6252 6431 6308
rect 15975 6362 16031 6418
rect 16079 6362 16135 6418
rect 16183 6362 16239 6418
rect 15975 6258 16031 6314
rect 16079 6258 16135 6314
rect 16183 6258 16239 6314
rect 6167 6148 6223 6204
rect 6271 6148 6327 6204
rect 6375 6148 6431 6204
rect 28120 731 28176 787
rect 28224 731 28280 787
rect 28328 731 28384 787
rect 28120 627 28176 683
rect 28224 627 28280 683
rect 28328 627 28384 683
rect 28120 523 28176 579
rect 28224 523 28280 579
rect 28328 523 28384 579
rect 13987 204 14043 206
rect 13987 152 13989 204
rect 13989 152 14041 204
rect 14041 152 14043 204
rect 13987 150 14043 152
rect 14091 204 14147 206
rect 14091 152 14093 204
rect 14093 152 14145 204
rect 14145 152 14147 204
rect 14091 150 14147 152
rect 14195 204 14251 206
rect 14195 152 14197 204
rect 14197 152 14249 204
rect 14249 152 14251 204
rect 14195 150 14251 152
rect 13987 100 14043 102
rect 13987 48 13989 100
rect 13989 48 14041 100
rect 14041 48 14043 100
rect 13987 46 14043 48
rect 14091 100 14147 102
rect 14091 48 14093 100
rect 14093 48 14145 100
rect 14145 48 14147 100
rect 14091 46 14147 48
rect 14195 100 14251 102
rect 14195 48 14197 100
rect 14197 48 14249 100
rect 14249 48 14251 100
rect 14195 46 14251 48
rect 13987 -4 14043 -2
rect 13987 -56 13989 -4
rect 13989 -56 14041 -4
rect 14041 -56 14043 -4
rect 13987 -58 14043 -56
rect 14091 -4 14147 -2
rect 14091 -56 14093 -4
rect 14093 -56 14145 -4
rect 14145 -56 14147 -4
rect 14091 -58 14147 -56
rect 14195 -4 14251 -2
rect 14195 -56 14197 -4
rect 14197 -56 14249 -4
rect 14249 -56 14251 -4
rect 14195 -58 14251 -56
rect 14385 215 14441 217
rect 14385 163 14387 215
rect 14387 163 14439 215
rect 14439 163 14441 215
rect 14385 161 14441 163
rect 14489 215 14545 217
rect 14489 163 14491 215
rect 14491 163 14543 215
rect 14543 163 14545 215
rect 14489 161 14545 163
rect 14593 215 14649 217
rect 14593 163 14595 215
rect 14595 163 14647 215
rect 14647 163 14649 215
rect 14593 161 14649 163
rect 14385 111 14441 113
rect 14385 59 14387 111
rect 14387 59 14439 111
rect 14439 59 14441 111
rect 14385 57 14441 59
rect 14489 111 14545 113
rect 14489 59 14491 111
rect 14491 59 14543 111
rect 14543 59 14545 111
rect 14489 57 14545 59
rect 14593 111 14649 113
rect 14593 59 14595 111
rect 14595 59 14647 111
rect 14647 59 14649 111
rect 14593 57 14649 59
rect 14385 7 14441 9
rect 14385 -45 14387 7
rect 14387 -45 14439 7
rect 14439 -45 14441 7
rect 14385 -47 14441 -45
rect 14489 7 14545 9
rect 14489 -45 14491 7
rect 14491 -45 14543 7
rect 14543 -45 14545 7
rect 14489 -47 14545 -45
rect 14593 7 14649 9
rect 14593 -45 14595 7
rect 14595 -45 14647 7
rect 14647 -45 14649 7
rect 14593 -47 14649 -45
rect 12133 -556 12189 -500
rect 12237 -556 12293 -500
rect 12341 -556 12397 -500
rect 15098 -603 15154 -547
rect 15202 -603 15258 -547
rect 15306 -603 15362 -547
rect 12133 -660 12189 -604
rect 12237 -660 12293 -604
rect 12341 -660 12397 -604
rect 15098 -707 15154 -651
rect 15202 -707 15258 -651
rect 15306 -707 15362 -651
rect 12133 -764 12189 -708
rect 12237 -764 12293 -708
rect 12341 -764 12397 -708
rect 15098 -811 15154 -755
rect 15202 -811 15258 -755
rect 15306 -811 15362 -755
rect 9517 -1165 9573 -1109
rect 9621 -1165 9677 -1109
rect 9725 -1165 9781 -1109
rect 17896 -1135 17952 -1079
rect 18000 -1135 18056 -1079
rect 18104 -1135 18160 -1079
rect 9517 -1269 9573 -1213
rect 9621 -1269 9677 -1213
rect 9725 -1269 9781 -1213
rect 17896 -1239 17952 -1183
rect 18000 -1239 18056 -1183
rect 18104 -1239 18160 -1183
rect 9517 -1373 9573 -1317
rect 9621 -1373 9677 -1317
rect 9725 -1373 9781 -1317
rect 17896 -1343 17952 -1287
rect 18000 -1343 18056 -1287
rect 18104 -1343 18160 -1287
rect 12133 -2606 12189 -2550
rect 12237 -2606 12293 -2550
rect 12341 -2606 12397 -2550
rect 12133 -2710 12189 -2654
rect 12237 -2710 12293 -2654
rect 12341 -2710 12397 -2654
rect 12133 -2814 12189 -2758
rect 12237 -2814 12293 -2758
rect 12341 -2814 12397 -2758
rect 9519 -3065 9575 -3009
rect 9623 -3065 9679 -3009
rect 9727 -3065 9783 -3009
rect 9519 -3169 9575 -3113
rect 9623 -3169 9679 -3113
rect 9727 -3169 9783 -3113
rect 9519 -3273 9575 -3217
rect 9623 -3273 9679 -3217
rect 9727 -3273 9783 -3217
rect -2742 -6451 -2686 -6395
rect -2638 -6451 -2582 -6395
rect -2534 -6451 -2478 -6395
rect -2343 -6454 -2287 -6398
rect -2239 -6454 -2183 -6398
rect -2135 -6454 -2079 -6398
rect -2742 -6555 -2686 -6499
rect -2638 -6555 -2582 -6499
rect -2534 -6555 -2478 -6499
rect -2343 -6558 -2287 -6502
rect -2239 -6558 -2183 -6502
rect -2135 -6558 -2079 -6502
rect -2742 -6659 -2686 -6603
rect -2638 -6659 -2582 -6603
rect -2534 -6659 -2478 -6603
rect -2343 -6662 -2287 -6606
rect -2239 -6662 -2183 -6606
rect -2135 -6662 -2079 -6606
rect 9967 -8465 10023 -8409
rect 10071 -8465 10127 -8409
rect 10175 -8465 10231 -8409
rect 14460 -3517 14516 -3515
rect 14128 -3522 14184 -3520
rect 14128 -3574 14130 -3522
rect 14130 -3574 14182 -3522
rect 14182 -3574 14184 -3522
rect 14128 -3576 14184 -3574
rect 14232 -3522 14288 -3520
rect 14232 -3574 14234 -3522
rect 14234 -3574 14286 -3522
rect 14286 -3574 14288 -3522
rect 14232 -3576 14288 -3574
rect 14336 -3522 14392 -3520
rect 14336 -3574 14338 -3522
rect 14338 -3574 14390 -3522
rect 14390 -3574 14392 -3522
rect 14460 -3569 14462 -3517
rect 14462 -3569 14514 -3517
rect 14514 -3569 14516 -3517
rect 14460 -3571 14516 -3569
rect 14564 -3517 14620 -3515
rect 14564 -3569 14566 -3517
rect 14566 -3569 14618 -3517
rect 14618 -3569 14620 -3517
rect 14564 -3571 14620 -3569
rect 14668 -3517 14724 -3515
rect 14668 -3569 14670 -3517
rect 14670 -3569 14722 -3517
rect 14722 -3569 14724 -3517
rect 14668 -3571 14724 -3569
rect 14336 -3576 14392 -3574
rect 14460 -3621 14516 -3619
rect 14128 -3626 14184 -3624
rect 14128 -3678 14130 -3626
rect 14130 -3678 14182 -3626
rect 14182 -3678 14184 -3626
rect 14128 -3680 14184 -3678
rect 14232 -3626 14288 -3624
rect 14232 -3678 14234 -3626
rect 14234 -3678 14286 -3626
rect 14286 -3678 14288 -3626
rect 14232 -3680 14288 -3678
rect 14336 -3626 14392 -3624
rect 14336 -3678 14338 -3626
rect 14338 -3678 14390 -3626
rect 14390 -3678 14392 -3626
rect 14460 -3673 14462 -3621
rect 14462 -3673 14514 -3621
rect 14514 -3673 14516 -3621
rect 14460 -3675 14516 -3673
rect 14564 -3621 14620 -3619
rect 14564 -3673 14566 -3621
rect 14566 -3673 14618 -3621
rect 14618 -3673 14620 -3621
rect 14564 -3675 14620 -3673
rect 14668 -3621 14724 -3619
rect 14668 -3673 14670 -3621
rect 14670 -3673 14722 -3621
rect 14722 -3673 14724 -3621
rect 14668 -3675 14724 -3673
rect 14336 -3680 14392 -3678
rect 14460 -3725 14516 -3723
rect 14128 -3730 14184 -3728
rect 14128 -3782 14130 -3730
rect 14130 -3782 14182 -3730
rect 14182 -3782 14184 -3730
rect 14128 -3784 14184 -3782
rect 14232 -3730 14288 -3728
rect 14232 -3782 14234 -3730
rect 14234 -3782 14286 -3730
rect 14286 -3782 14288 -3730
rect 14232 -3784 14288 -3782
rect 14336 -3730 14392 -3728
rect 14336 -3782 14338 -3730
rect 14338 -3782 14390 -3730
rect 14390 -3782 14392 -3730
rect 14460 -3777 14462 -3725
rect 14462 -3777 14514 -3725
rect 14514 -3777 14516 -3725
rect 14460 -3779 14516 -3777
rect 14564 -3725 14620 -3723
rect 14564 -3777 14566 -3725
rect 14566 -3777 14618 -3725
rect 14618 -3777 14620 -3725
rect 14564 -3779 14620 -3777
rect 14668 -3725 14724 -3723
rect 14668 -3777 14670 -3725
rect 14670 -3777 14722 -3725
rect 14722 -3777 14724 -3725
rect 14668 -3779 14724 -3777
rect 14336 -3784 14392 -3782
rect 14462 -3866 14518 -3864
rect 14462 -3918 14464 -3866
rect 14464 -3918 14516 -3866
rect 14516 -3918 14518 -3866
rect 14462 -3920 14518 -3918
rect 14566 -3866 14622 -3864
rect 14566 -3918 14568 -3866
rect 14568 -3918 14620 -3866
rect 14620 -3918 14622 -3866
rect 14566 -3920 14622 -3918
rect 14670 -3866 14726 -3864
rect 14670 -3918 14672 -3866
rect 14672 -3918 14724 -3866
rect 14724 -3918 14726 -3866
rect 14670 -3920 14726 -3918
rect 14462 -3970 14518 -3968
rect 14462 -4022 14464 -3970
rect 14464 -4022 14516 -3970
rect 14516 -4022 14518 -3970
rect 14462 -4024 14518 -4022
rect 14566 -3970 14622 -3968
rect 14566 -4022 14568 -3970
rect 14568 -4022 14620 -3970
rect 14620 -4022 14622 -3970
rect 14566 -4024 14622 -4022
rect 14670 -3970 14726 -3968
rect 14670 -4022 14672 -3970
rect 14672 -4022 14724 -3970
rect 14724 -4022 14726 -3970
rect 14670 -4024 14726 -4022
rect 14462 -4074 14518 -4072
rect 14462 -4126 14464 -4074
rect 14464 -4126 14516 -4074
rect 14516 -4126 14518 -4074
rect 14462 -4128 14518 -4126
rect 14566 -4074 14622 -4072
rect 14566 -4126 14568 -4074
rect 14568 -4126 14620 -4074
rect 14620 -4126 14622 -4074
rect 14566 -4128 14622 -4126
rect 14670 -4074 14726 -4072
rect 14670 -4126 14672 -4074
rect 14672 -4126 14724 -4074
rect 14724 -4126 14726 -4074
rect 14670 -4128 14726 -4126
rect 12226 -6540 12295 -6470
rect 12347 -6540 12416 -6470
rect 9967 -8569 10023 -8513
rect 10071 -8569 10127 -8513
rect 10175 -8569 10231 -8513
rect 9967 -8673 10023 -8617
rect 10071 -8673 10127 -8617
rect 10175 -8673 10231 -8617
rect 15101 -6064 15157 -6008
rect 15205 -6064 15261 -6008
rect 15309 -6064 15365 -6008
rect 15101 -6168 15157 -6112
rect 15205 -6168 15261 -6112
rect 15309 -6168 15365 -6112
rect 15223 -6535 15292 -6465
rect 15344 -6535 15413 -6465
rect 9293 -8965 9349 -8909
rect 9397 -8965 9453 -8909
rect 9501 -8965 9557 -8909
rect 9293 -9069 9349 -9013
rect 9397 -9069 9453 -9013
rect 9501 -9069 9557 -9013
rect 9293 -9173 9349 -9117
rect 9397 -9173 9453 -9117
rect 9501 -9173 9557 -9117
rect 10787 -9501 10857 -9432
rect 10912 -9502 10982 -9433
rect 10787 -9622 10857 -9553
rect 10912 -9623 10982 -9554
rect 17891 -6063 17947 -6007
rect 17995 -6063 18051 -6007
rect 18099 -6063 18155 -6007
rect 17891 -6167 17947 -6111
rect 17995 -6167 18051 -6111
rect 18099 -6167 18155 -6111
rect 18001 -6543 18070 -6473
rect 18122 -6543 18191 -6473
rect 28878 331 28934 387
rect 28982 331 29038 387
rect 29086 331 29142 387
rect 28878 227 28934 283
rect 28982 227 29038 283
rect 29086 227 29142 283
rect 28878 123 28934 179
rect 28982 123 29038 179
rect 29086 123 29142 179
rect 10799 -12040 10855 -11984
rect 10903 -12040 10959 -11984
rect 10799 -12144 10855 -12088
rect 10903 -12144 10959 -12088
rect 10799 -12248 10855 -12192
rect 10903 -12248 10959 -12192
<< metal3 >>
rect -35091 15219 -16674 15554
rect -35091 10171 -34756 15219
rect -34529 14729 -17140 15054
rect -34529 10282 -34204 14729
rect -36037 9836 -34205 10171
rect -17465 9418 -17140 14729
rect -17009 12568 -16674 15219
rect -1772 14386 -1488 14396
rect -1772 14330 -1762 14386
rect -1706 14330 -1658 14386
rect -1602 14330 -1554 14386
rect -1498 14349 -1488 14386
rect -1498 14330 3512 14349
rect -1772 14282 3512 14330
rect -1772 14226 -1762 14282
rect -1706 14226 -1658 14282
rect -1602 14226 -1554 14282
rect -1498 14226 3512 14282
rect -1772 14178 3512 14226
rect -1772 14122 -1762 14178
rect -1706 14122 -1658 14178
rect -1602 14122 -1554 14178
rect -1498 14148 3512 14178
rect -1498 14122 -1488 14148
rect -1772 14112 -1488 14122
rect -992 13250 -708 13260
rect -992 13229 -982 13250
rect -1046 13194 -982 13229
rect -926 13194 -878 13250
rect -822 13194 -774 13250
rect -718 13229 -708 13250
rect -718 13194 3240 13229
rect -1046 13146 3240 13194
rect -1046 13090 -982 13146
rect -926 13090 -878 13146
rect -822 13090 -774 13146
rect -718 13090 3240 13146
rect -1046 13042 3240 13090
rect -1046 13011 -982 13042
rect -992 12986 -982 13011
rect -926 12986 -878 13042
rect -822 12986 -774 13042
rect -718 13011 3240 13042
rect -718 12986 -708 13011
rect -992 12976 -708 12986
rect -17009 12525 -14283 12568
rect -17009 12469 -14608 12525
rect -14552 12469 -14504 12525
rect -14448 12469 -14400 12525
rect -14344 12469 -14283 12525
rect -17009 12421 -14283 12469
rect -17009 12365 -14608 12421
rect -14552 12365 -14504 12421
rect -14448 12365 -14400 12421
rect -14344 12365 -14283 12421
rect -17009 12317 -14283 12365
rect -17009 12261 -14608 12317
rect -14552 12261 -14504 12317
rect -14448 12261 -14400 12317
rect -14344 12261 -14283 12317
rect -17009 12233 -14283 12261
rect -9955 12004 -6953 12044
rect -9955 11997 -8890 12004
rect -9955 11937 -9917 11997
rect -9857 11996 -8890 11997
rect -9857 11937 -9804 11996
rect -9955 11936 -9804 11937
rect -9744 11936 -8890 11996
rect -9955 11926 -8890 11936
rect -8824 11926 -8755 12004
rect -8689 12001 -6953 12004
rect -8689 11941 -7165 12001
rect -7105 11941 -7051 12001
rect -6991 11941 -6953 12001
rect -8689 11926 -6953 11941
rect -9955 11902 -6953 11926
rect -19992 9375 -7398 9418
rect -19992 9319 -8056 9375
rect -8000 9319 -7952 9375
rect -7896 9319 -7848 9375
rect -7792 9374 -7398 9375
rect -7792 9319 -7720 9374
rect -19992 9318 -7720 9319
rect -7664 9318 -7616 9374
rect -7560 9318 -7512 9374
rect -7456 9318 -7398 9374
rect -19992 9271 -7398 9318
rect -19992 9215 -8056 9271
rect -8000 9215 -7952 9271
rect -7896 9215 -7848 9271
rect -7792 9270 -7398 9271
rect -7792 9215 -7720 9270
rect -19992 9214 -7720 9215
rect -7664 9214 -7616 9270
rect -7560 9214 -7512 9270
rect -7456 9214 -7398 9270
rect -19992 9167 -7398 9214
rect -19992 9111 -8056 9167
rect -8000 9111 -7952 9167
rect -7896 9111 -7848 9167
rect -7792 9166 -7398 9167
rect -7792 9111 -7720 9166
rect -19992 9110 -7720 9111
rect -7664 9110 -7616 9166
rect -7560 9110 -7512 9166
rect -7456 9110 -7398 9166
rect -19992 9093 -7398 9110
rect -7735 9092 -7431 9093
rect -8927 8735 -8646 8749
rect -8927 8657 -8884 8735
rect -8818 8657 -8764 8735
rect -8698 8657 -8646 8735
rect -8927 8605 -8646 8657
rect -8927 8527 -8884 8605
rect -8818 8527 -8764 8605
rect -8698 8527 -8646 8605
rect -8927 8475 -8646 8527
rect -8927 8397 -8884 8475
rect -8818 8397 -8764 8475
rect -8698 8397 -8646 8475
rect -35369 244 -16952 579
rect -35369 -4804 -35034 244
rect -34807 -246 -17418 79
rect -34807 -4693 -34482 -246
rect -36427 -5139 -34483 -4804
rect -17743 -5557 -17418 -246
rect -17287 -2407 -16952 244
rect -11553 -1803 -11119 -1681
rect -11553 -1859 -11405 -1803
rect -11349 -1859 -11301 -1803
rect -11245 -1859 -11197 -1803
rect -11141 -1859 -11119 -1803
rect -11553 -1907 -11119 -1859
rect -11553 -1963 -11405 -1907
rect -11349 -1963 -11301 -1907
rect -11245 -1963 -11197 -1907
rect -11141 -1963 -11119 -1907
rect -11553 -2011 -11119 -1963
rect -11553 -2067 -11405 -2011
rect -11349 -2067 -11301 -2011
rect -11245 -2067 -11197 -2011
rect -11141 -2067 -11119 -2011
rect -17287 -2450 -14561 -2407
rect -17287 -2506 -14886 -2450
rect -14830 -2506 -14782 -2450
rect -14726 -2506 -14678 -2450
rect -14622 -2506 -14561 -2450
rect -17287 -2554 -14561 -2506
rect -17287 -2610 -14886 -2554
rect -14830 -2610 -14782 -2554
rect -14726 -2610 -14678 -2554
rect -14622 -2610 -14561 -2554
rect -17287 -2658 -14561 -2610
rect -17287 -2714 -14886 -2658
rect -14830 -2714 -14782 -2658
rect -14726 -2714 -14678 -2658
rect -14622 -2714 -14561 -2658
rect -17287 -2742 -14561 -2714
rect -20270 -5562 -14242 -5557
rect -20270 -5588 -14241 -5562
rect -20270 -5590 -14531 -5588
rect -20270 -5646 -14913 -5590
rect -14857 -5646 -14809 -5590
rect -14753 -5646 -14705 -5590
rect -14649 -5644 -14531 -5590
rect -14475 -5644 -14427 -5588
rect -14371 -5644 -14323 -5588
rect -14267 -5644 -14241 -5588
rect -14649 -5646 -14241 -5644
rect -20270 -5692 -14241 -5646
rect -20270 -5694 -14531 -5692
rect -20270 -5750 -14913 -5694
rect -14857 -5750 -14809 -5694
rect -14753 -5750 -14705 -5694
rect -14649 -5748 -14531 -5694
rect -14475 -5748 -14427 -5692
rect -14371 -5748 -14323 -5692
rect -14267 -5748 -14241 -5692
rect -14649 -5750 -14241 -5748
rect -20270 -5796 -14241 -5750
rect -20270 -5798 -14531 -5796
rect -20270 -5854 -14913 -5798
rect -14857 -5854 -14809 -5798
rect -14753 -5854 -14705 -5798
rect -14649 -5852 -14531 -5798
rect -14475 -5852 -14427 -5796
rect -14371 -5852 -14323 -5796
rect -14267 -5852 -14241 -5796
rect -14649 -5854 -14241 -5852
rect -20270 -5874 -14241 -5854
rect -20270 -5882 -14242 -5874
rect -11553 -7077 -11119 -2067
rect -8927 -2976 -8646 8397
rect 6310 7113 6744 7114
rect 6310 7072 16699 7113
rect 6310 7016 6707 7072
rect 6763 7016 6811 7072
rect 6867 7016 6915 7072
rect 6971 7016 16699 7072
rect 6310 6977 16699 7016
rect 6310 6968 9832 6977
rect 6310 6912 6707 6968
rect 6763 6912 6811 6968
rect 6867 6912 6915 6968
rect 6971 6921 9832 6968
rect 9888 6921 9936 6977
rect 9992 6921 10040 6977
rect 10096 6960 16699 6977
rect 10096 6921 16395 6960
rect 6971 6912 16395 6921
rect 6310 6904 16395 6912
rect 16451 6904 16499 6960
rect 16555 6904 16603 6960
rect 16659 6904 16699 6960
rect 6310 6873 16699 6904
rect 6310 6864 9832 6873
rect 6310 6830 6707 6864
rect 6028 6828 6707 6830
rect -4409 6808 6707 6828
rect 6763 6808 6811 6864
rect 6867 6808 6915 6864
rect 6971 6817 9832 6864
rect 9888 6817 9936 6873
rect 9992 6817 10040 6873
rect 10096 6868 16699 6873
rect 10096 6817 15978 6868
rect 6971 6812 15978 6817
rect 16034 6812 16082 6868
rect 16138 6812 16186 6868
rect 16242 6856 16699 6868
rect 16242 6812 16395 6856
rect 6971 6808 16395 6812
rect -4409 6800 16395 6808
rect 16451 6800 16499 6856
rect 16555 6800 16603 6856
rect 16659 6800 16699 6856
rect -4409 6769 16699 6800
rect -4409 6755 9832 6769
rect -4409 6699 -4321 6755
rect -4265 6699 -4217 6755
rect -4161 6699 -4113 6755
rect -4057 6745 9832 6755
rect -4057 6741 6149 6745
rect -4057 6699 -3968 6741
rect -4409 6685 -3968 6699
rect -3912 6685 -3864 6741
rect -3808 6685 -3760 6741
rect -3704 6739 6149 6741
rect -3704 6685 -3552 6739
rect -4409 6683 -3552 6685
rect -3496 6683 -3448 6739
rect -3392 6683 -3344 6739
rect -3288 6689 6149 6739
rect 6205 6737 9832 6745
rect 6205 6689 6255 6737
rect -3288 6683 6255 6689
rect -4409 6681 6255 6683
rect 6311 6681 6359 6737
rect 6415 6681 6463 6737
rect 6519 6734 9832 6737
rect 6519 6681 6654 6734
rect -4409 6678 6654 6681
rect 6710 6678 6758 6734
rect 6814 6678 6862 6734
rect 6918 6713 9832 6734
rect 9888 6713 9936 6769
rect 9992 6713 10040 6769
rect 10096 6764 16699 6769
rect 10096 6713 15978 6764
rect 6918 6708 15978 6713
rect 16034 6708 16082 6764
rect 16138 6708 16186 6764
rect 16242 6752 16699 6764
rect 16242 6708 16395 6752
rect 6918 6696 16395 6708
rect 16451 6696 16499 6752
rect 16555 6696 16603 6752
rect 16659 6696 16699 6752
rect 6918 6678 16699 6696
rect -4409 6660 16699 6678
rect -4409 6651 7022 6660
rect -4409 6595 -4321 6651
rect -4265 6595 -4217 6651
rect -4161 6595 -4113 6651
rect -4057 6641 7022 6651
rect -4057 6637 6149 6641
rect -4057 6595 -3968 6637
rect -4409 6581 -3968 6595
rect -3912 6581 -3864 6637
rect -3808 6581 -3760 6637
rect -3704 6635 6149 6637
rect -3704 6581 -3552 6635
rect -4409 6579 -3552 6581
rect -3496 6579 -3448 6635
rect -3392 6579 -3344 6635
rect -3288 6585 6149 6635
rect 6205 6633 7022 6641
rect 6205 6585 6255 6633
rect -3288 6579 6255 6585
rect -4409 6577 6255 6579
rect 6311 6577 6359 6633
rect 6415 6577 6463 6633
rect 6519 6630 7022 6633
rect 6519 6577 6654 6630
rect -4409 6574 6654 6577
rect 6710 6574 6758 6630
rect 6814 6574 6862 6630
rect 6918 6574 7022 6630
rect -4409 6547 7022 6574
rect -4409 6491 -4321 6547
rect -4265 6491 -4217 6547
rect -4161 6491 -4113 6547
rect -4057 6537 7022 6547
rect -4057 6533 6149 6537
rect -4057 6491 -3968 6533
rect -4409 6477 -3968 6491
rect -3912 6477 -3864 6533
rect -3808 6477 -3760 6533
rect -3704 6531 6149 6533
rect -3704 6477 -3552 6531
rect -4409 6475 -3552 6477
rect -3496 6475 -3448 6531
rect -3392 6475 -3344 6531
rect -3288 6481 6149 6531
rect 6205 6529 7022 6537
rect 6205 6481 6255 6529
rect -3288 6475 6255 6481
rect -4409 6473 6255 6475
rect 6311 6473 6359 6529
rect 6415 6473 6463 6529
rect 6519 6526 7022 6529
rect 6519 6473 6654 6526
rect -4409 6470 6654 6473
rect 6710 6470 6758 6526
rect 6814 6470 6862 6526
rect 6918 6470 7022 6526
rect -4409 6412 7022 6470
rect -4409 6376 6167 6412
rect -4409 6320 -4289 6376
rect -4233 6320 -4185 6376
rect -4129 6374 6167 6376
rect -4129 6320 -4048 6374
rect -4409 6318 -4048 6320
rect -3992 6318 -3944 6374
rect -3888 6318 -3840 6374
rect -3784 6318 -3645 6374
rect -3589 6318 -3541 6374
rect -3485 6318 -3437 6374
rect -3381 6356 6167 6374
rect 6223 6356 6271 6412
rect 6327 6356 6375 6412
rect 6431 6394 7022 6412
rect 15879 6604 15978 6660
rect 16034 6604 16082 6660
rect 16138 6604 16186 6660
rect 16242 6604 16699 6660
rect 15879 6598 16699 6604
rect 15879 6522 16315 6598
rect 15879 6466 15975 6522
rect 16031 6466 16079 6522
rect 16135 6466 16183 6522
rect 16239 6466 16315 6522
rect 15879 6418 16315 6466
rect 6431 6356 7015 6394
rect -3381 6318 7015 6356
rect -4409 6308 7015 6318
rect -4409 6272 6167 6308
rect -4409 6216 -4289 6272
rect -4233 6216 -4185 6272
rect -4129 6270 6167 6272
rect -4129 6216 -4048 6270
rect -4409 6214 -4048 6216
rect -3992 6214 -3944 6270
rect -3888 6214 -3840 6270
rect -3784 6214 -3645 6270
rect -3589 6214 -3541 6270
rect -3485 6214 -3437 6270
rect -3381 6252 6167 6270
rect 6223 6252 6271 6308
rect 6327 6252 6375 6308
rect 6431 6252 7015 6308
rect -3381 6214 7015 6252
rect -4409 6204 7015 6214
rect -4409 6168 6167 6204
rect -4409 6112 -4289 6168
rect -4233 6112 -4185 6168
rect -4129 6166 6167 6168
rect -4129 6112 -4048 6166
rect -4409 6110 -4048 6112
rect -3992 6110 -3944 6166
rect -3888 6110 -3840 6166
rect -3784 6110 -3645 6166
rect -3589 6110 -3541 6166
rect -3485 6110 -3437 6166
rect -3381 6148 6167 6166
rect 6223 6148 6271 6204
rect 6327 6148 6375 6204
rect 6431 6148 7015 6204
rect 15879 6362 15975 6418
rect 16031 6362 16079 6418
rect 16135 6362 16183 6418
rect 16239 6362 16315 6418
rect 15879 6314 16315 6362
rect 15879 6258 15975 6314
rect 16031 6258 16079 6314
rect 16135 6258 16183 6314
rect 16239 6258 16315 6314
rect 15879 6170 16315 6258
rect -3381 6110 7015 6148
rect -4409 6041 7015 6110
rect -4409 6033 -3235 6041
rect -4409 5977 -4282 6033
rect -4226 5977 -4178 6033
rect -4122 6031 -3235 6033
rect -4122 5977 -4041 6031
rect -4409 5975 -4041 5977
rect -3985 5975 -3937 6031
rect -3881 5975 -3833 6031
rect -3777 5975 -3638 6031
rect -3582 5975 -3534 6031
rect -3478 5975 -3430 6031
rect -3374 5975 -3235 6031
rect -4409 5898 -3235 5975
rect -4409 5842 -4289 5898
rect -4233 5842 -4185 5898
rect -4129 5896 -3235 5898
rect -4129 5842 -4048 5896
rect -4409 5840 -4048 5842
rect -3992 5840 -3944 5896
rect -3888 5840 -3840 5896
rect -3784 5840 -3645 5896
rect -3589 5840 -3541 5896
rect -3485 5840 -3437 5896
rect -3381 5840 -3235 5896
rect -4409 5760 -3235 5840
rect 28110 787 28394 797
rect 28110 731 28120 787
rect 28176 731 28224 787
rect 28280 731 28328 787
rect 28384 731 28394 787
rect 28110 683 28394 731
rect 28110 627 28120 683
rect 28176 627 28224 683
rect 28280 627 28328 683
rect 28384 627 28394 683
rect 28110 579 28394 627
rect 28110 523 28120 579
rect 28176 523 28224 579
rect 28280 523 28328 579
rect 28384 523 28394 579
rect 28110 513 28394 523
rect 28868 387 29152 397
rect 28868 331 28878 387
rect 28934 331 28982 387
rect 29038 331 29086 387
rect 29142 331 29152 387
rect 28868 283 29152 331
rect 13962 217 14794 271
rect 13962 206 14385 217
rect 13962 150 13987 206
rect 14043 150 14091 206
rect 14147 150 14195 206
rect 14251 161 14385 206
rect 14441 161 14489 217
rect 14545 161 14593 217
rect 14649 161 14794 217
rect 14251 150 14794 161
rect 13962 113 14794 150
rect 28868 227 28878 283
rect 28934 227 28982 283
rect 29038 227 29086 283
rect 29142 227 29152 283
rect 28868 179 29152 227
rect 28868 123 28878 179
rect 28934 123 28982 179
rect 29038 123 29086 179
rect 29142 123 29152 179
rect 28868 113 29152 123
rect 13962 102 14385 113
rect 13962 46 13987 102
rect 14043 46 14091 102
rect 14147 46 14195 102
rect 14251 57 14385 102
rect 14441 57 14489 113
rect 14545 57 14593 113
rect 14649 57 14794 113
rect 14251 46 14794 57
rect 13962 9 14794 46
rect 13962 -2 14385 9
rect 13962 -58 13987 -2
rect 14043 -58 14091 -2
rect 14147 -58 14195 -2
rect 14251 -47 14385 -2
rect 14441 -47 14489 9
rect 14545 -47 14593 9
rect 14649 -47 14794 9
rect 14251 -58 14794 -47
rect 13962 -151 14794 -58
rect 12111 -500 12416 -433
rect 12111 -556 12133 -500
rect 12189 -556 12237 -500
rect 12293 -556 12341 -500
rect 12397 -556 12416 -500
rect 12111 -604 12416 -556
rect 12111 -660 12133 -604
rect 12189 -660 12237 -604
rect 12293 -660 12341 -604
rect 12397 -660 12416 -604
rect 12111 -708 12416 -660
rect 12111 -764 12133 -708
rect 12189 -764 12237 -708
rect 12293 -764 12341 -708
rect 12397 -764 12416 -708
rect 9497 -1090 9802 -1053
rect 9495 -1109 9802 -1090
rect 9495 -1165 9517 -1109
rect 9573 -1165 9621 -1109
rect 9677 -1165 9725 -1109
rect 9781 -1165 9802 -1109
rect 9495 -1213 9802 -1165
rect 9495 -1269 9517 -1213
rect 9573 -1269 9621 -1213
rect 9677 -1269 9725 -1213
rect 9781 -1269 9802 -1213
rect 9495 -1317 9802 -1269
rect 9495 -1373 9517 -1317
rect 9573 -1373 9621 -1317
rect 9677 -1373 9725 -1317
rect 9781 -1373 9802 -1317
rect 9495 -1391 9802 -1373
rect -8927 -2978 -8744 -2976
rect -8927 -3056 -8905 -2978
rect -8839 -3054 -8744 -2978
rect -8678 -3054 -8646 -2976
rect -8839 -3056 -8646 -3054
rect -8927 -3065 -8646 -3056
rect -7968 -2453 -7644 -2431
rect -7968 -2509 -7953 -2453
rect -7897 -2509 -7849 -2453
rect -7793 -2509 -7745 -2453
rect -7689 -2509 -7644 -2453
rect -7968 -2557 -7644 -2509
rect -7968 -2613 -7953 -2557
rect -7897 -2613 -7849 -2557
rect -7793 -2613 -7745 -2557
rect -7689 -2613 -7644 -2557
rect -7968 -2661 -7644 -2613
rect -7968 -2717 -7953 -2661
rect -7897 -2717 -7849 -2661
rect -7793 -2717 -7745 -2661
rect -7689 -2717 -7644 -2661
rect -7968 -5545 -7643 -2717
rect 9497 -3009 9802 -1391
rect 12111 -2550 12416 -764
rect 12111 -2606 12133 -2550
rect 12189 -2606 12237 -2550
rect 12293 -2606 12341 -2550
rect 12397 -2606 12416 -2550
rect 12111 -2654 12416 -2606
rect 12111 -2710 12133 -2654
rect 12189 -2710 12237 -2654
rect 12293 -2710 12341 -2654
rect 12397 -2710 12416 -2654
rect 12111 -2758 12416 -2710
rect 12111 -2814 12133 -2758
rect 12189 -2814 12237 -2758
rect 12293 -2814 12341 -2758
rect 12397 -2814 12416 -2758
rect 12111 -2832 12416 -2814
rect 9497 -3065 9519 -3009
rect 9575 -3065 9623 -3009
rect 9679 -3065 9727 -3009
rect 9783 -3065 9802 -3009
rect 9497 -3113 9802 -3065
rect 9497 -3169 9519 -3113
rect 9575 -3169 9623 -3113
rect 9679 -3169 9727 -3113
rect 9783 -3169 9802 -3113
rect 9497 -3217 9802 -3169
rect 9497 -3273 9519 -3217
rect 9575 -3273 9623 -3217
rect 9679 -3273 9727 -3217
rect 9783 -3273 9802 -3217
rect 9497 -3291 9802 -3273
rect 14036 -3515 14794 -151
rect 14036 -3520 14460 -3515
rect 14036 -3576 14128 -3520
rect 14184 -3576 14232 -3520
rect 14288 -3576 14336 -3520
rect 14392 -3571 14460 -3520
rect 14516 -3571 14564 -3515
rect 14620 -3571 14668 -3515
rect 14724 -3571 14794 -3515
rect 14392 -3576 14794 -3571
rect 14036 -3619 14794 -3576
rect 14036 -3624 14460 -3619
rect 14036 -3680 14128 -3624
rect 14184 -3680 14232 -3624
rect 14288 -3680 14336 -3624
rect 14392 -3675 14460 -3624
rect 14516 -3675 14564 -3619
rect 14620 -3675 14668 -3619
rect 14724 -3675 14794 -3619
rect 14392 -3680 14794 -3675
rect 14036 -3723 14794 -3680
rect 14036 -3728 14460 -3723
rect 14036 -3784 14128 -3728
rect 14184 -3784 14232 -3728
rect 14288 -3784 14336 -3728
rect 14392 -3779 14460 -3728
rect 14516 -3779 14564 -3723
rect 14620 -3779 14668 -3723
rect 14724 -3779 14794 -3723
rect 14392 -3784 14794 -3779
rect 14036 -3864 14794 -3784
rect 14036 -3920 14462 -3864
rect 14518 -3920 14566 -3864
rect 14622 -3920 14670 -3864
rect 14726 -3920 14794 -3864
rect 14036 -3968 14794 -3920
rect 14036 -3989 14462 -3968
rect 14372 -3993 14462 -3989
rect 14425 -4024 14462 -3993
rect 14518 -4024 14566 -3968
rect 14622 -4024 14670 -3968
rect 14726 -3993 14794 -3968
rect 15076 -547 15381 -528
rect 15076 -603 15098 -547
rect 15154 -603 15202 -547
rect 15258 -603 15306 -547
rect 15362 -603 15381 -547
rect 15076 -651 15381 -603
rect 15076 -707 15098 -651
rect 15154 -707 15202 -651
rect 15258 -707 15306 -651
rect 15362 -707 15381 -651
rect 15076 -755 15381 -707
rect 15076 -811 15098 -755
rect 15154 -811 15202 -755
rect 15258 -811 15306 -755
rect 15362 -811 15381 -755
rect 14726 -4024 14741 -3993
rect 14425 -4072 14741 -4024
rect 14425 -4128 14462 -4072
rect 14518 -4128 14566 -4072
rect 14622 -4128 14670 -4072
rect 14726 -4128 14741 -4072
rect 14425 -4160 14741 -4128
rect -8384 -5596 -7623 -5545
rect -8384 -5652 -8354 -5596
rect -8298 -5652 -8250 -5596
rect -8194 -5652 -8146 -5596
rect -8090 -5601 -7623 -5596
rect -8090 -5652 -7998 -5601
rect -8384 -5657 -7998 -5652
rect -7942 -5657 -7894 -5601
rect -7838 -5657 -7790 -5601
rect -7734 -5657 -7623 -5601
rect -8384 -5700 -7623 -5657
rect -8384 -5756 -8354 -5700
rect -8298 -5756 -8250 -5700
rect -8194 -5756 -8146 -5700
rect -8090 -5705 -7623 -5700
rect -8090 -5756 -7998 -5705
rect -8384 -5761 -7998 -5756
rect -7942 -5761 -7894 -5705
rect -7838 -5761 -7790 -5705
rect -7734 -5761 -7623 -5705
rect -8384 -5804 -7623 -5761
rect -8384 -5860 -8354 -5804
rect -8298 -5860 -8250 -5804
rect -8194 -5860 -8146 -5804
rect -8090 -5809 -7623 -5804
rect -8090 -5860 -7998 -5809
rect -8384 -5865 -7998 -5860
rect -7942 -5865 -7894 -5809
rect -7838 -5865 -7790 -5809
rect -7734 -5865 -7623 -5809
rect -8384 -5892 -7623 -5865
rect 15076 -6008 15381 -811
rect 17876 -1065 18179 -1060
rect 15076 -6064 15101 -6008
rect 15157 -6064 15205 -6008
rect 15261 -6064 15309 -6008
rect 15365 -6064 15381 -6008
rect 15076 -6112 15381 -6064
rect 15076 -6168 15101 -6112
rect 15157 -6168 15205 -6112
rect 15261 -6168 15309 -6112
rect 15365 -6168 15381 -6112
rect 15076 -6217 15381 -6168
rect 17875 -1079 18179 -1065
rect 17875 -1135 17896 -1079
rect 17952 -1135 18000 -1079
rect 18056 -1135 18104 -1079
rect 18160 -1135 18179 -1079
rect 17875 -1183 18179 -1135
rect 17875 -1239 17896 -1183
rect 17952 -1239 18000 -1183
rect 18056 -1239 18104 -1183
rect 18160 -1239 18179 -1183
rect 17875 -1287 18179 -1239
rect 17875 -1343 17896 -1287
rect 17952 -1343 18000 -1287
rect 18056 -1343 18104 -1287
rect 18160 -1343 18179 -1287
rect 17875 -1365 18179 -1343
rect 17875 -6007 18168 -1365
rect 17875 -6063 17891 -6007
rect 17947 -6063 17995 -6007
rect 18051 -6063 18099 -6007
rect 18155 -6063 18168 -6007
rect 17875 -6111 18168 -6063
rect 17875 -6167 17891 -6111
rect 17947 -6167 17995 -6111
rect 18051 -6167 18099 -6111
rect 18155 -6167 18168 -6111
rect 17875 -6184 18168 -6167
rect -2787 -6395 -643 -6283
rect -2787 -6451 -2742 -6395
rect -2686 -6451 -2638 -6395
rect -2582 -6451 -2534 -6395
rect -2478 -6398 -643 -6395
rect -2478 -6451 -2343 -6398
rect -2787 -6454 -2343 -6451
rect -2287 -6454 -2239 -6398
rect -2183 -6454 -2135 -6398
rect -2079 -6454 -643 -6398
rect -2787 -6499 -643 -6454
rect -2787 -6555 -2742 -6499
rect -2686 -6555 -2638 -6499
rect -2582 -6555 -2534 -6499
rect -2478 -6502 -643 -6499
rect -2478 -6555 -2343 -6502
rect -2787 -6558 -2343 -6555
rect -2287 -6558 -2239 -6502
rect -2183 -6558 -2135 -6502
rect -2079 -6558 -643 -6502
rect 12213 -6470 12429 -6458
rect 12213 -6540 12226 -6470
rect 12295 -6540 12347 -6470
rect 12416 -6540 12429 -6470
rect 12213 -6552 12429 -6540
rect 15210 -6465 15426 -6453
rect 15210 -6535 15223 -6465
rect 15292 -6535 15344 -6465
rect 15413 -6535 15426 -6465
rect 15210 -6547 15426 -6535
rect 17988 -6473 18204 -6461
rect 17988 -6543 18001 -6473
rect 18070 -6543 18122 -6473
rect 18191 -6543 18204 -6473
rect -2787 -6603 -643 -6558
rect -2787 -6659 -2742 -6603
rect -2686 -6659 -2638 -6603
rect -2582 -6659 -2534 -6603
rect -2478 -6606 -643 -6603
rect -2478 -6659 -2343 -6606
rect -2787 -6662 -2343 -6659
rect -2287 -6662 -2239 -6606
rect -2183 -6662 -2135 -6606
rect -2079 -6662 -643 -6606
rect -2787 -6717 -643 -6662
rect -11553 -7511 -1558 -7077
rect -1992 -10404 -1558 -7511
rect -1077 -9644 -643 -6717
rect 9912 -8409 10346 -8353
rect 9912 -8465 9967 -8409
rect 10023 -8465 10071 -8409
rect 10127 -8465 10175 -8409
rect 10231 -8465 10346 -8409
rect 9912 -8513 10346 -8465
rect 9912 -8569 9967 -8513
rect 10023 -8569 10071 -8513
rect 10127 -8569 10175 -8513
rect 10231 -8569 10346 -8513
rect 9912 -8617 10346 -8569
rect 9912 -8673 9967 -8617
rect 10023 -8673 10071 -8617
rect 10127 -8673 10175 -8617
rect 10231 -8673 10346 -8617
rect 9194 -8909 9628 -8838
rect 9194 -8965 9293 -8909
rect 9349 -8965 9397 -8909
rect 9453 -8965 9501 -8909
rect 9557 -8965 9628 -8909
rect 9194 -9013 9628 -8965
rect 9194 -9069 9293 -9013
rect 9349 -9069 9397 -9013
rect 9453 -9069 9501 -9013
rect 9557 -9069 9628 -9013
rect 9194 -9117 9628 -9069
rect 9194 -9173 9293 -9117
rect 9349 -9173 9397 -9117
rect 9453 -9173 9501 -9117
rect 9557 -9173 9628 -9117
rect 9194 -9644 9628 -9173
rect -1077 -10078 9628 -9644
rect 9912 -10404 10346 -8673
rect -1992 -10838 10346 -10404
rect 10731 -9432 11013 -9379
rect 10731 -9501 10787 -9432
rect 10857 -9433 11013 -9432
rect 10857 -9501 10912 -9433
rect 10731 -9502 10912 -9501
rect 10982 -9502 11013 -9433
rect 10731 -9526 11013 -9502
rect 12269 -9526 12378 -6552
rect 15266 -9526 15375 -6547
rect 17988 -6555 18204 -6543
rect 18036 -9526 18145 -6555
rect 10731 -9553 18145 -9526
rect 10731 -9622 10787 -9553
rect 10857 -9554 18145 -9553
rect 10857 -9622 10912 -9554
rect 10731 -9623 10912 -9622
rect 10982 -9623 18145 -9554
rect 10731 -9635 18145 -9623
rect 10731 -11984 11013 -9635
rect 10731 -12040 10799 -11984
rect 10855 -12040 10903 -11984
rect 10959 -12040 11013 -11984
rect 10731 -12088 11013 -12040
rect 10731 -12144 10799 -12088
rect 10855 -12144 10903 -12088
rect 10959 -12144 11013 -12088
rect 10731 -12192 11013 -12144
rect 10731 -12248 10799 -12192
rect 10855 -12248 10903 -12192
rect 10959 -12248 11013 -12192
rect 10731 -14224 11013 -12248
use fold_cascode_opamp_mag  fold_cascode_opamp_mag_0 ~/GF180Projects/Tapeout/Magic/Folded_single
timestamp 1699423855
transform 1 0 -30797 0 1 -2114
box -4063 -11248 17072 1731
use fold_cascode_opamp_mag  fold_cascode_opamp_mag_1
timestamp 1699423855
transform 1 0 -30519 0 1 12861
box -4063 -11248 17072 1731
use Folded_Diff_Op_Amp_Layout  Folded_Diff_Op_Amp_Layout_0 ~/GF180Projects/Tapeout/Magic/Op_Amp
timestamp 1699898304
transform 1 0 486 0 1 9157
box -486 -9157 66932 6239
use nfet_03v3_DNLN9V  nfet_03v3_DNLN9V_0
timestamp 1699541970
transform 1 0 -10708 0 1 -3680
box -140 -579 140 579
use pfet_03v3_9DZW5M  pfet_03v3_9DZW5M_0
timestamp 1699541970
transform 1 0 -10708 0 1 -2035
box -202 -1016 202 1016
use ppolyf_u_RKAYB7  ppolyf_u_RKAYB7_0
timestamp 1699111554
transform 1 0 24200 0 -1 -5724
box -3024 -1086 3024 1086
use ppolyf_u_RKAYB7  ppolyf_u_RKAYB7_1
timestamp 1699111554
transform 1 0 24200 0 1 -3174
box -3024 -1086 3024 1086
use ppolyf_u_RKAYB7  ppolyf_u_RKAYB7_2
timestamp 1699111554
transform 1 0 5930 0 -1 -7154
box -3024 -1086 3024 1086
use ppolyf_u_RKAYB7  ppolyf_u_RKAYB7_3
timestamp 1699111554
transform 1 0 24200 0 1 -8768
box -3024 -1086 3024 1086
use ppolyf_u_RKAYB7  ppolyf_u_RKAYB7_4
timestamp 1699111554
transform 1 0 5930 0 1 -4604
box -3024 -1086 3024 1086
use Transmission_Gate_Layout  Transmission_Gate_Layout_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/Transmission_Gate1
timestamp 1699271742
transform 1 0 10185 0 1 -7735
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_1
timestamp 1699271742
transform 1 0 18585 0 1 -7735
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_2
timestamp 1699271742
transform 1 0 12785 0 1 -7735
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_3
timestamp 1699271742
transform 1 0 15785 0 1 -7735
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_4
timestamp 1699271742
transform 1 0 -7031 0 1 -4234
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_5
timestamp 1699271742
transform 1 0 -13771 0 1 -4251
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_6
timestamp 1699271742
transform 1 0 -9765 0 1 -4237
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_7
timestamp 1699271742
transform 1 0 -6753 0 1 10741
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_8
timestamp 1699271742
transform 1 0 -13493 0 1 10724
box -350 -272 1471 3508
use Transmission_Gate_Layout  Transmission_Gate_Layout_9
timestamp 1699271742
transform 1 0 -9487 0 1 10738
box -350 -272 1471 3508
<< labels >>
flabel metal3 -8788 3390 -8788 3390 0 FreeSans 1600 0 0 0 SELB
port 0 nsew
flabel metal3 10895 -14040 10895 -14040 0 FreeSans 1600 0 0 0 SEL
port 1 nsew
flabel metal3 -35757 10008 -35757 10008 0 FreeSans 1600 0 0 0 VINP
port 2 nsew
flabel metal3 -36089 -4961 -36089 -4961 0 FreeSans 1600 0 0 0 VINN
port 3 nsew
flabel metal2 31360 15026 31360 15026 0 FreeSans 1600 0 0 0 OUTP
port 4 nsew
flabel metal2 32267 14476 32267 14476 0 FreeSans 1600 0 0 0 OUTN
port 5 nsew
flabel metal1 -4305 14455 -4305 14455 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
<< end >>
