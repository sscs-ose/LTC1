magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2169 -2045 2169 2045
<< psubdiff >>
rect -169 23 169 45
rect -169 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 169 23
rect -169 -45 169 -23
<< psubdiffcont >>
rect -147 -23 -101 23
rect -23 -23 23 23
rect 101 -23 147 23
<< metal1 >>
rect -158 23 158 34
rect -158 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 158 23
rect -158 -34 158 -23
<< end >>
