magic
tech gf180mcuC
magscale 1 10
timestamp 1693997255
<< pwell >>
rect -516 -804 516 804
<< nmos >>
rect -404 336 -204 736
rect -100 336 100 736
rect 204 336 404 736
rect -404 -200 -204 200
rect -100 -200 100 200
rect 204 -200 404 200
rect -404 -736 -204 -336
rect -100 -736 100 -336
rect 204 -736 404 -336
<< ndiff >>
rect -492 723 -404 736
rect -492 349 -479 723
rect -433 349 -404 723
rect -492 336 -404 349
rect -204 723 -100 736
rect -204 349 -175 723
rect -129 349 -100 723
rect -204 336 -100 349
rect 100 723 204 736
rect 100 349 129 723
rect 175 349 204 723
rect 100 336 204 349
rect 404 723 492 736
rect 404 349 433 723
rect 479 349 492 723
rect 404 336 492 349
rect -492 187 -404 200
rect -492 -187 -479 187
rect -433 -187 -404 187
rect -492 -200 -404 -187
rect -204 187 -100 200
rect -204 -187 -175 187
rect -129 -187 -100 187
rect -204 -200 -100 -187
rect 100 187 204 200
rect 100 -187 129 187
rect 175 -187 204 187
rect 100 -200 204 -187
rect 404 187 492 200
rect 404 -187 433 187
rect 479 -187 492 187
rect 404 -200 492 -187
rect -492 -349 -404 -336
rect -492 -723 -479 -349
rect -433 -723 -404 -349
rect -492 -736 -404 -723
rect -204 -349 -100 -336
rect -204 -723 -175 -349
rect -129 -723 -100 -349
rect -204 -736 -100 -723
rect 100 -349 204 -336
rect 100 -723 129 -349
rect 175 -723 204 -349
rect 100 -736 204 -723
rect 404 -349 492 -336
rect 404 -723 433 -349
rect 479 -723 492 -349
rect 404 -736 492 -723
<< ndiffc >>
rect -479 349 -433 723
rect -175 349 -129 723
rect 129 349 175 723
rect 433 349 479 723
rect -479 -187 -433 187
rect -175 -187 -129 187
rect 129 -187 175 187
rect 433 -187 479 187
rect -479 -723 -433 -349
rect -175 -723 -129 -349
rect 129 -723 175 -349
rect 433 -723 479 -349
<< polysilicon >>
rect -404 736 -204 780
rect -100 736 100 780
rect 204 736 404 780
rect -404 292 -204 336
rect -100 292 100 336
rect 204 292 404 336
rect -404 200 -204 244
rect -100 200 100 244
rect 204 200 404 244
rect -404 -244 -204 -200
rect -100 -244 100 -200
rect 204 -244 404 -200
rect -404 -336 -204 -292
rect -100 -336 100 -292
rect 204 -336 404 -292
rect -404 -780 -204 -736
rect -100 -780 100 -736
rect 204 -780 404 -736
<< metal1 >>
rect -479 723 -433 734
rect -479 338 -433 349
rect -175 723 -129 734
rect -175 338 -129 349
rect 129 723 175 734
rect 129 338 175 349
rect 433 723 479 734
rect 433 338 479 349
rect -479 187 -433 198
rect -479 -198 -433 -187
rect -175 187 -129 198
rect -175 -198 -129 -187
rect 129 187 175 198
rect 129 -198 175 -187
rect 433 187 479 198
rect 433 -198 479 -187
rect -479 -349 -433 -338
rect -479 -734 -433 -723
rect -175 -349 -129 -338
rect -175 -734 -129 -723
rect 129 -349 175 -338
rect 129 -734 175 -723
rect 433 -349 479 -338
rect 433 -734 479 -723
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 2 l 1 m 3 nf 3 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
