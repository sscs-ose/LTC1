magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1409 1045 1409
<< metal2 >>
rect -45 404 45 409
rect -45 -404 -40 404
rect 40 -404 45 404
rect -45 -409 45 -404
<< via2 >>
rect -40 -404 40 404
<< metal3 >>
rect -45 404 45 409
rect -45 -404 -40 404
rect 40 -404 45 404
rect -45 -409 45 -404
<< end >>
