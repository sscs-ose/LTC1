magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1331 1045 1331
<< metal2 >>
rect -45 326 45 331
rect -45 -326 -40 326
rect 40 -326 45 326
rect -45 -331 45 -326
<< via2 >>
rect -40 -326 40 326
<< metal3 >>
rect -45 326 45 331
rect -45 -326 -40 326
rect 40 -326 45 326
rect -45 -331 45 -326
<< end >>
