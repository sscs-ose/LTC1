magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2468 -2118 2468 2118
<< pwell >>
rect -468 -118 468 118
<< nmos >>
rect -356 -50 -256 50
rect -152 -50 -52 50
rect 52 -50 152 50
rect 256 -50 356 50
<< ndiff >>
rect -444 23 -356 50
rect -444 -23 -431 23
rect -385 -23 -356 23
rect -444 -50 -356 -23
rect -256 23 -152 50
rect -256 -23 -227 23
rect -181 -23 -152 23
rect -256 -50 -152 -23
rect -52 23 52 50
rect -52 -23 -23 23
rect 23 -23 52 23
rect -52 -50 52 -23
rect 152 23 256 50
rect 152 -23 181 23
rect 227 -23 256 23
rect 152 -50 256 -23
rect 356 23 444 50
rect 356 -23 385 23
rect 431 -23 444 23
rect 356 -50 444 -23
<< ndiffc >>
rect -431 -23 -385 23
rect -227 -23 -181 23
rect -23 -23 23 23
rect 181 -23 227 23
rect 385 -23 431 23
<< polysilicon >>
rect -356 50 -256 94
rect -152 50 -52 94
rect 52 50 152 94
rect 256 50 356 94
rect -356 -94 -256 -50
rect -152 -94 -52 -50
rect 52 -94 152 -50
rect 256 -94 356 -50
<< metal1 >>
rect -431 23 -385 48
rect -431 -48 -385 -23
rect -227 23 -181 48
rect -227 -48 -181 -23
rect -23 23 23 48
rect -23 -48 23 -23
rect 181 23 227 48
rect 181 -48 227 -23
rect 385 23 431 48
rect 385 -48 431 -23
<< end >>
