magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2195 -2995 2195 2995
<< ndiff >>
rect -195 973 195 995
rect -195 -973 -173 973
rect 173 -973 195 973
rect -195 -995 195 -973
<< ndiffc >>
rect -173 -973 173 973
<< metal1 >>
rect -184 973 184 984
rect -184 -973 -173 973
rect 173 -973 184 973
rect -184 -984 184 -973
<< end >>
