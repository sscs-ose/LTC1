magic
tech gf180mcuC
magscale 1 10
timestamp 1693226830
<< error_p >>
rect -2455 -58 -2409 58
rect -2151 -58 -2105 58
rect -1847 -58 -1801 58
rect -1543 -58 -1497 58
rect -1239 -58 -1193 58
rect -935 -58 -889 58
rect -631 -58 -585 58
rect -327 -58 -281 58
rect -23 -58 23 58
rect 281 -58 327 58
rect 585 -58 631 58
rect 889 -58 935 58
rect 1193 -58 1239 58
rect 1497 -58 1543 58
rect 1801 -58 1847 58
rect 2105 -58 2151 58
rect 2409 -58 2455 58
<< pwell >>
rect -2492 -128 2492 128
<< nmos >>
rect -2380 -60 -2180 60
rect -2076 -60 -1876 60
rect -1772 -60 -1572 60
rect -1468 -60 -1268 60
rect -1164 -60 -964 60
rect -860 -60 -660 60
rect -556 -60 -356 60
rect -252 -60 -52 60
rect 52 -60 252 60
rect 356 -60 556 60
rect 660 -60 860 60
rect 964 -60 1164 60
rect 1268 -60 1468 60
rect 1572 -60 1772 60
rect 1876 -60 2076 60
rect 2180 -60 2380 60
<< ndiff >>
rect -2468 47 -2380 60
rect -2468 -47 -2455 47
rect -2409 -47 -2380 47
rect -2468 -60 -2380 -47
rect -2180 47 -2076 60
rect -2180 -47 -2151 47
rect -2105 -47 -2076 47
rect -2180 -60 -2076 -47
rect -1876 47 -1772 60
rect -1876 -47 -1847 47
rect -1801 -47 -1772 47
rect -1876 -60 -1772 -47
rect -1572 47 -1468 60
rect -1572 -47 -1543 47
rect -1497 -47 -1468 47
rect -1572 -60 -1468 -47
rect -1268 47 -1164 60
rect -1268 -47 -1239 47
rect -1193 -47 -1164 47
rect -1268 -60 -1164 -47
rect -964 47 -860 60
rect -964 -47 -935 47
rect -889 -47 -860 47
rect -964 -60 -860 -47
rect -660 47 -556 60
rect -660 -47 -631 47
rect -585 -47 -556 47
rect -660 -60 -556 -47
rect -356 47 -252 60
rect -356 -47 -327 47
rect -281 -47 -252 47
rect -356 -60 -252 -47
rect -52 47 52 60
rect -52 -47 -23 47
rect 23 -47 52 47
rect -52 -60 52 -47
rect 252 47 356 60
rect 252 -47 281 47
rect 327 -47 356 47
rect 252 -60 356 -47
rect 556 47 660 60
rect 556 -47 585 47
rect 631 -47 660 47
rect 556 -60 660 -47
rect 860 47 964 60
rect 860 -47 889 47
rect 935 -47 964 47
rect 860 -60 964 -47
rect 1164 47 1268 60
rect 1164 -47 1193 47
rect 1239 -47 1268 47
rect 1164 -60 1268 -47
rect 1468 47 1572 60
rect 1468 -47 1497 47
rect 1543 -47 1572 47
rect 1468 -60 1572 -47
rect 1772 47 1876 60
rect 1772 -47 1801 47
rect 1847 -47 1876 47
rect 1772 -60 1876 -47
rect 2076 47 2180 60
rect 2076 -47 2105 47
rect 2151 -47 2180 47
rect 2076 -60 2180 -47
rect 2380 47 2468 60
rect 2380 -47 2409 47
rect 2455 -47 2468 47
rect 2380 -60 2468 -47
<< ndiffc >>
rect -2455 -47 -2409 47
rect -2151 -47 -2105 47
rect -1847 -47 -1801 47
rect -1543 -47 -1497 47
rect -1239 -47 -1193 47
rect -935 -47 -889 47
rect -631 -47 -585 47
rect -327 -47 -281 47
rect -23 -47 23 47
rect 281 -47 327 47
rect 585 -47 631 47
rect 889 -47 935 47
rect 1193 -47 1239 47
rect 1497 -47 1543 47
rect 1801 -47 1847 47
rect 2105 -47 2151 47
rect 2409 -47 2455 47
<< polysilicon >>
rect -2380 60 -2180 104
rect -2076 60 -1876 104
rect -1772 60 -1572 104
rect -1468 60 -1268 104
rect -1164 60 -964 104
rect -860 60 -660 104
rect -556 60 -356 104
rect -252 60 -52 104
rect 52 60 252 104
rect 356 60 556 104
rect 660 60 860 104
rect 964 60 1164 104
rect 1268 60 1468 104
rect 1572 60 1772 104
rect 1876 60 2076 104
rect 2180 60 2380 104
rect -2380 -104 -2180 -60
rect -2076 -104 -1876 -60
rect -1772 -104 -1572 -60
rect -1468 -104 -1268 -60
rect -1164 -104 -964 -60
rect -860 -104 -660 -60
rect -556 -104 -356 -60
rect -252 -104 -52 -60
rect 52 -104 252 -60
rect 356 -104 556 -60
rect 660 -104 860 -60
rect 964 -104 1164 -60
rect 1268 -104 1468 -60
rect 1572 -104 1772 -60
rect 1876 -104 2076 -60
rect 2180 -104 2380 -60
<< metal1 >>
rect -2455 47 -2409 58
rect -2455 -58 -2409 -47
rect -2151 47 -2105 58
rect -2151 -58 -2105 -47
rect -1847 47 -1801 58
rect -1847 -58 -1801 -47
rect -1543 47 -1497 58
rect -1543 -58 -1497 -47
rect -1239 47 -1193 58
rect -1239 -58 -1193 -47
rect -935 47 -889 58
rect -935 -58 -889 -47
rect -631 47 -585 58
rect -631 -58 -585 -47
rect -327 47 -281 58
rect -327 -58 -281 -47
rect -23 47 23 58
rect -23 -58 23 -47
rect 281 47 327 58
rect 281 -58 327 -47
rect 585 47 631 58
rect 585 -58 631 -47
rect 889 47 935 58
rect 889 -58 935 -47
rect 1193 47 1239 58
rect 1193 -58 1239 -47
rect 1497 47 1543 58
rect 1497 -58 1543 -47
rect 1801 47 1847 58
rect 1801 -58 1847 -47
rect 2105 47 2151 58
rect 2105 -58 2151 -47
rect 2409 47 2455 58
rect 2409 -58 2455 -47
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.6 l 1 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 0 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
