magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2400 -2000 15200 15065
<< metal2 >>
rect -400 12400 13200 13065
rect -400 400 400 12400
rect 668 400 1008 12400
rect 1068 400 1408 12400
rect 1468 400 1808 12400
rect 1868 400 2208 12400
rect 2268 400 2608 12400
rect 2668 400 3008 12400
rect 3068 400 3408 12400
rect 3468 400 3808 12400
rect 3868 400 4208 12400
rect 4268 400 4608 12400
rect 4668 400 5008 12400
rect 5068 400 5408 12400
rect 5468 400 5808 12400
rect 5868 400 6208 12400
rect 6268 400 6608 12400
rect 6668 400 7008 12400
rect 7068 400 7408 12400
rect 7468 400 7808 12400
rect 7868 400 8208 12400
rect 8268 400 8608 12400
rect 8668 400 9008 12400
rect 9068 400 9408 12400
rect 9468 400 9808 12400
rect 9868 400 10208 12400
rect 10268 400 10608 12400
rect 10668 400 11008 12400
rect 11068 400 11408 12400
rect 11468 400 11808 12400
rect 11868 400 12208 12400
rect 12400 400 13200 12400
rect -400 0 13200 400
<< metal3 >>
rect -400 12320 13200 13065
rect -400 458 400 12320
rect 668 458 1008 12320
rect 1068 458 1408 12320
rect 1468 458 1808 12320
rect 1868 458 2208 12320
rect 2268 458 2608 12320
rect 2668 458 3008 12320
rect 3068 458 3408 12320
rect 3468 458 3808 12320
rect 3868 458 4208 12320
rect 4268 458 4608 12320
rect 4668 458 5008 12320
rect 5068 458 5408 12320
rect 5468 458 5808 12320
rect 5868 458 6208 12320
rect 6268 458 6608 12320
rect 6668 458 7008 12320
rect 7068 458 7408 12320
rect 7468 458 7808 12320
rect 7868 458 8208 12320
rect 8268 458 8608 12320
rect 8668 458 9008 12320
rect 9068 458 9408 12320
rect 9468 458 9808 12320
rect 9868 458 10208 12320
rect 10268 458 10608 12320
rect 10668 458 11008 12320
rect 11068 458 11408 12320
rect 11468 458 11808 12320
rect 11868 458 12208 12320
rect 12400 458 13200 12320
rect -400 0 13200 458
<< metal4 >>
rect -400 12320 13200 13065
rect -400 458 400 12320
rect 668 458 1008 12320
rect 1068 458 1408 12320
rect 1468 458 1808 12320
rect 1868 458 2208 12320
rect 2268 458 2608 12320
rect 2668 458 3008 12320
rect 3068 458 3408 12320
rect 3468 458 3808 12320
rect 3868 458 4208 12320
rect 4268 458 4608 12320
rect 4668 458 5008 12320
rect 5068 458 5408 12320
rect 5468 458 5808 12320
rect 5868 458 6208 12320
rect 6268 458 6608 12320
rect 6668 458 7008 12320
rect 7068 458 7408 12320
rect 7468 458 7808 12320
rect 7868 458 8208 12320
rect 8268 458 8608 12320
rect 8668 458 9008 12320
rect 9068 458 9408 12320
rect 9468 458 9808 12320
rect 9868 458 10208 12320
rect 10268 458 10608 12320
rect 10668 458 11008 12320
rect 11068 458 11408 12320
rect 11468 458 11808 12320
rect 11868 458 12208 12320
rect 12400 458 13200 12320
rect -400 0 13200 458
<< metal5 >>
rect -400 0 13200 13065
<< glass >>
rect 400 400 12400 12400
use M3_M2_CDNS_6903358316516  M3_M2_CDNS_6903358316516_0
timestamp 1713338890
transform 0 -1 -10 1 0 6254
box -6114 -286 6114 286
use M3_M2_CDNS_6903358316516  M3_M2_CDNS_6903358316516_1
timestamp 1713338890
transform 0 -1 12802 1 0 6254
box -6114 -286 6114 286
use M3_M2_CDNS_6903358316517  M3_M2_CDNS_6903358316517_0
timestamp 1713338890
transform 1 0 6408 0 1 12735
box -6672 -224 6672 224
use M3_M2_CDNS_6903358316518  M3_M2_CDNS_6903358316518_0
timestamp 1713338890
transform 1 0 6407 0 1 203
box -6002 -109 6002 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_0
timestamp 1713338890
transform 0 -1 840 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_1
timestamp 1713338890
transform 0 -1 1241 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_2
timestamp 1713338890
transform 0 -1 2038 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_3
timestamp 1713338890
transform 0 -1 1641 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_4
timestamp 1713338890
transform 0 -1 2435 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_5
timestamp 1713338890
transform 0 -1 3235 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_6
timestamp 1713338890
transform 0 -1 2839 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_7
timestamp 1713338890
transform 0 -1 3635 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_8
timestamp 1713338890
transform 0 -1 4032 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_9
timestamp 1713338890
transform 0 -1 4437 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_10
timestamp 1713338890
transform 0 -1 4837 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_11
timestamp 1713338890
transform 0 -1 5242 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_12
timestamp 1713338890
transform 0 -1 5639 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_13
timestamp 1713338890
transform 0 -1 6036 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_14
timestamp 1713338890
transform 0 -1 6439 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_15
timestamp 1713338890
transform 0 -1 6841 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_16
timestamp 1713338890
transform 0 -1 7638 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_17
timestamp 1713338890
transform 0 -1 7244 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_18
timestamp 1713338890
transform 0 -1 8039 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_19
timestamp 1713338890
transform 0 -1 8836 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_20
timestamp 1713338890
transform 0 -1 8439 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_21
timestamp 1713338890
transform 0 -1 9233 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_22
timestamp 1713338890
transform 0 -1 9637 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_23
timestamp 1713338890
transform 0 -1 10033 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_24
timestamp 1713338890
transform 0 -1 10433 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_25
timestamp 1713338890
transform 0 -1 10830 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_26
timestamp 1713338890
transform 0 -1 11235 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_27
timestamp 1713338890
transform 0 -1 11635 1 0 6389
box -5931 -109 5931 109
use M3_M2_CDNS_6903358316519  M3_M2_CDNS_6903358316519_28
timestamp 1713338890
transform 0 -1 12040 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316512  M4_M3_CDNS_6903358316512_0
timestamp 1713338890
transform 1 0 6408 0 1 12735
box -6672 -224 6672 224
use M4_M3_CDNS_6903358316513  M4_M3_CDNS_6903358316513_0
timestamp 1713338890
transform 0 -1 -10 1 0 6254
box -6114 -286 6114 286
use M4_M3_CDNS_6903358316513  M4_M3_CDNS_6903358316513_1
timestamp 1713338890
transform 0 -1 12802 1 0 6254
box -6114 -286 6114 286
use M4_M3_CDNS_6903358316514  M4_M3_CDNS_6903358316514_0
timestamp 1713338890
transform 1 0 6407 0 1 203
box -6002 -109 6002 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_0
timestamp 1713338890
transform 0 -1 840 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_1
timestamp 1713338890
transform 0 -1 1241 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_2
timestamp 1713338890
transform 0 -1 2038 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_3
timestamp 1713338890
transform 0 -1 1641 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_4
timestamp 1713338890
transform 0 -1 2435 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_5
timestamp 1713338890
transform 0 -1 2839 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_6
timestamp 1713338890
transform 0 -1 3235 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_7
timestamp 1713338890
transform 0 -1 3635 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_8
timestamp 1713338890
transform 0 -1 4032 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_9
timestamp 1713338890
transform 0 -1 4437 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_10
timestamp 1713338890
transform 0 -1 4837 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_11
timestamp 1713338890
transform 0 -1 5242 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_12
timestamp 1713338890
transform 0 -1 5639 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_13
timestamp 1713338890
transform 0 -1 6036 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_14
timestamp 1713338890
transform 0 -1 6439 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_15
timestamp 1713338890
transform 0 -1 6841 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_16
timestamp 1713338890
transform 0 -1 7244 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_17
timestamp 1713338890
transform 0 -1 7638 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_18
timestamp 1713338890
transform 0 -1 8039 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_19
timestamp 1713338890
transform 0 -1 8439 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_20
timestamp 1713338890
transform 0 -1 8836 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_21
timestamp 1713338890
transform 0 -1 9233 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_22
timestamp 1713338890
transform 0 -1 9637 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_23
timestamp 1713338890
transform 0 -1 10033 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_24
timestamp 1713338890
transform 0 -1 10433 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_25
timestamp 1713338890
transform 0 -1 10830 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_26
timestamp 1713338890
transform 0 -1 11635 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_27
timestamp 1713338890
transform 0 -1 11235 1 0 6389
box -5931 -109 5931 109
use M4_M3_CDNS_6903358316515  M4_M3_CDNS_6903358316515_28
timestamp 1713338890
transform 0 -1 12040 1 0 6389
box -5931 -109 5931 109
use M5_M4_CDNS_690335831658  M5_M4_CDNS_690335831658_0
timestamp 1713338890
transform 1 0 6408 0 1 12735
box -6678 -230 6678 230
use M5_M4_CDNS_690335831659  M5_M4_CDNS_690335831659_0
timestamp 1713338890
transform 0 -1 -10 1 0 6254
box -6120 -292 6120 292
use M5_M4_CDNS_690335831659  M5_M4_CDNS_690335831659_1
timestamp 1713338890
transform 0 -1 12802 1 0 6254
box -6120 -292 6120 292
use M5_M4_CDNS_6903358316510  M5_M4_CDNS_6903358316510_0
timestamp 1713338890
transform 1 0 6407 0 1 203
box -6008 -115 6008 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_0
timestamp 1713338890
transform 0 -1 840 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_1
timestamp 1713338890
transform 0 -1 1241 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_2
timestamp 1713338890
transform 0 -1 2038 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_3
timestamp 1713338890
transform 0 -1 1641 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_4
timestamp 1713338890
transform 0 -1 2435 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_5
timestamp 1713338890
transform 0 -1 3235 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_6
timestamp 1713338890
transform 0 -1 2839 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_7
timestamp 1713338890
transform 0 -1 3635 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_8
timestamp 1713338890
transform 0 -1 4437 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_9
timestamp 1713338890
transform 0 -1 4032 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_10
timestamp 1713338890
transform 0 -1 4837 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_11
timestamp 1713338890
transform 0 -1 5639 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_12
timestamp 1713338890
transform 0 -1 5242 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_13
timestamp 1713338890
transform 0 -1 6036 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_14
timestamp 1713338890
transform 0 -1 6439 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_15
timestamp 1713338890
transform 0 -1 6841 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_16
timestamp 1713338890
transform 0 -1 7638 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_17
timestamp 1713338890
transform 0 -1 7244 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_18
timestamp 1713338890
transform 0 -1 8039 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_19
timestamp 1713338890
transform 0 -1 8836 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_20
timestamp 1713338890
transform 0 -1 8439 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_21
timestamp 1713338890
transform 0 -1 9233 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_22
timestamp 1713338890
transform 0 -1 9637 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_23
timestamp 1713338890
transform 0 -1 10433 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_24
timestamp 1713338890
transform 0 -1 10033 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_25
timestamp 1713338890
transform 0 -1 10830 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_26
timestamp 1713338890
transform 0 -1 11635 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_27
timestamp 1713338890
transform 0 -1 11235 1 0 6389
box -5937 -115 5937 115
use M5_M4_CDNS_6903358316511  M5_M4_CDNS_6903358316511_28
timestamp 1713338890
transform 0 -1 12040 1 0 6389
box -5937 -115 5937 115
<< end >>
