magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1409 1019 1409
<< metal2 >>
rect -19 404 19 409
rect -19 -404 -14 404
rect 14 -404 19 404
rect -19 -409 19 -404
<< via2 >>
rect -14 -404 14 404
<< metal3 >>
rect -19 404 19 409
rect -19 -404 -14 404
rect 14 -404 19 404
rect -19 -409 19 -404
<< end >>
