magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -4113 -2045 4113 2045
<< ndiff >>
rect -2113 23 2113 45
rect -2113 -23 -2091 23
rect 2091 -23 2113 23
rect -2113 -45 2113 -23
<< ndiffc >>
rect -2091 -23 2091 23
<< metal1 >>
rect -2102 23 2102 34
rect -2102 -23 -2091 23
rect 2091 -23 2102 23
rect -2102 -34 2102 -23
<< end >>
