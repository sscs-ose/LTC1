magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7204 -2128 7204 2128
<< nwell >>
rect -5204 -128 5204 128
<< nsubdiff >>
rect -5121 23 5121 45
rect -5121 -23 -5099 23
rect 5099 -23 5121 23
rect -5121 -45 5121 -23
<< nsubdiffcont >>
rect -5099 -23 5099 23
<< metal1 >>
rect -5110 23 5110 34
rect -5110 -23 -5099 23
rect 5099 -23 5110 23
rect -5110 -34 5110 -23
<< end >>
