magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 17032 71968
<< metal5 >>
rect 0 68400 15000 69678
rect 0 66800 15000 68200
rect 0 65200 15000 66600
rect 0 63600 15000 65000
rect 0 62000 15000 63400
rect 0 60400 15000 61800
rect 0 58800 15000 60200
rect 0 57200 15000 58600
rect 0 55600 15000 57000
rect 937 55400 3937 55600
rect 4337 55400 7337 55600
rect 7737 55400 10737 55600
rect 11137 55400 14137 55600
rect 0 54000 15000 55400
rect 937 53800 3937 54000
rect 4337 53800 7337 54000
rect 7737 53800 10737 54000
rect 11137 53800 14137 54000
rect 0 52400 15000 53800
rect 0 50800 15000 52200
rect 0 49200 15000 50600
rect 0 46000 15000 49000
rect 0 42800 15000 45800
rect 937 42600 3937 42800
rect 4337 42600 7337 42800
rect 7737 42600 10737 42800
rect 11137 42600 14137 42800
rect 0 41200 15000 42600
rect 0 39600 15000 41000
rect 0 36400 15000 39400
rect 937 36200 3937 36400
rect 4337 36200 7337 36400
rect 7737 36200 10737 36400
rect 11137 36200 14137 36400
rect 0 33200 15000 36200
rect 937 33000 3937 33200
rect 4337 33000 7337 33200
rect 7737 33000 10737 33200
rect 11137 33000 14137 33200
rect 0 30000 15000 33000
rect 937 29800 3937 30000
rect 4337 29800 7337 30000
rect 7737 29800 10737 30000
rect 11137 29800 14137 30000
rect 0 26800 15000 29800
rect 0 25200 15000 26600
rect 0 23600 15000 25000
rect 0 20400 15000 23400
rect 937 20200 3937 20400
rect 4337 20200 7337 20400
rect 7737 20200 10737 20400
rect 11137 20200 14137 20400
rect 0 17200 15000 20200
rect 937 17000 3937 17200
rect 4337 17000 7337 17200
rect 7737 17000 10737 17200
rect 11137 17000 14137 17200
rect 0 14000 15000 17000
use 4LM_METAL_RAIL  4LM_METAL_RAIL_0
timestamp 1713338890
transform 1 0 0 0 1 0
box -32 13097 15032 69968
use M4_M3_CDNS_690335831653  M4_M3_CDNS_690335831653_0
timestamp 1713338890
transform 1 0 7502 0 1 24296
box -7351 -677 7351 677
use M4_M3_CDNS_690335831653  M4_M3_CDNS_690335831653_1
timestamp 1713338890
transform 1 0 7502 0 1 41896
box -7351 -677 7351 677
use M4_M3_CDNS_690335831653  M4_M3_CDNS_690335831653_2
timestamp 1713338890
transform 1 0 7502 0 1 51496
box -7351 -677 7351 677
use M4_M3_CDNS_690335831653  M4_M3_CDNS_690335831653_3
timestamp 1713338890
transform 1 0 7502 0 1 54696
box -7351 -677 7351 677
use M4_M3_CDNS_690335831653  M4_M3_CDNS_690335831653_4
timestamp 1713338890
transform 1 0 7502 0 1 57896
box -7351 -677 7351 677
use M4_M3_CDNS_690335831653  M4_M3_CDNS_690335831653_5
timestamp 1713338890
transform 1 0 7502 0 1 61096
box -7351 -677 7351 677
use M4_M3_CDNS_690335831653  M4_M3_CDNS_690335831653_6
timestamp 1713338890
transform 1 0 7502 0 1 64296
box -7351 -677 7351 677
use M4_M3_CDNS_690335831653  M4_M3_CDNS_690335831653_7
timestamp 1713338890
transform 1 0 7502 0 1 67504
box -7351 -677 7351 677
use M4_M3_CDNS_690335831654  M4_M3_CDNS_690335831654_0
timestamp 1713338890
transform 1 0 7502 0 1 18693
box -7351 -1458 7351 1458
use M4_M3_CDNS_690335831654  M4_M3_CDNS_690335831654_1
timestamp 1713338890
transform 1 0 7502 0 1 31493
box -7351 -1458 7351 1458
use M4_M3_CDNS_690335831654  M4_M3_CDNS_690335831654_2
timestamp 1713338890
transform 1 0 7502 0 1 37894
box -7351 -1458 7351 1458
use M4_M3_CDNS_690335831654  M4_M3_CDNS_690335831654_3
timestamp 1713338890
transform 1 0 7502 0 1 47493
box -7351 -1458 7351 1458
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_0
timestamp 1713338890
transform 1 0 7502 0 1 15493
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_1
timestamp 1713338890
transform 1 0 7502 0 1 18693
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_2
timestamp 1713338890
transform 1 0 7502 0 1 21893
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_3
timestamp 1713338890
transform 1 0 7502 0 1 28293
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_4
timestamp 1713338890
transform 1 0 7502 0 1 31493
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_5
timestamp 1713338890
transform 1 0 7502 0 1 34694
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_6
timestamp 1713338890
transform 1 0 7502 0 1 37894
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_7
timestamp 1713338890
transform 1 0 7502 0 1 44293
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831650  M5_M4_CDNS_690335831650_8
timestamp 1713338890
transform 1 0 7502 0 1 47493
box -7357 -1464 7357 1464
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_0
timestamp 1713338890
transform 1 0 7502 0 1 24296
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_1
timestamp 1713338890
transform 1 0 7502 0 1 25896
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_2
timestamp 1713338890
transform 1 0 7502 0 1 41896
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_3
timestamp 1713338890
transform 1 0 7502 0 1 40296
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_4
timestamp 1713338890
transform 1 0 7502 0 1 49896
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_5
timestamp 1713338890
transform 1 0 7502 0 1 51496
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_6
timestamp 1713338890
transform 1 0 7502 0 1 53104
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_7
timestamp 1713338890
transform 1 0 7502 0 1 54696
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_8
timestamp 1713338890
transform 1 0 7502 0 1 56304
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_9
timestamp 1713338890
transform 1 0 7502 0 1 57896
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_10
timestamp 1713338890
transform 1 0 7502 0 1 59504
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_11
timestamp 1713338890
transform 1 0 7502 0 1 61096
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_12
timestamp 1713338890
transform 1 0 7502 0 1 62704
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_13
timestamp 1713338890
transform 1 0 7502 0 1 64296
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_14
timestamp 1713338890
transform 1 0 7502 0 1 67504
box -7357 -683 7357 683
use M5_M4_CDNS_690335831651  M5_M4_CDNS_690335831651_15
timestamp 1713338890
transform 1 0 7502 0 1 65904
box -7357 -683 7357 683
use M5_M4_CDNS_690335831652  M5_M4_CDNS_690335831652_0
timestamp 1713338890
transform 1 0 7502 0 1 69041
box -7357 -612 7357 612
<< labels >>
rlabel metal5 s 753 67369 753 67369 4 DVDD
port 1 nsew
rlabel metal5 s 753 59534 753 59534 4 DVDD
port 1 nsew
rlabel metal5 s 753 56334 753 56334 4 DVDD
port 1 nsew
rlabel metal5 s 753 54569 753 54569 4 DVDD
port 1 nsew
rlabel metal5 s 753 53134 753 53134 4 DVDD
port 1 nsew
rlabel metal5 s 753 44279 753 44279 4 DVDD
port 1 nsew
rlabel metal5 s 753 41888 753 41888 4 DVDD
port 1 nsew
rlabel metal5 s 753 37870 753 37870 4 DVDD
port 1 nsew
rlabel metal5 s 753 34634 753 34634 4 DVDD
port 1 nsew
rlabel metal5 s 753 31520 753 31520 4 DVDD
port 1 nsew
rlabel metal5 s 753 28305 753 28305 4 DVDD
port 1 nsew
rlabel metal5 s 753 24195 753 24195 4 DVDD
port 1 nsew
rlabel metal5 s 684 18832 684 18832 4 DVSS
port 2 nsew
rlabel metal5 s 731 15661 731 15661 4 DVSS
port 2 nsew
rlabel metal5 s 753 68960 753 68960 4 DVSS
port 2 nsew
rlabel metal5 s 753 65934 753 65934 4 DVSS
port 2 nsew
rlabel metal5 s 753 60969 753 60969 4 DVSS
port 2 nsew
rlabel metal5 s 753 57769 753 57769 4 DVSS
port 2 nsew
rlabel metal5 s 753 47506 753 47506 4 DVSS
port 2 nsew
rlabel metal5 s 753 40253 753 40253 4 DVSS
port 2 nsew
rlabel metal5 s 753 26011 753 26011 4 DVSS
port 2 nsew
rlabel metal5 s 753 21818 753 21818 4 DVSS
port 2 nsew
rlabel metal5 s 753 62734 753 62734 4 VDD
port 3 nsew
rlabel metal5 s 753 51369 753 51369 4 VDD
port 3 nsew
rlabel metal5 s 753 64169 753 64169 4 VSS
port 4 nsew
rlabel metal5 s 753 49934 753 49934 4 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 13097 15000 70000
<< end >>
