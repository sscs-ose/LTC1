* NGSPICE file created from OR_flat.ext - technology: gf180mcuC

.subckt OR_flat A B VSS VDD OUT
X0 a_230_424# A.t0 Inverter_0.IN VDD.t8 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 Inverter_0.IN A.t1 VSS.t5 VSS.t4 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X2 Inverter_0.IN B.t0 VSS.t3 VSS.t2 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X3 VDD B.t1 a_230_424# VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 OUT Inverter_0.IN VSS.t1 VSS.t0 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X5 OUT Inverter_0.IN VDD.t4 VDD.t3 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X6 Inverter_0.IN A.t2 a_230_424# VDD.t7 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X7 a_230_424# B.t2 VDD.t6 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 A.t2 A.t0 44.4957
R1 A.n0 A.t1 27.2239
R2 A.n0 A.t2 15.0244
R3 A A.n0 5.30993
R4 VDD.t8 VDD.n2 826.923
R5 VDD.n3 VDD.t7 448.719
R6 VDD.n3 VDD.t0 414.531
R7 VDD.t7 VDD.t8 341.88
R8 VDD.t0 VDD.t5 341.88
R9 VDD.n2 VDD.t3 36.3253
R10 VDD.n7 VDD.t6 6.90119
R11 VDD.n7 VDD.n6 6.61028
R12 VDD.n0 VDD.t4 6.40636
R13 VDD.n2 VDD 6.3005
R14 VDD.n5 VDD.n4 3.1505
R15 VDD.n4 VDD.n3 3.1505
R16 VDD.n5 VDD.n0 0.567623
R17 VDD VDD.n7 0.103227
R18 VDD VDD.n0 0.0319151
R19 VDD.n4 VDD.n1 0.0122537
R20 VDD VDD.n5 0.00140909
R21 VSS.t4 VSS.n0 2649.77
R22 VSS.n2 VSS.t4 1537.16
R23 VSS.n2 VSS.t2 1420.05
R24 VSS VSS.n0 992.072
R25 VSS.n0 VSS.t0 452.627
R26 VSS VSS.t3 9.22192
R27 VSS.n4 VSS.t5 9.0005
R28 VSS.n5 VSS.t1 8.96939
R29 VSS VSS.n3 2.6005
R30 VSS.n3 VSS.n2 2.6005
R31 VSS.n5 VSS.n4 0.445721
R32 VSS.n4 VSS 0.100854
R33 VSS VSS.n5 0.0689956
R34 VSS.n3 VSS.n1 0.00721141
R35 B.t1 B.t2 46.118
R36 B.n0 B.t1 30.0142
R37 B.n0 B.t0 12.341
R38 B B.n0 4.51075
R39 OUT.n2 OUT.n1 9.02722
R40 OUT.n2 OUT.n0 6.48941
R41 OUT OUT.n2 0.130713
C0 B a_230_424# 0.0242f
C1 a_230_424# VDD 0.886f
C2 OUT VDD 0.125f
C3 a_230_424# Inverter_0.IN 0.162f
C4 Inverter_0.IN OUT 0.116f
C5 B VDD 0.26f
C6 a_230_424# A 0.172f
C7 B Inverter_0.IN 0.0386f
C8 Inverter_0.IN VDD 0.305f
C9 OUT A 1.41e-19
C10 B A 0.241f
C11 A VDD 0.508f
C12 Inverter_0.IN A 0.258f
C13 A VSS 0.331f
C14 B VSS 0.497f
C15 OUT VSS 0.176f
C16 Inverter_0.IN VSS 0.769f
C17 a_230_424# VSS 0.167f
C18 VDD VSS 2.63f
.ends

