magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7578 -2492 7578 2492
<< nwell >>
rect -5578 -492 5578 492
<< nsubdiff >>
rect -5495 387 5495 409
rect -5495 341 -5428 387
rect 5428 341 5495 387
rect -5495 283 5495 341
rect -5495 237 -5428 283
rect 5428 237 5495 283
rect -5495 179 5495 237
rect -5495 133 -5428 179
rect 5428 133 5495 179
rect -5495 75 5495 133
rect -5495 29 -5428 75
rect 5428 29 5495 75
rect -5495 -29 5495 29
rect -5495 -75 -5428 -29
rect 5428 -75 5495 -29
rect -5495 -133 5495 -75
rect -5495 -179 -5428 -133
rect 5428 -179 5495 -133
rect -5495 -237 5495 -179
rect -5495 -283 -5428 -237
rect 5428 -283 5495 -237
rect -5495 -341 5495 -283
rect -5495 -387 -5428 -341
rect 5428 -387 5495 -341
rect -5495 -409 5495 -387
<< nsubdiffcont >>
rect -5428 341 5428 387
rect -5428 237 5428 283
rect -5428 133 5428 179
rect -5428 29 5428 75
rect -5428 -75 5428 -29
rect -5428 -179 5428 -133
rect -5428 -283 5428 -237
rect -5428 -387 5428 -341
<< metal1 >>
rect -5484 387 5484 398
rect -5484 341 -5428 387
rect 5428 341 5484 387
rect -5484 283 5484 341
rect -5484 237 -5428 283
rect 5428 237 5484 283
rect -5484 179 5484 237
rect -5484 133 -5428 179
rect 5428 133 5484 179
rect -5484 75 5484 133
rect -5484 29 -5428 75
rect 5428 29 5484 75
rect -5484 -29 5484 29
rect -5484 -75 -5428 -29
rect 5428 -75 5484 -29
rect -5484 -133 5484 -75
rect -5484 -179 -5428 -133
rect 5428 -179 5484 -133
rect -5484 -237 5484 -179
rect -5484 -283 -5428 -237
rect 5428 -283 5484 -237
rect -5484 -341 5484 -283
rect -5484 -387 -5428 -341
rect 5428 -387 5484 -341
rect -5484 -398 5484 -387
<< end >>
