magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2051 -1509 15725 19038
<< nwell >>
rect -51 491 13725 4487
<< psubdiff >>
rect 1565 17016 1901 17038
rect 1565 16970 1587 17016
rect 1633 16970 1701 17016
rect 1747 16970 1901 17016
rect 1565 16902 1901 16970
rect 1565 16856 1587 16902
rect 1633 16856 1701 16902
rect 1747 16856 1901 16902
rect 1565 16834 1901 16856
rect 1565 16788 1769 16834
rect 1565 16742 1587 16788
rect 1633 16742 1701 16788
rect 1747 16742 1769 16788
rect 1565 16218 1769 16742
rect 1565 16172 1587 16218
rect 1633 16172 1701 16218
rect 1747 16172 1769 16218
rect 1565 16104 1769 16172
rect 1565 16058 1587 16104
rect 1633 16058 1701 16104
rect 1747 16058 1769 16104
rect 1565 15990 1769 16058
rect 1565 15944 1587 15990
rect 1633 15944 1701 15990
rect 1747 15944 1769 15990
rect 1565 15876 1769 15944
rect 1565 15830 1587 15876
rect 1633 15830 1701 15876
rect 1747 15830 1769 15876
rect 1565 15762 1769 15830
rect 1565 15716 1587 15762
rect 1633 15716 1701 15762
rect 1747 15716 1769 15762
rect 1565 15648 1769 15716
rect 1565 15602 1587 15648
rect 1633 15602 1701 15648
rect 1747 15602 1769 15648
rect 1565 15534 1769 15602
rect 1565 15488 1587 15534
rect 1633 15488 1701 15534
rect 1747 15488 1769 15534
rect 1565 15420 1769 15488
rect 1565 15374 1587 15420
rect 1633 15374 1701 15420
rect 1747 15374 1769 15420
rect 1565 15306 1769 15374
rect 1565 15260 1587 15306
rect 1633 15260 1701 15306
rect 1747 15260 1769 15306
rect 1565 15192 1769 15260
rect 1565 15146 1587 15192
rect 1633 15146 1701 15192
rect 1747 15146 1769 15192
rect 1565 15078 1769 15146
rect 1565 15032 1587 15078
rect 1633 15032 1701 15078
rect 1747 15032 1769 15078
rect 1565 14964 1769 15032
rect 1565 14918 1587 14964
rect 1633 14918 1701 14964
rect 1747 14918 1769 14964
rect 1565 14850 1769 14918
rect 1565 14804 1587 14850
rect 1633 14804 1701 14850
rect 1747 14804 1769 14850
rect 1565 14736 1769 14804
rect 1565 14690 1587 14736
rect 1633 14690 1701 14736
rect 1747 14690 1769 14736
rect 1565 14622 1769 14690
rect 1565 14576 1587 14622
rect 1633 14576 1701 14622
rect 1747 14576 1769 14622
rect 1565 14508 1769 14576
rect 1565 14462 1587 14508
rect 1633 14462 1701 14508
rect 1747 14462 1769 14508
rect 1565 14394 1769 14462
rect 1565 14348 1587 14394
rect 1633 14348 1701 14394
rect 1747 14348 1769 14394
rect 1565 14280 1769 14348
rect 1565 14234 1587 14280
rect 1633 14234 1701 14280
rect 1747 14234 1769 14280
rect 1565 14166 1769 14234
rect 1565 14120 1587 14166
rect 1633 14120 1701 14166
rect 1747 14120 1769 14166
rect 1565 14052 1769 14120
rect 1565 14006 1587 14052
rect 1633 14006 1701 14052
rect 1747 14006 1769 14052
rect 1565 13938 1769 14006
rect 1565 13892 1587 13938
rect 1633 13892 1701 13938
rect 1747 13892 1769 13938
rect 1565 13824 1769 13892
rect 1565 13778 1587 13824
rect 1633 13778 1701 13824
rect 1747 13778 1769 13824
rect 1565 13710 1769 13778
rect 1565 13664 1587 13710
rect 1633 13664 1701 13710
rect 1747 13664 1769 13710
rect 1565 13596 1769 13664
rect 1565 13550 1587 13596
rect 1633 13550 1701 13596
rect 1747 13550 1769 13596
rect 1565 13482 1769 13550
rect 1565 13436 1587 13482
rect 1633 13436 1701 13482
rect 1747 13436 1769 13482
rect 1565 13368 1769 13436
rect 1565 13322 1587 13368
rect 1633 13322 1701 13368
rect 1747 13322 1769 13368
rect 1565 13254 1769 13322
rect 1565 13208 1587 13254
rect 1633 13208 1701 13254
rect 1747 13208 1769 13254
rect 1565 13140 1769 13208
rect 1565 13094 1587 13140
rect 1633 13094 1701 13140
rect 1747 13094 1769 13140
rect 1565 13026 1769 13094
rect 1565 12980 1587 13026
rect 1633 12980 1701 13026
rect 1747 12980 1769 13026
rect 1565 12912 1769 12980
rect 1565 12866 1587 12912
rect 1633 12866 1701 12912
rect 1747 12866 1769 12912
rect 1565 12798 1769 12866
rect 1565 12752 1587 12798
rect 1633 12752 1701 12798
rect 1747 12752 1769 12798
rect 1565 12684 1769 12752
rect 1565 12638 1587 12684
rect 1633 12638 1701 12684
rect 1747 12638 1769 12684
rect 1565 12570 1769 12638
rect 1565 12524 1587 12570
rect 1633 12524 1701 12570
rect 1747 12524 1769 12570
rect 1565 12456 1769 12524
rect 1565 12410 1587 12456
rect 1633 12410 1701 12456
rect 1747 12410 1769 12456
rect 1565 12342 1769 12410
rect 1565 12296 1587 12342
rect 1633 12296 1701 12342
rect 1747 12296 1769 12342
rect 1565 12228 1769 12296
rect 1565 12182 1587 12228
rect 1633 12182 1701 12228
rect 1747 12182 1769 12228
rect 1565 12114 1769 12182
rect 1565 12068 1587 12114
rect 1633 12068 1701 12114
rect 1747 12068 1769 12114
rect 1565 12000 1769 12068
rect 1565 11954 1587 12000
rect 1633 11954 1701 12000
rect 1747 11954 1769 12000
rect 1565 11886 1769 11954
rect 1565 11840 1587 11886
rect 1633 11840 1701 11886
rect 1747 11840 1769 11886
rect 1565 11772 1769 11840
rect 1565 11726 1587 11772
rect 1633 11726 1701 11772
rect 1747 11726 1769 11772
rect 1565 11658 1769 11726
rect 1565 11612 1587 11658
rect 1633 11612 1701 11658
rect 1747 11612 1769 11658
rect 1565 11544 1769 11612
rect 1565 11498 1587 11544
rect 1633 11498 1701 11544
rect 1747 11498 1769 11544
rect 1565 11430 1769 11498
rect 1565 11384 1587 11430
rect 1633 11384 1701 11430
rect 1747 11384 1769 11430
rect 1565 11316 1769 11384
rect 1565 11270 1587 11316
rect 1633 11270 1701 11316
rect 1747 11270 1769 11316
rect 1565 11202 1769 11270
rect 1565 11156 1587 11202
rect 1633 11156 1701 11202
rect 1747 11156 1769 11202
rect 1565 11088 1769 11156
rect 1565 11042 1587 11088
rect 1633 11042 1701 11088
rect 1747 11042 1769 11088
rect 1565 10974 1769 11042
rect 1565 10928 1587 10974
rect 1633 10928 1701 10974
rect 1747 10947 1769 10974
rect 1747 10928 1833 10947
rect 1565 10860 1833 10928
rect 1565 10814 1587 10860
rect 1633 10814 1701 10860
rect 1747 10814 1833 10860
rect 1565 10746 1833 10814
rect 1565 10700 1587 10746
rect 1633 10700 1701 10746
rect 1747 10743 1833 10746
rect 1747 10700 1769 10743
rect 1565 10632 1769 10700
rect 1565 10586 1587 10632
rect 1633 10586 1701 10632
rect 1747 10586 1769 10632
rect 1565 10518 1769 10586
rect 1565 10472 1587 10518
rect 1633 10472 1701 10518
rect 1747 10472 1769 10518
rect 1565 10404 1769 10472
rect 1565 10358 1587 10404
rect 1633 10358 1701 10404
rect 1747 10358 1769 10404
rect 1565 10290 1769 10358
rect 1565 10244 1587 10290
rect 1633 10244 1701 10290
rect 1747 10244 1769 10290
rect 1565 10176 1769 10244
rect 1565 10130 1587 10176
rect 1633 10130 1701 10176
rect 1747 10130 1769 10176
rect 1565 10062 1769 10130
rect 1565 10016 1587 10062
rect 1633 10016 1701 10062
rect 1747 10016 1769 10062
rect 1565 9948 1769 10016
rect 1565 9902 1587 9948
rect 1633 9902 1701 9948
rect 1747 9902 1769 9948
rect 1565 9834 1769 9902
rect 1565 9788 1587 9834
rect 1633 9788 1701 9834
rect 1747 9788 1769 9834
rect 1565 9720 1769 9788
rect 1565 9674 1587 9720
rect 1633 9674 1701 9720
rect 1747 9674 1769 9720
rect 1565 9606 1769 9674
rect 1565 9560 1587 9606
rect 1633 9560 1701 9606
rect 1747 9560 1769 9606
rect 1565 9492 1769 9560
rect 1565 9446 1587 9492
rect 1633 9446 1701 9492
rect 1747 9446 1769 9492
rect 1565 9378 1769 9446
rect 1565 9332 1587 9378
rect 1633 9332 1701 9378
rect 1747 9332 1769 9378
rect 1565 9264 1769 9332
rect 1565 9218 1587 9264
rect 1633 9218 1701 9264
rect 1747 9218 1769 9264
rect 1565 9150 1769 9218
rect 1565 9104 1587 9150
rect 1633 9104 1701 9150
rect 1747 9104 1769 9150
rect 1565 9036 1769 9104
rect 1565 8990 1587 9036
rect 1633 8990 1701 9036
rect 1747 8990 1769 9036
rect 1565 8922 1769 8990
rect 1565 8876 1587 8922
rect 1633 8876 1701 8922
rect 1747 8876 1769 8922
rect 1565 8808 1769 8876
rect 1565 8762 1587 8808
rect 1633 8762 1701 8808
rect 1747 8762 1769 8808
rect 1565 8694 1769 8762
rect 1565 8648 1587 8694
rect 1633 8648 1701 8694
rect 1747 8648 1769 8694
rect 1565 8580 1769 8648
rect 1565 8534 1587 8580
rect 1633 8534 1701 8580
rect 1747 8534 1769 8580
rect 1565 8466 1769 8534
rect 1565 8420 1587 8466
rect 1633 8420 1701 8466
rect 1747 8420 1769 8466
rect 1565 8352 1769 8420
rect 1565 8306 1587 8352
rect 1633 8306 1701 8352
rect 1747 8306 1769 8352
rect 1565 8238 1769 8306
rect 1565 8192 1587 8238
rect 1633 8192 1701 8238
rect 1747 8192 1769 8238
rect 1565 8124 1769 8192
rect 1565 8078 1587 8124
rect 1633 8078 1701 8124
rect 1747 8078 1769 8124
rect 1565 8010 1769 8078
rect 1565 7964 1587 8010
rect 1633 7964 1701 8010
rect 1747 7964 1769 8010
rect 1565 7896 1769 7964
rect 1565 7850 1587 7896
rect 1633 7850 1701 7896
rect 1747 7850 1769 7896
rect 1565 7782 1769 7850
rect 1565 7736 1587 7782
rect 1633 7736 1701 7782
rect 1747 7736 1769 7782
rect 1565 7668 1769 7736
rect 1565 7622 1587 7668
rect 1633 7622 1701 7668
rect 1747 7622 1769 7668
rect 1565 7554 1769 7622
rect 1565 7508 1587 7554
rect 1633 7508 1701 7554
rect 1747 7508 1769 7554
rect 1565 7440 1769 7508
rect 1565 7394 1587 7440
rect 1633 7394 1701 7440
rect 1747 7394 1769 7440
rect 1565 7326 1769 7394
rect 1565 7280 1587 7326
rect 1633 7280 1701 7326
rect 1747 7280 1769 7326
rect 1565 7212 1769 7280
rect 1565 7166 1587 7212
rect 1633 7166 1701 7212
rect 1747 7166 1769 7212
rect 1565 7098 1769 7166
rect 1565 7052 1587 7098
rect 1633 7052 1701 7098
rect 1747 7052 1769 7098
rect 1565 6984 1769 7052
rect 1565 6938 1587 6984
rect 1633 6938 1701 6984
rect 1747 6938 1769 6984
rect 1565 6870 1769 6938
rect 1565 6824 1587 6870
rect 1633 6824 1701 6870
rect 1747 6824 1769 6870
rect 1565 6756 1769 6824
rect 1565 6710 1587 6756
rect 1633 6710 1701 6756
rect 1747 6710 1769 6756
rect 1565 6642 1769 6710
rect 1565 6596 1587 6642
rect 1633 6596 1701 6642
rect 1747 6596 1769 6642
rect 1565 6528 1769 6596
rect 1565 6482 1587 6528
rect 1633 6482 1701 6528
rect 1747 6482 1769 6528
rect 1565 6414 1769 6482
rect 1565 6368 1587 6414
rect 1633 6368 1701 6414
rect 1747 6368 1769 6414
rect 1565 6300 1769 6368
rect 1565 6254 1587 6300
rect 1633 6254 1701 6300
rect 1747 6254 1769 6300
rect 1565 6186 1769 6254
rect 1565 6140 1587 6186
rect 1633 6140 1701 6186
rect 1747 6140 1769 6186
rect 1565 6072 1769 6140
rect 1565 6026 1587 6072
rect 1633 6026 1701 6072
rect 1747 6026 1769 6072
rect 1565 5958 1769 6026
rect 1565 5912 1587 5958
rect 1633 5912 1701 5958
rect 1747 5912 1769 5958
rect 1565 5844 1769 5912
rect 1565 5798 1587 5844
rect 1633 5798 1701 5844
rect 1747 5798 1769 5844
rect 1565 5730 1769 5798
rect 1565 5684 1587 5730
rect 1633 5684 1701 5730
rect 1747 5684 1769 5730
rect 1565 5616 1769 5684
rect 1565 5570 1587 5616
rect 1633 5570 1701 5616
rect 1747 5570 1769 5616
rect 1565 5502 1769 5570
rect 1565 5456 1587 5502
rect 1633 5456 1701 5502
rect 1747 5456 1769 5502
rect 1565 5046 1769 5456
rect 1565 5000 1587 5046
rect 1633 5000 1701 5046
rect 1747 5000 1769 5046
rect 1565 4954 1769 5000
rect 1565 4932 1901 4954
rect 1565 4886 1587 4932
rect 1633 4886 1701 4932
rect 1747 4886 1901 4932
rect 1565 4818 1901 4886
rect 1565 4772 1587 4818
rect 1633 4772 1701 4818
rect 1747 4772 1901 4818
rect 1565 4750 1901 4772
<< nsubdiff >>
rect 32 4382 13642 4404
rect 32 4336 54 4382
rect 100 4336 158 4382
rect 204 4336 574 4382
rect 620 4336 678 4382
rect 724 4336 782 4382
rect 828 4336 886 4382
rect 932 4336 990 4382
rect 1036 4336 1094 4382
rect 1140 4336 1198 4382
rect 1244 4336 1302 4382
rect 1348 4336 1406 4382
rect 1452 4336 1510 4382
rect 1556 4336 1614 4382
rect 1660 4336 1718 4382
rect 1764 4336 1822 4382
rect 1868 4336 1926 4382
rect 1972 4336 2030 4382
rect 2076 4336 2134 4382
rect 2180 4336 2238 4382
rect 2284 4336 2342 4382
rect 2388 4336 2446 4382
rect 2492 4336 2550 4382
rect 2596 4336 2654 4382
rect 2700 4336 2758 4382
rect 2804 4336 2862 4382
rect 2908 4336 2966 4382
rect 3012 4336 3070 4382
rect 3116 4336 3174 4382
rect 3220 4336 3278 4382
rect 3324 4336 3382 4382
rect 3428 4336 3486 4382
rect 3532 4336 3590 4382
rect 3636 4336 3694 4382
rect 3740 4336 3798 4382
rect 3844 4336 3902 4382
rect 3948 4336 4006 4382
rect 4052 4336 4110 4382
rect 4156 4336 4214 4382
rect 4260 4336 4318 4382
rect 4364 4336 4422 4382
rect 4468 4336 4526 4382
rect 4572 4336 4630 4382
rect 4676 4336 4734 4382
rect 4780 4336 4838 4382
rect 4884 4336 4942 4382
rect 4988 4336 5046 4382
rect 5092 4336 5150 4382
rect 5196 4336 5254 4382
rect 5300 4336 5358 4382
rect 5404 4336 5462 4382
rect 5508 4336 5566 4382
rect 5612 4336 5670 4382
rect 5716 4336 5774 4382
rect 5820 4336 5878 4382
rect 5924 4336 5982 4382
rect 6028 4336 6086 4382
rect 6132 4336 6190 4382
rect 6236 4336 6294 4382
rect 6340 4336 6398 4382
rect 6444 4336 6502 4382
rect 6548 4336 6606 4382
rect 6652 4336 6710 4382
rect 6756 4336 6814 4382
rect 6860 4336 6918 4382
rect 6964 4336 7022 4382
rect 7068 4336 7126 4382
rect 7172 4336 7230 4382
rect 7276 4336 7334 4382
rect 7380 4336 7438 4382
rect 7484 4336 7542 4382
rect 7588 4336 7646 4382
rect 7692 4336 7750 4382
rect 7796 4336 7854 4382
rect 7900 4336 7958 4382
rect 8004 4336 8062 4382
rect 8108 4336 8166 4382
rect 8212 4336 8270 4382
rect 8316 4336 8374 4382
rect 8420 4336 8478 4382
rect 8524 4336 8582 4382
rect 8628 4336 8686 4382
rect 8732 4336 8790 4382
rect 8836 4336 8894 4382
rect 8940 4336 8998 4382
rect 9044 4336 9102 4382
rect 9148 4336 9206 4382
rect 9252 4336 9310 4382
rect 9356 4336 9414 4382
rect 9460 4336 9518 4382
rect 9564 4336 9622 4382
rect 9668 4336 9726 4382
rect 9772 4336 9830 4382
rect 9876 4336 9934 4382
rect 9980 4336 10038 4382
rect 10084 4336 10142 4382
rect 10188 4336 10246 4382
rect 10292 4336 10350 4382
rect 10396 4336 10454 4382
rect 10500 4336 10558 4382
rect 10604 4336 10662 4382
rect 10708 4336 10766 4382
rect 10812 4336 10870 4382
rect 10916 4336 10974 4382
rect 11020 4336 11078 4382
rect 11124 4336 11182 4382
rect 11228 4336 11286 4382
rect 11332 4336 11390 4382
rect 11436 4336 11494 4382
rect 11540 4336 11598 4382
rect 11644 4336 11702 4382
rect 11748 4336 11806 4382
rect 11852 4336 11910 4382
rect 11956 4336 12014 4382
rect 12060 4336 12118 4382
rect 12164 4336 12222 4382
rect 12268 4336 12326 4382
rect 12372 4336 12430 4382
rect 12476 4336 12534 4382
rect 12580 4336 12638 4382
rect 12684 4336 12742 4382
rect 12788 4336 12846 4382
rect 12892 4336 12950 4382
rect 12996 4336 13054 4382
rect 13100 4336 13158 4382
rect 13204 4336 13262 4382
rect 13308 4336 13366 4382
rect 13412 4336 13470 4382
rect 13516 4336 13574 4382
rect 13620 4336 13642 4382
rect 32 4314 13642 4336
rect 32 4182 122 4314
rect 13552 4182 13642 4314
<< psubdiffcont >>
rect 1587 16970 1633 17016
rect 1701 16970 1747 17016
rect 1587 16856 1633 16902
rect 1701 16856 1747 16902
rect 1587 16742 1633 16788
rect 1701 16742 1747 16788
rect 1587 16172 1633 16218
rect 1701 16172 1747 16218
rect 1587 16058 1633 16104
rect 1701 16058 1747 16104
rect 1587 15944 1633 15990
rect 1701 15944 1747 15990
rect 1587 15830 1633 15876
rect 1701 15830 1747 15876
rect 1587 15716 1633 15762
rect 1701 15716 1747 15762
rect 1587 15602 1633 15648
rect 1701 15602 1747 15648
rect 1587 15488 1633 15534
rect 1701 15488 1747 15534
rect 1587 15374 1633 15420
rect 1701 15374 1747 15420
rect 1587 15260 1633 15306
rect 1701 15260 1747 15306
rect 1587 15146 1633 15192
rect 1701 15146 1747 15192
rect 1587 15032 1633 15078
rect 1701 15032 1747 15078
rect 1587 14918 1633 14964
rect 1701 14918 1747 14964
rect 1587 14804 1633 14850
rect 1701 14804 1747 14850
rect 1587 14690 1633 14736
rect 1701 14690 1747 14736
rect 1587 14576 1633 14622
rect 1701 14576 1747 14622
rect 1587 14462 1633 14508
rect 1701 14462 1747 14508
rect 1587 14348 1633 14394
rect 1701 14348 1747 14394
rect 1587 14234 1633 14280
rect 1701 14234 1747 14280
rect 1587 14120 1633 14166
rect 1701 14120 1747 14166
rect 1587 14006 1633 14052
rect 1701 14006 1747 14052
rect 1587 13892 1633 13938
rect 1701 13892 1747 13938
rect 1587 13778 1633 13824
rect 1701 13778 1747 13824
rect 1587 13664 1633 13710
rect 1701 13664 1747 13710
rect 1587 13550 1633 13596
rect 1701 13550 1747 13596
rect 1587 13436 1633 13482
rect 1701 13436 1747 13482
rect 1587 13322 1633 13368
rect 1701 13322 1747 13368
rect 1587 13208 1633 13254
rect 1701 13208 1747 13254
rect 1587 13094 1633 13140
rect 1701 13094 1747 13140
rect 1587 12980 1633 13026
rect 1701 12980 1747 13026
rect 1587 12866 1633 12912
rect 1701 12866 1747 12912
rect 1587 12752 1633 12798
rect 1701 12752 1747 12798
rect 1587 12638 1633 12684
rect 1701 12638 1747 12684
rect 1587 12524 1633 12570
rect 1701 12524 1747 12570
rect 1587 12410 1633 12456
rect 1701 12410 1747 12456
rect 1587 12296 1633 12342
rect 1701 12296 1747 12342
rect 1587 12182 1633 12228
rect 1701 12182 1747 12228
rect 1587 12068 1633 12114
rect 1701 12068 1747 12114
rect 1587 11954 1633 12000
rect 1701 11954 1747 12000
rect 1587 11840 1633 11886
rect 1701 11840 1747 11886
rect 1587 11726 1633 11772
rect 1701 11726 1747 11772
rect 1587 11612 1633 11658
rect 1701 11612 1747 11658
rect 1587 11498 1633 11544
rect 1701 11498 1747 11544
rect 1587 11384 1633 11430
rect 1701 11384 1747 11430
rect 1587 11270 1633 11316
rect 1701 11270 1747 11316
rect 1587 11156 1633 11202
rect 1701 11156 1747 11202
rect 1587 11042 1633 11088
rect 1701 11042 1747 11088
rect 1587 10928 1633 10974
rect 1701 10928 1747 10974
rect 1587 10814 1633 10860
rect 1701 10814 1747 10860
rect 1587 10700 1633 10746
rect 1701 10700 1747 10746
rect 1587 10586 1633 10632
rect 1701 10586 1747 10632
rect 1587 10472 1633 10518
rect 1701 10472 1747 10518
rect 1587 10358 1633 10404
rect 1701 10358 1747 10404
rect 1587 10244 1633 10290
rect 1701 10244 1747 10290
rect 1587 10130 1633 10176
rect 1701 10130 1747 10176
rect 1587 10016 1633 10062
rect 1701 10016 1747 10062
rect 1587 9902 1633 9948
rect 1701 9902 1747 9948
rect 1587 9788 1633 9834
rect 1701 9788 1747 9834
rect 1587 9674 1633 9720
rect 1701 9674 1747 9720
rect 1587 9560 1633 9606
rect 1701 9560 1747 9606
rect 1587 9446 1633 9492
rect 1701 9446 1747 9492
rect 1587 9332 1633 9378
rect 1701 9332 1747 9378
rect 1587 9218 1633 9264
rect 1701 9218 1747 9264
rect 1587 9104 1633 9150
rect 1701 9104 1747 9150
rect 1587 8990 1633 9036
rect 1701 8990 1747 9036
rect 1587 8876 1633 8922
rect 1701 8876 1747 8922
rect 1587 8762 1633 8808
rect 1701 8762 1747 8808
rect 1587 8648 1633 8694
rect 1701 8648 1747 8694
rect 1587 8534 1633 8580
rect 1701 8534 1747 8580
rect 1587 8420 1633 8466
rect 1701 8420 1747 8466
rect 1587 8306 1633 8352
rect 1701 8306 1747 8352
rect 1587 8192 1633 8238
rect 1701 8192 1747 8238
rect 1587 8078 1633 8124
rect 1701 8078 1747 8124
rect 1587 7964 1633 8010
rect 1701 7964 1747 8010
rect 1587 7850 1633 7896
rect 1701 7850 1747 7896
rect 1587 7736 1633 7782
rect 1701 7736 1747 7782
rect 1587 7622 1633 7668
rect 1701 7622 1747 7668
rect 1587 7508 1633 7554
rect 1701 7508 1747 7554
rect 1587 7394 1633 7440
rect 1701 7394 1747 7440
rect 1587 7280 1633 7326
rect 1701 7280 1747 7326
rect 1587 7166 1633 7212
rect 1701 7166 1747 7212
rect 1587 7052 1633 7098
rect 1701 7052 1747 7098
rect 1587 6938 1633 6984
rect 1701 6938 1747 6984
rect 1587 6824 1633 6870
rect 1701 6824 1747 6870
rect 1587 6710 1633 6756
rect 1701 6710 1747 6756
rect 1587 6596 1633 6642
rect 1701 6596 1747 6642
rect 1587 6482 1633 6528
rect 1701 6482 1747 6528
rect 1587 6368 1633 6414
rect 1701 6368 1747 6414
rect 1587 6254 1633 6300
rect 1701 6254 1747 6300
rect 1587 6140 1633 6186
rect 1701 6140 1747 6186
rect 1587 6026 1633 6072
rect 1701 6026 1747 6072
rect 1587 5912 1633 5958
rect 1701 5912 1747 5958
rect 1587 5798 1633 5844
rect 1701 5798 1747 5844
rect 1587 5684 1633 5730
rect 1701 5684 1747 5730
rect 1587 5570 1633 5616
rect 1701 5570 1747 5616
rect 1587 5456 1633 5502
rect 1701 5456 1747 5502
rect 1587 5000 1633 5046
rect 1701 5000 1747 5046
rect 1587 4886 1633 4932
rect 1701 4886 1747 4932
rect 1587 4772 1633 4818
rect 1701 4772 1747 4818
<< nsubdiffcont >>
rect 54 4336 100 4382
rect 158 4336 204 4382
rect 574 4336 620 4382
rect 678 4336 724 4382
rect 782 4336 828 4382
rect 886 4336 932 4382
rect 990 4336 1036 4382
rect 1094 4336 1140 4382
rect 1198 4336 1244 4382
rect 1302 4336 1348 4382
rect 1406 4336 1452 4382
rect 1510 4336 1556 4382
rect 1614 4336 1660 4382
rect 1718 4336 1764 4382
rect 1822 4336 1868 4382
rect 1926 4336 1972 4382
rect 2030 4336 2076 4382
rect 2134 4336 2180 4382
rect 2238 4336 2284 4382
rect 2342 4336 2388 4382
rect 2446 4336 2492 4382
rect 2550 4336 2596 4382
rect 2654 4336 2700 4382
rect 2758 4336 2804 4382
rect 2862 4336 2908 4382
rect 2966 4336 3012 4382
rect 3070 4336 3116 4382
rect 3174 4336 3220 4382
rect 3278 4336 3324 4382
rect 3382 4336 3428 4382
rect 3486 4336 3532 4382
rect 3590 4336 3636 4382
rect 3694 4336 3740 4382
rect 3798 4336 3844 4382
rect 3902 4336 3948 4382
rect 4006 4336 4052 4382
rect 4110 4336 4156 4382
rect 4214 4336 4260 4382
rect 4318 4336 4364 4382
rect 4422 4336 4468 4382
rect 4526 4336 4572 4382
rect 4630 4336 4676 4382
rect 4734 4336 4780 4382
rect 4838 4336 4884 4382
rect 4942 4336 4988 4382
rect 5046 4336 5092 4382
rect 5150 4336 5196 4382
rect 5254 4336 5300 4382
rect 5358 4336 5404 4382
rect 5462 4336 5508 4382
rect 5566 4336 5612 4382
rect 5670 4336 5716 4382
rect 5774 4336 5820 4382
rect 5878 4336 5924 4382
rect 5982 4336 6028 4382
rect 6086 4336 6132 4382
rect 6190 4336 6236 4382
rect 6294 4336 6340 4382
rect 6398 4336 6444 4382
rect 6502 4336 6548 4382
rect 6606 4336 6652 4382
rect 6710 4336 6756 4382
rect 6814 4336 6860 4382
rect 6918 4336 6964 4382
rect 7022 4336 7068 4382
rect 7126 4336 7172 4382
rect 7230 4336 7276 4382
rect 7334 4336 7380 4382
rect 7438 4336 7484 4382
rect 7542 4336 7588 4382
rect 7646 4336 7692 4382
rect 7750 4336 7796 4382
rect 7854 4336 7900 4382
rect 7958 4336 8004 4382
rect 8062 4336 8108 4382
rect 8166 4336 8212 4382
rect 8270 4336 8316 4382
rect 8374 4336 8420 4382
rect 8478 4336 8524 4382
rect 8582 4336 8628 4382
rect 8686 4336 8732 4382
rect 8790 4336 8836 4382
rect 8894 4336 8940 4382
rect 8998 4336 9044 4382
rect 9102 4336 9148 4382
rect 9206 4336 9252 4382
rect 9310 4336 9356 4382
rect 9414 4336 9460 4382
rect 9518 4336 9564 4382
rect 9622 4336 9668 4382
rect 9726 4336 9772 4382
rect 9830 4336 9876 4382
rect 9934 4336 9980 4382
rect 10038 4336 10084 4382
rect 10142 4336 10188 4382
rect 10246 4336 10292 4382
rect 10350 4336 10396 4382
rect 10454 4336 10500 4382
rect 10558 4336 10604 4382
rect 10662 4336 10708 4382
rect 10766 4336 10812 4382
rect 10870 4336 10916 4382
rect 10974 4336 11020 4382
rect 11078 4336 11124 4382
rect 11182 4336 11228 4382
rect 11286 4336 11332 4382
rect 11390 4336 11436 4382
rect 11494 4336 11540 4382
rect 11598 4336 11644 4382
rect 11702 4336 11748 4382
rect 11806 4336 11852 4382
rect 11910 4336 11956 4382
rect 12014 4336 12060 4382
rect 12118 4336 12164 4382
rect 12222 4336 12268 4382
rect 12326 4336 12372 4382
rect 12430 4336 12476 4382
rect 12534 4336 12580 4382
rect 12638 4336 12684 4382
rect 12742 4336 12788 4382
rect 12846 4336 12892 4382
rect 12950 4336 12996 4382
rect 13054 4336 13100 4382
rect 13158 4336 13204 4382
rect 13262 4336 13308 4382
rect 13366 4336 13412 4382
rect 13470 4336 13516 4382
rect 13574 4336 13620 4382
<< metal1 >>
rect 1576 17016 12098 17028
rect 1576 16970 1587 17016
rect 1633 16970 1701 17016
rect 1747 16970 12098 17016
rect 1576 16902 12098 16970
rect 1576 16856 1587 16902
rect 1633 16856 1701 16902
rect 1747 16856 12098 16902
rect 1576 16844 12098 16856
rect 1576 16788 1758 16844
rect 1576 16742 1587 16788
rect 1633 16742 1701 16788
rect 1747 16742 1758 16788
rect 1576 16681 1758 16742
rect 306 16441 11446 16573
rect 306 16411 4138 16441
rect 306 5279 466 16411
rect 2222 16373 4138 16411
rect 4658 16373 6574 16441
rect 7094 16373 9010 16441
rect 9530 16373 11446 16441
rect 1576 16218 1962 16351
rect 1576 16172 1587 16218
rect 1633 16172 1701 16218
rect 1747 16172 1962 16218
rect 1576 16104 1962 16172
rect 1576 16058 1587 16104
rect 1633 16058 1701 16104
rect 1747 16058 1962 16104
rect 1576 15990 1962 16058
rect 1576 15944 1587 15990
rect 1633 15944 1701 15990
rect 1747 15944 1962 15990
rect 1576 15876 1962 15944
rect 1576 15830 1587 15876
rect 1633 15830 1701 15876
rect 1747 15830 1962 15876
rect 1576 15762 1962 15830
rect 1576 15716 1587 15762
rect 1633 15716 1701 15762
rect 1747 15716 1962 15762
rect 1576 15648 1962 15716
rect 1576 15602 1587 15648
rect 1633 15602 1701 15648
rect 1747 15602 1962 15648
rect 1576 15534 1962 15602
rect 1576 15488 1587 15534
rect 1633 15488 1701 15534
rect 1747 15488 1962 15534
rect 1576 15420 1962 15488
rect 1576 15374 1587 15420
rect 1633 15374 1701 15420
rect 1747 15374 1962 15420
rect 1576 15306 1962 15374
rect 1576 15260 1587 15306
rect 1633 15260 1701 15306
rect 1747 15260 1962 15306
rect 1576 15192 1962 15260
rect 1576 15146 1587 15192
rect 1633 15146 1701 15192
rect 1747 15146 1962 15192
rect 1576 15078 1962 15146
rect 1576 15032 1587 15078
rect 1633 15032 1701 15078
rect 1747 15032 1962 15078
rect 1576 14964 1962 15032
rect 1576 14918 1587 14964
rect 1633 14918 1701 14964
rect 1747 14918 1962 14964
rect 1576 14850 1962 14918
rect 1576 14804 1587 14850
rect 1633 14804 1701 14850
rect 1747 14804 1962 14850
rect 1576 14736 1962 14804
rect 1576 14690 1587 14736
rect 1633 14690 1701 14736
rect 1747 14690 1962 14736
rect 1576 14622 1962 14690
rect 1576 14576 1587 14622
rect 1633 14576 1701 14622
rect 1747 14576 1962 14622
rect 1576 14508 1962 14576
rect 1576 14462 1587 14508
rect 1633 14462 1701 14508
rect 1747 14462 1962 14508
rect 1576 14394 1962 14462
rect 1576 14348 1587 14394
rect 1633 14348 1701 14394
rect 1747 14348 1962 14394
rect 1576 14280 1962 14348
rect 1576 14234 1587 14280
rect 1633 14234 1701 14280
rect 1747 14234 1962 14280
rect 1576 14166 1962 14234
rect 1576 14120 1587 14166
rect 1633 14120 1701 14166
rect 1747 14120 1962 14166
rect 1576 14052 1962 14120
rect 1576 14006 1587 14052
rect 1633 14006 1701 14052
rect 1747 14006 1962 14052
rect 1576 13938 1962 14006
rect 1576 13892 1587 13938
rect 1633 13892 1701 13938
rect 1747 13892 1962 13938
rect 1576 13824 1962 13892
rect 1576 13778 1587 13824
rect 1633 13778 1701 13824
rect 1747 13778 1962 13824
rect 1576 13710 1962 13778
rect 1576 13664 1587 13710
rect 1633 13664 1701 13710
rect 1747 13664 1962 13710
rect 1576 13596 1962 13664
rect 1576 13550 1587 13596
rect 1633 13550 1701 13596
rect 1747 13550 1962 13596
rect 1576 13482 1962 13550
rect 1576 13436 1587 13482
rect 1633 13436 1701 13482
rect 1747 13436 1962 13482
rect 1576 13368 1962 13436
rect 1576 13322 1587 13368
rect 1633 13322 1701 13368
rect 1747 13322 1962 13368
rect 1576 13254 1962 13322
rect 1576 13208 1587 13254
rect 1633 13208 1701 13254
rect 1747 13208 1962 13254
rect 1576 13140 1962 13208
rect 1576 13094 1587 13140
rect 1633 13094 1701 13140
rect 1747 13094 1962 13140
rect 1576 13026 1962 13094
rect 1576 12980 1587 13026
rect 1633 12980 1701 13026
rect 1747 12980 1962 13026
rect 1576 12912 1962 12980
rect 1576 12866 1587 12912
rect 1633 12866 1701 12912
rect 1747 12866 1962 12912
rect 1576 12798 1962 12866
rect 1576 12752 1587 12798
rect 1633 12752 1701 12798
rect 1747 12752 1962 12798
rect 1576 12684 1962 12752
rect 1576 12638 1587 12684
rect 1633 12638 1701 12684
rect 1747 12638 1962 12684
rect 1576 12570 1962 12638
rect 1576 12524 1587 12570
rect 1633 12524 1701 12570
rect 1747 12524 1962 12570
rect 1576 12456 1962 12524
rect 1576 12410 1587 12456
rect 1633 12410 1701 12456
rect 1747 12410 1962 12456
rect 1576 12342 1962 12410
rect 1576 12296 1587 12342
rect 1633 12296 1701 12342
rect 1747 12296 1962 12342
rect 1576 12228 1962 12296
rect 1576 12182 1587 12228
rect 1633 12182 1701 12228
rect 1747 12182 1962 12228
rect 1576 12114 1962 12182
rect 1576 12068 1587 12114
rect 1633 12068 1701 12114
rect 1747 12068 1962 12114
rect 1576 12000 1962 12068
rect 1576 11954 1587 12000
rect 1633 11954 1701 12000
rect 1747 11954 1962 12000
rect 1576 11886 1962 11954
rect 1576 11840 1587 11886
rect 1633 11840 1701 11886
rect 1747 11840 1962 11886
rect 1576 11772 1962 11840
rect 1576 11726 1587 11772
rect 1633 11726 1701 11772
rect 1747 11726 1962 11772
rect 1576 11658 1962 11726
rect 1576 11612 1587 11658
rect 1633 11612 1701 11658
rect 1747 11612 1962 11658
rect 1576 11544 1962 11612
rect 1576 11498 1587 11544
rect 1633 11498 1701 11544
rect 1747 11498 1962 11544
rect 1576 11430 1962 11498
rect 1576 11384 1587 11430
rect 1633 11384 1701 11430
rect 1747 11384 1962 11430
rect 1576 11316 1962 11384
rect 1576 11270 1587 11316
rect 1633 11270 1701 11316
rect 1747 11270 1962 11316
rect 1576 11202 1962 11270
rect 1576 11156 1587 11202
rect 1633 11156 1701 11202
rect 1747 11201 1962 11202
rect 11706 11201 11916 16351
rect 1747 11156 11916 11201
rect 1576 11088 11916 11156
rect 1576 11042 1587 11088
rect 1633 11042 1701 11088
rect 1747 11042 11916 11088
rect 1576 10974 11916 11042
rect 1576 10928 1587 10974
rect 1633 10928 1701 10974
rect 1747 10928 11916 10974
rect 1576 10860 11916 10928
rect 1576 10814 1587 10860
rect 1633 10814 1701 10860
rect 1747 10814 11916 10860
rect 1576 10746 11916 10814
rect 1576 10700 1587 10746
rect 1633 10700 1701 10746
rect 1747 10700 11916 10746
rect 1576 10632 11916 10700
rect 1576 10586 1587 10632
rect 1633 10586 1701 10632
rect 1747 10586 11916 10632
rect 1576 10518 11916 10586
rect 1576 10472 1587 10518
rect 1633 10472 1701 10518
rect 1747 10489 11916 10518
rect 1747 10472 1962 10489
rect 1576 10404 1962 10472
rect 1576 10358 1587 10404
rect 1633 10358 1701 10404
rect 1747 10358 1962 10404
rect 1576 10290 1962 10358
rect 1576 10244 1587 10290
rect 1633 10244 1701 10290
rect 1747 10244 1962 10290
rect 1576 10176 1962 10244
rect 1576 10130 1587 10176
rect 1633 10130 1701 10176
rect 1747 10130 1962 10176
rect 1576 10062 1962 10130
rect 1576 10016 1587 10062
rect 1633 10016 1701 10062
rect 1747 10016 1962 10062
rect 1576 9948 1962 10016
rect 1576 9902 1587 9948
rect 1633 9902 1701 9948
rect 1747 9902 1962 9948
rect 1576 9834 1962 9902
rect 1576 9788 1587 9834
rect 1633 9788 1701 9834
rect 1747 9788 1962 9834
rect 1576 9720 1962 9788
rect 1576 9674 1587 9720
rect 1633 9674 1701 9720
rect 1747 9674 1962 9720
rect 1576 9606 1962 9674
rect 1576 9560 1587 9606
rect 1633 9560 1701 9606
rect 1747 9560 1962 9606
rect 1576 9492 1962 9560
rect 1576 9446 1587 9492
rect 1633 9446 1701 9492
rect 1747 9446 1962 9492
rect 1576 9378 1962 9446
rect 1576 9332 1587 9378
rect 1633 9332 1701 9378
rect 1747 9332 1962 9378
rect 1576 9264 1962 9332
rect 1576 9218 1587 9264
rect 1633 9218 1701 9264
rect 1747 9218 1962 9264
rect 1576 9150 1962 9218
rect 1576 9104 1587 9150
rect 1633 9104 1701 9150
rect 1747 9104 1962 9150
rect 1576 9036 1962 9104
rect 1576 8990 1587 9036
rect 1633 8990 1701 9036
rect 1747 8990 1962 9036
rect 1576 8922 1962 8990
rect 1576 8876 1587 8922
rect 1633 8876 1701 8922
rect 1747 8876 1962 8922
rect 1576 8808 1962 8876
rect 1576 8762 1587 8808
rect 1633 8762 1701 8808
rect 1747 8762 1962 8808
rect 1576 8694 1962 8762
rect 1576 8648 1587 8694
rect 1633 8648 1701 8694
rect 1747 8648 1962 8694
rect 1576 8580 1962 8648
rect 1576 8534 1587 8580
rect 1633 8534 1701 8580
rect 1747 8534 1962 8580
rect 1576 8466 1962 8534
rect 1576 8420 1587 8466
rect 1633 8420 1701 8466
rect 1747 8420 1962 8466
rect 1576 8352 1962 8420
rect 1576 8306 1587 8352
rect 1633 8306 1701 8352
rect 1747 8306 1962 8352
rect 1576 8238 1962 8306
rect 1576 8192 1587 8238
rect 1633 8192 1701 8238
rect 1747 8192 1962 8238
rect 1576 8124 1962 8192
rect 1576 8078 1587 8124
rect 1633 8078 1701 8124
rect 1747 8078 1962 8124
rect 1576 8010 1962 8078
rect 1576 7964 1587 8010
rect 1633 7964 1701 8010
rect 1747 7964 1962 8010
rect 1576 7896 1962 7964
rect 1576 7850 1587 7896
rect 1633 7850 1701 7896
rect 1747 7850 1962 7896
rect 1576 7782 1962 7850
rect 1576 7736 1587 7782
rect 1633 7736 1701 7782
rect 1747 7736 1962 7782
rect 1576 7668 1962 7736
rect 1576 7622 1587 7668
rect 1633 7622 1701 7668
rect 1747 7622 1962 7668
rect 1576 7554 1962 7622
rect 1576 7508 1587 7554
rect 1633 7508 1701 7554
rect 1747 7508 1962 7554
rect 1576 7440 1962 7508
rect 1576 7394 1587 7440
rect 1633 7394 1701 7440
rect 1747 7394 1962 7440
rect 1576 7326 1962 7394
rect 1576 7280 1587 7326
rect 1633 7280 1701 7326
rect 1747 7280 1962 7326
rect 1576 7212 1962 7280
rect 1576 7166 1587 7212
rect 1633 7166 1701 7212
rect 1747 7166 1962 7212
rect 1576 7098 1962 7166
rect 1576 7052 1587 7098
rect 1633 7052 1701 7098
rect 1747 7052 1962 7098
rect 1576 6984 1962 7052
rect 1576 6938 1587 6984
rect 1633 6938 1701 6984
rect 1747 6938 1962 6984
rect 1576 6870 1962 6938
rect 1576 6824 1587 6870
rect 1633 6824 1701 6870
rect 1747 6824 1962 6870
rect 1576 6756 1962 6824
rect 1576 6710 1587 6756
rect 1633 6710 1701 6756
rect 1747 6710 1962 6756
rect 1576 6642 1962 6710
rect 1576 6596 1587 6642
rect 1633 6596 1701 6642
rect 1747 6596 1962 6642
rect 1576 6528 1962 6596
rect 1576 6482 1587 6528
rect 1633 6482 1701 6528
rect 1747 6482 1962 6528
rect 1576 6414 1962 6482
rect 1576 6368 1587 6414
rect 1633 6368 1701 6414
rect 1747 6368 1962 6414
rect 1576 6300 1962 6368
rect 1576 6254 1587 6300
rect 1633 6254 1701 6300
rect 1747 6254 1962 6300
rect 1576 6186 1962 6254
rect 1576 6140 1587 6186
rect 1633 6140 1701 6186
rect 1747 6140 1962 6186
rect 1576 6072 1962 6140
rect 1576 6026 1587 6072
rect 1633 6026 1701 6072
rect 1747 6026 1962 6072
rect 1576 5958 1962 6026
rect 1576 5912 1587 5958
rect 1633 5912 1701 5958
rect 1747 5912 1962 5958
rect 1576 5844 1962 5912
rect 1576 5798 1587 5844
rect 1633 5798 1701 5844
rect 1747 5798 1962 5844
rect 1576 5730 1962 5798
rect 1576 5684 1587 5730
rect 1633 5684 1701 5730
rect 1747 5684 1962 5730
rect 1576 5616 1962 5684
rect 1576 5570 1587 5616
rect 1633 5570 1701 5616
rect 1747 5570 1962 5616
rect 1576 5502 1962 5570
rect 1576 5456 1587 5502
rect 1633 5456 1701 5502
rect 1747 5456 1962 5502
rect 1576 5339 1962 5456
rect 11706 5339 11916 10489
rect 2222 5279 4138 5317
rect 306 5249 4138 5279
rect 4658 5249 6574 5317
rect 7094 5249 9010 5317
rect 9530 5249 11446 5317
rect 306 5117 11446 5249
rect 43 4382 233 4393
rect 43 4336 54 4382
rect 100 4336 158 4382
rect 204 4336 233 4382
rect 43 4325 233 4336
rect 43 657 111 4325
rect 306 3951 466 5117
rect 1576 5046 1758 5067
rect 1576 5000 1587 5046
rect 1633 5000 1701 5046
rect 1747 5000 1758 5046
rect 1576 4944 1758 5000
rect 1576 4932 12098 4944
rect 1576 4886 1587 4932
rect 1633 4886 1701 4932
rect 1747 4886 12098 4932
rect 1576 4818 12098 4886
rect 1576 4772 1587 4818
rect 1633 4772 1701 4818
rect 1747 4772 12098 4818
rect 1576 4760 12098 4772
rect 540 4382 13631 4397
rect 540 4336 574 4382
rect 620 4336 678 4382
rect 724 4336 782 4382
rect 828 4336 886 4382
rect 932 4336 990 4382
rect 1036 4336 1094 4382
rect 1140 4336 1198 4382
rect 1244 4336 1302 4382
rect 1348 4336 1406 4382
rect 1452 4336 1510 4382
rect 1556 4336 1614 4382
rect 1660 4336 1718 4382
rect 1764 4336 1822 4382
rect 1868 4336 1926 4382
rect 1972 4336 2030 4382
rect 2076 4336 2134 4382
rect 2180 4336 2238 4382
rect 2284 4336 2342 4382
rect 2388 4336 2446 4382
rect 2492 4336 2550 4382
rect 2596 4336 2654 4382
rect 2700 4336 2758 4382
rect 2804 4336 2862 4382
rect 2908 4336 2966 4382
rect 3012 4336 3070 4382
rect 3116 4336 3174 4382
rect 3220 4336 3278 4382
rect 3324 4336 3382 4382
rect 3428 4336 3486 4382
rect 3532 4336 3590 4382
rect 3636 4336 3694 4382
rect 3740 4336 3798 4382
rect 3844 4336 3902 4382
rect 3948 4336 4006 4382
rect 4052 4336 4110 4382
rect 4156 4336 4214 4382
rect 4260 4336 4318 4382
rect 4364 4336 4422 4382
rect 4468 4336 4526 4382
rect 4572 4336 4630 4382
rect 4676 4336 4734 4382
rect 4780 4336 4838 4382
rect 4884 4336 4942 4382
rect 4988 4336 5046 4382
rect 5092 4336 5150 4382
rect 5196 4336 5254 4382
rect 5300 4336 5358 4382
rect 5404 4336 5462 4382
rect 5508 4336 5566 4382
rect 5612 4336 5670 4382
rect 5716 4336 5774 4382
rect 5820 4336 5878 4382
rect 5924 4336 5982 4382
rect 6028 4336 6086 4382
rect 6132 4336 6190 4382
rect 6236 4336 6294 4382
rect 6340 4336 6398 4382
rect 6444 4336 6502 4382
rect 6548 4336 6606 4382
rect 6652 4336 6710 4382
rect 6756 4336 6814 4382
rect 6860 4336 6918 4382
rect 6964 4336 7022 4382
rect 7068 4336 7126 4382
rect 7172 4336 7230 4382
rect 7276 4336 7334 4382
rect 7380 4336 7438 4382
rect 7484 4336 7542 4382
rect 7588 4336 7646 4382
rect 7692 4336 7750 4382
rect 7796 4336 7854 4382
rect 7900 4336 7958 4382
rect 8004 4336 8062 4382
rect 8108 4336 8166 4382
rect 8212 4336 8270 4382
rect 8316 4336 8374 4382
rect 8420 4336 8478 4382
rect 8524 4336 8582 4382
rect 8628 4336 8686 4382
rect 8732 4336 8790 4382
rect 8836 4336 8894 4382
rect 8940 4336 8998 4382
rect 9044 4336 9102 4382
rect 9148 4336 9206 4382
rect 9252 4336 9310 4382
rect 9356 4336 9414 4382
rect 9460 4336 9518 4382
rect 9564 4336 9622 4382
rect 9668 4336 9726 4382
rect 9772 4336 9830 4382
rect 9876 4336 9934 4382
rect 9980 4336 10038 4382
rect 10084 4336 10142 4382
rect 10188 4336 10246 4382
rect 10292 4336 10350 4382
rect 10396 4336 10454 4382
rect 10500 4336 10558 4382
rect 10604 4336 10662 4382
rect 10708 4336 10766 4382
rect 10812 4336 10870 4382
rect 10916 4336 10974 4382
rect 11020 4336 11078 4382
rect 11124 4336 11182 4382
rect 11228 4336 11286 4382
rect 11332 4336 11390 4382
rect 11436 4336 11494 4382
rect 11540 4336 11598 4382
rect 11644 4336 11702 4382
rect 11748 4336 11806 4382
rect 11852 4336 11910 4382
rect 11956 4336 12014 4382
rect 12060 4336 12118 4382
rect 12164 4336 12222 4382
rect 12268 4336 12326 4382
rect 12372 4336 12430 4382
rect 12476 4336 12534 4382
rect 12580 4336 12638 4382
rect 12684 4336 12742 4382
rect 12788 4336 12846 4382
rect 12892 4336 12950 4382
rect 12996 4336 13054 4382
rect 13100 4336 13158 4382
rect 13204 4336 13262 4382
rect 13308 4336 13366 4382
rect 13412 4336 13470 4382
rect 13516 4336 13574 4382
rect 13620 4336 13631 4382
rect 540 4321 13631 4336
rect 13258 3821 13326 3956
rect 355 3534 423 3682
rect 13258 3263 13326 3398
rect 355 2975 423 3123
rect 13258 2705 13326 2840
rect 355 2415 423 2563
rect 13258 2141 13326 2276
rect 355 1856 423 2004
rect 13258 1581 13326 1716
rect 355 1307 423 1455
rect 13258 1027 13326 1162
rect 355 657 423 1027
rect 13563 657 13631 4321
rect 43 581 13631 657
use M1_NWELL_CDNS_40661953145127  M1_NWELL_CDNS_40661953145127_0
timestamp 1713338890
transform 0 -1 6837 -1 0 619
box -128 -6888 128 6888
use M1_NWELL_CDNS_40661953145128  M1_NWELL_CDNS_40661953145128_0
timestamp 1713338890
transform 1 0 77 0 -1 2489
box -128 -1844 128 1844
use M1_NWELL_CDNS_40661953145128  M1_NWELL_CDNS_40661953145128_1
timestamp 1713338890
transform 1 0 13597 0 -1 2489
box -128 -1844 128 1844
use M1_PSUB_CDNS_69033583165350  M1_PSUB_CDNS_69033583165350_0
timestamp 1713338890
transform 0 -1 6837 1 0 4852
box -102 -5004 102 5004
use M1_PSUB_CDNS_69033583165350  M1_PSUB_CDNS_69033583165350_1
timestamp 1713338890
transform 0 -1 6837 1 0 10845
box -102 -5004 102 5004
use M1_PSUB_CDNS_69033583165350  M1_PSUB_CDNS_69033583165350_2
timestamp 1713338890
transform 0 -1 6837 1 0 16936
box -102 -5004 102 5004
use M1_PSUB_CDNS_69033583165351  M1_PSUB_CDNS_69033583165351_0
timestamp 1713338890
transform 1 0 12007 0 1 10894
box -102 -6144 102 6144
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_0
timestamp 1713338890
transform 1 0 9488 0 -1 10339
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_1
timestamp 1713338890
transform 1 0 7052 0 -1 10339
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_2
timestamp 1713338890
transform 1 0 4616 0 -1 10339
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_3
timestamp 1713338890
transform 1 0 2180 0 -1 10339
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_4
timestamp 1713338890
transform 1 0 4616 0 1 11351
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_5
timestamp 1713338890
transform 1 0 7052 0 1 11351
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_6
timestamp 1713338890
transform 1 0 9488 0 1 11351
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_7
timestamp 1713338890
transform 1 0 2180 0 1 11351
box -218 -350 2218 5092
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_0
timestamp 1713338890
transform 1 0 353 0 1 1429
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_1
timestamp 1713338890
transform 1 0 353 0 1 1989
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_2
timestamp 1713338890
transform 1 0 353 0 1 2549
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_3
timestamp 1713338890
transform 1 0 353 0 -1 1029
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_4
timestamp 1713338890
transform -1 0 13328 0 1 2269
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_5
timestamp 1713338890
transform -1 0 13328 0 1 1709
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_6
timestamp 1713338890
transform -1 0 13328 0 1 1149
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_7
timestamp 1713338890
transform 1 0 353 0 1 3109
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_8
timestamp 1713338890
transform 1 0 353 0 1 3669
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_9
timestamp 1713338890
transform -1 0 13328 0 1 2829
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_10
timestamp 1713338890
transform -1 0 13328 0 1 3389
box 0 0 12975 160
use ppolyf_u_CDNS_406619531453  ppolyf_u_CDNS_406619531453_11
timestamp 1713338890
transform -1 0 13328 0 1 3949
box 0 0 12975 160
<< labels >>
rlabel metal1 s 6835 10844 6835 10844 4 VMINUS
port 1 nsew
rlabel metal1 s 475 619 475 619 4 VPLUS
port 2 nsew
rlabel metal1 s 984 16493 984 16493 4 VRC
port 3 nsew
<< end >>
