magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2208 -2120 2592 2720
<< nwell >>
rect -208 -120 592 720
<< mvpmos >>
rect 0 0 140 600
rect 244 0 384 600
<< mvpdiff >>
rect -88 587 0 600
rect -88 541 -75 587
rect -29 541 0 587
rect -88 482 0 541
rect -88 436 -75 482
rect -29 436 0 482
rect -88 377 0 436
rect -88 331 -75 377
rect -29 331 0 377
rect -88 271 0 331
rect -88 225 -75 271
rect -29 225 0 271
rect -88 165 0 225
rect -88 119 -75 165
rect -29 119 0 165
rect -88 59 0 119
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 587 244 600
rect 140 541 169 587
rect 215 541 244 587
rect 140 482 244 541
rect 140 436 169 482
rect 215 436 244 482
rect 140 377 244 436
rect 140 331 169 377
rect 215 331 244 377
rect 140 271 244 331
rect 140 225 169 271
rect 215 225 244 271
rect 140 165 244 225
rect 140 119 169 165
rect 215 119 244 165
rect 140 59 244 119
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 587 472 600
rect 384 541 413 587
rect 459 541 472 587
rect 384 482 472 541
rect 384 436 413 482
rect 459 436 472 482
rect 384 377 472 436
rect 384 331 413 377
rect 459 331 472 377
rect 384 271 472 331
rect 384 225 413 271
rect 459 225 472 271
rect 384 165 472 225
rect 384 119 413 165
rect 459 119 472 165
rect 384 59 472 119
rect 384 13 413 59
rect 459 13 472 59
rect 384 0 472 13
<< mvpdiffc >>
rect -75 541 -29 587
rect -75 436 -29 482
rect -75 331 -29 377
rect -75 225 -29 271
rect -75 119 -29 165
rect -75 13 -29 59
rect 169 541 215 587
rect 169 436 215 482
rect 169 331 215 377
rect 169 225 215 271
rect 169 119 215 165
rect 169 13 215 59
rect 413 541 459 587
rect 413 436 459 482
rect 413 331 459 377
rect 413 225 459 271
rect 413 119 459 165
rect 413 13 459 59
<< polysilicon >>
rect 0 600 140 644
rect 244 600 384 644
rect 0 -44 140 0
rect 244 -44 384 0
<< metal1 >>
rect -75 587 -29 600
rect -75 482 -29 541
rect -75 377 -29 436
rect -75 271 -29 331
rect -75 165 -29 225
rect -75 59 -29 119
rect -75 0 -29 13
rect 169 587 215 600
rect 169 482 215 541
rect 169 377 215 436
rect 169 271 215 331
rect 169 165 215 225
rect 169 59 215 119
rect 169 0 215 13
rect 413 587 459 600
rect 413 482 459 541
rect 413 377 459 436
rect 413 271 459 331
rect 413 165 459 225
rect 413 59 459 119
rect 413 0 459 13
<< labels >>
rlabel metal1 192 300 192 300 4 D
rlabel metal1 436 300 436 300 4 S
rlabel metal1 -52 300 -52 300 4 S
<< end >>
