magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2102 -5864 2102 5864
<< psubdiff >>
rect -102 3842 102 3864
rect -102 3796 -80 3842
rect -34 3796 34 3842
rect 80 3796 102 3842
rect -102 3728 102 3796
rect -102 3682 -80 3728
rect -34 3682 34 3728
rect 80 3682 102 3728
rect -102 3614 102 3682
rect -102 3568 -80 3614
rect -34 3568 34 3614
rect 80 3568 102 3614
rect -102 3500 102 3568
rect -102 3454 -80 3500
rect -34 3454 34 3500
rect 80 3454 102 3500
rect -102 3386 102 3454
rect -102 3340 -80 3386
rect -34 3340 34 3386
rect 80 3340 102 3386
rect -102 3272 102 3340
rect -102 3226 -80 3272
rect -34 3226 34 3272
rect 80 3226 102 3272
rect -102 3158 102 3226
rect -102 3112 -80 3158
rect -34 3112 34 3158
rect 80 3112 102 3158
rect -102 3044 102 3112
rect -102 2998 -80 3044
rect -34 2998 34 3044
rect 80 2998 102 3044
rect -102 2930 102 2998
rect -102 2884 -80 2930
rect -34 2884 34 2930
rect 80 2884 102 2930
rect -102 2816 102 2884
rect -102 2770 -80 2816
rect -34 2770 34 2816
rect 80 2770 102 2816
rect -102 2702 102 2770
rect -102 2656 -80 2702
rect -34 2656 34 2702
rect 80 2656 102 2702
rect -102 2588 102 2656
rect -102 2542 -80 2588
rect -34 2542 34 2588
rect 80 2542 102 2588
rect -102 2474 102 2542
rect -102 2428 -80 2474
rect -34 2428 34 2474
rect 80 2428 102 2474
rect -102 2360 102 2428
rect -102 2314 -80 2360
rect -34 2314 34 2360
rect 80 2314 102 2360
rect -102 2246 102 2314
rect -102 2200 -80 2246
rect -34 2200 34 2246
rect 80 2200 102 2246
rect -102 2132 102 2200
rect -102 2086 -80 2132
rect -34 2086 34 2132
rect 80 2086 102 2132
rect -102 2018 102 2086
rect -102 1972 -80 2018
rect -34 1972 34 2018
rect 80 1972 102 2018
rect -102 1904 102 1972
rect -102 1858 -80 1904
rect -34 1858 34 1904
rect 80 1858 102 1904
rect -102 1790 102 1858
rect -102 1744 -80 1790
rect -34 1744 34 1790
rect 80 1744 102 1790
rect -102 1676 102 1744
rect -102 1630 -80 1676
rect -34 1630 34 1676
rect 80 1630 102 1676
rect -102 1562 102 1630
rect -102 1516 -80 1562
rect -34 1516 34 1562
rect 80 1516 102 1562
rect -102 1448 102 1516
rect -102 1402 -80 1448
rect -34 1402 34 1448
rect 80 1402 102 1448
rect -102 1334 102 1402
rect -102 1288 -80 1334
rect -34 1288 34 1334
rect 80 1288 102 1334
rect -102 1220 102 1288
rect -102 1174 -80 1220
rect -34 1174 34 1220
rect 80 1174 102 1220
rect -102 1106 102 1174
rect -102 1060 -80 1106
rect -34 1060 34 1106
rect 80 1060 102 1106
rect -102 992 102 1060
rect -102 946 -80 992
rect -34 946 34 992
rect 80 946 102 992
rect -102 878 102 946
rect -102 832 -80 878
rect -34 832 34 878
rect 80 832 102 878
rect -102 764 102 832
rect -102 718 -80 764
rect -34 718 34 764
rect 80 718 102 764
rect -102 650 102 718
rect -102 604 -80 650
rect -34 604 34 650
rect 80 604 102 650
rect -102 536 102 604
rect -102 490 -80 536
rect -34 490 34 536
rect 80 490 102 536
rect -102 422 102 490
rect -102 376 -80 422
rect -34 376 34 422
rect 80 376 102 422
rect -102 308 102 376
rect -102 262 -80 308
rect -34 262 34 308
rect 80 262 102 308
rect -102 194 102 262
rect -102 148 -80 194
rect -34 148 34 194
rect 80 148 102 194
rect -102 80 102 148
rect -102 34 -80 80
rect -34 34 34 80
rect 80 34 102 80
rect -102 -34 102 34
rect -102 -80 -80 -34
rect -34 -80 34 -34
rect 80 -80 102 -34
rect -102 -148 102 -80
rect -102 -194 -80 -148
rect -34 -194 34 -148
rect 80 -194 102 -148
rect -102 -262 102 -194
rect -102 -308 -80 -262
rect -34 -308 34 -262
rect 80 -308 102 -262
rect -102 -376 102 -308
rect -102 -422 -80 -376
rect -34 -422 34 -376
rect 80 -422 102 -376
rect -102 -490 102 -422
rect -102 -536 -80 -490
rect -34 -536 34 -490
rect 80 -536 102 -490
rect -102 -604 102 -536
rect -102 -650 -80 -604
rect -34 -650 34 -604
rect 80 -650 102 -604
rect -102 -718 102 -650
rect -102 -764 -80 -718
rect -34 -764 34 -718
rect 80 -764 102 -718
rect -102 -832 102 -764
rect -102 -878 -80 -832
rect -34 -878 34 -832
rect 80 -878 102 -832
rect -102 -946 102 -878
rect -102 -992 -80 -946
rect -34 -992 34 -946
rect 80 -992 102 -946
rect -102 -1060 102 -992
rect -102 -1106 -80 -1060
rect -34 -1106 34 -1060
rect 80 -1106 102 -1060
rect -102 -1174 102 -1106
rect -102 -1220 -80 -1174
rect -34 -1220 34 -1174
rect 80 -1220 102 -1174
rect -102 -1288 102 -1220
rect -102 -1334 -80 -1288
rect -34 -1334 34 -1288
rect 80 -1334 102 -1288
rect -102 -1402 102 -1334
rect -102 -1448 -80 -1402
rect -34 -1448 34 -1402
rect 80 -1448 102 -1402
rect -102 -1516 102 -1448
rect -102 -1562 -80 -1516
rect -34 -1562 34 -1516
rect 80 -1562 102 -1516
rect -102 -1630 102 -1562
rect -102 -1676 -80 -1630
rect -34 -1676 34 -1630
rect 80 -1676 102 -1630
rect -102 -1744 102 -1676
rect -102 -1790 -80 -1744
rect -34 -1790 34 -1744
rect 80 -1790 102 -1744
rect -102 -1858 102 -1790
rect -102 -1904 -80 -1858
rect -34 -1904 34 -1858
rect 80 -1904 102 -1858
rect -102 -1972 102 -1904
rect -102 -2018 -80 -1972
rect -34 -2018 34 -1972
rect 80 -2018 102 -1972
rect -102 -2086 102 -2018
rect -102 -2132 -80 -2086
rect -34 -2132 34 -2086
rect 80 -2132 102 -2086
rect -102 -2200 102 -2132
rect -102 -2246 -80 -2200
rect -34 -2246 34 -2200
rect 80 -2246 102 -2200
rect -102 -2314 102 -2246
rect -102 -2360 -80 -2314
rect -34 -2360 34 -2314
rect 80 -2360 102 -2314
rect -102 -2428 102 -2360
rect -102 -2474 -80 -2428
rect -34 -2474 34 -2428
rect 80 -2474 102 -2428
rect -102 -2542 102 -2474
rect -102 -2588 -80 -2542
rect -34 -2588 34 -2542
rect 80 -2588 102 -2542
rect -102 -2656 102 -2588
rect -102 -2702 -80 -2656
rect -34 -2702 34 -2656
rect 80 -2702 102 -2656
rect -102 -2770 102 -2702
rect -102 -2816 -80 -2770
rect -34 -2816 34 -2770
rect 80 -2816 102 -2770
rect -102 -2884 102 -2816
rect -102 -2930 -80 -2884
rect -34 -2930 34 -2884
rect 80 -2930 102 -2884
rect -102 -2998 102 -2930
rect -102 -3044 -80 -2998
rect -34 -3044 34 -2998
rect 80 -3044 102 -2998
rect -102 -3112 102 -3044
rect -102 -3158 -80 -3112
rect -34 -3158 34 -3112
rect 80 -3158 102 -3112
rect -102 -3226 102 -3158
rect -102 -3272 -80 -3226
rect -34 -3272 34 -3226
rect 80 -3272 102 -3226
rect -102 -3340 102 -3272
rect -102 -3386 -80 -3340
rect -34 -3386 34 -3340
rect 80 -3386 102 -3340
rect -102 -3454 102 -3386
rect -102 -3500 -80 -3454
rect -34 -3500 34 -3454
rect 80 -3500 102 -3454
rect -102 -3568 102 -3500
rect -102 -3614 -80 -3568
rect -34 -3614 34 -3568
rect 80 -3614 102 -3568
rect -102 -3682 102 -3614
rect -102 -3728 -80 -3682
rect -34 -3728 34 -3682
rect 80 -3728 102 -3682
rect -102 -3796 102 -3728
rect -102 -3842 -80 -3796
rect -34 -3842 34 -3796
rect 80 -3842 102 -3796
rect -102 -3864 102 -3842
<< psubdiffcont >>
rect -80 3796 -34 3842
rect 34 3796 80 3842
rect -80 3682 -34 3728
rect 34 3682 80 3728
rect -80 3568 -34 3614
rect 34 3568 80 3614
rect -80 3454 -34 3500
rect 34 3454 80 3500
rect -80 3340 -34 3386
rect 34 3340 80 3386
rect -80 3226 -34 3272
rect 34 3226 80 3272
rect -80 3112 -34 3158
rect 34 3112 80 3158
rect -80 2998 -34 3044
rect 34 2998 80 3044
rect -80 2884 -34 2930
rect 34 2884 80 2930
rect -80 2770 -34 2816
rect 34 2770 80 2816
rect -80 2656 -34 2702
rect 34 2656 80 2702
rect -80 2542 -34 2588
rect 34 2542 80 2588
rect -80 2428 -34 2474
rect 34 2428 80 2474
rect -80 2314 -34 2360
rect 34 2314 80 2360
rect -80 2200 -34 2246
rect 34 2200 80 2246
rect -80 2086 -34 2132
rect 34 2086 80 2132
rect -80 1972 -34 2018
rect 34 1972 80 2018
rect -80 1858 -34 1904
rect 34 1858 80 1904
rect -80 1744 -34 1790
rect 34 1744 80 1790
rect -80 1630 -34 1676
rect 34 1630 80 1676
rect -80 1516 -34 1562
rect 34 1516 80 1562
rect -80 1402 -34 1448
rect 34 1402 80 1448
rect -80 1288 -34 1334
rect 34 1288 80 1334
rect -80 1174 -34 1220
rect 34 1174 80 1220
rect -80 1060 -34 1106
rect 34 1060 80 1106
rect -80 946 -34 992
rect 34 946 80 992
rect -80 832 -34 878
rect 34 832 80 878
rect -80 718 -34 764
rect 34 718 80 764
rect -80 604 -34 650
rect 34 604 80 650
rect -80 490 -34 536
rect 34 490 80 536
rect -80 376 -34 422
rect 34 376 80 422
rect -80 262 -34 308
rect 34 262 80 308
rect -80 148 -34 194
rect 34 148 80 194
rect -80 34 -34 80
rect 34 34 80 80
rect -80 -80 -34 -34
rect 34 -80 80 -34
rect -80 -194 -34 -148
rect 34 -194 80 -148
rect -80 -308 -34 -262
rect 34 -308 80 -262
rect -80 -422 -34 -376
rect 34 -422 80 -376
rect -80 -536 -34 -490
rect 34 -536 80 -490
rect -80 -650 -34 -604
rect 34 -650 80 -604
rect -80 -764 -34 -718
rect 34 -764 80 -718
rect -80 -878 -34 -832
rect 34 -878 80 -832
rect -80 -992 -34 -946
rect 34 -992 80 -946
rect -80 -1106 -34 -1060
rect 34 -1106 80 -1060
rect -80 -1220 -34 -1174
rect 34 -1220 80 -1174
rect -80 -1334 -34 -1288
rect 34 -1334 80 -1288
rect -80 -1448 -34 -1402
rect 34 -1448 80 -1402
rect -80 -1562 -34 -1516
rect 34 -1562 80 -1516
rect -80 -1676 -34 -1630
rect 34 -1676 80 -1630
rect -80 -1790 -34 -1744
rect 34 -1790 80 -1744
rect -80 -1904 -34 -1858
rect 34 -1904 80 -1858
rect -80 -2018 -34 -1972
rect 34 -2018 80 -1972
rect -80 -2132 -34 -2086
rect 34 -2132 80 -2086
rect -80 -2246 -34 -2200
rect 34 -2246 80 -2200
rect -80 -2360 -34 -2314
rect 34 -2360 80 -2314
rect -80 -2474 -34 -2428
rect 34 -2474 80 -2428
rect -80 -2588 -34 -2542
rect 34 -2588 80 -2542
rect -80 -2702 -34 -2656
rect 34 -2702 80 -2656
rect -80 -2816 -34 -2770
rect 34 -2816 80 -2770
rect -80 -2930 -34 -2884
rect 34 -2930 80 -2884
rect -80 -3044 -34 -2998
rect 34 -3044 80 -2998
rect -80 -3158 -34 -3112
rect 34 -3158 80 -3112
rect -80 -3272 -34 -3226
rect 34 -3272 80 -3226
rect -80 -3386 -34 -3340
rect 34 -3386 80 -3340
rect -80 -3500 -34 -3454
rect 34 -3500 80 -3454
rect -80 -3614 -34 -3568
rect 34 -3614 80 -3568
rect -80 -3728 -34 -3682
rect 34 -3728 80 -3682
rect -80 -3842 -34 -3796
rect 34 -3842 80 -3796
<< metal1 >>
rect -91 3842 91 3853
rect -91 3796 -80 3842
rect -34 3796 34 3842
rect 80 3796 91 3842
rect -91 3728 91 3796
rect -91 3682 -80 3728
rect -34 3682 34 3728
rect 80 3682 91 3728
rect -91 3614 91 3682
rect -91 3568 -80 3614
rect -34 3568 34 3614
rect 80 3568 91 3614
rect -91 3500 91 3568
rect -91 3454 -80 3500
rect -34 3454 34 3500
rect 80 3454 91 3500
rect -91 3386 91 3454
rect -91 3340 -80 3386
rect -34 3340 34 3386
rect 80 3340 91 3386
rect -91 3272 91 3340
rect -91 3226 -80 3272
rect -34 3226 34 3272
rect 80 3226 91 3272
rect -91 3158 91 3226
rect -91 3112 -80 3158
rect -34 3112 34 3158
rect 80 3112 91 3158
rect -91 3044 91 3112
rect -91 2998 -80 3044
rect -34 2998 34 3044
rect 80 2998 91 3044
rect -91 2930 91 2998
rect -91 2884 -80 2930
rect -34 2884 34 2930
rect 80 2884 91 2930
rect -91 2816 91 2884
rect -91 2770 -80 2816
rect -34 2770 34 2816
rect 80 2770 91 2816
rect -91 2702 91 2770
rect -91 2656 -80 2702
rect -34 2656 34 2702
rect 80 2656 91 2702
rect -91 2588 91 2656
rect -91 2542 -80 2588
rect -34 2542 34 2588
rect 80 2542 91 2588
rect -91 2474 91 2542
rect -91 2428 -80 2474
rect -34 2428 34 2474
rect 80 2428 91 2474
rect -91 2360 91 2428
rect -91 2314 -80 2360
rect -34 2314 34 2360
rect 80 2314 91 2360
rect -91 2246 91 2314
rect -91 2200 -80 2246
rect -34 2200 34 2246
rect 80 2200 91 2246
rect -91 2132 91 2200
rect -91 2086 -80 2132
rect -34 2086 34 2132
rect 80 2086 91 2132
rect -91 2018 91 2086
rect -91 1972 -80 2018
rect -34 1972 34 2018
rect 80 1972 91 2018
rect -91 1904 91 1972
rect -91 1858 -80 1904
rect -34 1858 34 1904
rect 80 1858 91 1904
rect -91 1790 91 1858
rect -91 1744 -80 1790
rect -34 1744 34 1790
rect 80 1744 91 1790
rect -91 1676 91 1744
rect -91 1630 -80 1676
rect -34 1630 34 1676
rect 80 1630 91 1676
rect -91 1562 91 1630
rect -91 1516 -80 1562
rect -34 1516 34 1562
rect 80 1516 91 1562
rect -91 1448 91 1516
rect -91 1402 -80 1448
rect -34 1402 34 1448
rect 80 1402 91 1448
rect -91 1334 91 1402
rect -91 1288 -80 1334
rect -34 1288 34 1334
rect 80 1288 91 1334
rect -91 1220 91 1288
rect -91 1174 -80 1220
rect -34 1174 34 1220
rect 80 1174 91 1220
rect -91 1106 91 1174
rect -91 1060 -80 1106
rect -34 1060 34 1106
rect 80 1060 91 1106
rect -91 992 91 1060
rect -91 946 -80 992
rect -34 946 34 992
rect 80 946 91 992
rect -91 878 91 946
rect -91 832 -80 878
rect -34 832 34 878
rect 80 832 91 878
rect -91 764 91 832
rect -91 718 -80 764
rect -34 718 34 764
rect 80 718 91 764
rect -91 650 91 718
rect -91 604 -80 650
rect -34 604 34 650
rect 80 604 91 650
rect -91 536 91 604
rect -91 490 -80 536
rect -34 490 34 536
rect 80 490 91 536
rect -91 422 91 490
rect -91 376 -80 422
rect -34 376 34 422
rect 80 376 91 422
rect -91 308 91 376
rect -91 262 -80 308
rect -34 262 34 308
rect 80 262 91 308
rect -91 194 91 262
rect -91 148 -80 194
rect -34 148 34 194
rect 80 148 91 194
rect -91 80 91 148
rect -91 34 -80 80
rect -34 34 34 80
rect 80 34 91 80
rect -91 -34 91 34
rect -91 -80 -80 -34
rect -34 -80 34 -34
rect 80 -80 91 -34
rect -91 -148 91 -80
rect -91 -194 -80 -148
rect -34 -194 34 -148
rect 80 -194 91 -148
rect -91 -262 91 -194
rect -91 -308 -80 -262
rect -34 -308 34 -262
rect 80 -308 91 -262
rect -91 -376 91 -308
rect -91 -422 -80 -376
rect -34 -422 34 -376
rect 80 -422 91 -376
rect -91 -490 91 -422
rect -91 -536 -80 -490
rect -34 -536 34 -490
rect 80 -536 91 -490
rect -91 -604 91 -536
rect -91 -650 -80 -604
rect -34 -650 34 -604
rect 80 -650 91 -604
rect -91 -718 91 -650
rect -91 -764 -80 -718
rect -34 -764 34 -718
rect 80 -764 91 -718
rect -91 -832 91 -764
rect -91 -878 -80 -832
rect -34 -878 34 -832
rect 80 -878 91 -832
rect -91 -946 91 -878
rect -91 -992 -80 -946
rect -34 -992 34 -946
rect 80 -992 91 -946
rect -91 -1060 91 -992
rect -91 -1106 -80 -1060
rect -34 -1106 34 -1060
rect 80 -1106 91 -1060
rect -91 -1174 91 -1106
rect -91 -1220 -80 -1174
rect -34 -1220 34 -1174
rect 80 -1220 91 -1174
rect -91 -1288 91 -1220
rect -91 -1334 -80 -1288
rect -34 -1334 34 -1288
rect 80 -1334 91 -1288
rect -91 -1402 91 -1334
rect -91 -1448 -80 -1402
rect -34 -1448 34 -1402
rect 80 -1448 91 -1402
rect -91 -1516 91 -1448
rect -91 -1562 -80 -1516
rect -34 -1562 34 -1516
rect 80 -1562 91 -1516
rect -91 -1630 91 -1562
rect -91 -1676 -80 -1630
rect -34 -1676 34 -1630
rect 80 -1676 91 -1630
rect -91 -1744 91 -1676
rect -91 -1790 -80 -1744
rect -34 -1790 34 -1744
rect 80 -1790 91 -1744
rect -91 -1858 91 -1790
rect -91 -1904 -80 -1858
rect -34 -1904 34 -1858
rect 80 -1904 91 -1858
rect -91 -1972 91 -1904
rect -91 -2018 -80 -1972
rect -34 -2018 34 -1972
rect 80 -2018 91 -1972
rect -91 -2086 91 -2018
rect -91 -2132 -80 -2086
rect -34 -2132 34 -2086
rect 80 -2132 91 -2086
rect -91 -2200 91 -2132
rect -91 -2246 -80 -2200
rect -34 -2246 34 -2200
rect 80 -2246 91 -2200
rect -91 -2314 91 -2246
rect -91 -2360 -80 -2314
rect -34 -2360 34 -2314
rect 80 -2360 91 -2314
rect -91 -2428 91 -2360
rect -91 -2474 -80 -2428
rect -34 -2474 34 -2428
rect 80 -2474 91 -2428
rect -91 -2542 91 -2474
rect -91 -2588 -80 -2542
rect -34 -2588 34 -2542
rect 80 -2588 91 -2542
rect -91 -2656 91 -2588
rect -91 -2702 -80 -2656
rect -34 -2702 34 -2656
rect 80 -2702 91 -2656
rect -91 -2770 91 -2702
rect -91 -2816 -80 -2770
rect -34 -2816 34 -2770
rect 80 -2816 91 -2770
rect -91 -2884 91 -2816
rect -91 -2930 -80 -2884
rect -34 -2930 34 -2884
rect 80 -2930 91 -2884
rect -91 -2998 91 -2930
rect -91 -3044 -80 -2998
rect -34 -3044 34 -2998
rect 80 -3044 91 -2998
rect -91 -3112 91 -3044
rect -91 -3158 -80 -3112
rect -34 -3158 34 -3112
rect 80 -3158 91 -3112
rect -91 -3226 91 -3158
rect -91 -3272 -80 -3226
rect -34 -3272 34 -3226
rect 80 -3272 91 -3226
rect -91 -3340 91 -3272
rect -91 -3386 -80 -3340
rect -34 -3386 34 -3340
rect 80 -3386 91 -3340
rect -91 -3454 91 -3386
rect -91 -3500 -80 -3454
rect -34 -3500 34 -3454
rect 80 -3500 91 -3454
rect -91 -3568 91 -3500
rect -91 -3614 -80 -3568
rect -34 -3614 34 -3568
rect 80 -3614 91 -3568
rect -91 -3682 91 -3614
rect -91 -3728 -80 -3682
rect -34 -3728 34 -3682
rect 80 -3728 91 -3682
rect -91 -3796 91 -3728
rect -91 -3842 -80 -3796
rect -34 -3842 34 -3796
rect 80 -3842 91 -3796
rect -91 -3853 91 -3842
<< end >>
