magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1484 -1050 1484 1050
<< metal1 >>
rect -484 44 484 50
rect -484 18 -478 44
rect -452 18 -416 44
rect -390 18 -354 44
rect -328 18 -292 44
rect -266 18 -230 44
rect -204 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 204 44
rect 230 18 266 44
rect 292 18 328 44
rect 354 18 390 44
rect 416 18 452 44
rect 478 18 484 44
rect -484 -18 484 18
rect -484 -44 -478 -18
rect -452 -44 -416 -18
rect -390 -44 -354 -18
rect -328 -44 -292 -18
rect -266 -44 -230 -18
rect -204 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 204 -18
rect 230 -44 266 -18
rect 292 -44 328 -18
rect 354 -44 390 -18
rect 416 -44 452 -18
rect 478 -44 484 -18
rect -484 -50 484 -44
<< via1 >>
rect -478 18 -452 44
rect -416 18 -390 44
rect -354 18 -328 44
rect -292 18 -266 44
rect -230 18 -204 44
rect -168 18 -142 44
rect -106 18 -80 44
rect -44 18 -18 44
rect 18 18 44 44
rect 80 18 106 44
rect 142 18 168 44
rect 204 18 230 44
rect 266 18 292 44
rect 328 18 354 44
rect 390 18 416 44
rect 452 18 478 44
rect -478 -44 -452 -18
rect -416 -44 -390 -18
rect -354 -44 -328 -18
rect -292 -44 -266 -18
rect -230 -44 -204 -18
rect -168 -44 -142 -18
rect -106 -44 -80 -18
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect 80 -44 106 -18
rect 142 -44 168 -18
rect 204 -44 230 -18
rect 266 -44 292 -18
rect 328 -44 354 -18
rect 390 -44 416 -18
rect 452 -44 478 -18
<< metal2 >>
rect -484 44 484 50
rect -484 18 -478 44
rect -452 18 -416 44
rect -390 18 -354 44
rect -328 18 -292 44
rect -266 18 -230 44
rect -204 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 204 44
rect 230 18 266 44
rect 292 18 328 44
rect 354 18 390 44
rect 416 18 452 44
rect 478 18 484 44
rect -484 -18 484 18
rect -484 -44 -478 -18
rect -452 -44 -416 -18
rect -390 -44 -354 -18
rect -328 -44 -292 -18
rect -266 -44 -230 -18
rect -204 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 204 -18
rect 230 -44 266 -18
rect 292 -44 328 -18
rect 354 -44 390 -18
rect 416 -44 452 -18
rect 478 -44 484 -18
rect -484 -50 484 -44
<< end >>
