magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1361 -1019 1361 1019
<< metal1 >>
rect -361 13 361 19
rect -361 -13 -355 13
rect -329 -13 -279 13
rect -253 -13 -203 13
rect -177 -13 -127 13
rect -101 -13 -51 13
rect -25 -13 25 13
rect 51 -13 101 13
rect 127 -13 177 13
rect 203 -13 253 13
rect 279 -13 329 13
rect 355 -13 361 13
rect -361 -19 361 -13
<< via1 >>
rect -355 -13 -329 13
rect -279 -13 -253 13
rect -203 -13 -177 13
rect -127 -13 -101 13
rect -51 -13 -25 13
rect 25 -13 51 13
rect 101 -13 127 13
rect 177 -13 203 13
rect 253 -13 279 13
rect 329 -13 355 13
<< metal2 >>
rect -361 13 361 19
rect -361 -13 -355 13
rect -329 -13 -279 13
rect -253 -13 -203 13
rect -177 -13 -127 13
rect -101 -13 -51 13
rect -25 -13 25 13
rect 51 -13 101 13
rect 127 -13 177 13
rect 203 -13 253 13
rect 279 -13 329 13
rect 355 -13 361 13
rect -361 -19 361 -13
<< end >>
