magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1513 -1019 1513 1019
<< metal1 >>
rect -513 13 513 19
rect -513 -13 -507 13
rect 507 -13 513 13
rect -513 -19 513 -13
<< via1 >>
rect -507 -13 507 13
<< metal2 >>
rect -513 13 513 19
rect -513 -13 -507 13
rect 507 -13 513 13
rect -513 -19 513 -13
<< end >>
