magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -30281 -2097 30281 2097
<< psubdiff >>
rect -28281 75 28281 97
rect -28281 29 -28259 75
rect -28213 29 -28155 75
rect -28109 29 -28051 75
rect -28005 29 -27947 75
rect -27901 29 -27843 75
rect -27797 29 -27739 75
rect -27693 29 -27635 75
rect -27589 29 -27531 75
rect -27485 29 -27427 75
rect -27381 29 -27323 75
rect -27277 29 -27219 75
rect -27173 29 -27115 75
rect -27069 29 -27011 75
rect -26965 29 -26907 75
rect -26861 29 -26803 75
rect -26757 29 -26699 75
rect -26653 29 -26595 75
rect -26549 29 -26491 75
rect -26445 29 -26387 75
rect -26341 29 -26283 75
rect -26237 29 -26179 75
rect -26133 29 -26075 75
rect -26029 29 -25971 75
rect -25925 29 -25867 75
rect -25821 29 -25763 75
rect -25717 29 -25659 75
rect -25613 29 -25555 75
rect -25509 29 -25451 75
rect -25405 29 -25347 75
rect -25301 29 -25243 75
rect -25197 29 -25139 75
rect -25093 29 -25035 75
rect -24989 29 -24931 75
rect -24885 29 -24827 75
rect -24781 29 -24723 75
rect -24677 29 -24619 75
rect -24573 29 -24515 75
rect -24469 29 -24411 75
rect -24365 29 -24307 75
rect -24261 29 -24203 75
rect -24157 29 -24099 75
rect -24053 29 -23995 75
rect -23949 29 -23891 75
rect -23845 29 -23787 75
rect -23741 29 -23683 75
rect -23637 29 -23579 75
rect -23533 29 -23475 75
rect -23429 29 -23371 75
rect -23325 29 -23267 75
rect -23221 29 -23163 75
rect -23117 29 -23059 75
rect -23013 29 -22955 75
rect -22909 29 -22851 75
rect -22805 29 -22747 75
rect -22701 29 -22643 75
rect -22597 29 -22539 75
rect -22493 29 -22435 75
rect -22389 29 -22331 75
rect -22285 29 -22227 75
rect -22181 29 -22123 75
rect -22077 29 -22019 75
rect -21973 29 -21915 75
rect -21869 29 -21811 75
rect -21765 29 -21707 75
rect -21661 29 -21603 75
rect -21557 29 -21499 75
rect -21453 29 -21395 75
rect -21349 29 -21291 75
rect -21245 29 -21187 75
rect -21141 29 -21083 75
rect -21037 29 -20979 75
rect -20933 29 -20875 75
rect -20829 29 -20771 75
rect -20725 29 -20667 75
rect -20621 29 -20563 75
rect -20517 29 -20459 75
rect -20413 29 -20355 75
rect -20309 29 -20251 75
rect -20205 29 -20147 75
rect -20101 29 -20043 75
rect -19997 29 -19939 75
rect -19893 29 -19835 75
rect -19789 29 -19731 75
rect -19685 29 -19627 75
rect -19581 29 -19523 75
rect -19477 29 -19419 75
rect -19373 29 -19315 75
rect -19269 29 -19211 75
rect -19165 29 -19107 75
rect -19061 29 -19003 75
rect -18957 29 -18899 75
rect -18853 29 -18795 75
rect -18749 29 -18691 75
rect -18645 29 -18587 75
rect -18541 29 -18483 75
rect -18437 29 -18379 75
rect -18333 29 -18275 75
rect -18229 29 -18171 75
rect -18125 29 -18067 75
rect -18021 29 -17963 75
rect -17917 29 -17859 75
rect -17813 29 -17755 75
rect -17709 29 -17651 75
rect -17605 29 -17547 75
rect -17501 29 -17443 75
rect -17397 29 -17339 75
rect -17293 29 -17235 75
rect -17189 29 -17131 75
rect -17085 29 -17027 75
rect -16981 29 -16923 75
rect -16877 29 -16819 75
rect -16773 29 -16715 75
rect -16669 29 -16611 75
rect -16565 29 -16507 75
rect -16461 29 -16403 75
rect -16357 29 -16299 75
rect -16253 29 -16195 75
rect -16149 29 -16091 75
rect -16045 29 -15987 75
rect -15941 29 -15883 75
rect -15837 29 -15779 75
rect -15733 29 -15675 75
rect -15629 29 -15571 75
rect -15525 29 -15467 75
rect -15421 29 -15363 75
rect -15317 29 -15259 75
rect -15213 29 -15155 75
rect -15109 29 -15051 75
rect -15005 29 -14947 75
rect -14901 29 -14843 75
rect -14797 29 -14739 75
rect -14693 29 -14635 75
rect -14589 29 -14531 75
rect -14485 29 -14427 75
rect -14381 29 -14323 75
rect -14277 29 -14219 75
rect -14173 29 -14115 75
rect -14069 29 -14011 75
rect -13965 29 -13907 75
rect -13861 29 -13803 75
rect -13757 29 -13699 75
rect -13653 29 -13595 75
rect -13549 29 -13491 75
rect -13445 29 -13387 75
rect -13341 29 -13283 75
rect -13237 29 -13179 75
rect -13133 29 -13075 75
rect -13029 29 -12971 75
rect -12925 29 -12867 75
rect -12821 29 -12763 75
rect -12717 29 -12659 75
rect -12613 29 -12555 75
rect -12509 29 -12451 75
rect -12405 29 -12347 75
rect -12301 29 -12243 75
rect -12197 29 -12139 75
rect -12093 29 -12035 75
rect -11989 29 -11931 75
rect -11885 29 -11827 75
rect -11781 29 -11723 75
rect -11677 29 -11619 75
rect -11573 29 -11515 75
rect -11469 29 -11411 75
rect -11365 29 -11307 75
rect -11261 29 -11203 75
rect -11157 29 -11099 75
rect -11053 29 -10995 75
rect -10949 29 -10891 75
rect -10845 29 -10787 75
rect -10741 29 -10683 75
rect -10637 29 -10579 75
rect -10533 29 -10475 75
rect -10429 29 -10371 75
rect -10325 29 -10267 75
rect -10221 29 -10163 75
rect -10117 29 -10059 75
rect -10013 29 -9955 75
rect -9909 29 -9851 75
rect -9805 29 -9747 75
rect -9701 29 -9643 75
rect -9597 29 -9539 75
rect -9493 29 -9435 75
rect -9389 29 -9331 75
rect -9285 29 -9227 75
rect -9181 29 -9123 75
rect -9077 29 -9019 75
rect -8973 29 -8915 75
rect -8869 29 -8811 75
rect -8765 29 -8707 75
rect -8661 29 -8603 75
rect -8557 29 -8499 75
rect -8453 29 -8395 75
rect -8349 29 -8291 75
rect -8245 29 -8187 75
rect -8141 29 -8083 75
rect -8037 29 -7979 75
rect -7933 29 -7875 75
rect -7829 29 -7771 75
rect -7725 29 -7667 75
rect -7621 29 -7563 75
rect -7517 29 -7459 75
rect -7413 29 -7355 75
rect -7309 29 -7251 75
rect -7205 29 -7147 75
rect -7101 29 -7043 75
rect -6997 29 -6939 75
rect -6893 29 -6835 75
rect -6789 29 -6731 75
rect -6685 29 -6627 75
rect -6581 29 -6523 75
rect -6477 29 -6419 75
rect -6373 29 -6315 75
rect -6269 29 -6211 75
rect -6165 29 -6107 75
rect -6061 29 -6003 75
rect -5957 29 -5899 75
rect -5853 29 -5795 75
rect -5749 29 -5691 75
rect -5645 29 -5587 75
rect -5541 29 -5483 75
rect -5437 29 -5379 75
rect -5333 29 -5275 75
rect -5229 29 -5171 75
rect -5125 29 -5067 75
rect -5021 29 -4963 75
rect -4917 29 -4859 75
rect -4813 29 -4755 75
rect -4709 29 -4651 75
rect -4605 29 -4547 75
rect -4501 29 -4443 75
rect -4397 29 -4339 75
rect -4293 29 -4235 75
rect -4189 29 -4131 75
rect -4085 29 -4027 75
rect -3981 29 -3923 75
rect -3877 29 -3819 75
rect -3773 29 -3715 75
rect -3669 29 -3611 75
rect -3565 29 -3507 75
rect -3461 29 -3403 75
rect -3357 29 -3299 75
rect -3253 29 -3195 75
rect -3149 29 -3091 75
rect -3045 29 -2987 75
rect -2941 29 -2883 75
rect -2837 29 -2779 75
rect -2733 29 -2675 75
rect -2629 29 -2571 75
rect -2525 29 -2467 75
rect -2421 29 -2363 75
rect -2317 29 -2259 75
rect -2213 29 -2155 75
rect -2109 29 -2051 75
rect -2005 29 -1947 75
rect -1901 29 -1843 75
rect -1797 29 -1739 75
rect -1693 29 -1635 75
rect -1589 29 -1531 75
rect -1485 29 -1427 75
rect -1381 29 -1323 75
rect -1277 29 -1219 75
rect -1173 29 -1115 75
rect -1069 29 -1011 75
rect -965 29 -907 75
rect -861 29 -803 75
rect -757 29 -699 75
rect -653 29 -595 75
rect -549 29 -491 75
rect -445 29 -387 75
rect -341 29 -283 75
rect -237 29 -179 75
rect -133 29 -75 75
rect -29 29 29 75
rect 75 29 133 75
rect 179 29 237 75
rect 283 29 341 75
rect 387 29 445 75
rect 491 29 549 75
rect 595 29 653 75
rect 699 29 757 75
rect 803 29 861 75
rect 907 29 965 75
rect 1011 29 1069 75
rect 1115 29 1173 75
rect 1219 29 1277 75
rect 1323 29 1381 75
rect 1427 29 1485 75
rect 1531 29 1589 75
rect 1635 29 1693 75
rect 1739 29 1797 75
rect 1843 29 1901 75
rect 1947 29 2005 75
rect 2051 29 2109 75
rect 2155 29 2213 75
rect 2259 29 2317 75
rect 2363 29 2421 75
rect 2467 29 2525 75
rect 2571 29 2629 75
rect 2675 29 2733 75
rect 2779 29 2837 75
rect 2883 29 2941 75
rect 2987 29 3045 75
rect 3091 29 3149 75
rect 3195 29 3253 75
rect 3299 29 3357 75
rect 3403 29 3461 75
rect 3507 29 3565 75
rect 3611 29 3669 75
rect 3715 29 3773 75
rect 3819 29 3877 75
rect 3923 29 3981 75
rect 4027 29 4085 75
rect 4131 29 4189 75
rect 4235 29 4293 75
rect 4339 29 4397 75
rect 4443 29 4501 75
rect 4547 29 4605 75
rect 4651 29 4709 75
rect 4755 29 4813 75
rect 4859 29 4917 75
rect 4963 29 5021 75
rect 5067 29 5125 75
rect 5171 29 5229 75
rect 5275 29 5333 75
rect 5379 29 5437 75
rect 5483 29 5541 75
rect 5587 29 5645 75
rect 5691 29 5749 75
rect 5795 29 5853 75
rect 5899 29 5957 75
rect 6003 29 6061 75
rect 6107 29 6165 75
rect 6211 29 6269 75
rect 6315 29 6373 75
rect 6419 29 6477 75
rect 6523 29 6581 75
rect 6627 29 6685 75
rect 6731 29 6789 75
rect 6835 29 6893 75
rect 6939 29 6997 75
rect 7043 29 7101 75
rect 7147 29 7205 75
rect 7251 29 7309 75
rect 7355 29 7413 75
rect 7459 29 7517 75
rect 7563 29 7621 75
rect 7667 29 7725 75
rect 7771 29 7829 75
rect 7875 29 7933 75
rect 7979 29 8037 75
rect 8083 29 8141 75
rect 8187 29 8245 75
rect 8291 29 8349 75
rect 8395 29 8453 75
rect 8499 29 8557 75
rect 8603 29 8661 75
rect 8707 29 8765 75
rect 8811 29 8869 75
rect 8915 29 8973 75
rect 9019 29 9077 75
rect 9123 29 9181 75
rect 9227 29 9285 75
rect 9331 29 9389 75
rect 9435 29 9493 75
rect 9539 29 9597 75
rect 9643 29 9701 75
rect 9747 29 9805 75
rect 9851 29 9909 75
rect 9955 29 10013 75
rect 10059 29 10117 75
rect 10163 29 10221 75
rect 10267 29 10325 75
rect 10371 29 10429 75
rect 10475 29 10533 75
rect 10579 29 10637 75
rect 10683 29 10741 75
rect 10787 29 10845 75
rect 10891 29 10949 75
rect 10995 29 11053 75
rect 11099 29 11157 75
rect 11203 29 11261 75
rect 11307 29 11365 75
rect 11411 29 11469 75
rect 11515 29 11573 75
rect 11619 29 11677 75
rect 11723 29 11781 75
rect 11827 29 11885 75
rect 11931 29 11989 75
rect 12035 29 12093 75
rect 12139 29 12197 75
rect 12243 29 12301 75
rect 12347 29 12405 75
rect 12451 29 12509 75
rect 12555 29 12613 75
rect 12659 29 12717 75
rect 12763 29 12821 75
rect 12867 29 12925 75
rect 12971 29 13029 75
rect 13075 29 13133 75
rect 13179 29 13237 75
rect 13283 29 13341 75
rect 13387 29 13445 75
rect 13491 29 13549 75
rect 13595 29 13653 75
rect 13699 29 13757 75
rect 13803 29 13861 75
rect 13907 29 13965 75
rect 14011 29 14069 75
rect 14115 29 14173 75
rect 14219 29 14277 75
rect 14323 29 14381 75
rect 14427 29 14485 75
rect 14531 29 14589 75
rect 14635 29 14693 75
rect 14739 29 14797 75
rect 14843 29 14901 75
rect 14947 29 15005 75
rect 15051 29 15109 75
rect 15155 29 15213 75
rect 15259 29 15317 75
rect 15363 29 15421 75
rect 15467 29 15525 75
rect 15571 29 15629 75
rect 15675 29 15733 75
rect 15779 29 15837 75
rect 15883 29 15941 75
rect 15987 29 16045 75
rect 16091 29 16149 75
rect 16195 29 16253 75
rect 16299 29 16357 75
rect 16403 29 16461 75
rect 16507 29 16565 75
rect 16611 29 16669 75
rect 16715 29 16773 75
rect 16819 29 16877 75
rect 16923 29 16981 75
rect 17027 29 17085 75
rect 17131 29 17189 75
rect 17235 29 17293 75
rect 17339 29 17397 75
rect 17443 29 17501 75
rect 17547 29 17605 75
rect 17651 29 17709 75
rect 17755 29 17813 75
rect 17859 29 17917 75
rect 17963 29 18021 75
rect 18067 29 18125 75
rect 18171 29 18229 75
rect 18275 29 18333 75
rect 18379 29 18437 75
rect 18483 29 18541 75
rect 18587 29 18645 75
rect 18691 29 18749 75
rect 18795 29 18853 75
rect 18899 29 18957 75
rect 19003 29 19061 75
rect 19107 29 19165 75
rect 19211 29 19269 75
rect 19315 29 19373 75
rect 19419 29 19477 75
rect 19523 29 19581 75
rect 19627 29 19685 75
rect 19731 29 19789 75
rect 19835 29 19893 75
rect 19939 29 19997 75
rect 20043 29 20101 75
rect 20147 29 20205 75
rect 20251 29 20309 75
rect 20355 29 20413 75
rect 20459 29 20517 75
rect 20563 29 20621 75
rect 20667 29 20725 75
rect 20771 29 20829 75
rect 20875 29 20933 75
rect 20979 29 21037 75
rect 21083 29 21141 75
rect 21187 29 21245 75
rect 21291 29 21349 75
rect 21395 29 21453 75
rect 21499 29 21557 75
rect 21603 29 21661 75
rect 21707 29 21765 75
rect 21811 29 21869 75
rect 21915 29 21973 75
rect 22019 29 22077 75
rect 22123 29 22181 75
rect 22227 29 22285 75
rect 22331 29 22389 75
rect 22435 29 22493 75
rect 22539 29 22597 75
rect 22643 29 22701 75
rect 22747 29 22805 75
rect 22851 29 22909 75
rect 22955 29 23013 75
rect 23059 29 23117 75
rect 23163 29 23221 75
rect 23267 29 23325 75
rect 23371 29 23429 75
rect 23475 29 23533 75
rect 23579 29 23637 75
rect 23683 29 23741 75
rect 23787 29 23845 75
rect 23891 29 23949 75
rect 23995 29 24053 75
rect 24099 29 24157 75
rect 24203 29 24261 75
rect 24307 29 24365 75
rect 24411 29 24469 75
rect 24515 29 24573 75
rect 24619 29 24677 75
rect 24723 29 24781 75
rect 24827 29 24885 75
rect 24931 29 24989 75
rect 25035 29 25093 75
rect 25139 29 25197 75
rect 25243 29 25301 75
rect 25347 29 25405 75
rect 25451 29 25509 75
rect 25555 29 25613 75
rect 25659 29 25717 75
rect 25763 29 25821 75
rect 25867 29 25925 75
rect 25971 29 26029 75
rect 26075 29 26133 75
rect 26179 29 26237 75
rect 26283 29 26341 75
rect 26387 29 26445 75
rect 26491 29 26549 75
rect 26595 29 26653 75
rect 26699 29 26757 75
rect 26803 29 26861 75
rect 26907 29 26965 75
rect 27011 29 27069 75
rect 27115 29 27173 75
rect 27219 29 27277 75
rect 27323 29 27381 75
rect 27427 29 27485 75
rect 27531 29 27589 75
rect 27635 29 27693 75
rect 27739 29 27797 75
rect 27843 29 27901 75
rect 27947 29 28005 75
rect 28051 29 28109 75
rect 28155 29 28213 75
rect 28259 29 28281 75
rect -28281 -29 28281 29
rect -28281 -75 -28259 -29
rect -28213 -75 -28155 -29
rect -28109 -75 -28051 -29
rect -28005 -75 -27947 -29
rect -27901 -75 -27843 -29
rect -27797 -75 -27739 -29
rect -27693 -75 -27635 -29
rect -27589 -75 -27531 -29
rect -27485 -75 -27427 -29
rect -27381 -75 -27323 -29
rect -27277 -75 -27219 -29
rect -27173 -75 -27115 -29
rect -27069 -75 -27011 -29
rect -26965 -75 -26907 -29
rect -26861 -75 -26803 -29
rect -26757 -75 -26699 -29
rect -26653 -75 -26595 -29
rect -26549 -75 -26491 -29
rect -26445 -75 -26387 -29
rect -26341 -75 -26283 -29
rect -26237 -75 -26179 -29
rect -26133 -75 -26075 -29
rect -26029 -75 -25971 -29
rect -25925 -75 -25867 -29
rect -25821 -75 -25763 -29
rect -25717 -75 -25659 -29
rect -25613 -75 -25555 -29
rect -25509 -75 -25451 -29
rect -25405 -75 -25347 -29
rect -25301 -75 -25243 -29
rect -25197 -75 -25139 -29
rect -25093 -75 -25035 -29
rect -24989 -75 -24931 -29
rect -24885 -75 -24827 -29
rect -24781 -75 -24723 -29
rect -24677 -75 -24619 -29
rect -24573 -75 -24515 -29
rect -24469 -75 -24411 -29
rect -24365 -75 -24307 -29
rect -24261 -75 -24203 -29
rect -24157 -75 -24099 -29
rect -24053 -75 -23995 -29
rect -23949 -75 -23891 -29
rect -23845 -75 -23787 -29
rect -23741 -75 -23683 -29
rect -23637 -75 -23579 -29
rect -23533 -75 -23475 -29
rect -23429 -75 -23371 -29
rect -23325 -75 -23267 -29
rect -23221 -75 -23163 -29
rect -23117 -75 -23059 -29
rect -23013 -75 -22955 -29
rect -22909 -75 -22851 -29
rect -22805 -75 -22747 -29
rect -22701 -75 -22643 -29
rect -22597 -75 -22539 -29
rect -22493 -75 -22435 -29
rect -22389 -75 -22331 -29
rect -22285 -75 -22227 -29
rect -22181 -75 -22123 -29
rect -22077 -75 -22019 -29
rect -21973 -75 -21915 -29
rect -21869 -75 -21811 -29
rect -21765 -75 -21707 -29
rect -21661 -75 -21603 -29
rect -21557 -75 -21499 -29
rect -21453 -75 -21395 -29
rect -21349 -75 -21291 -29
rect -21245 -75 -21187 -29
rect -21141 -75 -21083 -29
rect -21037 -75 -20979 -29
rect -20933 -75 -20875 -29
rect -20829 -75 -20771 -29
rect -20725 -75 -20667 -29
rect -20621 -75 -20563 -29
rect -20517 -75 -20459 -29
rect -20413 -75 -20355 -29
rect -20309 -75 -20251 -29
rect -20205 -75 -20147 -29
rect -20101 -75 -20043 -29
rect -19997 -75 -19939 -29
rect -19893 -75 -19835 -29
rect -19789 -75 -19731 -29
rect -19685 -75 -19627 -29
rect -19581 -75 -19523 -29
rect -19477 -75 -19419 -29
rect -19373 -75 -19315 -29
rect -19269 -75 -19211 -29
rect -19165 -75 -19107 -29
rect -19061 -75 -19003 -29
rect -18957 -75 -18899 -29
rect -18853 -75 -18795 -29
rect -18749 -75 -18691 -29
rect -18645 -75 -18587 -29
rect -18541 -75 -18483 -29
rect -18437 -75 -18379 -29
rect -18333 -75 -18275 -29
rect -18229 -75 -18171 -29
rect -18125 -75 -18067 -29
rect -18021 -75 -17963 -29
rect -17917 -75 -17859 -29
rect -17813 -75 -17755 -29
rect -17709 -75 -17651 -29
rect -17605 -75 -17547 -29
rect -17501 -75 -17443 -29
rect -17397 -75 -17339 -29
rect -17293 -75 -17235 -29
rect -17189 -75 -17131 -29
rect -17085 -75 -17027 -29
rect -16981 -75 -16923 -29
rect -16877 -75 -16819 -29
rect -16773 -75 -16715 -29
rect -16669 -75 -16611 -29
rect -16565 -75 -16507 -29
rect -16461 -75 -16403 -29
rect -16357 -75 -16299 -29
rect -16253 -75 -16195 -29
rect -16149 -75 -16091 -29
rect -16045 -75 -15987 -29
rect -15941 -75 -15883 -29
rect -15837 -75 -15779 -29
rect -15733 -75 -15675 -29
rect -15629 -75 -15571 -29
rect -15525 -75 -15467 -29
rect -15421 -75 -15363 -29
rect -15317 -75 -15259 -29
rect -15213 -75 -15155 -29
rect -15109 -75 -15051 -29
rect -15005 -75 -14947 -29
rect -14901 -75 -14843 -29
rect -14797 -75 -14739 -29
rect -14693 -75 -14635 -29
rect -14589 -75 -14531 -29
rect -14485 -75 -14427 -29
rect -14381 -75 -14323 -29
rect -14277 -75 -14219 -29
rect -14173 -75 -14115 -29
rect -14069 -75 -14011 -29
rect -13965 -75 -13907 -29
rect -13861 -75 -13803 -29
rect -13757 -75 -13699 -29
rect -13653 -75 -13595 -29
rect -13549 -75 -13491 -29
rect -13445 -75 -13387 -29
rect -13341 -75 -13283 -29
rect -13237 -75 -13179 -29
rect -13133 -75 -13075 -29
rect -13029 -75 -12971 -29
rect -12925 -75 -12867 -29
rect -12821 -75 -12763 -29
rect -12717 -75 -12659 -29
rect -12613 -75 -12555 -29
rect -12509 -75 -12451 -29
rect -12405 -75 -12347 -29
rect -12301 -75 -12243 -29
rect -12197 -75 -12139 -29
rect -12093 -75 -12035 -29
rect -11989 -75 -11931 -29
rect -11885 -75 -11827 -29
rect -11781 -75 -11723 -29
rect -11677 -75 -11619 -29
rect -11573 -75 -11515 -29
rect -11469 -75 -11411 -29
rect -11365 -75 -11307 -29
rect -11261 -75 -11203 -29
rect -11157 -75 -11099 -29
rect -11053 -75 -10995 -29
rect -10949 -75 -10891 -29
rect -10845 -75 -10787 -29
rect -10741 -75 -10683 -29
rect -10637 -75 -10579 -29
rect -10533 -75 -10475 -29
rect -10429 -75 -10371 -29
rect -10325 -75 -10267 -29
rect -10221 -75 -10163 -29
rect -10117 -75 -10059 -29
rect -10013 -75 -9955 -29
rect -9909 -75 -9851 -29
rect -9805 -75 -9747 -29
rect -9701 -75 -9643 -29
rect -9597 -75 -9539 -29
rect -9493 -75 -9435 -29
rect -9389 -75 -9331 -29
rect -9285 -75 -9227 -29
rect -9181 -75 -9123 -29
rect -9077 -75 -9019 -29
rect -8973 -75 -8915 -29
rect -8869 -75 -8811 -29
rect -8765 -75 -8707 -29
rect -8661 -75 -8603 -29
rect -8557 -75 -8499 -29
rect -8453 -75 -8395 -29
rect -8349 -75 -8291 -29
rect -8245 -75 -8187 -29
rect -8141 -75 -8083 -29
rect -8037 -75 -7979 -29
rect -7933 -75 -7875 -29
rect -7829 -75 -7771 -29
rect -7725 -75 -7667 -29
rect -7621 -75 -7563 -29
rect -7517 -75 -7459 -29
rect -7413 -75 -7355 -29
rect -7309 -75 -7251 -29
rect -7205 -75 -7147 -29
rect -7101 -75 -7043 -29
rect -6997 -75 -6939 -29
rect -6893 -75 -6835 -29
rect -6789 -75 -6731 -29
rect -6685 -75 -6627 -29
rect -6581 -75 -6523 -29
rect -6477 -75 -6419 -29
rect -6373 -75 -6315 -29
rect -6269 -75 -6211 -29
rect -6165 -75 -6107 -29
rect -6061 -75 -6003 -29
rect -5957 -75 -5899 -29
rect -5853 -75 -5795 -29
rect -5749 -75 -5691 -29
rect -5645 -75 -5587 -29
rect -5541 -75 -5483 -29
rect -5437 -75 -5379 -29
rect -5333 -75 -5275 -29
rect -5229 -75 -5171 -29
rect -5125 -75 -5067 -29
rect -5021 -75 -4963 -29
rect -4917 -75 -4859 -29
rect -4813 -75 -4755 -29
rect -4709 -75 -4651 -29
rect -4605 -75 -4547 -29
rect -4501 -75 -4443 -29
rect -4397 -75 -4339 -29
rect -4293 -75 -4235 -29
rect -4189 -75 -4131 -29
rect -4085 -75 -4027 -29
rect -3981 -75 -3923 -29
rect -3877 -75 -3819 -29
rect -3773 -75 -3715 -29
rect -3669 -75 -3611 -29
rect -3565 -75 -3507 -29
rect -3461 -75 -3403 -29
rect -3357 -75 -3299 -29
rect -3253 -75 -3195 -29
rect -3149 -75 -3091 -29
rect -3045 -75 -2987 -29
rect -2941 -75 -2883 -29
rect -2837 -75 -2779 -29
rect -2733 -75 -2675 -29
rect -2629 -75 -2571 -29
rect -2525 -75 -2467 -29
rect -2421 -75 -2363 -29
rect -2317 -75 -2259 -29
rect -2213 -75 -2155 -29
rect -2109 -75 -2051 -29
rect -2005 -75 -1947 -29
rect -1901 -75 -1843 -29
rect -1797 -75 -1739 -29
rect -1693 -75 -1635 -29
rect -1589 -75 -1531 -29
rect -1485 -75 -1427 -29
rect -1381 -75 -1323 -29
rect -1277 -75 -1219 -29
rect -1173 -75 -1115 -29
rect -1069 -75 -1011 -29
rect -965 -75 -907 -29
rect -861 -75 -803 -29
rect -757 -75 -699 -29
rect -653 -75 -595 -29
rect -549 -75 -491 -29
rect -445 -75 -387 -29
rect -341 -75 -283 -29
rect -237 -75 -179 -29
rect -133 -75 -75 -29
rect -29 -75 29 -29
rect 75 -75 133 -29
rect 179 -75 237 -29
rect 283 -75 341 -29
rect 387 -75 445 -29
rect 491 -75 549 -29
rect 595 -75 653 -29
rect 699 -75 757 -29
rect 803 -75 861 -29
rect 907 -75 965 -29
rect 1011 -75 1069 -29
rect 1115 -75 1173 -29
rect 1219 -75 1277 -29
rect 1323 -75 1381 -29
rect 1427 -75 1485 -29
rect 1531 -75 1589 -29
rect 1635 -75 1693 -29
rect 1739 -75 1797 -29
rect 1843 -75 1901 -29
rect 1947 -75 2005 -29
rect 2051 -75 2109 -29
rect 2155 -75 2213 -29
rect 2259 -75 2317 -29
rect 2363 -75 2421 -29
rect 2467 -75 2525 -29
rect 2571 -75 2629 -29
rect 2675 -75 2733 -29
rect 2779 -75 2837 -29
rect 2883 -75 2941 -29
rect 2987 -75 3045 -29
rect 3091 -75 3149 -29
rect 3195 -75 3253 -29
rect 3299 -75 3357 -29
rect 3403 -75 3461 -29
rect 3507 -75 3565 -29
rect 3611 -75 3669 -29
rect 3715 -75 3773 -29
rect 3819 -75 3877 -29
rect 3923 -75 3981 -29
rect 4027 -75 4085 -29
rect 4131 -75 4189 -29
rect 4235 -75 4293 -29
rect 4339 -75 4397 -29
rect 4443 -75 4501 -29
rect 4547 -75 4605 -29
rect 4651 -75 4709 -29
rect 4755 -75 4813 -29
rect 4859 -75 4917 -29
rect 4963 -75 5021 -29
rect 5067 -75 5125 -29
rect 5171 -75 5229 -29
rect 5275 -75 5333 -29
rect 5379 -75 5437 -29
rect 5483 -75 5541 -29
rect 5587 -75 5645 -29
rect 5691 -75 5749 -29
rect 5795 -75 5853 -29
rect 5899 -75 5957 -29
rect 6003 -75 6061 -29
rect 6107 -75 6165 -29
rect 6211 -75 6269 -29
rect 6315 -75 6373 -29
rect 6419 -75 6477 -29
rect 6523 -75 6581 -29
rect 6627 -75 6685 -29
rect 6731 -75 6789 -29
rect 6835 -75 6893 -29
rect 6939 -75 6997 -29
rect 7043 -75 7101 -29
rect 7147 -75 7205 -29
rect 7251 -75 7309 -29
rect 7355 -75 7413 -29
rect 7459 -75 7517 -29
rect 7563 -75 7621 -29
rect 7667 -75 7725 -29
rect 7771 -75 7829 -29
rect 7875 -75 7933 -29
rect 7979 -75 8037 -29
rect 8083 -75 8141 -29
rect 8187 -75 8245 -29
rect 8291 -75 8349 -29
rect 8395 -75 8453 -29
rect 8499 -75 8557 -29
rect 8603 -75 8661 -29
rect 8707 -75 8765 -29
rect 8811 -75 8869 -29
rect 8915 -75 8973 -29
rect 9019 -75 9077 -29
rect 9123 -75 9181 -29
rect 9227 -75 9285 -29
rect 9331 -75 9389 -29
rect 9435 -75 9493 -29
rect 9539 -75 9597 -29
rect 9643 -75 9701 -29
rect 9747 -75 9805 -29
rect 9851 -75 9909 -29
rect 9955 -75 10013 -29
rect 10059 -75 10117 -29
rect 10163 -75 10221 -29
rect 10267 -75 10325 -29
rect 10371 -75 10429 -29
rect 10475 -75 10533 -29
rect 10579 -75 10637 -29
rect 10683 -75 10741 -29
rect 10787 -75 10845 -29
rect 10891 -75 10949 -29
rect 10995 -75 11053 -29
rect 11099 -75 11157 -29
rect 11203 -75 11261 -29
rect 11307 -75 11365 -29
rect 11411 -75 11469 -29
rect 11515 -75 11573 -29
rect 11619 -75 11677 -29
rect 11723 -75 11781 -29
rect 11827 -75 11885 -29
rect 11931 -75 11989 -29
rect 12035 -75 12093 -29
rect 12139 -75 12197 -29
rect 12243 -75 12301 -29
rect 12347 -75 12405 -29
rect 12451 -75 12509 -29
rect 12555 -75 12613 -29
rect 12659 -75 12717 -29
rect 12763 -75 12821 -29
rect 12867 -75 12925 -29
rect 12971 -75 13029 -29
rect 13075 -75 13133 -29
rect 13179 -75 13237 -29
rect 13283 -75 13341 -29
rect 13387 -75 13445 -29
rect 13491 -75 13549 -29
rect 13595 -75 13653 -29
rect 13699 -75 13757 -29
rect 13803 -75 13861 -29
rect 13907 -75 13965 -29
rect 14011 -75 14069 -29
rect 14115 -75 14173 -29
rect 14219 -75 14277 -29
rect 14323 -75 14381 -29
rect 14427 -75 14485 -29
rect 14531 -75 14589 -29
rect 14635 -75 14693 -29
rect 14739 -75 14797 -29
rect 14843 -75 14901 -29
rect 14947 -75 15005 -29
rect 15051 -75 15109 -29
rect 15155 -75 15213 -29
rect 15259 -75 15317 -29
rect 15363 -75 15421 -29
rect 15467 -75 15525 -29
rect 15571 -75 15629 -29
rect 15675 -75 15733 -29
rect 15779 -75 15837 -29
rect 15883 -75 15941 -29
rect 15987 -75 16045 -29
rect 16091 -75 16149 -29
rect 16195 -75 16253 -29
rect 16299 -75 16357 -29
rect 16403 -75 16461 -29
rect 16507 -75 16565 -29
rect 16611 -75 16669 -29
rect 16715 -75 16773 -29
rect 16819 -75 16877 -29
rect 16923 -75 16981 -29
rect 17027 -75 17085 -29
rect 17131 -75 17189 -29
rect 17235 -75 17293 -29
rect 17339 -75 17397 -29
rect 17443 -75 17501 -29
rect 17547 -75 17605 -29
rect 17651 -75 17709 -29
rect 17755 -75 17813 -29
rect 17859 -75 17917 -29
rect 17963 -75 18021 -29
rect 18067 -75 18125 -29
rect 18171 -75 18229 -29
rect 18275 -75 18333 -29
rect 18379 -75 18437 -29
rect 18483 -75 18541 -29
rect 18587 -75 18645 -29
rect 18691 -75 18749 -29
rect 18795 -75 18853 -29
rect 18899 -75 18957 -29
rect 19003 -75 19061 -29
rect 19107 -75 19165 -29
rect 19211 -75 19269 -29
rect 19315 -75 19373 -29
rect 19419 -75 19477 -29
rect 19523 -75 19581 -29
rect 19627 -75 19685 -29
rect 19731 -75 19789 -29
rect 19835 -75 19893 -29
rect 19939 -75 19997 -29
rect 20043 -75 20101 -29
rect 20147 -75 20205 -29
rect 20251 -75 20309 -29
rect 20355 -75 20413 -29
rect 20459 -75 20517 -29
rect 20563 -75 20621 -29
rect 20667 -75 20725 -29
rect 20771 -75 20829 -29
rect 20875 -75 20933 -29
rect 20979 -75 21037 -29
rect 21083 -75 21141 -29
rect 21187 -75 21245 -29
rect 21291 -75 21349 -29
rect 21395 -75 21453 -29
rect 21499 -75 21557 -29
rect 21603 -75 21661 -29
rect 21707 -75 21765 -29
rect 21811 -75 21869 -29
rect 21915 -75 21973 -29
rect 22019 -75 22077 -29
rect 22123 -75 22181 -29
rect 22227 -75 22285 -29
rect 22331 -75 22389 -29
rect 22435 -75 22493 -29
rect 22539 -75 22597 -29
rect 22643 -75 22701 -29
rect 22747 -75 22805 -29
rect 22851 -75 22909 -29
rect 22955 -75 23013 -29
rect 23059 -75 23117 -29
rect 23163 -75 23221 -29
rect 23267 -75 23325 -29
rect 23371 -75 23429 -29
rect 23475 -75 23533 -29
rect 23579 -75 23637 -29
rect 23683 -75 23741 -29
rect 23787 -75 23845 -29
rect 23891 -75 23949 -29
rect 23995 -75 24053 -29
rect 24099 -75 24157 -29
rect 24203 -75 24261 -29
rect 24307 -75 24365 -29
rect 24411 -75 24469 -29
rect 24515 -75 24573 -29
rect 24619 -75 24677 -29
rect 24723 -75 24781 -29
rect 24827 -75 24885 -29
rect 24931 -75 24989 -29
rect 25035 -75 25093 -29
rect 25139 -75 25197 -29
rect 25243 -75 25301 -29
rect 25347 -75 25405 -29
rect 25451 -75 25509 -29
rect 25555 -75 25613 -29
rect 25659 -75 25717 -29
rect 25763 -75 25821 -29
rect 25867 -75 25925 -29
rect 25971 -75 26029 -29
rect 26075 -75 26133 -29
rect 26179 -75 26237 -29
rect 26283 -75 26341 -29
rect 26387 -75 26445 -29
rect 26491 -75 26549 -29
rect 26595 -75 26653 -29
rect 26699 -75 26757 -29
rect 26803 -75 26861 -29
rect 26907 -75 26965 -29
rect 27011 -75 27069 -29
rect 27115 -75 27173 -29
rect 27219 -75 27277 -29
rect 27323 -75 27381 -29
rect 27427 -75 27485 -29
rect 27531 -75 27589 -29
rect 27635 -75 27693 -29
rect 27739 -75 27797 -29
rect 27843 -75 27901 -29
rect 27947 -75 28005 -29
rect 28051 -75 28109 -29
rect 28155 -75 28213 -29
rect 28259 -75 28281 -29
rect -28281 -97 28281 -75
<< psubdiffcont >>
rect -28259 29 -28213 75
rect -28155 29 -28109 75
rect -28051 29 -28005 75
rect -27947 29 -27901 75
rect -27843 29 -27797 75
rect -27739 29 -27693 75
rect -27635 29 -27589 75
rect -27531 29 -27485 75
rect -27427 29 -27381 75
rect -27323 29 -27277 75
rect -27219 29 -27173 75
rect -27115 29 -27069 75
rect -27011 29 -26965 75
rect -26907 29 -26861 75
rect -26803 29 -26757 75
rect -26699 29 -26653 75
rect -26595 29 -26549 75
rect -26491 29 -26445 75
rect -26387 29 -26341 75
rect -26283 29 -26237 75
rect -26179 29 -26133 75
rect -26075 29 -26029 75
rect -25971 29 -25925 75
rect -25867 29 -25821 75
rect -25763 29 -25717 75
rect -25659 29 -25613 75
rect -25555 29 -25509 75
rect -25451 29 -25405 75
rect -25347 29 -25301 75
rect -25243 29 -25197 75
rect -25139 29 -25093 75
rect -25035 29 -24989 75
rect -24931 29 -24885 75
rect -24827 29 -24781 75
rect -24723 29 -24677 75
rect -24619 29 -24573 75
rect -24515 29 -24469 75
rect -24411 29 -24365 75
rect -24307 29 -24261 75
rect -24203 29 -24157 75
rect -24099 29 -24053 75
rect -23995 29 -23949 75
rect -23891 29 -23845 75
rect -23787 29 -23741 75
rect -23683 29 -23637 75
rect -23579 29 -23533 75
rect -23475 29 -23429 75
rect -23371 29 -23325 75
rect -23267 29 -23221 75
rect -23163 29 -23117 75
rect -23059 29 -23013 75
rect -22955 29 -22909 75
rect -22851 29 -22805 75
rect -22747 29 -22701 75
rect -22643 29 -22597 75
rect -22539 29 -22493 75
rect -22435 29 -22389 75
rect -22331 29 -22285 75
rect -22227 29 -22181 75
rect -22123 29 -22077 75
rect -22019 29 -21973 75
rect -21915 29 -21869 75
rect -21811 29 -21765 75
rect -21707 29 -21661 75
rect -21603 29 -21557 75
rect -21499 29 -21453 75
rect -21395 29 -21349 75
rect -21291 29 -21245 75
rect -21187 29 -21141 75
rect -21083 29 -21037 75
rect -20979 29 -20933 75
rect -20875 29 -20829 75
rect -20771 29 -20725 75
rect -20667 29 -20621 75
rect -20563 29 -20517 75
rect -20459 29 -20413 75
rect -20355 29 -20309 75
rect -20251 29 -20205 75
rect -20147 29 -20101 75
rect -20043 29 -19997 75
rect -19939 29 -19893 75
rect -19835 29 -19789 75
rect -19731 29 -19685 75
rect -19627 29 -19581 75
rect -19523 29 -19477 75
rect -19419 29 -19373 75
rect -19315 29 -19269 75
rect -19211 29 -19165 75
rect -19107 29 -19061 75
rect -19003 29 -18957 75
rect -18899 29 -18853 75
rect -18795 29 -18749 75
rect -18691 29 -18645 75
rect -18587 29 -18541 75
rect -18483 29 -18437 75
rect -18379 29 -18333 75
rect -18275 29 -18229 75
rect -18171 29 -18125 75
rect -18067 29 -18021 75
rect -17963 29 -17917 75
rect -17859 29 -17813 75
rect -17755 29 -17709 75
rect -17651 29 -17605 75
rect -17547 29 -17501 75
rect -17443 29 -17397 75
rect -17339 29 -17293 75
rect -17235 29 -17189 75
rect -17131 29 -17085 75
rect -17027 29 -16981 75
rect -16923 29 -16877 75
rect -16819 29 -16773 75
rect -16715 29 -16669 75
rect -16611 29 -16565 75
rect -16507 29 -16461 75
rect -16403 29 -16357 75
rect -16299 29 -16253 75
rect -16195 29 -16149 75
rect -16091 29 -16045 75
rect -15987 29 -15941 75
rect -15883 29 -15837 75
rect -15779 29 -15733 75
rect -15675 29 -15629 75
rect -15571 29 -15525 75
rect -15467 29 -15421 75
rect -15363 29 -15317 75
rect -15259 29 -15213 75
rect -15155 29 -15109 75
rect -15051 29 -15005 75
rect -14947 29 -14901 75
rect -14843 29 -14797 75
rect -14739 29 -14693 75
rect -14635 29 -14589 75
rect -14531 29 -14485 75
rect -14427 29 -14381 75
rect -14323 29 -14277 75
rect -14219 29 -14173 75
rect -14115 29 -14069 75
rect -14011 29 -13965 75
rect -13907 29 -13861 75
rect -13803 29 -13757 75
rect -13699 29 -13653 75
rect -13595 29 -13549 75
rect -13491 29 -13445 75
rect -13387 29 -13341 75
rect -13283 29 -13237 75
rect -13179 29 -13133 75
rect -13075 29 -13029 75
rect -12971 29 -12925 75
rect -12867 29 -12821 75
rect -12763 29 -12717 75
rect -12659 29 -12613 75
rect -12555 29 -12509 75
rect -12451 29 -12405 75
rect -12347 29 -12301 75
rect -12243 29 -12197 75
rect -12139 29 -12093 75
rect -12035 29 -11989 75
rect -11931 29 -11885 75
rect -11827 29 -11781 75
rect -11723 29 -11677 75
rect -11619 29 -11573 75
rect -11515 29 -11469 75
rect -11411 29 -11365 75
rect -11307 29 -11261 75
rect -11203 29 -11157 75
rect -11099 29 -11053 75
rect -10995 29 -10949 75
rect -10891 29 -10845 75
rect -10787 29 -10741 75
rect -10683 29 -10637 75
rect -10579 29 -10533 75
rect -10475 29 -10429 75
rect -10371 29 -10325 75
rect -10267 29 -10221 75
rect -10163 29 -10117 75
rect -10059 29 -10013 75
rect -9955 29 -9909 75
rect -9851 29 -9805 75
rect -9747 29 -9701 75
rect -9643 29 -9597 75
rect -9539 29 -9493 75
rect -9435 29 -9389 75
rect -9331 29 -9285 75
rect -9227 29 -9181 75
rect -9123 29 -9077 75
rect -9019 29 -8973 75
rect -8915 29 -8869 75
rect -8811 29 -8765 75
rect -8707 29 -8661 75
rect -8603 29 -8557 75
rect -8499 29 -8453 75
rect -8395 29 -8349 75
rect -8291 29 -8245 75
rect -8187 29 -8141 75
rect -8083 29 -8037 75
rect -7979 29 -7933 75
rect -7875 29 -7829 75
rect -7771 29 -7725 75
rect -7667 29 -7621 75
rect -7563 29 -7517 75
rect -7459 29 -7413 75
rect -7355 29 -7309 75
rect -7251 29 -7205 75
rect -7147 29 -7101 75
rect -7043 29 -6997 75
rect -6939 29 -6893 75
rect -6835 29 -6789 75
rect -6731 29 -6685 75
rect -6627 29 -6581 75
rect -6523 29 -6477 75
rect -6419 29 -6373 75
rect -6315 29 -6269 75
rect -6211 29 -6165 75
rect -6107 29 -6061 75
rect -6003 29 -5957 75
rect -5899 29 -5853 75
rect -5795 29 -5749 75
rect -5691 29 -5645 75
rect -5587 29 -5541 75
rect -5483 29 -5437 75
rect -5379 29 -5333 75
rect -5275 29 -5229 75
rect -5171 29 -5125 75
rect -5067 29 -5021 75
rect -4963 29 -4917 75
rect -4859 29 -4813 75
rect -4755 29 -4709 75
rect -4651 29 -4605 75
rect -4547 29 -4501 75
rect -4443 29 -4397 75
rect -4339 29 -4293 75
rect -4235 29 -4189 75
rect -4131 29 -4085 75
rect -4027 29 -3981 75
rect -3923 29 -3877 75
rect -3819 29 -3773 75
rect -3715 29 -3669 75
rect -3611 29 -3565 75
rect -3507 29 -3461 75
rect -3403 29 -3357 75
rect -3299 29 -3253 75
rect -3195 29 -3149 75
rect -3091 29 -3045 75
rect -2987 29 -2941 75
rect -2883 29 -2837 75
rect -2779 29 -2733 75
rect -2675 29 -2629 75
rect -2571 29 -2525 75
rect -2467 29 -2421 75
rect -2363 29 -2317 75
rect -2259 29 -2213 75
rect -2155 29 -2109 75
rect -2051 29 -2005 75
rect -1947 29 -1901 75
rect -1843 29 -1797 75
rect -1739 29 -1693 75
rect -1635 29 -1589 75
rect -1531 29 -1485 75
rect -1427 29 -1381 75
rect -1323 29 -1277 75
rect -1219 29 -1173 75
rect -1115 29 -1069 75
rect -1011 29 -965 75
rect -907 29 -861 75
rect -803 29 -757 75
rect -699 29 -653 75
rect -595 29 -549 75
rect -491 29 -445 75
rect -387 29 -341 75
rect -283 29 -237 75
rect -179 29 -133 75
rect -75 29 -29 75
rect 29 29 75 75
rect 133 29 179 75
rect 237 29 283 75
rect 341 29 387 75
rect 445 29 491 75
rect 549 29 595 75
rect 653 29 699 75
rect 757 29 803 75
rect 861 29 907 75
rect 965 29 1011 75
rect 1069 29 1115 75
rect 1173 29 1219 75
rect 1277 29 1323 75
rect 1381 29 1427 75
rect 1485 29 1531 75
rect 1589 29 1635 75
rect 1693 29 1739 75
rect 1797 29 1843 75
rect 1901 29 1947 75
rect 2005 29 2051 75
rect 2109 29 2155 75
rect 2213 29 2259 75
rect 2317 29 2363 75
rect 2421 29 2467 75
rect 2525 29 2571 75
rect 2629 29 2675 75
rect 2733 29 2779 75
rect 2837 29 2883 75
rect 2941 29 2987 75
rect 3045 29 3091 75
rect 3149 29 3195 75
rect 3253 29 3299 75
rect 3357 29 3403 75
rect 3461 29 3507 75
rect 3565 29 3611 75
rect 3669 29 3715 75
rect 3773 29 3819 75
rect 3877 29 3923 75
rect 3981 29 4027 75
rect 4085 29 4131 75
rect 4189 29 4235 75
rect 4293 29 4339 75
rect 4397 29 4443 75
rect 4501 29 4547 75
rect 4605 29 4651 75
rect 4709 29 4755 75
rect 4813 29 4859 75
rect 4917 29 4963 75
rect 5021 29 5067 75
rect 5125 29 5171 75
rect 5229 29 5275 75
rect 5333 29 5379 75
rect 5437 29 5483 75
rect 5541 29 5587 75
rect 5645 29 5691 75
rect 5749 29 5795 75
rect 5853 29 5899 75
rect 5957 29 6003 75
rect 6061 29 6107 75
rect 6165 29 6211 75
rect 6269 29 6315 75
rect 6373 29 6419 75
rect 6477 29 6523 75
rect 6581 29 6627 75
rect 6685 29 6731 75
rect 6789 29 6835 75
rect 6893 29 6939 75
rect 6997 29 7043 75
rect 7101 29 7147 75
rect 7205 29 7251 75
rect 7309 29 7355 75
rect 7413 29 7459 75
rect 7517 29 7563 75
rect 7621 29 7667 75
rect 7725 29 7771 75
rect 7829 29 7875 75
rect 7933 29 7979 75
rect 8037 29 8083 75
rect 8141 29 8187 75
rect 8245 29 8291 75
rect 8349 29 8395 75
rect 8453 29 8499 75
rect 8557 29 8603 75
rect 8661 29 8707 75
rect 8765 29 8811 75
rect 8869 29 8915 75
rect 8973 29 9019 75
rect 9077 29 9123 75
rect 9181 29 9227 75
rect 9285 29 9331 75
rect 9389 29 9435 75
rect 9493 29 9539 75
rect 9597 29 9643 75
rect 9701 29 9747 75
rect 9805 29 9851 75
rect 9909 29 9955 75
rect 10013 29 10059 75
rect 10117 29 10163 75
rect 10221 29 10267 75
rect 10325 29 10371 75
rect 10429 29 10475 75
rect 10533 29 10579 75
rect 10637 29 10683 75
rect 10741 29 10787 75
rect 10845 29 10891 75
rect 10949 29 10995 75
rect 11053 29 11099 75
rect 11157 29 11203 75
rect 11261 29 11307 75
rect 11365 29 11411 75
rect 11469 29 11515 75
rect 11573 29 11619 75
rect 11677 29 11723 75
rect 11781 29 11827 75
rect 11885 29 11931 75
rect 11989 29 12035 75
rect 12093 29 12139 75
rect 12197 29 12243 75
rect 12301 29 12347 75
rect 12405 29 12451 75
rect 12509 29 12555 75
rect 12613 29 12659 75
rect 12717 29 12763 75
rect 12821 29 12867 75
rect 12925 29 12971 75
rect 13029 29 13075 75
rect 13133 29 13179 75
rect 13237 29 13283 75
rect 13341 29 13387 75
rect 13445 29 13491 75
rect 13549 29 13595 75
rect 13653 29 13699 75
rect 13757 29 13803 75
rect 13861 29 13907 75
rect 13965 29 14011 75
rect 14069 29 14115 75
rect 14173 29 14219 75
rect 14277 29 14323 75
rect 14381 29 14427 75
rect 14485 29 14531 75
rect 14589 29 14635 75
rect 14693 29 14739 75
rect 14797 29 14843 75
rect 14901 29 14947 75
rect 15005 29 15051 75
rect 15109 29 15155 75
rect 15213 29 15259 75
rect 15317 29 15363 75
rect 15421 29 15467 75
rect 15525 29 15571 75
rect 15629 29 15675 75
rect 15733 29 15779 75
rect 15837 29 15883 75
rect 15941 29 15987 75
rect 16045 29 16091 75
rect 16149 29 16195 75
rect 16253 29 16299 75
rect 16357 29 16403 75
rect 16461 29 16507 75
rect 16565 29 16611 75
rect 16669 29 16715 75
rect 16773 29 16819 75
rect 16877 29 16923 75
rect 16981 29 17027 75
rect 17085 29 17131 75
rect 17189 29 17235 75
rect 17293 29 17339 75
rect 17397 29 17443 75
rect 17501 29 17547 75
rect 17605 29 17651 75
rect 17709 29 17755 75
rect 17813 29 17859 75
rect 17917 29 17963 75
rect 18021 29 18067 75
rect 18125 29 18171 75
rect 18229 29 18275 75
rect 18333 29 18379 75
rect 18437 29 18483 75
rect 18541 29 18587 75
rect 18645 29 18691 75
rect 18749 29 18795 75
rect 18853 29 18899 75
rect 18957 29 19003 75
rect 19061 29 19107 75
rect 19165 29 19211 75
rect 19269 29 19315 75
rect 19373 29 19419 75
rect 19477 29 19523 75
rect 19581 29 19627 75
rect 19685 29 19731 75
rect 19789 29 19835 75
rect 19893 29 19939 75
rect 19997 29 20043 75
rect 20101 29 20147 75
rect 20205 29 20251 75
rect 20309 29 20355 75
rect 20413 29 20459 75
rect 20517 29 20563 75
rect 20621 29 20667 75
rect 20725 29 20771 75
rect 20829 29 20875 75
rect 20933 29 20979 75
rect 21037 29 21083 75
rect 21141 29 21187 75
rect 21245 29 21291 75
rect 21349 29 21395 75
rect 21453 29 21499 75
rect 21557 29 21603 75
rect 21661 29 21707 75
rect 21765 29 21811 75
rect 21869 29 21915 75
rect 21973 29 22019 75
rect 22077 29 22123 75
rect 22181 29 22227 75
rect 22285 29 22331 75
rect 22389 29 22435 75
rect 22493 29 22539 75
rect 22597 29 22643 75
rect 22701 29 22747 75
rect 22805 29 22851 75
rect 22909 29 22955 75
rect 23013 29 23059 75
rect 23117 29 23163 75
rect 23221 29 23267 75
rect 23325 29 23371 75
rect 23429 29 23475 75
rect 23533 29 23579 75
rect 23637 29 23683 75
rect 23741 29 23787 75
rect 23845 29 23891 75
rect 23949 29 23995 75
rect 24053 29 24099 75
rect 24157 29 24203 75
rect 24261 29 24307 75
rect 24365 29 24411 75
rect 24469 29 24515 75
rect 24573 29 24619 75
rect 24677 29 24723 75
rect 24781 29 24827 75
rect 24885 29 24931 75
rect 24989 29 25035 75
rect 25093 29 25139 75
rect 25197 29 25243 75
rect 25301 29 25347 75
rect 25405 29 25451 75
rect 25509 29 25555 75
rect 25613 29 25659 75
rect 25717 29 25763 75
rect 25821 29 25867 75
rect 25925 29 25971 75
rect 26029 29 26075 75
rect 26133 29 26179 75
rect 26237 29 26283 75
rect 26341 29 26387 75
rect 26445 29 26491 75
rect 26549 29 26595 75
rect 26653 29 26699 75
rect 26757 29 26803 75
rect 26861 29 26907 75
rect 26965 29 27011 75
rect 27069 29 27115 75
rect 27173 29 27219 75
rect 27277 29 27323 75
rect 27381 29 27427 75
rect 27485 29 27531 75
rect 27589 29 27635 75
rect 27693 29 27739 75
rect 27797 29 27843 75
rect 27901 29 27947 75
rect 28005 29 28051 75
rect 28109 29 28155 75
rect 28213 29 28259 75
rect -28259 -75 -28213 -29
rect -28155 -75 -28109 -29
rect -28051 -75 -28005 -29
rect -27947 -75 -27901 -29
rect -27843 -75 -27797 -29
rect -27739 -75 -27693 -29
rect -27635 -75 -27589 -29
rect -27531 -75 -27485 -29
rect -27427 -75 -27381 -29
rect -27323 -75 -27277 -29
rect -27219 -75 -27173 -29
rect -27115 -75 -27069 -29
rect -27011 -75 -26965 -29
rect -26907 -75 -26861 -29
rect -26803 -75 -26757 -29
rect -26699 -75 -26653 -29
rect -26595 -75 -26549 -29
rect -26491 -75 -26445 -29
rect -26387 -75 -26341 -29
rect -26283 -75 -26237 -29
rect -26179 -75 -26133 -29
rect -26075 -75 -26029 -29
rect -25971 -75 -25925 -29
rect -25867 -75 -25821 -29
rect -25763 -75 -25717 -29
rect -25659 -75 -25613 -29
rect -25555 -75 -25509 -29
rect -25451 -75 -25405 -29
rect -25347 -75 -25301 -29
rect -25243 -75 -25197 -29
rect -25139 -75 -25093 -29
rect -25035 -75 -24989 -29
rect -24931 -75 -24885 -29
rect -24827 -75 -24781 -29
rect -24723 -75 -24677 -29
rect -24619 -75 -24573 -29
rect -24515 -75 -24469 -29
rect -24411 -75 -24365 -29
rect -24307 -75 -24261 -29
rect -24203 -75 -24157 -29
rect -24099 -75 -24053 -29
rect -23995 -75 -23949 -29
rect -23891 -75 -23845 -29
rect -23787 -75 -23741 -29
rect -23683 -75 -23637 -29
rect -23579 -75 -23533 -29
rect -23475 -75 -23429 -29
rect -23371 -75 -23325 -29
rect -23267 -75 -23221 -29
rect -23163 -75 -23117 -29
rect -23059 -75 -23013 -29
rect -22955 -75 -22909 -29
rect -22851 -75 -22805 -29
rect -22747 -75 -22701 -29
rect -22643 -75 -22597 -29
rect -22539 -75 -22493 -29
rect -22435 -75 -22389 -29
rect -22331 -75 -22285 -29
rect -22227 -75 -22181 -29
rect -22123 -75 -22077 -29
rect -22019 -75 -21973 -29
rect -21915 -75 -21869 -29
rect -21811 -75 -21765 -29
rect -21707 -75 -21661 -29
rect -21603 -75 -21557 -29
rect -21499 -75 -21453 -29
rect -21395 -75 -21349 -29
rect -21291 -75 -21245 -29
rect -21187 -75 -21141 -29
rect -21083 -75 -21037 -29
rect -20979 -75 -20933 -29
rect -20875 -75 -20829 -29
rect -20771 -75 -20725 -29
rect -20667 -75 -20621 -29
rect -20563 -75 -20517 -29
rect -20459 -75 -20413 -29
rect -20355 -75 -20309 -29
rect -20251 -75 -20205 -29
rect -20147 -75 -20101 -29
rect -20043 -75 -19997 -29
rect -19939 -75 -19893 -29
rect -19835 -75 -19789 -29
rect -19731 -75 -19685 -29
rect -19627 -75 -19581 -29
rect -19523 -75 -19477 -29
rect -19419 -75 -19373 -29
rect -19315 -75 -19269 -29
rect -19211 -75 -19165 -29
rect -19107 -75 -19061 -29
rect -19003 -75 -18957 -29
rect -18899 -75 -18853 -29
rect -18795 -75 -18749 -29
rect -18691 -75 -18645 -29
rect -18587 -75 -18541 -29
rect -18483 -75 -18437 -29
rect -18379 -75 -18333 -29
rect -18275 -75 -18229 -29
rect -18171 -75 -18125 -29
rect -18067 -75 -18021 -29
rect -17963 -75 -17917 -29
rect -17859 -75 -17813 -29
rect -17755 -75 -17709 -29
rect -17651 -75 -17605 -29
rect -17547 -75 -17501 -29
rect -17443 -75 -17397 -29
rect -17339 -75 -17293 -29
rect -17235 -75 -17189 -29
rect -17131 -75 -17085 -29
rect -17027 -75 -16981 -29
rect -16923 -75 -16877 -29
rect -16819 -75 -16773 -29
rect -16715 -75 -16669 -29
rect -16611 -75 -16565 -29
rect -16507 -75 -16461 -29
rect -16403 -75 -16357 -29
rect -16299 -75 -16253 -29
rect -16195 -75 -16149 -29
rect -16091 -75 -16045 -29
rect -15987 -75 -15941 -29
rect -15883 -75 -15837 -29
rect -15779 -75 -15733 -29
rect -15675 -75 -15629 -29
rect -15571 -75 -15525 -29
rect -15467 -75 -15421 -29
rect -15363 -75 -15317 -29
rect -15259 -75 -15213 -29
rect -15155 -75 -15109 -29
rect -15051 -75 -15005 -29
rect -14947 -75 -14901 -29
rect -14843 -75 -14797 -29
rect -14739 -75 -14693 -29
rect -14635 -75 -14589 -29
rect -14531 -75 -14485 -29
rect -14427 -75 -14381 -29
rect -14323 -75 -14277 -29
rect -14219 -75 -14173 -29
rect -14115 -75 -14069 -29
rect -14011 -75 -13965 -29
rect -13907 -75 -13861 -29
rect -13803 -75 -13757 -29
rect -13699 -75 -13653 -29
rect -13595 -75 -13549 -29
rect -13491 -75 -13445 -29
rect -13387 -75 -13341 -29
rect -13283 -75 -13237 -29
rect -13179 -75 -13133 -29
rect -13075 -75 -13029 -29
rect -12971 -75 -12925 -29
rect -12867 -75 -12821 -29
rect -12763 -75 -12717 -29
rect -12659 -75 -12613 -29
rect -12555 -75 -12509 -29
rect -12451 -75 -12405 -29
rect -12347 -75 -12301 -29
rect -12243 -75 -12197 -29
rect -12139 -75 -12093 -29
rect -12035 -75 -11989 -29
rect -11931 -75 -11885 -29
rect -11827 -75 -11781 -29
rect -11723 -75 -11677 -29
rect -11619 -75 -11573 -29
rect -11515 -75 -11469 -29
rect -11411 -75 -11365 -29
rect -11307 -75 -11261 -29
rect -11203 -75 -11157 -29
rect -11099 -75 -11053 -29
rect -10995 -75 -10949 -29
rect -10891 -75 -10845 -29
rect -10787 -75 -10741 -29
rect -10683 -75 -10637 -29
rect -10579 -75 -10533 -29
rect -10475 -75 -10429 -29
rect -10371 -75 -10325 -29
rect -10267 -75 -10221 -29
rect -10163 -75 -10117 -29
rect -10059 -75 -10013 -29
rect -9955 -75 -9909 -29
rect -9851 -75 -9805 -29
rect -9747 -75 -9701 -29
rect -9643 -75 -9597 -29
rect -9539 -75 -9493 -29
rect -9435 -75 -9389 -29
rect -9331 -75 -9285 -29
rect -9227 -75 -9181 -29
rect -9123 -75 -9077 -29
rect -9019 -75 -8973 -29
rect -8915 -75 -8869 -29
rect -8811 -75 -8765 -29
rect -8707 -75 -8661 -29
rect -8603 -75 -8557 -29
rect -8499 -75 -8453 -29
rect -8395 -75 -8349 -29
rect -8291 -75 -8245 -29
rect -8187 -75 -8141 -29
rect -8083 -75 -8037 -29
rect -7979 -75 -7933 -29
rect -7875 -75 -7829 -29
rect -7771 -75 -7725 -29
rect -7667 -75 -7621 -29
rect -7563 -75 -7517 -29
rect -7459 -75 -7413 -29
rect -7355 -75 -7309 -29
rect -7251 -75 -7205 -29
rect -7147 -75 -7101 -29
rect -7043 -75 -6997 -29
rect -6939 -75 -6893 -29
rect -6835 -75 -6789 -29
rect -6731 -75 -6685 -29
rect -6627 -75 -6581 -29
rect -6523 -75 -6477 -29
rect -6419 -75 -6373 -29
rect -6315 -75 -6269 -29
rect -6211 -75 -6165 -29
rect -6107 -75 -6061 -29
rect -6003 -75 -5957 -29
rect -5899 -75 -5853 -29
rect -5795 -75 -5749 -29
rect -5691 -75 -5645 -29
rect -5587 -75 -5541 -29
rect -5483 -75 -5437 -29
rect -5379 -75 -5333 -29
rect -5275 -75 -5229 -29
rect -5171 -75 -5125 -29
rect -5067 -75 -5021 -29
rect -4963 -75 -4917 -29
rect -4859 -75 -4813 -29
rect -4755 -75 -4709 -29
rect -4651 -75 -4605 -29
rect -4547 -75 -4501 -29
rect -4443 -75 -4397 -29
rect -4339 -75 -4293 -29
rect -4235 -75 -4189 -29
rect -4131 -75 -4085 -29
rect -4027 -75 -3981 -29
rect -3923 -75 -3877 -29
rect -3819 -75 -3773 -29
rect -3715 -75 -3669 -29
rect -3611 -75 -3565 -29
rect -3507 -75 -3461 -29
rect -3403 -75 -3357 -29
rect -3299 -75 -3253 -29
rect -3195 -75 -3149 -29
rect -3091 -75 -3045 -29
rect -2987 -75 -2941 -29
rect -2883 -75 -2837 -29
rect -2779 -75 -2733 -29
rect -2675 -75 -2629 -29
rect -2571 -75 -2525 -29
rect -2467 -75 -2421 -29
rect -2363 -75 -2317 -29
rect -2259 -75 -2213 -29
rect -2155 -75 -2109 -29
rect -2051 -75 -2005 -29
rect -1947 -75 -1901 -29
rect -1843 -75 -1797 -29
rect -1739 -75 -1693 -29
rect -1635 -75 -1589 -29
rect -1531 -75 -1485 -29
rect -1427 -75 -1381 -29
rect -1323 -75 -1277 -29
rect -1219 -75 -1173 -29
rect -1115 -75 -1069 -29
rect -1011 -75 -965 -29
rect -907 -75 -861 -29
rect -803 -75 -757 -29
rect -699 -75 -653 -29
rect -595 -75 -549 -29
rect -491 -75 -445 -29
rect -387 -75 -341 -29
rect -283 -75 -237 -29
rect -179 -75 -133 -29
rect -75 -75 -29 -29
rect 29 -75 75 -29
rect 133 -75 179 -29
rect 237 -75 283 -29
rect 341 -75 387 -29
rect 445 -75 491 -29
rect 549 -75 595 -29
rect 653 -75 699 -29
rect 757 -75 803 -29
rect 861 -75 907 -29
rect 965 -75 1011 -29
rect 1069 -75 1115 -29
rect 1173 -75 1219 -29
rect 1277 -75 1323 -29
rect 1381 -75 1427 -29
rect 1485 -75 1531 -29
rect 1589 -75 1635 -29
rect 1693 -75 1739 -29
rect 1797 -75 1843 -29
rect 1901 -75 1947 -29
rect 2005 -75 2051 -29
rect 2109 -75 2155 -29
rect 2213 -75 2259 -29
rect 2317 -75 2363 -29
rect 2421 -75 2467 -29
rect 2525 -75 2571 -29
rect 2629 -75 2675 -29
rect 2733 -75 2779 -29
rect 2837 -75 2883 -29
rect 2941 -75 2987 -29
rect 3045 -75 3091 -29
rect 3149 -75 3195 -29
rect 3253 -75 3299 -29
rect 3357 -75 3403 -29
rect 3461 -75 3507 -29
rect 3565 -75 3611 -29
rect 3669 -75 3715 -29
rect 3773 -75 3819 -29
rect 3877 -75 3923 -29
rect 3981 -75 4027 -29
rect 4085 -75 4131 -29
rect 4189 -75 4235 -29
rect 4293 -75 4339 -29
rect 4397 -75 4443 -29
rect 4501 -75 4547 -29
rect 4605 -75 4651 -29
rect 4709 -75 4755 -29
rect 4813 -75 4859 -29
rect 4917 -75 4963 -29
rect 5021 -75 5067 -29
rect 5125 -75 5171 -29
rect 5229 -75 5275 -29
rect 5333 -75 5379 -29
rect 5437 -75 5483 -29
rect 5541 -75 5587 -29
rect 5645 -75 5691 -29
rect 5749 -75 5795 -29
rect 5853 -75 5899 -29
rect 5957 -75 6003 -29
rect 6061 -75 6107 -29
rect 6165 -75 6211 -29
rect 6269 -75 6315 -29
rect 6373 -75 6419 -29
rect 6477 -75 6523 -29
rect 6581 -75 6627 -29
rect 6685 -75 6731 -29
rect 6789 -75 6835 -29
rect 6893 -75 6939 -29
rect 6997 -75 7043 -29
rect 7101 -75 7147 -29
rect 7205 -75 7251 -29
rect 7309 -75 7355 -29
rect 7413 -75 7459 -29
rect 7517 -75 7563 -29
rect 7621 -75 7667 -29
rect 7725 -75 7771 -29
rect 7829 -75 7875 -29
rect 7933 -75 7979 -29
rect 8037 -75 8083 -29
rect 8141 -75 8187 -29
rect 8245 -75 8291 -29
rect 8349 -75 8395 -29
rect 8453 -75 8499 -29
rect 8557 -75 8603 -29
rect 8661 -75 8707 -29
rect 8765 -75 8811 -29
rect 8869 -75 8915 -29
rect 8973 -75 9019 -29
rect 9077 -75 9123 -29
rect 9181 -75 9227 -29
rect 9285 -75 9331 -29
rect 9389 -75 9435 -29
rect 9493 -75 9539 -29
rect 9597 -75 9643 -29
rect 9701 -75 9747 -29
rect 9805 -75 9851 -29
rect 9909 -75 9955 -29
rect 10013 -75 10059 -29
rect 10117 -75 10163 -29
rect 10221 -75 10267 -29
rect 10325 -75 10371 -29
rect 10429 -75 10475 -29
rect 10533 -75 10579 -29
rect 10637 -75 10683 -29
rect 10741 -75 10787 -29
rect 10845 -75 10891 -29
rect 10949 -75 10995 -29
rect 11053 -75 11099 -29
rect 11157 -75 11203 -29
rect 11261 -75 11307 -29
rect 11365 -75 11411 -29
rect 11469 -75 11515 -29
rect 11573 -75 11619 -29
rect 11677 -75 11723 -29
rect 11781 -75 11827 -29
rect 11885 -75 11931 -29
rect 11989 -75 12035 -29
rect 12093 -75 12139 -29
rect 12197 -75 12243 -29
rect 12301 -75 12347 -29
rect 12405 -75 12451 -29
rect 12509 -75 12555 -29
rect 12613 -75 12659 -29
rect 12717 -75 12763 -29
rect 12821 -75 12867 -29
rect 12925 -75 12971 -29
rect 13029 -75 13075 -29
rect 13133 -75 13179 -29
rect 13237 -75 13283 -29
rect 13341 -75 13387 -29
rect 13445 -75 13491 -29
rect 13549 -75 13595 -29
rect 13653 -75 13699 -29
rect 13757 -75 13803 -29
rect 13861 -75 13907 -29
rect 13965 -75 14011 -29
rect 14069 -75 14115 -29
rect 14173 -75 14219 -29
rect 14277 -75 14323 -29
rect 14381 -75 14427 -29
rect 14485 -75 14531 -29
rect 14589 -75 14635 -29
rect 14693 -75 14739 -29
rect 14797 -75 14843 -29
rect 14901 -75 14947 -29
rect 15005 -75 15051 -29
rect 15109 -75 15155 -29
rect 15213 -75 15259 -29
rect 15317 -75 15363 -29
rect 15421 -75 15467 -29
rect 15525 -75 15571 -29
rect 15629 -75 15675 -29
rect 15733 -75 15779 -29
rect 15837 -75 15883 -29
rect 15941 -75 15987 -29
rect 16045 -75 16091 -29
rect 16149 -75 16195 -29
rect 16253 -75 16299 -29
rect 16357 -75 16403 -29
rect 16461 -75 16507 -29
rect 16565 -75 16611 -29
rect 16669 -75 16715 -29
rect 16773 -75 16819 -29
rect 16877 -75 16923 -29
rect 16981 -75 17027 -29
rect 17085 -75 17131 -29
rect 17189 -75 17235 -29
rect 17293 -75 17339 -29
rect 17397 -75 17443 -29
rect 17501 -75 17547 -29
rect 17605 -75 17651 -29
rect 17709 -75 17755 -29
rect 17813 -75 17859 -29
rect 17917 -75 17963 -29
rect 18021 -75 18067 -29
rect 18125 -75 18171 -29
rect 18229 -75 18275 -29
rect 18333 -75 18379 -29
rect 18437 -75 18483 -29
rect 18541 -75 18587 -29
rect 18645 -75 18691 -29
rect 18749 -75 18795 -29
rect 18853 -75 18899 -29
rect 18957 -75 19003 -29
rect 19061 -75 19107 -29
rect 19165 -75 19211 -29
rect 19269 -75 19315 -29
rect 19373 -75 19419 -29
rect 19477 -75 19523 -29
rect 19581 -75 19627 -29
rect 19685 -75 19731 -29
rect 19789 -75 19835 -29
rect 19893 -75 19939 -29
rect 19997 -75 20043 -29
rect 20101 -75 20147 -29
rect 20205 -75 20251 -29
rect 20309 -75 20355 -29
rect 20413 -75 20459 -29
rect 20517 -75 20563 -29
rect 20621 -75 20667 -29
rect 20725 -75 20771 -29
rect 20829 -75 20875 -29
rect 20933 -75 20979 -29
rect 21037 -75 21083 -29
rect 21141 -75 21187 -29
rect 21245 -75 21291 -29
rect 21349 -75 21395 -29
rect 21453 -75 21499 -29
rect 21557 -75 21603 -29
rect 21661 -75 21707 -29
rect 21765 -75 21811 -29
rect 21869 -75 21915 -29
rect 21973 -75 22019 -29
rect 22077 -75 22123 -29
rect 22181 -75 22227 -29
rect 22285 -75 22331 -29
rect 22389 -75 22435 -29
rect 22493 -75 22539 -29
rect 22597 -75 22643 -29
rect 22701 -75 22747 -29
rect 22805 -75 22851 -29
rect 22909 -75 22955 -29
rect 23013 -75 23059 -29
rect 23117 -75 23163 -29
rect 23221 -75 23267 -29
rect 23325 -75 23371 -29
rect 23429 -75 23475 -29
rect 23533 -75 23579 -29
rect 23637 -75 23683 -29
rect 23741 -75 23787 -29
rect 23845 -75 23891 -29
rect 23949 -75 23995 -29
rect 24053 -75 24099 -29
rect 24157 -75 24203 -29
rect 24261 -75 24307 -29
rect 24365 -75 24411 -29
rect 24469 -75 24515 -29
rect 24573 -75 24619 -29
rect 24677 -75 24723 -29
rect 24781 -75 24827 -29
rect 24885 -75 24931 -29
rect 24989 -75 25035 -29
rect 25093 -75 25139 -29
rect 25197 -75 25243 -29
rect 25301 -75 25347 -29
rect 25405 -75 25451 -29
rect 25509 -75 25555 -29
rect 25613 -75 25659 -29
rect 25717 -75 25763 -29
rect 25821 -75 25867 -29
rect 25925 -75 25971 -29
rect 26029 -75 26075 -29
rect 26133 -75 26179 -29
rect 26237 -75 26283 -29
rect 26341 -75 26387 -29
rect 26445 -75 26491 -29
rect 26549 -75 26595 -29
rect 26653 -75 26699 -29
rect 26757 -75 26803 -29
rect 26861 -75 26907 -29
rect 26965 -75 27011 -29
rect 27069 -75 27115 -29
rect 27173 -75 27219 -29
rect 27277 -75 27323 -29
rect 27381 -75 27427 -29
rect 27485 -75 27531 -29
rect 27589 -75 27635 -29
rect 27693 -75 27739 -29
rect 27797 -75 27843 -29
rect 27901 -75 27947 -29
rect 28005 -75 28051 -29
rect 28109 -75 28155 -29
rect 28213 -75 28259 -29
<< metal1 >>
rect -28270 75 28270 86
rect -28270 29 -28259 75
rect -28213 29 -28155 75
rect -28109 29 -28051 75
rect -28005 29 -27947 75
rect -27901 29 -27843 75
rect -27797 29 -27739 75
rect -27693 29 -27635 75
rect -27589 29 -27531 75
rect -27485 29 -27427 75
rect -27381 29 -27323 75
rect -27277 29 -27219 75
rect -27173 29 -27115 75
rect -27069 29 -27011 75
rect -26965 29 -26907 75
rect -26861 29 -26803 75
rect -26757 29 -26699 75
rect -26653 29 -26595 75
rect -26549 29 -26491 75
rect -26445 29 -26387 75
rect -26341 29 -26283 75
rect -26237 29 -26179 75
rect -26133 29 -26075 75
rect -26029 29 -25971 75
rect -25925 29 -25867 75
rect -25821 29 -25763 75
rect -25717 29 -25659 75
rect -25613 29 -25555 75
rect -25509 29 -25451 75
rect -25405 29 -25347 75
rect -25301 29 -25243 75
rect -25197 29 -25139 75
rect -25093 29 -25035 75
rect -24989 29 -24931 75
rect -24885 29 -24827 75
rect -24781 29 -24723 75
rect -24677 29 -24619 75
rect -24573 29 -24515 75
rect -24469 29 -24411 75
rect -24365 29 -24307 75
rect -24261 29 -24203 75
rect -24157 29 -24099 75
rect -24053 29 -23995 75
rect -23949 29 -23891 75
rect -23845 29 -23787 75
rect -23741 29 -23683 75
rect -23637 29 -23579 75
rect -23533 29 -23475 75
rect -23429 29 -23371 75
rect -23325 29 -23267 75
rect -23221 29 -23163 75
rect -23117 29 -23059 75
rect -23013 29 -22955 75
rect -22909 29 -22851 75
rect -22805 29 -22747 75
rect -22701 29 -22643 75
rect -22597 29 -22539 75
rect -22493 29 -22435 75
rect -22389 29 -22331 75
rect -22285 29 -22227 75
rect -22181 29 -22123 75
rect -22077 29 -22019 75
rect -21973 29 -21915 75
rect -21869 29 -21811 75
rect -21765 29 -21707 75
rect -21661 29 -21603 75
rect -21557 29 -21499 75
rect -21453 29 -21395 75
rect -21349 29 -21291 75
rect -21245 29 -21187 75
rect -21141 29 -21083 75
rect -21037 29 -20979 75
rect -20933 29 -20875 75
rect -20829 29 -20771 75
rect -20725 29 -20667 75
rect -20621 29 -20563 75
rect -20517 29 -20459 75
rect -20413 29 -20355 75
rect -20309 29 -20251 75
rect -20205 29 -20147 75
rect -20101 29 -20043 75
rect -19997 29 -19939 75
rect -19893 29 -19835 75
rect -19789 29 -19731 75
rect -19685 29 -19627 75
rect -19581 29 -19523 75
rect -19477 29 -19419 75
rect -19373 29 -19315 75
rect -19269 29 -19211 75
rect -19165 29 -19107 75
rect -19061 29 -19003 75
rect -18957 29 -18899 75
rect -18853 29 -18795 75
rect -18749 29 -18691 75
rect -18645 29 -18587 75
rect -18541 29 -18483 75
rect -18437 29 -18379 75
rect -18333 29 -18275 75
rect -18229 29 -18171 75
rect -18125 29 -18067 75
rect -18021 29 -17963 75
rect -17917 29 -17859 75
rect -17813 29 -17755 75
rect -17709 29 -17651 75
rect -17605 29 -17547 75
rect -17501 29 -17443 75
rect -17397 29 -17339 75
rect -17293 29 -17235 75
rect -17189 29 -17131 75
rect -17085 29 -17027 75
rect -16981 29 -16923 75
rect -16877 29 -16819 75
rect -16773 29 -16715 75
rect -16669 29 -16611 75
rect -16565 29 -16507 75
rect -16461 29 -16403 75
rect -16357 29 -16299 75
rect -16253 29 -16195 75
rect -16149 29 -16091 75
rect -16045 29 -15987 75
rect -15941 29 -15883 75
rect -15837 29 -15779 75
rect -15733 29 -15675 75
rect -15629 29 -15571 75
rect -15525 29 -15467 75
rect -15421 29 -15363 75
rect -15317 29 -15259 75
rect -15213 29 -15155 75
rect -15109 29 -15051 75
rect -15005 29 -14947 75
rect -14901 29 -14843 75
rect -14797 29 -14739 75
rect -14693 29 -14635 75
rect -14589 29 -14531 75
rect -14485 29 -14427 75
rect -14381 29 -14323 75
rect -14277 29 -14219 75
rect -14173 29 -14115 75
rect -14069 29 -14011 75
rect -13965 29 -13907 75
rect -13861 29 -13803 75
rect -13757 29 -13699 75
rect -13653 29 -13595 75
rect -13549 29 -13491 75
rect -13445 29 -13387 75
rect -13341 29 -13283 75
rect -13237 29 -13179 75
rect -13133 29 -13075 75
rect -13029 29 -12971 75
rect -12925 29 -12867 75
rect -12821 29 -12763 75
rect -12717 29 -12659 75
rect -12613 29 -12555 75
rect -12509 29 -12451 75
rect -12405 29 -12347 75
rect -12301 29 -12243 75
rect -12197 29 -12139 75
rect -12093 29 -12035 75
rect -11989 29 -11931 75
rect -11885 29 -11827 75
rect -11781 29 -11723 75
rect -11677 29 -11619 75
rect -11573 29 -11515 75
rect -11469 29 -11411 75
rect -11365 29 -11307 75
rect -11261 29 -11203 75
rect -11157 29 -11099 75
rect -11053 29 -10995 75
rect -10949 29 -10891 75
rect -10845 29 -10787 75
rect -10741 29 -10683 75
rect -10637 29 -10579 75
rect -10533 29 -10475 75
rect -10429 29 -10371 75
rect -10325 29 -10267 75
rect -10221 29 -10163 75
rect -10117 29 -10059 75
rect -10013 29 -9955 75
rect -9909 29 -9851 75
rect -9805 29 -9747 75
rect -9701 29 -9643 75
rect -9597 29 -9539 75
rect -9493 29 -9435 75
rect -9389 29 -9331 75
rect -9285 29 -9227 75
rect -9181 29 -9123 75
rect -9077 29 -9019 75
rect -8973 29 -8915 75
rect -8869 29 -8811 75
rect -8765 29 -8707 75
rect -8661 29 -8603 75
rect -8557 29 -8499 75
rect -8453 29 -8395 75
rect -8349 29 -8291 75
rect -8245 29 -8187 75
rect -8141 29 -8083 75
rect -8037 29 -7979 75
rect -7933 29 -7875 75
rect -7829 29 -7771 75
rect -7725 29 -7667 75
rect -7621 29 -7563 75
rect -7517 29 -7459 75
rect -7413 29 -7355 75
rect -7309 29 -7251 75
rect -7205 29 -7147 75
rect -7101 29 -7043 75
rect -6997 29 -6939 75
rect -6893 29 -6835 75
rect -6789 29 -6731 75
rect -6685 29 -6627 75
rect -6581 29 -6523 75
rect -6477 29 -6419 75
rect -6373 29 -6315 75
rect -6269 29 -6211 75
rect -6165 29 -6107 75
rect -6061 29 -6003 75
rect -5957 29 -5899 75
rect -5853 29 -5795 75
rect -5749 29 -5691 75
rect -5645 29 -5587 75
rect -5541 29 -5483 75
rect -5437 29 -5379 75
rect -5333 29 -5275 75
rect -5229 29 -5171 75
rect -5125 29 -5067 75
rect -5021 29 -4963 75
rect -4917 29 -4859 75
rect -4813 29 -4755 75
rect -4709 29 -4651 75
rect -4605 29 -4547 75
rect -4501 29 -4443 75
rect -4397 29 -4339 75
rect -4293 29 -4235 75
rect -4189 29 -4131 75
rect -4085 29 -4027 75
rect -3981 29 -3923 75
rect -3877 29 -3819 75
rect -3773 29 -3715 75
rect -3669 29 -3611 75
rect -3565 29 -3507 75
rect -3461 29 -3403 75
rect -3357 29 -3299 75
rect -3253 29 -3195 75
rect -3149 29 -3091 75
rect -3045 29 -2987 75
rect -2941 29 -2883 75
rect -2837 29 -2779 75
rect -2733 29 -2675 75
rect -2629 29 -2571 75
rect -2525 29 -2467 75
rect -2421 29 -2363 75
rect -2317 29 -2259 75
rect -2213 29 -2155 75
rect -2109 29 -2051 75
rect -2005 29 -1947 75
rect -1901 29 -1843 75
rect -1797 29 -1739 75
rect -1693 29 -1635 75
rect -1589 29 -1531 75
rect -1485 29 -1427 75
rect -1381 29 -1323 75
rect -1277 29 -1219 75
rect -1173 29 -1115 75
rect -1069 29 -1011 75
rect -965 29 -907 75
rect -861 29 -803 75
rect -757 29 -699 75
rect -653 29 -595 75
rect -549 29 -491 75
rect -445 29 -387 75
rect -341 29 -283 75
rect -237 29 -179 75
rect -133 29 -75 75
rect -29 29 29 75
rect 75 29 133 75
rect 179 29 237 75
rect 283 29 341 75
rect 387 29 445 75
rect 491 29 549 75
rect 595 29 653 75
rect 699 29 757 75
rect 803 29 861 75
rect 907 29 965 75
rect 1011 29 1069 75
rect 1115 29 1173 75
rect 1219 29 1277 75
rect 1323 29 1381 75
rect 1427 29 1485 75
rect 1531 29 1589 75
rect 1635 29 1693 75
rect 1739 29 1797 75
rect 1843 29 1901 75
rect 1947 29 2005 75
rect 2051 29 2109 75
rect 2155 29 2213 75
rect 2259 29 2317 75
rect 2363 29 2421 75
rect 2467 29 2525 75
rect 2571 29 2629 75
rect 2675 29 2733 75
rect 2779 29 2837 75
rect 2883 29 2941 75
rect 2987 29 3045 75
rect 3091 29 3149 75
rect 3195 29 3253 75
rect 3299 29 3357 75
rect 3403 29 3461 75
rect 3507 29 3565 75
rect 3611 29 3669 75
rect 3715 29 3773 75
rect 3819 29 3877 75
rect 3923 29 3981 75
rect 4027 29 4085 75
rect 4131 29 4189 75
rect 4235 29 4293 75
rect 4339 29 4397 75
rect 4443 29 4501 75
rect 4547 29 4605 75
rect 4651 29 4709 75
rect 4755 29 4813 75
rect 4859 29 4917 75
rect 4963 29 5021 75
rect 5067 29 5125 75
rect 5171 29 5229 75
rect 5275 29 5333 75
rect 5379 29 5437 75
rect 5483 29 5541 75
rect 5587 29 5645 75
rect 5691 29 5749 75
rect 5795 29 5853 75
rect 5899 29 5957 75
rect 6003 29 6061 75
rect 6107 29 6165 75
rect 6211 29 6269 75
rect 6315 29 6373 75
rect 6419 29 6477 75
rect 6523 29 6581 75
rect 6627 29 6685 75
rect 6731 29 6789 75
rect 6835 29 6893 75
rect 6939 29 6997 75
rect 7043 29 7101 75
rect 7147 29 7205 75
rect 7251 29 7309 75
rect 7355 29 7413 75
rect 7459 29 7517 75
rect 7563 29 7621 75
rect 7667 29 7725 75
rect 7771 29 7829 75
rect 7875 29 7933 75
rect 7979 29 8037 75
rect 8083 29 8141 75
rect 8187 29 8245 75
rect 8291 29 8349 75
rect 8395 29 8453 75
rect 8499 29 8557 75
rect 8603 29 8661 75
rect 8707 29 8765 75
rect 8811 29 8869 75
rect 8915 29 8973 75
rect 9019 29 9077 75
rect 9123 29 9181 75
rect 9227 29 9285 75
rect 9331 29 9389 75
rect 9435 29 9493 75
rect 9539 29 9597 75
rect 9643 29 9701 75
rect 9747 29 9805 75
rect 9851 29 9909 75
rect 9955 29 10013 75
rect 10059 29 10117 75
rect 10163 29 10221 75
rect 10267 29 10325 75
rect 10371 29 10429 75
rect 10475 29 10533 75
rect 10579 29 10637 75
rect 10683 29 10741 75
rect 10787 29 10845 75
rect 10891 29 10949 75
rect 10995 29 11053 75
rect 11099 29 11157 75
rect 11203 29 11261 75
rect 11307 29 11365 75
rect 11411 29 11469 75
rect 11515 29 11573 75
rect 11619 29 11677 75
rect 11723 29 11781 75
rect 11827 29 11885 75
rect 11931 29 11989 75
rect 12035 29 12093 75
rect 12139 29 12197 75
rect 12243 29 12301 75
rect 12347 29 12405 75
rect 12451 29 12509 75
rect 12555 29 12613 75
rect 12659 29 12717 75
rect 12763 29 12821 75
rect 12867 29 12925 75
rect 12971 29 13029 75
rect 13075 29 13133 75
rect 13179 29 13237 75
rect 13283 29 13341 75
rect 13387 29 13445 75
rect 13491 29 13549 75
rect 13595 29 13653 75
rect 13699 29 13757 75
rect 13803 29 13861 75
rect 13907 29 13965 75
rect 14011 29 14069 75
rect 14115 29 14173 75
rect 14219 29 14277 75
rect 14323 29 14381 75
rect 14427 29 14485 75
rect 14531 29 14589 75
rect 14635 29 14693 75
rect 14739 29 14797 75
rect 14843 29 14901 75
rect 14947 29 15005 75
rect 15051 29 15109 75
rect 15155 29 15213 75
rect 15259 29 15317 75
rect 15363 29 15421 75
rect 15467 29 15525 75
rect 15571 29 15629 75
rect 15675 29 15733 75
rect 15779 29 15837 75
rect 15883 29 15941 75
rect 15987 29 16045 75
rect 16091 29 16149 75
rect 16195 29 16253 75
rect 16299 29 16357 75
rect 16403 29 16461 75
rect 16507 29 16565 75
rect 16611 29 16669 75
rect 16715 29 16773 75
rect 16819 29 16877 75
rect 16923 29 16981 75
rect 17027 29 17085 75
rect 17131 29 17189 75
rect 17235 29 17293 75
rect 17339 29 17397 75
rect 17443 29 17501 75
rect 17547 29 17605 75
rect 17651 29 17709 75
rect 17755 29 17813 75
rect 17859 29 17917 75
rect 17963 29 18021 75
rect 18067 29 18125 75
rect 18171 29 18229 75
rect 18275 29 18333 75
rect 18379 29 18437 75
rect 18483 29 18541 75
rect 18587 29 18645 75
rect 18691 29 18749 75
rect 18795 29 18853 75
rect 18899 29 18957 75
rect 19003 29 19061 75
rect 19107 29 19165 75
rect 19211 29 19269 75
rect 19315 29 19373 75
rect 19419 29 19477 75
rect 19523 29 19581 75
rect 19627 29 19685 75
rect 19731 29 19789 75
rect 19835 29 19893 75
rect 19939 29 19997 75
rect 20043 29 20101 75
rect 20147 29 20205 75
rect 20251 29 20309 75
rect 20355 29 20413 75
rect 20459 29 20517 75
rect 20563 29 20621 75
rect 20667 29 20725 75
rect 20771 29 20829 75
rect 20875 29 20933 75
rect 20979 29 21037 75
rect 21083 29 21141 75
rect 21187 29 21245 75
rect 21291 29 21349 75
rect 21395 29 21453 75
rect 21499 29 21557 75
rect 21603 29 21661 75
rect 21707 29 21765 75
rect 21811 29 21869 75
rect 21915 29 21973 75
rect 22019 29 22077 75
rect 22123 29 22181 75
rect 22227 29 22285 75
rect 22331 29 22389 75
rect 22435 29 22493 75
rect 22539 29 22597 75
rect 22643 29 22701 75
rect 22747 29 22805 75
rect 22851 29 22909 75
rect 22955 29 23013 75
rect 23059 29 23117 75
rect 23163 29 23221 75
rect 23267 29 23325 75
rect 23371 29 23429 75
rect 23475 29 23533 75
rect 23579 29 23637 75
rect 23683 29 23741 75
rect 23787 29 23845 75
rect 23891 29 23949 75
rect 23995 29 24053 75
rect 24099 29 24157 75
rect 24203 29 24261 75
rect 24307 29 24365 75
rect 24411 29 24469 75
rect 24515 29 24573 75
rect 24619 29 24677 75
rect 24723 29 24781 75
rect 24827 29 24885 75
rect 24931 29 24989 75
rect 25035 29 25093 75
rect 25139 29 25197 75
rect 25243 29 25301 75
rect 25347 29 25405 75
rect 25451 29 25509 75
rect 25555 29 25613 75
rect 25659 29 25717 75
rect 25763 29 25821 75
rect 25867 29 25925 75
rect 25971 29 26029 75
rect 26075 29 26133 75
rect 26179 29 26237 75
rect 26283 29 26341 75
rect 26387 29 26445 75
rect 26491 29 26549 75
rect 26595 29 26653 75
rect 26699 29 26757 75
rect 26803 29 26861 75
rect 26907 29 26965 75
rect 27011 29 27069 75
rect 27115 29 27173 75
rect 27219 29 27277 75
rect 27323 29 27381 75
rect 27427 29 27485 75
rect 27531 29 27589 75
rect 27635 29 27693 75
rect 27739 29 27797 75
rect 27843 29 27901 75
rect 27947 29 28005 75
rect 28051 29 28109 75
rect 28155 29 28213 75
rect 28259 29 28270 75
rect -28270 -29 28270 29
rect -28270 -75 -28259 -29
rect -28213 -75 -28155 -29
rect -28109 -75 -28051 -29
rect -28005 -75 -27947 -29
rect -27901 -75 -27843 -29
rect -27797 -75 -27739 -29
rect -27693 -75 -27635 -29
rect -27589 -75 -27531 -29
rect -27485 -75 -27427 -29
rect -27381 -75 -27323 -29
rect -27277 -75 -27219 -29
rect -27173 -75 -27115 -29
rect -27069 -75 -27011 -29
rect -26965 -75 -26907 -29
rect -26861 -75 -26803 -29
rect -26757 -75 -26699 -29
rect -26653 -75 -26595 -29
rect -26549 -75 -26491 -29
rect -26445 -75 -26387 -29
rect -26341 -75 -26283 -29
rect -26237 -75 -26179 -29
rect -26133 -75 -26075 -29
rect -26029 -75 -25971 -29
rect -25925 -75 -25867 -29
rect -25821 -75 -25763 -29
rect -25717 -75 -25659 -29
rect -25613 -75 -25555 -29
rect -25509 -75 -25451 -29
rect -25405 -75 -25347 -29
rect -25301 -75 -25243 -29
rect -25197 -75 -25139 -29
rect -25093 -75 -25035 -29
rect -24989 -75 -24931 -29
rect -24885 -75 -24827 -29
rect -24781 -75 -24723 -29
rect -24677 -75 -24619 -29
rect -24573 -75 -24515 -29
rect -24469 -75 -24411 -29
rect -24365 -75 -24307 -29
rect -24261 -75 -24203 -29
rect -24157 -75 -24099 -29
rect -24053 -75 -23995 -29
rect -23949 -75 -23891 -29
rect -23845 -75 -23787 -29
rect -23741 -75 -23683 -29
rect -23637 -75 -23579 -29
rect -23533 -75 -23475 -29
rect -23429 -75 -23371 -29
rect -23325 -75 -23267 -29
rect -23221 -75 -23163 -29
rect -23117 -75 -23059 -29
rect -23013 -75 -22955 -29
rect -22909 -75 -22851 -29
rect -22805 -75 -22747 -29
rect -22701 -75 -22643 -29
rect -22597 -75 -22539 -29
rect -22493 -75 -22435 -29
rect -22389 -75 -22331 -29
rect -22285 -75 -22227 -29
rect -22181 -75 -22123 -29
rect -22077 -75 -22019 -29
rect -21973 -75 -21915 -29
rect -21869 -75 -21811 -29
rect -21765 -75 -21707 -29
rect -21661 -75 -21603 -29
rect -21557 -75 -21499 -29
rect -21453 -75 -21395 -29
rect -21349 -75 -21291 -29
rect -21245 -75 -21187 -29
rect -21141 -75 -21083 -29
rect -21037 -75 -20979 -29
rect -20933 -75 -20875 -29
rect -20829 -75 -20771 -29
rect -20725 -75 -20667 -29
rect -20621 -75 -20563 -29
rect -20517 -75 -20459 -29
rect -20413 -75 -20355 -29
rect -20309 -75 -20251 -29
rect -20205 -75 -20147 -29
rect -20101 -75 -20043 -29
rect -19997 -75 -19939 -29
rect -19893 -75 -19835 -29
rect -19789 -75 -19731 -29
rect -19685 -75 -19627 -29
rect -19581 -75 -19523 -29
rect -19477 -75 -19419 -29
rect -19373 -75 -19315 -29
rect -19269 -75 -19211 -29
rect -19165 -75 -19107 -29
rect -19061 -75 -19003 -29
rect -18957 -75 -18899 -29
rect -18853 -75 -18795 -29
rect -18749 -75 -18691 -29
rect -18645 -75 -18587 -29
rect -18541 -75 -18483 -29
rect -18437 -75 -18379 -29
rect -18333 -75 -18275 -29
rect -18229 -75 -18171 -29
rect -18125 -75 -18067 -29
rect -18021 -75 -17963 -29
rect -17917 -75 -17859 -29
rect -17813 -75 -17755 -29
rect -17709 -75 -17651 -29
rect -17605 -75 -17547 -29
rect -17501 -75 -17443 -29
rect -17397 -75 -17339 -29
rect -17293 -75 -17235 -29
rect -17189 -75 -17131 -29
rect -17085 -75 -17027 -29
rect -16981 -75 -16923 -29
rect -16877 -75 -16819 -29
rect -16773 -75 -16715 -29
rect -16669 -75 -16611 -29
rect -16565 -75 -16507 -29
rect -16461 -75 -16403 -29
rect -16357 -75 -16299 -29
rect -16253 -75 -16195 -29
rect -16149 -75 -16091 -29
rect -16045 -75 -15987 -29
rect -15941 -75 -15883 -29
rect -15837 -75 -15779 -29
rect -15733 -75 -15675 -29
rect -15629 -75 -15571 -29
rect -15525 -75 -15467 -29
rect -15421 -75 -15363 -29
rect -15317 -75 -15259 -29
rect -15213 -75 -15155 -29
rect -15109 -75 -15051 -29
rect -15005 -75 -14947 -29
rect -14901 -75 -14843 -29
rect -14797 -75 -14739 -29
rect -14693 -75 -14635 -29
rect -14589 -75 -14531 -29
rect -14485 -75 -14427 -29
rect -14381 -75 -14323 -29
rect -14277 -75 -14219 -29
rect -14173 -75 -14115 -29
rect -14069 -75 -14011 -29
rect -13965 -75 -13907 -29
rect -13861 -75 -13803 -29
rect -13757 -75 -13699 -29
rect -13653 -75 -13595 -29
rect -13549 -75 -13491 -29
rect -13445 -75 -13387 -29
rect -13341 -75 -13283 -29
rect -13237 -75 -13179 -29
rect -13133 -75 -13075 -29
rect -13029 -75 -12971 -29
rect -12925 -75 -12867 -29
rect -12821 -75 -12763 -29
rect -12717 -75 -12659 -29
rect -12613 -75 -12555 -29
rect -12509 -75 -12451 -29
rect -12405 -75 -12347 -29
rect -12301 -75 -12243 -29
rect -12197 -75 -12139 -29
rect -12093 -75 -12035 -29
rect -11989 -75 -11931 -29
rect -11885 -75 -11827 -29
rect -11781 -75 -11723 -29
rect -11677 -75 -11619 -29
rect -11573 -75 -11515 -29
rect -11469 -75 -11411 -29
rect -11365 -75 -11307 -29
rect -11261 -75 -11203 -29
rect -11157 -75 -11099 -29
rect -11053 -75 -10995 -29
rect -10949 -75 -10891 -29
rect -10845 -75 -10787 -29
rect -10741 -75 -10683 -29
rect -10637 -75 -10579 -29
rect -10533 -75 -10475 -29
rect -10429 -75 -10371 -29
rect -10325 -75 -10267 -29
rect -10221 -75 -10163 -29
rect -10117 -75 -10059 -29
rect -10013 -75 -9955 -29
rect -9909 -75 -9851 -29
rect -9805 -75 -9747 -29
rect -9701 -75 -9643 -29
rect -9597 -75 -9539 -29
rect -9493 -75 -9435 -29
rect -9389 -75 -9331 -29
rect -9285 -75 -9227 -29
rect -9181 -75 -9123 -29
rect -9077 -75 -9019 -29
rect -8973 -75 -8915 -29
rect -8869 -75 -8811 -29
rect -8765 -75 -8707 -29
rect -8661 -75 -8603 -29
rect -8557 -75 -8499 -29
rect -8453 -75 -8395 -29
rect -8349 -75 -8291 -29
rect -8245 -75 -8187 -29
rect -8141 -75 -8083 -29
rect -8037 -75 -7979 -29
rect -7933 -75 -7875 -29
rect -7829 -75 -7771 -29
rect -7725 -75 -7667 -29
rect -7621 -75 -7563 -29
rect -7517 -75 -7459 -29
rect -7413 -75 -7355 -29
rect -7309 -75 -7251 -29
rect -7205 -75 -7147 -29
rect -7101 -75 -7043 -29
rect -6997 -75 -6939 -29
rect -6893 -75 -6835 -29
rect -6789 -75 -6731 -29
rect -6685 -75 -6627 -29
rect -6581 -75 -6523 -29
rect -6477 -75 -6419 -29
rect -6373 -75 -6315 -29
rect -6269 -75 -6211 -29
rect -6165 -75 -6107 -29
rect -6061 -75 -6003 -29
rect -5957 -75 -5899 -29
rect -5853 -75 -5795 -29
rect -5749 -75 -5691 -29
rect -5645 -75 -5587 -29
rect -5541 -75 -5483 -29
rect -5437 -75 -5379 -29
rect -5333 -75 -5275 -29
rect -5229 -75 -5171 -29
rect -5125 -75 -5067 -29
rect -5021 -75 -4963 -29
rect -4917 -75 -4859 -29
rect -4813 -75 -4755 -29
rect -4709 -75 -4651 -29
rect -4605 -75 -4547 -29
rect -4501 -75 -4443 -29
rect -4397 -75 -4339 -29
rect -4293 -75 -4235 -29
rect -4189 -75 -4131 -29
rect -4085 -75 -4027 -29
rect -3981 -75 -3923 -29
rect -3877 -75 -3819 -29
rect -3773 -75 -3715 -29
rect -3669 -75 -3611 -29
rect -3565 -75 -3507 -29
rect -3461 -75 -3403 -29
rect -3357 -75 -3299 -29
rect -3253 -75 -3195 -29
rect -3149 -75 -3091 -29
rect -3045 -75 -2987 -29
rect -2941 -75 -2883 -29
rect -2837 -75 -2779 -29
rect -2733 -75 -2675 -29
rect -2629 -75 -2571 -29
rect -2525 -75 -2467 -29
rect -2421 -75 -2363 -29
rect -2317 -75 -2259 -29
rect -2213 -75 -2155 -29
rect -2109 -75 -2051 -29
rect -2005 -75 -1947 -29
rect -1901 -75 -1843 -29
rect -1797 -75 -1739 -29
rect -1693 -75 -1635 -29
rect -1589 -75 -1531 -29
rect -1485 -75 -1427 -29
rect -1381 -75 -1323 -29
rect -1277 -75 -1219 -29
rect -1173 -75 -1115 -29
rect -1069 -75 -1011 -29
rect -965 -75 -907 -29
rect -861 -75 -803 -29
rect -757 -75 -699 -29
rect -653 -75 -595 -29
rect -549 -75 -491 -29
rect -445 -75 -387 -29
rect -341 -75 -283 -29
rect -237 -75 -179 -29
rect -133 -75 -75 -29
rect -29 -75 29 -29
rect 75 -75 133 -29
rect 179 -75 237 -29
rect 283 -75 341 -29
rect 387 -75 445 -29
rect 491 -75 549 -29
rect 595 -75 653 -29
rect 699 -75 757 -29
rect 803 -75 861 -29
rect 907 -75 965 -29
rect 1011 -75 1069 -29
rect 1115 -75 1173 -29
rect 1219 -75 1277 -29
rect 1323 -75 1381 -29
rect 1427 -75 1485 -29
rect 1531 -75 1589 -29
rect 1635 -75 1693 -29
rect 1739 -75 1797 -29
rect 1843 -75 1901 -29
rect 1947 -75 2005 -29
rect 2051 -75 2109 -29
rect 2155 -75 2213 -29
rect 2259 -75 2317 -29
rect 2363 -75 2421 -29
rect 2467 -75 2525 -29
rect 2571 -75 2629 -29
rect 2675 -75 2733 -29
rect 2779 -75 2837 -29
rect 2883 -75 2941 -29
rect 2987 -75 3045 -29
rect 3091 -75 3149 -29
rect 3195 -75 3253 -29
rect 3299 -75 3357 -29
rect 3403 -75 3461 -29
rect 3507 -75 3565 -29
rect 3611 -75 3669 -29
rect 3715 -75 3773 -29
rect 3819 -75 3877 -29
rect 3923 -75 3981 -29
rect 4027 -75 4085 -29
rect 4131 -75 4189 -29
rect 4235 -75 4293 -29
rect 4339 -75 4397 -29
rect 4443 -75 4501 -29
rect 4547 -75 4605 -29
rect 4651 -75 4709 -29
rect 4755 -75 4813 -29
rect 4859 -75 4917 -29
rect 4963 -75 5021 -29
rect 5067 -75 5125 -29
rect 5171 -75 5229 -29
rect 5275 -75 5333 -29
rect 5379 -75 5437 -29
rect 5483 -75 5541 -29
rect 5587 -75 5645 -29
rect 5691 -75 5749 -29
rect 5795 -75 5853 -29
rect 5899 -75 5957 -29
rect 6003 -75 6061 -29
rect 6107 -75 6165 -29
rect 6211 -75 6269 -29
rect 6315 -75 6373 -29
rect 6419 -75 6477 -29
rect 6523 -75 6581 -29
rect 6627 -75 6685 -29
rect 6731 -75 6789 -29
rect 6835 -75 6893 -29
rect 6939 -75 6997 -29
rect 7043 -75 7101 -29
rect 7147 -75 7205 -29
rect 7251 -75 7309 -29
rect 7355 -75 7413 -29
rect 7459 -75 7517 -29
rect 7563 -75 7621 -29
rect 7667 -75 7725 -29
rect 7771 -75 7829 -29
rect 7875 -75 7933 -29
rect 7979 -75 8037 -29
rect 8083 -75 8141 -29
rect 8187 -75 8245 -29
rect 8291 -75 8349 -29
rect 8395 -75 8453 -29
rect 8499 -75 8557 -29
rect 8603 -75 8661 -29
rect 8707 -75 8765 -29
rect 8811 -75 8869 -29
rect 8915 -75 8973 -29
rect 9019 -75 9077 -29
rect 9123 -75 9181 -29
rect 9227 -75 9285 -29
rect 9331 -75 9389 -29
rect 9435 -75 9493 -29
rect 9539 -75 9597 -29
rect 9643 -75 9701 -29
rect 9747 -75 9805 -29
rect 9851 -75 9909 -29
rect 9955 -75 10013 -29
rect 10059 -75 10117 -29
rect 10163 -75 10221 -29
rect 10267 -75 10325 -29
rect 10371 -75 10429 -29
rect 10475 -75 10533 -29
rect 10579 -75 10637 -29
rect 10683 -75 10741 -29
rect 10787 -75 10845 -29
rect 10891 -75 10949 -29
rect 10995 -75 11053 -29
rect 11099 -75 11157 -29
rect 11203 -75 11261 -29
rect 11307 -75 11365 -29
rect 11411 -75 11469 -29
rect 11515 -75 11573 -29
rect 11619 -75 11677 -29
rect 11723 -75 11781 -29
rect 11827 -75 11885 -29
rect 11931 -75 11989 -29
rect 12035 -75 12093 -29
rect 12139 -75 12197 -29
rect 12243 -75 12301 -29
rect 12347 -75 12405 -29
rect 12451 -75 12509 -29
rect 12555 -75 12613 -29
rect 12659 -75 12717 -29
rect 12763 -75 12821 -29
rect 12867 -75 12925 -29
rect 12971 -75 13029 -29
rect 13075 -75 13133 -29
rect 13179 -75 13237 -29
rect 13283 -75 13341 -29
rect 13387 -75 13445 -29
rect 13491 -75 13549 -29
rect 13595 -75 13653 -29
rect 13699 -75 13757 -29
rect 13803 -75 13861 -29
rect 13907 -75 13965 -29
rect 14011 -75 14069 -29
rect 14115 -75 14173 -29
rect 14219 -75 14277 -29
rect 14323 -75 14381 -29
rect 14427 -75 14485 -29
rect 14531 -75 14589 -29
rect 14635 -75 14693 -29
rect 14739 -75 14797 -29
rect 14843 -75 14901 -29
rect 14947 -75 15005 -29
rect 15051 -75 15109 -29
rect 15155 -75 15213 -29
rect 15259 -75 15317 -29
rect 15363 -75 15421 -29
rect 15467 -75 15525 -29
rect 15571 -75 15629 -29
rect 15675 -75 15733 -29
rect 15779 -75 15837 -29
rect 15883 -75 15941 -29
rect 15987 -75 16045 -29
rect 16091 -75 16149 -29
rect 16195 -75 16253 -29
rect 16299 -75 16357 -29
rect 16403 -75 16461 -29
rect 16507 -75 16565 -29
rect 16611 -75 16669 -29
rect 16715 -75 16773 -29
rect 16819 -75 16877 -29
rect 16923 -75 16981 -29
rect 17027 -75 17085 -29
rect 17131 -75 17189 -29
rect 17235 -75 17293 -29
rect 17339 -75 17397 -29
rect 17443 -75 17501 -29
rect 17547 -75 17605 -29
rect 17651 -75 17709 -29
rect 17755 -75 17813 -29
rect 17859 -75 17917 -29
rect 17963 -75 18021 -29
rect 18067 -75 18125 -29
rect 18171 -75 18229 -29
rect 18275 -75 18333 -29
rect 18379 -75 18437 -29
rect 18483 -75 18541 -29
rect 18587 -75 18645 -29
rect 18691 -75 18749 -29
rect 18795 -75 18853 -29
rect 18899 -75 18957 -29
rect 19003 -75 19061 -29
rect 19107 -75 19165 -29
rect 19211 -75 19269 -29
rect 19315 -75 19373 -29
rect 19419 -75 19477 -29
rect 19523 -75 19581 -29
rect 19627 -75 19685 -29
rect 19731 -75 19789 -29
rect 19835 -75 19893 -29
rect 19939 -75 19997 -29
rect 20043 -75 20101 -29
rect 20147 -75 20205 -29
rect 20251 -75 20309 -29
rect 20355 -75 20413 -29
rect 20459 -75 20517 -29
rect 20563 -75 20621 -29
rect 20667 -75 20725 -29
rect 20771 -75 20829 -29
rect 20875 -75 20933 -29
rect 20979 -75 21037 -29
rect 21083 -75 21141 -29
rect 21187 -75 21245 -29
rect 21291 -75 21349 -29
rect 21395 -75 21453 -29
rect 21499 -75 21557 -29
rect 21603 -75 21661 -29
rect 21707 -75 21765 -29
rect 21811 -75 21869 -29
rect 21915 -75 21973 -29
rect 22019 -75 22077 -29
rect 22123 -75 22181 -29
rect 22227 -75 22285 -29
rect 22331 -75 22389 -29
rect 22435 -75 22493 -29
rect 22539 -75 22597 -29
rect 22643 -75 22701 -29
rect 22747 -75 22805 -29
rect 22851 -75 22909 -29
rect 22955 -75 23013 -29
rect 23059 -75 23117 -29
rect 23163 -75 23221 -29
rect 23267 -75 23325 -29
rect 23371 -75 23429 -29
rect 23475 -75 23533 -29
rect 23579 -75 23637 -29
rect 23683 -75 23741 -29
rect 23787 -75 23845 -29
rect 23891 -75 23949 -29
rect 23995 -75 24053 -29
rect 24099 -75 24157 -29
rect 24203 -75 24261 -29
rect 24307 -75 24365 -29
rect 24411 -75 24469 -29
rect 24515 -75 24573 -29
rect 24619 -75 24677 -29
rect 24723 -75 24781 -29
rect 24827 -75 24885 -29
rect 24931 -75 24989 -29
rect 25035 -75 25093 -29
rect 25139 -75 25197 -29
rect 25243 -75 25301 -29
rect 25347 -75 25405 -29
rect 25451 -75 25509 -29
rect 25555 -75 25613 -29
rect 25659 -75 25717 -29
rect 25763 -75 25821 -29
rect 25867 -75 25925 -29
rect 25971 -75 26029 -29
rect 26075 -75 26133 -29
rect 26179 -75 26237 -29
rect 26283 -75 26341 -29
rect 26387 -75 26445 -29
rect 26491 -75 26549 -29
rect 26595 -75 26653 -29
rect 26699 -75 26757 -29
rect 26803 -75 26861 -29
rect 26907 -75 26965 -29
rect 27011 -75 27069 -29
rect 27115 -75 27173 -29
rect 27219 -75 27277 -29
rect 27323 -75 27381 -29
rect 27427 -75 27485 -29
rect 27531 -75 27589 -29
rect 27635 -75 27693 -29
rect 27739 -75 27797 -29
rect 27843 -75 27901 -29
rect 27947 -75 28005 -29
rect 28051 -75 28109 -29
rect 28155 -75 28213 -29
rect 28259 -75 28270 -29
rect -28270 -86 28270 -75
<< end >>
