magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2216 -2216 2312 2312
<< nwell >>
rect -216 -216 312 312
<< mvnsubdiff >>
rect -168 251 264 264
rect -168 205 -155 251
rect -109 205 -35 251
rect 11 205 85 251
rect 131 205 205 251
rect 251 205 264 251
rect -168 192 264 205
rect -168 131 -96 192
rect -168 85 -155 131
rect -109 85 -96 131
rect 192 131 264 192
rect -168 11 -96 85
rect -168 -35 -155 11
rect -109 -35 -96 11
rect 192 85 205 131
rect 251 85 264 131
rect 192 11 264 85
rect -168 -96 -96 -35
rect 192 -35 205 11
rect 251 -35 264 11
rect 192 -96 264 -35
rect -168 -109 264 -96
rect -168 -155 -155 -109
rect -109 -155 -35 -109
rect 11 -155 85 -109
rect 131 -155 205 -109
rect 251 -155 264 -109
rect -168 -168 264 -155
<< mvnsubdiffcont >>
rect -155 205 -109 251
rect -35 205 11 251
rect 85 205 131 251
rect 205 205 251 251
rect -155 85 -109 131
rect -155 -35 -109 11
rect 205 85 251 131
rect 205 -35 251 11
rect -155 -155 -109 -109
rect -35 -155 11 -109
rect 85 -155 131 -109
rect 205 -155 251 -109
<< mvpdiode >>
rect 0 71 96 96
rect 0 25 25 71
rect 71 25 96 71
rect 0 0 96 25
<< mvpdiodec >>
rect 25 25 71 71
<< metal1 >>
rect -168 251 264 264
rect -168 205 -155 251
rect -109 205 -35 251
rect 11 205 85 251
rect 131 205 205 251
rect 251 205 264 251
rect -168 192 264 205
rect -168 131 -96 192
rect -168 85 -155 131
rect -109 85 -96 131
rect 192 131 264 192
rect -168 11 -96 85
rect -168 -35 -155 11
rect -109 -35 -96 11
rect 0 71 96 96
rect 0 25 25 71
rect 71 25 96 71
rect 0 0 96 25
rect 192 85 205 131
rect 251 85 264 131
rect 192 11 264 85
rect -168 -96 -96 -35
rect 192 -35 205 11
rect 251 -35 264 11
rect 192 -96 264 -35
rect -168 -109 264 -96
rect -168 -155 -155 -109
rect -109 -155 -35 -109
rect 11 -155 85 -109
rect 131 -155 205 -109
rect 251 -155 264 -109
rect -168 -168 264 -155
<< labels >>
rlabel metal1 48 -132 48 -132 4 MINUS
rlabel metal1 48 228 48 228 4 MINUS
rlabel metal1 228 48 228 48 4 MINUS
rlabel metal1 -132 48 -132 48 4 MINUS
rlabel mvpdiodec 48 48 48 48 4 PLUS
<< end >>
