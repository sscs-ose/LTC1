magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1050 -1794 1050 1794
<< metal1 >>
rect -50 788 50 794
rect -50 762 -44 788
rect -18 762 18 788
rect 44 762 50 788
rect -50 726 50 762
rect -50 700 -44 726
rect -18 700 18 726
rect 44 700 50 726
rect -50 664 50 700
rect -50 638 -44 664
rect -18 638 18 664
rect 44 638 50 664
rect -50 602 50 638
rect -50 576 -44 602
rect -18 576 18 602
rect 44 576 50 602
rect -50 540 50 576
rect -50 514 -44 540
rect -18 514 18 540
rect 44 514 50 540
rect -50 478 50 514
rect -50 452 -44 478
rect -18 452 18 478
rect 44 452 50 478
rect -50 416 50 452
rect -50 390 -44 416
rect -18 390 18 416
rect 44 390 50 416
rect -50 354 50 390
rect -50 328 -44 354
rect -18 328 18 354
rect 44 328 50 354
rect -50 292 50 328
rect -50 266 -44 292
rect -18 266 18 292
rect 44 266 50 292
rect -50 230 50 266
rect -50 204 -44 230
rect -18 204 18 230
rect 44 204 50 230
rect -50 168 50 204
rect -50 142 -44 168
rect -18 142 18 168
rect 44 142 50 168
rect -50 106 50 142
rect -50 80 -44 106
rect -18 80 18 106
rect 44 80 50 106
rect -50 44 50 80
rect -50 18 -44 44
rect -18 18 18 44
rect 44 18 50 44
rect -50 -18 50 18
rect -50 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 50 -18
rect -50 -80 50 -44
rect -50 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 50 -80
rect -50 -142 50 -106
rect -50 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 50 -142
rect -50 -204 50 -168
rect -50 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 50 -204
rect -50 -266 50 -230
rect -50 -292 -44 -266
rect -18 -292 18 -266
rect 44 -292 50 -266
rect -50 -328 50 -292
rect -50 -354 -44 -328
rect -18 -354 18 -328
rect 44 -354 50 -328
rect -50 -390 50 -354
rect -50 -416 -44 -390
rect -18 -416 18 -390
rect 44 -416 50 -390
rect -50 -452 50 -416
rect -50 -478 -44 -452
rect -18 -478 18 -452
rect 44 -478 50 -452
rect -50 -514 50 -478
rect -50 -540 -44 -514
rect -18 -540 18 -514
rect 44 -540 50 -514
rect -50 -576 50 -540
rect -50 -602 -44 -576
rect -18 -602 18 -576
rect 44 -602 50 -576
rect -50 -638 50 -602
rect -50 -664 -44 -638
rect -18 -664 18 -638
rect 44 -664 50 -638
rect -50 -700 50 -664
rect -50 -726 -44 -700
rect -18 -726 18 -700
rect 44 -726 50 -700
rect -50 -762 50 -726
rect -50 -788 -44 -762
rect -18 -788 18 -762
rect 44 -788 50 -762
rect -50 -794 50 -788
<< via1 >>
rect -44 762 -18 788
rect 18 762 44 788
rect -44 700 -18 726
rect 18 700 44 726
rect -44 638 -18 664
rect 18 638 44 664
rect -44 576 -18 602
rect 18 576 44 602
rect -44 514 -18 540
rect 18 514 44 540
rect -44 452 -18 478
rect 18 452 44 478
rect -44 390 -18 416
rect 18 390 44 416
rect -44 328 -18 354
rect 18 328 44 354
rect -44 266 -18 292
rect 18 266 44 292
rect -44 204 -18 230
rect 18 204 44 230
rect -44 142 -18 168
rect 18 142 44 168
rect -44 80 -18 106
rect 18 80 44 106
rect -44 18 -18 44
rect 18 18 44 44
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect -44 -106 -18 -80
rect 18 -106 44 -80
rect -44 -168 -18 -142
rect 18 -168 44 -142
rect -44 -230 -18 -204
rect 18 -230 44 -204
rect -44 -292 -18 -266
rect 18 -292 44 -266
rect -44 -354 -18 -328
rect 18 -354 44 -328
rect -44 -416 -18 -390
rect 18 -416 44 -390
rect -44 -478 -18 -452
rect 18 -478 44 -452
rect -44 -540 -18 -514
rect 18 -540 44 -514
rect -44 -602 -18 -576
rect 18 -602 44 -576
rect -44 -664 -18 -638
rect 18 -664 44 -638
rect -44 -726 -18 -700
rect 18 -726 44 -700
rect -44 -788 -18 -762
rect 18 -788 44 -762
<< metal2 >>
rect -50 788 50 794
rect -50 762 -44 788
rect -18 762 18 788
rect 44 762 50 788
rect -50 726 50 762
rect -50 700 -44 726
rect -18 700 18 726
rect 44 700 50 726
rect -50 664 50 700
rect -50 638 -44 664
rect -18 638 18 664
rect 44 638 50 664
rect -50 602 50 638
rect -50 576 -44 602
rect -18 576 18 602
rect 44 576 50 602
rect -50 540 50 576
rect -50 514 -44 540
rect -18 514 18 540
rect 44 514 50 540
rect -50 478 50 514
rect -50 452 -44 478
rect -18 452 18 478
rect 44 452 50 478
rect -50 416 50 452
rect -50 390 -44 416
rect -18 390 18 416
rect 44 390 50 416
rect -50 354 50 390
rect -50 328 -44 354
rect -18 328 18 354
rect 44 328 50 354
rect -50 292 50 328
rect -50 266 -44 292
rect -18 266 18 292
rect 44 266 50 292
rect -50 230 50 266
rect -50 204 -44 230
rect -18 204 18 230
rect 44 204 50 230
rect -50 168 50 204
rect -50 142 -44 168
rect -18 142 18 168
rect 44 142 50 168
rect -50 106 50 142
rect -50 80 -44 106
rect -18 80 18 106
rect 44 80 50 106
rect -50 44 50 80
rect -50 18 -44 44
rect -18 18 18 44
rect 44 18 50 44
rect -50 -18 50 18
rect -50 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 50 -18
rect -50 -80 50 -44
rect -50 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 50 -80
rect -50 -142 50 -106
rect -50 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 50 -142
rect -50 -204 50 -168
rect -50 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 50 -204
rect -50 -266 50 -230
rect -50 -292 -44 -266
rect -18 -292 18 -266
rect 44 -292 50 -266
rect -50 -328 50 -292
rect -50 -354 -44 -328
rect -18 -354 18 -328
rect 44 -354 50 -328
rect -50 -390 50 -354
rect -50 -416 -44 -390
rect -18 -416 18 -390
rect 44 -416 50 -390
rect -50 -452 50 -416
rect -50 -478 -44 -452
rect -18 -478 18 -452
rect 44 -478 50 -452
rect -50 -514 50 -478
rect -50 -540 -44 -514
rect -18 -540 18 -514
rect 44 -540 50 -514
rect -50 -576 50 -540
rect -50 -602 -44 -576
rect -18 -602 18 -576
rect 44 -602 50 -576
rect -50 -638 50 -602
rect -50 -664 -44 -638
rect -18 -664 18 -638
rect 44 -664 50 -638
rect -50 -700 50 -664
rect -50 -726 -44 -700
rect -18 -726 18 -700
rect 44 -726 50 -700
rect -50 -762 50 -726
rect -50 -788 -44 -762
rect -18 -788 18 -762
rect 44 -788 50 -762
rect -50 -794 50 -788
<< end >>
