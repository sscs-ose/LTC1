magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 3032 71968
<< metal4 >>
rect 0 68400 1000 69678
rect 0 66800 1000 68200
rect 0 65200 1000 66600
rect 0 63600 1000 65000
rect 0 62000 1000 63400
rect 0 60400 1000 61800
rect 0 58800 1000 60200
rect 0 57200 1000 58600
rect 0 55600 1000 57000
rect 0 54000 1000 55400
rect 0 52400 1000 53800
rect 0 50800 1000 52200
rect 0 49200 1000 50600
rect 0 46000 1000 49000
rect 0 42800 1000 45800
rect 0 41200 1000 42600
rect 0 39600 1000 41000
rect 0 36400 1000 39400
rect 0 33200 1000 36200
rect 0 30000 1000 33000
rect 0 26800 1000 29800
rect 0 25200 1000 26600
rect 0 23600 1000 25000
rect 0 20400 1000 23400
rect 0 17200 1000 20200
rect 0 14000 1000 17000
<< metal5 >>
rect 0 68400 1000 69678
rect 0 66800 1000 68200
rect 0 65200 1000 66600
rect 0 63600 1000 65000
rect 0 62000 1000 63400
rect 0 60400 1000 61800
rect 0 58800 1000 60200
rect 0 57200 1000 58600
rect 0 55600 1000 57000
rect 0 54000 1000 55400
rect 0 52400 1000 53800
rect 0 50800 1000 52200
rect 0 49200 1000 50600
rect 0 46000 1000 49000
rect 0 42800 1000 45800
rect 0 41200 1000 42600
rect 0 39600 1000 41000
rect 0 36400 1000 39400
rect 0 33200 1000 36200
rect 0 30000 1000 33000
rect 0 26800 1000 29800
rect 0 25200 1000 26600
rect 0 23600 1000 25000
rect 0 20400 1000 23400
rect 0 17200 1000 20200
rect 0 14000 1000 17000
use GF_NI_FILL5_0  GF_NI_FILL5_0_0
timestamp 1713338890
transform 1 0 0 0 1 0
box -32 13097 1032 69968
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_0
timestamp 1713338890
transform 1 0 494 0 1 15521
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_1
timestamp 1713338890
transform 1 0 494 0 1 18694
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_2
timestamp 1713338890
transform 1 0 494 0 1 21905
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_3
timestamp 1713338890
transform 1 0 494 0 1 28293
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_4
timestamp 1713338890
transform 1 0 494 0 1 31510
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_5
timestamp 1713338890
transform 1 0 494 0 1 34702
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_6
timestamp 1713338890
transform 1 0 494 0 1 37912
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_7
timestamp 1713338890
transform 1 0 494 0 1 44305
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316572  M4_M3_CDNS_6903358316572_8
timestamp 1713338890
transform 1 0 494 0 1 47501
box -410 -1402 410 1402
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_0
timestamp 1713338890
transform 1 0 495 0 1 24298
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_1
timestamp 1713338890
transform 1 0 495 0 1 25910
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_2
timestamp 1713338890
transform 1 0 495 0 1 40310
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_3
timestamp 1713338890
transform 1 0 495 0 1 41898
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_4
timestamp 1713338890
transform 1 0 495 0 1 49894
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_5
timestamp 1713338890
transform 1 0 494 0 1 51493
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_6
timestamp 1713338890
transform 1 0 494 0 1 53096
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_7
timestamp 1713338890
transform 1 0 494 0 1 54702
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_8
timestamp 1713338890
transform 1 0 494 0 1 57899
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_9
timestamp 1713338890
transform 1 0 494 0 1 56306
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_10
timestamp 1713338890
transform 1 0 494 0 1 59516
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_11
timestamp 1713338890
transform 1 0 494 0 1 61108
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_12
timestamp 1713338890
transform 1 0 494 0 1 64300
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_13
timestamp 1713338890
transform 1 0 494 0 1 62694
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_14
timestamp 1713338890
transform 1 0 494 0 1 65891
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_15
timestamp 1713338890
transform 1 0 494 0 1 69043
box -410 -596 410 596
use M4_M3_CDNS_6903358316574  M4_M3_CDNS_6903358316574_16
timestamp 1713338890
transform 1 0 494 0 1 67498
box -410 -596 410 596
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_0
timestamp 1713338890
transform 1 0 494 0 1 15521
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_1
timestamp 1713338890
transform 1 0 494 0 1 18694
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_2
timestamp 1713338890
transform 1 0 494 0 1 21905
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_3
timestamp 1713338890
transform 1 0 494 0 1 28293
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_4
timestamp 1713338890
transform 1 0 494 0 1 31510
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_5
timestamp 1713338890
transform 1 0 494 0 1 34702
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_6
timestamp 1713338890
transform 1 0 494 0 1 37912
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_7
timestamp 1713338890
transform 1 0 494 0 1 44305
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316573  M5_M4_CDNS_6903358316573_8
timestamp 1713338890
transform 1 0 494 0 1 47501
box -416 -1408 416 1408
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_0
timestamp 1713338890
transform 1 0 495 0 1 24298
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_1
timestamp 1713338890
transform 1 0 495 0 1 25910
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_2
timestamp 1713338890
transform 1 0 495 0 1 40310
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_3
timestamp 1713338890
transform 1 0 495 0 1 41898
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_4
timestamp 1713338890
transform 1 0 495 0 1 49894
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_5
timestamp 1713338890
transform 1 0 494 0 1 51493
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_6
timestamp 1713338890
transform 1 0 494 0 1 53096
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_7
timestamp 1713338890
transform 1 0 494 0 1 54702
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_8
timestamp 1713338890
transform 1 0 494 0 1 57899
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_9
timestamp 1713338890
transform 1 0 494 0 1 56306
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_10
timestamp 1713338890
transform 1 0 494 0 1 61108
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_11
timestamp 1713338890
transform 1 0 494 0 1 59516
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_12
timestamp 1713338890
transform 1 0 494 0 1 64300
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_13
timestamp 1713338890
transform 1 0 494 0 1 62694
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_14
timestamp 1713338890
transform 1 0 494 0 1 65891
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_15
timestamp 1713338890
transform 1 0 494 0 1 67498
box -416 -602 416 602
use M5_M4_CDNS_6903358316575  M5_M4_CDNS_6903358316575_16
timestamp 1713338890
transform 1 0 494 0 1 69043
box -416 -602 416 602
<< labels >>
rlabel metal5 s 480 69049 480 69049 4 DVSS
port 1 nsew
rlabel metal5 s 480 15750 480 15750 4 DVSS
port 1 nsew
rlabel metal5 s 480 18921 480 18921 4 DVSS
port 1 nsew
rlabel metal5 s 480 21907 480 21907 4 DVSS
port 1 nsew
rlabel metal5 s 480 26100 480 26100 4 DVSS
port 1 nsew
rlabel metal5 s 480 40342 480 40342 4 DVSS
port 1 nsew
rlabel metal5 s 480 47595 480 47595 4 DVSS
port 1 nsew
rlabel metal5 s 480 57858 480 57858 4 DVSS
port 1 nsew
rlabel metal5 s 480 61058 480 61058 4 DVSS
port 1 nsew
rlabel metal5 s 480 66023 480 66023 4 DVSS
port 1 nsew
rlabel metal5 s 480 69049 480 69049 4 DVSS
port 1 nsew
rlabel metal4 s 480 69049 480 69049 4 DVSS
port 1 nsew
rlabel metal4 s 480 18921 480 18921 4 DVSS
port 1 nsew
rlabel metal4 s 480 15750 480 15750 4 DVSS
port 1 nsew
rlabel metal4 s 480 66023 480 66023 4 DVSS
port 1 nsew
rlabel metal4 s 480 57858 480 57858 4 DVSS
port 1 nsew
rlabel metal4 s 480 61058 480 61058 4 DVSS
port 1 nsew
rlabel metal4 s 480 47595 480 47595 4 DVSS
port 1 nsew
rlabel metal4 s 480 40342 480 40342 4 DVSS
port 1 nsew
rlabel metal4 s 480 69049 480 69049 4 DVSS
port 1 nsew
rlabel metal4 s 480 26100 480 26100 4 DVSS
port 1 nsew
rlabel metal4 s 480 21907 480 21907 4 DVSS
port 1 nsew
rlabel metal3 s 480 26100 480 26100 4 DVSS
port 1 nsew
rlabel metal3 s 480 69049 480 69049 4 DVSS
port 1 nsew
rlabel metal3 s 480 66023 480 66023 4 DVSS
port 1 nsew
rlabel metal3 s 480 61058 480 61058 4 DVSS
port 1 nsew
rlabel metal3 s 480 47595 480 47595 4 DVSS
port 1 nsew
rlabel metal3 s 480 15750 480 15750 4 DVSS
port 1 nsew
rlabel metal3 s 480 18921 480 18921 4 DVSS
port 1 nsew
rlabel metal3 s 480 21907 480 21907 4 DVSS
port 1 nsew
rlabel metal3 s 480 40342 480 40342 4 DVSS
port 1 nsew
rlabel metal3 s 480 57858 480 57858 4 DVSS
port 1 nsew
rlabel metal5 s 480 24284 480 24284 4 DVDD
port 2 nsew
rlabel metal5 s 480 28394 480 28394 4 DVDD
port 2 nsew
rlabel metal5 s 480 31609 480 31609 4 DVDD
port 2 nsew
rlabel metal5 s 480 34723 480 34723 4 DVDD
port 2 nsew
rlabel metal5 s 480 37959 480 37959 4 DVDD
port 2 nsew
rlabel metal5 s 480 41977 480 41977 4 DVDD
port 2 nsew
rlabel metal5 s 480 44368 480 44368 4 DVDD
port 2 nsew
rlabel metal5 s 480 53223 480 53223 4 DVDD
port 2 nsew
rlabel metal5 s 480 54658 480 54658 4 DVDD
port 2 nsew
rlabel metal5 s 480 56423 480 56423 4 DVDD
port 2 nsew
rlabel metal5 s 480 59623 480 59623 4 DVDD
port 2 nsew
rlabel metal5 s 480 67458 480 67458 4 DVDD
port 2 nsew
rlabel metal4 s 480 67458 480 67458 4 DVDD
port 2 nsew
rlabel metal4 s 480 59623 480 59623 4 DVDD
port 2 nsew
rlabel metal4 s 480 54658 480 54658 4 DVDD
port 2 nsew
rlabel metal4 s 480 53223 480 53223 4 DVDD
port 2 nsew
rlabel metal4 s 480 44368 480 44368 4 DVDD
port 2 nsew
rlabel metal4 s 480 41977 480 41977 4 DVDD
port 2 nsew
rlabel metal4 s 480 31609 480 31609 4 DVDD
port 2 nsew
rlabel metal4 s 480 37959 480 37959 4 DVDD
port 2 nsew
rlabel metal4 s 480 34723 480 34723 4 DVDD
port 2 nsew
rlabel metal4 s 480 28394 480 28394 4 DVDD
port 2 nsew
rlabel metal4 s 480 24284 480 24284 4 DVDD
port 2 nsew
rlabel metal4 s 480 56423 480 56423 4 DVDD
port 2 nsew
rlabel metal3 s 480 56423 480 56423 4 DVDD
port 2 nsew
rlabel metal3 s 480 24284 480 24284 4 DVDD
port 2 nsew
rlabel metal3 s 480 54658 480 54658 4 DVDD
port 2 nsew
rlabel metal3 s 480 53223 480 53223 4 DVDD
port 2 nsew
rlabel metal3 s 480 37959 480 37959 4 DVDD
port 2 nsew
rlabel metal3 s 480 28394 480 28394 4 DVDD
port 2 nsew
rlabel metal3 s 480 44368 480 44368 4 DVDD
port 2 nsew
rlabel metal3 s 480 67458 480 67458 4 DVDD
port 2 nsew
rlabel metal3 s 480 31609 480 31609 4 DVDD
port 2 nsew
rlabel metal3 s 480 34723 480 34723 4 DVDD
port 2 nsew
rlabel metal3 s 480 41977 480 41977 4 DVDD
port 2 nsew
rlabel metal3 s 480 59623 480 59623 4 DVDD
port 2 nsew
rlabel metal5 s 480 51458 480 51458 4 VDD
port 3 nsew
rlabel metal5 s 480 62823 480 62823 4 VDD
port 3 nsew
rlabel metal4 s 480 62823 480 62823 4 VDD
port 3 nsew
rlabel metal4 s 480 51458 480 51458 4 VDD
port 3 nsew
rlabel metal3 s 480 62823 480 62823 4 VDD
port 3 nsew
rlabel metal3 s 480 51458 480 51458 4 VDD
port 3 nsew
rlabel metal5 s 480 50023 480 50023 4 VSS
port 4 nsew
rlabel metal5 s 480 64258 480 64258 4 VSS
port 4 nsew
rlabel metal4 s 480 50023 480 50023 4 VSS
port 4 nsew
rlabel metal4 s 480 64258 480 64258 4 VSS
port 4 nsew
rlabel metal3 s 480 64258 480 64258 4 VSS
port 4 nsew
rlabel metal3 s 480 50023 480 50023 4 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1000 70000
<< end >>
