* NGSPICE file created from Balance_Inverter_flat.ext - technology: gf180mcuC

.subckt Balance_Inverter_flat VSS OUT OUT_B VIN VDD
X0 Inverter_0.OUT VIN.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X1 VDD OUT_B.t2 OUT.t1 VDD.t2 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2 OUT_B OUT.t2 VDD.t6 VDD.t5 pfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3 OUT_B VIN.t1 VSS.t3 VSS.t2 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X4 Inverter_0.OUT VIN.t2 VSS.t1 VSS.t0 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X5 VSS Inverter_0.OUT OUT.t0 VSS.t4 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
R0 VIN VIN.t1 48.6474
R1 VIN.n0 VIN.t2 19.0247
R2 VIN.n0 VIN.t0 17.3935
R3 VIN.n1 VIN.n0 4.12942
R4 VIN.n1 VIN 2.25699
R5 VIN.n2 VIN.n1 0.00437931
R6 VIN VIN.n2 0.00282759
R7 VDD.n1 VDD.t2 490.522
R8 VDD.n1 VDD.t5 485.783
R9 VDD VDD.t0 432.043
R10 VDD.n4 VDD.t6 9.56883
R11 VDD.n5 VDD.n0 9.47246
R12 VDD VDD.t1 6.4653
R13 VDD.n4 VDD.n3 3.1505
R14 VDD.n3 VDD.n1 3.1505
R15 VDD.n3 VDD.n2 1.4478
R16 VDD VDD.n5 0.510235
R17 VDD.n5 VDD 0.0857212
R18 VDD VDD.n4 0.0140398
R19 OUT_B OUT_B.t2 19.4226
R20 OUT_B.n3 OUT_B.n0 9.49418
R21 OUT_B.n2 OUT_B.n1 9.38848
R22 OUT_B OUT_B.n3 2.25319
R23 OUT_B.n3 OUT_B.n2 0.0122391
R24 OUT.n1 OUT.t2 49.5502
R25 OUT.n2 OUT.t0 9.49371
R26 OUT.n2 OUT.t1 9.3756
R27 OUT OUT.n2 3.6563
R28 OUT OUT.n1 2.25981
R29 OUT.n1 OUT.n0 0.00981034
R30 VSS.n6 VSS.t4 3956.52
R31 VSS.n5 VSS.t2 2285.81
R32 VSS.t4 VSS.n5 2169.44
R33 VSS VSS.n6 1909.39
R34 VSS.n6 VSS.t0 16.314
R35 VSS.n3 VSS.t3 9.48597
R36 VSS.n1 VSS.n0 9.32914
R37 VSS VSS.t1 9.03788
R38 VSS.n4 VSS.n3 2.6005
R39 VSS.n5 VSS.n4 2.6005
R40 VSS VSS.n1 0.451296
R41 VSS VSS.n1 0.139881
R42 VSS.n4 VSS.n2 0.0640538
R43 VSS.n3 VSS 0.00129646
C0 VDD VIN 0.268f
C1 OUT_B VIN 0.156f
C2 VIN Inverter_0.OUT 0.158f
C3 VDD OUT_B 0.313f
C4 VDD Inverter_0.OUT 0.14f
C5 OUT_B Inverter_0.OUT 0.00424f
C6 OUT VIN 0.087f
C7 OUT VDD 0.602f
C8 OUT OUT_B 0.268f
C9 OUT Inverter_0.OUT 0.219f
C10 OUT_B VSS 0.295f
C11 OUT VSS 0.556f
C12 Inverter_0.OUT VSS 0.565f
C13 VIN VSS 1.36f
C14 VDD VSS 1.98f
.ends

