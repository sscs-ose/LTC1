magic
tech gf180mcuC
magscale 1 10
timestamp 1695100097
<< nwell >>
rect -4444 -386 4444 386
<< nsubdiff >>
rect -4420 290 4420 362
rect -4420 -290 -4348 290
rect 4348 -290 4420 290
rect -4420 -362 4420 -290
<< polysilicon >>
rect -4260 189 -3480 202
rect -4260 143 -4247 189
rect -3493 143 -3480 189
rect -4260 100 -3480 143
rect -4260 -143 -3480 -100
rect -4260 -189 -4247 -143
rect -3493 -189 -3480 -143
rect -4260 -202 -3480 -189
rect -3400 189 -2620 202
rect -3400 143 -3387 189
rect -2633 143 -2620 189
rect -3400 100 -2620 143
rect -3400 -143 -2620 -100
rect -3400 -189 -3387 -143
rect -2633 -189 -2620 -143
rect -3400 -202 -2620 -189
rect -2540 189 -1760 202
rect -2540 143 -2527 189
rect -1773 143 -1760 189
rect -2540 100 -1760 143
rect -2540 -143 -1760 -100
rect -2540 -189 -2527 -143
rect -1773 -189 -1760 -143
rect -2540 -202 -1760 -189
rect -1680 189 -900 202
rect -1680 143 -1667 189
rect -913 143 -900 189
rect -1680 100 -900 143
rect -1680 -143 -900 -100
rect -1680 -189 -1667 -143
rect -913 -189 -900 -143
rect -1680 -202 -900 -189
rect -820 189 -40 202
rect -820 143 -807 189
rect -53 143 -40 189
rect -820 100 -40 143
rect -820 -143 -40 -100
rect -820 -189 -807 -143
rect -53 -189 -40 -143
rect -820 -202 -40 -189
rect 40 189 820 202
rect 40 143 53 189
rect 807 143 820 189
rect 40 100 820 143
rect 40 -143 820 -100
rect 40 -189 53 -143
rect 807 -189 820 -143
rect 40 -202 820 -189
rect 900 189 1680 202
rect 900 143 913 189
rect 1667 143 1680 189
rect 900 100 1680 143
rect 900 -143 1680 -100
rect 900 -189 913 -143
rect 1667 -189 1680 -143
rect 900 -202 1680 -189
rect 1760 189 2540 202
rect 1760 143 1773 189
rect 2527 143 2540 189
rect 1760 100 2540 143
rect 1760 -143 2540 -100
rect 1760 -189 1773 -143
rect 2527 -189 2540 -143
rect 1760 -202 2540 -189
rect 2620 189 3400 202
rect 2620 143 2633 189
rect 3387 143 3400 189
rect 2620 100 3400 143
rect 2620 -143 3400 -100
rect 2620 -189 2633 -143
rect 3387 -189 3400 -143
rect 2620 -202 3400 -189
rect 3480 189 4260 202
rect 3480 143 3493 189
rect 4247 143 4260 189
rect 3480 100 4260 143
rect 3480 -143 4260 -100
rect 3480 -189 3493 -143
rect 4247 -189 4260 -143
rect 3480 -202 4260 -189
<< polycontact >>
rect -4247 143 -3493 189
rect -4247 -189 -3493 -143
rect -3387 143 -2633 189
rect -3387 -189 -2633 -143
rect -2527 143 -1773 189
rect -2527 -189 -1773 -143
rect -1667 143 -913 189
rect -1667 -189 -913 -143
rect -807 143 -53 189
rect -807 -189 -53 -143
rect 53 143 807 189
rect 53 -189 807 -143
rect 913 143 1667 189
rect 913 -189 1667 -143
rect 1773 143 2527 189
rect 1773 -189 2527 -143
rect 2633 143 3387 189
rect 2633 -189 3387 -143
rect 3493 143 4247 189
rect 3493 -189 4247 -143
<< ppolyres >>
rect -4260 -100 -3480 100
rect -3400 -100 -2620 100
rect -2540 -100 -1760 100
rect -1680 -100 -900 100
rect -820 -100 -40 100
rect 40 -100 820 100
rect 900 -100 1680 100
rect 1760 -100 2540 100
rect 2620 -100 3400 100
rect 3480 -100 4260 100
<< metal1 >>
rect -4258 143 -4247 189
rect -3493 143 -3482 189
rect -3398 143 -3387 189
rect -2633 143 -2622 189
rect -2538 143 -2527 189
rect -1773 143 -1762 189
rect -1678 143 -1667 189
rect -913 143 -902 189
rect -818 143 -807 189
rect -53 143 -42 189
rect 42 143 53 189
rect 807 143 818 189
rect 902 143 913 189
rect 1667 143 1678 189
rect 1762 143 1773 189
rect 2527 143 2538 189
rect 2622 143 2633 189
rect 3387 143 3398 189
rect 3482 143 3493 189
rect 4247 143 4258 189
rect -4258 -189 -4247 -143
rect -3493 -189 -3482 -143
rect -3398 -189 -3387 -143
rect -2633 -189 -2622 -143
rect -2538 -189 -2527 -143
rect -1773 -189 -1762 -143
rect -1678 -189 -1667 -143
rect -913 -189 -902 -143
rect -818 -189 -807 -143
rect -53 -189 -42 -143
rect 42 -189 53 -143
rect 807 -189 818 -143
rect 902 -189 913 -143
rect 1667 -189 1678 -143
rect 1762 -189 1773 -143
rect 2527 -189 2538 -143
rect 2622 -189 2633 -143
rect 3387 -189 3398 -143
rect 3482 -189 3493 -143
rect 4247 -189 4258 -143
<< properties >>
string FIXED_BBOX -4384 -326 4384 326
string gencell ppolyf_u
string library gf180mcu
string parameters w 3.9 l 1.0 m 1 nx 10 wmin 0.80 lmin 1.00 rho 315 val 82.245 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
