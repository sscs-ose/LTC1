magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2913 -2045 2913 2045
<< psubdiff >>
rect -913 23 913 45
rect -913 -23 -891 23
rect -845 -23 -767 23
rect -721 -23 -643 23
rect -597 -23 -519 23
rect -473 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 597 23
rect 643 -23 721 23
rect 767 -23 845 23
rect 891 -23 913 23
rect -913 -45 913 -23
<< psubdiffcont >>
rect -891 -23 -845 23
rect -767 -23 -721 23
rect -643 -23 -597 23
rect -519 -23 -473 23
rect -395 -23 -349 23
rect -271 -23 -225 23
rect -147 -23 -101 23
rect -23 -23 23 23
rect 101 -23 147 23
rect 225 -23 271 23
rect 349 -23 395 23
rect 473 -23 519 23
rect 597 -23 643 23
rect 721 -23 767 23
rect 845 -23 891 23
<< metal1 >>
rect -902 23 902 34
rect -902 -23 -891 23
rect -845 -23 -767 23
rect -721 -23 -643 23
rect -597 -23 -519 23
rect -473 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 597 23
rect 643 -23 721 23
rect 767 -23 845 23
rect 891 -23 902 23
rect -902 -34 902 -23
<< end >>
