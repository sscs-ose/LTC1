magic
tech gf180mcuC
magscale 1 10
timestamp 1693552597
<< error_p >>
rect -874 -23 -863 23
rect -706 -23 -695 23
rect -538 -23 -527 23
rect -370 -23 -359 23
rect -202 -23 -191 23
rect -34 -23 -23 23
rect 134 -23 145 23
rect 302 -23 313 23
rect 470 -23 481 23
rect 638 -23 649 23
rect 806 -23 817 23
<< pwell >>
rect -900 -97 900 97
<< nmos >>
rect -784 -22 -728 22
rect -616 -22 -560 22
rect -448 -22 -392 22
rect -280 -22 -224 22
rect -112 -22 -56 22
rect 56 -22 112 22
rect 224 -22 280 22
rect 392 -22 448 22
rect 560 -22 616 22
rect 728 -22 784 22
<< ndiff >>
rect -876 23 -804 36
rect -876 -23 -863 23
rect -817 22 -804 23
rect -708 23 -636 36
rect -708 22 -695 23
rect -817 -22 -784 22
rect -728 -22 -695 22
rect -817 -23 -804 -22
rect -876 -36 -804 -23
rect -708 -23 -695 -22
rect -649 22 -636 23
rect -540 23 -468 36
rect -540 22 -527 23
rect -649 -22 -616 22
rect -560 -22 -527 22
rect -649 -23 -636 -22
rect -708 -36 -636 -23
rect -540 -23 -527 -22
rect -481 22 -468 23
rect -372 23 -300 36
rect -372 22 -359 23
rect -481 -22 -448 22
rect -392 -22 -359 22
rect -481 -23 -468 -22
rect -540 -36 -468 -23
rect -372 -23 -359 -22
rect -313 22 -300 23
rect -204 23 -132 36
rect -204 22 -191 23
rect -313 -22 -280 22
rect -224 -22 -191 22
rect -313 -23 -300 -22
rect -372 -36 -300 -23
rect -204 -23 -191 -22
rect -145 22 -132 23
rect -36 23 36 36
rect -36 22 -23 23
rect -145 -22 -112 22
rect -56 -22 -23 22
rect -145 -23 -132 -22
rect -204 -36 -132 -23
rect -36 -23 -23 -22
rect 23 22 36 23
rect 132 23 204 36
rect 132 22 145 23
rect 23 -22 56 22
rect 112 -22 145 22
rect 23 -23 36 -22
rect -36 -36 36 -23
rect 132 -23 145 -22
rect 191 22 204 23
rect 300 23 372 36
rect 300 22 313 23
rect 191 -22 224 22
rect 280 -22 313 22
rect 191 -23 204 -22
rect 132 -36 204 -23
rect 300 -23 313 -22
rect 359 22 372 23
rect 468 23 540 36
rect 468 22 481 23
rect 359 -22 392 22
rect 448 -22 481 22
rect 359 -23 372 -22
rect 300 -36 372 -23
rect 468 -23 481 -22
rect 527 22 540 23
rect 636 23 708 36
rect 636 22 649 23
rect 527 -22 560 22
rect 616 -22 649 22
rect 527 -23 540 -22
rect 468 -36 540 -23
rect 636 -23 649 -22
rect 695 22 708 23
rect 804 23 876 36
rect 804 22 817 23
rect 695 -22 728 22
rect 784 -22 817 22
rect 695 -23 708 -22
rect 636 -36 708 -23
rect 804 -23 817 -22
rect 863 -23 876 23
rect 804 -36 876 -23
<< ndiffc >>
rect -863 -23 -817 23
rect -695 -23 -649 23
rect -527 -23 -481 23
rect -359 -23 -313 23
rect -191 -23 -145 23
rect -23 -23 23 23
rect 145 -23 191 23
rect 313 -23 359 23
rect 481 -23 527 23
rect 649 -23 695 23
rect 817 -23 863 23
<< polysilicon >>
rect -784 22 -728 66
rect -784 -66 -728 -22
rect -616 22 -560 66
rect -616 -66 -560 -22
rect -448 22 -392 66
rect -448 -66 -392 -22
rect -280 22 -224 66
rect -280 -66 -224 -22
rect -112 22 -56 66
rect -112 -66 -56 -22
rect 56 22 112 66
rect 56 -66 112 -22
rect 224 22 280 66
rect 224 -66 280 -22
rect 392 22 448 66
rect 392 -66 448 -22
rect 560 22 616 66
rect 560 -66 616 -22
rect 728 22 784 66
rect 728 -66 784 -22
<< metal1 >>
rect -874 -23 -863 23
rect -817 -23 -806 23
rect -706 -23 -695 23
rect -649 -23 -638 23
rect -538 -23 -527 23
rect -481 -23 -470 23
rect -370 -23 -359 23
rect -313 -23 -302 23
rect -202 -23 -191 23
rect -145 -23 -134 23
rect -34 -23 -23 23
rect 23 -23 34 23
rect 134 -23 145 23
rect 191 -23 202 23
rect 302 -23 313 23
rect 359 -23 370 23
rect 470 -23 481 23
rect 527 -23 538 23
rect 638 -23 649 23
rect 695 -23 706 23
rect 806 -23 817 23
rect 863 -23 874 23
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.22 l 0.280 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
