* NGSPICE file created from pga_res_magice_parallel.ext - technology: gf180mcuC

.subckt ppolyf_u_VRC5QE a_2280_n202# a_4240_100# a_1720_n202# a_2560_100# a_n2200_n202#
+ a_n1640_n202# a_n4160_100# a_3120_n202# a_n2480_100# a_2560_n202# a_n3040_n202#
+ a_880_100# a_n2480_n202# a_n1920_n202# a_n2200_100# a_600_100# a_3680_100# w_n4904_n386#
+ a_3400_n202# a_2840_n202# a_n3320_n202# a_n520_100# a_n2760_n202# a_3400_100# a_1720_100#
+ a_4240_n202# a_3680_n202# a_n4160_n202# a_n3320_100# a_n1640_100# a_n3600_n202#
+ a_40_n202# a_4520_100# a_4520_n202# a_2840_100# a_3960_n202# a_320_n202# a_n4440_n202#
+ a_n3880_n202# a_n4440_100# a_1160_100# a_40_100# a_n2760_100# a_600_n202# a_n1080_100#
+ a_n4720_n202# a_3960_100# a_n800_100# a_880_n202# a_2280_100# a_n240_n202# a_n3880_100#
+ a_2000_100# a_n3600_100# a_n1920_100# a_n520_n202# a_1160_n202# a_320_100# a_n1080_n202#
+ a_n240_100# a_3120_100# a_n4720_100# a_1440_100# a_n800_n202# a_2000_n202# a_1440_n202#
+ a_n1360_n202# a_n3040_100# a_n1360_100#
X0 a_600_100# a_600_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X1 a_2280_100# a_2280_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X2 a_n800_100# a_n800_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X3 a_1160_100# a_1160_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X4 a_n4160_100# a_n4160_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X5 a_n240_100# a_n240_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X6 a_n3600_100# a_n3600_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X7 a_40_100# a_40_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X8 a_n3040_100# a_n3040_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X9 a_4520_100# a_4520_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X10 a_n2480_100# a_n2480_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X11 a_3960_100# a_3960_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X12 a_n1360_100# a_n1360_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X13 a_3400_100# a_3400_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X14 a_2840_100# a_2840_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X15 a_1720_100# a_1720_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X16 a_n4720_100# a_n4720_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X17 a_880_100# a_880_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X18 a_320_100# a_320_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X19 a_n1920_100# a_n1920_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X20 a_4240_100# a_4240_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X21 a_n2200_100# a_n2200_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X22 a_3680_100# a_3680_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X23 a_3120_100# a_3120_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X24 a_n1080_100# a_n1080_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X25 a_2560_100# a_2560_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X26 a_2000_100# a_2000_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X27 a_1440_100# a_1440_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X28 a_n4440_100# a_n4440_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X29 a_n520_100# a_n520_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X30 a_n3880_100# a_n3880_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X31 a_n3320_100# a_n3320_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X32 a_n2760_100# a_n2760_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X33 a_n1640_100# a_n1640_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
.ends

.subckt pag_res_magic A B G E C H F D VDD
Xppolyf_u_VRC5QE_0 m1_7017_3724# F m1_5335_5023# m1_7297_4056# m1_2973_3724# m1_6642_3724#
+ m1_577_3724# m1_8322_3724# m1_2680_4056# m1_7575_3720# C m1_5335_4371# m1_2973_3724#
+ m1_3095_3720# m1_2973_4056# m1_6642_4376# m1_8882_4056# VDD H D m1_3842_3724# m1_3095_5024#
+ m1_855_5023# m1_8415_4029# m1_6737_4056# m1_8977_3724# F m1_577_3724# m1_1695_4029#
+ m1_3512_4056# G m1_5057_3724# VDD VDD m1_7992_4056# m1_8977_3724# m1_5057_3724#
+ m1_577_3724# G E m1_6175_4029# m1_5242_4056# m1_2680_4056# m1_5802_3724# m1_3935_4029#
+ VDD m1_7575_5024# m1_4402_4056# m1_6082_3724# m1_7297_4056# m1_4497_3724# m1_2162_4376#
+ m1_6737_4056# G m1_2973_4056# m1_4497_3724# m1_8322_3724# m1_5335_4029# m1_6082_3724#
+ m1_5242_4056# m1_7575_4371# VDD m1_6642_4056# m1_5802_3724# m1_7017_3724# m1_6642_3724#
+ m1_3842_3724# m1_2162_4056# m1_3095_4371# ppolyf_u_VRC5QE
Xppolyf_u_VRC5QE_1 m1_7017_5028# m1_8966_5360# m1_5335_4029# m1_7297_5360# m1_2537_5028#
+ m1_3512_4920# E m1_7575_4677# m1_2257_5360# m1_7575_5024# m1_2162_5028# m1_6036_5360#
+ m1_2537_5028# m1_3095_5024# m1_2817_5360# m1_8882_5360# m1_8882_5360# VDD m1_9442_4708#
+ m1_7992_4920# m1_1695_5024# m1_4486_5360# m1_577_3724# m1_8602_5360# m1_6737_5360#
+ D m1_8882_5028# m1_855_5023# G m1_3562_5360# m1_714_4708# m1_5242_5028# VDD VDD
+ m1_8042_5360# m1_7575_3720# m1_5335_5023# E m1_2162_4708# E a_5435_4665# m1_5057_5360#
+ m1_2257_5360# m1_6642_4708# m1_4122_5360# VDD m1_8966_5360# m1_4402_5360# m1_5194_4708#
+ m1_7297_5360# m1_5242_5028# m1_4402_5360# m1_6737_5360# m1_4122_5360# m1_2817_5360#
+ m1_3095_3720# m1_6175_5024# m1_5057_5360# m1_4962_4708# m1_4486_5360# m1_8135_5333#
+ VDD m1_8042_5360# m1_4402_5028# m1_7017_5028# m1_6642_5028# m1_3095_4677# m1_3562_5360#
+ m1_3655_5333# ppolyf_u_VRC5QE
Xppolyf_u_VRC5QE_2 m1_7017_4376# m1_9442_4708# m1_6175_4029# m1_7575_4677# m1_4122_5360#
+ m1_4402_4056# G m1_8137_4376# m1_4122_5360# m1_7575_4371# m1_2162_4376# m1_6082_4708#
+ m1_4122_5360# m1_3095_4371# m1_4122_5360# m1_6642_5028# m1_7992_4920# VDD m1_8137_4376#
+ m1_8882_4056# m1_1417_4376# m1_3655_5333# m1_1695_4029# B m1_6175_5024# B m1_7992_4056#
+ G m1_3842_4708# m1_4402_5028# m1_1417_4376# m1_5242_4376# VDD VDD m1_8882_5028#
+ m1_8415_4029# m1_5335_4371# A m1_2162_4056# m1_714_4708# m1_8322_4708# m1_5194_4708#
+ m1_1695_5024# m1_6642_4056# m1_6082_4708# VDD m1_8135_5333# m1_3512_4920# m1_5897_4376#
+ m1_8602_5360# m1_5242_4376# m1_2162_5028# m1_6036_5360# C m1_3095_4677# m1_3935_4029#
+ m1_5897_4376# a_5435_4665# m1_3657_4376# m1_4962_4708# m1_8322_4708# VDD m1_6642_4708#
+ m1_3512_4056# m1_7017_4376# m1_6642_4376# m1_3657_4376# m1_2162_4708# m1_3842_4708#
+ ppolyf_u_VRC5QE
.ends

.subckt pga_res_magice_parallel VDD A C E G B D F H
Xpag_res_magic_0 A B G E C H F D VDD pag_res_magic
Xpag_res_magic_1 A B G E C H F D VDD pag_res_magic
.ends

