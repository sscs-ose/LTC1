magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2417 -2045 2417 2045
<< psubdiff >>
rect -417 23 417 45
rect -417 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 417 23
rect -417 -45 417 -23
<< psubdiffcont >>
rect -395 -23 -349 23
rect -271 -23 -225 23
rect -147 -23 -101 23
rect -23 -23 23 23
rect 101 -23 147 23
rect 225 -23 271 23
rect 349 -23 395 23
<< metal1 >>
rect -406 23 406 34
rect -406 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 406 23
rect -406 -34 406 -23
<< end >>
