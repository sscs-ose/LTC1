magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6678 -2278 6678 2278
<< nwell >>
rect -4678 -278 4678 278
<< nsubdiff >>
rect -4595 173 4595 195
rect -4595 -173 -4573 173
rect 4573 -173 4595 173
rect -4595 -195 4595 -173
<< nsubdiffcont >>
rect -4573 -173 4573 173
<< metal1 >>
rect -4584 173 4584 184
rect -4584 -173 -4573 173
rect 4573 -173 4584 173
rect -4584 -184 4584 -173
<< end >>
