magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2083 -2803 4795 4911
<< isosubstrate >>
rect 1479 -83 2795 2911
<< nwell >>
rect -83 1213 1139 2911
rect 1479 1213 2795 2911
<< polysilicon >>
rect 354 914 494 1914
rect 598 914 738 1914
rect 1999 1213 2139 1314
rect 1783 1002 2139 1213
rect 1999 914 2139 1002
rect 2243 914 2383 1314
<< metal1 >>
rect 79 2749 165 2817
rect 264 1958 340 2787
rect 508 1794 584 2558
rect 752 1958 828 2787
rect 891 2749 977 2817
rect 1641 2749 1727 2817
rect 508 1718 828 1794
rect 752 1197 828 1718
rect 1909 1197 1985 2558
rect 2153 1358 2229 2787
rect 2547 2749 2633 2817
rect 752 1019 1804 1197
rect 1909 1019 2347 1197
rect 79 11 165 79
rect 264 11 340 870
rect 752 270 828 1019
rect 1909 270 1985 1019
rect 891 11 977 79
rect 1115 -81 1191 106
rect 1641 11 1727 79
rect 2153 39 2229 870
rect 2397 270 2473 2558
rect 2547 11 2633 79
rect 1115 -157 1671 -81
rect 386 -411 789 -231
rect 1595 -282 1671 -157
rect 895 -803 1953 -727
<< metal2 >>
rect 386 -411 462 1556
rect 630 1376 1191 1556
rect 895 -803 971 77
rect 1115 11 1191 1376
rect 1773 -803 1849 -409
use M1_NWELL_CDNS_40661953145218  M1_NWELL_CDNS_40661953145218_0
timestamp 1713338890
transform 1 0 528 0 1 2783
box -457 -128 457 128
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_0
timestamp 1713338890
transform 1 0 1011 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_1
timestamp 1713338890
transform 1 0 45 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_2
timestamp 1713338890
transform 1 0 1607 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_3
timestamp 1713338890
transform 1 0 2667 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145225  M1_NWELL_CDNS_40661953145225_0
timestamp 1713338890
transform 1 0 2137 0 1 2783
box -504 -128 504 128
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform -1 0 668 0 1 1467
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform -1 0 424 0 1 1467
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_2
timestamp 1713338890
transform 1 0 1825 0 1 1108
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_3
timestamp 1713338890
transform 1 0 2305 0 1 1108
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 1 0 45 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 1 0 2667 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165611  M1_PSUB_CDNS_69033583165611_0
timestamp 1713338890
transform 1 0 1011 0 -1 468
box -45 -468 45 468
use M1_PSUB_CDNS_69033583165611  M1_PSUB_CDNS_69033583165611_1
timestamp 1713338890
transform 1 0 1607 0 -1 468
box -45 -468 45 468
use M1_PSUB_CDNS_69033583165612  M1_PSUB_CDNS_69033583165612_0
timestamp 1713338890
transform 1 0 2137 0 -1 45
box -421 -45 421 45
use M1_PSUB_CDNS_69033583165613  M1_PSUB_CDNS_69033583165613_0
timestamp 1713338890
transform 1 0 528 0 -1 45
box -374 -45 374 45
use M2_M1_CDNS_6903358316579  M2_M1_CDNS_6903358316579_0
timestamp 1713338890
transform 1 0 933 0 1 -447
box -38 -38 38 38
use M2_M1_CDNS_6903358316579  M2_M1_CDNS_6903358316579_1
timestamp 1713338890
transform 1 0 1811 0 1 -447
box -38 -38 38 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_0
timestamp 1713338890
transform 1 0 955 0 1 49
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_1
timestamp 1713338890
transform 1 0 985 0 1 -765
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_2
timestamp 1713338890
transform 1 0 1863 0 1 -765
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_3
timestamp 1713338890
transform 0 -1 1153 1 0 101
box -90 -38 90 38
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_0
timestamp 1713338890
transform 1 0 424 0 1 -321
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_1
timestamp 1713338890
transform 1 0 424 0 1 1466
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_2
timestamp 1713338890
transform 1 0 668 0 1 1466
box -38 -90 38 90
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_0
timestamp 1713338890
transform -1 0 738 0 1 270
box -88 -44 228 644
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_1
timestamp 1713338890
transform -1 0 494 0 1 270
box -88 -44 228 644
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_2
timestamp 1713338890
transform 1 0 1999 0 1 270
box -88 -44 228 644
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_3
timestamp 1713338890
transform 1 0 2243 0 1 270
box -88 -44 228 644
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1713338890
transform 1 0 598 0 1 1958
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_1
timestamp 1713338890
transform 1 0 354 0 1 1958
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314513  pmos_6p0_CDNS_4066195314513_0
timestamp 1713338890
transform -1 0 2139 0 1 1358
box -208 -120 348 1320
use pmos_6p0_CDNS_4066195314513  pmos_6p0_CDNS_4066195314513_1
timestamp 1713338890
transform -1 0 2383 0 1 1358
box -208 -120 348 1320
use pn_6p0_CDNS_4066195314510  pn_6p0_CDNS_4066195314510_0
timestamp 1713338890
transform -1 0 981 0 -1 -399
box -216 -216 312 312
use pn_6p0_CDNS_4066195314510  pn_6p0_CDNS_4066195314510_1
timestamp 1713338890
transform -1 0 1859 0 -1 -399
box -216 -216 312 312
<< labels >>
rlabel metal1 s 2112 1100 2112 1100 4 EN
port 1 nsew
rlabel metal1 s 2290 45 2290 45 4 DVSS
port 2 nsew
rlabel metal1 s 2283 2788 2283 2788 4 DVDD
port 3 nsew
rlabel metal1 s 256 45 256 45 4 VSS
port 4 nsew
rlabel metal1 s 75 2788 75 2788 4 VDD
port 5 nsew
rlabel metal1 s 2435 1100 2435 1100 4 ENB
port 6 nsew
rlabel metal1 s 421 1468 421 1468 4 PDRV
port 7 nsew
rlabel metal1 s 667 1468 667 1468 4 OE
port 8 nsew
<< end >>
