magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1487 -1019 1487 1019
<< metal1 >>
rect -487 13 487 19
rect -487 -13 -481 13
rect 481 -13 487 13
rect -487 -19 487 -13
<< via1 >>
rect -481 -13 481 13
<< metal2 >>
rect -487 13 487 19
rect -487 -13 -481 13
rect 481 -13 487 13
rect -487 -19 487 -13
<< end >>
