magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1484 -1019 1484 1019
<< metal2 >>
rect -484 14 484 19
rect -484 -14 -479 14
rect -451 -14 -417 14
rect -389 -14 -355 14
rect -327 -14 -293 14
rect -265 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 265 14
rect 293 -14 327 14
rect 355 -14 389 14
rect 417 -14 451 14
rect 479 -14 484 14
rect -484 -19 484 -14
<< via2 >>
rect -479 -14 -451 14
rect -417 -14 -389 14
rect -355 -14 -327 14
rect -293 -14 -265 14
rect -231 -14 -203 14
rect -169 -14 -141 14
rect -107 -14 -79 14
rect -45 -14 -17 14
rect 17 -14 45 14
rect 79 -14 107 14
rect 141 -14 169 14
rect 203 -14 231 14
rect 265 -14 293 14
rect 327 -14 355 14
rect 389 -14 417 14
rect 451 -14 479 14
<< metal3 >>
rect -484 14 484 19
rect -484 -14 -479 14
rect -451 -14 -417 14
rect -389 -14 -355 14
rect -327 -14 -293 14
rect -265 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 265 14
rect 293 -14 327 14
rect 355 -14 389 14
rect 417 -14 451 14
rect 479 -14 484 14
rect -484 -19 484 -14
<< end >>
