magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1073 -7013 1073 7013
<< metal1 >>
rect -73 6007 73 6013
rect -73 5981 -67 6007
rect -41 5981 -13 6007
rect 13 5981 41 6007
rect 67 5981 73 6007
rect -73 5953 73 5981
rect -73 5927 -67 5953
rect -41 5927 -13 5953
rect 13 5927 41 5953
rect 67 5927 73 5953
rect -73 5899 73 5927
rect -73 5873 -67 5899
rect -41 5873 -13 5899
rect 13 5873 41 5899
rect 67 5873 73 5899
rect -73 5845 73 5873
rect -73 5819 -67 5845
rect -41 5819 -13 5845
rect 13 5819 41 5845
rect 67 5819 73 5845
rect -73 5791 73 5819
rect -73 5765 -67 5791
rect -41 5765 -13 5791
rect 13 5765 41 5791
rect 67 5765 73 5791
rect -73 5737 73 5765
rect -73 5711 -67 5737
rect -41 5711 -13 5737
rect 13 5711 41 5737
rect 67 5711 73 5737
rect -73 5683 73 5711
rect -73 5657 -67 5683
rect -41 5657 -13 5683
rect 13 5657 41 5683
rect 67 5657 73 5683
rect -73 5629 73 5657
rect -73 5603 -67 5629
rect -41 5603 -13 5629
rect 13 5603 41 5629
rect 67 5603 73 5629
rect -73 5575 73 5603
rect -73 5549 -67 5575
rect -41 5549 -13 5575
rect 13 5549 41 5575
rect 67 5549 73 5575
rect -73 5521 73 5549
rect -73 5495 -67 5521
rect -41 5495 -13 5521
rect 13 5495 41 5521
rect 67 5495 73 5521
rect -73 5467 73 5495
rect -73 5441 -67 5467
rect -41 5441 -13 5467
rect 13 5441 41 5467
rect 67 5441 73 5467
rect -73 5413 73 5441
rect -73 5387 -67 5413
rect -41 5387 -13 5413
rect 13 5387 41 5413
rect 67 5387 73 5413
rect -73 5359 73 5387
rect -73 5333 -67 5359
rect -41 5333 -13 5359
rect 13 5333 41 5359
rect 67 5333 73 5359
rect -73 5305 73 5333
rect -73 5279 -67 5305
rect -41 5279 -13 5305
rect 13 5279 41 5305
rect 67 5279 73 5305
rect -73 5251 73 5279
rect -73 5225 -67 5251
rect -41 5225 -13 5251
rect 13 5225 41 5251
rect 67 5225 73 5251
rect -73 5197 73 5225
rect -73 5171 -67 5197
rect -41 5171 -13 5197
rect 13 5171 41 5197
rect 67 5171 73 5197
rect -73 5143 73 5171
rect -73 5117 -67 5143
rect -41 5117 -13 5143
rect 13 5117 41 5143
rect 67 5117 73 5143
rect -73 5089 73 5117
rect -73 5063 -67 5089
rect -41 5063 -13 5089
rect 13 5063 41 5089
rect 67 5063 73 5089
rect -73 5035 73 5063
rect -73 5009 -67 5035
rect -41 5009 -13 5035
rect 13 5009 41 5035
rect 67 5009 73 5035
rect -73 4981 73 5009
rect -73 4955 -67 4981
rect -41 4955 -13 4981
rect 13 4955 41 4981
rect 67 4955 73 4981
rect -73 4927 73 4955
rect -73 4901 -67 4927
rect -41 4901 -13 4927
rect 13 4901 41 4927
rect 67 4901 73 4927
rect -73 4873 73 4901
rect -73 4847 -67 4873
rect -41 4847 -13 4873
rect 13 4847 41 4873
rect 67 4847 73 4873
rect -73 4819 73 4847
rect -73 4793 -67 4819
rect -41 4793 -13 4819
rect 13 4793 41 4819
rect 67 4793 73 4819
rect -73 4765 73 4793
rect -73 4739 -67 4765
rect -41 4739 -13 4765
rect 13 4739 41 4765
rect 67 4739 73 4765
rect -73 4711 73 4739
rect -73 4685 -67 4711
rect -41 4685 -13 4711
rect 13 4685 41 4711
rect 67 4685 73 4711
rect -73 4657 73 4685
rect -73 4631 -67 4657
rect -41 4631 -13 4657
rect 13 4631 41 4657
rect 67 4631 73 4657
rect -73 4603 73 4631
rect -73 4577 -67 4603
rect -41 4577 -13 4603
rect 13 4577 41 4603
rect 67 4577 73 4603
rect -73 4549 73 4577
rect -73 4523 -67 4549
rect -41 4523 -13 4549
rect 13 4523 41 4549
rect 67 4523 73 4549
rect -73 4495 73 4523
rect -73 4469 -67 4495
rect -41 4469 -13 4495
rect 13 4469 41 4495
rect 67 4469 73 4495
rect -73 4441 73 4469
rect -73 4415 -67 4441
rect -41 4415 -13 4441
rect 13 4415 41 4441
rect 67 4415 73 4441
rect -73 4387 73 4415
rect -73 4361 -67 4387
rect -41 4361 -13 4387
rect 13 4361 41 4387
rect 67 4361 73 4387
rect -73 4333 73 4361
rect -73 4307 -67 4333
rect -41 4307 -13 4333
rect 13 4307 41 4333
rect 67 4307 73 4333
rect -73 4279 73 4307
rect -73 4253 -67 4279
rect -41 4253 -13 4279
rect 13 4253 41 4279
rect 67 4253 73 4279
rect -73 4225 73 4253
rect -73 4199 -67 4225
rect -41 4199 -13 4225
rect 13 4199 41 4225
rect 67 4199 73 4225
rect -73 4171 73 4199
rect -73 4145 -67 4171
rect -41 4145 -13 4171
rect 13 4145 41 4171
rect 67 4145 73 4171
rect -73 4117 73 4145
rect -73 4091 -67 4117
rect -41 4091 -13 4117
rect 13 4091 41 4117
rect 67 4091 73 4117
rect -73 4063 73 4091
rect -73 4037 -67 4063
rect -41 4037 -13 4063
rect 13 4037 41 4063
rect 67 4037 73 4063
rect -73 4009 73 4037
rect -73 3983 -67 4009
rect -41 3983 -13 4009
rect 13 3983 41 4009
rect 67 3983 73 4009
rect -73 3955 73 3983
rect -73 3929 -67 3955
rect -41 3929 -13 3955
rect 13 3929 41 3955
rect 67 3929 73 3955
rect -73 3901 73 3929
rect -73 3875 -67 3901
rect -41 3875 -13 3901
rect 13 3875 41 3901
rect 67 3875 73 3901
rect -73 3847 73 3875
rect -73 3821 -67 3847
rect -41 3821 -13 3847
rect 13 3821 41 3847
rect 67 3821 73 3847
rect -73 3793 73 3821
rect -73 3767 -67 3793
rect -41 3767 -13 3793
rect 13 3767 41 3793
rect 67 3767 73 3793
rect -73 3739 73 3767
rect -73 3713 -67 3739
rect -41 3713 -13 3739
rect 13 3713 41 3739
rect 67 3713 73 3739
rect -73 3685 73 3713
rect -73 3659 -67 3685
rect -41 3659 -13 3685
rect 13 3659 41 3685
rect 67 3659 73 3685
rect -73 3631 73 3659
rect -73 3605 -67 3631
rect -41 3605 -13 3631
rect 13 3605 41 3631
rect 67 3605 73 3631
rect -73 3577 73 3605
rect -73 3551 -67 3577
rect -41 3551 -13 3577
rect 13 3551 41 3577
rect 67 3551 73 3577
rect -73 3523 73 3551
rect -73 3497 -67 3523
rect -41 3497 -13 3523
rect 13 3497 41 3523
rect 67 3497 73 3523
rect -73 3469 73 3497
rect -73 3443 -67 3469
rect -41 3443 -13 3469
rect 13 3443 41 3469
rect 67 3443 73 3469
rect -73 3415 73 3443
rect -73 3389 -67 3415
rect -41 3389 -13 3415
rect 13 3389 41 3415
rect 67 3389 73 3415
rect -73 3361 73 3389
rect -73 3335 -67 3361
rect -41 3335 -13 3361
rect 13 3335 41 3361
rect 67 3335 73 3361
rect -73 3307 73 3335
rect -73 3281 -67 3307
rect -41 3281 -13 3307
rect 13 3281 41 3307
rect 67 3281 73 3307
rect -73 3253 73 3281
rect -73 3227 -67 3253
rect -41 3227 -13 3253
rect 13 3227 41 3253
rect 67 3227 73 3253
rect -73 3199 73 3227
rect -73 3173 -67 3199
rect -41 3173 -13 3199
rect 13 3173 41 3199
rect 67 3173 73 3199
rect -73 3145 73 3173
rect -73 3119 -67 3145
rect -41 3119 -13 3145
rect 13 3119 41 3145
rect 67 3119 73 3145
rect -73 3091 73 3119
rect -73 3065 -67 3091
rect -41 3065 -13 3091
rect 13 3065 41 3091
rect 67 3065 73 3091
rect -73 3037 73 3065
rect -73 3011 -67 3037
rect -41 3011 -13 3037
rect 13 3011 41 3037
rect 67 3011 73 3037
rect -73 2983 73 3011
rect -73 2957 -67 2983
rect -41 2957 -13 2983
rect 13 2957 41 2983
rect 67 2957 73 2983
rect -73 2929 73 2957
rect -73 2903 -67 2929
rect -41 2903 -13 2929
rect 13 2903 41 2929
rect 67 2903 73 2929
rect -73 2875 73 2903
rect -73 2849 -67 2875
rect -41 2849 -13 2875
rect 13 2849 41 2875
rect 67 2849 73 2875
rect -73 2821 73 2849
rect -73 2795 -67 2821
rect -41 2795 -13 2821
rect 13 2795 41 2821
rect 67 2795 73 2821
rect -73 2767 73 2795
rect -73 2741 -67 2767
rect -41 2741 -13 2767
rect 13 2741 41 2767
rect 67 2741 73 2767
rect -73 2713 73 2741
rect -73 2687 -67 2713
rect -41 2687 -13 2713
rect 13 2687 41 2713
rect 67 2687 73 2713
rect -73 2659 73 2687
rect -73 2633 -67 2659
rect -41 2633 -13 2659
rect 13 2633 41 2659
rect 67 2633 73 2659
rect -73 2605 73 2633
rect -73 2579 -67 2605
rect -41 2579 -13 2605
rect 13 2579 41 2605
rect 67 2579 73 2605
rect -73 2551 73 2579
rect -73 2525 -67 2551
rect -41 2525 -13 2551
rect 13 2525 41 2551
rect 67 2525 73 2551
rect -73 2497 73 2525
rect -73 2471 -67 2497
rect -41 2471 -13 2497
rect 13 2471 41 2497
rect 67 2471 73 2497
rect -73 2443 73 2471
rect -73 2417 -67 2443
rect -41 2417 -13 2443
rect 13 2417 41 2443
rect 67 2417 73 2443
rect -73 2389 73 2417
rect -73 2363 -67 2389
rect -41 2363 -13 2389
rect 13 2363 41 2389
rect 67 2363 73 2389
rect -73 2335 73 2363
rect -73 2309 -67 2335
rect -41 2309 -13 2335
rect 13 2309 41 2335
rect 67 2309 73 2335
rect -73 2281 73 2309
rect -73 2255 -67 2281
rect -41 2255 -13 2281
rect 13 2255 41 2281
rect 67 2255 73 2281
rect -73 2227 73 2255
rect -73 2201 -67 2227
rect -41 2201 -13 2227
rect 13 2201 41 2227
rect 67 2201 73 2227
rect -73 2173 73 2201
rect -73 2147 -67 2173
rect -41 2147 -13 2173
rect 13 2147 41 2173
rect 67 2147 73 2173
rect -73 2119 73 2147
rect -73 2093 -67 2119
rect -41 2093 -13 2119
rect 13 2093 41 2119
rect 67 2093 73 2119
rect -73 2065 73 2093
rect -73 2039 -67 2065
rect -41 2039 -13 2065
rect 13 2039 41 2065
rect 67 2039 73 2065
rect -73 2011 73 2039
rect -73 1985 -67 2011
rect -41 1985 -13 2011
rect 13 1985 41 2011
rect 67 1985 73 2011
rect -73 1957 73 1985
rect -73 1931 -67 1957
rect -41 1931 -13 1957
rect 13 1931 41 1957
rect 67 1931 73 1957
rect -73 1903 73 1931
rect -73 1877 -67 1903
rect -41 1877 -13 1903
rect 13 1877 41 1903
rect 67 1877 73 1903
rect -73 1849 73 1877
rect -73 1823 -67 1849
rect -41 1823 -13 1849
rect 13 1823 41 1849
rect 67 1823 73 1849
rect -73 1795 73 1823
rect -73 1769 -67 1795
rect -41 1769 -13 1795
rect 13 1769 41 1795
rect 67 1769 73 1795
rect -73 1741 73 1769
rect -73 1715 -67 1741
rect -41 1715 -13 1741
rect 13 1715 41 1741
rect 67 1715 73 1741
rect -73 1687 73 1715
rect -73 1661 -67 1687
rect -41 1661 -13 1687
rect 13 1661 41 1687
rect 67 1661 73 1687
rect -73 1633 73 1661
rect -73 1607 -67 1633
rect -41 1607 -13 1633
rect 13 1607 41 1633
rect 67 1607 73 1633
rect -73 1579 73 1607
rect -73 1553 -67 1579
rect -41 1553 -13 1579
rect 13 1553 41 1579
rect 67 1553 73 1579
rect -73 1525 73 1553
rect -73 1499 -67 1525
rect -41 1499 -13 1525
rect 13 1499 41 1525
rect 67 1499 73 1525
rect -73 1471 73 1499
rect -73 1445 -67 1471
rect -41 1445 -13 1471
rect 13 1445 41 1471
rect 67 1445 73 1471
rect -73 1417 73 1445
rect -73 1391 -67 1417
rect -41 1391 -13 1417
rect 13 1391 41 1417
rect 67 1391 73 1417
rect -73 1363 73 1391
rect -73 1337 -67 1363
rect -41 1337 -13 1363
rect 13 1337 41 1363
rect 67 1337 73 1363
rect -73 1309 73 1337
rect -73 1283 -67 1309
rect -41 1283 -13 1309
rect 13 1283 41 1309
rect 67 1283 73 1309
rect -73 1255 73 1283
rect -73 1229 -67 1255
rect -41 1229 -13 1255
rect 13 1229 41 1255
rect 67 1229 73 1255
rect -73 1201 73 1229
rect -73 1175 -67 1201
rect -41 1175 -13 1201
rect 13 1175 41 1201
rect 67 1175 73 1201
rect -73 1147 73 1175
rect -73 1121 -67 1147
rect -41 1121 -13 1147
rect 13 1121 41 1147
rect 67 1121 73 1147
rect -73 1093 73 1121
rect -73 1067 -67 1093
rect -41 1067 -13 1093
rect 13 1067 41 1093
rect 67 1067 73 1093
rect -73 1039 73 1067
rect -73 1013 -67 1039
rect -41 1013 -13 1039
rect 13 1013 41 1039
rect 67 1013 73 1039
rect -73 985 73 1013
rect -73 959 -67 985
rect -41 959 -13 985
rect 13 959 41 985
rect 67 959 73 985
rect -73 931 73 959
rect -73 905 -67 931
rect -41 905 -13 931
rect 13 905 41 931
rect 67 905 73 931
rect -73 877 73 905
rect -73 851 -67 877
rect -41 851 -13 877
rect 13 851 41 877
rect 67 851 73 877
rect -73 823 73 851
rect -73 797 -67 823
rect -41 797 -13 823
rect 13 797 41 823
rect 67 797 73 823
rect -73 769 73 797
rect -73 743 -67 769
rect -41 743 -13 769
rect 13 743 41 769
rect 67 743 73 769
rect -73 715 73 743
rect -73 689 -67 715
rect -41 689 -13 715
rect 13 689 41 715
rect 67 689 73 715
rect -73 661 73 689
rect -73 635 -67 661
rect -41 635 -13 661
rect 13 635 41 661
rect 67 635 73 661
rect -73 607 73 635
rect -73 581 -67 607
rect -41 581 -13 607
rect 13 581 41 607
rect 67 581 73 607
rect -73 553 73 581
rect -73 527 -67 553
rect -41 527 -13 553
rect 13 527 41 553
rect 67 527 73 553
rect -73 499 73 527
rect -73 473 -67 499
rect -41 473 -13 499
rect 13 473 41 499
rect 67 473 73 499
rect -73 445 73 473
rect -73 419 -67 445
rect -41 419 -13 445
rect 13 419 41 445
rect 67 419 73 445
rect -73 391 73 419
rect -73 365 -67 391
rect -41 365 -13 391
rect 13 365 41 391
rect 67 365 73 391
rect -73 337 73 365
rect -73 311 -67 337
rect -41 311 -13 337
rect 13 311 41 337
rect 67 311 73 337
rect -73 283 73 311
rect -73 257 -67 283
rect -41 257 -13 283
rect 13 257 41 283
rect 67 257 73 283
rect -73 229 73 257
rect -73 203 -67 229
rect -41 203 -13 229
rect 13 203 41 229
rect 67 203 73 229
rect -73 175 73 203
rect -73 149 -67 175
rect -41 149 -13 175
rect 13 149 41 175
rect 67 149 73 175
rect -73 121 73 149
rect -73 95 -67 121
rect -41 95 -13 121
rect 13 95 41 121
rect 67 95 73 121
rect -73 67 73 95
rect -73 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 73 67
rect -73 13 73 41
rect -73 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 73 13
rect -73 -41 73 -13
rect -73 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 73 -41
rect -73 -95 73 -67
rect -73 -121 -67 -95
rect -41 -121 -13 -95
rect 13 -121 41 -95
rect 67 -121 73 -95
rect -73 -149 73 -121
rect -73 -175 -67 -149
rect -41 -175 -13 -149
rect 13 -175 41 -149
rect 67 -175 73 -149
rect -73 -203 73 -175
rect -73 -229 -67 -203
rect -41 -229 -13 -203
rect 13 -229 41 -203
rect 67 -229 73 -203
rect -73 -257 73 -229
rect -73 -283 -67 -257
rect -41 -283 -13 -257
rect 13 -283 41 -257
rect 67 -283 73 -257
rect -73 -311 73 -283
rect -73 -337 -67 -311
rect -41 -337 -13 -311
rect 13 -337 41 -311
rect 67 -337 73 -311
rect -73 -365 73 -337
rect -73 -391 -67 -365
rect -41 -391 -13 -365
rect 13 -391 41 -365
rect 67 -391 73 -365
rect -73 -419 73 -391
rect -73 -445 -67 -419
rect -41 -445 -13 -419
rect 13 -445 41 -419
rect 67 -445 73 -419
rect -73 -473 73 -445
rect -73 -499 -67 -473
rect -41 -499 -13 -473
rect 13 -499 41 -473
rect 67 -499 73 -473
rect -73 -527 73 -499
rect -73 -553 -67 -527
rect -41 -553 -13 -527
rect 13 -553 41 -527
rect 67 -553 73 -527
rect -73 -581 73 -553
rect -73 -607 -67 -581
rect -41 -607 -13 -581
rect 13 -607 41 -581
rect 67 -607 73 -581
rect -73 -635 73 -607
rect -73 -661 -67 -635
rect -41 -661 -13 -635
rect 13 -661 41 -635
rect 67 -661 73 -635
rect -73 -689 73 -661
rect -73 -715 -67 -689
rect -41 -715 -13 -689
rect 13 -715 41 -689
rect 67 -715 73 -689
rect -73 -743 73 -715
rect -73 -769 -67 -743
rect -41 -769 -13 -743
rect 13 -769 41 -743
rect 67 -769 73 -743
rect -73 -797 73 -769
rect -73 -823 -67 -797
rect -41 -823 -13 -797
rect 13 -823 41 -797
rect 67 -823 73 -797
rect -73 -851 73 -823
rect -73 -877 -67 -851
rect -41 -877 -13 -851
rect 13 -877 41 -851
rect 67 -877 73 -851
rect -73 -905 73 -877
rect -73 -931 -67 -905
rect -41 -931 -13 -905
rect 13 -931 41 -905
rect 67 -931 73 -905
rect -73 -959 73 -931
rect -73 -985 -67 -959
rect -41 -985 -13 -959
rect 13 -985 41 -959
rect 67 -985 73 -959
rect -73 -1013 73 -985
rect -73 -1039 -67 -1013
rect -41 -1039 -13 -1013
rect 13 -1039 41 -1013
rect 67 -1039 73 -1013
rect -73 -1067 73 -1039
rect -73 -1093 -67 -1067
rect -41 -1093 -13 -1067
rect 13 -1093 41 -1067
rect 67 -1093 73 -1067
rect -73 -1121 73 -1093
rect -73 -1147 -67 -1121
rect -41 -1147 -13 -1121
rect 13 -1147 41 -1121
rect 67 -1147 73 -1121
rect -73 -1175 73 -1147
rect -73 -1201 -67 -1175
rect -41 -1201 -13 -1175
rect 13 -1201 41 -1175
rect 67 -1201 73 -1175
rect -73 -1229 73 -1201
rect -73 -1255 -67 -1229
rect -41 -1255 -13 -1229
rect 13 -1255 41 -1229
rect 67 -1255 73 -1229
rect -73 -1283 73 -1255
rect -73 -1309 -67 -1283
rect -41 -1309 -13 -1283
rect 13 -1309 41 -1283
rect 67 -1309 73 -1283
rect -73 -1337 73 -1309
rect -73 -1363 -67 -1337
rect -41 -1363 -13 -1337
rect 13 -1363 41 -1337
rect 67 -1363 73 -1337
rect -73 -1391 73 -1363
rect -73 -1417 -67 -1391
rect -41 -1417 -13 -1391
rect 13 -1417 41 -1391
rect 67 -1417 73 -1391
rect -73 -1445 73 -1417
rect -73 -1471 -67 -1445
rect -41 -1471 -13 -1445
rect 13 -1471 41 -1445
rect 67 -1471 73 -1445
rect -73 -1499 73 -1471
rect -73 -1525 -67 -1499
rect -41 -1525 -13 -1499
rect 13 -1525 41 -1499
rect 67 -1525 73 -1499
rect -73 -1553 73 -1525
rect -73 -1579 -67 -1553
rect -41 -1579 -13 -1553
rect 13 -1579 41 -1553
rect 67 -1579 73 -1553
rect -73 -1607 73 -1579
rect -73 -1633 -67 -1607
rect -41 -1633 -13 -1607
rect 13 -1633 41 -1607
rect 67 -1633 73 -1607
rect -73 -1661 73 -1633
rect -73 -1687 -67 -1661
rect -41 -1687 -13 -1661
rect 13 -1687 41 -1661
rect 67 -1687 73 -1661
rect -73 -1715 73 -1687
rect -73 -1741 -67 -1715
rect -41 -1741 -13 -1715
rect 13 -1741 41 -1715
rect 67 -1741 73 -1715
rect -73 -1769 73 -1741
rect -73 -1795 -67 -1769
rect -41 -1795 -13 -1769
rect 13 -1795 41 -1769
rect 67 -1795 73 -1769
rect -73 -1823 73 -1795
rect -73 -1849 -67 -1823
rect -41 -1849 -13 -1823
rect 13 -1849 41 -1823
rect 67 -1849 73 -1823
rect -73 -1877 73 -1849
rect -73 -1903 -67 -1877
rect -41 -1903 -13 -1877
rect 13 -1903 41 -1877
rect 67 -1903 73 -1877
rect -73 -1931 73 -1903
rect -73 -1957 -67 -1931
rect -41 -1957 -13 -1931
rect 13 -1957 41 -1931
rect 67 -1957 73 -1931
rect -73 -1985 73 -1957
rect -73 -2011 -67 -1985
rect -41 -2011 -13 -1985
rect 13 -2011 41 -1985
rect 67 -2011 73 -1985
rect -73 -2039 73 -2011
rect -73 -2065 -67 -2039
rect -41 -2065 -13 -2039
rect 13 -2065 41 -2039
rect 67 -2065 73 -2039
rect -73 -2093 73 -2065
rect -73 -2119 -67 -2093
rect -41 -2119 -13 -2093
rect 13 -2119 41 -2093
rect 67 -2119 73 -2093
rect -73 -2147 73 -2119
rect -73 -2173 -67 -2147
rect -41 -2173 -13 -2147
rect 13 -2173 41 -2147
rect 67 -2173 73 -2147
rect -73 -2201 73 -2173
rect -73 -2227 -67 -2201
rect -41 -2227 -13 -2201
rect 13 -2227 41 -2201
rect 67 -2227 73 -2201
rect -73 -2255 73 -2227
rect -73 -2281 -67 -2255
rect -41 -2281 -13 -2255
rect 13 -2281 41 -2255
rect 67 -2281 73 -2255
rect -73 -2309 73 -2281
rect -73 -2335 -67 -2309
rect -41 -2335 -13 -2309
rect 13 -2335 41 -2309
rect 67 -2335 73 -2309
rect -73 -2363 73 -2335
rect -73 -2389 -67 -2363
rect -41 -2389 -13 -2363
rect 13 -2389 41 -2363
rect 67 -2389 73 -2363
rect -73 -2417 73 -2389
rect -73 -2443 -67 -2417
rect -41 -2443 -13 -2417
rect 13 -2443 41 -2417
rect 67 -2443 73 -2417
rect -73 -2471 73 -2443
rect -73 -2497 -67 -2471
rect -41 -2497 -13 -2471
rect 13 -2497 41 -2471
rect 67 -2497 73 -2471
rect -73 -2525 73 -2497
rect -73 -2551 -67 -2525
rect -41 -2551 -13 -2525
rect 13 -2551 41 -2525
rect 67 -2551 73 -2525
rect -73 -2579 73 -2551
rect -73 -2605 -67 -2579
rect -41 -2605 -13 -2579
rect 13 -2605 41 -2579
rect 67 -2605 73 -2579
rect -73 -2633 73 -2605
rect -73 -2659 -67 -2633
rect -41 -2659 -13 -2633
rect 13 -2659 41 -2633
rect 67 -2659 73 -2633
rect -73 -2687 73 -2659
rect -73 -2713 -67 -2687
rect -41 -2713 -13 -2687
rect 13 -2713 41 -2687
rect 67 -2713 73 -2687
rect -73 -2741 73 -2713
rect -73 -2767 -67 -2741
rect -41 -2767 -13 -2741
rect 13 -2767 41 -2741
rect 67 -2767 73 -2741
rect -73 -2795 73 -2767
rect -73 -2821 -67 -2795
rect -41 -2821 -13 -2795
rect 13 -2821 41 -2795
rect 67 -2821 73 -2795
rect -73 -2849 73 -2821
rect -73 -2875 -67 -2849
rect -41 -2875 -13 -2849
rect 13 -2875 41 -2849
rect 67 -2875 73 -2849
rect -73 -2903 73 -2875
rect -73 -2929 -67 -2903
rect -41 -2929 -13 -2903
rect 13 -2929 41 -2903
rect 67 -2929 73 -2903
rect -73 -2957 73 -2929
rect -73 -2983 -67 -2957
rect -41 -2983 -13 -2957
rect 13 -2983 41 -2957
rect 67 -2983 73 -2957
rect -73 -3011 73 -2983
rect -73 -3037 -67 -3011
rect -41 -3037 -13 -3011
rect 13 -3037 41 -3011
rect 67 -3037 73 -3011
rect -73 -3065 73 -3037
rect -73 -3091 -67 -3065
rect -41 -3091 -13 -3065
rect 13 -3091 41 -3065
rect 67 -3091 73 -3065
rect -73 -3119 73 -3091
rect -73 -3145 -67 -3119
rect -41 -3145 -13 -3119
rect 13 -3145 41 -3119
rect 67 -3145 73 -3119
rect -73 -3173 73 -3145
rect -73 -3199 -67 -3173
rect -41 -3199 -13 -3173
rect 13 -3199 41 -3173
rect 67 -3199 73 -3173
rect -73 -3227 73 -3199
rect -73 -3253 -67 -3227
rect -41 -3253 -13 -3227
rect 13 -3253 41 -3227
rect 67 -3253 73 -3227
rect -73 -3281 73 -3253
rect -73 -3307 -67 -3281
rect -41 -3307 -13 -3281
rect 13 -3307 41 -3281
rect 67 -3307 73 -3281
rect -73 -3335 73 -3307
rect -73 -3361 -67 -3335
rect -41 -3361 -13 -3335
rect 13 -3361 41 -3335
rect 67 -3361 73 -3335
rect -73 -3389 73 -3361
rect -73 -3415 -67 -3389
rect -41 -3415 -13 -3389
rect 13 -3415 41 -3389
rect 67 -3415 73 -3389
rect -73 -3443 73 -3415
rect -73 -3469 -67 -3443
rect -41 -3469 -13 -3443
rect 13 -3469 41 -3443
rect 67 -3469 73 -3443
rect -73 -3497 73 -3469
rect -73 -3523 -67 -3497
rect -41 -3523 -13 -3497
rect 13 -3523 41 -3497
rect 67 -3523 73 -3497
rect -73 -3551 73 -3523
rect -73 -3577 -67 -3551
rect -41 -3577 -13 -3551
rect 13 -3577 41 -3551
rect 67 -3577 73 -3551
rect -73 -3605 73 -3577
rect -73 -3631 -67 -3605
rect -41 -3631 -13 -3605
rect 13 -3631 41 -3605
rect 67 -3631 73 -3605
rect -73 -3659 73 -3631
rect -73 -3685 -67 -3659
rect -41 -3685 -13 -3659
rect 13 -3685 41 -3659
rect 67 -3685 73 -3659
rect -73 -3713 73 -3685
rect -73 -3739 -67 -3713
rect -41 -3739 -13 -3713
rect 13 -3739 41 -3713
rect 67 -3739 73 -3713
rect -73 -3767 73 -3739
rect -73 -3793 -67 -3767
rect -41 -3793 -13 -3767
rect 13 -3793 41 -3767
rect 67 -3793 73 -3767
rect -73 -3821 73 -3793
rect -73 -3847 -67 -3821
rect -41 -3847 -13 -3821
rect 13 -3847 41 -3821
rect 67 -3847 73 -3821
rect -73 -3875 73 -3847
rect -73 -3901 -67 -3875
rect -41 -3901 -13 -3875
rect 13 -3901 41 -3875
rect 67 -3901 73 -3875
rect -73 -3929 73 -3901
rect -73 -3955 -67 -3929
rect -41 -3955 -13 -3929
rect 13 -3955 41 -3929
rect 67 -3955 73 -3929
rect -73 -3983 73 -3955
rect -73 -4009 -67 -3983
rect -41 -4009 -13 -3983
rect 13 -4009 41 -3983
rect 67 -4009 73 -3983
rect -73 -4037 73 -4009
rect -73 -4063 -67 -4037
rect -41 -4063 -13 -4037
rect 13 -4063 41 -4037
rect 67 -4063 73 -4037
rect -73 -4091 73 -4063
rect -73 -4117 -67 -4091
rect -41 -4117 -13 -4091
rect 13 -4117 41 -4091
rect 67 -4117 73 -4091
rect -73 -4145 73 -4117
rect -73 -4171 -67 -4145
rect -41 -4171 -13 -4145
rect 13 -4171 41 -4145
rect 67 -4171 73 -4145
rect -73 -4199 73 -4171
rect -73 -4225 -67 -4199
rect -41 -4225 -13 -4199
rect 13 -4225 41 -4199
rect 67 -4225 73 -4199
rect -73 -4253 73 -4225
rect -73 -4279 -67 -4253
rect -41 -4279 -13 -4253
rect 13 -4279 41 -4253
rect 67 -4279 73 -4253
rect -73 -4307 73 -4279
rect -73 -4333 -67 -4307
rect -41 -4333 -13 -4307
rect 13 -4333 41 -4307
rect 67 -4333 73 -4307
rect -73 -4361 73 -4333
rect -73 -4387 -67 -4361
rect -41 -4387 -13 -4361
rect 13 -4387 41 -4361
rect 67 -4387 73 -4361
rect -73 -4415 73 -4387
rect -73 -4441 -67 -4415
rect -41 -4441 -13 -4415
rect 13 -4441 41 -4415
rect 67 -4441 73 -4415
rect -73 -4469 73 -4441
rect -73 -4495 -67 -4469
rect -41 -4495 -13 -4469
rect 13 -4495 41 -4469
rect 67 -4495 73 -4469
rect -73 -4523 73 -4495
rect -73 -4549 -67 -4523
rect -41 -4549 -13 -4523
rect 13 -4549 41 -4523
rect 67 -4549 73 -4523
rect -73 -4577 73 -4549
rect -73 -4603 -67 -4577
rect -41 -4603 -13 -4577
rect 13 -4603 41 -4577
rect 67 -4603 73 -4577
rect -73 -4631 73 -4603
rect -73 -4657 -67 -4631
rect -41 -4657 -13 -4631
rect 13 -4657 41 -4631
rect 67 -4657 73 -4631
rect -73 -4685 73 -4657
rect -73 -4711 -67 -4685
rect -41 -4711 -13 -4685
rect 13 -4711 41 -4685
rect 67 -4711 73 -4685
rect -73 -4739 73 -4711
rect -73 -4765 -67 -4739
rect -41 -4765 -13 -4739
rect 13 -4765 41 -4739
rect 67 -4765 73 -4739
rect -73 -4793 73 -4765
rect -73 -4819 -67 -4793
rect -41 -4819 -13 -4793
rect 13 -4819 41 -4793
rect 67 -4819 73 -4793
rect -73 -4847 73 -4819
rect -73 -4873 -67 -4847
rect -41 -4873 -13 -4847
rect 13 -4873 41 -4847
rect 67 -4873 73 -4847
rect -73 -4901 73 -4873
rect -73 -4927 -67 -4901
rect -41 -4927 -13 -4901
rect 13 -4927 41 -4901
rect 67 -4927 73 -4901
rect -73 -4955 73 -4927
rect -73 -4981 -67 -4955
rect -41 -4981 -13 -4955
rect 13 -4981 41 -4955
rect 67 -4981 73 -4955
rect -73 -5009 73 -4981
rect -73 -5035 -67 -5009
rect -41 -5035 -13 -5009
rect 13 -5035 41 -5009
rect 67 -5035 73 -5009
rect -73 -5063 73 -5035
rect -73 -5089 -67 -5063
rect -41 -5089 -13 -5063
rect 13 -5089 41 -5063
rect 67 -5089 73 -5063
rect -73 -5117 73 -5089
rect -73 -5143 -67 -5117
rect -41 -5143 -13 -5117
rect 13 -5143 41 -5117
rect 67 -5143 73 -5117
rect -73 -5171 73 -5143
rect -73 -5197 -67 -5171
rect -41 -5197 -13 -5171
rect 13 -5197 41 -5171
rect 67 -5197 73 -5171
rect -73 -5225 73 -5197
rect -73 -5251 -67 -5225
rect -41 -5251 -13 -5225
rect 13 -5251 41 -5225
rect 67 -5251 73 -5225
rect -73 -5279 73 -5251
rect -73 -5305 -67 -5279
rect -41 -5305 -13 -5279
rect 13 -5305 41 -5279
rect 67 -5305 73 -5279
rect -73 -5333 73 -5305
rect -73 -5359 -67 -5333
rect -41 -5359 -13 -5333
rect 13 -5359 41 -5333
rect 67 -5359 73 -5333
rect -73 -5387 73 -5359
rect -73 -5413 -67 -5387
rect -41 -5413 -13 -5387
rect 13 -5413 41 -5387
rect 67 -5413 73 -5387
rect -73 -5441 73 -5413
rect -73 -5467 -67 -5441
rect -41 -5467 -13 -5441
rect 13 -5467 41 -5441
rect 67 -5467 73 -5441
rect -73 -5495 73 -5467
rect -73 -5521 -67 -5495
rect -41 -5521 -13 -5495
rect 13 -5521 41 -5495
rect 67 -5521 73 -5495
rect -73 -5549 73 -5521
rect -73 -5575 -67 -5549
rect -41 -5575 -13 -5549
rect 13 -5575 41 -5549
rect 67 -5575 73 -5549
rect -73 -5603 73 -5575
rect -73 -5629 -67 -5603
rect -41 -5629 -13 -5603
rect 13 -5629 41 -5603
rect 67 -5629 73 -5603
rect -73 -5657 73 -5629
rect -73 -5683 -67 -5657
rect -41 -5683 -13 -5657
rect 13 -5683 41 -5657
rect 67 -5683 73 -5657
rect -73 -5711 73 -5683
rect -73 -5737 -67 -5711
rect -41 -5737 -13 -5711
rect 13 -5737 41 -5711
rect 67 -5737 73 -5711
rect -73 -5765 73 -5737
rect -73 -5791 -67 -5765
rect -41 -5791 -13 -5765
rect 13 -5791 41 -5765
rect 67 -5791 73 -5765
rect -73 -5819 73 -5791
rect -73 -5845 -67 -5819
rect -41 -5845 -13 -5819
rect 13 -5845 41 -5819
rect 67 -5845 73 -5819
rect -73 -5873 73 -5845
rect -73 -5899 -67 -5873
rect -41 -5899 -13 -5873
rect 13 -5899 41 -5873
rect 67 -5899 73 -5873
rect -73 -5927 73 -5899
rect -73 -5953 -67 -5927
rect -41 -5953 -13 -5927
rect 13 -5953 41 -5927
rect 67 -5953 73 -5927
rect -73 -5981 73 -5953
rect -73 -6007 -67 -5981
rect -41 -6007 -13 -5981
rect 13 -6007 41 -5981
rect 67 -6007 73 -5981
rect -73 -6013 73 -6007
<< via1 >>
rect -67 5981 -41 6007
rect -13 5981 13 6007
rect 41 5981 67 6007
rect -67 5927 -41 5953
rect -13 5927 13 5953
rect 41 5927 67 5953
rect -67 5873 -41 5899
rect -13 5873 13 5899
rect 41 5873 67 5899
rect -67 5819 -41 5845
rect -13 5819 13 5845
rect 41 5819 67 5845
rect -67 5765 -41 5791
rect -13 5765 13 5791
rect 41 5765 67 5791
rect -67 5711 -41 5737
rect -13 5711 13 5737
rect 41 5711 67 5737
rect -67 5657 -41 5683
rect -13 5657 13 5683
rect 41 5657 67 5683
rect -67 5603 -41 5629
rect -13 5603 13 5629
rect 41 5603 67 5629
rect -67 5549 -41 5575
rect -13 5549 13 5575
rect 41 5549 67 5575
rect -67 5495 -41 5521
rect -13 5495 13 5521
rect 41 5495 67 5521
rect -67 5441 -41 5467
rect -13 5441 13 5467
rect 41 5441 67 5467
rect -67 5387 -41 5413
rect -13 5387 13 5413
rect 41 5387 67 5413
rect -67 5333 -41 5359
rect -13 5333 13 5359
rect 41 5333 67 5359
rect -67 5279 -41 5305
rect -13 5279 13 5305
rect 41 5279 67 5305
rect -67 5225 -41 5251
rect -13 5225 13 5251
rect 41 5225 67 5251
rect -67 5171 -41 5197
rect -13 5171 13 5197
rect 41 5171 67 5197
rect -67 5117 -41 5143
rect -13 5117 13 5143
rect 41 5117 67 5143
rect -67 5063 -41 5089
rect -13 5063 13 5089
rect 41 5063 67 5089
rect -67 5009 -41 5035
rect -13 5009 13 5035
rect 41 5009 67 5035
rect -67 4955 -41 4981
rect -13 4955 13 4981
rect 41 4955 67 4981
rect -67 4901 -41 4927
rect -13 4901 13 4927
rect 41 4901 67 4927
rect -67 4847 -41 4873
rect -13 4847 13 4873
rect 41 4847 67 4873
rect -67 4793 -41 4819
rect -13 4793 13 4819
rect 41 4793 67 4819
rect -67 4739 -41 4765
rect -13 4739 13 4765
rect 41 4739 67 4765
rect -67 4685 -41 4711
rect -13 4685 13 4711
rect 41 4685 67 4711
rect -67 4631 -41 4657
rect -13 4631 13 4657
rect 41 4631 67 4657
rect -67 4577 -41 4603
rect -13 4577 13 4603
rect 41 4577 67 4603
rect -67 4523 -41 4549
rect -13 4523 13 4549
rect 41 4523 67 4549
rect -67 4469 -41 4495
rect -13 4469 13 4495
rect 41 4469 67 4495
rect -67 4415 -41 4441
rect -13 4415 13 4441
rect 41 4415 67 4441
rect -67 4361 -41 4387
rect -13 4361 13 4387
rect 41 4361 67 4387
rect -67 4307 -41 4333
rect -13 4307 13 4333
rect 41 4307 67 4333
rect -67 4253 -41 4279
rect -13 4253 13 4279
rect 41 4253 67 4279
rect -67 4199 -41 4225
rect -13 4199 13 4225
rect 41 4199 67 4225
rect -67 4145 -41 4171
rect -13 4145 13 4171
rect 41 4145 67 4171
rect -67 4091 -41 4117
rect -13 4091 13 4117
rect 41 4091 67 4117
rect -67 4037 -41 4063
rect -13 4037 13 4063
rect 41 4037 67 4063
rect -67 3983 -41 4009
rect -13 3983 13 4009
rect 41 3983 67 4009
rect -67 3929 -41 3955
rect -13 3929 13 3955
rect 41 3929 67 3955
rect -67 3875 -41 3901
rect -13 3875 13 3901
rect 41 3875 67 3901
rect -67 3821 -41 3847
rect -13 3821 13 3847
rect 41 3821 67 3847
rect -67 3767 -41 3793
rect -13 3767 13 3793
rect 41 3767 67 3793
rect -67 3713 -41 3739
rect -13 3713 13 3739
rect 41 3713 67 3739
rect -67 3659 -41 3685
rect -13 3659 13 3685
rect 41 3659 67 3685
rect -67 3605 -41 3631
rect -13 3605 13 3631
rect 41 3605 67 3631
rect -67 3551 -41 3577
rect -13 3551 13 3577
rect 41 3551 67 3577
rect -67 3497 -41 3523
rect -13 3497 13 3523
rect 41 3497 67 3523
rect -67 3443 -41 3469
rect -13 3443 13 3469
rect 41 3443 67 3469
rect -67 3389 -41 3415
rect -13 3389 13 3415
rect 41 3389 67 3415
rect -67 3335 -41 3361
rect -13 3335 13 3361
rect 41 3335 67 3361
rect -67 3281 -41 3307
rect -13 3281 13 3307
rect 41 3281 67 3307
rect -67 3227 -41 3253
rect -13 3227 13 3253
rect 41 3227 67 3253
rect -67 3173 -41 3199
rect -13 3173 13 3199
rect 41 3173 67 3199
rect -67 3119 -41 3145
rect -13 3119 13 3145
rect 41 3119 67 3145
rect -67 3065 -41 3091
rect -13 3065 13 3091
rect 41 3065 67 3091
rect -67 3011 -41 3037
rect -13 3011 13 3037
rect 41 3011 67 3037
rect -67 2957 -41 2983
rect -13 2957 13 2983
rect 41 2957 67 2983
rect -67 2903 -41 2929
rect -13 2903 13 2929
rect 41 2903 67 2929
rect -67 2849 -41 2875
rect -13 2849 13 2875
rect 41 2849 67 2875
rect -67 2795 -41 2821
rect -13 2795 13 2821
rect 41 2795 67 2821
rect -67 2741 -41 2767
rect -13 2741 13 2767
rect 41 2741 67 2767
rect -67 2687 -41 2713
rect -13 2687 13 2713
rect 41 2687 67 2713
rect -67 2633 -41 2659
rect -13 2633 13 2659
rect 41 2633 67 2659
rect -67 2579 -41 2605
rect -13 2579 13 2605
rect 41 2579 67 2605
rect -67 2525 -41 2551
rect -13 2525 13 2551
rect 41 2525 67 2551
rect -67 2471 -41 2497
rect -13 2471 13 2497
rect 41 2471 67 2497
rect -67 2417 -41 2443
rect -13 2417 13 2443
rect 41 2417 67 2443
rect -67 2363 -41 2389
rect -13 2363 13 2389
rect 41 2363 67 2389
rect -67 2309 -41 2335
rect -13 2309 13 2335
rect 41 2309 67 2335
rect -67 2255 -41 2281
rect -13 2255 13 2281
rect 41 2255 67 2281
rect -67 2201 -41 2227
rect -13 2201 13 2227
rect 41 2201 67 2227
rect -67 2147 -41 2173
rect -13 2147 13 2173
rect 41 2147 67 2173
rect -67 2093 -41 2119
rect -13 2093 13 2119
rect 41 2093 67 2119
rect -67 2039 -41 2065
rect -13 2039 13 2065
rect 41 2039 67 2065
rect -67 1985 -41 2011
rect -13 1985 13 2011
rect 41 1985 67 2011
rect -67 1931 -41 1957
rect -13 1931 13 1957
rect 41 1931 67 1957
rect -67 1877 -41 1903
rect -13 1877 13 1903
rect 41 1877 67 1903
rect -67 1823 -41 1849
rect -13 1823 13 1849
rect 41 1823 67 1849
rect -67 1769 -41 1795
rect -13 1769 13 1795
rect 41 1769 67 1795
rect -67 1715 -41 1741
rect -13 1715 13 1741
rect 41 1715 67 1741
rect -67 1661 -41 1687
rect -13 1661 13 1687
rect 41 1661 67 1687
rect -67 1607 -41 1633
rect -13 1607 13 1633
rect 41 1607 67 1633
rect -67 1553 -41 1579
rect -13 1553 13 1579
rect 41 1553 67 1579
rect -67 1499 -41 1525
rect -13 1499 13 1525
rect 41 1499 67 1525
rect -67 1445 -41 1471
rect -13 1445 13 1471
rect 41 1445 67 1471
rect -67 1391 -41 1417
rect -13 1391 13 1417
rect 41 1391 67 1417
rect -67 1337 -41 1363
rect -13 1337 13 1363
rect 41 1337 67 1363
rect -67 1283 -41 1309
rect -13 1283 13 1309
rect 41 1283 67 1309
rect -67 1229 -41 1255
rect -13 1229 13 1255
rect 41 1229 67 1255
rect -67 1175 -41 1201
rect -13 1175 13 1201
rect 41 1175 67 1201
rect -67 1121 -41 1147
rect -13 1121 13 1147
rect 41 1121 67 1147
rect -67 1067 -41 1093
rect -13 1067 13 1093
rect 41 1067 67 1093
rect -67 1013 -41 1039
rect -13 1013 13 1039
rect 41 1013 67 1039
rect -67 959 -41 985
rect -13 959 13 985
rect 41 959 67 985
rect -67 905 -41 931
rect -13 905 13 931
rect 41 905 67 931
rect -67 851 -41 877
rect -13 851 13 877
rect 41 851 67 877
rect -67 797 -41 823
rect -13 797 13 823
rect 41 797 67 823
rect -67 743 -41 769
rect -13 743 13 769
rect 41 743 67 769
rect -67 689 -41 715
rect -13 689 13 715
rect 41 689 67 715
rect -67 635 -41 661
rect -13 635 13 661
rect 41 635 67 661
rect -67 581 -41 607
rect -13 581 13 607
rect 41 581 67 607
rect -67 527 -41 553
rect -13 527 13 553
rect 41 527 67 553
rect -67 473 -41 499
rect -13 473 13 499
rect 41 473 67 499
rect -67 419 -41 445
rect -13 419 13 445
rect 41 419 67 445
rect -67 365 -41 391
rect -13 365 13 391
rect 41 365 67 391
rect -67 311 -41 337
rect -13 311 13 337
rect 41 311 67 337
rect -67 257 -41 283
rect -13 257 13 283
rect 41 257 67 283
rect -67 203 -41 229
rect -13 203 13 229
rect 41 203 67 229
rect -67 149 -41 175
rect -13 149 13 175
rect 41 149 67 175
rect -67 95 -41 121
rect -13 95 13 121
rect 41 95 67 121
rect -67 41 -41 67
rect -13 41 13 67
rect 41 41 67 67
rect -67 -13 -41 13
rect -13 -13 13 13
rect 41 -13 67 13
rect -67 -67 -41 -41
rect -13 -67 13 -41
rect 41 -67 67 -41
rect -67 -121 -41 -95
rect -13 -121 13 -95
rect 41 -121 67 -95
rect -67 -175 -41 -149
rect -13 -175 13 -149
rect 41 -175 67 -149
rect -67 -229 -41 -203
rect -13 -229 13 -203
rect 41 -229 67 -203
rect -67 -283 -41 -257
rect -13 -283 13 -257
rect 41 -283 67 -257
rect -67 -337 -41 -311
rect -13 -337 13 -311
rect 41 -337 67 -311
rect -67 -391 -41 -365
rect -13 -391 13 -365
rect 41 -391 67 -365
rect -67 -445 -41 -419
rect -13 -445 13 -419
rect 41 -445 67 -419
rect -67 -499 -41 -473
rect -13 -499 13 -473
rect 41 -499 67 -473
rect -67 -553 -41 -527
rect -13 -553 13 -527
rect 41 -553 67 -527
rect -67 -607 -41 -581
rect -13 -607 13 -581
rect 41 -607 67 -581
rect -67 -661 -41 -635
rect -13 -661 13 -635
rect 41 -661 67 -635
rect -67 -715 -41 -689
rect -13 -715 13 -689
rect 41 -715 67 -689
rect -67 -769 -41 -743
rect -13 -769 13 -743
rect 41 -769 67 -743
rect -67 -823 -41 -797
rect -13 -823 13 -797
rect 41 -823 67 -797
rect -67 -877 -41 -851
rect -13 -877 13 -851
rect 41 -877 67 -851
rect -67 -931 -41 -905
rect -13 -931 13 -905
rect 41 -931 67 -905
rect -67 -985 -41 -959
rect -13 -985 13 -959
rect 41 -985 67 -959
rect -67 -1039 -41 -1013
rect -13 -1039 13 -1013
rect 41 -1039 67 -1013
rect -67 -1093 -41 -1067
rect -13 -1093 13 -1067
rect 41 -1093 67 -1067
rect -67 -1147 -41 -1121
rect -13 -1147 13 -1121
rect 41 -1147 67 -1121
rect -67 -1201 -41 -1175
rect -13 -1201 13 -1175
rect 41 -1201 67 -1175
rect -67 -1255 -41 -1229
rect -13 -1255 13 -1229
rect 41 -1255 67 -1229
rect -67 -1309 -41 -1283
rect -13 -1309 13 -1283
rect 41 -1309 67 -1283
rect -67 -1363 -41 -1337
rect -13 -1363 13 -1337
rect 41 -1363 67 -1337
rect -67 -1417 -41 -1391
rect -13 -1417 13 -1391
rect 41 -1417 67 -1391
rect -67 -1471 -41 -1445
rect -13 -1471 13 -1445
rect 41 -1471 67 -1445
rect -67 -1525 -41 -1499
rect -13 -1525 13 -1499
rect 41 -1525 67 -1499
rect -67 -1579 -41 -1553
rect -13 -1579 13 -1553
rect 41 -1579 67 -1553
rect -67 -1633 -41 -1607
rect -13 -1633 13 -1607
rect 41 -1633 67 -1607
rect -67 -1687 -41 -1661
rect -13 -1687 13 -1661
rect 41 -1687 67 -1661
rect -67 -1741 -41 -1715
rect -13 -1741 13 -1715
rect 41 -1741 67 -1715
rect -67 -1795 -41 -1769
rect -13 -1795 13 -1769
rect 41 -1795 67 -1769
rect -67 -1849 -41 -1823
rect -13 -1849 13 -1823
rect 41 -1849 67 -1823
rect -67 -1903 -41 -1877
rect -13 -1903 13 -1877
rect 41 -1903 67 -1877
rect -67 -1957 -41 -1931
rect -13 -1957 13 -1931
rect 41 -1957 67 -1931
rect -67 -2011 -41 -1985
rect -13 -2011 13 -1985
rect 41 -2011 67 -1985
rect -67 -2065 -41 -2039
rect -13 -2065 13 -2039
rect 41 -2065 67 -2039
rect -67 -2119 -41 -2093
rect -13 -2119 13 -2093
rect 41 -2119 67 -2093
rect -67 -2173 -41 -2147
rect -13 -2173 13 -2147
rect 41 -2173 67 -2147
rect -67 -2227 -41 -2201
rect -13 -2227 13 -2201
rect 41 -2227 67 -2201
rect -67 -2281 -41 -2255
rect -13 -2281 13 -2255
rect 41 -2281 67 -2255
rect -67 -2335 -41 -2309
rect -13 -2335 13 -2309
rect 41 -2335 67 -2309
rect -67 -2389 -41 -2363
rect -13 -2389 13 -2363
rect 41 -2389 67 -2363
rect -67 -2443 -41 -2417
rect -13 -2443 13 -2417
rect 41 -2443 67 -2417
rect -67 -2497 -41 -2471
rect -13 -2497 13 -2471
rect 41 -2497 67 -2471
rect -67 -2551 -41 -2525
rect -13 -2551 13 -2525
rect 41 -2551 67 -2525
rect -67 -2605 -41 -2579
rect -13 -2605 13 -2579
rect 41 -2605 67 -2579
rect -67 -2659 -41 -2633
rect -13 -2659 13 -2633
rect 41 -2659 67 -2633
rect -67 -2713 -41 -2687
rect -13 -2713 13 -2687
rect 41 -2713 67 -2687
rect -67 -2767 -41 -2741
rect -13 -2767 13 -2741
rect 41 -2767 67 -2741
rect -67 -2821 -41 -2795
rect -13 -2821 13 -2795
rect 41 -2821 67 -2795
rect -67 -2875 -41 -2849
rect -13 -2875 13 -2849
rect 41 -2875 67 -2849
rect -67 -2929 -41 -2903
rect -13 -2929 13 -2903
rect 41 -2929 67 -2903
rect -67 -2983 -41 -2957
rect -13 -2983 13 -2957
rect 41 -2983 67 -2957
rect -67 -3037 -41 -3011
rect -13 -3037 13 -3011
rect 41 -3037 67 -3011
rect -67 -3091 -41 -3065
rect -13 -3091 13 -3065
rect 41 -3091 67 -3065
rect -67 -3145 -41 -3119
rect -13 -3145 13 -3119
rect 41 -3145 67 -3119
rect -67 -3199 -41 -3173
rect -13 -3199 13 -3173
rect 41 -3199 67 -3173
rect -67 -3253 -41 -3227
rect -13 -3253 13 -3227
rect 41 -3253 67 -3227
rect -67 -3307 -41 -3281
rect -13 -3307 13 -3281
rect 41 -3307 67 -3281
rect -67 -3361 -41 -3335
rect -13 -3361 13 -3335
rect 41 -3361 67 -3335
rect -67 -3415 -41 -3389
rect -13 -3415 13 -3389
rect 41 -3415 67 -3389
rect -67 -3469 -41 -3443
rect -13 -3469 13 -3443
rect 41 -3469 67 -3443
rect -67 -3523 -41 -3497
rect -13 -3523 13 -3497
rect 41 -3523 67 -3497
rect -67 -3577 -41 -3551
rect -13 -3577 13 -3551
rect 41 -3577 67 -3551
rect -67 -3631 -41 -3605
rect -13 -3631 13 -3605
rect 41 -3631 67 -3605
rect -67 -3685 -41 -3659
rect -13 -3685 13 -3659
rect 41 -3685 67 -3659
rect -67 -3739 -41 -3713
rect -13 -3739 13 -3713
rect 41 -3739 67 -3713
rect -67 -3793 -41 -3767
rect -13 -3793 13 -3767
rect 41 -3793 67 -3767
rect -67 -3847 -41 -3821
rect -13 -3847 13 -3821
rect 41 -3847 67 -3821
rect -67 -3901 -41 -3875
rect -13 -3901 13 -3875
rect 41 -3901 67 -3875
rect -67 -3955 -41 -3929
rect -13 -3955 13 -3929
rect 41 -3955 67 -3929
rect -67 -4009 -41 -3983
rect -13 -4009 13 -3983
rect 41 -4009 67 -3983
rect -67 -4063 -41 -4037
rect -13 -4063 13 -4037
rect 41 -4063 67 -4037
rect -67 -4117 -41 -4091
rect -13 -4117 13 -4091
rect 41 -4117 67 -4091
rect -67 -4171 -41 -4145
rect -13 -4171 13 -4145
rect 41 -4171 67 -4145
rect -67 -4225 -41 -4199
rect -13 -4225 13 -4199
rect 41 -4225 67 -4199
rect -67 -4279 -41 -4253
rect -13 -4279 13 -4253
rect 41 -4279 67 -4253
rect -67 -4333 -41 -4307
rect -13 -4333 13 -4307
rect 41 -4333 67 -4307
rect -67 -4387 -41 -4361
rect -13 -4387 13 -4361
rect 41 -4387 67 -4361
rect -67 -4441 -41 -4415
rect -13 -4441 13 -4415
rect 41 -4441 67 -4415
rect -67 -4495 -41 -4469
rect -13 -4495 13 -4469
rect 41 -4495 67 -4469
rect -67 -4549 -41 -4523
rect -13 -4549 13 -4523
rect 41 -4549 67 -4523
rect -67 -4603 -41 -4577
rect -13 -4603 13 -4577
rect 41 -4603 67 -4577
rect -67 -4657 -41 -4631
rect -13 -4657 13 -4631
rect 41 -4657 67 -4631
rect -67 -4711 -41 -4685
rect -13 -4711 13 -4685
rect 41 -4711 67 -4685
rect -67 -4765 -41 -4739
rect -13 -4765 13 -4739
rect 41 -4765 67 -4739
rect -67 -4819 -41 -4793
rect -13 -4819 13 -4793
rect 41 -4819 67 -4793
rect -67 -4873 -41 -4847
rect -13 -4873 13 -4847
rect 41 -4873 67 -4847
rect -67 -4927 -41 -4901
rect -13 -4927 13 -4901
rect 41 -4927 67 -4901
rect -67 -4981 -41 -4955
rect -13 -4981 13 -4955
rect 41 -4981 67 -4955
rect -67 -5035 -41 -5009
rect -13 -5035 13 -5009
rect 41 -5035 67 -5009
rect -67 -5089 -41 -5063
rect -13 -5089 13 -5063
rect 41 -5089 67 -5063
rect -67 -5143 -41 -5117
rect -13 -5143 13 -5117
rect 41 -5143 67 -5117
rect -67 -5197 -41 -5171
rect -13 -5197 13 -5171
rect 41 -5197 67 -5171
rect -67 -5251 -41 -5225
rect -13 -5251 13 -5225
rect 41 -5251 67 -5225
rect -67 -5305 -41 -5279
rect -13 -5305 13 -5279
rect 41 -5305 67 -5279
rect -67 -5359 -41 -5333
rect -13 -5359 13 -5333
rect 41 -5359 67 -5333
rect -67 -5413 -41 -5387
rect -13 -5413 13 -5387
rect 41 -5413 67 -5387
rect -67 -5467 -41 -5441
rect -13 -5467 13 -5441
rect 41 -5467 67 -5441
rect -67 -5521 -41 -5495
rect -13 -5521 13 -5495
rect 41 -5521 67 -5495
rect -67 -5575 -41 -5549
rect -13 -5575 13 -5549
rect 41 -5575 67 -5549
rect -67 -5629 -41 -5603
rect -13 -5629 13 -5603
rect 41 -5629 67 -5603
rect -67 -5683 -41 -5657
rect -13 -5683 13 -5657
rect 41 -5683 67 -5657
rect -67 -5737 -41 -5711
rect -13 -5737 13 -5711
rect 41 -5737 67 -5711
rect -67 -5791 -41 -5765
rect -13 -5791 13 -5765
rect 41 -5791 67 -5765
rect -67 -5845 -41 -5819
rect -13 -5845 13 -5819
rect 41 -5845 67 -5819
rect -67 -5899 -41 -5873
rect -13 -5899 13 -5873
rect 41 -5899 67 -5873
rect -67 -5953 -41 -5927
rect -13 -5953 13 -5927
rect 41 -5953 67 -5927
rect -67 -6007 -41 -5981
rect -13 -6007 13 -5981
rect 41 -6007 67 -5981
<< metal2 >>
rect -73 6007 73 6013
rect -73 5981 -67 6007
rect -41 5981 -13 6007
rect 13 5981 41 6007
rect 67 5981 73 6007
rect -73 5953 73 5981
rect -73 5927 -67 5953
rect -41 5927 -13 5953
rect 13 5927 41 5953
rect 67 5927 73 5953
rect -73 5899 73 5927
rect -73 5873 -67 5899
rect -41 5873 -13 5899
rect 13 5873 41 5899
rect 67 5873 73 5899
rect -73 5845 73 5873
rect -73 5819 -67 5845
rect -41 5819 -13 5845
rect 13 5819 41 5845
rect 67 5819 73 5845
rect -73 5791 73 5819
rect -73 5765 -67 5791
rect -41 5765 -13 5791
rect 13 5765 41 5791
rect 67 5765 73 5791
rect -73 5737 73 5765
rect -73 5711 -67 5737
rect -41 5711 -13 5737
rect 13 5711 41 5737
rect 67 5711 73 5737
rect -73 5683 73 5711
rect -73 5657 -67 5683
rect -41 5657 -13 5683
rect 13 5657 41 5683
rect 67 5657 73 5683
rect -73 5629 73 5657
rect -73 5603 -67 5629
rect -41 5603 -13 5629
rect 13 5603 41 5629
rect 67 5603 73 5629
rect -73 5575 73 5603
rect -73 5549 -67 5575
rect -41 5549 -13 5575
rect 13 5549 41 5575
rect 67 5549 73 5575
rect -73 5521 73 5549
rect -73 5495 -67 5521
rect -41 5495 -13 5521
rect 13 5495 41 5521
rect 67 5495 73 5521
rect -73 5467 73 5495
rect -73 5441 -67 5467
rect -41 5441 -13 5467
rect 13 5441 41 5467
rect 67 5441 73 5467
rect -73 5413 73 5441
rect -73 5387 -67 5413
rect -41 5387 -13 5413
rect 13 5387 41 5413
rect 67 5387 73 5413
rect -73 5359 73 5387
rect -73 5333 -67 5359
rect -41 5333 -13 5359
rect 13 5333 41 5359
rect 67 5333 73 5359
rect -73 5305 73 5333
rect -73 5279 -67 5305
rect -41 5279 -13 5305
rect 13 5279 41 5305
rect 67 5279 73 5305
rect -73 5251 73 5279
rect -73 5225 -67 5251
rect -41 5225 -13 5251
rect 13 5225 41 5251
rect 67 5225 73 5251
rect -73 5197 73 5225
rect -73 5171 -67 5197
rect -41 5171 -13 5197
rect 13 5171 41 5197
rect 67 5171 73 5197
rect -73 5143 73 5171
rect -73 5117 -67 5143
rect -41 5117 -13 5143
rect 13 5117 41 5143
rect 67 5117 73 5143
rect -73 5089 73 5117
rect -73 5063 -67 5089
rect -41 5063 -13 5089
rect 13 5063 41 5089
rect 67 5063 73 5089
rect -73 5035 73 5063
rect -73 5009 -67 5035
rect -41 5009 -13 5035
rect 13 5009 41 5035
rect 67 5009 73 5035
rect -73 4981 73 5009
rect -73 4955 -67 4981
rect -41 4955 -13 4981
rect 13 4955 41 4981
rect 67 4955 73 4981
rect -73 4927 73 4955
rect -73 4901 -67 4927
rect -41 4901 -13 4927
rect 13 4901 41 4927
rect 67 4901 73 4927
rect -73 4873 73 4901
rect -73 4847 -67 4873
rect -41 4847 -13 4873
rect 13 4847 41 4873
rect 67 4847 73 4873
rect -73 4819 73 4847
rect -73 4793 -67 4819
rect -41 4793 -13 4819
rect 13 4793 41 4819
rect 67 4793 73 4819
rect -73 4765 73 4793
rect -73 4739 -67 4765
rect -41 4739 -13 4765
rect 13 4739 41 4765
rect 67 4739 73 4765
rect -73 4711 73 4739
rect -73 4685 -67 4711
rect -41 4685 -13 4711
rect 13 4685 41 4711
rect 67 4685 73 4711
rect -73 4657 73 4685
rect -73 4631 -67 4657
rect -41 4631 -13 4657
rect 13 4631 41 4657
rect 67 4631 73 4657
rect -73 4603 73 4631
rect -73 4577 -67 4603
rect -41 4577 -13 4603
rect 13 4577 41 4603
rect 67 4577 73 4603
rect -73 4549 73 4577
rect -73 4523 -67 4549
rect -41 4523 -13 4549
rect 13 4523 41 4549
rect 67 4523 73 4549
rect -73 4495 73 4523
rect -73 4469 -67 4495
rect -41 4469 -13 4495
rect 13 4469 41 4495
rect 67 4469 73 4495
rect -73 4441 73 4469
rect -73 4415 -67 4441
rect -41 4415 -13 4441
rect 13 4415 41 4441
rect 67 4415 73 4441
rect -73 4387 73 4415
rect -73 4361 -67 4387
rect -41 4361 -13 4387
rect 13 4361 41 4387
rect 67 4361 73 4387
rect -73 4333 73 4361
rect -73 4307 -67 4333
rect -41 4307 -13 4333
rect 13 4307 41 4333
rect 67 4307 73 4333
rect -73 4279 73 4307
rect -73 4253 -67 4279
rect -41 4253 -13 4279
rect 13 4253 41 4279
rect 67 4253 73 4279
rect -73 4225 73 4253
rect -73 4199 -67 4225
rect -41 4199 -13 4225
rect 13 4199 41 4225
rect 67 4199 73 4225
rect -73 4171 73 4199
rect -73 4145 -67 4171
rect -41 4145 -13 4171
rect 13 4145 41 4171
rect 67 4145 73 4171
rect -73 4117 73 4145
rect -73 4091 -67 4117
rect -41 4091 -13 4117
rect 13 4091 41 4117
rect 67 4091 73 4117
rect -73 4063 73 4091
rect -73 4037 -67 4063
rect -41 4037 -13 4063
rect 13 4037 41 4063
rect 67 4037 73 4063
rect -73 4009 73 4037
rect -73 3983 -67 4009
rect -41 3983 -13 4009
rect 13 3983 41 4009
rect 67 3983 73 4009
rect -73 3955 73 3983
rect -73 3929 -67 3955
rect -41 3929 -13 3955
rect 13 3929 41 3955
rect 67 3929 73 3955
rect -73 3901 73 3929
rect -73 3875 -67 3901
rect -41 3875 -13 3901
rect 13 3875 41 3901
rect 67 3875 73 3901
rect -73 3847 73 3875
rect -73 3821 -67 3847
rect -41 3821 -13 3847
rect 13 3821 41 3847
rect 67 3821 73 3847
rect -73 3793 73 3821
rect -73 3767 -67 3793
rect -41 3767 -13 3793
rect 13 3767 41 3793
rect 67 3767 73 3793
rect -73 3739 73 3767
rect -73 3713 -67 3739
rect -41 3713 -13 3739
rect 13 3713 41 3739
rect 67 3713 73 3739
rect -73 3685 73 3713
rect -73 3659 -67 3685
rect -41 3659 -13 3685
rect 13 3659 41 3685
rect 67 3659 73 3685
rect -73 3631 73 3659
rect -73 3605 -67 3631
rect -41 3605 -13 3631
rect 13 3605 41 3631
rect 67 3605 73 3631
rect -73 3577 73 3605
rect -73 3551 -67 3577
rect -41 3551 -13 3577
rect 13 3551 41 3577
rect 67 3551 73 3577
rect -73 3523 73 3551
rect -73 3497 -67 3523
rect -41 3497 -13 3523
rect 13 3497 41 3523
rect 67 3497 73 3523
rect -73 3469 73 3497
rect -73 3443 -67 3469
rect -41 3443 -13 3469
rect 13 3443 41 3469
rect 67 3443 73 3469
rect -73 3415 73 3443
rect -73 3389 -67 3415
rect -41 3389 -13 3415
rect 13 3389 41 3415
rect 67 3389 73 3415
rect -73 3361 73 3389
rect -73 3335 -67 3361
rect -41 3335 -13 3361
rect 13 3335 41 3361
rect 67 3335 73 3361
rect -73 3307 73 3335
rect -73 3281 -67 3307
rect -41 3281 -13 3307
rect 13 3281 41 3307
rect 67 3281 73 3307
rect -73 3253 73 3281
rect -73 3227 -67 3253
rect -41 3227 -13 3253
rect 13 3227 41 3253
rect 67 3227 73 3253
rect -73 3199 73 3227
rect -73 3173 -67 3199
rect -41 3173 -13 3199
rect 13 3173 41 3199
rect 67 3173 73 3199
rect -73 3145 73 3173
rect -73 3119 -67 3145
rect -41 3119 -13 3145
rect 13 3119 41 3145
rect 67 3119 73 3145
rect -73 3091 73 3119
rect -73 3065 -67 3091
rect -41 3065 -13 3091
rect 13 3065 41 3091
rect 67 3065 73 3091
rect -73 3037 73 3065
rect -73 3011 -67 3037
rect -41 3011 -13 3037
rect 13 3011 41 3037
rect 67 3011 73 3037
rect -73 2983 73 3011
rect -73 2957 -67 2983
rect -41 2957 -13 2983
rect 13 2957 41 2983
rect 67 2957 73 2983
rect -73 2929 73 2957
rect -73 2903 -67 2929
rect -41 2903 -13 2929
rect 13 2903 41 2929
rect 67 2903 73 2929
rect -73 2875 73 2903
rect -73 2849 -67 2875
rect -41 2849 -13 2875
rect 13 2849 41 2875
rect 67 2849 73 2875
rect -73 2821 73 2849
rect -73 2795 -67 2821
rect -41 2795 -13 2821
rect 13 2795 41 2821
rect 67 2795 73 2821
rect -73 2767 73 2795
rect -73 2741 -67 2767
rect -41 2741 -13 2767
rect 13 2741 41 2767
rect 67 2741 73 2767
rect -73 2713 73 2741
rect -73 2687 -67 2713
rect -41 2687 -13 2713
rect 13 2687 41 2713
rect 67 2687 73 2713
rect -73 2659 73 2687
rect -73 2633 -67 2659
rect -41 2633 -13 2659
rect 13 2633 41 2659
rect 67 2633 73 2659
rect -73 2605 73 2633
rect -73 2579 -67 2605
rect -41 2579 -13 2605
rect 13 2579 41 2605
rect 67 2579 73 2605
rect -73 2551 73 2579
rect -73 2525 -67 2551
rect -41 2525 -13 2551
rect 13 2525 41 2551
rect 67 2525 73 2551
rect -73 2497 73 2525
rect -73 2471 -67 2497
rect -41 2471 -13 2497
rect 13 2471 41 2497
rect 67 2471 73 2497
rect -73 2443 73 2471
rect -73 2417 -67 2443
rect -41 2417 -13 2443
rect 13 2417 41 2443
rect 67 2417 73 2443
rect -73 2389 73 2417
rect -73 2363 -67 2389
rect -41 2363 -13 2389
rect 13 2363 41 2389
rect 67 2363 73 2389
rect -73 2335 73 2363
rect -73 2309 -67 2335
rect -41 2309 -13 2335
rect 13 2309 41 2335
rect 67 2309 73 2335
rect -73 2281 73 2309
rect -73 2255 -67 2281
rect -41 2255 -13 2281
rect 13 2255 41 2281
rect 67 2255 73 2281
rect -73 2227 73 2255
rect -73 2201 -67 2227
rect -41 2201 -13 2227
rect 13 2201 41 2227
rect 67 2201 73 2227
rect -73 2173 73 2201
rect -73 2147 -67 2173
rect -41 2147 -13 2173
rect 13 2147 41 2173
rect 67 2147 73 2173
rect -73 2119 73 2147
rect -73 2093 -67 2119
rect -41 2093 -13 2119
rect 13 2093 41 2119
rect 67 2093 73 2119
rect -73 2065 73 2093
rect -73 2039 -67 2065
rect -41 2039 -13 2065
rect 13 2039 41 2065
rect 67 2039 73 2065
rect -73 2011 73 2039
rect -73 1985 -67 2011
rect -41 1985 -13 2011
rect 13 1985 41 2011
rect 67 1985 73 2011
rect -73 1957 73 1985
rect -73 1931 -67 1957
rect -41 1931 -13 1957
rect 13 1931 41 1957
rect 67 1931 73 1957
rect -73 1903 73 1931
rect -73 1877 -67 1903
rect -41 1877 -13 1903
rect 13 1877 41 1903
rect 67 1877 73 1903
rect -73 1849 73 1877
rect -73 1823 -67 1849
rect -41 1823 -13 1849
rect 13 1823 41 1849
rect 67 1823 73 1849
rect -73 1795 73 1823
rect -73 1769 -67 1795
rect -41 1769 -13 1795
rect 13 1769 41 1795
rect 67 1769 73 1795
rect -73 1741 73 1769
rect -73 1715 -67 1741
rect -41 1715 -13 1741
rect 13 1715 41 1741
rect 67 1715 73 1741
rect -73 1687 73 1715
rect -73 1661 -67 1687
rect -41 1661 -13 1687
rect 13 1661 41 1687
rect 67 1661 73 1687
rect -73 1633 73 1661
rect -73 1607 -67 1633
rect -41 1607 -13 1633
rect 13 1607 41 1633
rect 67 1607 73 1633
rect -73 1579 73 1607
rect -73 1553 -67 1579
rect -41 1553 -13 1579
rect 13 1553 41 1579
rect 67 1553 73 1579
rect -73 1525 73 1553
rect -73 1499 -67 1525
rect -41 1499 -13 1525
rect 13 1499 41 1525
rect 67 1499 73 1525
rect -73 1471 73 1499
rect -73 1445 -67 1471
rect -41 1445 -13 1471
rect 13 1445 41 1471
rect 67 1445 73 1471
rect -73 1417 73 1445
rect -73 1391 -67 1417
rect -41 1391 -13 1417
rect 13 1391 41 1417
rect 67 1391 73 1417
rect -73 1363 73 1391
rect -73 1337 -67 1363
rect -41 1337 -13 1363
rect 13 1337 41 1363
rect 67 1337 73 1363
rect -73 1309 73 1337
rect -73 1283 -67 1309
rect -41 1283 -13 1309
rect 13 1283 41 1309
rect 67 1283 73 1309
rect -73 1255 73 1283
rect -73 1229 -67 1255
rect -41 1229 -13 1255
rect 13 1229 41 1255
rect 67 1229 73 1255
rect -73 1201 73 1229
rect -73 1175 -67 1201
rect -41 1175 -13 1201
rect 13 1175 41 1201
rect 67 1175 73 1201
rect -73 1147 73 1175
rect -73 1121 -67 1147
rect -41 1121 -13 1147
rect 13 1121 41 1147
rect 67 1121 73 1147
rect -73 1093 73 1121
rect -73 1067 -67 1093
rect -41 1067 -13 1093
rect 13 1067 41 1093
rect 67 1067 73 1093
rect -73 1039 73 1067
rect -73 1013 -67 1039
rect -41 1013 -13 1039
rect 13 1013 41 1039
rect 67 1013 73 1039
rect -73 985 73 1013
rect -73 959 -67 985
rect -41 959 -13 985
rect 13 959 41 985
rect 67 959 73 985
rect -73 931 73 959
rect -73 905 -67 931
rect -41 905 -13 931
rect 13 905 41 931
rect 67 905 73 931
rect -73 877 73 905
rect -73 851 -67 877
rect -41 851 -13 877
rect 13 851 41 877
rect 67 851 73 877
rect -73 823 73 851
rect -73 797 -67 823
rect -41 797 -13 823
rect 13 797 41 823
rect 67 797 73 823
rect -73 769 73 797
rect -73 743 -67 769
rect -41 743 -13 769
rect 13 743 41 769
rect 67 743 73 769
rect -73 715 73 743
rect -73 689 -67 715
rect -41 689 -13 715
rect 13 689 41 715
rect 67 689 73 715
rect -73 661 73 689
rect -73 635 -67 661
rect -41 635 -13 661
rect 13 635 41 661
rect 67 635 73 661
rect -73 607 73 635
rect -73 581 -67 607
rect -41 581 -13 607
rect 13 581 41 607
rect 67 581 73 607
rect -73 553 73 581
rect -73 527 -67 553
rect -41 527 -13 553
rect 13 527 41 553
rect 67 527 73 553
rect -73 499 73 527
rect -73 473 -67 499
rect -41 473 -13 499
rect 13 473 41 499
rect 67 473 73 499
rect -73 445 73 473
rect -73 419 -67 445
rect -41 419 -13 445
rect 13 419 41 445
rect 67 419 73 445
rect -73 391 73 419
rect -73 365 -67 391
rect -41 365 -13 391
rect 13 365 41 391
rect 67 365 73 391
rect -73 337 73 365
rect -73 311 -67 337
rect -41 311 -13 337
rect 13 311 41 337
rect 67 311 73 337
rect -73 283 73 311
rect -73 257 -67 283
rect -41 257 -13 283
rect 13 257 41 283
rect 67 257 73 283
rect -73 229 73 257
rect -73 203 -67 229
rect -41 203 -13 229
rect 13 203 41 229
rect 67 203 73 229
rect -73 175 73 203
rect -73 149 -67 175
rect -41 149 -13 175
rect 13 149 41 175
rect 67 149 73 175
rect -73 121 73 149
rect -73 95 -67 121
rect -41 95 -13 121
rect 13 95 41 121
rect 67 95 73 121
rect -73 67 73 95
rect -73 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 73 67
rect -73 13 73 41
rect -73 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 73 13
rect -73 -41 73 -13
rect -73 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 73 -41
rect -73 -95 73 -67
rect -73 -121 -67 -95
rect -41 -121 -13 -95
rect 13 -121 41 -95
rect 67 -121 73 -95
rect -73 -149 73 -121
rect -73 -175 -67 -149
rect -41 -175 -13 -149
rect 13 -175 41 -149
rect 67 -175 73 -149
rect -73 -203 73 -175
rect -73 -229 -67 -203
rect -41 -229 -13 -203
rect 13 -229 41 -203
rect 67 -229 73 -203
rect -73 -257 73 -229
rect -73 -283 -67 -257
rect -41 -283 -13 -257
rect 13 -283 41 -257
rect 67 -283 73 -257
rect -73 -311 73 -283
rect -73 -337 -67 -311
rect -41 -337 -13 -311
rect 13 -337 41 -311
rect 67 -337 73 -311
rect -73 -365 73 -337
rect -73 -391 -67 -365
rect -41 -391 -13 -365
rect 13 -391 41 -365
rect 67 -391 73 -365
rect -73 -419 73 -391
rect -73 -445 -67 -419
rect -41 -445 -13 -419
rect 13 -445 41 -419
rect 67 -445 73 -419
rect -73 -473 73 -445
rect -73 -499 -67 -473
rect -41 -499 -13 -473
rect 13 -499 41 -473
rect 67 -499 73 -473
rect -73 -527 73 -499
rect -73 -553 -67 -527
rect -41 -553 -13 -527
rect 13 -553 41 -527
rect 67 -553 73 -527
rect -73 -581 73 -553
rect -73 -607 -67 -581
rect -41 -607 -13 -581
rect 13 -607 41 -581
rect 67 -607 73 -581
rect -73 -635 73 -607
rect -73 -661 -67 -635
rect -41 -661 -13 -635
rect 13 -661 41 -635
rect 67 -661 73 -635
rect -73 -689 73 -661
rect -73 -715 -67 -689
rect -41 -715 -13 -689
rect 13 -715 41 -689
rect 67 -715 73 -689
rect -73 -743 73 -715
rect -73 -769 -67 -743
rect -41 -769 -13 -743
rect 13 -769 41 -743
rect 67 -769 73 -743
rect -73 -797 73 -769
rect -73 -823 -67 -797
rect -41 -823 -13 -797
rect 13 -823 41 -797
rect 67 -823 73 -797
rect -73 -851 73 -823
rect -73 -877 -67 -851
rect -41 -877 -13 -851
rect 13 -877 41 -851
rect 67 -877 73 -851
rect -73 -905 73 -877
rect -73 -931 -67 -905
rect -41 -931 -13 -905
rect 13 -931 41 -905
rect 67 -931 73 -905
rect -73 -959 73 -931
rect -73 -985 -67 -959
rect -41 -985 -13 -959
rect 13 -985 41 -959
rect 67 -985 73 -959
rect -73 -1013 73 -985
rect -73 -1039 -67 -1013
rect -41 -1039 -13 -1013
rect 13 -1039 41 -1013
rect 67 -1039 73 -1013
rect -73 -1067 73 -1039
rect -73 -1093 -67 -1067
rect -41 -1093 -13 -1067
rect 13 -1093 41 -1067
rect 67 -1093 73 -1067
rect -73 -1121 73 -1093
rect -73 -1147 -67 -1121
rect -41 -1147 -13 -1121
rect 13 -1147 41 -1121
rect 67 -1147 73 -1121
rect -73 -1175 73 -1147
rect -73 -1201 -67 -1175
rect -41 -1201 -13 -1175
rect 13 -1201 41 -1175
rect 67 -1201 73 -1175
rect -73 -1229 73 -1201
rect -73 -1255 -67 -1229
rect -41 -1255 -13 -1229
rect 13 -1255 41 -1229
rect 67 -1255 73 -1229
rect -73 -1283 73 -1255
rect -73 -1309 -67 -1283
rect -41 -1309 -13 -1283
rect 13 -1309 41 -1283
rect 67 -1309 73 -1283
rect -73 -1337 73 -1309
rect -73 -1363 -67 -1337
rect -41 -1363 -13 -1337
rect 13 -1363 41 -1337
rect 67 -1363 73 -1337
rect -73 -1391 73 -1363
rect -73 -1417 -67 -1391
rect -41 -1417 -13 -1391
rect 13 -1417 41 -1391
rect 67 -1417 73 -1391
rect -73 -1445 73 -1417
rect -73 -1471 -67 -1445
rect -41 -1471 -13 -1445
rect 13 -1471 41 -1445
rect 67 -1471 73 -1445
rect -73 -1499 73 -1471
rect -73 -1525 -67 -1499
rect -41 -1525 -13 -1499
rect 13 -1525 41 -1499
rect 67 -1525 73 -1499
rect -73 -1553 73 -1525
rect -73 -1579 -67 -1553
rect -41 -1579 -13 -1553
rect 13 -1579 41 -1553
rect 67 -1579 73 -1553
rect -73 -1607 73 -1579
rect -73 -1633 -67 -1607
rect -41 -1633 -13 -1607
rect 13 -1633 41 -1607
rect 67 -1633 73 -1607
rect -73 -1661 73 -1633
rect -73 -1687 -67 -1661
rect -41 -1687 -13 -1661
rect 13 -1687 41 -1661
rect 67 -1687 73 -1661
rect -73 -1715 73 -1687
rect -73 -1741 -67 -1715
rect -41 -1741 -13 -1715
rect 13 -1741 41 -1715
rect 67 -1741 73 -1715
rect -73 -1769 73 -1741
rect -73 -1795 -67 -1769
rect -41 -1795 -13 -1769
rect 13 -1795 41 -1769
rect 67 -1795 73 -1769
rect -73 -1823 73 -1795
rect -73 -1849 -67 -1823
rect -41 -1849 -13 -1823
rect 13 -1849 41 -1823
rect 67 -1849 73 -1823
rect -73 -1877 73 -1849
rect -73 -1903 -67 -1877
rect -41 -1903 -13 -1877
rect 13 -1903 41 -1877
rect 67 -1903 73 -1877
rect -73 -1931 73 -1903
rect -73 -1957 -67 -1931
rect -41 -1957 -13 -1931
rect 13 -1957 41 -1931
rect 67 -1957 73 -1931
rect -73 -1985 73 -1957
rect -73 -2011 -67 -1985
rect -41 -2011 -13 -1985
rect 13 -2011 41 -1985
rect 67 -2011 73 -1985
rect -73 -2039 73 -2011
rect -73 -2065 -67 -2039
rect -41 -2065 -13 -2039
rect 13 -2065 41 -2039
rect 67 -2065 73 -2039
rect -73 -2093 73 -2065
rect -73 -2119 -67 -2093
rect -41 -2119 -13 -2093
rect 13 -2119 41 -2093
rect 67 -2119 73 -2093
rect -73 -2147 73 -2119
rect -73 -2173 -67 -2147
rect -41 -2173 -13 -2147
rect 13 -2173 41 -2147
rect 67 -2173 73 -2147
rect -73 -2201 73 -2173
rect -73 -2227 -67 -2201
rect -41 -2227 -13 -2201
rect 13 -2227 41 -2201
rect 67 -2227 73 -2201
rect -73 -2255 73 -2227
rect -73 -2281 -67 -2255
rect -41 -2281 -13 -2255
rect 13 -2281 41 -2255
rect 67 -2281 73 -2255
rect -73 -2309 73 -2281
rect -73 -2335 -67 -2309
rect -41 -2335 -13 -2309
rect 13 -2335 41 -2309
rect 67 -2335 73 -2309
rect -73 -2363 73 -2335
rect -73 -2389 -67 -2363
rect -41 -2389 -13 -2363
rect 13 -2389 41 -2363
rect 67 -2389 73 -2363
rect -73 -2417 73 -2389
rect -73 -2443 -67 -2417
rect -41 -2443 -13 -2417
rect 13 -2443 41 -2417
rect 67 -2443 73 -2417
rect -73 -2471 73 -2443
rect -73 -2497 -67 -2471
rect -41 -2497 -13 -2471
rect 13 -2497 41 -2471
rect 67 -2497 73 -2471
rect -73 -2525 73 -2497
rect -73 -2551 -67 -2525
rect -41 -2551 -13 -2525
rect 13 -2551 41 -2525
rect 67 -2551 73 -2525
rect -73 -2579 73 -2551
rect -73 -2605 -67 -2579
rect -41 -2605 -13 -2579
rect 13 -2605 41 -2579
rect 67 -2605 73 -2579
rect -73 -2633 73 -2605
rect -73 -2659 -67 -2633
rect -41 -2659 -13 -2633
rect 13 -2659 41 -2633
rect 67 -2659 73 -2633
rect -73 -2687 73 -2659
rect -73 -2713 -67 -2687
rect -41 -2713 -13 -2687
rect 13 -2713 41 -2687
rect 67 -2713 73 -2687
rect -73 -2741 73 -2713
rect -73 -2767 -67 -2741
rect -41 -2767 -13 -2741
rect 13 -2767 41 -2741
rect 67 -2767 73 -2741
rect -73 -2795 73 -2767
rect -73 -2821 -67 -2795
rect -41 -2821 -13 -2795
rect 13 -2821 41 -2795
rect 67 -2821 73 -2795
rect -73 -2849 73 -2821
rect -73 -2875 -67 -2849
rect -41 -2875 -13 -2849
rect 13 -2875 41 -2849
rect 67 -2875 73 -2849
rect -73 -2903 73 -2875
rect -73 -2929 -67 -2903
rect -41 -2929 -13 -2903
rect 13 -2929 41 -2903
rect 67 -2929 73 -2903
rect -73 -2957 73 -2929
rect -73 -2983 -67 -2957
rect -41 -2983 -13 -2957
rect 13 -2983 41 -2957
rect 67 -2983 73 -2957
rect -73 -3011 73 -2983
rect -73 -3037 -67 -3011
rect -41 -3037 -13 -3011
rect 13 -3037 41 -3011
rect 67 -3037 73 -3011
rect -73 -3065 73 -3037
rect -73 -3091 -67 -3065
rect -41 -3091 -13 -3065
rect 13 -3091 41 -3065
rect 67 -3091 73 -3065
rect -73 -3119 73 -3091
rect -73 -3145 -67 -3119
rect -41 -3145 -13 -3119
rect 13 -3145 41 -3119
rect 67 -3145 73 -3119
rect -73 -3173 73 -3145
rect -73 -3199 -67 -3173
rect -41 -3199 -13 -3173
rect 13 -3199 41 -3173
rect 67 -3199 73 -3173
rect -73 -3227 73 -3199
rect -73 -3253 -67 -3227
rect -41 -3253 -13 -3227
rect 13 -3253 41 -3227
rect 67 -3253 73 -3227
rect -73 -3281 73 -3253
rect -73 -3307 -67 -3281
rect -41 -3307 -13 -3281
rect 13 -3307 41 -3281
rect 67 -3307 73 -3281
rect -73 -3335 73 -3307
rect -73 -3361 -67 -3335
rect -41 -3361 -13 -3335
rect 13 -3361 41 -3335
rect 67 -3361 73 -3335
rect -73 -3389 73 -3361
rect -73 -3415 -67 -3389
rect -41 -3415 -13 -3389
rect 13 -3415 41 -3389
rect 67 -3415 73 -3389
rect -73 -3443 73 -3415
rect -73 -3469 -67 -3443
rect -41 -3469 -13 -3443
rect 13 -3469 41 -3443
rect 67 -3469 73 -3443
rect -73 -3497 73 -3469
rect -73 -3523 -67 -3497
rect -41 -3523 -13 -3497
rect 13 -3523 41 -3497
rect 67 -3523 73 -3497
rect -73 -3551 73 -3523
rect -73 -3577 -67 -3551
rect -41 -3577 -13 -3551
rect 13 -3577 41 -3551
rect 67 -3577 73 -3551
rect -73 -3605 73 -3577
rect -73 -3631 -67 -3605
rect -41 -3631 -13 -3605
rect 13 -3631 41 -3605
rect 67 -3631 73 -3605
rect -73 -3659 73 -3631
rect -73 -3685 -67 -3659
rect -41 -3685 -13 -3659
rect 13 -3685 41 -3659
rect 67 -3685 73 -3659
rect -73 -3713 73 -3685
rect -73 -3739 -67 -3713
rect -41 -3739 -13 -3713
rect 13 -3739 41 -3713
rect 67 -3739 73 -3713
rect -73 -3767 73 -3739
rect -73 -3793 -67 -3767
rect -41 -3793 -13 -3767
rect 13 -3793 41 -3767
rect 67 -3793 73 -3767
rect -73 -3821 73 -3793
rect -73 -3847 -67 -3821
rect -41 -3847 -13 -3821
rect 13 -3847 41 -3821
rect 67 -3847 73 -3821
rect -73 -3875 73 -3847
rect -73 -3901 -67 -3875
rect -41 -3901 -13 -3875
rect 13 -3901 41 -3875
rect 67 -3901 73 -3875
rect -73 -3929 73 -3901
rect -73 -3955 -67 -3929
rect -41 -3955 -13 -3929
rect 13 -3955 41 -3929
rect 67 -3955 73 -3929
rect -73 -3983 73 -3955
rect -73 -4009 -67 -3983
rect -41 -4009 -13 -3983
rect 13 -4009 41 -3983
rect 67 -4009 73 -3983
rect -73 -4037 73 -4009
rect -73 -4063 -67 -4037
rect -41 -4063 -13 -4037
rect 13 -4063 41 -4037
rect 67 -4063 73 -4037
rect -73 -4091 73 -4063
rect -73 -4117 -67 -4091
rect -41 -4117 -13 -4091
rect 13 -4117 41 -4091
rect 67 -4117 73 -4091
rect -73 -4145 73 -4117
rect -73 -4171 -67 -4145
rect -41 -4171 -13 -4145
rect 13 -4171 41 -4145
rect 67 -4171 73 -4145
rect -73 -4199 73 -4171
rect -73 -4225 -67 -4199
rect -41 -4225 -13 -4199
rect 13 -4225 41 -4199
rect 67 -4225 73 -4199
rect -73 -4253 73 -4225
rect -73 -4279 -67 -4253
rect -41 -4279 -13 -4253
rect 13 -4279 41 -4253
rect 67 -4279 73 -4253
rect -73 -4307 73 -4279
rect -73 -4333 -67 -4307
rect -41 -4333 -13 -4307
rect 13 -4333 41 -4307
rect 67 -4333 73 -4307
rect -73 -4361 73 -4333
rect -73 -4387 -67 -4361
rect -41 -4387 -13 -4361
rect 13 -4387 41 -4361
rect 67 -4387 73 -4361
rect -73 -4415 73 -4387
rect -73 -4441 -67 -4415
rect -41 -4441 -13 -4415
rect 13 -4441 41 -4415
rect 67 -4441 73 -4415
rect -73 -4469 73 -4441
rect -73 -4495 -67 -4469
rect -41 -4495 -13 -4469
rect 13 -4495 41 -4469
rect 67 -4495 73 -4469
rect -73 -4523 73 -4495
rect -73 -4549 -67 -4523
rect -41 -4549 -13 -4523
rect 13 -4549 41 -4523
rect 67 -4549 73 -4523
rect -73 -4577 73 -4549
rect -73 -4603 -67 -4577
rect -41 -4603 -13 -4577
rect 13 -4603 41 -4577
rect 67 -4603 73 -4577
rect -73 -4631 73 -4603
rect -73 -4657 -67 -4631
rect -41 -4657 -13 -4631
rect 13 -4657 41 -4631
rect 67 -4657 73 -4631
rect -73 -4685 73 -4657
rect -73 -4711 -67 -4685
rect -41 -4711 -13 -4685
rect 13 -4711 41 -4685
rect 67 -4711 73 -4685
rect -73 -4739 73 -4711
rect -73 -4765 -67 -4739
rect -41 -4765 -13 -4739
rect 13 -4765 41 -4739
rect 67 -4765 73 -4739
rect -73 -4793 73 -4765
rect -73 -4819 -67 -4793
rect -41 -4819 -13 -4793
rect 13 -4819 41 -4793
rect 67 -4819 73 -4793
rect -73 -4847 73 -4819
rect -73 -4873 -67 -4847
rect -41 -4873 -13 -4847
rect 13 -4873 41 -4847
rect 67 -4873 73 -4847
rect -73 -4901 73 -4873
rect -73 -4927 -67 -4901
rect -41 -4927 -13 -4901
rect 13 -4927 41 -4901
rect 67 -4927 73 -4901
rect -73 -4955 73 -4927
rect -73 -4981 -67 -4955
rect -41 -4981 -13 -4955
rect 13 -4981 41 -4955
rect 67 -4981 73 -4955
rect -73 -5009 73 -4981
rect -73 -5035 -67 -5009
rect -41 -5035 -13 -5009
rect 13 -5035 41 -5009
rect 67 -5035 73 -5009
rect -73 -5063 73 -5035
rect -73 -5089 -67 -5063
rect -41 -5089 -13 -5063
rect 13 -5089 41 -5063
rect 67 -5089 73 -5063
rect -73 -5117 73 -5089
rect -73 -5143 -67 -5117
rect -41 -5143 -13 -5117
rect 13 -5143 41 -5117
rect 67 -5143 73 -5117
rect -73 -5171 73 -5143
rect -73 -5197 -67 -5171
rect -41 -5197 -13 -5171
rect 13 -5197 41 -5171
rect 67 -5197 73 -5171
rect -73 -5225 73 -5197
rect -73 -5251 -67 -5225
rect -41 -5251 -13 -5225
rect 13 -5251 41 -5225
rect 67 -5251 73 -5225
rect -73 -5279 73 -5251
rect -73 -5305 -67 -5279
rect -41 -5305 -13 -5279
rect 13 -5305 41 -5279
rect 67 -5305 73 -5279
rect -73 -5333 73 -5305
rect -73 -5359 -67 -5333
rect -41 -5359 -13 -5333
rect 13 -5359 41 -5333
rect 67 -5359 73 -5333
rect -73 -5387 73 -5359
rect -73 -5413 -67 -5387
rect -41 -5413 -13 -5387
rect 13 -5413 41 -5387
rect 67 -5413 73 -5387
rect -73 -5441 73 -5413
rect -73 -5467 -67 -5441
rect -41 -5467 -13 -5441
rect 13 -5467 41 -5441
rect 67 -5467 73 -5441
rect -73 -5495 73 -5467
rect -73 -5521 -67 -5495
rect -41 -5521 -13 -5495
rect 13 -5521 41 -5495
rect 67 -5521 73 -5495
rect -73 -5549 73 -5521
rect -73 -5575 -67 -5549
rect -41 -5575 -13 -5549
rect 13 -5575 41 -5549
rect 67 -5575 73 -5549
rect -73 -5603 73 -5575
rect -73 -5629 -67 -5603
rect -41 -5629 -13 -5603
rect 13 -5629 41 -5603
rect 67 -5629 73 -5603
rect -73 -5657 73 -5629
rect -73 -5683 -67 -5657
rect -41 -5683 -13 -5657
rect 13 -5683 41 -5657
rect 67 -5683 73 -5657
rect -73 -5711 73 -5683
rect -73 -5737 -67 -5711
rect -41 -5737 -13 -5711
rect 13 -5737 41 -5711
rect 67 -5737 73 -5711
rect -73 -5765 73 -5737
rect -73 -5791 -67 -5765
rect -41 -5791 -13 -5765
rect 13 -5791 41 -5765
rect 67 -5791 73 -5765
rect -73 -5819 73 -5791
rect -73 -5845 -67 -5819
rect -41 -5845 -13 -5819
rect 13 -5845 41 -5819
rect 67 -5845 73 -5819
rect -73 -5873 73 -5845
rect -73 -5899 -67 -5873
rect -41 -5899 -13 -5873
rect 13 -5899 41 -5873
rect 67 -5899 73 -5873
rect -73 -5927 73 -5899
rect -73 -5953 -67 -5927
rect -41 -5953 -13 -5927
rect 13 -5953 41 -5927
rect 67 -5953 73 -5927
rect -73 -5981 73 -5953
rect -73 -6007 -67 -5981
rect -41 -6007 -13 -5981
rect 13 -6007 41 -5981
rect 67 -6007 73 -5981
rect -73 -6013 73 -6007
<< end >>
