magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1721 1019 1721
<< metal1 >>
rect -19 715 19 721
rect -19 -715 -13 715
rect 13 -715 19 715
rect -19 -721 19 -715
<< via1 >>
rect -13 -715 13 715
<< metal2 >>
rect -19 715 19 721
rect -19 -715 -13 715
rect 13 -715 19 715
rect -19 -721 19 -715
<< end >>
