magic
tech gf180mcuC
magscale 1 10
timestamp 1694675087
<< nwell >>
rect -282 -365 282 365
<< pmos >>
rect -108 -235 -52 235
rect 52 -235 108 235
<< pdiff >>
rect -196 222 -108 235
rect -196 -222 -183 222
rect -137 -222 -108 222
rect -196 -235 -108 -222
rect -52 222 52 235
rect -52 -222 -23 222
rect 23 -222 52 222
rect -52 -235 52 -222
rect 108 222 196 235
rect 108 -222 137 222
rect 183 -222 196 222
rect 108 -235 196 -222
<< pdiffc >>
rect -183 -222 -137 222
rect -23 -222 23 222
rect 137 -222 183 222
<< polysilicon >>
rect -108 235 -52 279
rect 52 235 108 279
rect -108 -279 -52 -235
rect 52 -279 108 -235
<< metal1 >>
rect -183 222 -137 233
rect -183 -233 -137 -222
rect -23 222 23 233
rect -23 -233 23 -222
rect 137 222 183 233
rect 137 -233 183 -222
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2.35 l 0.280 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
