magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1539 1019 1539
<< metal2 >>
rect -19 534 19 539
rect -19 -534 -14 534
rect 14 -534 19 534
rect -19 -539 19 -534
<< via2 >>
rect -14 -534 14 534
<< metal3 >>
rect -19 534 19 539
rect -19 -534 -14 534
rect 14 -534 19 534
rect -19 -539 19 -534
<< end >>
