magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1374 1019 1374
<< metal2 >>
rect -19 369 19 374
rect -19 341 -14 369
rect 14 341 19 369
rect -19 298 19 341
rect -19 270 -14 298
rect 14 270 19 298
rect -19 227 19 270
rect -19 199 -14 227
rect 14 199 19 227
rect -19 156 19 199
rect -19 128 -14 156
rect 14 128 19 156
rect -19 85 19 128
rect -19 57 -14 85
rect 14 57 19 85
rect -19 14 19 57
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -57 19 -14
rect -19 -85 -14 -57
rect 14 -85 19 -57
rect -19 -128 19 -85
rect -19 -156 -14 -128
rect 14 -156 19 -128
rect -19 -199 19 -156
rect -19 -227 -14 -199
rect 14 -227 19 -199
rect -19 -270 19 -227
rect -19 -298 -14 -270
rect 14 -298 19 -270
rect -19 -341 19 -298
rect -19 -369 -14 -341
rect 14 -369 19 -341
rect -19 -374 19 -369
<< via2 >>
rect -14 341 14 369
rect -14 270 14 298
rect -14 199 14 227
rect -14 128 14 156
rect -14 57 14 85
rect -14 -14 14 14
rect -14 -85 14 -57
rect -14 -156 14 -128
rect -14 -227 14 -199
rect -14 -298 14 -270
rect -14 -369 14 -341
<< metal3 >>
rect -19 369 19 374
rect -19 341 -14 369
rect 14 341 19 369
rect -19 298 19 341
rect -19 270 -14 298
rect 14 270 19 298
rect -19 227 19 270
rect -19 199 -14 227
rect 14 199 19 227
rect -19 156 19 199
rect -19 128 -14 156
rect 14 128 19 156
rect -19 85 19 128
rect -19 57 -14 85
rect 14 57 19 85
rect -19 14 19 57
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -57 19 -14
rect -19 -85 -14 -57
rect 14 -85 19 -57
rect -19 -128 19 -85
rect -19 -156 -14 -128
rect 14 -156 19 -128
rect -19 -199 19 -156
rect -19 -227 -14 -199
rect 14 -227 19 -199
rect -19 -270 19 -227
rect -19 -298 -14 -270
rect 14 -298 19 -270
rect -19 -341 19 -298
rect -19 -369 -14 -341
rect 14 -369 19 -341
rect -19 -374 19 -369
<< end >>
