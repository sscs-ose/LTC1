* NGSPICE file created from Inv_16x_Layout_flat.ext - technology: gf180mcuC

.subckt Inv_16x_Layout_flat IN OUT VSS VDD
X0 OUT IN.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.194p pd=1.76u as=0.194p ps=1.76u w=0.44u l=2.24u
X1 OUT IN.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=2.24u
R0 IN.n0 IN.t1 17.8546
R1 IN IN.n0 14.0337
R2 IN.n0 IN.t0 13.5862
R3 VDD.n8 VDD.t0 282.663
R4 VDD.n0 VDD.t1 7.06752
R5 VDD.n4 VDD.n3 3.1505
R6 VDD.n2 VDD.n1 3.1505
R7 VDD.n9 VDD.n5 2.18581
R8 VDD.n7 VDD.n5 1.78473
R9 VDD.n9 VDD.n8 1.44481
R10 VDD.n8 VDD.n7 0.684132
R11 VDD.n8 VDD.n6 0.684132
R12 VDD VDD.n9 0.215997
R13 VDD VDD.n4 0.0760357
R14 VDD.n4 VDD.n2 0.0760357
R15 VDD.n2 VDD.n0 0.0366607
R16 OUT OUT.n1 9.60502
R17 OUT OUT.n0 7.16491
R18 VSS.n1 VSS.t0 604.271
R19 VSS.n5 VSS.t1 9.32958
R20 VSS.n8 VSS.n3 9.13939
R21 VSS VSS.n3 5.2005
R22 VSS VSS.n3 5.2005
R23 VSS.n5 VSS.n4 2.60371
R24 VSS.n9 VSS.n8 2.6005
R25 VSS.n7 VSS.n6 2.6005
R26 VSS.n3 VSS.n2 1.92228
R27 VSS VSS.n2 1.62146
R28 VSS.n1 VSS.n0 0.472445
R29 VSS.n2 VSS.n1 0.173689
R30 VSS VSS.n9 0.0760357
R31 VSS.n9 VSS.n7 0.0760357
R32 VSS.n7 VSS.n5 0.0728214
C0 OUT VDD 0.0656f
C1 OUT IN 0.0486f
C2 VDD IN 0.429f
.ends

