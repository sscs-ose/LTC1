magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2478 -2278 2478 2278
<< nwell >>
rect -478 -278 478 278
<< nsubdiff >>
rect -395 173 395 195
rect -395 -173 -373 173
rect 373 -173 395 173
rect -395 -195 395 -173
<< nsubdiffcont >>
rect -373 -173 373 173
<< metal1 >>
rect -384 173 384 184
rect -384 -173 -373 173
rect 373 -173 384 173
rect -384 -184 384 -173
<< end >>
