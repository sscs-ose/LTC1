magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1267 -1174 1267 1174
<< metal1 >>
rect -267 168 267 174
rect -267 142 -261 168
rect -235 142 -199 168
rect -173 142 -137 168
rect -111 142 -75 168
rect -49 142 -13 168
rect 13 142 49 168
rect 75 142 111 168
rect 137 142 173 168
rect 199 142 235 168
rect 261 142 267 168
rect -267 106 267 142
rect -267 80 -261 106
rect -235 80 -199 106
rect -173 80 -137 106
rect -111 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 111 106
rect 137 80 173 106
rect 199 80 235 106
rect 261 80 267 106
rect -267 44 267 80
rect -267 18 -261 44
rect -235 18 -199 44
rect -173 18 -137 44
rect -111 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 111 44
rect 137 18 173 44
rect 199 18 235 44
rect 261 18 267 44
rect -267 -18 267 18
rect -267 -44 -261 -18
rect -235 -44 -199 -18
rect -173 -44 -137 -18
rect -111 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 111 -18
rect 137 -44 173 -18
rect 199 -44 235 -18
rect 261 -44 267 -18
rect -267 -80 267 -44
rect -267 -106 -261 -80
rect -235 -106 -199 -80
rect -173 -106 -137 -80
rect -111 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 111 -80
rect 137 -106 173 -80
rect 199 -106 235 -80
rect 261 -106 267 -80
rect -267 -142 267 -106
rect -267 -168 -261 -142
rect -235 -168 -199 -142
rect -173 -168 -137 -142
rect -111 -168 -75 -142
rect -49 -168 -13 -142
rect 13 -168 49 -142
rect 75 -168 111 -142
rect 137 -168 173 -142
rect 199 -168 235 -142
rect 261 -168 267 -142
rect -267 -174 267 -168
<< via1 >>
rect -261 142 -235 168
rect -199 142 -173 168
rect -137 142 -111 168
rect -75 142 -49 168
rect -13 142 13 168
rect 49 142 75 168
rect 111 142 137 168
rect 173 142 199 168
rect 235 142 261 168
rect -261 80 -235 106
rect -199 80 -173 106
rect -137 80 -111 106
rect -75 80 -49 106
rect -13 80 13 106
rect 49 80 75 106
rect 111 80 137 106
rect 173 80 199 106
rect 235 80 261 106
rect -261 18 -235 44
rect -199 18 -173 44
rect -137 18 -111 44
rect -75 18 -49 44
rect -13 18 13 44
rect 49 18 75 44
rect 111 18 137 44
rect 173 18 199 44
rect 235 18 261 44
rect -261 -44 -235 -18
rect -199 -44 -173 -18
rect -137 -44 -111 -18
rect -75 -44 -49 -18
rect -13 -44 13 -18
rect 49 -44 75 -18
rect 111 -44 137 -18
rect 173 -44 199 -18
rect 235 -44 261 -18
rect -261 -106 -235 -80
rect -199 -106 -173 -80
rect -137 -106 -111 -80
rect -75 -106 -49 -80
rect -13 -106 13 -80
rect 49 -106 75 -80
rect 111 -106 137 -80
rect 173 -106 199 -80
rect 235 -106 261 -80
rect -261 -168 -235 -142
rect -199 -168 -173 -142
rect -137 -168 -111 -142
rect -75 -168 -49 -142
rect -13 -168 13 -142
rect 49 -168 75 -142
rect 111 -168 137 -142
rect 173 -168 199 -142
rect 235 -168 261 -142
<< metal2 >>
rect -267 168 267 174
rect -267 142 -261 168
rect -235 142 -199 168
rect -173 142 -137 168
rect -111 142 -75 168
rect -49 142 -13 168
rect 13 142 49 168
rect 75 142 111 168
rect 137 142 173 168
rect 199 142 235 168
rect 261 142 267 168
rect -267 106 267 142
rect -267 80 -261 106
rect -235 80 -199 106
rect -173 80 -137 106
rect -111 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 111 106
rect 137 80 173 106
rect 199 80 235 106
rect 261 80 267 106
rect -267 44 267 80
rect -267 18 -261 44
rect -235 18 -199 44
rect -173 18 -137 44
rect -111 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 111 44
rect 137 18 173 44
rect 199 18 235 44
rect 261 18 267 44
rect -267 -18 267 18
rect -267 -44 -261 -18
rect -235 -44 -199 -18
rect -173 -44 -137 -18
rect -111 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 111 -18
rect 137 -44 173 -18
rect 199 -44 235 -18
rect 261 -44 267 -18
rect -267 -80 267 -44
rect -267 -106 -261 -80
rect -235 -106 -199 -80
rect -173 -106 -137 -80
rect -111 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 111 -80
rect 137 -106 173 -80
rect 199 -106 235 -80
rect 261 -106 267 -80
rect -267 -142 267 -106
rect -267 -168 -261 -142
rect -235 -168 -199 -142
rect -173 -168 -137 -142
rect -111 -168 -75 -142
rect -49 -168 -13 -142
rect 13 -168 49 -142
rect 75 -168 111 -142
rect 137 -168 173 -142
rect 199 -168 235 -142
rect 261 -168 267 -142
rect -267 -174 267 -168
<< end >>
