magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2109 -2677 2109 2677
<< metal2 >>
rect -109 667 109 677
rect -109 611 -99 667
rect -43 611 43 667
rect 99 611 109 667
rect -109 525 109 611
rect -109 469 -99 525
rect -43 469 43 525
rect 99 469 109 525
rect -109 383 109 469
rect -109 327 -99 383
rect -43 327 43 383
rect 99 327 109 383
rect -109 241 109 327
rect -109 185 -99 241
rect -43 185 43 241
rect 99 185 109 241
rect -109 99 109 185
rect -109 43 -99 99
rect -43 43 43 99
rect 99 43 109 99
rect -109 -43 109 43
rect -109 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 109 -43
rect -109 -185 109 -99
rect -109 -241 -99 -185
rect -43 -241 43 -185
rect 99 -241 109 -185
rect -109 -327 109 -241
rect -109 -383 -99 -327
rect -43 -383 43 -327
rect 99 -383 109 -327
rect -109 -469 109 -383
rect -109 -525 -99 -469
rect -43 -525 43 -469
rect 99 -525 109 -469
rect -109 -611 109 -525
rect -109 -667 -99 -611
rect -43 -667 43 -611
rect 99 -667 109 -611
rect -109 -677 109 -667
<< via2 >>
rect -99 611 -43 667
rect 43 611 99 667
rect -99 469 -43 525
rect 43 469 99 525
rect -99 327 -43 383
rect 43 327 99 383
rect -99 185 -43 241
rect 43 185 99 241
rect -99 43 -43 99
rect 43 43 99 99
rect -99 -99 -43 -43
rect 43 -99 99 -43
rect -99 -241 -43 -185
rect 43 -241 99 -185
rect -99 -383 -43 -327
rect 43 -383 99 -327
rect -99 -525 -43 -469
rect 43 -525 99 -469
rect -99 -667 -43 -611
rect 43 -667 99 -611
<< metal3 >>
rect -109 667 109 677
rect -109 611 -99 667
rect -43 611 43 667
rect 99 611 109 667
rect -109 525 109 611
rect -109 469 -99 525
rect -43 469 43 525
rect 99 469 109 525
rect -109 383 109 469
rect -109 327 -99 383
rect -43 327 43 383
rect 99 327 109 383
rect -109 241 109 327
rect -109 185 -99 241
rect -43 185 43 241
rect 99 185 109 241
rect -109 99 109 185
rect -109 43 -99 99
rect -43 43 43 99
rect 99 43 109 99
rect -109 -43 109 43
rect -109 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 109 -43
rect -109 -185 109 -99
rect -109 -241 -99 -185
rect -43 -241 43 -185
rect 99 -241 109 -185
rect -109 -327 109 -241
rect -109 -383 -99 -327
rect -43 -383 43 -327
rect 99 -383 109 -327
rect -109 -469 109 -383
rect -109 -525 -99 -469
rect -43 -525 43 -469
rect 99 -525 109 -469
rect -109 -611 109 -525
rect -109 -667 -99 -611
rect -43 -667 43 -611
rect 99 -667 109 -611
rect -109 -677 109 -667
<< end >>
