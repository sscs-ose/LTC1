* NGSPICE file created from INVERTER_MUX_flat.ext - technology: gf180mcuC

.subckt INVERTER_MUX_flat VDD VSS IN OUT
X0 OUT IN.t0 VDD.t15 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 OUT IN.t1 VSS.t15 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 OUT IN.t2 VDD.t14 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 VDD IN.t3 OUT.t5 VDD.t7 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X4 VSS IN.t4 OUT.t15 VSS.t10 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 OUT IN.t5 VDD.t11 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 VDD IN.t6 OUT.t3 VDD.t7 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X7 VSS IN.t7 OUT.t14 VSS.t10 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X8 OUT IN.t8 VSS.t9 VSS.t5 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X9 VSS IN.t9 OUT.t13 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X10 VDD IN.t10 OUT.t2 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X11 OUT IN.t11 VSS.t6 VSS.t5 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X12 OUT IN.t12 VDD.t4 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X13 VSS IN.t13 OUT.t12 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X14 VDD IN.t14 OUT.t0 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X15 OUT IN.t15 VSS.t1 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 IN.t3 IN.t6 43.8005
R1 IN.t12 IN.t0 43.8005
R2 IN.t10 IN.t14 43.8005
R3 IN.t2 IN.t5 43.8005
R4 IN.t7 IN.t4 30.7648
R5 IN.t11 IN.t8 30.7648
R6 IN.t13 IN.t9 30.7648
R7 IN.t1 IN.t15 30.7648
R8 IN.n0 IN.t7 30.3737
R9 IN.n1 IN.t11 30.3737
R10 IN.n2 IN.t13 30.3737
R11 IN.n0 IN.t3 21.6398
R12 IN.n1 IN.t12 21.6398
R13 IN.n2 IN.t10 21.6398
R14 IN.n3 IN.t2 21.6398
R15 IN.n4 IN.t1 17.7827
R16 IN.n1 IN.n0 17.255
R17 IN.n2 IN.n1 17.255
R18 IN.n3 IN.n2 17.255
R19 IN.n4 IN.n3 8.06475
R20 IN IN.n4 4.24369
R21 VDD.t3 VDD.t7 171.124
R22 VDD.t0 VDD.t10 171.124
R23 VDD.n9 VDD.t3 91.9791
R24 VDD.n9 VDD.t0 79.1449
R25 VDD.n13 VDD.t14 5.07789
R26 VDD.n7 VDD.n6 5.07789
R27 VDD.n13 VDD.t11 4.4205
R28 VDD.n7 VDD.n5 4.4205
R29 VDD.n4 VDD.n3 3.25789
R30 VDD.n12 VDD.n11 3.1505
R31 VDD.n11 VDD.n9 3.1505
R32 VDD.n4 VDD.n1 2.6005
R33 VDD.n1 VDD.t15 1.8205
R34 VDD.n1 VDD.n0 1.8205
R35 VDD.n3 VDD.t4 1.8205
R36 VDD.n3 VDD.n2 1.8205
R37 VDD.n8 VDD.n7 0.657694
R38 VDD VDD.n13 0.652514
R39 VDD.n8 VDD.n4 0.4505
R40 VDD.n11 VDD.n10 0.1405
R41 VDD.n12 VDD.n8 0.00438489
R42 VDD VDD.n12 0.00179496
R43 OUT.n9 OUT.n8 3.61224
R44 OUT.n19 OUT.n18 3.61224
R45 OUT.n6 OUT.t14 3.2765
R46 OUT.n6 OUT.n5 3.2765
R47 OUT.n8 OUT.t15 3.2765
R48 OUT.n8 OUT.n7 3.2765
R49 OUT.n16 OUT.t12 3.2765
R50 OUT.n16 OUT.n15 3.2765
R51 OUT.n18 OUT.t13 3.2765
R52 OUT.n18 OUT.n17 3.2765
R53 OUT.n4 OUT.n1 3.25789
R54 OUT.n14 OUT.n11 3.25789
R55 OUT.n9 OUT.n6 3.1505
R56 OUT.n19 OUT.n16 3.1505
R57 OUT.n4 OUT.n3 2.6005
R58 OUT.n14 OUT.n13 2.6005
R59 OUT.n3 OUT.t5 1.8205
R60 OUT.n3 OUT.n2 1.8205
R61 OUT.n1 OUT.t3 1.8205
R62 OUT.n1 OUT.n0 1.8205
R63 OUT.n11 OUT.t0 1.8205
R64 OUT.n11 OUT.n10 1.8205
R65 OUT.n13 OUT.t2 1.8205
R66 OUT.n13 OUT.n12 1.8205
R67 OUT.n21 OUT.n20 0.626587
R68 OUT OUT.n21 0.487674
R69 OUT.n21 OUT.n4 0.427022
R70 OUT.n20 OUT.n14 0.427022
R71 OUT.n21 OUT.n9 0.26463
R72 OUT.n20 OUT.n19 0.26463
R73 VSS.t5 VSS.t10 771.514
R74 VSS.t2 VSS.t0 771.514
R75 VSS.n9 VSS.t5 414.688
R76 VSS.n9 VSS.t2 356.825
R77 VSS.n7 VSS.n5 6.88824
R78 VSS.n13 VSS.t15 6.88824
R79 VSS.n7 VSS.n6 6.4265
R80 VSS.n13 VSS.t1 6.4265
R81 VSS.n4 VSS.n1 3.61224
R82 VSS.n3 VSS.t9 3.2765
R83 VSS.n3 VSS.n2 3.2765
R84 VSS.n1 VSS.t6 3.2765
R85 VSS.n1 VSS.n0 3.2765
R86 VSS.n4 VSS.n3 3.1505
R87 VSS.n12 VSS.n11 2.6005
R88 VSS.n11 VSS.n9 2.6005
R89 VSS.n11 VSS.n10 0.846654
R90 VSS.n8 VSS.n7 0.462042
R91 VSS VSS.n13 0.451035
R92 VSS.n8 VSS.n4 0.254848
R93 VSS VSS.n12 0.0076223
R94 VSS.n12 VSS.n8 0.00438489
C0 VDD OUT 1.02f
C1 VDD IN 0.852f
C2 IN OUT 0.307f
.ends

