* NGSPICE file created from folded_cascode_check1_flat.ext - technology: gf180mcuC

.subckt folded_cascode_check1_flat VDD
X0 VDD a_n2679_n1703# a_n2983_n1659.t30 VDD.t2 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X1 a_n2983_n1659.t15 a_n2983_n1659.t14 a_n2983_n1659.t15 VDD.t1 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X2 VDD a_n2679_n1703# a_n2983_n1659.t26 VDD.t4 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X3 VDD a_n2679_n1703# a_n2983_n1659.t25 VDD.t4 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X4 a_n2983_n1659.t13 a_n2983_n1659.t12 a_n2983_n1659.t13 VDD.t1 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X5 a_n2983_n1659.t11 a_n2983_n1659.t10 a_n2983_n1659.t11 VDD.t1 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X6 VDD a_n2679_n1703# a_n2983_n1659.t24 VDD.t4 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X7 a_n2983_n1659.t9 a_n2983_n1659.t8 a_n2983_n1659.t9 VDD.t1 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X8 a_n2983_n1659.t7 a_n2983_n1659.t6 a_n2983_n1659.t7 VDD.t0 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X9 VDD a_n2679_n1703# a_n2983_n1659.t19 VDD.t2 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X10 a_n2983_n1659.t5 a_n2983_n1659.t4 a_n2983_n1659.t5 VDD.t0 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X11 a_n2983_n1659.t3 a_n2983_n1659.t2 a_n2983_n1659.t3 VDD.t0 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
X12 VDD a_n2679_n1703# a_n2983_n1659.t18 VDD.t4 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X13 VDD a_n2679_n1703# a_n2983_n1659.t17 VDD.t2 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X14 VDD a_n2679_n1703# a_n2983_n1659.t16 VDD.t2 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X15 a_n2983_n1659.t1 a_n2983_n1659.t0 a_n2983_n1659.t1 VDD.t0 pfet_03v3 ad=0 pd=0 as=1.32p ps=6.88u w=3u l=0.56u
R0 VDD.n126 VDD.t4 12.698
R1 VDD.n107 VDD.t0 11.005
R2 VDD.n136 VDD.t15 5.92601
R3 VDD.n120 VDD.t8 4.79734
R4 VDD.n241 VDD.n240 3.1505
R5 VDD.n243 VDD.n242 3.1505
R6 VDD.n196 VDD.n195 3.1505
R7 VDD.n79 VDD.n78 3.1505
R8 VDD.n76 VDD.n75 3.1505
R9 VDD.n73 VDD.n72 3.1505
R10 VDD.n71 VDD.n70 3.1505
R11 VDD.n68 VDD.n67 3.1505
R12 VDD.n66 VDD.n65 3.1505
R13 VDD.n63 VDD.n62 3.1505
R14 VDD.n61 VDD.n60 3.1505
R15 VDD.n58 VDD.n57 3.1505
R16 VDD.n56 VDD.n55 3.1505
R17 VDD.n53 VDD.n52 3.1505
R18 VDD.n51 VDD.n50 3.1505
R19 VDD.n48 VDD.n47 3.1505
R20 VDD.n46 VDD.n45 3.1505
R21 VDD.n43 VDD.n42 3.1505
R22 VDD.n41 VDD.n40 3.1505
R23 VDD.n39 VDD.n38 3.1505
R24 VDD.n37 VDD.n36 3.1505
R25 VDD.n35 VDD.n34 3.1505
R26 VDD.n33 VDD.n32 3.1505
R27 VDD.n31 VDD.n30 3.1505
R28 VDD.n29 VDD.n28 3.1505
R29 VDD.n27 VDD.n26 3.1505
R30 VDD.n25 VDD.n24 3.1505
R31 VDD.n23 VDD.n22 3.1505
R32 VDD.n21 VDD.n20 3.1505
R33 VDD.n19 VDD.n18 3.1505
R34 VDD.n182 VDD.n181 3.1505
R35 VDD.n184 VDD.n183 3.1505
R36 VDD.n186 VDD.n185 3.1505
R37 VDD.n188 VDD.n187 3.1505
R38 VDD.n191 VDD.n190 3.1505
R39 VDD.n193 VDD.n192 3.1505
R40 VDD.n81 VDD.n80 3.1505
R41 VDD.n239 VDD.n238 3.1505
R42 VDD.n237 VDD.n236 3.1505
R43 VDD.n235 VDD.n234 3.1505
R44 VDD.n233 VDD.n232 3.1505
R45 VDD.n231 VDD.n230 3.1505
R46 VDD.n229 VDD.n228 3.1505
R47 VDD.n223 VDD.n222 3.1505
R48 VDD.n221 VDD.n220 3.1505
R49 VDD.n219 VDD.n218 3.1505
R50 VDD.n217 VDD.n216 3.1505
R51 VDD.n214 VDD.n213 3.1505
R52 VDD.n212 VDD.n211 3.1505
R53 VDD.n210 VDD.n209 3.1505
R54 VDD.n208 VDD.n207 3.1505
R55 VDD.n206 VDD.n205 3.1505
R56 VDD.n204 VDD.n203 3.1505
R57 VDD.n202 VDD.n201 3.1505
R58 VDD.n200 VDD.n199 3.1505
R59 VDD.n198 VDD.n197 3.1505
R60 VDD.n152 VDD.n151 3.1505
R61 VDD.n97 VDD.n96 3.1505
R62 VDD.n96 VDD.n95 3.1505
R63 VDD.n100 VDD.n99 3.1505
R64 VDD.n99 VDD.n98 3.1505
R65 VDD.n103 VDD.n102 3.1505
R66 VDD.n102 VDD.n101 3.1505
R67 VDD.n106 VDD.n105 3.1505
R68 VDD.n105 VDD.n104 3.1505
R69 VDD.n109 VDD.n108 3.1505
R70 VDD.n108 VDD.n107 3.1505
R71 VDD.n112 VDD.n111 3.1505
R72 VDD.n111 VDD.n110 3.1505
R73 VDD.n115 VDD.n114 3.1505
R74 VDD.n114 VDD.n113 3.1505
R75 VDD.n118 VDD.n117 3.1505
R76 VDD.n117 VDD.n116 3.1505
R77 VDD.n122 VDD.n121 3.1505
R78 VDD.n121 VDD.n120 3.1505
R79 VDD.n125 VDD.n124 3.1505
R80 VDD.n124 VDD.n123 3.1505
R81 VDD.n128 VDD.n127 3.1505
R82 VDD.n127 VDD.n126 3.1505
R83 VDD.n131 VDD.n130 3.1505
R84 VDD.n130 VDD.n129 3.1505
R85 VDD.n135 VDD.n134 3.1505
R86 VDD.n134 VDD.n133 3.1505
R87 VDD.n138 VDD.n137 3.1505
R88 VDD.n137 VDD.n136 3.1505
R89 VDD.n141 VDD.n140 3.1505
R90 VDD.n140 VDD.n139 3.1505
R91 VDD.n144 VDD.n143 3.1505
R92 VDD.n143 VDD.n142 3.1505
R93 VDD.n147 VDD.n146 3.1505
R94 VDD.n146 VDD.n145 3.1505
R95 VDD.n150 VDD.n149 3.1505
R96 VDD.n149 VDD.n148 3.1505
R97 VDD.n153 VDD.n152 3.1505
R98 VDD.n156 VDD.n155 3.1505
R99 VDD.n155 VDD.n154 3.1505
R100 VDD.n158 VDD.n157 3.1505
R101 VDD.n94 VDD.n93 3.1505
R102 VDD.n248 VDD.n247 3.1505
R103 VDD.n250 VDD.n249 3.1505
R104 VDD.n253 VDD.n252 3.1505
R105 VDD.n256 VDD.n255 3.1505
R106 VDD.n259 VDD.n258 3.1505
R107 VDD.n262 VDD.n261 3.1505
R108 VDD.n265 VDD.n264 3.1505
R109 VDD.n268 VDD.n267 3.1505
R110 VDD.n271 VDD.n270 3.1505
R111 VDD.n274 VDD.n273 3.1505
R112 VDD.n277 VDD.n276 3.1505
R113 VDD.n280 VDD.n279 3.1505
R114 VDD.n283 VDD.n282 3.1505
R115 VDD.n286 VDD.n285 3.1505
R116 VDD.n289 VDD.n288 3.1505
R117 VDD.n292 VDD.n291 3.1505
R118 VDD.n295 VDD.n294 3.1505
R119 VDD.n298 VDD.n297 3.1505
R120 VDD.n301 VDD.n300 3.1505
R121 VDD.n304 VDD.n303 3.1505
R122 VDD.n307 VDD.n306 3.1505
R123 VDD.n310 VDD.n309 3.1505
R124 VDD.n313 VDD.n312 3.1505
R125 VDD.n316 VDD.n315 3.1505
R126 VDD.n319 VDD.n318 3.1505
R127 VDD.n322 VDD.n321 3.1505
R128 VDD.n325 VDD.n324 3.1505
R129 VDD.n328 VDD.n327 3.1505
R130 VDD.n332 VDD.n331 3.1505
R131 VDD.n177 VDD.n176 3.1505
R132 VDD.n174 VDD.n173 3.1505
R133 VDD.n171 VDD.n170 3.1505
R134 VDD.n168 VDD.n167 3.1505
R135 VDD.n165 VDD.n164 3.1505
R136 VDD.n163 VDD.n162 3.1505
R137 VDD.n245 VDD.n244 3.1505
R138 VDD.n113 VDD.t2 3.10434
R139 VDD.n180 VDD.n179 2.6005
R140 VDD.n15 VDD.n14 2.6005
R141 VDD.n16 VDD.n12 2.6005
R142 VDD.n17 VDD.n10 2.6005
R143 VDD.n226 VDD.n225 2.6005
R144 VDD.n6 VDD.n5 2.6005
R145 VDD.n7 VDD.n3 2.6005
R146 VDD.n8 VDD.n1 2.6005
R147 VDD.n167 VDD.n166 2.40832
R148 VDD.n170 VDD.n169 2.40832
R149 VDD.n173 VDD.n172 2.40832
R150 VDD.n176 VDD.n175 2.40832
R151 VDD.n331 VDD.n329 2.40832
R152 VDD.n331 VDD.n330 2.40832
R153 VDD.n327 VDD.n326 2.40832
R154 VDD.n324 VDD.n323 2.40832
R155 VDD.n321 VDD.n320 2.40832
R156 VDD.n318 VDD.n317 2.40832
R157 VDD.n315 VDD.n314 2.40832
R158 VDD.n312 VDD.n311 2.40832
R159 VDD.n309 VDD.n308 2.40832
R160 VDD.n306 VDD.n305 2.40832
R161 VDD.n303 VDD.n302 2.40832
R162 VDD.n300 VDD.n299 2.40832
R163 VDD.n297 VDD.n296 2.40832
R164 VDD.n294 VDD.n293 2.40832
R165 VDD.n291 VDD.n290 2.40832
R166 VDD.n288 VDD.n287 2.40832
R167 VDD.n285 VDD.n284 2.40832
R168 VDD.n282 VDD.n281 2.40832
R169 VDD.n279 VDD.n278 2.40832
R170 VDD.n276 VDD.n275 2.40832
R171 VDD.n273 VDD.n272 2.40832
R172 VDD.n270 VDD.n269 2.40832
R173 VDD.n267 VDD.n266 2.40832
R174 VDD.n264 VDD.n263 2.40832
R175 VDD.n261 VDD.n260 2.40832
R176 VDD.n258 VDD.n257 2.40832
R177 VDD.n255 VDD.n254 2.40832
R178 VDD.n252 VDD.n251 2.40832
R179 VDD.n142 VDD.t1 1.97567
R180 VDD.n75 VDD.n74 1.74343
R181 VDD.n70 VDD.n69 1.74343
R182 VDD.n65 VDD.n64 1.74343
R183 VDD.n60 VDD.n59 1.74343
R184 VDD.n55 VDD.n54 1.74343
R185 VDD.n50 VDD.n49 1.74343
R186 VDD.n45 VDD.n44 1.74343
R187 VDD.n162 VDD.n161 1.42472
R188 VDD.n247 VDD.n246 1.42456
R189 VDD.n78 VDD.n77 1.42456
R190 VDD.n190 VDD.n189 1.42456
R191 VDD.n195 VDD.n194 1.42456
R192 VDD.n92 VDD.n91 1.40117
R193 VDD.n17 VDD.n16 1.27435
R194 VDD.n16 VDD.n15 1.27435
R195 VDD.n8 VDD.n7 1.27435
R196 VDD.n7 VDD.n6 1.27435
R197 VDD.n161 VDD.n160 1.15215
R198 VDD.n93 VDD.n92 1.0512
R199 VDD.n215 VDD.n180 0.968
R200 VDD.n227 VDD.n226 0.968
R201 VDD.n119 VDD.n17 0.9005
R202 VDD.n132 VDD.n8 0.9005
R203 VDD.n91 VDD.n90 0.705355
R204 VDD.n91 VDD.n89 0.705355
R205 VDD.n91 VDD.n88 0.705355
R206 VDD.n91 VDD.n87 0.705355
R207 VDD.n91 VDD.n86 0.705355
R208 VDD.n91 VDD.n85 0.705355
R209 VDD.n91 VDD.n84 0.705355
R210 VDD.n91 VDD.n83 0.705355
R211 VDD.n1 VDD.t26 0.607167
R212 VDD.n1 VDD.n0 0.607167
R213 VDD.n3 VDD.t17 0.607167
R214 VDD.n3 VDD.n2 0.607167
R215 VDD.n5 VDD.t16 0.607167
R216 VDD.n5 VDD.n4 0.607167
R217 VDD.n225 VDD.t29 0.607167
R218 VDD.n225 VDD.n224 0.607167
R219 VDD.n10 VDD.t18 0.607167
R220 VDD.n10 VDD.n9 0.607167
R221 VDD.n12 VDD.t25 0.607167
R222 VDD.n12 VDD.n11 0.607167
R223 VDD.n14 VDD.t24 0.607167
R224 VDD.n14 VDD.n13 0.607167
R225 VDD.n179 VDD.t9 0.607167
R226 VDD.n179 VDD.n178 0.607167
R227 VDD.n160 VDD.n159 0.282667
R228 VDD.n91 VDD.n82 0.282667
R229 VDD VDD.n333 0.121376
R230 VDD.n97 VDD.n94 0.0877449
R231 VDD.n307 VDD.n304 0.0868265
R232 VDD.n81 VDD.n79 0.0868265
R233 VDD.n79 VDD.n76 0.0868265
R234 VDD.n76 VDD.n73 0.0868265
R235 VDD.n73 VDD.n71 0.0868265
R236 VDD.n71 VDD.n68 0.0868265
R237 VDD.n68 VDD.n66 0.0868265
R238 VDD.n66 VDD.n63 0.0868265
R239 VDD.n63 VDD.n61 0.0868265
R240 VDD.n61 VDD.n58 0.0868265
R241 VDD.n58 VDD.n56 0.0868265
R242 VDD.n56 VDD.n53 0.0868265
R243 VDD.n53 VDD.n51 0.0868265
R244 VDD.n51 VDD.n48 0.0868265
R245 VDD.n48 VDD.n46 0.0868265
R246 VDD.n46 VDD.n43 0.0868265
R247 VDD.n43 VDD.n41 0.0868265
R248 VDD.n41 VDD.n39 0.0868265
R249 VDD.n39 VDD.n37 0.0868265
R250 VDD.n37 VDD.n35 0.0868265
R251 VDD.n35 VDD.n33 0.0868265
R252 VDD.n33 VDD.n31 0.0868265
R253 VDD.n31 VDD.n29 0.0868265
R254 VDD.n29 VDD.n27 0.0868265
R255 VDD.n27 VDD.n25 0.0868265
R256 VDD.n25 VDD.n23 0.0868265
R257 VDD.n23 VDD.n21 0.0868265
R258 VDD.n21 VDD.n19 0.0868265
R259 VDD.n184 VDD.n182 0.0868265
R260 VDD.n186 VDD.n184 0.0868265
R261 VDD.n188 VDD.n186 0.0868265
R262 VDD.n191 VDD.n188 0.0868265
R263 VDD.n193 VDD.n191 0.0868265
R264 VDD.n196 VDD.n193 0.0868265
R265 VDD.n239 VDD.n237 0.0868265
R266 VDD.n237 VDD.n235 0.0868265
R267 VDD.n235 VDD.n233 0.0868265
R268 VDD.n233 VDD.n231 0.0868265
R269 VDD.n231 VDD.n229 0.0868265
R270 VDD.n223 VDD.n221 0.0868265
R271 VDD.n221 VDD.n219 0.0868265
R272 VDD.n219 VDD.n217 0.0868265
R273 VDD.n214 VDD.n212 0.0868265
R274 VDD.n212 VDD.n210 0.0868265
R275 VDD.n210 VDD.n208 0.0868265
R276 VDD.n208 VDD.n206 0.0868265
R277 VDD.n206 VDD.n204 0.0868265
R278 VDD.n204 VDD.n202 0.0868265
R279 VDD.n202 VDD.n200 0.0868265
R280 VDD.n200 VDD.n198 0.0868265
R281 VDD.n158 VDD.n156 0.0868265
R282 VDD.n156 VDD.n153 0.0868265
R283 VDD.n153 VDD.n150 0.0868265
R284 VDD.n150 VDD.n147 0.0868265
R285 VDD.n147 VDD.n144 0.0868265
R286 VDD.n144 VDD.n141 0.0868265
R287 VDD.n141 VDD.n138 0.0868265
R288 VDD.n138 VDD.n135 0.0868265
R289 VDD.n131 VDD.n128 0.0868265
R290 VDD.n128 VDD.n125 0.0868265
R291 VDD.n125 VDD.n122 0.0868265
R292 VDD.n118 VDD.n115 0.0868265
R293 VDD.n115 VDD.n112 0.0868265
R294 VDD.n112 VDD.n109 0.0868265
R295 VDD.n109 VDD.n106 0.0868265
R296 VDD.n106 VDD.n103 0.0868265
R297 VDD.n103 VDD.n100 0.0868265
R298 VDD.n100 VDD.n97 0.0868265
R299 VDD.n165 VDD.n163 0.0868265
R300 VDD.n168 VDD.n165 0.0868265
R301 VDD.n171 VDD.n168 0.0868265
R302 VDD.n174 VDD.n171 0.0868265
R303 VDD.n177 VDD.n174 0.0868265
R304 VDD.n332 VDD.n328 0.0868265
R305 VDD.n328 VDD.n325 0.0868265
R306 VDD.n325 VDD.n322 0.0868265
R307 VDD.n322 VDD.n319 0.0868265
R308 VDD.n319 VDD.n316 0.0868265
R309 VDD.n316 VDD.n313 0.0868265
R310 VDD.n313 VDD.n310 0.0868265
R311 VDD.n310 VDD.n307 0.0868265
R312 VDD.n304 VDD.n301 0.0868265
R313 VDD.n301 VDD.n298 0.0868265
R314 VDD.n298 VDD.n295 0.0868265
R315 VDD.n295 VDD.n292 0.0868265
R316 VDD.n292 VDD.n289 0.0868265
R317 VDD.n289 VDD.n286 0.0868265
R318 VDD.n286 VDD.n283 0.0868265
R319 VDD.n283 VDD.n280 0.0868265
R320 VDD.n280 VDD.n277 0.0868265
R321 VDD.n277 VDD.n274 0.0868265
R322 VDD.n274 VDD.n271 0.0868265
R323 VDD.n271 VDD.n268 0.0868265
R324 VDD.n268 VDD.n265 0.0868265
R325 VDD.n265 VDD.n262 0.0868265
R326 VDD.n262 VDD.n259 0.0868265
R327 VDD.n259 VDD.n256 0.0868265
R328 VDD.n256 VDD.n253 0.0868265
R329 VDD.n253 VDD.n250 0.0868265
R330 VDD.n250 VDD.n248 0.0868265
R331 VDD.n248 VDD.n245 0.0868265
R332 VDD.n217 VDD.n215 0.0840714
R333 VDD.n122 VDD.n119 0.0840714
R334 VDD.n333 VDD.n177 0.0712143
R335 VDD.n227 VDD.n223 0.0546837
R336 VDD.n132 VDD.n131 0.0546837
R337 VDD.n241 VDD.n239 0.0482121
R338 VDD.n163 VDD.n158 0.0436633
R339 VDD.n94 VDD.n81 0.0427449
R340 VDD.n198 VDD.n196 0.0427449
R341 VDD.n229 VDD.n227 0.0326429
R342 VDD.n135 VDD.n132 0.0326429
R343 VDD.n245 VDD.n243 0.0293783
R344 VDD.n243 VDD.n241 0.0170234
R345 VDD.n333 VDD.n332 0.0161122
R346 VDD.n215 VDD.n214 0.0032551
R347 VDD.n119 VDD.n118 0.0032551
R348 a_n2983_n1659.n27 a_n2983_n1659.t0 23.9862
R349 a_n2983_n1659.n42 a_n2983_n1659.t6 23.9862
R350 a_n2983_n1659.n42 a_n2983_n1659.t2 23.9862
R351 a_n2983_n1659.n32 a_n2983_n1659.t4 23.9862
R352 a_n2983_n1659.n53 a_n2983_n1659.t14 23.9862
R353 a_n2983_n1659.n53 a_n2983_n1659.t12 23.9862
R354 a_n2983_n1659.n4 a_n2983_n1659.t10 23.9862
R355 a_n2983_n1659.n0 a_n2983_n1659.t8 23.9862
R356 a_n2983_n1659.n48 a_n2983_n1659.n47 6.23075
R357 a_n2983_n1659.n47 a_n2983_n1659.n46 6.22569
R358 a_n2983_n1659.n47 a_n2983_n1659.n25 5.8995
R359 a_n2983_n1659.n28 a_n2983_n1659.n27 4.0005
R360 a_n2983_n1659.n33 a_n2983_n1659.n32 4.0005
R361 a_n2983_n1659.n43 a_n2983_n1659.n42 4.0005
R362 a_n2983_n1659.n1 a_n2983_n1659.n0 4.0005
R363 a_n2983_n1659.n5 a_n2983_n1659.n4 4.0005
R364 a_n2983_n1659.n54 a_n2983_n1659.n53 4.0005
R365 a_n2983_n1659.n19 a_n2983_n1659.n16 3.87435
R366 a_n2983_n1659.t15 a_n2983_n1659.n8 3.79909
R367 a_n2983_n1659.n57 a_n2983_n1659.n55 3.19242
R368 a_n2983_n1659.n29 a_n2983_n1659.n26 3.19069
R369 a_n2983_n1659.n31 a_n2983_n1659.n30 2.6005
R370 a_n2983_n1659.n36 a_n2983_n1659.n35 2.6005
R371 a_n2983_n1659.n46 a_n2983_n1659.n45 2.6005
R372 a_n2983_n1659.n25 a_n2983_n1659.n24 2.6005
R373 a_n2983_n1659.n22 a_n2983_n1659.n21 2.6005
R374 a_n2983_n1659.n19 a_n2983_n1659.n18 2.6005
R375 a_n2983_n1659.n48 a_n2983_n1659.n14 2.6005
R376 a_n2983_n1659.n52 a_n2983_n1659.n10 2.6005
R377 a_n2983_n1659.n50 a_n2983_n1659.n12 2.6005
R378 a_n2983_n1659.n22 a_n2983_n1659.n19 1.27435
R379 a_n2983_n1659.n25 a_n2983_n1659.n22 1.27435
R380 a_n2983_n1659.n12 a_n2983_n1659.t11 0.607167
R381 a_n2983_n1659.n12 a_n2983_n1659.n11 0.607167
R382 a_n2983_n1659.n14 a_n2983_n1659.t9 0.607167
R383 a_n2983_n1659.n14 a_n2983_n1659.n13 0.607167
R384 a_n2983_n1659.n45 a_n2983_n1659.t30 0.607167
R385 a_n2983_n1659.n45 a_n2983_n1659.t7 0.607167
R386 a_n2983_n1659.n35 a_n2983_n1659.t16 0.607167
R387 a_n2983_n1659.n35 a_n2983_n1659.t3 0.607167
R388 a_n2983_n1659.n30 a_n2983_n1659.t17 0.607167
R389 a_n2983_n1659.n30 a_n2983_n1659.t5 0.607167
R390 a_n2983_n1659.n26 a_n2983_n1659.t19 0.607167
R391 a_n2983_n1659.n26 a_n2983_n1659.t1 0.607167
R392 a_n2983_n1659.n16 a_n2983_n1659.t24 0.607167
R393 a_n2983_n1659.n16 a_n2983_n1659.n15 0.607167
R394 a_n2983_n1659.n18 a_n2983_n1659.t26 0.607167
R395 a_n2983_n1659.n18 a_n2983_n1659.n17 0.607167
R396 a_n2983_n1659.n21 a_n2983_n1659.t25 0.607167
R397 a_n2983_n1659.n21 a_n2983_n1659.n20 0.607167
R398 a_n2983_n1659.n24 a_n2983_n1659.t18 0.607167
R399 a_n2983_n1659.n24 a_n2983_n1659.n23 0.607167
R400 a_n2983_n1659.n10 a_n2983_n1659.t13 0.607167
R401 a_n2983_n1659.n10 a_n2983_n1659.n9 0.607167
R402 a_n2983_n1659.t15 a_n2983_n1659.n57 0.607167
R403 a_n2983_n1659.n57 a_n2983_n1659.n56 0.607167
R404 a_n2983_n1659.n38 a_n2983_n1659.n37 0.590692
R405 a_n2983_n1659.n39 a_n2983_n1659.n38 0.590692
R406 a_n2983_n1659.n31 a_n2983_n1659.n29 0.590692
R407 a_n2983_n1659.n34 a_n2983_n1659.n31 0.590692
R408 a_n2983_n1659.n36 a_n2983_n1659.n34 0.590692
R409 a_n2983_n1659.n44 a_n2983_n1659.n36 0.590692
R410 a_n2983_n1659.n40 a_n2983_n1659.n39 0.590692
R411 a_n2983_n1659.n41 a_n2983_n1659.n40 0.590692
R412 a_n2983_n1659.n46 a_n2983_n1659.n44 0.590692
R413 a_n2983_n1659.n49 a_n2983_n1659.n48 0.590692
R414 a_n2983_n1659.n6 a_n2983_n1659.n3 0.590692
R415 a_n2983_n1659.n3 a_n2983_n1659.n2 0.590692
R416 a_n2983_n1659.n52 a_n2983_n1659.n51 0.590692
R417 a_n2983_n1659.n51 a_n2983_n1659.n50 0.590692
R418 a_n2983_n1659.n50 a_n2983_n1659.n49 0.590692
R419 a_n2983_n1659.n7 a_n2983_n1659.n6 0.590692
R420 a_n2983_n1659.n55 a_n2983_n1659.n52 0.588962
R421 a_n2983_n1659.n8 a_n2983_n1659.n7 0.588962
R422 a_n2983_n1659.n29 a_n2983_n1659.n28 0.183833
R423 a_n2983_n1659.n34 a_n2983_n1659.n33 0.183833
R424 a_n2983_n1659.n44 a_n2983_n1659.n43 0.182167
R425 a_n2983_n1659.n55 a_n2983_n1659.n54 0.1805
R426 a_n2983_n1659.n43 a_n2983_n1659.n41 0.178833
R427 a_n2983_n1659.n2 a_n2983_n1659.n1 0.178833
R428 a_n2983_n1659.n6 a_n2983_n1659.n5 0.178833
C0 a_n2679_n1703# VDD 7.64f
C1 VDD VSUBS 24.6f
C2 a_n2679_n1703# VSUBS 1.32f
C3 a_n2983_n1659.t8 VSUBS 0.174f
C4 a_n2983_n1659.n0 VSUBS 0.146f
C5 a_n2983_n1659.n1 VSUBS 0.0206f
C6 a_n2983_n1659.n2 VSUBS 0.172f
C7 a_n2983_n1659.n3 VSUBS 0.0875f
C8 a_n2983_n1659.t10 VSUBS 0.146f
C9 a_n2983_n1659.n4 VSUBS 0.146f
C10 a_n2983_n1659.n5 VSUBS 0.0206f
C11 a_n2983_n1659.n6 VSUBS 0.0778f
C12 a_n2983_n1659.n7 VSUBS 0.0874f
C13 a_n2983_n1659.n8 VSUBS 0.172f
C14 a_n2983_n1659.t13 VSUBS 0.217f
C15 a_n2983_n1659.n9 VSUBS 0.0551f
C16 a_n2983_n1659.n10 VSUBS 0.11f
C17 a_n2983_n1659.t11 VSUBS 0.217f
C18 a_n2983_n1659.n11 VSUBS 0.0551f
C19 a_n2983_n1659.n12 VSUBS 0.11f
C20 a_n2983_n1659.t9 VSUBS 0.234f
C21 a_n2983_n1659.n13 VSUBS 0.0551f
C22 a_n2983_n1659.n14 VSUBS 0.11f
C23 a_n2983_n1659.t24 VSUBS 0.0551f
C24 a_n2983_n1659.n15 VSUBS 0.0551f
C25 a_n2983_n1659.n16 VSUBS 0.151f
C26 a_n2983_n1659.t26 VSUBS 0.0551f
C27 a_n2983_n1659.n17 VSUBS 0.0551f
C28 a_n2983_n1659.n18 VSUBS 0.11f
C29 a_n2983_n1659.n19 VSUBS 0.218f
C30 a_n2983_n1659.t25 VSUBS 0.0551f
C31 a_n2983_n1659.n20 VSUBS 0.0551f
C32 a_n2983_n1659.n21 VSUBS 0.11f
C33 a_n2983_n1659.n22 VSUBS 0.135f
C34 a_n2983_n1659.t18 VSUBS 0.0551f
C35 a_n2983_n1659.n23 VSUBS 0.0551f
C36 a_n2983_n1659.n24 VSUBS 0.11f
C37 a_n2983_n1659.n25 VSUBS 0.209f
C38 a_n2983_n1659.t19 VSUBS 0.0551f
C39 a_n2983_n1659.t1 VSUBS 0.234f
C40 a_n2983_n1659.n26 VSUBS 0.126f
C41 a_n2983_n1659.t0 VSUBS 0.174f
C42 a_n2983_n1659.n27 VSUBS 0.146f
C43 a_n2983_n1659.n28 VSUBS 0.0206f
C44 a_n2983_n1659.n29 VSUBS 0.149f
C45 a_n2983_n1659.t17 VSUBS 0.0551f
C46 a_n2983_n1659.t5 VSUBS 0.217f
C47 a_n2983_n1659.n30 VSUBS 0.11f
C48 a_n2983_n1659.n31 VSUBS 0.0626f
C49 a_n2983_n1659.t4 VSUBS 0.146f
C50 a_n2983_n1659.n32 VSUBS 0.146f
C51 a_n2983_n1659.n33 VSUBS 0.0206f
C52 a_n2983_n1659.n34 VSUBS 0.0781f
C53 a_n2983_n1659.t16 VSUBS 0.0551f
C54 a_n2983_n1659.t3 VSUBS 0.217f
C55 a_n2983_n1659.n35 VSUBS 0.11f
C56 a_n2983_n1659.n36 VSUBS 0.0626f
C57 a_n2983_n1659.n37 VSUBS 0.172f
C58 a_n2983_n1659.n38 VSUBS 0.0875f
C59 a_n2983_n1659.n39 VSUBS 0.0777f
C60 a_n2983_n1659.n40 VSUBS 0.0875f
C61 a_n2983_n1659.n41 VSUBS 0.172f
C62 a_n2983_n1659.t2 VSUBS 0.146f
C63 a_n2983_n1659.t6 VSUBS 0.174f
C64 a_n2983_n1659.n42 VSUBS 0.146f
C65 a_n2983_n1659.n43 VSUBS 0.0206f
C66 a_n2983_n1659.n44 VSUBS 0.078f
C67 a_n2983_n1659.t30 VSUBS 0.0551f
C68 a_n2983_n1659.t7 VSUBS 0.234f
C69 a_n2983_n1659.n45 VSUBS 0.11f
C70 a_n2983_n1659.n46 VSUBS 0.21f
C71 a_n2983_n1659.n47 VSUBS 1.14f
C72 a_n2983_n1659.n48 VSUBS 0.184f
C73 a_n2983_n1659.n49 VSUBS 0.078f
C74 a_n2983_n1659.n50 VSUBS 0.0626f
C75 a_n2983_n1659.n51 VSUBS 0.078f
C76 a_n2983_n1659.n52 VSUBS 0.0625f
C77 a_n2983_n1659.t14 VSUBS 0.174f
C78 a_n2983_n1659.t12 VSUBS 0.146f
C79 a_n2983_n1659.n53 VSUBS 0.146f
C80 a_n2983_n1659.n54 VSUBS 0.0206f
C81 a_n2983_n1659.n55 VSUBS 0.148f
C82 a_n2983_n1659.n56 VSUBS 0.0551f
C83 a_n2983_n1659.n57 VSUBS 0.126f
C84 a_n2983_n1659.t15 VSUBS 0.234f
C85 VDD.t26 VSUBS 0.0201f
C86 VDD.n0 VSUBS 0.0201f
C87 VDD.n1 VSUBS 0.0403f
C88 VDD.t17 VSUBS 0.0201f
C89 VDD.n2 VSUBS 0.0201f
C90 VDD.n3 VSUBS 0.0403f
C91 VDD.t16 VSUBS 0.0201f
C92 VDD.n4 VSUBS 0.0201f
C93 VDD.n5 VSUBS 0.0403f
C94 VDD.n6 VSUBS 0.0494f
C95 VDD.n7 VSUBS 0.0494f
C96 VDD.n8 VSUBS 0.0422f
C97 VDD.t18 VSUBS 0.0201f
C98 VDD.n9 VSUBS 0.0201f
C99 VDD.n10 VSUBS 0.0403f
C100 VDD.t25 VSUBS 0.0201f
C101 VDD.n11 VSUBS 0.0201f
C102 VDD.n12 VSUBS 0.0403f
C103 VDD.t24 VSUBS 0.0201f
C104 VDD.n13 VSUBS 0.0201f
C105 VDD.n14 VSUBS 0.0403f
C106 VDD.n15 VSUBS 0.0494f
C107 VDD.n16 VSUBS 0.0494f
C108 VDD.n17 VSUBS 0.0422f
C109 VDD.n18 VSUBS 0.00922f
C110 VDD.n19 VSUBS 0.0119f
C111 VDD.n20 VSUBS 0.00922f
C112 VDD.n21 VSUBS 0.0119f
C113 VDD.n22 VSUBS 0.00922f
C114 VDD.n23 VSUBS 0.0119f
C115 VDD.n24 VSUBS 0.00922f
C116 VDD.n25 VSUBS 0.0119f
C117 VDD.n26 VSUBS 0.00922f
C118 VDD.n27 VSUBS 0.0119f
C119 VDD.n28 VSUBS 0.00922f
C120 VDD.n29 VSUBS 0.0119f
C121 VDD.n30 VSUBS 0.00922f
C122 VDD.n31 VSUBS 0.0119f
C123 VDD.n32 VSUBS 0.00922f
C124 VDD.n33 VSUBS 0.0119f
C125 VDD.n34 VSUBS 0.00922f
C126 VDD.n35 VSUBS 0.0119f
C127 VDD.n36 VSUBS 0.00922f
C128 VDD.n37 VSUBS 0.0119f
C129 VDD.n38 VSUBS 0.00922f
C130 VDD.n39 VSUBS 0.0119f
C131 VDD.n40 VSUBS 0.00922f
C132 VDD.n41 VSUBS 0.0119f
C133 VDD.n42 VSUBS 0.00922f
C134 VDD.n43 VSUBS 0.0119f
C135 VDD.n45 VSUBS 0.00922f
C136 VDD.n46 VSUBS 0.0119f
C137 VDD.n47 VSUBS 0.00922f
C138 VDD.n48 VSUBS 0.0119f
C139 VDD.n50 VSUBS 0.00922f
C140 VDD.n51 VSUBS 0.0119f
C141 VDD.n52 VSUBS 0.00922f
C142 VDD.n53 VSUBS 0.0119f
C143 VDD.n55 VSUBS 0.00922f
C144 VDD.n56 VSUBS 0.0119f
C145 VDD.n57 VSUBS 0.00922f
C146 VDD.n58 VSUBS 0.0119f
C147 VDD.n60 VSUBS 0.00922f
C148 VDD.n61 VSUBS 0.0119f
C149 VDD.n62 VSUBS 0.00922f
C150 VDD.n63 VSUBS 0.0119f
C151 VDD.n65 VSUBS 0.00922f
C152 VDD.n66 VSUBS 0.0119f
C153 VDD.n67 VSUBS 0.00922f
C154 VDD.n68 VSUBS 0.0119f
C155 VDD.n70 VSUBS 0.00922f
C156 VDD.n71 VSUBS 0.0119f
C157 VDD.n72 VSUBS 0.00922f
C158 VDD.n73 VSUBS 0.0119f
C159 VDD.n75 VSUBS 0.00922f
C160 VDD.n76 VSUBS 0.0119f
C161 VDD.n78 VSUBS 0.00922f
C162 VDD.n79 VSUBS 0.0119f
C163 VDD.n80 VSUBS 0.00741f
C164 VDD.n81 VSUBS 0.00886f
C165 VDD.n82 VSUBS 0.217f
C166 VDD.n91 VSUBS 0.391f
C167 VDD.n93 VSUBS 0.0112f
C168 VDD.n94 VSUBS 0.0151f
C169 VDD.n95 VSUBS 0.43f
C170 VDD.n96 VSUBS 0.00927f
C171 VDD.n97 VSUBS 0.012f
C172 VDD.n98 VSUBS 0.43f
C173 VDD.n99 VSUBS 0.00922f
C174 VDD.n100 VSUBS 0.0119f
C175 VDD.n101 VSUBS 0.43f
C176 VDD.n102 VSUBS 0.00922f
C177 VDD.n103 VSUBS 0.0119f
C178 VDD.n104 VSUBS 0.341f
C179 VDD.n105 VSUBS 0.00922f
C180 VDD.n106 VSUBS 0.0119f
C181 VDD.t0 VSUBS 0.215f
C182 VDD.n107 VSUBS 0.304f
C183 VDD.n108 VSUBS 0.00922f
C184 VDD.n109 VSUBS 0.0119f
C185 VDD.n110 VSUBS 0.405f
C186 VDD.n111 VSUBS 0.00922f
C187 VDD.n112 VSUBS 0.0119f
C188 VDD.t2 VSUBS 0.215f
C189 VDD.n113 VSUBS 0.24f
C190 VDD.n114 VSUBS 0.00922f
C191 VDD.n115 VSUBS 0.0119f
C192 VDD.n116 VSUBS 0.43f
C193 VDD.n117 VSUBS 0.00922f
C194 VDD.n118 VSUBS 0.00614f
C195 VDD.n119 VSUBS 0.0234f
C196 VDD.t8 VSUBS 0.215f
C197 VDD.n120 VSUBS 0.254f
C198 VDD.n121 VSUBS 0.00922f
C199 VDD.n122 VSUBS 0.0117f
C200 VDD.n123 VSUBS 0.391f
C201 VDD.n124 VSUBS 0.00922f
C202 VDD.n125 VSUBS 0.0119f
C203 VDD.t4 VSUBS 0.215f
C204 VDD.n126 VSUBS 0.318f
C205 VDD.n127 VSUBS 0.00922f
C206 VDD.n128 VSUBS 0.0119f
C207 VDD.n129 VSUBS 0.327f
C208 VDD.n130 VSUBS 0.00922f
C209 VDD.n131 VSUBS 0.00968f
C210 VDD.n132 VSUBS 0.0234f
C211 VDD.n133 VSUBS 0.382f
C212 VDD.n134 VSUBS 0.00922f
C213 VDD.n135 VSUBS 0.00816f
C214 VDD.t15 VSUBS 0.215f
C215 VDD.n136 VSUBS 0.263f
C216 VDD.n137 VSUBS 0.00922f
C217 VDD.n138 VSUBS 0.0119f
C218 VDD.n139 VSUBS 0.43f
C219 VDD.n140 VSUBS 0.00922f
C220 VDD.n141 VSUBS 0.0119f
C221 VDD.t1 VSUBS 0.215f
C222 VDD.n142 VSUBS 0.231f
C223 VDD.n143 VSUBS 0.00922f
C224 VDD.n144 VSUBS 0.0119f
C225 VDD.n145 VSUBS 0.414f
C226 VDD.n146 VSUBS 0.00922f
C227 VDD.n147 VSUBS 0.0119f
C228 VDD.n148 VSUBS 0.43f
C229 VDD.n149 VSUBS 0.00922f
C230 VDD.n150 VSUBS 0.0119f
C231 VDD.n151 VSUBS 0.43f
C232 VDD.n152 VSUBS 0.00922f
C233 VDD.n153 VSUBS 0.0119f
C234 VDD.n154 VSUBS 0.43f
C235 VDD.n155 VSUBS 0.00922f
C236 VDD.n156 VSUBS 0.0119f
C237 VDD.n157 VSUBS 0.0111f
C238 VDD.n158 VSUBS 0.015f
C239 VDD.n159 VSUBS 0.217f
C240 VDD.n160 VSUBS 0.332f
C241 VDD.n162 VSUBS 0.00752f
C242 VDD.n163 VSUBS 0.00905f
C243 VDD.n164 VSUBS 0.00922f
C244 VDD.n165 VSUBS 0.0119f
C245 VDD.n167 VSUBS 0.00922f
C246 VDD.n168 VSUBS 0.0119f
C247 VDD.n170 VSUBS 0.00922f
C248 VDD.n171 VSUBS 0.0119f
C249 VDD.n173 VSUBS 0.00922f
C250 VDD.n174 VSUBS 0.0119f
C251 VDD.n176 VSUBS 0.00922f
C252 VDD.n177 VSUBS 0.0108f
C253 VDD.t9 VSUBS 0.0201f
C254 VDD.n178 VSUBS 0.0201f
C255 VDD.n179 VSUBS 0.0403f
C256 VDD.n180 VSUBS 0.0435f
C257 VDD.n181 VSUBS 0.00922f
C258 VDD.n182 VSUBS 0.0119f
C259 VDD.n183 VSUBS 0.00922f
C260 VDD.n184 VSUBS 0.0119f
C261 VDD.n185 VSUBS 0.00922f
C262 VDD.n186 VSUBS 0.0119f
C263 VDD.n187 VSUBS 0.00922f
C264 VDD.n188 VSUBS 0.0119f
C265 VDD.n190 VSUBS 0.00922f
C266 VDD.n191 VSUBS 0.0119f
C267 VDD.n192 VSUBS 0.00922f
C268 VDD.n193 VSUBS 0.0119f
C269 VDD.n195 VSUBS 0.00747f
C270 VDD.n196 VSUBS 0.00899f
C271 VDD.n197 VSUBS 0.0111f
C272 VDD.n198 VSUBS 0.0149f
C273 VDD.n199 VSUBS 0.00922f
C274 VDD.n200 VSUBS 0.0119f
C275 VDD.n201 VSUBS 0.00922f
C276 VDD.n202 VSUBS 0.0119f
C277 VDD.n203 VSUBS 0.00922f
C278 VDD.n204 VSUBS 0.0119f
C279 VDD.n205 VSUBS 0.00922f
C280 VDD.n206 VSUBS 0.0119f
C281 VDD.n207 VSUBS 0.00922f
C282 VDD.n208 VSUBS 0.0119f
C283 VDD.n209 VSUBS 0.00922f
C284 VDD.n210 VSUBS 0.0119f
C285 VDD.n211 VSUBS 0.00922f
C286 VDD.n212 VSUBS 0.0119f
C287 VDD.n213 VSUBS 0.00922f
C288 VDD.n214 VSUBS 0.00614f
C289 VDD.n215 VSUBS 0.0247f
C290 VDD.n216 VSUBS 0.00922f
C291 VDD.n217 VSUBS 0.0117f
C292 VDD.n218 VSUBS 0.00922f
C293 VDD.n219 VSUBS 0.0119f
C294 VDD.n220 VSUBS 0.00922f
C295 VDD.n221 VSUBS 0.0119f
C296 VDD.n222 VSUBS 0.00922f
C297 VDD.n223 VSUBS 0.00968f
C298 VDD.t29 VSUBS 0.0201f
C299 VDD.n224 VSUBS 0.0201f
C300 VDD.n225 VSUBS 0.0403f
C301 VDD.n226 VSUBS 0.0435f
C302 VDD.n227 VSUBS 0.0247f
C303 VDD.n228 VSUBS 0.00922f
C304 VDD.n229 VSUBS 0.00816f
C305 VDD.n230 VSUBS 0.00922f
C306 VDD.n231 VSUBS 0.0119f
C307 VDD.n232 VSUBS 0.00922f
C308 VDD.n233 VSUBS 0.0119f
C309 VDD.n234 VSUBS 0.00922f
C310 VDD.n235 VSUBS 0.0119f
C311 VDD.n236 VSUBS 0.00922f
C312 VDD.n237 VSUBS 0.0119f
C313 VDD.n238 VSUBS 0.00922f
C314 VDD.n239 VSUBS 0.0124f
C315 VDD.n240 VSUBS 0.00922f
C316 VDD.n241 VSUBS 0.0643f
C317 VDD.n242 VSUBS 0.00922f
C318 VDD.n243 VSUBS 0.0439f
C319 VDD.n244 VSUBS 0.0111f
C320 VDD.n245 VSUBS 0.0103f
C321 VDD.n247 VSUBS 0.00747f
C322 VDD.n248 VSUBS -0.0306f
C323 VDD.n249 VSUBS 0.00922f
C324 VDD.n250 VSUBS 0.0119f
C325 VDD.n252 VSUBS 0.00922f
C326 VDD.n253 VSUBS 0.0119f
C327 VDD.n255 VSUBS 0.00922f
C328 VDD.n256 VSUBS 0.0119f
C329 VDD.n258 VSUBS 0.00922f
C330 VDD.n259 VSUBS 0.0119f
C331 VDD.n261 VSUBS 0.00922f
C332 VDD.n262 VSUBS 0.0119f
C333 VDD.n264 VSUBS 0.00922f
C334 VDD.n265 VSUBS -0.0342f
C335 VDD.n267 VSUBS 0.00922f
C336 VDD.n268 VSUBS 0.0109f
C337 VDD.n270 VSUBS 0.00922f
C338 VDD.n271 VSUBS 0.0119f
C339 VDD.n273 VSUBS 0.00922f
C340 VDD.n274 VSUBS 0.0119f
C341 VDD.n276 VSUBS 0.00922f
C342 VDD.n277 VSUBS 0.0119f
C343 VDD.n279 VSUBS 0.00922f
C344 VDD.n280 VSUBS 0.0119f
C345 VDD.n282 VSUBS 0.00922f
C346 VDD.n283 VSUBS -0.00412f
C347 VDD.n285 VSUBS 0.00922f
C348 VDD.n286 VSUBS -0.0191f
C349 VDD.n288 VSUBS 0.00922f
C350 VDD.n289 VSUBS 0.0119f
C351 VDD.n291 VSUBS 0.00922f
C352 VDD.n292 VSUBS 0.0119f
C353 VDD.n294 VSUBS 0.00922f
C354 VDD.n295 VSUBS 0.0119f
C355 VDD.n297 VSUBS 0.00922f
C356 VDD.n298 VSUBS 0.0119f
C357 VDD.n300 VSUBS 0.00922f
C358 VDD.n301 VSUBS 0.0119f
C359 VDD.n303 VSUBS 0.00922f
C360 VDD.n304 VSUBS 0.00288f
C361 VDD.n306 VSUBS 0.00922f
C362 VDD.n307 VSUBS -0.0261f
C363 VDD.n309 VSUBS 0.00922f
C364 VDD.n310 VSUBS 0.0119f
C365 VDD.n312 VSUBS 0.00922f
C366 VDD.n313 VSUBS 0.0119f
C367 VDD.n315 VSUBS 0.00922f
C368 VDD.n316 VSUBS 0.0119f
C369 VDD.n318 VSUBS 0.00922f
C370 VDD.n319 VSUBS 0.0119f
C371 VDD.n321 VSUBS 0.00922f
C372 VDD.n322 VSUBS 0.0119f
C373 VDD.n324 VSUBS 0.00922f
C374 VDD.n325 VSUBS 0.0119f
C375 VDD.n327 VSUBS 0.00922f
C376 VDD.n328 VSUBS 0.0119f
C377 VDD.n331 VSUBS 0.00922f
C378 VDD.n332 VSUBS 0.00702f
C379 VDD.n333 VSUBS 0.0222f
.ends

