* NGSPICE file created from nand_5_mag_flat.ext - technology: gf180mcuC

.subckt nand_5_mag_flat VSS A C B D E OUT VDD
X0 and_5_mag_0.and2_mag_3.IN2 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t20 VDD.t19 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 VDD E.t0 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2 OUT GF_INV_MAG_0.IN VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3 and_5_mag_0.and2_mag_1.IN2 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t26 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_2.IN2 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X5 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t8 VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_1.IN2 VDD.t24 VDD.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN A.t0 a_352_340# VSS.t14 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X8 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN B.t0 VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X9 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN E.t1 a_3213_335# VSS.t7 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X10 a_2249_324# and_5_mag_0.and2_mag_2.IN2 VSS.t16 VSS.t15 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X11 and_5_mag_0.and2_mag_3.IN2 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t13 VSS.t12 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X12 OUT GF_INV_MAG_0.IN VSS.t3 VSS.t2 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X13 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t5 VSS.t4 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X14 a_1298_335# and_5_mag_0.and2_mag_1.IN2 VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X15 VDD D.t0 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t9 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X16 GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t16 VDD.t15 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X17 VDD C.t0 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t27 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X18 VDD A.t1 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t12 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X19 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.IN2 VDD.t18 VDD.t17 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 and_5_mag_0.and2_mag_1.IN2 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t20 VSS.t19 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X21 a_352_340# B.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X22 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN D.t1 a_2249_324# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X23 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN C.t1 a_1298_335# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X24 GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t9 VSS.t8 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X25 a_3213_335# and_5_mag_0.and2_mag_3.IN2 VSS.t11 VSS.t10 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
R0 VDD.n10 VDD.t23 13882.6
R1 VDD.n7 VDD.t21 12382.6
R2 VDD.n4 VDD.t17 7208.33
R3 VDD.t15 VDD.n0 848.615
R4 VDD.t4 VDD.n1 809.492
R5 VDD VDD.n10 451.327
R6 VDD VDD.n7 445.577
R7 VDD VDD.n4 431.3
R8 VDD.t9 VDD.n4 378.788
R9 VDD.t27 VDD.n7 378.788
R10 VDD.t12 VDD.n10 378.788
R11 VDD.n3 VDD.t4 193.183
R12 VDD.n6 VDD.t9 193.183
R13 VDD.n9 VDD.t27 193.183
R14 VDD.n12 VDD.t12 193.183
R15 VDD.t17 VDD.n3 109.849
R16 VDD.t21 VDD.n6 109.849
R17 VDD.t23 VDD.n9 109.849
R18 VDD.n12 VDD.t2 109.849
R19 VDD.n10 VDD.t25 62.8277
R20 VDD.n7 VDD.t7 62.016
R21 VDD.n4 VDD.t19 60.0005
R22 VDD.n13 VDD.n12 6.3005
R23 VDD.n17 VDD.n9 6.3005
R24 VDD.n21 VDD.n6 6.3005
R25 VDD.n25 VDD.n3 6.3005
R26 VDD VDD.n0 6.3005
R27 VDD VDD.n1 6.3005
R28 VDD VDD.t3 5.1878
R29 VDD.n14 VDD.n11 5.13287
R30 VDD.n16 VDD.t24 5.13287
R31 VDD.n18 VDD.n8 5.13287
R32 VDD.n20 VDD.t22 5.13287
R33 VDD.n22 VDD.n5 5.13287
R34 VDD.n24 VDD.t18 5.13287
R35 VDD.n26 VDD.n2 5.13287
R36 VDD.n15 VDD.t26 5.09407
R37 VDD.n19 VDD.t8 5.09407
R38 VDD.n23 VDD.t20 5.09407
R39 VDD.n27 VDD.t16 5.09407
R40 VDD.n28 VDD.t1 5.09407
R41 VDD.n0 VDD.t0 4.26489
R42 VDD.n1 VDD.t15 4.26489
R43 VDD.n24 VDD 0.126036
R44 VDD.n28 VDD 0.125632
R45 VDD.n20 VDD 0.12226
R46 VDD.n16 VDD 0.11887
R47 VDD.n15 VDD.n14 0.0984239
R48 VDD.n19 VDD.n18 0.0962255
R49 VDD.n27 VDD.n26 0.0962255
R50 VDD.n23 VDD.n22 0.0917202
R51 VDD.n14 VDD.n13 0.0782465
R52 VDD.n18 VDD.n17 0.0764633
R53 VDD.n26 VDD.n25 0.0764633
R54 VDD.n22 VDD.n21 0.0728144
R55 VDD VDD.n16 0.0541697
R56 VDD VDD.n24 0.0541697
R57 VDD VDD.n20 0.0515917
R58 VDD VDD.n15 0.0339978
R59 VDD VDD.n19 0.0332632
R60 VDD VDD.n27 0.0332632
R61 VDD VDD.n23 0.0317552
R62 VDD VDD.n28 0.00839474
R63 VDD.n13 VDD 0.00388028
R64 VDD.n17 VDD 0.00380275
R65 VDD.n25 VDD 0.00380275
R66 VDD.n21 VDD 0.0036441
R67 E.n0 E.t1 31.528
R68 E.n0 E.t0 15.3826
R69 E.n1 E.n0 7.622
R70 E.n2 E.n1 5.05815
R71 E.n2 E 2.25844
R72 E.n1 E 0.0323803
R73 E E.n2 0.0095
R74 OUT.n2 OUT.n1 9.33985
R75 OUT.n2 OUT.n0 5.17836
R76 OUT OUT.n2 0.115328
R77 A.n0 A.t0 31.528
R78 A.n0 A.t1 15.3826
R79 A.n1 A.n0 7.63442
R80 A.n2 A 2.26567
R81 A.n2 A.n1 1.48351
R82 A.n1 A 0.0831009
R83 A A.n2 0.00322727
R84 VSS.t12 VSS.t10 2176.12
R85 VSS.t8 VSS.n0 2123.55
R86 VSS.t4 VSS.t15 2106.05
R87 VSS.t19 VSS.t17 2050.89
R88 VSS.n4 VSS.t21 527.028
R89 VSS.n6 VSS.t6 517.413
R90 VSS.n2 VSS.t7 517.413
R91 VSS.n8 VSS.t14 513.159
R92 VSS.t15 VSS.n4 351.351
R93 VSS.t17 VSS.n6 344.942
R94 VSS.t10 VSS.n2 344.942
R95 VSS.n8 VSS.t0 342.106
R96 VSS.n3 VSS.t12 32.9397
R97 VSS.n5 VSS.t4 32.3388
R98 VSS.n0 VSS.t2 32.3388
R99 VSS.n1 VSS.t8 32.3388
R100 VSS.n7 VSS.t19 32.0729
R101 VSS.n10 VSS.t20 9.30652
R102 VSS.n14 VSS.t5 9.30652
R103 VSS.n18 VSS.t13 9.30652
R104 VSS.n22 VSS.t9 9.30652
R105 VSS.n24 VSS.t3 9.30652
R106 VSS VSS.t1 7.20535
R107 VSS.n12 VSS.t18 7.13989
R108 VSS.n20 VSS.t11 7.13989
R109 VSS.n16 VSS.t16 7.12156
R110 VSS.n9 VSS.n8 5.2005
R111 VSS.n11 VSS.n7 5.2005
R112 VSS.n13 VSS.n6 5.2005
R113 VSS.n15 VSS.n5 5.2005
R114 VSS.n17 VSS.n4 5.2005
R115 VSS.n19 VSS.n3 5.2005
R116 VSS.n21 VSS.n2 5.2005
R117 VSS.n23 VSS.n1 5.2005
R118 VSS.n25 VSS.n0 5.2005
R119 VSS.n18 VSS.n17 0.152216
R120 VSS.n14 VSS.n13 0.151517
R121 VSS.n22 VSS.n21 0.151517
R122 VSS.n10 VSS.n9 0.151143
R123 VSS.n20 VSS 0.100904
R124 VSS.n16 VSS 0.0940347
R125 VSS.n12 VSS 0.0799976
R126 VSS.n24 VSS 0.0777785
R127 VSS VSS.n12 0.0576233
R128 VSS VSS.n16 0.0576233
R129 VSS VSS.n20 0.0576233
R130 VSS.n19 VSS.n18 0.02025
R131 VSS.n15 VSS.n14 0.0196644
R132 VSS.n23 VSS.n22 0.0196644
R133 VSS.n11 VSS.n10 0.0194096
R134 VSS VSS.n24 0.0135645
R135 VSS.n25 VSS 0.00654839
R136 VSS.n9 VSS 0.00214384
R137 VSS.n13 VSS 0.00214384
R138 VSS.n17 VSS 0.00214384
R139 VSS.n21 VSS 0.00214384
R140 VSS VSS.n19 0.001
R141 VSS VSS.n15 0.000985175
R142 VSS VSS.n23 0.000985175
R143 VSS VSS.n25 0.000983871
R144 VSS VSS.n11 0.000978723
R145 B.n0 B.t0 30.9379
R146 B.n0 B.t1 21.6422
R147 B B.n0 4.11094
R148 D.n0 D.t1 31.528
R149 D.n0 D.t0 15.3826
R150 D.n1 D.n0 7.63656
R151 D.n2 D.n1 4.925
R152 D.n2 D 2.26759
R153 D.n1 D 0.0809204
R154 D D.n2 0.0153101
R155 C.n2 C.t1 31.528
R156 C.n2 C.t0 15.3826
R157 C.n3 C.n2 5.75592
R158 C.n6 C.n5 2.52047
R159 C.n6 C 2.26388
R160 C.n1 C.n0 2.24713
R161 C.n5 C.n4 2.24658
R162 C.n0 C 0.0565142
R163 C C.n6 0.0199595
R164 C.n4 C.n3 0.0191207
R165 C.n5 C.n1 0.0105495
C0 and_5_mag_0.and2_mag_1.IN2 D 0.0053f
C1 a_1298_335# and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 4.56e-21
C2 C VDD 0.254f
C3 a_3213_335# E 0.00479f
C4 C and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0724f
C5 C a_2249_324# 9.22e-21
C6 VDD and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.43f
C7 VDD and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.429f
C8 a_1298_335# A 3.11e-21
C9 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.23e-19
C10 C and_5_mag_0.and2_mag_3.IN2 1.05e-20
C11 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_2249_324# 1.05e-20
C12 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.119f
C13 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.IN2 1.97e-19
C14 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.IN2 0.118f
C15 GF_INV_MAG_0.IN and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 5.82e-21
C16 C D 0.713f
C17 VDD B 0.174f
C18 VDD OUT 0.154f
C19 B and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0929f
C20 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN D 0.0263f
C21 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN D 0.00164f
C22 E and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.046f
C23 and_5_mag_0.and2_mag_2.IN2 A 9.39e-21
C24 C a_352_340# 0.00632f
C25 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_352_340# 4.6e-21
C26 E A 0.287f
C27 and_5_mag_0.and2_mag_2.IN2 E 0.0512f
C28 GF_INV_MAG_0.IN E 0.0103f
C29 B D 0.00833f
C30 VDD and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.428f
C31 VDD a_2249_324# 3.14e-19
C32 B a_352_340# 0.00347f
C33 a_1298_335# and_5_mag_0.and2_mag_1.IN2 0.00347f
C34 VDD and_5_mag_0.and2_mag_3.IN2 0.384f
C35 a_2249_324# and_5_mag_0.and2_mag_3.IN2 8.97e-21
C36 VDD D 0.252f
C37 a_3213_335# and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.069f
C38 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN D 0.0126f
C39 a_2249_324# D 0.0193f
C40 and_5_mag_0.and2_mag_1.IN2 A 0.00841f
C41 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_1.IN2 5.06e-21
C42 VDD a_352_340# 3.14e-19
C43 D and_5_mag_0.and2_mag_3.IN2 0.0127f
C44 C a_1298_335# 0.00943f
C45 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_352_340# 0.069f
C46 and_5_mag_0.and2_mag_1.IN2 E 0.0502f
C47 C and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 5.23e-19
C48 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_1298_335# 0.069f
C49 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.17e-19
C50 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.8e-19
C51 a_352_340# D 0.0108f
C52 C A 0.164f
C53 C and_5_mag_0.and2_mag_2.IN2 0.0122f
C54 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN A 1.88e-19
C55 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_2.IN2 0.128f
C56 VDD a_3213_335# 3.14e-19
C57 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN GF_INV_MAG_0.IN 0.128f
C58 C E 0.176f
C59 OUT and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 3.06e-21
C60 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN E 0.0477f
C61 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN E 0.3f
C62 a_3213_335# and_5_mag_0.and2_mag_3.IN2 0.00347f
C63 B A 0.169f
C64 GF_INV_MAG_0.IN OUT 0.122f
C65 VDD a_1298_335# 3.14e-19
C66 a_3213_335# D 4.35e-19
C67 a_1298_335# and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.85e-20
C68 B E 0.0106f
C69 VDD and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.429f
C70 E OUT 8.28e-19
C71 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1.9e-21
C72 a_2249_324# and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C73 C and_5_mag_0.and2_mag_1.IN2 0.101f
C74 VDD A 0.257f
C75 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.IN2 0.127f
C76 VDD and_5_mag_0.and2_mag_2.IN2 0.388f
C77 a_1298_335# D 0.0114f
C78 VDD GF_INV_MAG_0.IN 0.407f
C79 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN A 0.298f
C80 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.34e-21
C81 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_1.IN2 0.12f
C82 and_5_mag_0.and2_mag_2.IN2 a_2249_324# 0.00347f
C83 D and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.314f
C84 VDD E 0.974f
C85 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_3.IN2 4.92e-21
C86 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN E 0.0441f
C87 a_2249_324# E 7.37e-19
C88 A D 0.00372f
C89 and_5_mag_0.and2_mag_2.IN2 D 0.0782f
C90 GF_INV_MAG_0.IN D 3.08e-19
C91 E and_5_mag_0.and2_mag_3.IN2 0.101f
C92 A a_352_340# 0.00353f
C93 E D 0.143f
C94 C and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.318f
C95 VDD and_5_mag_0.and2_mag_1.IN2 0.387f
C96 C B 0.15f
C97 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_1.IN2 0.129f
C98 a_3213_335# and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.67e-20
C99 a_3213_335# VSS 0.073f
C100 a_2249_324# VSS 0.0757f
C101 a_1298_335# VSS 0.073f
C102 OUT VSS 0.204f
C103 a_352_340# VSS 0.072f
C104 GF_INV_MAG_0.IN VSS 0.418f
C105 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.446f
C106 E VSS 0.867f
C107 and_5_mag_0.and2_mag_3.IN2 VSS 0.401f
C108 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.451f
C109 D VSS 1.22f
C110 and_5_mag_0.and2_mag_2.IN2 VSS 0.399f
C111 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.446f
C112 C VSS 0.372f
C113 and_5_mag_0.and2_mag_1.IN2 VSS 0.396f
C114 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.45f
C115 A VSS 0.276f
C116 B VSS 0.337f
C117 VDD VSS 7.42f
.ends

