* NGSPICE file created from and2_mag_flat.ext - technology: gf180mcuC

.subckt and2_mag_flat IN2 IN1 OUT VDD VSS
X0 GF_INV_MAG_0.IN IN1.t0 a_168_68# VSS.t4 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1 GF_INV_MAG_0.IN IN2.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 OUT GF_INV_MAG_0.IN VSS.t3 VSS.t2 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3 a_168_68# IN2.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X4 VDD IN1.t1 GF_INV_MAG_0.IN VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X5 OUT GF_INV_MAG_0.IN VDD.t3 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 IN1.n0 IN1.t0 31.528
R1 IN1.n0 IN1.t1 15.3826
R2 IN1 IN1.n0 8.83438
R3 VSS.n4 VSS.t4 596.558
R4 VSS.n4 VSS.t0 397.707
R5 VSS.n0 VSS.t2 37.2854
R6 VSS.n2 VSS.t3 9.30652
R7 VSS VSS.t1 7.30633
R8 VSS.n1 VSS.n0 5.2005
R9 VSS.n6 VSS.n5 2.6005
R10 VSS.n5 VSS.n4 2.6005
R11 VSS.n6 VSS.n2 0.396455
R12 VSS.n5 VSS.n3 0.368921
R13 VSS.n2 VSS.n1 0.0675755
R14 VSS VSS.n6 0.00380275
R15 VSS.n1 VSS 0.00219811
R16 IN2.n0 IN2.t0 30.9379
R17 IN2.n0 IN2.t1 21.6422
R18 IN2 IN2.n0 4.11094
R19 VDD.n4 VDD 425.019
R20 VDD.t4 VDD.n4 378.788
R21 VDD.n5 VDD.t4 193.183
R22 VDD.n5 VDD.t0 109.849
R23 VDD.n4 VDD.t2 59.1138
R24 VDD VDD.t1 5.20835
R25 VDD.n1 VDD.n0 5.13287
R26 VDD.n3 VDD.t3 5.09407
R27 VDD.n7 VDD.n6 3.1505
R28 VDD.n6 VDD.n5 3.1505
R29 VDD.n3 VDD.n1 0.170231
R30 VDD.n6 VDD.n2 0.160669
R31 VDD.n7 VDD.n1 0.107339
R32 VDD VDD.n3 0.0709717
R33 VDD VDD.n7 0.00514516
R34 OUT.n2 OUT.n1 9.33985
R35 OUT.n2 OUT.n0 5.17836
R36 OUT OUT.n2 0.0594655
C0 GF_INV_MAG_0.IN IN2 0.0929f
C1 GF_INV_MAG_0.IN OUT 0.116f
C2 VDD IN1 0.229f
C3 a_168_68# IN2 0.00347f
C4 GF_INV_MAG_0.IN IN1 0.251f
C5 GF_INV_MAG_0.IN VDD 0.42f
C6 a_168_68# IN1 0.00348f
C7 VDD a_168_68# 3.14e-19
C8 IN2 IN1 0.0466f
C9 OUT IN1 0.00639f
C10 VDD IN2 0.158f
C11 VDD OUT 0.154f
C12 GF_INV_MAG_0.IN a_168_68# 0.069f
C13 IN1 VSS 0.218f
C14 IN2 VSS 0.307f
C15 a_168_68# VSS 0.0678f
C16 OUT VSS 0.175f
C17 GF_INV_MAG_0.IN VSS 0.48f
C18 VDD VSS 1.74f
.ends

