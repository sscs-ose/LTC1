magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -4649 -2975 4649 2975
<< psubdiff >>
rect -2649 953 2649 975
rect -2649 907 -2627 953
rect -2581 907 -2503 953
rect -2457 907 -2379 953
rect -2333 907 -2255 953
rect -2209 907 -2131 953
rect -2085 907 -2007 953
rect -1961 907 -1883 953
rect -1837 907 -1759 953
rect -1713 907 -1635 953
rect -1589 907 -1511 953
rect -1465 907 -1387 953
rect -1341 907 -1263 953
rect -1217 907 -1139 953
rect -1093 907 -1015 953
rect -969 907 -891 953
rect -845 907 -767 953
rect -721 907 -643 953
rect -597 907 -519 953
rect -473 907 -395 953
rect -349 907 -271 953
rect -225 907 -147 953
rect -101 907 -23 953
rect 23 907 101 953
rect 147 907 225 953
rect 271 907 349 953
rect 395 907 473 953
rect 519 907 597 953
rect 643 907 721 953
rect 767 907 845 953
rect 891 907 969 953
rect 1015 907 1093 953
rect 1139 907 1217 953
rect 1263 907 1341 953
rect 1387 907 1465 953
rect 1511 907 1589 953
rect 1635 907 1713 953
rect 1759 907 1837 953
rect 1883 907 1961 953
rect 2007 907 2085 953
rect 2131 907 2209 953
rect 2255 907 2333 953
rect 2379 907 2457 953
rect 2503 907 2581 953
rect 2627 907 2649 953
rect -2649 829 2649 907
rect -2649 783 -2627 829
rect -2581 783 -2503 829
rect -2457 783 -2379 829
rect -2333 783 -2255 829
rect -2209 783 -2131 829
rect -2085 783 -2007 829
rect -1961 783 -1883 829
rect -1837 783 -1759 829
rect -1713 783 -1635 829
rect -1589 783 -1511 829
rect -1465 783 -1387 829
rect -1341 783 -1263 829
rect -1217 783 -1139 829
rect -1093 783 -1015 829
rect -969 783 -891 829
rect -845 783 -767 829
rect -721 783 -643 829
rect -597 783 -519 829
rect -473 783 -395 829
rect -349 783 -271 829
rect -225 783 -147 829
rect -101 783 -23 829
rect 23 783 101 829
rect 147 783 225 829
rect 271 783 349 829
rect 395 783 473 829
rect 519 783 597 829
rect 643 783 721 829
rect 767 783 845 829
rect 891 783 969 829
rect 1015 783 1093 829
rect 1139 783 1217 829
rect 1263 783 1341 829
rect 1387 783 1465 829
rect 1511 783 1589 829
rect 1635 783 1713 829
rect 1759 783 1837 829
rect 1883 783 1961 829
rect 2007 783 2085 829
rect 2131 783 2209 829
rect 2255 783 2333 829
rect 2379 783 2457 829
rect 2503 783 2581 829
rect 2627 783 2649 829
rect -2649 705 2649 783
rect -2649 659 -2627 705
rect -2581 659 -2503 705
rect -2457 659 -2379 705
rect -2333 659 -2255 705
rect -2209 659 -2131 705
rect -2085 659 -2007 705
rect -1961 659 -1883 705
rect -1837 659 -1759 705
rect -1713 659 -1635 705
rect -1589 659 -1511 705
rect -1465 659 -1387 705
rect -1341 659 -1263 705
rect -1217 659 -1139 705
rect -1093 659 -1015 705
rect -969 659 -891 705
rect -845 659 -767 705
rect -721 659 -643 705
rect -597 659 -519 705
rect -473 659 -395 705
rect -349 659 -271 705
rect -225 659 -147 705
rect -101 659 -23 705
rect 23 659 101 705
rect 147 659 225 705
rect 271 659 349 705
rect 395 659 473 705
rect 519 659 597 705
rect 643 659 721 705
rect 767 659 845 705
rect 891 659 969 705
rect 1015 659 1093 705
rect 1139 659 1217 705
rect 1263 659 1341 705
rect 1387 659 1465 705
rect 1511 659 1589 705
rect 1635 659 1713 705
rect 1759 659 1837 705
rect 1883 659 1961 705
rect 2007 659 2085 705
rect 2131 659 2209 705
rect 2255 659 2333 705
rect 2379 659 2457 705
rect 2503 659 2581 705
rect 2627 659 2649 705
rect -2649 581 2649 659
rect -2649 535 -2627 581
rect -2581 535 -2503 581
rect -2457 535 -2379 581
rect -2333 535 -2255 581
rect -2209 535 -2131 581
rect -2085 535 -2007 581
rect -1961 535 -1883 581
rect -1837 535 -1759 581
rect -1713 535 -1635 581
rect -1589 535 -1511 581
rect -1465 535 -1387 581
rect -1341 535 -1263 581
rect -1217 535 -1139 581
rect -1093 535 -1015 581
rect -969 535 -891 581
rect -845 535 -767 581
rect -721 535 -643 581
rect -597 535 -519 581
rect -473 535 -395 581
rect -349 535 -271 581
rect -225 535 -147 581
rect -101 535 -23 581
rect 23 535 101 581
rect 147 535 225 581
rect 271 535 349 581
rect 395 535 473 581
rect 519 535 597 581
rect 643 535 721 581
rect 767 535 845 581
rect 891 535 969 581
rect 1015 535 1093 581
rect 1139 535 1217 581
rect 1263 535 1341 581
rect 1387 535 1465 581
rect 1511 535 1589 581
rect 1635 535 1713 581
rect 1759 535 1837 581
rect 1883 535 1961 581
rect 2007 535 2085 581
rect 2131 535 2209 581
rect 2255 535 2333 581
rect 2379 535 2457 581
rect 2503 535 2581 581
rect 2627 535 2649 581
rect -2649 457 2649 535
rect -2649 411 -2627 457
rect -2581 411 -2503 457
rect -2457 411 -2379 457
rect -2333 411 -2255 457
rect -2209 411 -2131 457
rect -2085 411 -2007 457
rect -1961 411 -1883 457
rect -1837 411 -1759 457
rect -1713 411 -1635 457
rect -1589 411 -1511 457
rect -1465 411 -1387 457
rect -1341 411 -1263 457
rect -1217 411 -1139 457
rect -1093 411 -1015 457
rect -969 411 -891 457
rect -845 411 -767 457
rect -721 411 -643 457
rect -597 411 -519 457
rect -473 411 -395 457
rect -349 411 -271 457
rect -225 411 -147 457
rect -101 411 -23 457
rect 23 411 101 457
rect 147 411 225 457
rect 271 411 349 457
rect 395 411 473 457
rect 519 411 597 457
rect 643 411 721 457
rect 767 411 845 457
rect 891 411 969 457
rect 1015 411 1093 457
rect 1139 411 1217 457
rect 1263 411 1341 457
rect 1387 411 1465 457
rect 1511 411 1589 457
rect 1635 411 1713 457
rect 1759 411 1837 457
rect 1883 411 1961 457
rect 2007 411 2085 457
rect 2131 411 2209 457
rect 2255 411 2333 457
rect 2379 411 2457 457
rect 2503 411 2581 457
rect 2627 411 2649 457
rect -2649 333 2649 411
rect -2649 287 -2627 333
rect -2581 287 -2503 333
rect -2457 287 -2379 333
rect -2333 287 -2255 333
rect -2209 287 -2131 333
rect -2085 287 -2007 333
rect -1961 287 -1883 333
rect -1837 287 -1759 333
rect -1713 287 -1635 333
rect -1589 287 -1511 333
rect -1465 287 -1387 333
rect -1341 287 -1263 333
rect -1217 287 -1139 333
rect -1093 287 -1015 333
rect -969 287 -891 333
rect -845 287 -767 333
rect -721 287 -643 333
rect -597 287 -519 333
rect -473 287 -395 333
rect -349 287 -271 333
rect -225 287 -147 333
rect -101 287 -23 333
rect 23 287 101 333
rect 147 287 225 333
rect 271 287 349 333
rect 395 287 473 333
rect 519 287 597 333
rect 643 287 721 333
rect 767 287 845 333
rect 891 287 969 333
rect 1015 287 1093 333
rect 1139 287 1217 333
rect 1263 287 1341 333
rect 1387 287 1465 333
rect 1511 287 1589 333
rect 1635 287 1713 333
rect 1759 287 1837 333
rect 1883 287 1961 333
rect 2007 287 2085 333
rect 2131 287 2209 333
rect 2255 287 2333 333
rect 2379 287 2457 333
rect 2503 287 2581 333
rect 2627 287 2649 333
rect -2649 209 2649 287
rect -2649 163 -2627 209
rect -2581 163 -2503 209
rect -2457 163 -2379 209
rect -2333 163 -2255 209
rect -2209 163 -2131 209
rect -2085 163 -2007 209
rect -1961 163 -1883 209
rect -1837 163 -1759 209
rect -1713 163 -1635 209
rect -1589 163 -1511 209
rect -1465 163 -1387 209
rect -1341 163 -1263 209
rect -1217 163 -1139 209
rect -1093 163 -1015 209
rect -969 163 -891 209
rect -845 163 -767 209
rect -721 163 -643 209
rect -597 163 -519 209
rect -473 163 -395 209
rect -349 163 -271 209
rect -225 163 -147 209
rect -101 163 -23 209
rect 23 163 101 209
rect 147 163 225 209
rect 271 163 349 209
rect 395 163 473 209
rect 519 163 597 209
rect 643 163 721 209
rect 767 163 845 209
rect 891 163 969 209
rect 1015 163 1093 209
rect 1139 163 1217 209
rect 1263 163 1341 209
rect 1387 163 1465 209
rect 1511 163 1589 209
rect 1635 163 1713 209
rect 1759 163 1837 209
rect 1883 163 1961 209
rect 2007 163 2085 209
rect 2131 163 2209 209
rect 2255 163 2333 209
rect 2379 163 2457 209
rect 2503 163 2581 209
rect 2627 163 2649 209
rect -2649 85 2649 163
rect -2649 39 -2627 85
rect -2581 39 -2503 85
rect -2457 39 -2379 85
rect -2333 39 -2255 85
rect -2209 39 -2131 85
rect -2085 39 -2007 85
rect -1961 39 -1883 85
rect -1837 39 -1759 85
rect -1713 39 -1635 85
rect -1589 39 -1511 85
rect -1465 39 -1387 85
rect -1341 39 -1263 85
rect -1217 39 -1139 85
rect -1093 39 -1015 85
rect -969 39 -891 85
rect -845 39 -767 85
rect -721 39 -643 85
rect -597 39 -519 85
rect -473 39 -395 85
rect -349 39 -271 85
rect -225 39 -147 85
rect -101 39 -23 85
rect 23 39 101 85
rect 147 39 225 85
rect 271 39 349 85
rect 395 39 473 85
rect 519 39 597 85
rect 643 39 721 85
rect 767 39 845 85
rect 891 39 969 85
rect 1015 39 1093 85
rect 1139 39 1217 85
rect 1263 39 1341 85
rect 1387 39 1465 85
rect 1511 39 1589 85
rect 1635 39 1713 85
rect 1759 39 1837 85
rect 1883 39 1961 85
rect 2007 39 2085 85
rect 2131 39 2209 85
rect 2255 39 2333 85
rect 2379 39 2457 85
rect 2503 39 2581 85
rect 2627 39 2649 85
rect -2649 -39 2649 39
rect -2649 -85 -2627 -39
rect -2581 -85 -2503 -39
rect -2457 -85 -2379 -39
rect -2333 -85 -2255 -39
rect -2209 -85 -2131 -39
rect -2085 -85 -2007 -39
rect -1961 -85 -1883 -39
rect -1837 -85 -1759 -39
rect -1713 -85 -1635 -39
rect -1589 -85 -1511 -39
rect -1465 -85 -1387 -39
rect -1341 -85 -1263 -39
rect -1217 -85 -1139 -39
rect -1093 -85 -1015 -39
rect -969 -85 -891 -39
rect -845 -85 -767 -39
rect -721 -85 -643 -39
rect -597 -85 -519 -39
rect -473 -85 -395 -39
rect -349 -85 -271 -39
rect -225 -85 -147 -39
rect -101 -85 -23 -39
rect 23 -85 101 -39
rect 147 -85 225 -39
rect 271 -85 349 -39
rect 395 -85 473 -39
rect 519 -85 597 -39
rect 643 -85 721 -39
rect 767 -85 845 -39
rect 891 -85 969 -39
rect 1015 -85 1093 -39
rect 1139 -85 1217 -39
rect 1263 -85 1341 -39
rect 1387 -85 1465 -39
rect 1511 -85 1589 -39
rect 1635 -85 1713 -39
rect 1759 -85 1837 -39
rect 1883 -85 1961 -39
rect 2007 -85 2085 -39
rect 2131 -85 2209 -39
rect 2255 -85 2333 -39
rect 2379 -85 2457 -39
rect 2503 -85 2581 -39
rect 2627 -85 2649 -39
rect -2649 -163 2649 -85
rect -2649 -209 -2627 -163
rect -2581 -209 -2503 -163
rect -2457 -209 -2379 -163
rect -2333 -209 -2255 -163
rect -2209 -209 -2131 -163
rect -2085 -209 -2007 -163
rect -1961 -209 -1883 -163
rect -1837 -209 -1759 -163
rect -1713 -209 -1635 -163
rect -1589 -209 -1511 -163
rect -1465 -209 -1387 -163
rect -1341 -209 -1263 -163
rect -1217 -209 -1139 -163
rect -1093 -209 -1015 -163
rect -969 -209 -891 -163
rect -845 -209 -767 -163
rect -721 -209 -643 -163
rect -597 -209 -519 -163
rect -473 -209 -395 -163
rect -349 -209 -271 -163
rect -225 -209 -147 -163
rect -101 -209 -23 -163
rect 23 -209 101 -163
rect 147 -209 225 -163
rect 271 -209 349 -163
rect 395 -209 473 -163
rect 519 -209 597 -163
rect 643 -209 721 -163
rect 767 -209 845 -163
rect 891 -209 969 -163
rect 1015 -209 1093 -163
rect 1139 -209 1217 -163
rect 1263 -209 1341 -163
rect 1387 -209 1465 -163
rect 1511 -209 1589 -163
rect 1635 -209 1713 -163
rect 1759 -209 1837 -163
rect 1883 -209 1961 -163
rect 2007 -209 2085 -163
rect 2131 -209 2209 -163
rect 2255 -209 2333 -163
rect 2379 -209 2457 -163
rect 2503 -209 2581 -163
rect 2627 -209 2649 -163
rect -2649 -287 2649 -209
rect -2649 -333 -2627 -287
rect -2581 -333 -2503 -287
rect -2457 -333 -2379 -287
rect -2333 -333 -2255 -287
rect -2209 -333 -2131 -287
rect -2085 -333 -2007 -287
rect -1961 -333 -1883 -287
rect -1837 -333 -1759 -287
rect -1713 -333 -1635 -287
rect -1589 -333 -1511 -287
rect -1465 -333 -1387 -287
rect -1341 -333 -1263 -287
rect -1217 -333 -1139 -287
rect -1093 -333 -1015 -287
rect -969 -333 -891 -287
rect -845 -333 -767 -287
rect -721 -333 -643 -287
rect -597 -333 -519 -287
rect -473 -333 -395 -287
rect -349 -333 -271 -287
rect -225 -333 -147 -287
rect -101 -333 -23 -287
rect 23 -333 101 -287
rect 147 -333 225 -287
rect 271 -333 349 -287
rect 395 -333 473 -287
rect 519 -333 597 -287
rect 643 -333 721 -287
rect 767 -333 845 -287
rect 891 -333 969 -287
rect 1015 -333 1093 -287
rect 1139 -333 1217 -287
rect 1263 -333 1341 -287
rect 1387 -333 1465 -287
rect 1511 -333 1589 -287
rect 1635 -333 1713 -287
rect 1759 -333 1837 -287
rect 1883 -333 1961 -287
rect 2007 -333 2085 -287
rect 2131 -333 2209 -287
rect 2255 -333 2333 -287
rect 2379 -333 2457 -287
rect 2503 -333 2581 -287
rect 2627 -333 2649 -287
rect -2649 -411 2649 -333
rect -2649 -457 -2627 -411
rect -2581 -457 -2503 -411
rect -2457 -457 -2379 -411
rect -2333 -457 -2255 -411
rect -2209 -457 -2131 -411
rect -2085 -457 -2007 -411
rect -1961 -457 -1883 -411
rect -1837 -457 -1759 -411
rect -1713 -457 -1635 -411
rect -1589 -457 -1511 -411
rect -1465 -457 -1387 -411
rect -1341 -457 -1263 -411
rect -1217 -457 -1139 -411
rect -1093 -457 -1015 -411
rect -969 -457 -891 -411
rect -845 -457 -767 -411
rect -721 -457 -643 -411
rect -597 -457 -519 -411
rect -473 -457 -395 -411
rect -349 -457 -271 -411
rect -225 -457 -147 -411
rect -101 -457 -23 -411
rect 23 -457 101 -411
rect 147 -457 225 -411
rect 271 -457 349 -411
rect 395 -457 473 -411
rect 519 -457 597 -411
rect 643 -457 721 -411
rect 767 -457 845 -411
rect 891 -457 969 -411
rect 1015 -457 1093 -411
rect 1139 -457 1217 -411
rect 1263 -457 1341 -411
rect 1387 -457 1465 -411
rect 1511 -457 1589 -411
rect 1635 -457 1713 -411
rect 1759 -457 1837 -411
rect 1883 -457 1961 -411
rect 2007 -457 2085 -411
rect 2131 -457 2209 -411
rect 2255 -457 2333 -411
rect 2379 -457 2457 -411
rect 2503 -457 2581 -411
rect 2627 -457 2649 -411
rect -2649 -535 2649 -457
rect -2649 -581 -2627 -535
rect -2581 -581 -2503 -535
rect -2457 -581 -2379 -535
rect -2333 -581 -2255 -535
rect -2209 -581 -2131 -535
rect -2085 -581 -2007 -535
rect -1961 -581 -1883 -535
rect -1837 -581 -1759 -535
rect -1713 -581 -1635 -535
rect -1589 -581 -1511 -535
rect -1465 -581 -1387 -535
rect -1341 -581 -1263 -535
rect -1217 -581 -1139 -535
rect -1093 -581 -1015 -535
rect -969 -581 -891 -535
rect -845 -581 -767 -535
rect -721 -581 -643 -535
rect -597 -581 -519 -535
rect -473 -581 -395 -535
rect -349 -581 -271 -535
rect -225 -581 -147 -535
rect -101 -581 -23 -535
rect 23 -581 101 -535
rect 147 -581 225 -535
rect 271 -581 349 -535
rect 395 -581 473 -535
rect 519 -581 597 -535
rect 643 -581 721 -535
rect 767 -581 845 -535
rect 891 -581 969 -535
rect 1015 -581 1093 -535
rect 1139 -581 1217 -535
rect 1263 -581 1341 -535
rect 1387 -581 1465 -535
rect 1511 -581 1589 -535
rect 1635 -581 1713 -535
rect 1759 -581 1837 -535
rect 1883 -581 1961 -535
rect 2007 -581 2085 -535
rect 2131 -581 2209 -535
rect 2255 -581 2333 -535
rect 2379 -581 2457 -535
rect 2503 -581 2581 -535
rect 2627 -581 2649 -535
rect -2649 -659 2649 -581
rect -2649 -705 -2627 -659
rect -2581 -705 -2503 -659
rect -2457 -705 -2379 -659
rect -2333 -705 -2255 -659
rect -2209 -705 -2131 -659
rect -2085 -705 -2007 -659
rect -1961 -705 -1883 -659
rect -1837 -705 -1759 -659
rect -1713 -705 -1635 -659
rect -1589 -705 -1511 -659
rect -1465 -705 -1387 -659
rect -1341 -705 -1263 -659
rect -1217 -705 -1139 -659
rect -1093 -705 -1015 -659
rect -969 -705 -891 -659
rect -845 -705 -767 -659
rect -721 -705 -643 -659
rect -597 -705 -519 -659
rect -473 -705 -395 -659
rect -349 -705 -271 -659
rect -225 -705 -147 -659
rect -101 -705 -23 -659
rect 23 -705 101 -659
rect 147 -705 225 -659
rect 271 -705 349 -659
rect 395 -705 473 -659
rect 519 -705 597 -659
rect 643 -705 721 -659
rect 767 -705 845 -659
rect 891 -705 969 -659
rect 1015 -705 1093 -659
rect 1139 -705 1217 -659
rect 1263 -705 1341 -659
rect 1387 -705 1465 -659
rect 1511 -705 1589 -659
rect 1635 -705 1713 -659
rect 1759 -705 1837 -659
rect 1883 -705 1961 -659
rect 2007 -705 2085 -659
rect 2131 -705 2209 -659
rect 2255 -705 2333 -659
rect 2379 -705 2457 -659
rect 2503 -705 2581 -659
rect 2627 -705 2649 -659
rect -2649 -783 2649 -705
rect -2649 -829 -2627 -783
rect -2581 -829 -2503 -783
rect -2457 -829 -2379 -783
rect -2333 -829 -2255 -783
rect -2209 -829 -2131 -783
rect -2085 -829 -2007 -783
rect -1961 -829 -1883 -783
rect -1837 -829 -1759 -783
rect -1713 -829 -1635 -783
rect -1589 -829 -1511 -783
rect -1465 -829 -1387 -783
rect -1341 -829 -1263 -783
rect -1217 -829 -1139 -783
rect -1093 -829 -1015 -783
rect -969 -829 -891 -783
rect -845 -829 -767 -783
rect -721 -829 -643 -783
rect -597 -829 -519 -783
rect -473 -829 -395 -783
rect -349 -829 -271 -783
rect -225 -829 -147 -783
rect -101 -829 -23 -783
rect 23 -829 101 -783
rect 147 -829 225 -783
rect 271 -829 349 -783
rect 395 -829 473 -783
rect 519 -829 597 -783
rect 643 -829 721 -783
rect 767 -829 845 -783
rect 891 -829 969 -783
rect 1015 -829 1093 -783
rect 1139 -829 1217 -783
rect 1263 -829 1341 -783
rect 1387 -829 1465 -783
rect 1511 -829 1589 -783
rect 1635 -829 1713 -783
rect 1759 -829 1837 -783
rect 1883 -829 1961 -783
rect 2007 -829 2085 -783
rect 2131 -829 2209 -783
rect 2255 -829 2333 -783
rect 2379 -829 2457 -783
rect 2503 -829 2581 -783
rect 2627 -829 2649 -783
rect -2649 -907 2649 -829
rect -2649 -953 -2627 -907
rect -2581 -953 -2503 -907
rect -2457 -953 -2379 -907
rect -2333 -953 -2255 -907
rect -2209 -953 -2131 -907
rect -2085 -953 -2007 -907
rect -1961 -953 -1883 -907
rect -1837 -953 -1759 -907
rect -1713 -953 -1635 -907
rect -1589 -953 -1511 -907
rect -1465 -953 -1387 -907
rect -1341 -953 -1263 -907
rect -1217 -953 -1139 -907
rect -1093 -953 -1015 -907
rect -969 -953 -891 -907
rect -845 -953 -767 -907
rect -721 -953 -643 -907
rect -597 -953 -519 -907
rect -473 -953 -395 -907
rect -349 -953 -271 -907
rect -225 -953 -147 -907
rect -101 -953 -23 -907
rect 23 -953 101 -907
rect 147 -953 225 -907
rect 271 -953 349 -907
rect 395 -953 473 -907
rect 519 -953 597 -907
rect 643 -953 721 -907
rect 767 -953 845 -907
rect 891 -953 969 -907
rect 1015 -953 1093 -907
rect 1139 -953 1217 -907
rect 1263 -953 1341 -907
rect 1387 -953 1465 -907
rect 1511 -953 1589 -907
rect 1635 -953 1713 -907
rect 1759 -953 1837 -907
rect 1883 -953 1961 -907
rect 2007 -953 2085 -907
rect 2131 -953 2209 -907
rect 2255 -953 2333 -907
rect 2379 -953 2457 -907
rect 2503 -953 2581 -907
rect 2627 -953 2649 -907
rect -2649 -975 2649 -953
<< psubdiffcont >>
rect -2627 907 -2581 953
rect -2503 907 -2457 953
rect -2379 907 -2333 953
rect -2255 907 -2209 953
rect -2131 907 -2085 953
rect -2007 907 -1961 953
rect -1883 907 -1837 953
rect -1759 907 -1713 953
rect -1635 907 -1589 953
rect -1511 907 -1465 953
rect -1387 907 -1341 953
rect -1263 907 -1217 953
rect -1139 907 -1093 953
rect -1015 907 -969 953
rect -891 907 -845 953
rect -767 907 -721 953
rect -643 907 -597 953
rect -519 907 -473 953
rect -395 907 -349 953
rect -271 907 -225 953
rect -147 907 -101 953
rect -23 907 23 953
rect 101 907 147 953
rect 225 907 271 953
rect 349 907 395 953
rect 473 907 519 953
rect 597 907 643 953
rect 721 907 767 953
rect 845 907 891 953
rect 969 907 1015 953
rect 1093 907 1139 953
rect 1217 907 1263 953
rect 1341 907 1387 953
rect 1465 907 1511 953
rect 1589 907 1635 953
rect 1713 907 1759 953
rect 1837 907 1883 953
rect 1961 907 2007 953
rect 2085 907 2131 953
rect 2209 907 2255 953
rect 2333 907 2379 953
rect 2457 907 2503 953
rect 2581 907 2627 953
rect -2627 783 -2581 829
rect -2503 783 -2457 829
rect -2379 783 -2333 829
rect -2255 783 -2209 829
rect -2131 783 -2085 829
rect -2007 783 -1961 829
rect -1883 783 -1837 829
rect -1759 783 -1713 829
rect -1635 783 -1589 829
rect -1511 783 -1465 829
rect -1387 783 -1341 829
rect -1263 783 -1217 829
rect -1139 783 -1093 829
rect -1015 783 -969 829
rect -891 783 -845 829
rect -767 783 -721 829
rect -643 783 -597 829
rect -519 783 -473 829
rect -395 783 -349 829
rect -271 783 -225 829
rect -147 783 -101 829
rect -23 783 23 829
rect 101 783 147 829
rect 225 783 271 829
rect 349 783 395 829
rect 473 783 519 829
rect 597 783 643 829
rect 721 783 767 829
rect 845 783 891 829
rect 969 783 1015 829
rect 1093 783 1139 829
rect 1217 783 1263 829
rect 1341 783 1387 829
rect 1465 783 1511 829
rect 1589 783 1635 829
rect 1713 783 1759 829
rect 1837 783 1883 829
rect 1961 783 2007 829
rect 2085 783 2131 829
rect 2209 783 2255 829
rect 2333 783 2379 829
rect 2457 783 2503 829
rect 2581 783 2627 829
rect -2627 659 -2581 705
rect -2503 659 -2457 705
rect -2379 659 -2333 705
rect -2255 659 -2209 705
rect -2131 659 -2085 705
rect -2007 659 -1961 705
rect -1883 659 -1837 705
rect -1759 659 -1713 705
rect -1635 659 -1589 705
rect -1511 659 -1465 705
rect -1387 659 -1341 705
rect -1263 659 -1217 705
rect -1139 659 -1093 705
rect -1015 659 -969 705
rect -891 659 -845 705
rect -767 659 -721 705
rect -643 659 -597 705
rect -519 659 -473 705
rect -395 659 -349 705
rect -271 659 -225 705
rect -147 659 -101 705
rect -23 659 23 705
rect 101 659 147 705
rect 225 659 271 705
rect 349 659 395 705
rect 473 659 519 705
rect 597 659 643 705
rect 721 659 767 705
rect 845 659 891 705
rect 969 659 1015 705
rect 1093 659 1139 705
rect 1217 659 1263 705
rect 1341 659 1387 705
rect 1465 659 1511 705
rect 1589 659 1635 705
rect 1713 659 1759 705
rect 1837 659 1883 705
rect 1961 659 2007 705
rect 2085 659 2131 705
rect 2209 659 2255 705
rect 2333 659 2379 705
rect 2457 659 2503 705
rect 2581 659 2627 705
rect -2627 535 -2581 581
rect -2503 535 -2457 581
rect -2379 535 -2333 581
rect -2255 535 -2209 581
rect -2131 535 -2085 581
rect -2007 535 -1961 581
rect -1883 535 -1837 581
rect -1759 535 -1713 581
rect -1635 535 -1589 581
rect -1511 535 -1465 581
rect -1387 535 -1341 581
rect -1263 535 -1217 581
rect -1139 535 -1093 581
rect -1015 535 -969 581
rect -891 535 -845 581
rect -767 535 -721 581
rect -643 535 -597 581
rect -519 535 -473 581
rect -395 535 -349 581
rect -271 535 -225 581
rect -147 535 -101 581
rect -23 535 23 581
rect 101 535 147 581
rect 225 535 271 581
rect 349 535 395 581
rect 473 535 519 581
rect 597 535 643 581
rect 721 535 767 581
rect 845 535 891 581
rect 969 535 1015 581
rect 1093 535 1139 581
rect 1217 535 1263 581
rect 1341 535 1387 581
rect 1465 535 1511 581
rect 1589 535 1635 581
rect 1713 535 1759 581
rect 1837 535 1883 581
rect 1961 535 2007 581
rect 2085 535 2131 581
rect 2209 535 2255 581
rect 2333 535 2379 581
rect 2457 535 2503 581
rect 2581 535 2627 581
rect -2627 411 -2581 457
rect -2503 411 -2457 457
rect -2379 411 -2333 457
rect -2255 411 -2209 457
rect -2131 411 -2085 457
rect -2007 411 -1961 457
rect -1883 411 -1837 457
rect -1759 411 -1713 457
rect -1635 411 -1589 457
rect -1511 411 -1465 457
rect -1387 411 -1341 457
rect -1263 411 -1217 457
rect -1139 411 -1093 457
rect -1015 411 -969 457
rect -891 411 -845 457
rect -767 411 -721 457
rect -643 411 -597 457
rect -519 411 -473 457
rect -395 411 -349 457
rect -271 411 -225 457
rect -147 411 -101 457
rect -23 411 23 457
rect 101 411 147 457
rect 225 411 271 457
rect 349 411 395 457
rect 473 411 519 457
rect 597 411 643 457
rect 721 411 767 457
rect 845 411 891 457
rect 969 411 1015 457
rect 1093 411 1139 457
rect 1217 411 1263 457
rect 1341 411 1387 457
rect 1465 411 1511 457
rect 1589 411 1635 457
rect 1713 411 1759 457
rect 1837 411 1883 457
rect 1961 411 2007 457
rect 2085 411 2131 457
rect 2209 411 2255 457
rect 2333 411 2379 457
rect 2457 411 2503 457
rect 2581 411 2627 457
rect -2627 287 -2581 333
rect -2503 287 -2457 333
rect -2379 287 -2333 333
rect -2255 287 -2209 333
rect -2131 287 -2085 333
rect -2007 287 -1961 333
rect -1883 287 -1837 333
rect -1759 287 -1713 333
rect -1635 287 -1589 333
rect -1511 287 -1465 333
rect -1387 287 -1341 333
rect -1263 287 -1217 333
rect -1139 287 -1093 333
rect -1015 287 -969 333
rect -891 287 -845 333
rect -767 287 -721 333
rect -643 287 -597 333
rect -519 287 -473 333
rect -395 287 -349 333
rect -271 287 -225 333
rect -147 287 -101 333
rect -23 287 23 333
rect 101 287 147 333
rect 225 287 271 333
rect 349 287 395 333
rect 473 287 519 333
rect 597 287 643 333
rect 721 287 767 333
rect 845 287 891 333
rect 969 287 1015 333
rect 1093 287 1139 333
rect 1217 287 1263 333
rect 1341 287 1387 333
rect 1465 287 1511 333
rect 1589 287 1635 333
rect 1713 287 1759 333
rect 1837 287 1883 333
rect 1961 287 2007 333
rect 2085 287 2131 333
rect 2209 287 2255 333
rect 2333 287 2379 333
rect 2457 287 2503 333
rect 2581 287 2627 333
rect -2627 163 -2581 209
rect -2503 163 -2457 209
rect -2379 163 -2333 209
rect -2255 163 -2209 209
rect -2131 163 -2085 209
rect -2007 163 -1961 209
rect -1883 163 -1837 209
rect -1759 163 -1713 209
rect -1635 163 -1589 209
rect -1511 163 -1465 209
rect -1387 163 -1341 209
rect -1263 163 -1217 209
rect -1139 163 -1093 209
rect -1015 163 -969 209
rect -891 163 -845 209
rect -767 163 -721 209
rect -643 163 -597 209
rect -519 163 -473 209
rect -395 163 -349 209
rect -271 163 -225 209
rect -147 163 -101 209
rect -23 163 23 209
rect 101 163 147 209
rect 225 163 271 209
rect 349 163 395 209
rect 473 163 519 209
rect 597 163 643 209
rect 721 163 767 209
rect 845 163 891 209
rect 969 163 1015 209
rect 1093 163 1139 209
rect 1217 163 1263 209
rect 1341 163 1387 209
rect 1465 163 1511 209
rect 1589 163 1635 209
rect 1713 163 1759 209
rect 1837 163 1883 209
rect 1961 163 2007 209
rect 2085 163 2131 209
rect 2209 163 2255 209
rect 2333 163 2379 209
rect 2457 163 2503 209
rect 2581 163 2627 209
rect -2627 39 -2581 85
rect -2503 39 -2457 85
rect -2379 39 -2333 85
rect -2255 39 -2209 85
rect -2131 39 -2085 85
rect -2007 39 -1961 85
rect -1883 39 -1837 85
rect -1759 39 -1713 85
rect -1635 39 -1589 85
rect -1511 39 -1465 85
rect -1387 39 -1341 85
rect -1263 39 -1217 85
rect -1139 39 -1093 85
rect -1015 39 -969 85
rect -891 39 -845 85
rect -767 39 -721 85
rect -643 39 -597 85
rect -519 39 -473 85
rect -395 39 -349 85
rect -271 39 -225 85
rect -147 39 -101 85
rect -23 39 23 85
rect 101 39 147 85
rect 225 39 271 85
rect 349 39 395 85
rect 473 39 519 85
rect 597 39 643 85
rect 721 39 767 85
rect 845 39 891 85
rect 969 39 1015 85
rect 1093 39 1139 85
rect 1217 39 1263 85
rect 1341 39 1387 85
rect 1465 39 1511 85
rect 1589 39 1635 85
rect 1713 39 1759 85
rect 1837 39 1883 85
rect 1961 39 2007 85
rect 2085 39 2131 85
rect 2209 39 2255 85
rect 2333 39 2379 85
rect 2457 39 2503 85
rect 2581 39 2627 85
rect -2627 -85 -2581 -39
rect -2503 -85 -2457 -39
rect -2379 -85 -2333 -39
rect -2255 -85 -2209 -39
rect -2131 -85 -2085 -39
rect -2007 -85 -1961 -39
rect -1883 -85 -1837 -39
rect -1759 -85 -1713 -39
rect -1635 -85 -1589 -39
rect -1511 -85 -1465 -39
rect -1387 -85 -1341 -39
rect -1263 -85 -1217 -39
rect -1139 -85 -1093 -39
rect -1015 -85 -969 -39
rect -891 -85 -845 -39
rect -767 -85 -721 -39
rect -643 -85 -597 -39
rect -519 -85 -473 -39
rect -395 -85 -349 -39
rect -271 -85 -225 -39
rect -147 -85 -101 -39
rect -23 -85 23 -39
rect 101 -85 147 -39
rect 225 -85 271 -39
rect 349 -85 395 -39
rect 473 -85 519 -39
rect 597 -85 643 -39
rect 721 -85 767 -39
rect 845 -85 891 -39
rect 969 -85 1015 -39
rect 1093 -85 1139 -39
rect 1217 -85 1263 -39
rect 1341 -85 1387 -39
rect 1465 -85 1511 -39
rect 1589 -85 1635 -39
rect 1713 -85 1759 -39
rect 1837 -85 1883 -39
rect 1961 -85 2007 -39
rect 2085 -85 2131 -39
rect 2209 -85 2255 -39
rect 2333 -85 2379 -39
rect 2457 -85 2503 -39
rect 2581 -85 2627 -39
rect -2627 -209 -2581 -163
rect -2503 -209 -2457 -163
rect -2379 -209 -2333 -163
rect -2255 -209 -2209 -163
rect -2131 -209 -2085 -163
rect -2007 -209 -1961 -163
rect -1883 -209 -1837 -163
rect -1759 -209 -1713 -163
rect -1635 -209 -1589 -163
rect -1511 -209 -1465 -163
rect -1387 -209 -1341 -163
rect -1263 -209 -1217 -163
rect -1139 -209 -1093 -163
rect -1015 -209 -969 -163
rect -891 -209 -845 -163
rect -767 -209 -721 -163
rect -643 -209 -597 -163
rect -519 -209 -473 -163
rect -395 -209 -349 -163
rect -271 -209 -225 -163
rect -147 -209 -101 -163
rect -23 -209 23 -163
rect 101 -209 147 -163
rect 225 -209 271 -163
rect 349 -209 395 -163
rect 473 -209 519 -163
rect 597 -209 643 -163
rect 721 -209 767 -163
rect 845 -209 891 -163
rect 969 -209 1015 -163
rect 1093 -209 1139 -163
rect 1217 -209 1263 -163
rect 1341 -209 1387 -163
rect 1465 -209 1511 -163
rect 1589 -209 1635 -163
rect 1713 -209 1759 -163
rect 1837 -209 1883 -163
rect 1961 -209 2007 -163
rect 2085 -209 2131 -163
rect 2209 -209 2255 -163
rect 2333 -209 2379 -163
rect 2457 -209 2503 -163
rect 2581 -209 2627 -163
rect -2627 -333 -2581 -287
rect -2503 -333 -2457 -287
rect -2379 -333 -2333 -287
rect -2255 -333 -2209 -287
rect -2131 -333 -2085 -287
rect -2007 -333 -1961 -287
rect -1883 -333 -1837 -287
rect -1759 -333 -1713 -287
rect -1635 -333 -1589 -287
rect -1511 -333 -1465 -287
rect -1387 -333 -1341 -287
rect -1263 -333 -1217 -287
rect -1139 -333 -1093 -287
rect -1015 -333 -969 -287
rect -891 -333 -845 -287
rect -767 -333 -721 -287
rect -643 -333 -597 -287
rect -519 -333 -473 -287
rect -395 -333 -349 -287
rect -271 -333 -225 -287
rect -147 -333 -101 -287
rect -23 -333 23 -287
rect 101 -333 147 -287
rect 225 -333 271 -287
rect 349 -333 395 -287
rect 473 -333 519 -287
rect 597 -333 643 -287
rect 721 -333 767 -287
rect 845 -333 891 -287
rect 969 -333 1015 -287
rect 1093 -333 1139 -287
rect 1217 -333 1263 -287
rect 1341 -333 1387 -287
rect 1465 -333 1511 -287
rect 1589 -333 1635 -287
rect 1713 -333 1759 -287
rect 1837 -333 1883 -287
rect 1961 -333 2007 -287
rect 2085 -333 2131 -287
rect 2209 -333 2255 -287
rect 2333 -333 2379 -287
rect 2457 -333 2503 -287
rect 2581 -333 2627 -287
rect -2627 -457 -2581 -411
rect -2503 -457 -2457 -411
rect -2379 -457 -2333 -411
rect -2255 -457 -2209 -411
rect -2131 -457 -2085 -411
rect -2007 -457 -1961 -411
rect -1883 -457 -1837 -411
rect -1759 -457 -1713 -411
rect -1635 -457 -1589 -411
rect -1511 -457 -1465 -411
rect -1387 -457 -1341 -411
rect -1263 -457 -1217 -411
rect -1139 -457 -1093 -411
rect -1015 -457 -969 -411
rect -891 -457 -845 -411
rect -767 -457 -721 -411
rect -643 -457 -597 -411
rect -519 -457 -473 -411
rect -395 -457 -349 -411
rect -271 -457 -225 -411
rect -147 -457 -101 -411
rect -23 -457 23 -411
rect 101 -457 147 -411
rect 225 -457 271 -411
rect 349 -457 395 -411
rect 473 -457 519 -411
rect 597 -457 643 -411
rect 721 -457 767 -411
rect 845 -457 891 -411
rect 969 -457 1015 -411
rect 1093 -457 1139 -411
rect 1217 -457 1263 -411
rect 1341 -457 1387 -411
rect 1465 -457 1511 -411
rect 1589 -457 1635 -411
rect 1713 -457 1759 -411
rect 1837 -457 1883 -411
rect 1961 -457 2007 -411
rect 2085 -457 2131 -411
rect 2209 -457 2255 -411
rect 2333 -457 2379 -411
rect 2457 -457 2503 -411
rect 2581 -457 2627 -411
rect -2627 -581 -2581 -535
rect -2503 -581 -2457 -535
rect -2379 -581 -2333 -535
rect -2255 -581 -2209 -535
rect -2131 -581 -2085 -535
rect -2007 -581 -1961 -535
rect -1883 -581 -1837 -535
rect -1759 -581 -1713 -535
rect -1635 -581 -1589 -535
rect -1511 -581 -1465 -535
rect -1387 -581 -1341 -535
rect -1263 -581 -1217 -535
rect -1139 -581 -1093 -535
rect -1015 -581 -969 -535
rect -891 -581 -845 -535
rect -767 -581 -721 -535
rect -643 -581 -597 -535
rect -519 -581 -473 -535
rect -395 -581 -349 -535
rect -271 -581 -225 -535
rect -147 -581 -101 -535
rect -23 -581 23 -535
rect 101 -581 147 -535
rect 225 -581 271 -535
rect 349 -581 395 -535
rect 473 -581 519 -535
rect 597 -581 643 -535
rect 721 -581 767 -535
rect 845 -581 891 -535
rect 969 -581 1015 -535
rect 1093 -581 1139 -535
rect 1217 -581 1263 -535
rect 1341 -581 1387 -535
rect 1465 -581 1511 -535
rect 1589 -581 1635 -535
rect 1713 -581 1759 -535
rect 1837 -581 1883 -535
rect 1961 -581 2007 -535
rect 2085 -581 2131 -535
rect 2209 -581 2255 -535
rect 2333 -581 2379 -535
rect 2457 -581 2503 -535
rect 2581 -581 2627 -535
rect -2627 -705 -2581 -659
rect -2503 -705 -2457 -659
rect -2379 -705 -2333 -659
rect -2255 -705 -2209 -659
rect -2131 -705 -2085 -659
rect -2007 -705 -1961 -659
rect -1883 -705 -1837 -659
rect -1759 -705 -1713 -659
rect -1635 -705 -1589 -659
rect -1511 -705 -1465 -659
rect -1387 -705 -1341 -659
rect -1263 -705 -1217 -659
rect -1139 -705 -1093 -659
rect -1015 -705 -969 -659
rect -891 -705 -845 -659
rect -767 -705 -721 -659
rect -643 -705 -597 -659
rect -519 -705 -473 -659
rect -395 -705 -349 -659
rect -271 -705 -225 -659
rect -147 -705 -101 -659
rect -23 -705 23 -659
rect 101 -705 147 -659
rect 225 -705 271 -659
rect 349 -705 395 -659
rect 473 -705 519 -659
rect 597 -705 643 -659
rect 721 -705 767 -659
rect 845 -705 891 -659
rect 969 -705 1015 -659
rect 1093 -705 1139 -659
rect 1217 -705 1263 -659
rect 1341 -705 1387 -659
rect 1465 -705 1511 -659
rect 1589 -705 1635 -659
rect 1713 -705 1759 -659
rect 1837 -705 1883 -659
rect 1961 -705 2007 -659
rect 2085 -705 2131 -659
rect 2209 -705 2255 -659
rect 2333 -705 2379 -659
rect 2457 -705 2503 -659
rect 2581 -705 2627 -659
rect -2627 -829 -2581 -783
rect -2503 -829 -2457 -783
rect -2379 -829 -2333 -783
rect -2255 -829 -2209 -783
rect -2131 -829 -2085 -783
rect -2007 -829 -1961 -783
rect -1883 -829 -1837 -783
rect -1759 -829 -1713 -783
rect -1635 -829 -1589 -783
rect -1511 -829 -1465 -783
rect -1387 -829 -1341 -783
rect -1263 -829 -1217 -783
rect -1139 -829 -1093 -783
rect -1015 -829 -969 -783
rect -891 -829 -845 -783
rect -767 -829 -721 -783
rect -643 -829 -597 -783
rect -519 -829 -473 -783
rect -395 -829 -349 -783
rect -271 -829 -225 -783
rect -147 -829 -101 -783
rect -23 -829 23 -783
rect 101 -829 147 -783
rect 225 -829 271 -783
rect 349 -829 395 -783
rect 473 -829 519 -783
rect 597 -829 643 -783
rect 721 -829 767 -783
rect 845 -829 891 -783
rect 969 -829 1015 -783
rect 1093 -829 1139 -783
rect 1217 -829 1263 -783
rect 1341 -829 1387 -783
rect 1465 -829 1511 -783
rect 1589 -829 1635 -783
rect 1713 -829 1759 -783
rect 1837 -829 1883 -783
rect 1961 -829 2007 -783
rect 2085 -829 2131 -783
rect 2209 -829 2255 -783
rect 2333 -829 2379 -783
rect 2457 -829 2503 -783
rect 2581 -829 2627 -783
rect -2627 -953 -2581 -907
rect -2503 -953 -2457 -907
rect -2379 -953 -2333 -907
rect -2255 -953 -2209 -907
rect -2131 -953 -2085 -907
rect -2007 -953 -1961 -907
rect -1883 -953 -1837 -907
rect -1759 -953 -1713 -907
rect -1635 -953 -1589 -907
rect -1511 -953 -1465 -907
rect -1387 -953 -1341 -907
rect -1263 -953 -1217 -907
rect -1139 -953 -1093 -907
rect -1015 -953 -969 -907
rect -891 -953 -845 -907
rect -767 -953 -721 -907
rect -643 -953 -597 -907
rect -519 -953 -473 -907
rect -395 -953 -349 -907
rect -271 -953 -225 -907
rect -147 -953 -101 -907
rect -23 -953 23 -907
rect 101 -953 147 -907
rect 225 -953 271 -907
rect 349 -953 395 -907
rect 473 -953 519 -907
rect 597 -953 643 -907
rect 721 -953 767 -907
rect 845 -953 891 -907
rect 969 -953 1015 -907
rect 1093 -953 1139 -907
rect 1217 -953 1263 -907
rect 1341 -953 1387 -907
rect 1465 -953 1511 -907
rect 1589 -953 1635 -907
rect 1713 -953 1759 -907
rect 1837 -953 1883 -907
rect 1961 -953 2007 -907
rect 2085 -953 2131 -907
rect 2209 -953 2255 -907
rect 2333 -953 2379 -907
rect 2457 -953 2503 -907
rect 2581 -953 2627 -907
<< metal1 >>
rect -2638 953 2638 964
rect -2638 907 -2627 953
rect -2581 907 -2503 953
rect -2457 907 -2379 953
rect -2333 907 -2255 953
rect -2209 907 -2131 953
rect -2085 907 -2007 953
rect -1961 907 -1883 953
rect -1837 907 -1759 953
rect -1713 907 -1635 953
rect -1589 907 -1511 953
rect -1465 907 -1387 953
rect -1341 907 -1263 953
rect -1217 907 -1139 953
rect -1093 907 -1015 953
rect -969 907 -891 953
rect -845 907 -767 953
rect -721 907 -643 953
rect -597 907 -519 953
rect -473 907 -395 953
rect -349 907 -271 953
rect -225 907 -147 953
rect -101 907 -23 953
rect 23 907 101 953
rect 147 907 225 953
rect 271 907 349 953
rect 395 907 473 953
rect 519 907 597 953
rect 643 907 721 953
rect 767 907 845 953
rect 891 907 969 953
rect 1015 907 1093 953
rect 1139 907 1217 953
rect 1263 907 1341 953
rect 1387 907 1465 953
rect 1511 907 1589 953
rect 1635 907 1713 953
rect 1759 907 1837 953
rect 1883 907 1961 953
rect 2007 907 2085 953
rect 2131 907 2209 953
rect 2255 907 2333 953
rect 2379 907 2457 953
rect 2503 907 2581 953
rect 2627 907 2638 953
rect -2638 829 2638 907
rect -2638 783 -2627 829
rect -2581 783 -2503 829
rect -2457 783 -2379 829
rect -2333 783 -2255 829
rect -2209 783 -2131 829
rect -2085 783 -2007 829
rect -1961 783 -1883 829
rect -1837 783 -1759 829
rect -1713 783 -1635 829
rect -1589 783 -1511 829
rect -1465 783 -1387 829
rect -1341 783 -1263 829
rect -1217 783 -1139 829
rect -1093 783 -1015 829
rect -969 783 -891 829
rect -845 783 -767 829
rect -721 783 -643 829
rect -597 783 -519 829
rect -473 783 -395 829
rect -349 783 -271 829
rect -225 783 -147 829
rect -101 783 -23 829
rect 23 783 101 829
rect 147 783 225 829
rect 271 783 349 829
rect 395 783 473 829
rect 519 783 597 829
rect 643 783 721 829
rect 767 783 845 829
rect 891 783 969 829
rect 1015 783 1093 829
rect 1139 783 1217 829
rect 1263 783 1341 829
rect 1387 783 1465 829
rect 1511 783 1589 829
rect 1635 783 1713 829
rect 1759 783 1837 829
rect 1883 783 1961 829
rect 2007 783 2085 829
rect 2131 783 2209 829
rect 2255 783 2333 829
rect 2379 783 2457 829
rect 2503 783 2581 829
rect 2627 783 2638 829
rect -2638 705 2638 783
rect -2638 659 -2627 705
rect -2581 659 -2503 705
rect -2457 659 -2379 705
rect -2333 659 -2255 705
rect -2209 659 -2131 705
rect -2085 659 -2007 705
rect -1961 659 -1883 705
rect -1837 659 -1759 705
rect -1713 659 -1635 705
rect -1589 659 -1511 705
rect -1465 659 -1387 705
rect -1341 659 -1263 705
rect -1217 659 -1139 705
rect -1093 659 -1015 705
rect -969 659 -891 705
rect -845 659 -767 705
rect -721 659 -643 705
rect -597 659 -519 705
rect -473 659 -395 705
rect -349 659 -271 705
rect -225 659 -147 705
rect -101 659 -23 705
rect 23 659 101 705
rect 147 659 225 705
rect 271 659 349 705
rect 395 659 473 705
rect 519 659 597 705
rect 643 659 721 705
rect 767 659 845 705
rect 891 659 969 705
rect 1015 659 1093 705
rect 1139 659 1217 705
rect 1263 659 1341 705
rect 1387 659 1465 705
rect 1511 659 1589 705
rect 1635 659 1713 705
rect 1759 659 1837 705
rect 1883 659 1961 705
rect 2007 659 2085 705
rect 2131 659 2209 705
rect 2255 659 2333 705
rect 2379 659 2457 705
rect 2503 659 2581 705
rect 2627 659 2638 705
rect -2638 581 2638 659
rect -2638 535 -2627 581
rect -2581 535 -2503 581
rect -2457 535 -2379 581
rect -2333 535 -2255 581
rect -2209 535 -2131 581
rect -2085 535 -2007 581
rect -1961 535 -1883 581
rect -1837 535 -1759 581
rect -1713 535 -1635 581
rect -1589 535 -1511 581
rect -1465 535 -1387 581
rect -1341 535 -1263 581
rect -1217 535 -1139 581
rect -1093 535 -1015 581
rect -969 535 -891 581
rect -845 535 -767 581
rect -721 535 -643 581
rect -597 535 -519 581
rect -473 535 -395 581
rect -349 535 -271 581
rect -225 535 -147 581
rect -101 535 -23 581
rect 23 535 101 581
rect 147 535 225 581
rect 271 535 349 581
rect 395 535 473 581
rect 519 535 597 581
rect 643 535 721 581
rect 767 535 845 581
rect 891 535 969 581
rect 1015 535 1093 581
rect 1139 535 1217 581
rect 1263 535 1341 581
rect 1387 535 1465 581
rect 1511 535 1589 581
rect 1635 535 1713 581
rect 1759 535 1837 581
rect 1883 535 1961 581
rect 2007 535 2085 581
rect 2131 535 2209 581
rect 2255 535 2333 581
rect 2379 535 2457 581
rect 2503 535 2581 581
rect 2627 535 2638 581
rect -2638 457 2638 535
rect -2638 411 -2627 457
rect -2581 411 -2503 457
rect -2457 411 -2379 457
rect -2333 411 -2255 457
rect -2209 411 -2131 457
rect -2085 411 -2007 457
rect -1961 411 -1883 457
rect -1837 411 -1759 457
rect -1713 411 -1635 457
rect -1589 411 -1511 457
rect -1465 411 -1387 457
rect -1341 411 -1263 457
rect -1217 411 -1139 457
rect -1093 411 -1015 457
rect -969 411 -891 457
rect -845 411 -767 457
rect -721 411 -643 457
rect -597 411 -519 457
rect -473 411 -395 457
rect -349 411 -271 457
rect -225 411 -147 457
rect -101 411 -23 457
rect 23 411 101 457
rect 147 411 225 457
rect 271 411 349 457
rect 395 411 473 457
rect 519 411 597 457
rect 643 411 721 457
rect 767 411 845 457
rect 891 411 969 457
rect 1015 411 1093 457
rect 1139 411 1217 457
rect 1263 411 1341 457
rect 1387 411 1465 457
rect 1511 411 1589 457
rect 1635 411 1713 457
rect 1759 411 1837 457
rect 1883 411 1961 457
rect 2007 411 2085 457
rect 2131 411 2209 457
rect 2255 411 2333 457
rect 2379 411 2457 457
rect 2503 411 2581 457
rect 2627 411 2638 457
rect -2638 333 2638 411
rect -2638 287 -2627 333
rect -2581 287 -2503 333
rect -2457 287 -2379 333
rect -2333 287 -2255 333
rect -2209 287 -2131 333
rect -2085 287 -2007 333
rect -1961 287 -1883 333
rect -1837 287 -1759 333
rect -1713 287 -1635 333
rect -1589 287 -1511 333
rect -1465 287 -1387 333
rect -1341 287 -1263 333
rect -1217 287 -1139 333
rect -1093 287 -1015 333
rect -969 287 -891 333
rect -845 287 -767 333
rect -721 287 -643 333
rect -597 287 -519 333
rect -473 287 -395 333
rect -349 287 -271 333
rect -225 287 -147 333
rect -101 287 -23 333
rect 23 287 101 333
rect 147 287 225 333
rect 271 287 349 333
rect 395 287 473 333
rect 519 287 597 333
rect 643 287 721 333
rect 767 287 845 333
rect 891 287 969 333
rect 1015 287 1093 333
rect 1139 287 1217 333
rect 1263 287 1341 333
rect 1387 287 1465 333
rect 1511 287 1589 333
rect 1635 287 1713 333
rect 1759 287 1837 333
rect 1883 287 1961 333
rect 2007 287 2085 333
rect 2131 287 2209 333
rect 2255 287 2333 333
rect 2379 287 2457 333
rect 2503 287 2581 333
rect 2627 287 2638 333
rect -2638 209 2638 287
rect -2638 163 -2627 209
rect -2581 163 -2503 209
rect -2457 163 -2379 209
rect -2333 163 -2255 209
rect -2209 163 -2131 209
rect -2085 163 -2007 209
rect -1961 163 -1883 209
rect -1837 163 -1759 209
rect -1713 163 -1635 209
rect -1589 163 -1511 209
rect -1465 163 -1387 209
rect -1341 163 -1263 209
rect -1217 163 -1139 209
rect -1093 163 -1015 209
rect -969 163 -891 209
rect -845 163 -767 209
rect -721 163 -643 209
rect -597 163 -519 209
rect -473 163 -395 209
rect -349 163 -271 209
rect -225 163 -147 209
rect -101 163 -23 209
rect 23 163 101 209
rect 147 163 225 209
rect 271 163 349 209
rect 395 163 473 209
rect 519 163 597 209
rect 643 163 721 209
rect 767 163 845 209
rect 891 163 969 209
rect 1015 163 1093 209
rect 1139 163 1217 209
rect 1263 163 1341 209
rect 1387 163 1465 209
rect 1511 163 1589 209
rect 1635 163 1713 209
rect 1759 163 1837 209
rect 1883 163 1961 209
rect 2007 163 2085 209
rect 2131 163 2209 209
rect 2255 163 2333 209
rect 2379 163 2457 209
rect 2503 163 2581 209
rect 2627 163 2638 209
rect -2638 85 2638 163
rect -2638 39 -2627 85
rect -2581 39 -2503 85
rect -2457 39 -2379 85
rect -2333 39 -2255 85
rect -2209 39 -2131 85
rect -2085 39 -2007 85
rect -1961 39 -1883 85
rect -1837 39 -1759 85
rect -1713 39 -1635 85
rect -1589 39 -1511 85
rect -1465 39 -1387 85
rect -1341 39 -1263 85
rect -1217 39 -1139 85
rect -1093 39 -1015 85
rect -969 39 -891 85
rect -845 39 -767 85
rect -721 39 -643 85
rect -597 39 -519 85
rect -473 39 -395 85
rect -349 39 -271 85
rect -225 39 -147 85
rect -101 39 -23 85
rect 23 39 101 85
rect 147 39 225 85
rect 271 39 349 85
rect 395 39 473 85
rect 519 39 597 85
rect 643 39 721 85
rect 767 39 845 85
rect 891 39 969 85
rect 1015 39 1093 85
rect 1139 39 1217 85
rect 1263 39 1341 85
rect 1387 39 1465 85
rect 1511 39 1589 85
rect 1635 39 1713 85
rect 1759 39 1837 85
rect 1883 39 1961 85
rect 2007 39 2085 85
rect 2131 39 2209 85
rect 2255 39 2333 85
rect 2379 39 2457 85
rect 2503 39 2581 85
rect 2627 39 2638 85
rect -2638 -39 2638 39
rect -2638 -85 -2627 -39
rect -2581 -85 -2503 -39
rect -2457 -85 -2379 -39
rect -2333 -85 -2255 -39
rect -2209 -85 -2131 -39
rect -2085 -85 -2007 -39
rect -1961 -85 -1883 -39
rect -1837 -85 -1759 -39
rect -1713 -85 -1635 -39
rect -1589 -85 -1511 -39
rect -1465 -85 -1387 -39
rect -1341 -85 -1263 -39
rect -1217 -85 -1139 -39
rect -1093 -85 -1015 -39
rect -969 -85 -891 -39
rect -845 -85 -767 -39
rect -721 -85 -643 -39
rect -597 -85 -519 -39
rect -473 -85 -395 -39
rect -349 -85 -271 -39
rect -225 -85 -147 -39
rect -101 -85 -23 -39
rect 23 -85 101 -39
rect 147 -85 225 -39
rect 271 -85 349 -39
rect 395 -85 473 -39
rect 519 -85 597 -39
rect 643 -85 721 -39
rect 767 -85 845 -39
rect 891 -85 969 -39
rect 1015 -85 1093 -39
rect 1139 -85 1217 -39
rect 1263 -85 1341 -39
rect 1387 -85 1465 -39
rect 1511 -85 1589 -39
rect 1635 -85 1713 -39
rect 1759 -85 1837 -39
rect 1883 -85 1961 -39
rect 2007 -85 2085 -39
rect 2131 -85 2209 -39
rect 2255 -85 2333 -39
rect 2379 -85 2457 -39
rect 2503 -85 2581 -39
rect 2627 -85 2638 -39
rect -2638 -163 2638 -85
rect -2638 -209 -2627 -163
rect -2581 -209 -2503 -163
rect -2457 -209 -2379 -163
rect -2333 -209 -2255 -163
rect -2209 -209 -2131 -163
rect -2085 -209 -2007 -163
rect -1961 -209 -1883 -163
rect -1837 -209 -1759 -163
rect -1713 -209 -1635 -163
rect -1589 -209 -1511 -163
rect -1465 -209 -1387 -163
rect -1341 -209 -1263 -163
rect -1217 -209 -1139 -163
rect -1093 -209 -1015 -163
rect -969 -209 -891 -163
rect -845 -209 -767 -163
rect -721 -209 -643 -163
rect -597 -209 -519 -163
rect -473 -209 -395 -163
rect -349 -209 -271 -163
rect -225 -209 -147 -163
rect -101 -209 -23 -163
rect 23 -209 101 -163
rect 147 -209 225 -163
rect 271 -209 349 -163
rect 395 -209 473 -163
rect 519 -209 597 -163
rect 643 -209 721 -163
rect 767 -209 845 -163
rect 891 -209 969 -163
rect 1015 -209 1093 -163
rect 1139 -209 1217 -163
rect 1263 -209 1341 -163
rect 1387 -209 1465 -163
rect 1511 -209 1589 -163
rect 1635 -209 1713 -163
rect 1759 -209 1837 -163
rect 1883 -209 1961 -163
rect 2007 -209 2085 -163
rect 2131 -209 2209 -163
rect 2255 -209 2333 -163
rect 2379 -209 2457 -163
rect 2503 -209 2581 -163
rect 2627 -209 2638 -163
rect -2638 -287 2638 -209
rect -2638 -333 -2627 -287
rect -2581 -333 -2503 -287
rect -2457 -333 -2379 -287
rect -2333 -333 -2255 -287
rect -2209 -333 -2131 -287
rect -2085 -333 -2007 -287
rect -1961 -333 -1883 -287
rect -1837 -333 -1759 -287
rect -1713 -333 -1635 -287
rect -1589 -333 -1511 -287
rect -1465 -333 -1387 -287
rect -1341 -333 -1263 -287
rect -1217 -333 -1139 -287
rect -1093 -333 -1015 -287
rect -969 -333 -891 -287
rect -845 -333 -767 -287
rect -721 -333 -643 -287
rect -597 -333 -519 -287
rect -473 -333 -395 -287
rect -349 -333 -271 -287
rect -225 -333 -147 -287
rect -101 -333 -23 -287
rect 23 -333 101 -287
rect 147 -333 225 -287
rect 271 -333 349 -287
rect 395 -333 473 -287
rect 519 -333 597 -287
rect 643 -333 721 -287
rect 767 -333 845 -287
rect 891 -333 969 -287
rect 1015 -333 1093 -287
rect 1139 -333 1217 -287
rect 1263 -333 1341 -287
rect 1387 -333 1465 -287
rect 1511 -333 1589 -287
rect 1635 -333 1713 -287
rect 1759 -333 1837 -287
rect 1883 -333 1961 -287
rect 2007 -333 2085 -287
rect 2131 -333 2209 -287
rect 2255 -333 2333 -287
rect 2379 -333 2457 -287
rect 2503 -333 2581 -287
rect 2627 -333 2638 -287
rect -2638 -411 2638 -333
rect -2638 -457 -2627 -411
rect -2581 -457 -2503 -411
rect -2457 -457 -2379 -411
rect -2333 -457 -2255 -411
rect -2209 -457 -2131 -411
rect -2085 -457 -2007 -411
rect -1961 -457 -1883 -411
rect -1837 -457 -1759 -411
rect -1713 -457 -1635 -411
rect -1589 -457 -1511 -411
rect -1465 -457 -1387 -411
rect -1341 -457 -1263 -411
rect -1217 -457 -1139 -411
rect -1093 -457 -1015 -411
rect -969 -457 -891 -411
rect -845 -457 -767 -411
rect -721 -457 -643 -411
rect -597 -457 -519 -411
rect -473 -457 -395 -411
rect -349 -457 -271 -411
rect -225 -457 -147 -411
rect -101 -457 -23 -411
rect 23 -457 101 -411
rect 147 -457 225 -411
rect 271 -457 349 -411
rect 395 -457 473 -411
rect 519 -457 597 -411
rect 643 -457 721 -411
rect 767 -457 845 -411
rect 891 -457 969 -411
rect 1015 -457 1093 -411
rect 1139 -457 1217 -411
rect 1263 -457 1341 -411
rect 1387 -457 1465 -411
rect 1511 -457 1589 -411
rect 1635 -457 1713 -411
rect 1759 -457 1837 -411
rect 1883 -457 1961 -411
rect 2007 -457 2085 -411
rect 2131 -457 2209 -411
rect 2255 -457 2333 -411
rect 2379 -457 2457 -411
rect 2503 -457 2581 -411
rect 2627 -457 2638 -411
rect -2638 -535 2638 -457
rect -2638 -581 -2627 -535
rect -2581 -581 -2503 -535
rect -2457 -581 -2379 -535
rect -2333 -581 -2255 -535
rect -2209 -581 -2131 -535
rect -2085 -581 -2007 -535
rect -1961 -581 -1883 -535
rect -1837 -581 -1759 -535
rect -1713 -581 -1635 -535
rect -1589 -581 -1511 -535
rect -1465 -581 -1387 -535
rect -1341 -581 -1263 -535
rect -1217 -581 -1139 -535
rect -1093 -581 -1015 -535
rect -969 -581 -891 -535
rect -845 -581 -767 -535
rect -721 -581 -643 -535
rect -597 -581 -519 -535
rect -473 -581 -395 -535
rect -349 -581 -271 -535
rect -225 -581 -147 -535
rect -101 -581 -23 -535
rect 23 -581 101 -535
rect 147 -581 225 -535
rect 271 -581 349 -535
rect 395 -581 473 -535
rect 519 -581 597 -535
rect 643 -581 721 -535
rect 767 -581 845 -535
rect 891 -581 969 -535
rect 1015 -581 1093 -535
rect 1139 -581 1217 -535
rect 1263 -581 1341 -535
rect 1387 -581 1465 -535
rect 1511 -581 1589 -535
rect 1635 -581 1713 -535
rect 1759 -581 1837 -535
rect 1883 -581 1961 -535
rect 2007 -581 2085 -535
rect 2131 -581 2209 -535
rect 2255 -581 2333 -535
rect 2379 -581 2457 -535
rect 2503 -581 2581 -535
rect 2627 -581 2638 -535
rect -2638 -659 2638 -581
rect -2638 -705 -2627 -659
rect -2581 -705 -2503 -659
rect -2457 -705 -2379 -659
rect -2333 -705 -2255 -659
rect -2209 -705 -2131 -659
rect -2085 -705 -2007 -659
rect -1961 -705 -1883 -659
rect -1837 -705 -1759 -659
rect -1713 -705 -1635 -659
rect -1589 -705 -1511 -659
rect -1465 -705 -1387 -659
rect -1341 -705 -1263 -659
rect -1217 -705 -1139 -659
rect -1093 -705 -1015 -659
rect -969 -705 -891 -659
rect -845 -705 -767 -659
rect -721 -705 -643 -659
rect -597 -705 -519 -659
rect -473 -705 -395 -659
rect -349 -705 -271 -659
rect -225 -705 -147 -659
rect -101 -705 -23 -659
rect 23 -705 101 -659
rect 147 -705 225 -659
rect 271 -705 349 -659
rect 395 -705 473 -659
rect 519 -705 597 -659
rect 643 -705 721 -659
rect 767 -705 845 -659
rect 891 -705 969 -659
rect 1015 -705 1093 -659
rect 1139 -705 1217 -659
rect 1263 -705 1341 -659
rect 1387 -705 1465 -659
rect 1511 -705 1589 -659
rect 1635 -705 1713 -659
rect 1759 -705 1837 -659
rect 1883 -705 1961 -659
rect 2007 -705 2085 -659
rect 2131 -705 2209 -659
rect 2255 -705 2333 -659
rect 2379 -705 2457 -659
rect 2503 -705 2581 -659
rect 2627 -705 2638 -659
rect -2638 -783 2638 -705
rect -2638 -829 -2627 -783
rect -2581 -829 -2503 -783
rect -2457 -829 -2379 -783
rect -2333 -829 -2255 -783
rect -2209 -829 -2131 -783
rect -2085 -829 -2007 -783
rect -1961 -829 -1883 -783
rect -1837 -829 -1759 -783
rect -1713 -829 -1635 -783
rect -1589 -829 -1511 -783
rect -1465 -829 -1387 -783
rect -1341 -829 -1263 -783
rect -1217 -829 -1139 -783
rect -1093 -829 -1015 -783
rect -969 -829 -891 -783
rect -845 -829 -767 -783
rect -721 -829 -643 -783
rect -597 -829 -519 -783
rect -473 -829 -395 -783
rect -349 -829 -271 -783
rect -225 -829 -147 -783
rect -101 -829 -23 -783
rect 23 -829 101 -783
rect 147 -829 225 -783
rect 271 -829 349 -783
rect 395 -829 473 -783
rect 519 -829 597 -783
rect 643 -829 721 -783
rect 767 -829 845 -783
rect 891 -829 969 -783
rect 1015 -829 1093 -783
rect 1139 -829 1217 -783
rect 1263 -829 1341 -783
rect 1387 -829 1465 -783
rect 1511 -829 1589 -783
rect 1635 -829 1713 -783
rect 1759 -829 1837 -783
rect 1883 -829 1961 -783
rect 2007 -829 2085 -783
rect 2131 -829 2209 -783
rect 2255 -829 2333 -783
rect 2379 -829 2457 -783
rect 2503 -829 2581 -783
rect 2627 -829 2638 -783
rect -2638 -907 2638 -829
rect -2638 -953 -2627 -907
rect -2581 -953 -2503 -907
rect -2457 -953 -2379 -907
rect -2333 -953 -2255 -907
rect -2209 -953 -2131 -907
rect -2085 -953 -2007 -907
rect -1961 -953 -1883 -907
rect -1837 -953 -1759 -907
rect -1713 -953 -1635 -907
rect -1589 -953 -1511 -907
rect -1465 -953 -1387 -907
rect -1341 -953 -1263 -907
rect -1217 -953 -1139 -907
rect -1093 -953 -1015 -907
rect -969 -953 -891 -907
rect -845 -953 -767 -907
rect -721 -953 -643 -907
rect -597 -953 -519 -907
rect -473 -953 -395 -907
rect -349 -953 -271 -907
rect -225 -953 -147 -907
rect -101 -953 -23 -907
rect 23 -953 101 -907
rect 147 -953 225 -907
rect 271 -953 349 -907
rect 395 -953 473 -907
rect 519 -953 597 -907
rect 643 -953 721 -907
rect 767 -953 845 -907
rect 891 -953 969 -907
rect 1015 -953 1093 -907
rect 1139 -953 1217 -907
rect 1263 -953 1341 -907
rect 1387 -953 1465 -907
rect 1511 -953 1589 -907
rect 1635 -953 1713 -907
rect 1759 -953 1837 -907
rect 1883 -953 1961 -907
rect 2007 -953 2085 -907
rect 2131 -953 2209 -907
rect 2255 -953 2333 -907
rect 2379 -953 2457 -907
rect 2503 -953 2581 -907
rect 2627 -953 2638 -907
rect -2638 -964 2638 -953
<< end >>
