magic
tech gf180mcuD
magscale 1 10
timestamp 1713530186
<< checkpaint >>
rect 15348 402 844842 4646
rect 1168852 4159 1366706 4563
rect 978500 877 1366706 4159
rect 978500 402 1394912 877
rect 15348 -3363 1394912 402
rect -2000 -10400 1394912 -3363
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
use x7b_counter  X7b_counter_0
timestamp 1713530185
transform 1 0 17348 0 1 -400
box 0 -8000 825494 3046
use DFF_magic  XDFF_magic_0
timestamp 1713530183
transform 1 0 940250 0 1 -5445
box -5636 -2955 40250 3847
use divide_by_2  Xdivide_by_2_0
timestamp 1713530185
transform 1 0 848478 0 1 -5445
box -5636 -2955 40250 3847
use divide_by_2  Xdivide_by_2_1
timestamp 1713530185
transform 1 0 894364 0 1 -5445
box -5636 -2955 40250 3847
use mux_magic  Xmux_magic_0
timestamp 1713530184
transform 1 0 1366530 0 1 -2671
box -1824 -5729 26382 1548
use OR_magic  XOR_magic_1
timestamp 1713530181
transform 1 0 812 0 1 -5974
box -812 -2426 7862 611
use OR_magic  XOR_magic_2
timestamp 1713530181
transform 1 0 9486 0 1 -5974
box -812 -2426 7862 611
use p2_gen_magic  Xp2_gen_magic_0
timestamp 1713530185
transform 1 0 980938 0 1 -2000
box -438 -6400 189914 4159
use p3_gen_magic  Xp3_gen_magic_0
timestamp 1713530186
transform 1 0 1171290 0 1 -1600
box -438 -6800 193416 4163
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 1280 0 0 0 P2
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 1280 0 0 0 OUT1
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 1280 0 0 0 VDD
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 1280 0 0 0 Q1
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 1280 0 0 0 Q2
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 1280 0 0 0 Q3
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 1280 0 0 0 D2_3
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 1280 0 0 0 D2_6
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 1280 0 0 0 D2_7
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 1280 0 0 0 LD
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 1280 0 0 0 D2_5
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 1280 0 0 0 D2_4
port 11 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 1280 0 0 0 {}
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 1280 0 0 0 D2_1
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 1280 0 0 0 CLK
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 1280 0 0 0 Q6
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 1280 0 0 0 Q7
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 1280 0 0 0 Q5
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 1280 0 0 0 VSS
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 1280 0 0 0 Q4
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 1280 0 0 0 D2_2
port 21 nsew
<< end >>
