magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -2636 -1151 2636 1151
<< metal1 >>
rect -1636 145 1636 151
rect -1636 119 -1630 145
rect -1604 119 -1564 145
rect -1538 119 -1498 145
rect -1472 119 -1432 145
rect -1406 119 -1366 145
rect -1340 119 -1300 145
rect -1274 119 -1234 145
rect -1208 119 -1168 145
rect -1142 119 -1102 145
rect -1076 119 -1036 145
rect -1010 119 -970 145
rect -944 119 -904 145
rect -878 119 -838 145
rect -812 119 -772 145
rect -746 119 -706 145
rect -680 119 -640 145
rect -614 119 -574 145
rect -548 119 -508 145
rect -482 119 -442 145
rect -416 119 -376 145
rect -350 119 -310 145
rect -284 119 -244 145
rect -218 119 -178 145
rect -152 119 -112 145
rect -86 119 -46 145
rect -20 119 20 145
rect 46 119 86 145
rect 112 119 152 145
rect 178 119 218 145
rect 244 119 284 145
rect 310 119 350 145
rect 376 119 416 145
rect 442 119 482 145
rect 508 119 548 145
rect 574 119 614 145
rect 640 119 680 145
rect 706 119 746 145
rect 772 119 812 145
rect 838 119 878 145
rect 904 119 944 145
rect 970 119 1010 145
rect 1036 119 1076 145
rect 1102 119 1142 145
rect 1168 119 1208 145
rect 1234 119 1274 145
rect 1300 119 1340 145
rect 1366 119 1406 145
rect 1432 119 1472 145
rect 1498 119 1538 145
rect 1564 119 1604 145
rect 1630 119 1636 145
rect -1636 79 1636 119
rect -1636 53 -1630 79
rect -1604 53 -1564 79
rect -1538 53 -1498 79
rect -1472 53 -1432 79
rect -1406 53 -1366 79
rect -1340 53 -1300 79
rect -1274 53 -1234 79
rect -1208 53 -1168 79
rect -1142 53 -1102 79
rect -1076 53 -1036 79
rect -1010 53 -970 79
rect -944 53 -904 79
rect -878 53 -838 79
rect -812 53 -772 79
rect -746 53 -706 79
rect -680 53 -640 79
rect -614 53 -574 79
rect -548 53 -508 79
rect -482 53 -442 79
rect -416 53 -376 79
rect -350 53 -310 79
rect -284 53 -244 79
rect -218 53 -178 79
rect -152 53 -112 79
rect -86 53 -46 79
rect -20 53 20 79
rect 46 53 86 79
rect 112 53 152 79
rect 178 53 218 79
rect 244 53 284 79
rect 310 53 350 79
rect 376 53 416 79
rect 442 53 482 79
rect 508 53 548 79
rect 574 53 614 79
rect 640 53 680 79
rect 706 53 746 79
rect 772 53 812 79
rect 838 53 878 79
rect 904 53 944 79
rect 970 53 1010 79
rect 1036 53 1076 79
rect 1102 53 1142 79
rect 1168 53 1208 79
rect 1234 53 1274 79
rect 1300 53 1340 79
rect 1366 53 1406 79
rect 1432 53 1472 79
rect 1498 53 1538 79
rect 1564 53 1604 79
rect 1630 53 1636 79
rect -1636 13 1636 53
rect -1636 -13 -1630 13
rect -1604 -13 -1564 13
rect -1538 -13 -1498 13
rect -1472 -13 -1432 13
rect -1406 -13 -1366 13
rect -1340 -13 -1300 13
rect -1274 -13 -1234 13
rect -1208 -13 -1168 13
rect -1142 -13 -1102 13
rect -1076 -13 -1036 13
rect -1010 -13 -970 13
rect -944 -13 -904 13
rect -878 -13 -838 13
rect -812 -13 -772 13
rect -746 -13 -706 13
rect -680 -13 -640 13
rect -614 -13 -574 13
rect -548 -13 -508 13
rect -482 -13 -442 13
rect -416 -13 -376 13
rect -350 -13 -310 13
rect -284 -13 -244 13
rect -218 -13 -178 13
rect -152 -13 -112 13
rect -86 -13 -46 13
rect -20 -13 20 13
rect 46 -13 86 13
rect 112 -13 152 13
rect 178 -13 218 13
rect 244 -13 284 13
rect 310 -13 350 13
rect 376 -13 416 13
rect 442 -13 482 13
rect 508 -13 548 13
rect 574 -13 614 13
rect 640 -13 680 13
rect 706 -13 746 13
rect 772 -13 812 13
rect 838 -13 878 13
rect 904 -13 944 13
rect 970 -13 1010 13
rect 1036 -13 1076 13
rect 1102 -13 1142 13
rect 1168 -13 1208 13
rect 1234 -13 1274 13
rect 1300 -13 1340 13
rect 1366 -13 1406 13
rect 1432 -13 1472 13
rect 1498 -13 1538 13
rect 1564 -13 1604 13
rect 1630 -13 1636 13
rect -1636 -53 1636 -13
rect -1636 -79 -1630 -53
rect -1604 -79 -1564 -53
rect -1538 -79 -1498 -53
rect -1472 -79 -1432 -53
rect -1406 -79 -1366 -53
rect -1340 -79 -1300 -53
rect -1274 -79 -1234 -53
rect -1208 -79 -1168 -53
rect -1142 -79 -1102 -53
rect -1076 -79 -1036 -53
rect -1010 -79 -970 -53
rect -944 -79 -904 -53
rect -878 -79 -838 -53
rect -812 -79 -772 -53
rect -746 -79 -706 -53
rect -680 -79 -640 -53
rect -614 -79 -574 -53
rect -548 -79 -508 -53
rect -482 -79 -442 -53
rect -416 -79 -376 -53
rect -350 -79 -310 -53
rect -284 -79 -244 -53
rect -218 -79 -178 -53
rect -152 -79 -112 -53
rect -86 -79 -46 -53
rect -20 -79 20 -53
rect 46 -79 86 -53
rect 112 -79 152 -53
rect 178 -79 218 -53
rect 244 -79 284 -53
rect 310 -79 350 -53
rect 376 -79 416 -53
rect 442 -79 482 -53
rect 508 -79 548 -53
rect 574 -79 614 -53
rect 640 -79 680 -53
rect 706 -79 746 -53
rect 772 -79 812 -53
rect 838 -79 878 -53
rect 904 -79 944 -53
rect 970 -79 1010 -53
rect 1036 -79 1076 -53
rect 1102 -79 1142 -53
rect 1168 -79 1208 -53
rect 1234 -79 1274 -53
rect 1300 -79 1340 -53
rect 1366 -79 1406 -53
rect 1432 -79 1472 -53
rect 1498 -79 1538 -53
rect 1564 -79 1604 -53
rect 1630 -79 1636 -53
rect -1636 -119 1636 -79
rect -1636 -145 -1630 -119
rect -1604 -145 -1564 -119
rect -1538 -145 -1498 -119
rect -1472 -145 -1432 -119
rect -1406 -145 -1366 -119
rect -1340 -145 -1300 -119
rect -1274 -145 -1234 -119
rect -1208 -145 -1168 -119
rect -1142 -145 -1102 -119
rect -1076 -145 -1036 -119
rect -1010 -145 -970 -119
rect -944 -145 -904 -119
rect -878 -145 -838 -119
rect -812 -145 -772 -119
rect -746 -145 -706 -119
rect -680 -145 -640 -119
rect -614 -145 -574 -119
rect -548 -145 -508 -119
rect -482 -145 -442 -119
rect -416 -145 -376 -119
rect -350 -145 -310 -119
rect -284 -145 -244 -119
rect -218 -145 -178 -119
rect -152 -145 -112 -119
rect -86 -145 -46 -119
rect -20 -145 20 -119
rect 46 -145 86 -119
rect 112 -145 152 -119
rect 178 -145 218 -119
rect 244 -145 284 -119
rect 310 -145 350 -119
rect 376 -145 416 -119
rect 442 -145 482 -119
rect 508 -145 548 -119
rect 574 -145 614 -119
rect 640 -145 680 -119
rect 706 -145 746 -119
rect 772 -145 812 -119
rect 838 -145 878 -119
rect 904 -145 944 -119
rect 970 -145 1010 -119
rect 1036 -145 1076 -119
rect 1102 -145 1142 -119
rect 1168 -145 1208 -119
rect 1234 -145 1274 -119
rect 1300 -145 1340 -119
rect 1366 -145 1406 -119
rect 1432 -145 1472 -119
rect 1498 -145 1538 -119
rect 1564 -145 1604 -119
rect 1630 -145 1636 -119
rect -1636 -151 1636 -145
<< via1 >>
rect -1630 119 -1604 145
rect -1564 119 -1538 145
rect -1498 119 -1472 145
rect -1432 119 -1406 145
rect -1366 119 -1340 145
rect -1300 119 -1274 145
rect -1234 119 -1208 145
rect -1168 119 -1142 145
rect -1102 119 -1076 145
rect -1036 119 -1010 145
rect -970 119 -944 145
rect -904 119 -878 145
rect -838 119 -812 145
rect -772 119 -746 145
rect -706 119 -680 145
rect -640 119 -614 145
rect -574 119 -548 145
rect -508 119 -482 145
rect -442 119 -416 145
rect -376 119 -350 145
rect -310 119 -284 145
rect -244 119 -218 145
rect -178 119 -152 145
rect -112 119 -86 145
rect -46 119 -20 145
rect 20 119 46 145
rect 86 119 112 145
rect 152 119 178 145
rect 218 119 244 145
rect 284 119 310 145
rect 350 119 376 145
rect 416 119 442 145
rect 482 119 508 145
rect 548 119 574 145
rect 614 119 640 145
rect 680 119 706 145
rect 746 119 772 145
rect 812 119 838 145
rect 878 119 904 145
rect 944 119 970 145
rect 1010 119 1036 145
rect 1076 119 1102 145
rect 1142 119 1168 145
rect 1208 119 1234 145
rect 1274 119 1300 145
rect 1340 119 1366 145
rect 1406 119 1432 145
rect 1472 119 1498 145
rect 1538 119 1564 145
rect 1604 119 1630 145
rect -1630 53 -1604 79
rect -1564 53 -1538 79
rect -1498 53 -1472 79
rect -1432 53 -1406 79
rect -1366 53 -1340 79
rect -1300 53 -1274 79
rect -1234 53 -1208 79
rect -1168 53 -1142 79
rect -1102 53 -1076 79
rect -1036 53 -1010 79
rect -970 53 -944 79
rect -904 53 -878 79
rect -838 53 -812 79
rect -772 53 -746 79
rect -706 53 -680 79
rect -640 53 -614 79
rect -574 53 -548 79
rect -508 53 -482 79
rect -442 53 -416 79
rect -376 53 -350 79
rect -310 53 -284 79
rect -244 53 -218 79
rect -178 53 -152 79
rect -112 53 -86 79
rect -46 53 -20 79
rect 20 53 46 79
rect 86 53 112 79
rect 152 53 178 79
rect 218 53 244 79
rect 284 53 310 79
rect 350 53 376 79
rect 416 53 442 79
rect 482 53 508 79
rect 548 53 574 79
rect 614 53 640 79
rect 680 53 706 79
rect 746 53 772 79
rect 812 53 838 79
rect 878 53 904 79
rect 944 53 970 79
rect 1010 53 1036 79
rect 1076 53 1102 79
rect 1142 53 1168 79
rect 1208 53 1234 79
rect 1274 53 1300 79
rect 1340 53 1366 79
rect 1406 53 1432 79
rect 1472 53 1498 79
rect 1538 53 1564 79
rect 1604 53 1630 79
rect -1630 -13 -1604 13
rect -1564 -13 -1538 13
rect -1498 -13 -1472 13
rect -1432 -13 -1406 13
rect -1366 -13 -1340 13
rect -1300 -13 -1274 13
rect -1234 -13 -1208 13
rect -1168 -13 -1142 13
rect -1102 -13 -1076 13
rect -1036 -13 -1010 13
rect -970 -13 -944 13
rect -904 -13 -878 13
rect -838 -13 -812 13
rect -772 -13 -746 13
rect -706 -13 -680 13
rect -640 -13 -614 13
rect -574 -13 -548 13
rect -508 -13 -482 13
rect -442 -13 -416 13
rect -376 -13 -350 13
rect -310 -13 -284 13
rect -244 -13 -218 13
rect -178 -13 -152 13
rect -112 -13 -86 13
rect -46 -13 -20 13
rect 20 -13 46 13
rect 86 -13 112 13
rect 152 -13 178 13
rect 218 -13 244 13
rect 284 -13 310 13
rect 350 -13 376 13
rect 416 -13 442 13
rect 482 -13 508 13
rect 548 -13 574 13
rect 614 -13 640 13
rect 680 -13 706 13
rect 746 -13 772 13
rect 812 -13 838 13
rect 878 -13 904 13
rect 944 -13 970 13
rect 1010 -13 1036 13
rect 1076 -13 1102 13
rect 1142 -13 1168 13
rect 1208 -13 1234 13
rect 1274 -13 1300 13
rect 1340 -13 1366 13
rect 1406 -13 1432 13
rect 1472 -13 1498 13
rect 1538 -13 1564 13
rect 1604 -13 1630 13
rect -1630 -79 -1604 -53
rect -1564 -79 -1538 -53
rect -1498 -79 -1472 -53
rect -1432 -79 -1406 -53
rect -1366 -79 -1340 -53
rect -1300 -79 -1274 -53
rect -1234 -79 -1208 -53
rect -1168 -79 -1142 -53
rect -1102 -79 -1076 -53
rect -1036 -79 -1010 -53
rect -970 -79 -944 -53
rect -904 -79 -878 -53
rect -838 -79 -812 -53
rect -772 -79 -746 -53
rect -706 -79 -680 -53
rect -640 -79 -614 -53
rect -574 -79 -548 -53
rect -508 -79 -482 -53
rect -442 -79 -416 -53
rect -376 -79 -350 -53
rect -310 -79 -284 -53
rect -244 -79 -218 -53
rect -178 -79 -152 -53
rect -112 -79 -86 -53
rect -46 -79 -20 -53
rect 20 -79 46 -53
rect 86 -79 112 -53
rect 152 -79 178 -53
rect 218 -79 244 -53
rect 284 -79 310 -53
rect 350 -79 376 -53
rect 416 -79 442 -53
rect 482 -79 508 -53
rect 548 -79 574 -53
rect 614 -79 640 -53
rect 680 -79 706 -53
rect 746 -79 772 -53
rect 812 -79 838 -53
rect 878 -79 904 -53
rect 944 -79 970 -53
rect 1010 -79 1036 -53
rect 1076 -79 1102 -53
rect 1142 -79 1168 -53
rect 1208 -79 1234 -53
rect 1274 -79 1300 -53
rect 1340 -79 1366 -53
rect 1406 -79 1432 -53
rect 1472 -79 1498 -53
rect 1538 -79 1564 -53
rect 1604 -79 1630 -53
rect -1630 -145 -1604 -119
rect -1564 -145 -1538 -119
rect -1498 -145 -1472 -119
rect -1432 -145 -1406 -119
rect -1366 -145 -1340 -119
rect -1300 -145 -1274 -119
rect -1234 -145 -1208 -119
rect -1168 -145 -1142 -119
rect -1102 -145 -1076 -119
rect -1036 -145 -1010 -119
rect -970 -145 -944 -119
rect -904 -145 -878 -119
rect -838 -145 -812 -119
rect -772 -145 -746 -119
rect -706 -145 -680 -119
rect -640 -145 -614 -119
rect -574 -145 -548 -119
rect -508 -145 -482 -119
rect -442 -145 -416 -119
rect -376 -145 -350 -119
rect -310 -145 -284 -119
rect -244 -145 -218 -119
rect -178 -145 -152 -119
rect -112 -145 -86 -119
rect -46 -145 -20 -119
rect 20 -145 46 -119
rect 86 -145 112 -119
rect 152 -145 178 -119
rect 218 -145 244 -119
rect 284 -145 310 -119
rect 350 -145 376 -119
rect 416 -145 442 -119
rect 482 -145 508 -119
rect 548 -145 574 -119
rect 614 -145 640 -119
rect 680 -145 706 -119
rect 746 -145 772 -119
rect 812 -145 838 -119
rect 878 -145 904 -119
rect 944 -145 970 -119
rect 1010 -145 1036 -119
rect 1076 -145 1102 -119
rect 1142 -145 1168 -119
rect 1208 -145 1234 -119
rect 1274 -145 1300 -119
rect 1340 -145 1366 -119
rect 1406 -145 1432 -119
rect 1472 -145 1498 -119
rect 1538 -145 1564 -119
rect 1604 -145 1630 -119
<< metal2 >>
rect -1636 145 1636 151
rect -1636 119 -1630 145
rect -1604 119 -1564 145
rect -1538 119 -1498 145
rect -1472 119 -1432 145
rect -1406 119 -1366 145
rect -1340 119 -1300 145
rect -1274 119 -1234 145
rect -1208 119 -1168 145
rect -1142 119 -1102 145
rect -1076 119 -1036 145
rect -1010 119 -970 145
rect -944 119 -904 145
rect -878 119 -838 145
rect -812 119 -772 145
rect -746 119 -706 145
rect -680 119 -640 145
rect -614 119 -574 145
rect -548 119 -508 145
rect -482 119 -442 145
rect -416 119 -376 145
rect -350 119 -310 145
rect -284 119 -244 145
rect -218 119 -178 145
rect -152 119 -112 145
rect -86 119 -46 145
rect -20 119 20 145
rect 46 119 86 145
rect 112 119 152 145
rect 178 119 218 145
rect 244 119 284 145
rect 310 119 350 145
rect 376 119 416 145
rect 442 119 482 145
rect 508 119 548 145
rect 574 119 614 145
rect 640 119 680 145
rect 706 119 746 145
rect 772 119 812 145
rect 838 119 878 145
rect 904 119 944 145
rect 970 119 1010 145
rect 1036 119 1076 145
rect 1102 119 1142 145
rect 1168 119 1208 145
rect 1234 119 1274 145
rect 1300 119 1340 145
rect 1366 119 1406 145
rect 1432 119 1472 145
rect 1498 119 1538 145
rect 1564 119 1604 145
rect 1630 119 1636 145
rect -1636 79 1636 119
rect -1636 53 -1630 79
rect -1604 53 -1564 79
rect -1538 53 -1498 79
rect -1472 53 -1432 79
rect -1406 53 -1366 79
rect -1340 53 -1300 79
rect -1274 53 -1234 79
rect -1208 53 -1168 79
rect -1142 53 -1102 79
rect -1076 53 -1036 79
rect -1010 53 -970 79
rect -944 53 -904 79
rect -878 53 -838 79
rect -812 53 -772 79
rect -746 53 -706 79
rect -680 53 -640 79
rect -614 53 -574 79
rect -548 53 -508 79
rect -482 53 -442 79
rect -416 53 -376 79
rect -350 53 -310 79
rect -284 53 -244 79
rect -218 53 -178 79
rect -152 53 -112 79
rect -86 53 -46 79
rect -20 53 20 79
rect 46 53 86 79
rect 112 53 152 79
rect 178 53 218 79
rect 244 53 284 79
rect 310 53 350 79
rect 376 53 416 79
rect 442 53 482 79
rect 508 53 548 79
rect 574 53 614 79
rect 640 53 680 79
rect 706 53 746 79
rect 772 53 812 79
rect 838 53 878 79
rect 904 53 944 79
rect 970 53 1010 79
rect 1036 53 1076 79
rect 1102 53 1142 79
rect 1168 53 1208 79
rect 1234 53 1274 79
rect 1300 53 1340 79
rect 1366 53 1406 79
rect 1432 53 1472 79
rect 1498 53 1538 79
rect 1564 53 1604 79
rect 1630 53 1636 79
rect -1636 13 1636 53
rect -1636 -13 -1630 13
rect -1604 -13 -1564 13
rect -1538 -13 -1498 13
rect -1472 -13 -1432 13
rect -1406 -13 -1366 13
rect -1340 -13 -1300 13
rect -1274 -13 -1234 13
rect -1208 -13 -1168 13
rect -1142 -13 -1102 13
rect -1076 -13 -1036 13
rect -1010 -13 -970 13
rect -944 -13 -904 13
rect -878 -13 -838 13
rect -812 -13 -772 13
rect -746 -13 -706 13
rect -680 -13 -640 13
rect -614 -13 -574 13
rect -548 -13 -508 13
rect -482 -13 -442 13
rect -416 -13 -376 13
rect -350 -13 -310 13
rect -284 -13 -244 13
rect -218 -13 -178 13
rect -152 -13 -112 13
rect -86 -13 -46 13
rect -20 -13 20 13
rect 46 -13 86 13
rect 112 -13 152 13
rect 178 -13 218 13
rect 244 -13 284 13
rect 310 -13 350 13
rect 376 -13 416 13
rect 442 -13 482 13
rect 508 -13 548 13
rect 574 -13 614 13
rect 640 -13 680 13
rect 706 -13 746 13
rect 772 -13 812 13
rect 838 -13 878 13
rect 904 -13 944 13
rect 970 -13 1010 13
rect 1036 -13 1076 13
rect 1102 -13 1142 13
rect 1168 -13 1208 13
rect 1234 -13 1274 13
rect 1300 -13 1340 13
rect 1366 -13 1406 13
rect 1432 -13 1472 13
rect 1498 -13 1538 13
rect 1564 -13 1604 13
rect 1630 -13 1636 13
rect -1636 -53 1636 -13
rect -1636 -79 -1630 -53
rect -1604 -79 -1564 -53
rect -1538 -79 -1498 -53
rect -1472 -79 -1432 -53
rect -1406 -79 -1366 -53
rect -1340 -79 -1300 -53
rect -1274 -79 -1234 -53
rect -1208 -79 -1168 -53
rect -1142 -79 -1102 -53
rect -1076 -79 -1036 -53
rect -1010 -79 -970 -53
rect -944 -79 -904 -53
rect -878 -79 -838 -53
rect -812 -79 -772 -53
rect -746 -79 -706 -53
rect -680 -79 -640 -53
rect -614 -79 -574 -53
rect -548 -79 -508 -53
rect -482 -79 -442 -53
rect -416 -79 -376 -53
rect -350 -79 -310 -53
rect -284 -79 -244 -53
rect -218 -79 -178 -53
rect -152 -79 -112 -53
rect -86 -79 -46 -53
rect -20 -79 20 -53
rect 46 -79 86 -53
rect 112 -79 152 -53
rect 178 -79 218 -53
rect 244 -79 284 -53
rect 310 -79 350 -53
rect 376 -79 416 -53
rect 442 -79 482 -53
rect 508 -79 548 -53
rect 574 -79 614 -53
rect 640 -79 680 -53
rect 706 -79 746 -53
rect 772 -79 812 -53
rect 838 -79 878 -53
rect 904 -79 944 -53
rect 970 -79 1010 -53
rect 1036 -79 1076 -53
rect 1102 -79 1142 -53
rect 1168 -79 1208 -53
rect 1234 -79 1274 -53
rect 1300 -79 1340 -53
rect 1366 -79 1406 -53
rect 1432 -79 1472 -53
rect 1498 -79 1538 -53
rect 1564 -79 1604 -53
rect 1630 -79 1636 -53
rect -1636 -119 1636 -79
rect -1636 -145 -1630 -119
rect -1604 -145 -1564 -119
rect -1538 -145 -1498 -119
rect -1472 -145 -1432 -119
rect -1406 -145 -1366 -119
rect -1340 -145 -1300 -119
rect -1274 -145 -1234 -119
rect -1208 -145 -1168 -119
rect -1142 -145 -1102 -119
rect -1076 -145 -1036 -119
rect -1010 -145 -970 -119
rect -944 -145 -904 -119
rect -878 -145 -838 -119
rect -812 -145 -772 -119
rect -746 -145 -706 -119
rect -680 -145 -640 -119
rect -614 -145 -574 -119
rect -548 -145 -508 -119
rect -482 -145 -442 -119
rect -416 -145 -376 -119
rect -350 -145 -310 -119
rect -284 -145 -244 -119
rect -218 -145 -178 -119
rect -152 -145 -112 -119
rect -86 -145 -46 -119
rect -20 -145 20 -119
rect 46 -145 86 -119
rect 112 -145 152 -119
rect 178 -145 218 -119
rect 244 -145 284 -119
rect 310 -145 350 -119
rect 376 -145 416 -119
rect 442 -145 482 -119
rect 508 -145 548 -119
rect 574 -145 614 -119
rect 640 -145 680 -119
rect 706 -145 746 -119
rect 772 -145 812 -119
rect 838 -145 878 -119
rect 904 -145 944 -119
rect 970 -145 1010 -119
rect 1036 -145 1076 -119
rect 1102 -145 1142 -119
rect 1168 -145 1208 -119
rect 1234 -145 1274 -119
rect 1300 -145 1340 -119
rect 1366 -145 1406 -119
rect 1432 -145 1472 -119
rect 1498 -145 1538 -119
rect 1564 -145 1604 -119
rect 1630 -145 1636 -119
rect -1636 -151 1636 -145
<< end >>
