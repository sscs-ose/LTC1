magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2042 -2089 2042 2089
<< polysilicon >>
rect -42 70 42 89
rect -42 -70 -23 70
rect 23 -70 42 70
rect -42 -89 42 -70
<< polycontact >>
rect -23 -70 23 70
<< metal1 >>
rect -34 70 34 81
rect -34 -70 -23 70
rect 23 -70 34 70
rect -34 -81 34 -70
<< end >>
