magic
tech gf180mcuC
magscale 1 10
timestamp 1694765517
<< metal1 >>
rect 56075 46987 67056 47998
rect 59407 41842 59720 46987
rect 58483 41792 59720 41842
rect 58483 41693 59368 41792
rect 59635 41693 59720 41792
rect 58483 41666 59720 41693
rect 58483 41662 59409 41666
rect 59540 41662 59718 41666
rect 55974 21282 56130 39904
rect 59223 27012 59786 27051
rect 58616 26694 59037 26872
rect 59223 26834 59324 27012
rect 59718 26834 59786 27012
rect 59223 26777 59786 26834
rect 64823 25513 66673 25694
rect 64823 25415 65004 25513
rect 66328 25271 66428 25363
rect 65883 25176 65977 25184
rect 65883 25122 65896 25176
rect 65962 25172 65977 25176
rect 65962 25122 66376 25172
rect 65883 25120 66376 25122
rect 65883 25115 65977 25120
rect 58166 24948 58331 25024
rect 65878 24948 65972 24956
rect 58166 24898 58591 24948
rect 65878 24947 65888 24948
rect 58166 24847 58331 24898
rect 65373 24896 65888 24947
rect 65958 24896 65972 24948
rect 65373 24895 65972 24896
rect 65878 24887 65972 24895
rect 66328 24854 66430 24951
rect 65881 24764 65958 24770
rect 65881 24712 65894 24764
rect 65946 24762 65958 24764
rect 65946 24712 66423 24762
rect 65881 24710 66423 24712
rect 65881 24698 65958 24710
rect 65283 24373 68806 24641
rect 65271 23577 65681 23614
rect 65271 23406 65582 23577
rect 65660 23406 65681 23577
rect 65271 23342 65681 23406
rect 57645 23078 58421 23080
rect 57645 23028 58501 23078
rect 57645 22966 58421 23028
rect 68929 23004 69086 23093
rect 68932 22987 69086 23004
rect 55926 21206 56211 21282
rect 55926 21052 55993 21206
rect 56135 21052 56211 21206
rect 55926 20990 56211 21052
rect 57645 10767 57832 22966
rect 65874 22911 65960 22913
rect 65874 22899 65961 22911
rect 65874 22898 65887 22899
rect 65448 22846 65887 22898
rect 65874 22844 65887 22846
rect 65950 22844 65961 22899
rect 65874 22830 65961 22844
rect 65545 22769 65691 22778
rect 65545 22753 66351 22769
rect 65545 22629 65569 22753
rect 65676 22629 66351 22753
rect 65545 22624 66351 22629
rect 65545 22609 65691 22624
rect 69190 22623 69320 22637
rect 69190 22616 69203 22623
rect 68924 22546 69203 22616
rect 69305 22546 69320 22623
rect 68924 22540 69320 22546
rect 69190 22530 69320 22540
rect 69070 22137 69193 22153
rect 69070 22127 69086 22137
rect 69057 22124 69086 22127
rect 68844 22065 69086 22124
rect 69180 22065 69193 22137
rect 68844 22056 69193 22065
rect 69070 22052 69193 22056
rect 60529 20706 60919 21748
rect 65096 21359 66157 21748
rect 58050 20607 58267 20649
rect 58050 20453 58083 20607
rect 58234 20453 58267 20607
rect 58675 20566 58829 20589
rect 58675 20509 58700 20566
rect 58788 20509 58829 20566
rect 58675 20476 58829 20509
rect 58050 20420 58267 20453
rect 58040 18703 58248 18758
rect 58040 18600 58099 18703
rect 58197 18600 58248 18703
rect 58040 18556 58248 18600
rect 59369 17342 59499 17350
rect 58258 17317 59499 17342
rect 58258 17190 59389 17317
rect 59474 17190 59499 17317
rect 58258 17182 59499 17190
rect 59369 17169 59499 17182
rect 67600 17222 68729 17233
rect 67600 17154 67618 17222
rect 67676 17154 68729 17222
rect 67600 17141 68729 17154
rect 62603 17034 62708 17055
rect 62603 16969 62624 17034
rect 62689 16969 62708 17034
rect 62603 16950 62708 16969
rect 64509 17042 64600 17054
rect 64509 16972 64519 17042
rect 64587 16972 64600 17042
rect 64509 16963 64600 16972
rect 57973 16271 58167 16307
rect 57973 16175 58028 16271
rect 58125 16175 58167 16271
rect 57973 16131 58167 16175
rect 58906 16153 59007 16288
rect 57619 10738 57864 10767
rect 57619 10597 57647 10738
rect 57837 10597 57864 10738
rect 57619 10576 57864 10597
rect 58005 9460 58154 16131
rect 62571 13175 62900 13811
rect 68812 13643 68942 13675
rect 68812 13575 68839 13643
rect 68913 13575 68942 13643
rect 68812 13549 68942 13575
rect 58575 10663 58653 10675
rect 58575 10601 58587 10663
rect 58642 10601 58653 10663
rect 58575 10590 58653 10601
rect 57985 9436 58197 9460
rect 57985 9315 58012 9436
rect 58171 9315 58197 9436
rect 57985 9288 58197 9315
rect 59580 7678 59748 7700
rect 59580 7599 59609 7678
rect 59717 7599 59748 7678
rect 59580 7580 59748 7599
rect 56871 1165 70990 1240
rect 56871 1086 59614 1165
rect 59722 1086 70990 1165
rect 56871 450 70990 1086
<< via1 >>
rect 59368 41693 59635 41792
rect 59324 26834 59718 27012
rect 65896 25122 65962 25176
rect 65888 24896 65958 24948
rect 65894 24712 65946 24764
rect 65582 23406 65660 23577
rect 55993 21052 56135 21206
rect 65887 22844 65950 22899
rect 65569 22629 65676 22753
rect 69203 22546 69305 22623
rect 69086 22065 69180 22137
rect 58083 20453 58234 20607
rect 58700 20509 58788 20566
rect 58099 18600 58197 18703
rect 59389 17190 59474 17317
rect 67618 17154 67676 17222
rect 62624 16969 62689 17034
rect 64519 16972 64587 17042
rect 58028 16175 58125 16271
rect 57647 10597 57837 10738
rect 68839 13575 68913 13643
rect 58614 12215 58685 12286
rect 58587 10601 58642 10663
rect 58012 9315 58171 9436
rect 59609 7599 59717 7678
rect 59614 1086 59722 1165
<< metal2 >>
rect 59325 41792 59670 41815
rect 59325 41693 59368 41792
rect 59635 41693 59670 41792
rect 59325 27051 59670 41693
rect 59223 27012 59786 27051
rect 59223 26966 59324 27012
rect 56398 26843 59324 26966
rect 55926 21240 56211 21282
rect 55926 21018 55960 21240
rect 56177 21018 56211 21240
rect 55926 20990 56211 21018
rect 56398 12311 56521 26843
rect 58616 26694 59037 26843
rect 59223 26834 59324 26843
rect 59718 26834 59786 27012
rect 59223 26777 59786 26834
rect 68725 25289 69297 25293
rect 68725 25221 69308 25289
rect 65883 25176 65977 25184
rect 65883 25122 65896 25176
rect 65962 25122 65977 25176
rect 65883 25115 65977 25122
rect 65891 24956 65962 25115
rect 65878 24948 65972 24956
rect 65878 24896 65888 24948
rect 65958 24896 65972 24948
rect 65878 24887 65972 24896
rect 65881 24764 65958 24770
rect 65881 24712 65894 24764
rect 65946 24712 65958 24764
rect 65881 24698 65958 24712
rect 65560 23577 65681 23614
rect 65560 23406 65582 23577
rect 65660 23406 65681 23577
rect 65560 22778 65681 23406
rect 65890 22913 65951 24698
rect 65874 22911 65960 22913
rect 65874 22899 65961 22911
rect 65874 22844 65887 22899
rect 65950 22844 65961 22899
rect 65874 22830 65961 22844
rect 65545 22753 65691 22778
rect 65545 22629 65569 22753
rect 65676 22629 65691 22753
rect 69200 22637 69308 25221
rect 65545 22609 65691 22629
rect 69190 22632 69320 22637
rect 69190 22623 69406 22632
rect 69190 22546 69203 22623
rect 69305 22546 69406 22623
rect 69190 22530 69406 22546
rect 69070 22137 69193 22153
rect 69070 22065 69086 22137
rect 69180 22065 69193 22137
rect 69070 22052 69193 22065
rect 69080 21250 69191 22052
rect 69070 21216 69203 21250
rect 69070 21052 69096 21216
rect 69179 21052 69203 21216
rect 69070 21014 69203 21052
rect 58050 20621 58267 20649
rect 58050 20444 58066 20621
rect 58246 20444 58267 20621
rect 58675 20576 58829 20589
rect 58675 20490 58689 20576
rect 58809 20490 58829 20576
rect 58675 20476 58829 20490
rect 58050 20420 58267 20444
rect 69302 18853 69406 22530
rect 69289 18835 69427 18853
rect 58040 18732 58248 18758
rect 58040 18582 58072 18732
rect 58218 18582 58248 18732
rect 69289 18708 69309 18835
rect 69414 18708 69427 18835
rect 69289 18688 69427 18708
rect 58040 18556 58248 18582
rect 59369 17317 59499 17350
rect 59369 17190 59389 17317
rect 59474 17190 59499 17317
rect 59369 17169 59499 17190
rect 67608 17222 67700 17234
rect 67608 17154 67618 17222
rect 67676 17154 67700 17222
rect 67608 17142 67700 17154
rect 62603 17034 62708 17055
rect 62603 16969 62624 17034
rect 62689 16969 62708 17034
rect 62603 16950 62708 16969
rect 64509 17042 64600 17054
rect 64509 16972 64519 17042
rect 64587 16972 64600 17042
rect 64509 16963 64600 16972
rect 57973 16287 58167 16307
rect 57973 16153 57998 16287
rect 58146 16153 58167 16287
rect 58906 16256 59007 16288
rect 58906 16176 58925 16256
rect 58987 16176 59007 16256
rect 58906 16153 59007 16176
rect 57973 16131 58167 16153
rect 68812 13662 68942 13675
rect 68812 13571 68824 13662
rect 68928 13571 68942 13662
rect 68812 13549 68942 13571
rect 56398 12286 58706 12311
rect 56398 12215 58614 12286
rect 58685 12215 58706 12286
rect 56398 12188 58706 12215
rect 57619 10738 57864 10767
rect 57619 10597 57647 10738
rect 57837 10668 57864 10738
rect 58575 10668 58653 10675
rect 57837 10663 58653 10668
rect 57837 10601 58587 10663
rect 58642 10601 58653 10663
rect 57837 10597 58653 10601
rect 57619 10596 58653 10597
rect 57619 10576 57864 10596
rect 58575 10590 58653 10596
rect 57985 9436 58197 9460
rect 57985 9315 58012 9436
rect 58171 9381 58197 9436
rect 58171 9324 58810 9381
rect 58171 9315 58197 9324
rect 57985 9288 58197 9315
rect 59580 7678 59902 7700
rect 59580 7599 59609 7678
rect 59717 7599 59902 7678
rect 59580 7554 59902 7599
rect 59590 1395 59901 7554
rect 59590 1235 59904 1395
rect 59565 1165 59904 1235
rect 59565 1086 59614 1165
rect 59722 1086 59904 1165
rect 59565 1085 59904 1086
rect 59590 1050 59740 1085
<< via2 >>
rect 55960 21206 56177 21240
rect 55960 21052 55993 21206
rect 55993 21052 56135 21206
rect 56135 21052 56177 21206
rect 55960 21018 56177 21052
rect 69096 21052 69179 21216
rect 58066 20607 58246 20621
rect 58066 20453 58083 20607
rect 58083 20453 58234 20607
rect 58234 20453 58246 20607
rect 58066 20444 58246 20453
rect 58689 20566 58809 20576
rect 58689 20509 58700 20566
rect 58700 20509 58788 20566
rect 58788 20509 58809 20566
rect 58689 20490 58809 20509
rect 58072 18703 58218 18732
rect 58072 18600 58099 18703
rect 58099 18600 58197 18703
rect 58197 18600 58218 18703
rect 58072 18582 58218 18600
rect 69309 18708 69414 18835
rect 59389 17190 59474 17317
rect 67618 17154 67676 17222
rect 62624 16969 62689 17034
rect 64519 16972 64587 17042
rect 57998 16271 58146 16287
rect 57998 16175 58028 16271
rect 58028 16175 58125 16271
rect 58125 16175 58146 16271
rect 57998 16153 58146 16175
rect 58925 16176 58987 16256
rect 68824 13643 68928 13662
rect 68824 13575 68839 13643
rect 68839 13575 68913 13643
rect 68913 13575 68928 13643
rect 68824 13571 68928 13575
<< metal3 >>
rect 55926 21240 56211 21282
rect 69070 21242 69203 21250
rect 55926 21018 55960 21240
rect 56177 21239 56211 21240
rect 69057 21239 69203 21242
rect 56177 21216 69203 21239
rect 56177 21052 69096 21216
rect 69179 21052 69203 21216
rect 56177 21018 69203 21052
rect 55926 21014 69203 21018
rect 55926 20990 56211 21014
rect 58050 20621 58267 20649
rect 58050 20444 58066 20621
rect 58246 20589 58267 20621
rect 58246 20576 58828 20589
rect 58246 20490 58689 20576
rect 58809 20490 58828 20576
rect 58246 20472 58828 20490
rect 58246 20444 58267 20472
rect 58050 20420 58267 20444
rect 69289 18837 69427 18853
rect 67744 18835 69427 18837
rect 58040 18732 58248 18758
rect 58040 18582 58072 18732
rect 58218 18721 58248 18732
rect 58218 18582 59208 18721
rect 67744 18708 69309 18835
rect 69414 18708 69427 18835
rect 67744 18703 69427 18708
rect 69289 18688 69427 18703
rect 58040 18579 59208 18582
rect 58040 18556 58248 18579
rect 59066 18495 59208 18579
rect 59369 17317 59499 17350
rect 59369 17190 59389 17317
rect 59474 17316 59499 17317
rect 59474 17211 62347 17316
rect 59474 17190 59499 17211
rect 59369 17169 59499 17190
rect 62242 17055 62347 17211
rect 64601 17222 67686 17232
rect 64601 17154 67618 17222
rect 67676 17154 67686 17222
rect 64601 17143 67686 17154
rect 64601 17055 64690 17143
rect 62242 17034 62708 17055
rect 64521 17054 64690 17055
rect 62242 16969 62624 17034
rect 62689 16969 62708 17034
rect 62242 16950 62708 16969
rect 64509 17042 64690 17054
rect 64509 16972 64519 17042
rect 64587 16972 64690 17042
rect 64509 16966 64690 16972
rect 64509 16963 64600 16966
rect 57973 16291 58167 16307
rect 57973 16289 58986 16291
rect 57973 16288 59006 16289
rect 57973 16287 59007 16288
rect 57973 16153 57998 16287
rect 58146 16256 59007 16287
rect 58146 16176 58925 16256
rect 58987 16176 59007 16256
rect 58146 16153 59007 16176
rect 57973 16152 59006 16153
rect 57973 16131 58167 16152
rect 68810 13662 68943 13679
rect 68810 13571 68824 13662
rect 68928 13571 68943 13662
rect 68810 13539 68943 13571
rect 68833 12601 68910 13539
use a2x1mux_mag  a2x1mux_mag_0
timestamp 1694760847
transform 1 0 66622 0 1 22687
box -615 -1160 2414 924
use CLK_div_100_mag  CLK_div_100_mag_0
timestamp 1694693600
transform 1 0 58542 0 1 7660
box -125 0 12197 5567
use CP_mag  CP_mag_0
timestamp 1694750549
transform 1 0 66253 0 1 23857
box 76 665 2629 1837
use LF_mag  LF_mag_0
timestamp 1694765517
transform 1 0 10937 0 1 291
box -85 43 54977 46220
use PFD_layout  PFD_layout_0
timestamp 1694755381
transform 1 0 58974 0 1 21506
box -555 -148 6587 5567
<< labels >>
flabel via2 58142 18646 58142 18646 0 FreeSans 1600 0 0 0 EN
port 0 nsew
flabel via2 58149 20529 58149 20529 0 FreeSans 1600 0 0 0 VDD_VCO
port 2 nsew
flabel metal1 58241 24941 58241 24941 0 FreeSans 1600 0 0 0 Vref
port 3 nsew
flabel metal1 66339 25284 66339 25284 0 FreeSans 1600 0 0 0 IPD_
port 4 nsew
flabel metal1 66336 24875 66336 24875 0 FreeSans 1600 0 0 0 IPD+
port 5 nsew
flabel metal1 69049 23035 69049 23035 0 FreeSans 1600 0 0 0 LP_ext
port 6 nsew
flabel via2 68871 13612 68871 13612 0 FreeSans 1600 0 0 0 RST_DIV
port 7 nsew
flabel metal1 65648 24927 65648 24927 0 FreeSans 800 0 0 0 pu
port 9 nsew
flabel metal1 66023 24730 66023 24730 0 FreeSans 800 0 0 0 pd
port 10 nsew
flabel metal1 63232 703 63232 703 0 FreeSans 1600 0 0 0 VSS
port 11 nsew
flabel metal1 61439 47505 61439 47505 0 FreeSans 1600 0 0 0 VDD
port 12 nsew
flabel metal1 68680 17189 68680 17189 0 FreeSans 1600 0 0 0 VCO_op
port 14 nsew
flabel metal1 58326 17258 58326 17258 0 FreeSans 1600 0 0 0 VCO_op_bar
port 15 nsew
<< end >>
