magic
tech gf180mcuD
magscale 1 10
timestamp 1713866589
<< error_p >>
rect 77983 453525 77993 453535
rect 78106 453525 78116 453535
rect 77973 453515 77983 453525
rect 78116 453515 78126 453525
rect 77973 453392 77983 453402
rect 78116 453392 78126 453402
rect 77983 453382 77993 453392
rect 78106 453382 78116 453392
rect 126959 453359 126960 453369
rect 78123 453263 78124 453273
rect 78123 453140 78124 453150
rect 77991 452882 78001 452892
rect 78114 452882 78124 452892
rect 77981 452872 77991 452882
rect 78124 452872 78134 452882
rect 77981 452749 77991 452759
rect 78124 452749 78134 452759
rect 77991 452739 78001 452749
rect 78114 452739 78124 452749
rect 126959 452148 126960 452158
rect 126959 447184 126960 447194
rect 126959 445973 126960 445983
rect 126940 445963 126950 445964
<< error_s >>
rect 75060 577769 75113 577963
rect 75060 521247 75113 577761
rect 81937 577198 82064 577281
rect 93054 577198 93182 577281
rect 141937 577228 142064 577311
rect 153054 577228 153182 577311
rect 161937 577228 162064 577311
rect 173054 577228 173182 577311
rect 82023 576797 82024 577198
rect 82064 576797 93054 577198
rect 93096 576797 93182 577198
rect 142023 576827 142024 577228
rect 142064 576827 153054 577228
rect 153096 576827 153182 577228
rect 142023 576826 153182 576827
rect 162023 576827 162024 577228
rect 162064 576827 173054 577228
rect 173096 576827 173182 577228
rect 162023 576826 173182 576827
rect 82023 576796 93182 576797
rect 141937 567231 142023 567234
rect 153096 567231 153182 567234
rect 81937 567201 82023 567204
rect 93096 567201 93182 567204
rect 81937 567118 82118 567201
rect 93000 567118 93182 567201
rect 141937 567148 142118 567231
rect 153000 567148 153182 567231
rect 161937 567231 162023 567234
rect 173096 567231 173182 567234
rect 161937 567148 162118 567231
rect 173000 567148 173182 567231
rect 82023 566301 82024 567118
rect 82032 566301 82118 567118
rect 82023 566300 82118 566301
rect 93086 566300 93182 567118
rect 142023 566331 142024 567148
rect 142032 566331 142118 567148
rect 142023 566330 142118 566331
rect 153086 566330 153182 567148
rect 162023 566331 162024 567148
rect 162032 566331 162118 567148
rect 162023 566330 162118 566331
rect 173086 566330 173182 567148
rect 142338 561964 142377 561966
rect 142517 561964 142549 561966
rect 143724 561964 143761 561966
rect 143901 561964 143935 561966
rect 144111 561964 144145 561966
rect 144285 561964 144322 561966
rect 145490 561964 145529 561966
rect 145669 561964 145701 561966
rect 145877 561964 145913 561966
rect 146053 561964 146088 561966
rect 147259 561964 147297 561966
rect 147437 561964 147470 561966
rect 147647 561964 147681 561966
rect 147821 561964 147858 561966
rect 149028 561964 149065 561966
rect 149205 561964 149239 561966
rect 149419 561964 149449 561966
rect 149589 561964 149630 561966
rect 150793 561964 150833 561966
rect 150973 561964 151004 561966
rect 151179 561964 151217 561966
rect 151357 561964 151390 561966
rect 152565 561964 152601 561966
rect 152741 561964 152776 561966
rect 162338 561964 162377 561966
rect 162517 561964 162549 561966
rect 163724 561964 163761 561966
rect 163901 561964 163935 561966
rect 164111 561964 164145 561966
rect 164285 561964 164322 561966
rect 165490 561964 165529 561966
rect 165669 561964 165701 561966
rect 165877 561964 165913 561966
rect 166053 561964 166088 561966
rect 167259 561964 167297 561966
rect 167437 561964 167470 561966
rect 167647 561964 167681 561966
rect 167821 561964 167858 561966
rect 169028 561964 169065 561966
rect 169205 561964 169239 561966
rect 169419 561964 169449 561966
rect 169589 561964 169630 561966
rect 170793 561964 170833 561966
rect 170973 561964 171004 561966
rect 171179 561964 171217 561966
rect 171357 561964 171390 561966
rect 172565 561964 172601 561966
rect 172741 561964 172776 561966
rect 82338 561934 82377 561936
rect 82517 561934 82549 561936
rect 83724 561934 83761 561936
rect 83901 561934 83935 561936
rect 84111 561934 84145 561936
rect 84285 561934 84322 561936
rect 85490 561934 85529 561936
rect 85669 561934 85701 561936
rect 85877 561934 85913 561936
rect 86053 561934 86088 561936
rect 87259 561934 87297 561936
rect 87437 561934 87470 561936
rect 87647 561934 87681 561936
rect 87821 561934 87858 561936
rect 89028 561934 89065 561936
rect 89205 561934 89239 561936
rect 89419 561934 89449 561936
rect 89589 561934 89630 561936
rect 90793 561934 90833 561936
rect 90973 561934 91004 561936
rect 91179 561934 91217 561936
rect 91357 561934 91390 561936
rect 92565 561934 92601 561936
rect 92741 561934 92776 561936
rect 142321 561874 142377 561876
rect 142517 561874 142639 561876
rect 143634 561874 143761 561876
rect 143901 561874 143957 561876
rect 144089 561874 144145 561876
rect 144285 561874 144412 561876
rect 145400 561874 145529 561876
rect 145669 561874 145725 561876
rect 145857 561874 145913 561876
rect 146053 561874 146178 561876
rect 147169 561874 147297 561876
rect 147437 561874 147493 561876
rect 147625 561874 147681 561876
rect 147821 561874 147948 561876
rect 148938 561874 149065 561876
rect 149205 561874 149261 561876
rect 149393 561874 149449 561876
rect 149589 561874 149720 561876
rect 150703 561874 150833 561876
rect 150973 561874 151029 561876
rect 151161 561874 151217 561876
rect 151357 561874 151480 561876
rect 152475 561874 152601 561876
rect 152741 561874 152797 561876
rect 162321 561874 162377 561876
rect 162517 561874 162639 561876
rect 163634 561874 163761 561876
rect 163901 561874 163957 561876
rect 164089 561874 164145 561876
rect 164285 561874 164412 561876
rect 165400 561874 165529 561876
rect 165669 561874 165725 561876
rect 165857 561874 165913 561876
rect 166053 561874 166178 561876
rect 167169 561874 167297 561876
rect 167437 561874 167493 561876
rect 167625 561874 167681 561876
rect 167821 561874 167948 561876
rect 168938 561874 169065 561876
rect 169205 561874 169261 561876
rect 169393 561874 169449 561876
rect 169589 561874 169720 561876
rect 170703 561874 170833 561876
rect 170973 561874 171029 561876
rect 171161 561874 171217 561876
rect 171357 561874 171480 561876
rect 172475 561874 172601 561876
rect 172741 561874 172797 561876
rect 82321 561844 82377 561846
rect 82517 561844 82639 561846
rect 83634 561844 83761 561846
rect 83901 561844 83957 561846
rect 84089 561844 84145 561846
rect 84285 561844 84412 561846
rect 85400 561844 85529 561846
rect 85669 561844 85725 561846
rect 85857 561844 85913 561846
rect 86053 561844 86178 561846
rect 87169 561844 87297 561846
rect 87437 561844 87493 561846
rect 87625 561844 87681 561846
rect 87821 561844 87948 561846
rect 88938 561844 89065 561846
rect 89205 561844 89261 561846
rect 89393 561844 89449 561846
rect 89589 561844 89720 561846
rect 90703 561844 90833 561846
rect 90973 561844 91029 561846
rect 91161 561844 91217 561846
rect 91357 561844 91480 561846
rect 92475 561844 92601 561846
rect 92741 561844 92797 561846
rect 142321 553876 142377 553878
rect 142517 553876 142639 553878
rect 143634 553876 143761 553878
rect 143901 553876 143957 553878
rect 144089 553876 144145 553878
rect 144285 553876 144412 553878
rect 145400 553876 145529 553878
rect 145669 553876 145725 553878
rect 145857 553876 145913 553878
rect 146053 553876 146178 553878
rect 147169 553876 147297 553878
rect 147437 553876 147493 553878
rect 147625 553876 147681 553878
rect 147821 553876 147948 553878
rect 148938 553876 149065 553878
rect 149205 553876 149261 553878
rect 149393 553876 149449 553878
rect 149589 553876 149720 553878
rect 150703 553876 150833 553878
rect 150973 553876 151029 553878
rect 151161 553876 151217 553878
rect 151357 553876 151480 553878
rect 152475 553876 152601 553878
rect 152741 553876 152797 553878
rect 162321 553876 162377 553878
rect 162517 553876 162639 553878
rect 163634 553876 163761 553878
rect 163901 553876 163957 553878
rect 164089 553876 164145 553878
rect 164285 553876 164412 553878
rect 165400 553876 165529 553878
rect 165669 553876 165725 553878
rect 165857 553876 165913 553878
rect 166053 553876 166178 553878
rect 167169 553876 167297 553878
rect 167437 553876 167493 553878
rect 167625 553876 167681 553878
rect 167821 553876 167948 553878
rect 168938 553876 169065 553878
rect 169205 553876 169261 553878
rect 169393 553876 169449 553878
rect 169589 553876 169720 553878
rect 170703 553876 170833 553878
rect 170973 553876 171029 553878
rect 171161 553876 171217 553878
rect 171357 553876 171480 553878
rect 172475 553876 172601 553878
rect 172741 553876 172797 553878
rect 82321 553846 82377 553848
rect 82517 553846 82639 553848
rect 83634 553846 83761 553848
rect 83901 553846 83957 553848
rect 84089 553846 84145 553848
rect 84285 553846 84412 553848
rect 85400 553846 85529 553848
rect 85669 553846 85725 553848
rect 85857 553846 85913 553848
rect 86053 553846 86178 553848
rect 87169 553846 87297 553848
rect 87437 553846 87493 553848
rect 87625 553846 87681 553848
rect 87821 553846 87948 553848
rect 88938 553846 89065 553848
rect 89205 553846 89261 553848
rect 89393 553846 89449 553848
rect 89589 553846 89720 553848
rect 90703 553846 90833 553848
rect 90973 553846 91029 553848
rect 91161 553846 91217 553848
rect 91357 553846 91480 553848
rect 92475 553846 92601 553848
rect 92741 553846 92797 553848
rect 142338 553786 142377 553788
rect 142517 553786 142549 553788
rect 143724 553786 143761 553788
rect 143901 553786 143935 553788
rect 144111 553786 144145 553788
rect 144285 553786 144322 553788
rect 145490 553786 145529 553788
rect 145669 553786 145701 553788
rect 145877 553786 145913 553788
rect 146053 553786 146088 553788
rect 147259 553786 147297 553788
rect 147437 553786 147470 553788
rect 147647 553786 147681 553788
rect 147821 553786 147858 553788
rect 149028 553786 149065 553788
rect 149205 553786 149239 553788
rect 149419 553786 149449 553788
rect 149589 553786 149630 553788
rect 150793 553786 150833 553788
rect 150973 553786 151004 553788
rect 151179 553786 151217 553788
rect 151357 553786 151390 553788
rect 152565 553786 152601 553788
rect 152741 553786 152776 553788
rect 162338 553786 162377 553788
rect 162517 553786 162549 553788
rect 163724 553786 163761 553788
rect 163901 553786 163935 553788
rect 164111 553786 164145 553788
rect 164285 553786 164322 553788
rect 165490 553786 165529 553788
rect 165669 553786 165701 553788
rect 165877 553786 165913 553788
rect 166053 553786 166088 553788
rect 167259 553786 167297 553788
rect 167437 553786 167470 553788
rect 167647 553786 167681 553788
rect 167821 553786 167858 553788
rect 169028 553786 169065 553788
rect 169205 553786 169239 553788
rect 169419 553786 169449 553788
rect 169589 553786 169630 553788
rect 170793 553786 170833 553788
rect 170973 553786 171004 553788
rect 171179 553786 171217 553788
rect 171357 553786 171390 553788
rect 172565 553786 172601 553788
rect 172741 553786 172776 553788
rect 82338 553756 82377 553758
rect 82517 553756 82549 553758
rect 83724 553756 83761 553758
rect 83901 553756 83935 553758
rect 84111 553756 84145 553758
rect 84285 553756 84322 553758
rect 85490 553756 85529 553758
rect 85669 553756 85701 553758
rect 85877 553756 85913 553758
rect 86053 553756 86088 553758
rect 87259 553756 87297 553758
rect 87437 553756 87470 553758
rect 87647 553756 87681 553758
rect 87821 553756 87858 553758
rect 89028 553756 89065 553758
rect 89205 553756 89239 553758
rect 89419 553756 89449 553758
rect 89589 553756 89630 553758
rect 90793 553756 90833 553758
rect 90973 553756 91004 553758
rect 91179 553756 91217 553758
rect 91357 553756 91390 553758
rect 92565 553756 92601 553758
rect 92741 553756 92776 553758
rect 81314 548328 81322 548360
rect 86790 548328 86798 548360
rect 88322 548328 88330 548360
rect 93798 548328 93806 548360
rect 141314 548358 141322 548390
rect 146790 548358 146798 548390
rect 148322 548358 148330 548390
rect 153798 548358 153806 548390
rect 161314 548358 161322 548390
rect 166790 548358 166798 548390
rect 168322 548358 168330 548390
rect 173798 548358 173806 548390
rect 80754 548268 81802 548328
rect 80754 545988 81314 548268
rect 81322 545988 81802 548268
rect 86310 548268 87358 548328
rect 83792 545990 83844 547602
rect 84268 545990 84320 547602
rect 80754 545928 81802 545988
rect 86310 545988 86790 548268
rect 86798 545988 87358 548268
rect 86310 545928 87358 545988
rect 87762 548268 88810 548328
rect 87762 545988 88322 548268
rect 88330 545988 88810 548268
rect 93318 548268 94366 548328
rect 90800 545990 90852 547602
rect 91276 545990 91328 547602
rect 87762 545928 88810 545988
rect 93318 545988 93798 548268
rect 93806 545988 94366 548268
rect 93318 545928 94366 545988
rect 140754 548298 141802 548358
rect 140754 546018 141314 548298
rect 141322 546018 141802 548298
rect 146310 548298 147358 548358
rect 143792 546020 143844 547632
rect 144268 546020 144320 547632
rect 140754 545958 141802 546018
rect 146310 546018 146790 548298
rect 146798 546018 147358 548298
rect 146310 545958 147358 546018
rect 147762 548298 148810 548358
rect 147762 546018 148322 548298
rect 148330 546018 148810 548298
rect 153318 548298 154366 548358
rect 150800 546020 150852 547632
rect 151276 546020 151328 547632
rect 147762 545958 148810 546018
rect 153318 546018 153798 548298
rect 153806 546018 154366 548298
rect 153318 545958 154366 546018
rect 160754 548298 161802 548358
rect 160754 546018 161314 548298
rect 161322 546018 161802 548298
rect 166310 548298 167358 548358
rect 163792 546020 163844 547632
rect 164268 546020 164320 547632
rect 160754 545958 161802 546018
rect 166310 546018 166790 548298
rect 166798 546018 167358 548298
rect 166310 545958 167358 546018
rect 167762 548298 168810 548358
rect 167762 546018 168322 548298
rect 168330 546018 168810 548298
rect 173318 548298 174366 548358
rect 170800 546020 170852 547632
rect 171276 546020 171328 547632
rect 167762 545958 168810 546018
rect 173318 546018 173798 548298
rect 173806 546018 174366 548298
rect 173318 545958 174366 546018
rect 84528 537635 90592 537718
rect 144528 537665 150592 537748
rect 164528 537665 170592 537748
rect 82949 537475 82988 537565
rect 84611 535646 84612 537635
rect 85001 537246 85087 537635
rect 90055 537246 90141 537635
rect 85001 537245 90141 537246
rect 85001 536121 85087 537245
rect 90119 536121 90120 537245
rect 84979 536035 90141 536121
rect 85001 535646 85087 536035
rect 90055 535646 90141 536035
rect 90509 535646 90592 537635
rect 142949 537505 142988 537595
rect 144611 535676 144612 537665
rect 145001 537276 145087 537665
rect 150055 537276 150141 537665
rect 145001 537275 150141 537276
rect 145001 536151 145087 537275
rect 150119 536151 150120 537275
rect 144979 536065 150141 536151
rect 145001 535676 145087 536065
rect 150055 535676 150141 536065
rect 150509 535676 150592 537665
rect 162949 537505 162988 537595
rect 144611 535675 150592 535676
rect 164611 535676 164612 537665
rect 165001 537276 165087 537665
rect 170055 537276 170141 537665
rect 165001 537275 170141 537276
rect 165001 536151 165087 537275
rect 170119 536151 170120 537275
rect 164979 536065 170141 536151
rect 165001 535676 165087 536065
rect 170055 535676 170141 536065
rect 170509 535676 170592 537665
rect 164611 535675 170592 535676
rect 84611 535645 90592 535646
rect 82949 535031 82988 535177
rect 142949 535061 142988 535207
rect 162949 535061 162988 535207
rect 85165 534842 89955 534932
rect 145165 534872 149955 534962
rect 165165 534872 169955 534962
rect 85148 533156 85238 534750
rect 85302 534096 85392 534750
rect 85447 534688 89673 534778
rect 85447 534062 89673 534152
rect 89728 534096 89818 534750
rect 85306 533908 89814 533998
rect 85302 533162 85392 533816
rect 85447 533754 89673 533844
rect 85447 533128 89673 533218
rect 89728 533162 89818 533816
rect 89882 533156 89972 534750
rect 145148 533186 145238 534780
rect 145302 534126 145392 534780
rect 145447 534718 149673 534808
rect 145447 534092 149673 534182
rect 149728 534126 149818 534780
rect 145306 533938 149814 534028
rect 145302 533192 145392 533846
rect 145447 533784 149673 533874
rect 145447 533158 149673 533248
rect 149728 533192 149818 533846
rect 149882 533186 149972 534780
rect 165148 533186 165238 534780
rect 165302 534126 165392 534780
rect 165447 534718 169673 534808
rect 165447 534092 169673 534182
rect 169728 534126 169818 534780
rect 165306 533938 169814 534028
rect 165302 533192 165392 533846
rect 165447 533784 169673 533874
rect 165447 533158 169673 533248
rect 169728 533192 169818 533846
rect 169882 533186 169972 534780
rect 85165 532974 89955 533064
rect 145165 533004 149955 533094
rect 165165 533004 169955 533094
rect 84528 532261 90592 532344
rect 144528 532291 150592 532374
rect 164528 532291 170592 532374
rect 84611 529172 84612 532261
rect 85001 531872 85087 532261
rect 90055 531872 90141 532261
rect 85001 531871 90141 531872
rect 85001 531788 85087 531871
rect 85001 529647 85084 531788
rect 90119 529647 90120 531871
rect 84979 529644 85084 529647
rect 90036 529644 90141 529647
rect 84979 529561 90141 529644
rect 85001 529172 85087 529561
rect 90055 529172 90141 529561
rect 90509 529172 90592 532261
rect 144611 529202 144612 532291
rect 145001 531902 145087 532291
rect 150055 531902 150141 532291
rect 145001 531901 150141 531902
rect 145001 531818 145087 531901
rect 145001 529677 145084 531818
rect 150119 529677 150120 531901
rect 144979 529674 145084 529677
rect 150036 529674 150141 529677
rect 144979 529591 150141 529674
rect 145001 529202 145087 529591
rect 150055 529202 150141 529591
rect 150509 529202 150592 532291
rect 144611 529201 150592 529202
rect 164611 529202 164612 532291
rect 165001 531902 165087 532291
rect 170055 531902 170141 532291
rect 165001 531901 170141 531902
rect 165001 531818 165087 531901
rect 165001 529677 165084 531818
rect 170119 529677 170120 531901
rect 164979 529674 165084 529677
rect 170036 529674 170141 529677
rect 164979 529591 170141 529674
rect 165001 529202 165087 529591
rect 170055 529202 170141 529591
rect 170509 529202 170592 532291
rect 164611 529201 170592 529202
rect 84611 529171 90592 529172
rect 84138 528338 84162 528428
rect 144138 528368 144162 528458
rect 164138 528368 164162 528458
rect 84795 526026 84824 526082
rect 84851 525936 84880 526026
rect 85697 525936 85749 526082
rect 144795 526056 144824 526112
rect 144851 525966 144880 526056
rect 145697 525966 145749 526112
rect 164795 526056 164824 526112
rect 164851 525966 164880 526056
rect 165697 525966 165749 526112
rect 520064 521418 520116 577624
rect 17496 520064 73702 520116
rect 521247 520063 577705 520116
rect 577769 520063 577963 520116
rect 46792 513806 49192 514366
rect 46792 513798 46852 513806
rect 49132 513798 49224 513806
rect 46792 513318 49192 513798
rect 17839 513096 18410 513182
rect 27916 513096 28903 513182
rect 17922 513054 17923 513096
rect 18324 513054 18407 513096
rect 28002 513086 28903 513096
rect 17922 511028 18324 513054
rect 17922 502064 18324 504092
rect 17922 502024 17923 502064
rect 18324 502024 18407 502064
rect 27919 502032 28903 502092
rect 17922 502023 18407 502024
rect 28002 502024 28003 502032
rect 28820 502024 28903 502032
rect 28002 502023 28903 502024
rect 46792 501322 49192 501802
rect 46792 501314 46852 501322
rect 49132 501314 49224 501322
rect 46792 500754 49192 501314
rect 46792 493806 49192 494366
rect 46792 493798 46852 493806
rect 49132 493798 49224 493806
rect 46792 493318 49192 493798
rect 17839 493096 18410 493182
rect 27916 493096 28903 493182
rect 17922 493054 17923 493096
rect 18324 493054 18407 493096
rect 28002 493086 28903 493096
rect 17922 482064 18324 493054
rect 33184 492741 33186 492776
rect 33274 492741 33276 492797
rect 41272 492741 41274 492797
rect 41362 492741 41364 492776
rect 33184 492565 33186 492601
rect 33274 492475 33276 492601
rect 41272 492475 41274 492601
rect 41362 492565 41364 492601
rect 33184 491357 33186 491390
rect 33274 491357 33276 491480
rect 41272 491357 41274 491480
rect 41362 491357 41364 491390
rect 47518 491276 49130 491328
rect 33184 491179 33186 491217
rect 33274 491161 33276 491217
rect 41272 491161 41274 491217
rect 41362 491179 41364 491217
rect 33184 490973 33186 491004
rect 33274 490973 33276 491029
rect 41272 490973 41274 491029
rect 41362 490973 41364 491004
rect 33184 490793 33186 490833
rect 33274 490703 33276 490833
rect 41272 490703 41274 490833
rect 41362 490793 41364 490833
rect 47518 490800 49130 490852
rect 57402 490509 59558 490592
rect 62776 490509 66032 490592
rect 57485 490141 57486 490509
rect 59475 490141 59558 490509
rect 62859 490141 62860 490509
rect 65949 490141 66032 490509
rect 57402 490120 57961 490141
rect 58999 490120 59558 490141
rect 57402 490119 59558 490120
rect 57402 490055 57961 490119
rect 58999 490055 59558 490119
rect 62776 490120 63335 490141
rect 65473 490120 66032 490141
rect 62776 490119 66032 490120
rect 62776 490055 63335 490119
rect 65473 490055 66032 490119
rect 33184 489589 33186 489630
rect 33274 489589 33276 489720
rect 41272 489589 41274 489720
rect 41362 489589 41364 489630
rect 33184 489419 33186 489449
rect 33274 489393 33276 489449
rect 41272 489393 41274 489449
rect 41362 489419 41364 489449
rect 33184 489205 33186 489239
rect 33274 489205 33276 489261
rect 41272 489205 41274 489261
rect 41362 489205 41364 489239
rect 33184 489028 33186 489065
rect 33274 488938 33276 489065
rect 41272 488938 41274 489065
rect 41362 489028 41364 489065
rect 46792 488330 49192 488810
rect 46792 488322 46852 488330
rect 49132 488322 49224 488330
rect 33184 487821 33186 487858
rect 33274 487821 33276 487948
rect 41272 487821 41274 487948
rect 41362 487821 41364 487858
rect 46792 487762 49192 488322
rect 33184 487647 33186 487681
rect 33274 487625 33276 487681
rect 41272 487625 41274 487681
rect 41362 487647 41364 487681
rect 33184 487437 33186 487470
rect 33274 487437 33276 487493
rect 41272 487437 41274 487493
rect 41362 487437 41364 487470
rect 33184 487259 33186 487297
rect 33274 487169 33276 487297
rect 41272 487169 41274 487297
rect 41362 487259 41364 487297
rect 46792 486798 49192 487358
rect 46792 486790 46852 486798
rect 49132 486790 49224 486798
rect 46792 486310 49192 486790
rect 33184 486053 33186 486088
rect 33274 486053 33276 486178
rect 41272 486053 41274 486178
rect 41362 486053 41364 486088
rect 33184 485877 33186 485913
rect 33274 485857 33276 485913
rect 41272 485857 41274 485913
rect 41362 485877 41364 485913
rect 33184 485669 33186 485701
rect 33274 485669 33276 485725
rect 41272 485669 41274 485725
rect 41362 485669 41364 485701
rect 33184 485490 33186 485529
rect 33274 485400 33276 485529
rect 41272 485400 41274 485529
rect 41362 485490 41364 485529
rect 57485 485087 57486 490055
rect 57875 485087 57961 490055
rect 59085 485087 59086 490055
rect 59475 485087 59558 490055
rect 60188 485165 60278 489955
rect 60370 489882 61964 489972
rect 60370 489728 61024 489818
rect 60342 485447 60432 489673
rect 60968 485447 61058 489673
rect 60370 485302 61024 485392
rect 61122 485306 61212 489814
rect 61304 489728 61958 489818
rect 61276 485447 61366 489673
rect 61902 485447 61992 489673
rect 61304 485302 61958 485392
rect 60370 485148 61964 485238
rect 62056 485165 62146 489955
rect 62859 485087 62860 490055
rect 63249 490036 63335 490055
rect 63249 485087 63332 490036
rect 65559 485087 65560 490055
rect 65949 485087 66032 490055
rect 69038 485697 69184 485749
rect 57402 485001 59558 485087
rect 62776 485084 63332 485087
rect 65476 485084 66032 485087
rect 62776 485001 66032 485084
rect 57485 484612 57486 485001
rect 59475 484612 59558 485001
rect 57485 484611 59558 484612
rect 62859 484612 62860 485001
rect 65949 484612 66032 485001
rect 69094 484851 69184 484880
rect 62859 484611 66032 484612
rect 33184 484285 33186 484322
rect 33274 484285 33276 484412
rect 41272 484285 41274 484412
rect 41362 484285 41364 484322
rect 47518 484268 49130 484320
rect 33184 484111 33186 484145
rect 33274 484089 33276 484145
rect 41272 484089 41274 484145
rect 41362 484111 41364 484145
rect 66692 484138 66838 484162
rect 33184 483901 33186 483935
rect 33274 483901 33276 483957
rect 41272 483901 41274 483957
rect 41362 483901 41364 483935
rect 47518 483792 49130 483844
rect 33184 483724 33186 483761
rect 33274 483634 33276 483761
rect 41272 483634 41274 483761
rect 41362 483724 41364 483761
rect 57555 482949 57701 482988
rect 59943 482949 60089 482988
rect 33184 482517 33186 482549
rect 33274 482517 33276 482639
rect 41272 482517 41274 482639
rect 41362 482517 41364 482549
rect 33184 482338 33186 482377
rect 33274 482321 33276 482377
rect 41272 482321 41274 482377
rect 41362 482338 41364 482377
rect 17922 482024 17923 482064
rect 18324 482024 18407 482064
rect 27919 482032 28903 482118
rect 17922 482023 18407 482024
rect 28002 482024 28003 482032
rect 28820 482024 28903 482032
rect 28002 482023 28903 482024
rect 46792 481322 49192 481802
rect 46792 481314 46852 481322
rect 49132 481314 49224 481322
rect 46792 480754 49192 481314
rect 46792 453806 49192 454366
rect 46792 453798 46852 453806
rect 49132 453798 49224 453806
rect 46792 453318 49192 453798
rect 17839 453096 18410 453182
rect 27916 453096 28903 453182
rect 17922 453054 17923 453096
rect 18324 453054 18407 453096
rect 28002 453086 28903 453096
rect 17922 451028 18324 453054
rect 17922 442064 18324 444092
rect 17922 442024 17923 442064
rect 18324 442024 18407 442064
rect 27919 442032 28903 442092
rect 17922 442023 18407 442024
rect 28002 442024 28003 442032
rect 28820 442024 28903 442032
rect 28002 442023 28903 442024
rect 46792 441322 49192 441802
rect 46792 441314 46852 441322
rect 49132 441314 49224 441322
rect 46792 440754 49192 441314
rect 46792 433806 49192 434366
rect 46792 433798 46852 433806
rect 49132 433798 49224 433806
rect 46792 433318 49192 433798
rect 75954 433754 75955 433788
rect 17839 433096 18410 433182
rect 27916 433096 28903 433182
rect 17922 433054 17923 433096
rect 18324 433054 18407 433096
rect 28002 433086 28903 433096
rect 17922 422064 18324 433054
rect 33184 432741 33186 432776
rect 33274 432741 33276 432797
rect 41272 432741 41274 432797
rect 41362 432741 41364 432776
rect 33184 432565 33186 432601
rect 33274 432475 33276 432601
rect 41272 432475 41274 432601
rect 41362 432565 41364 432601
rect 33184 431357 33186 431390
rect 33274 431357 33276 431480
rect 41272 431357 41274 431480
rect 41362 431357 41364 431390
rect 47518 431276 49130 431328
rect 33184 431179 33186 431217
rect 33274 431161 33276 431217
rect 41272 431161 41274 431217
rect 41362 431179 41364 431217
rect 33184 430973 33186 431004
rect 33274 430973 33276 431029
rect 41272 430973 41274 431029
rect 41362 430973 41364 431004
rect 33184 430793 33186 430833
rect 33274 430703 33276 430833
rect 41272 430703 41274 430833
rect 41362 430793 41364 430833
rect 47518 430800 49130 430852
rect 57402 430509 59558 430592
rect 62776 430509 66032 430592
rect 57485 430141 57486 430509
rect 59475 430141 59558 430509
rect 62859 430141 62860 430509
rect 65949 430141 66032 430509
rect 57402 430120 57961 430141
rect 58999 430120 59558 430141
rect 57402 430119 59558 430120
rect 57402 430055 57961 430119
rect 58999 430055 59558 430119
rect 62776 430120 63335 430141
rect 65473 430120 66032 430141
rect 62776 430119 66032 430120
rect 62776 430055 63335 430119
rect 65473 430055 66032 430119
rect 33184 429589 33186 429630
rect 33274 429589 33276 429720
rect 41272 429589 41274 429720
rect 41362 429589 41364 429630
rect 33184 429419 33186 429449
rect 33274 429393 33276 429449
rect 41272 429393 41274 429449
rect 41362 429419 41364 429449
rect 33184 429205 33186 429239
rect 33274 429205 33276 429261
rect 41272 429205 41274 429261
rect 41362 429205 41364 429239
rect 33184 429028 33186 429065
rect 33274 428938 33276 429065
rect 41272 428938 41274 429065
rect 41362 429028 41364 429065
rect 46792 428330 49192 428810
rect 46792 428322 46852 428330
rect 49132 428322 49224 428330
rect 33184 427821 33186 427858
rect 33274 427821 33276 427948
rect 41272 427821 41274 427948
rect 41362 427821 41364 427858
rect 46792 427762 49192 428322
rect 33184 427647 33186 427681
rect 33274 427625 33276 427681
rect 41272 427625 41274 427681
rect 41362 427647 41364 427681
rect 33184 427437 33186 427470
rect 33274 427437 33276 427493
rect 41272 427437 41274 427493
rect 41362 427437 41364 427470
rect 33184 427259 33186 427297
rect 33274 427169 33276 427297
rect 41272 427169 41274 427297
rect 41362 427259 41364 427297
rect 46792 426798 49192 427358
rect 46792 426790 46852 426798
rect 49132 426790 49224 426798
rect 46792 426310 49192 426790
rect 33184 426053 33186 426088
rect 33274 426053 33276 426178
rect 41272 426053 41274 426178
rect 41362 426053 41364 426088
rect 33184 425877 33186 425913
rect 33274 425857 33276 425913
rect 41272 425857 41274 425913
rect 41362 425877 41364 425913
rect 33184 425669 33186 425701
rect 33274 425669 33276 425725
rect 41272 425669 41274 425725
rect 41362 425669 41364 425701
rect 33184 425490 33186 425529
rect 33274 425400 33276 425529
rect 41272 425400 41274 425529
rect 41362 425490 41364 425529
rect 57485 425087 57486 430055
rect 57875 425087 57961 430055
rect 59085 425087 59086 430055
rect 59475 425087 59558 430055
rect 60188 425165 60278 429955
rect 60370 429882 61964 429972
rect 60370 429728 61024 429818
rect 60342 425447 60432 429673
rect 60968 425447 61058 429673
rect 60370 425302 61024 425392
rect 61122 425306 61212 429814
rect 61304 429728 61958 429818
rect 61276 425447 61366 429673
rect 61902 425447 61992 429673
rect 61304 425302 61958 425392
rect 60370 425148 61964 425238
rect 62056 425165 62146 429955
rect 62859 425087 62860 430055
rect 63249 430036 63335 430055
rect 63249 425087 63332 430036
rect 65559 425087 65560 430055
rect 65949 425087 66032 430055
rect 69038 425697 69184 425749
rect 57402 425001 59558 425087
rect 62776 425084 63332 425087
rect 65476 425084 66032 425087
rect 62776 425001 66032 425084
rect 57485 424612 57486 425001
rect 59475 424612 59558 425001
rect 57485 424611 59558 424612
rect 62859 424612 62860 425001
rect 65949 424612 66032 425001
rect 69094 424851 69184 424880
rect 62859 424611 66032 424612
rect 33184 424285 33186 424322
rect 33274 424285 33276 424412
rect 41272 424285 41274 424412
rect 41362 424285 41364 424322
rect 47518 424268 49130 424320
rect 33184 424111 33186 424145
rect 33274 424089 33276 424145
rect 41272 424089 41274 424145
rect 41362 424111 41364 424145
rect 66692 424138 66838 424162
rect 33184 423901 33186 423935
rect 33274 423901 33276 423957
rect 41272 423901 41274 423957
rect 41362 423901 41364 423935
rect 47518 423792 49130 423844
rect 33184 423724 33186 423761
rect 33274 423634 33276 423761
rect 41272 423634 41274 423761
rect 41362 423724 41364 423761
rect 57555 422949 57701 422988
rect 59943 422949 60089 422988
rect 33184 422517 33186 422549
rect 33274 422517 33276 422639
rect 41272 422517 41274 422639
rect 41362 422517 41364 422549
rect 33184 422338 33186 422377
rect 33274 422321 33276 422377
rect 41272 422321 41274 422377
rect 41362 422338 41364 422377
rect 17922 422024 17923 422064
rect 18324 422024 18407 422064
rect 27919 422032 28903 422118
rect 17922 422023 18407 422024
rect 28002 422024 28003 422032
rect 28820 422024 28903 422032
rect 28002 422023 28903 422024
rect 46792 421322 49192 421802
rect 46792 421314 46852 421322
rect 49132 421314 49224 421322
rect 46792 420754 49192 421314
rect 46792 413806 49192 414366
rect 46792 413798 46852 413806
rect 49132 413798 49224 413806
rect 46792 413318 49192 413798
rect 17839 413096 18410 413182
rect 27916 413096 28903 413182
rect 17922 413054 17923 413096
rect 18324 413054 18407 413096
rect 28002 413086 28903 413096
rect 17922 402064 18324 413054
rect 33184 412741 33186 412776
rect 33274 412741 33276 412797
rect 41272 412741 41274 412797
rect 41362 412741 41364 412776
rect 33184 412565 33186 412601
rect 33274 412475 33276 412601
rect 41272 412475 41274 412601
rect 41362 412565 41364 412601
rect 33184 411357 33186 411390
rect 33274 411357 33276 411480
rect 41272 411357 41274 411480
rect 41362 411357 41364 411390
rect 47518 411276 49130 411328
rect 33184 411179 33186 411217
rect 33274 411161 33276 411217
rect 41272 411161 41274 411217
rect 41362 411179 41364 411217
rect 33184 410973 33186 411004
rect 33274 410973 33276 411029
rect 41272 410973 41274 411029
rect 41362 410973 41364 411004
rect 33184 410793 33186 410833
rect 33274 410703 33276 410833
rect 41272 410703 41274 410833
rect 41362 410793 41364 410833
rect 47518 410800 49130 410852
rect 57402 410509 59558 410592
rect 62776 410509 66032 410592
rect 57485 410141 57486 410509
rect 59475 410141 59558 410509
rect 62859 410141 62860 410509
rect 65949 410141 66032 410509
rect 57402 410120 57961 410141
rect 58999 410120 59558 410141
rect 57402 410119 59558 410120
rect 57402 410055 57961 410119
rect 58999 410055 59558 410119
rect 62776 410120 63335 410141
rect 65473 410120 66032 410141
rect 62776 410119 66032 410120
rect 62776 410055 63335 410119
rect 65473 410055 66032 410119
rect 33184 409589 33186 409630
rect 33274 409589 33276 409720
rect 41272 409589 41274 409720
rect 41362 409589 41364 409630
rect 33184 409419 33186 409449
rect 33274 409393 33276 409449
rect 41272 409393 41274 409449
rect 41362 409419 41364 409449
rect 33184 409205 33186 409239
rect 33274 409205 33276 409261
rect 41272 409205 41274 409261
rect 41362 409205 41364 409239
rect 33184 409028 33186 409065
rect 33274 408938 33276 409065
rect 41272 408938 41274 409065
rect 41362 409028 41364 409065
rect 46792 408330 49192 408810
rect 46792 408322 46852 408330
rect 49132 408322 49224 408330
rect 33184 407821 33186 407858
rect 33274 407821 33276 407948
rect 41272 407821 41274 407948
rect 41362 407821 41364 407858
rect 46792 407762 49192 408322
rect 33184 407647 33186 407681
rect 33274 407625 33276 407681
rect 41272 407625 41274 407681
rect 41362 407647 41364 407681
rect 33184 407437 33186 407470
rect 33274 407437 33276 407493
rect 41272 407437 41274 407493
rect 41362 407437 41364 407470
rect 33184 407259 33186 407297
rect 33274 407169 33276 407297
rect 41272 407169 41274 407297
rect 41362 407259 41364 407297
rect 46792 406798 49192 407358
rect 46792 406790 46852 406798
rect 49132 406790 49224 406798
rect 46792 406310 49192 406790
rect 33184 406053 33186 406088
rect 33274 406053 33276 406178
rect 41272 406053 41274 406178
rect 41362 406053 41364 406088
rect 33184 405877 33186 405913
rect 33274 405857 33276 405913
rect 41272 405857 41274 405913
rect 41362 405877 41364 405913
rect 33184 405669 33186 405701
rect 33274 405669 33276 405725
rect 41272 405669 41274 405725
rect 41362 405669 41364 405701
rect 33184 405490 33186 405529
rect 33274 405400 33276 405529
rect 41272 405400 41274 405529
rect 41362 405490 41364 405529
rect 57485 405087 57486 410055
rect 57875 405087 57961 410055
rect 59085 405087 59086 410055
rect 59475 405087 59558 410055
rect 60188 405165 60278 409955
rect 60370 409882 61964 409972
rect 60370 409728 61024 409818
rect 60342 405447 60432 409673
rect 60968 405447 61058 409673
rect 60370 405302 61024 405392
rect 61122 405306 61212 409814
rect 61304 409728 61958 409818
rect 61276 405447 61366 409673
rect 61902 405447 61992 409673
rect 61304 405302 61958 405392
rect 60370 405148 61964 405238
rect 62056 405165 62146 409955
rect 62859 405087 62860 410055
rect 63249 410036 63335 410055
rect 63249 405087 63332 410036
rect 65559 405087 65560 410055
rect 65949 405087 66032 410055
rect 69038 405697 69184 405749
rect 57402 405001 59558 405087
rect 62776 405084 63332 405087
rect 65476 405084 66032 405087
rect 62776 405001 66032 405084
rect 57485 404612 57486 405001
rect 59475 404612 59558 405001
rect 57485 404611 59558 404612
rect 62859 404612 62860 405001
rect 65949 404612 66032 405001
rect 69094 404851 69184 404880
rect 62859 404611 66032 404612
rect 33184 404285 33186 404322
rect 33274 404285 33276 404412
rect 41272 404285 41274 404412
rect 41362 404285 41364 404322
rect 47518 404268 49130 404320
rect 33184 404111 33186 404145
rect 33274 404089 33276 404145
rect 41272 404089 41274 404145
rect 41362 404111 41364 404145
rect 66692 404138 66838 404162
rect 33184 403901 33186 403935
rect 33274 403901 33276 403957
rect 41272 403901 41274 403957
rect 41362 403901 41364 403935
rect 47518 403792 49130 403844
rect 33184 403724 33186 403761
rect 33274 403634 33276 403761
rect 41272 403634 41274 403761
rect 41362 403724 41364 403761
rect 57555 402949 57701 402988
rect 59943 402949 60089 402988
rect 33184 402517 33186 402549
rect 33274 402517 33276 402639
rect 41272 402517 41274 402639
rect 41362 402517 41364 402549
rect 33184 402338 33186 402377
rect 33274 402321 33276 402377
rect 41272 402321 41274 402377
rect 41362 402338 41364 402377
rect 17922 402024 17923 402064
rect 18324 402024 18407 402064
rect 27919 402032 28903 402118
rect 17922 402023 18407 402024
rect 28002 402024 28003 402032
rect 28820 402024 28903 402032
rect 28002 402023 28903 402024
rect 46792 401322 49192 401802
rect 46792 401314 46852 401322
rect 49132 401314 49224 401322
rect 46792 400754 49192 401314
rect 46792 393806 49192 394366
rect 46792 393798 46852 393806
rect 49132 393798 49224 393806
rect 46792 393318 49192 393798
rect 17839 393096 18410 393182
rect 27916 393096 28903 393182
rect 17922 393054 17923 393096
rect 18324 393054 18407 393096
rect 28002 393086 28903 393096
rect 17922 391028 18324 393054
rect 17922 382064 18324 384000
rect 17922 382024 17923 382064
rect 18324 382024 18407 382064
rect 27919 382032 28903 382092
rect 17922 382023 18407 382024
rect 28002 382024 28003 382032
rect 28820 382024 28903 382032
rect 28002 382023 28903 382024
rect 46792 381322 49192 381802
rect 46792 381314 46852 381322
rect 49132 381314 49224 381322
rect 46792 380754 49192 381314
rect 46792 353806 49192 354366
rect 46792 353798 46852 353806
rect 49132 353798 49224 353806
rect 46792 353318 49192 353798
rect 17839 353096 18410 353182
rect 27916 353096 28903 353182
rect 17922 353054 17923 353096
rect 18324 353054 18407 353096
rect 28002 353086 28903 353096
rect 17922 351028 18324 353054
rect 17922 342064 18324 344092
rect 17922 342024 17923 342064
rect 18324 342024 18407 342064
rect 27919 342032 28903 342092
rect 17922 342023 18407 342024
rect 28002 342024 28003 342032
rect 28820 342024 28903 342032
rect 28002 342023 28903 342024
rect 46792 341322 49192 341802
rect 46792 341314 46852 341322
rect 49132 341314 49224 341322
rect 46792 340754 49192 341314
rect 46792 333806 49192 334366
rect 46792 333798 46852 333806
rect 49132 333798 49224 333806
rect 46792 333318 49192 333798
rect 17839 333096 18410 333182
rect 27916 333096 28903 333182
rect 17922 333054 17923 333096
rect 18324 333054 18407 333096
rect 28002 333086 28903 333096
rect 17922 322064 18324 333054
rect 33184 332741 33186 332776
rect 33274 332741 33276 332797
rect 41272 332741 41274 332797
rect 41362 332741 41364 332776
rect 33184 332565 33186 332601
rect 33274 332475 33276 332601
rect 41272 332475 41274 332601
rect 41362 332565 41364 332601
rect 33184 331357 33186 331390
rect 33274 331357 33276 331480
rect 41272 331357 41274 331480
rect 41362 331357 41364 331390
rect 47518 331276 49130 331328
rect 33184 331179 33186 331217
rect 33274 331161 33276 331217
rect 41272 331161 41274 331217
rect 41362 331179 41364 331217
rect 33184 330973 33186 331004
rect 33274 330973 33276 331029
rect 41272 330973 41274 331029
rect 41362 330973 41364 331004
rect 33184 330793 33186 330833
rect 33274 330703 33276 330833
rect 41272 330703 41274 330833
rect 41362 330793 41364 330833
rect 47518 330800 49130 330852
rect 57402 330509 59558 330592
rect 62776 330509 66032 330592
rect 57485 330141 57486 330509
rect 59475 330141 59558 330509
rect 62859 330141 62860 330509
rect 65949 330141 66032 330509
rect 57402 330120 57961 330141
rect 58999 330120 59558 330141
rect 57402 330119 59558 330120
rect 57402 330055 57961 330119
rect 58999 330055 59558 330119
rect 62776 330120 63335 330141
rect 65473 330120 66032 330141
rect 62776 330119 66032 330120
rect 62776 330055 63335 330119
rect 65473 330055 66032 330119
rect 33184 329589 33186 329630
rect 33274 329589 33276 329720
rect 41272 329589 41274 329720
rect 41362 329589 41364 329630
rect 33184 329419 33186 329449
rect 33274 329393 33276 329449
rect 41272 329393 41274 329449
rect 41362 329419 41364 329449
rect 33184 329205 33186 329239
rect 33274 329205 33276 329261
rect 41272 329205 41274 329261
rect 41362 329205 41364 329239
rect 33184 329028 33186 329065
rect 33274 328938 33276 329065
rect 41272 328938 41274 329065
rect 41362 329028 41364 329065
rect 46792 328330 49192 328810
rect 46792 328322 46852 328330
rect 49132 328322 49224 328330
rect 33184 327821 33186 327858
rect 33274 327821 33276 327948
rect 41272 327821 41274 327948
rect 41362 327821 41364 327858
rect 46792 327762 49192 328322
rect 33184 327647 33186 327681
rect 33274 327625 33276 327681
rect 41272 327625 41274 327681
rect 41362 327647 41364 327681
rect 33184 327437 33186 327470
rect 33274 327437 33276 327493
rect 41272 327437 41274 327493
rect 41362 327437 41364 327470
rect 33184 327259 33186 327297
rect 33274 327169 33276 327297
rect 41272 327169 41274 327297
rect 41362 327259 41364 327297
rect 46792 326798 49192 327358
rect 46792 326790 46852 326798
rect 49132 326790 49224 326798
rect 46792 326310 49192 326790
rect 33184 326053 33186 326088
rect 33274 326053 33276 326178
rect 41272 326053 41274 326178
rect 41362 326053 41364 326088
rect 33184 325877 33186 325913
rect 33274 325857 33276 325913
rect 41272 325857 41274 325913
rect 41362 325877 41364 325913
rect 33184 325669 33186 325701
rect 33274 325669 33276 325725
rect 41272 325669 41274 325725
rect 41362 325669 41364 325701
rect 33184 325490 33186 325529
rect 33274 325400 33276 325529
rect 41272 325400 41274 325529
rect 41362 325490 41364 325529
rect 57485 325087 57486 330055
rect 57875 325087 57961 330055
rect 59085 325087 59086 330055
rect 59475 325087 59558 330055
rect 60188 325165 60278 329955
rect 60370 329882 61964 329972
rect 60370 329728 61024 329818
rect 60342 325447 60432 329673
rect 60968 325447 61058 329673
rect 60370 325302 61024 325392
rect 61122 325306 61212 329814
rect 61304 329728 61958 329818
rect 61276 325447 61366 329673
rect 61902 325447 61992 329673
rect 61304 325302 61958 325392
rect 60370 325148 61964 325238
rect 62056 325165 62146 329955
rect 62859 325087 62860 330055
rect 63249 330036 63335 330055
rect 63249 325087 63332 330036
rect 65559 325087 65560 330055
rect 65949 325087 66032 330055
rect 69038 325697 69184 325749
rect 57402 325001 59558 325087
rect 62776 325084 63332 325087
rect 65476 325084 66032 325087
rect 62776 325001 66032 325084
rect 57485 324612 57486 325001
rect 59475 324612 59558 325001
rect 57485 324611 59558 324612
rect 62859 324612 62860 325001
rect 65949 324612 66032 325001
rect 69094 324851 69184 324880
rect 62859 324611 66032 324612
rect 33184 324285 33186 324322
rect 33274 324285 33276 324412
rect 41272 324285 41274 324412
rect 41362 324285 41364 324322
rect 47518 324268 49130 324320
rect 33184 324111 33186 324145
rect 33274 324089 33276 324145
rect 41272 324089 41274 324145
rect 41362 324111 41364 324145
rect 66692 324138 66838 324162
rect 33184 323901 33186 323935
rect 33274 323901 33276 323957
rect 41272 323901 41274 323957
rect 41362 323901 41364 323935
rect 47518 323792 49130 323844
rect 33184 323724 33186 323761
rect 33274 323634 33276 323761
rect 41272 323634 41274 323761
rect 41362 323724 41364 323761
rect 57555 322949 57701 322988
rect 59943 322949 60089 322988
rect 33184 322517 33186 322549
rect 33274 322517 33276 322639
rect 41272 322517 41274 322639
rect 41362 322517 41364 322549
rect 33184 322338 33186 322377
rect 33274 322321 33276 322377
rect 41272 322321 41274 322377
rect 41362 322338 41364 322377
rect 17922 322024 17923 322064
rect 18324 322024 18407 322064
rect 27919 322032 28903 322118
rect 17922 322023 18407 322024
rect 28002 322024 28003 322032
rect 28820 322024 28903 322032
rect 28002 322023 28903 322024
rect 46792 321322 49192 321802
rect 46792 321314 46852 321322
rect 49132 321314 49224 321322
rect 46792 320754 49192 321314
rect 46792 313806 49192 314366
rect 46792 313798 46852 313806
rect 49132 313798 49224 313806
rect 46792 313318 49192 313798
rect 17839 313096 18410 313182
rect 27916 313096 28903 313182
rect 17922 313054 17923 313096
rect 18324 313054 18407 313096
rect 28002 313086 28903 313096
rect 17922 302064 18324 313054
rect 33184 312741 33186 312776
rect 33274 312741 33276 312797
rect 41272 312741 41274 312797
rect 41362 312741 41364 312776
rect 33184 312565 33186 312601
rect 33274 312475 33276 312601
rect 41272 312475 41274 312601
rect 41362 312565 41364 312601
rect 33184 311357 33186 311390
rect 33274 311357 33276 311480
rect 41272 311357 41274 311480
rect 41362 311357 41364 311390
rect 47518 311276 49130 311328
rect 33184 311179 33186 311217
rect 33274 311161 33276 311217
rect 41272 311161 41274 311217
rect 41362 311179 41364 311217
rect 33184 310973 33186 311004
rect 33274 310973 33276 311029
rect 41272 310973 41274 311029
rect 41362 310973 41364 311004
rect 33184 310793 33186 310833
rect 33274 310703 33276 310833
rect 41272 310703 41274 310833
rect 41362 310793 41364 310833
rect 47518 310800 49130 310852
rect 57402 310509 59558 310592
rect 62776 310509 66032 310592
rect 57485 310141 57486 310509
rect 59475 310141 59558 310509
rect 62859 310141 62860 310509
rect 65949 310141 66032 310509
rect 57402 310120 57961 310141
rect 58999 310120 59558 310141
rect 57402 310119 59558 310120
rect 57402 310055 57961 310119
rect 58999 310055 59558 310119
rect 62776 310120 63335 310141
rect 65473 310120 66032 310141
rect 62776 310119 66032 310120
rect 62776 310055 63335 310119
rect 65473 310055 66032 310119
rect 33184 309589 33186 309630
rect 33274 309589 33276 309720
rect 41272 309589 41274 309720
rect 41362 309589 41364 309630
rect 33184 309419 33186 309449
rect 33274 309393 33276 309449
rect 41272 309393 41274 309449
rect 41362 309419 41364 309449
rect 33184 309205 33186 309239
rect 33274 309205 33276 309261
rect 41272 309205 41274 309261
rect 41362 309205 41364 309239
rect 33184 309028 33186 309065
rect 33274 308938 33276 309065
rect 41272 308938 41274 309065
rect 41362 309028 41364 309065
rect 46792 308330 49192 308810
rect 46792 308322 46852 308330
rect 49132 308322 49224 308330
rect 33184 307821 33186 307858
rect 33274 307821 33276 307948
rect 41272 307821 41274 307948
rect 41362 307821 41364 307858
rect 46792 307762 49192 308322
rect 33184 307647 33186 307681
rect 33274 307625 33276 307681
rect 41272 307625 41274 307681
rect 41362 307647 41364 307681
rect 33184 307437 33186 307470
rect 33274 307437 33276 307493
rect 41272 307437 41274 307493
rect 41362 307437 41364 307470
rect 33184 307259 33186 307297
rect 33274 307169 33276 307297
rect 41272 307169 41274 307297
rect 41362 307259 41364 307297
rect 46792 306798 49192 307358
rect 46792 306790 46852 306798
rect 49132 306790 49224 306798
rect 46792 306310 49192 306790
rect 33184 306053 33186 306088
rect 33274 306053 33276 306178
rect 41272 306053 41274 306178
rect 41362 306053 41364 306088
rect 33184 305877 33186 305913
rect 33274 305857 33276 305913
rect 41272 305857 41274 305913
rect 41362 305877 41364 305913
rect 33184 305669 33186 305701
rect 33274 305669 33276 305725
rect 41272 305669 41274 305725
rect 41362 305669 41364 305701
rect 33184 305490 33186 305529
rect 33274 305400 33276 305529
rect 41272 305400 41274 305529
rect 41362 305490 41364 305529
rect 57485 305087 57486 310055
rect 57875 305087 57961 310055
rect 59085 305087 59086 310055
rect 59475 305087 59558 310055
rect 60188 305165 60278 309955
rect 60370 309882 61964 309972
rect 60370 309728 61024 309818
rect 60342 305447 60432 309673
rect 60968 305447 61058 309673
rect 60370 305302 61024 305392
rect 61122 305306 61212 309814
rect 61304 309728 61958 309818
rect 61276 305447 61366 309673
rect 61902 305447 61992 309673
rect 61304 305302 61958 305392
rect 60370 305148 61964 305238
rect 62056 305165 62146 309955
rect 62859 305087 62860 310055
rect 63249 310036 63335 310055
rect 63249 305087 63332 310036
rect 65559 305087 65560 310055
rect 65949 305087 66032 310055
rect 69038 305697 69184 305749
rect 57402 305001 59558 305087
rect 62776 305084 63332 305087
rect 65476 305084 66032 305087
rect 62776 305001 66032 305084
rect 57485 304612 57486 305001
rect 59475 304612 59558 305001
rect 57485 304611 59558 304612
rect 62859 304612 62860 305001
rect 65949 304612 66032 305001
rect 69094 304851 69184 304880
rect 62859 304611 66032 304612
rect 33184 304285 33186 304322
rect 33274 304285 33276 304412
rect 41272 304285 41274 304412
rect 41362 304285 41364 304322
rect 47518 304268 49130 304320
rect 33184 304111 33186 304145
rect 33274 304089 33276 304145
rect 41272 304089 41274 304145
rect 41362 304111 41364 304145
rect 66692 304138 66838 304162
rect 33184 303901 33186 303935
rect 33274 303901 33276 303957
rect 41272 303901 41274 303957
rect 41362 303901 41364 303935
rect 47518 303792 49130 303844
rect 33184 303724 33186 303761
rect 33274 303634 33276 303761
rect 41272 303634 41274 303761
rect 41362 303724 41364 303761
rect 57555 302949 57701 302988
rect 59943 302949 60089 302988
rect 33184 302517 33186 302549
rect 33274 302517 33276 302639
rect 41272 302517 41274 302639
rect 41362 302517 41364 302549
rect 33184 302338 33186 302377
rect 33274 302321 33276 302377
rect 41272 302321 41274 302377
rect 41362 302338 41364 302377
rect 17922 302024 17923 302064
rect 18324 302024 18407 302064
rect 27919 302032 28903 302118
rect 17922 302023 18407 302024
rect 28002 302024 28003 302032
rect 28820 302024 28903 302032
rect 28002 302023 28903 302024
rect 46792 301322 49192 301802
rect 46792 301314 46852 301322
rect 49132 301314 49224 301322
rect 46792 300754 49192 301314
rect 46792 293806 49192 294366
rect 46792 293798 46852 293806
rect 49132 293798 49224 293806
rect 46792 293318 49192 293798
rect 17839 293096 18410 293182
rect 27916 293096 28903 293182
rect 17922 293054 17923 293096
rect 18324 293054 18407 293096
rect 28002 293086 28903 293096
rect 17922 291028 18324 293054
rect 17922 282064 18324 284092
rect 17922 282024 17923 282064
rect 18324 282024 18407 282064
rect 27919 282032 28903 282092
rect 17922 282023 18407 282024
rect 28002 282024 28003 282032
rect 28820 282024 28903 282032
rect 28002 282023 28903 282024
rect 46792 281322 49192 281802
rect 46792 281314 46852 281322
rect 49132 281314 49224 281322
rect 46792 280754 49192 281314
rect 545958 273806 548358 274366
rect 545958 273798 546018 273806
rect 548298 273798 548390 273806
rect 545958 273318 548358 273798
rect 566247 273097 567234 273183
rect 576740 273097 577311 273183
rect 566330 273088 567231 273097
rect 576826 273056 576827 273097
rect 577228 273056 577311 273097
rect 553786 272743 553788 272782
rect 553876 272743 553878 272799
rect 561874 272743 561876 272799
rect 561964 272743 561966 272782
rect 553786 272571 553788 272603
rect 553876 272481 553878 272603
rect 561874 272481 561876 272603
rect 561964 272571 561966 272603
rect 535061 272188 535151 272227
rect 537505 272188 537595 272227
rect 553786 271359 553788 271396
rect 553876 271359 553878 271486
rect 561874 271359 561876 271486
rect 561964 271359 561966 271396
rect 546020 271276 547632 271328
rect 553786 271185 553788 271219
rect 553876 271163 553878 271219
rect 561874 271163 561876 271219
rect 561964 271185 561966 271219
rect 528368 271014 528458 271038
rect 553786 270975 553788 271009
rect 553876 270975 553878 271031
rect 561874 270975 561876 271031
rect 561964 270975 561966 271009
rect 546020 270800 547632 270852
rect 553786 270798 553788 270835
rect 553876 270708 553878 270835
rect 561874 270708 561876 270835
rect 561964 270798 561966 270835
rect 530544 270592 531740 270595
rect 529118 270509 532374 270592
rect 535592 270509 537748 270592
rect 525966 270296 526112 270325
rect 529201 270141 529202 270509
rect 532291 270141 532374 270509
rect 535675 270141 535676 270509
rect 537665 270141 537748 270509
rect 529118 270120 529677 270141
rect 531815 270120 532374 270141
rect 529118 270119 532374 270120
rect 529118 270055 529677 270119
rect 531815 270055 532374 270119
rect 535592 270120 536151 270141
rect 537189 270120 537748 270141
rect 535592 270119 537748 270120
rect 535592 270055 536151 270119
rect 537189 270055 537748 270119
rect 525966 269427 526056 269479
rect 529201 265087 529202 270055
rect 529591 270036 529677 270055
rect 529591 265087 529674 270036
rect 531901 265087 531902 270055
rect 532291 265087 532374 270055
rect 533004 265165 533094 269955
rect 533186 269882 534780 269972
rect 533192 269728 533846 269818
rect 533158 265447 533248 269673
rect 533784 265447 533874 269673
rect 533192 265302 533846 265392
rect 533938 265306 534028 269814
rect 534126 269728 534780 269818
rect 534092 265447 534182 269673
rect 534718 265447 534808 269673
rect 534126 265302 534780 265392
rect 533186 265148 534780 265238
rect 534872 265165 534962 269955
rect 535675 265087 535676 270055
rect 536065 265087 536151 270055
rect 537275 265087 537276 270055
rect 537665 265087 537748 270055
rect 553786 269591 553788 269630
rect 553876 269591 553878 269720
rect 561874 269591 561876 269720
rect 561964 269591 561966 269630
rect 553786 269419 553788 269451
rect 553876 269395 553878 269451
rect 561874 269395 561876 269451
rect 561964 269419 561966 269451
rect 553786 269207 553788 269243
rect 553876 269207 553878 269263
rect 561874 269207 561876 269263
rect 561964 269207 561966 269243
rect 553786 269032 553788 269067
rect 553876 268942 553878 269067
rect 561874 268942 561876 269067
rect 561964 269032 561966 269067
rect 545958 268330 548358 268810
rect 545958 268322 546018 268330
rect 548298 268322 548390 268330
rect 545958 267762 548358 268322
rect 553786 267823 553788 267861
rect 553876 267823 553878 267951
rect 561874 267823 561876 267951
rect 561964 267823 561966 267861
rect 553786 267650 553788 267683
rect 553876 267627 553878 267683
rect 561874 267627 561876 267683
rect 561964 267650 561966 267683
rect 553786 267439 553788 267473
rect 553876 267439 553878 267495
rect 561874 267439 561876 267495
rect 561964 267439 561966 267473
rect 545958 266798 548358 267358
rect 553786 267262 553788 267299
rect 553876 267172 553878 267299
rect 561874 267172 561876 267299
rect 561964 267262 561966 267299
rect 545958 266790 546018 266798
rect 548298 266790 548390 266798
rect 545958 266310 548358 266790
rect 553786 266055 553788 266092
rect 553876 266055 553878 266182
rect 561874 266055 561876 266182
rect 561964 266055 561966 266092
rect 553786 265881 553788 265915
rect 553876 265859 553878 265915
rect 561874 265859 561876 265915
rect 561964 265881 561966 265915
rect 553786 265671 553788 265701
rect 553876 265671 553878 265727
rect 561874 265671 561876 265727
rect 561964 265671 561966 265701
rect 553786 265490 553788 265531
rect 553876 265400 553878 265531
rect 561874 265400 561876 265531
rect 561964 265490 561966 265531
rect 529118 265084 529674 265087
rect 531818 265084 532374 265087
rect 529118 265001 532374 265084
rect 535592 265001 537748 265087
rect 529201 264612 529202 265001
rect 532291 264612 532374 265001
rect 529201 264611 532374 264612
rect 535675 264612 535676 265001
rect 537665 264612 537748 265001
rect 535675 264611 537748 264612
rect 546020 264268 547632 264320
rect 553786 264287 553788 264327
rect 553876 264287 553878 264417
rect 561874 264287 561876 264417
rect 561964 264287 561966 264327
rect 553786 264116 553788 264147
rect 553876 264091 553878 264147
rect 561874 264091 561876 264147
rect 561964 264116 561966 264147
rect 553786 263903 553788 263941
rect 553876 263903 553878 263959
rect 561874 263903 561876 263959
rect 561964 263903 561966 263941
rect 546020 263792 547632 263844
rect 553786 263730 553788 263763
rect 553876 263640 553878 263763
rect 561874 263640 561876 263763
rect 561964 263730 561966 263763
rect 553786 262519 553788 262555
rect 553876 262519 553878 262645
rect 561874 262519 561876 262645
rect 561964 262519 561966 262555
rect 553786 262344 553788 262379
rect 553876 262323 553878 262379
rect 561874 262323 561876 262379
rect 561964 262344 561966 262379
rect 566247 262034 567231 262120
rect 566330 262025 566331 262034
rect 567148 262025 567231 262034
rect 566330 262024 567231 262025
rect 576826 262066 577228 273056
rect 576826 262025 576827 262066
rect 577228 262025 577311 262066
rect 576826 262024 577311 262025
rect 545958 261322 548358 261802
rect 545958 261314 546018 261322
rect 548298 261314 548390 261322
rect 545958 260754 548358 261314
rect 46792 253806 49192 254366
rect 545958 253806 548358 254366
rect 46792 253798 46852 253806
rect 49132 253798 49224 253806
rect 545958 253798 546018 253806
rect 548298 253798 548390 253806
rect 46792 253318 49192 253798
rect 545958 253318 548358 253798
rect 17839 253096 18410 253182
rect 27916 253096 28903 253182
rect 566247 253097 567234 253183
rect 576740 253097 577311 253183
rect 17922 253054 17923 253096
rect 18324 253054 18407 253096
rect 28002 253086 28903 253096
rect 566330 253088 567231 253097
rect 576826 253056 576827 253097
rect 577228 253056 577311 253097
rect 17922 242064 18324 253054
rect 33184 252741 33186 252776
rect 33274 252741 33276 252797
rect 41272 252741 41274 252797
rect 41362 252741 41364 252776
rect 553786 252743 553788 252782
rect 553876 252743 553878 252799
rect 561874 252743 561876 252799
rect 561964 252743 561966 252782
rect 33184 252565 33186 252601
rect 33274 252475 33276 252601
rect 41272 252475 41274 252601
rect 41362 252565 41364 252601
rect 553786 252571 553788 252603
rect 553876 252481 553878 252603
rect 561874 252481 561876 252603
rect 561964 252571 561966 252603
rect 535061 252188 535151 252227
rect 537505 252188 537595 252227
rect 33184 251357 33186 251390
rect 33274 251357 33276 251480
rect 41272 251357 41274 251480
rect 41362 251357 41364 251390
rect 553786 251359 553788 251396
rect 553876 251359 553878 251486
rect 561874 251359 561876 251486
rect 561964 251359 561966 251396
rect 47518 251276 49130 251328
rect 546020 251276 547632 251328
rect 33184 251179 33186 251217
rect 33274 251161 33276 251217
rect 41272 251161 41274 251217
rect 41362 251179 41364 251217
rect 553786 251185 553788 251219
rect 553876 251163 553878 251219
rect 561874 251163 561876 251219
rect 561964 251185 561966 251219
rect 33184 250973 33186 251004
rect 33274 250973 33276 251029
rect 41272 250973 41274 251029
rect 528368 251014 528458 251038
rect 41362 250973 41364 251004
rect 553786 250975 553788 251009
rect 553876 250975 553878 251031
rect 561874 250975 561876 251031
rect 561964 250975 561966 251009
rect 33184 250793 33186 250833
rect 33274 250703 33276 250833
rect 41272 250703 41274 250833
rect 41362 250793 41364 250833
rect 47518 250800 49130 250852
rect 546020 250800 547632 250852
rect 553786 250798 553788 250835
rect 553876 250708 553878 250835
rect 561874 250708 561876 250835
rect 561964 250798 561966 250835
rect 530544 250592 531740 250595
rect 57402 250509 59558 250592
rect 62776 250509 66032 250592
rect 529118 250509 532374 250592
rect 535592 250509 537748 250592
rect 57485 250141 57486 250509
rect 59475 250141 59558 250509
rect 62859 250141 62860 250509
rect 65949 250141 66032 250509
rect 525966 250296 526112 250325
rect 529201 250141 529202 250509
rect 532291 250141 532374 250509
rect 535675 250141 535676 250509
rect 537665 250141 537748 250509
rect 57402 250120 57961 250141
rect 58999 250120 59558 250141
rect 57402 250119 59558 250120
rect 57402 250055 57961 250119
rect 58999 250055 59558 250119
rect 62776 250120 63335 250141
rect 65473 250120 66032 250141
rect 62776 250119 66032 250120
rect 62776 250055 63335 250119
rect 65473 250055 66032 250119
rect 529118 250120 529677 250141
rect 531815 250120 532374 250141
rect 529118 250119 532374 250120
rect 529118 250055 529677 250119
rect 531815 250055 532374 250119
rect 535592 250120 536151 250141
rect 537189 250120 537748 250141
rect 535592 250119 537748 250120
rect 535592 250055 536151 250119
rect 537189 250055 537748 250119
rect 33184 249589 33186 249630
rect 33274 249589 33276 249720
rect 41272 249589 41274 249720
rect 41362 249589 41364 249630
rect 33184 249419 33186 249449
rect 33274 249393 33276 249449
rect 41272 249393 41274 249449
rect 41362 249419 41364 249449
rect 33184 249205 33186 249239
rect 33274 249205 33276 249261
rect 41272 249205 41274 249261
rect 41362 249205 41364 249239
rect 33184 249028 33186 249065
rect 33274 248938 33276 249065
rect 41272 248938 41274 249065
rect 41362 249028 41364 249065
rect 46792 248330 49192 248810
rect 46792 248322 46852 248330
rect 49132 248322 49224 248330
rect 33184 247821 33186 247858
rect 33274 247821 33276 247948
rect 41272 247821 41274 247948
rect 41362 247821 41364 247858
rect 46792 247762 49192 248322
rect 33184 247647 33186 247681
rect 33274 247625 33276 247681
rect 41272 247625 41274 247681
rect 41362 247647 41364 247681
rect 33184 247437 33186 247470
rect 33274 247437 33276 247493
rect 41272 247437 41274 247493
rect 41362 247437 41364 247470
rect 33184 247259 33186 247297
rect 33274 247169 33276 247297
rect 41272 247169 41274 247297
rect 41362 247259 41364 247297
rect 46792 246798 49192 247358
rect 46792 246790 46852 246798
rect 49132 246790 49224 246798
rect 46792 246310 49192 246790
rect 33184 246053 33186 246088
rect 33274 246053 33276 246178
rect 41272 246053 41274 246178
rect 41362 246053 41364 246088
rect 33184 245877 33186 245913
rect 33274 245857 33276 245913
rect 41272 245857 41274 245913
rect 41362 245877 41364 245913
rect 33184 245669 33186 245701
rect 33274 245669 33276 245725
rect 41272 245669 41274 245725
rect 41362 245669 41364 245701
rect 33184 245490 33186 245529
rect 33274 245400 33276 245529
rect 41272 245400 41274 245529
rect 41362 245490 41364 245529
rect 57485 245087 57486 250055
rect 57875 245087 57961 250055
rect 59085 245087 59086 250055
rect 59475 245087 59558 250055
rect 60188 245165 60278 249955
rect 60370 249882 61964 249972
rect 60370 249728 61024 249818
rect 60342 245447 60432 249673
rect 60968 245447 61058 249673
rect 60370 245302 61024 245392
rect 61122 245306 61212 249814
rect 61304 249728 61958 249818
rect 61276 245447 61366 249673
rect 61902 245447 61992 249673
rect 61304 245302 61958 245392
rect 60370 245148 61964 245238
rect 62056 245165 62146 249955
rect 62859 245087 62860 250055
rect 63249 250036 63335 250055
rect 63249 245087 63332 250036
rect 65559 245087 65560 250055
rect 65949 245087 66032 250055
rect 525966 249427 526056 249479
rect 69038 245697 69184 245749
rect 529201 245087 529202 250055
rect 529591 250036 529677 250055
rect 529591 245087 529674 250036
rect 531901 245087 531902 250055
rect 532291 245087 532374 250055
rect 533004 245165 533094 249955
rect 533186 249882 534780 249972
rect 533192 249728 533846 249818
rect 533158 245447 533248 249673
rect 533784 245447 533874 249673
rect 533192 245302 533846 245392
rect 533938 245306 534028 249814
rect 534126 249728 534780 249818
rect 534092 245447 534182 249673
rect 534718 245447 534808 249673
rect 534126 245302 534780 245392
rect 533186 245148 534780 245238
rect 534872 245165 534962 249955
rect 535675 245087 535676 250055
rect 536065 245087 536151 250055
rect 537275 245087 537276 250055
rect 537665 245087 537748 250055
rect 553786 249591 553788 249630
rect 553876 249591 553878 249720
rect 561874 249591 561876 249720
rect 561964 249591 561966 249630
rect 553786 249419 553788 249451
rect 553876 249395 553878 249451
rect 561874 249395 561876 249451
rect 561964 249419 561966 249451
rect 553786 249207 553788 249243
rect 553876 249207 553878 249263
rect 561874 249207 561876 249263
rect 561964 249207 561966 249243
rect 553786 249032 553788 249067
rect 553876 248942 553878 249067
rect 561874 248942 561876 249067
rect 561964 249032 561966 249067
rect 545958 248330 548358 248810
rect 545958 248322 546018 248330
rect 548298 248322 548390 248330
rect 545958 247762 548358 248322
rect 553786 247823 553788 247861
rect 553876 247823 553878 247951
rect 561874 247823 561876 247951
rect 561964 247823 561966 247861
rect 553786 247650 553788 247683
rect 553876 247627 553878 247683
rect 561874 247627 561876 247683
rect 561964 247650 561966 247683
rect 553786 247439 553788 247473
rect 553876 247439 553878 247495
rect 561874 247439 561876 247495
rect 561964 247439 561966 247473
rect 545958 246798 548358 247358
rect 553786 247262 553788 247299
rect 553876 247172 553878 247299
rect 561874 247172 561876 247299
rect 561964 247262 561966 247299
rect 545958 246790 546018 246798
rect 548298 246790 548390 246798
rect 545958 246310 548358 246790
rect 553786 246055 553788 246092
rect 553876 246055 553878 246182
rect 561874 246055 561876 246182
rect 561964 246055 561966 246092
rect 553786 245881 553788 245915
rect 553876 245859 553878 245915
rect 561874 245859 561876 245915
rect 561964 245881 561966 245915
rect 553786 245671 553788 245701
rect 553876 245671 553878 245727
rect 561874 245671 561876 245727
rect 561964 245671 561966 245701
rect 553786 245490 553788 245531
rect 553876 245400 553878 245531
rect 561874 245400 561876 245531
rect 561964 245490 561966 245531
rect 57402 245001 59558 245087
rect 62776 245084 63332 245087
rect 65476 245084 66032 245087
rect 62776 245001 66032 245084
rect 529118 245084 529674 245087
rect 531818 245084 532374 245087
rect 529118 245001 532374 245084
rect 535592 245001 537748 245087
rect 57485 244612 57486 245001
rect 59475 244612 59558 245001
rect 57485 244611 59558 244612
rect 62859 244612 62860 245001
rect 65949 244612 66032 245001
rect 69094 244851 69184 244880
rect 62859 244611 66032 244612
rect 529201 244612 529202 245001
rect 532291 244612 532374 245001
rect 529201 244611 532374 244612
rect 535675 244612 535676 245001
rect 537665 244612 537748 245001
rect 535675 244611 537748 244612
rect 33184 244285 33186 244322
rect 33274 244285 33276 244412
rect 41272 244285 41274 244412
rect 41362 244285 41364 244322
rect 47518 244268 49130 244320
rect 546020 244268 547632 244320
rect 553786 244287 553788 244327
rect 553876 244287 553878 244417
rect 561874 244287 561876 244417
rect 561964 244287 561966 244327
rect 33184 244111 33186 244145
rect 33274 244089 33276 244145
rect 41272 244089 41274 244145
rect 41362 244111 41364 244145
rect 66692 244138 66838 244162
rect 553786 244116 553788 244147
rect 553876 244091 553878 244147
rect 561874 244091 561876 244147
rect 561964 244116 561966 244147
rect 33184 243901 33186 243935
rect 33274 243901 33276 243957
rect 41272 243901 41274 243957
rect 41362 243901 41364 243935
rect 553786 243903 553788 243941
rect 553876 243903 553878 243959
rect 561874 243903 561876 243959
rect 561964 243903 561966 243941
rect 47518 243792 49130 243844
rect 546020 243792 547632 243844
rect 33184 243724 33186 243761
rect 33274 243634 33276 243761
rect 41272 243634 41274 243761
rect 41362 243724 41364 243761
rect 553786 243730 553788 243763
rect 553876 243640 553878 243763
rect 561874 243640 561876 243763
rect 561964 243730 561966 243763
rect 57555 242949 57701 242988
rect 59943 242949 60089 242988
rect 33184 242517 33186 242549
rect 33274 242517 33276 242639
rect 41272 242517 41274 242639
rect 41362 242517 41364 242549
rect 553786 242519 553788 242555
rect 553876 242519 553878 242645
rect 561874 242519 561876 242645
rect 561964 242519 561966 242555
rect 33184 242338 33186 242377
rect 33274 242321 33276 242377
rect 41272 242321 41274 242377
rect 41362 242338 41364 242377
rect 553786 242344 553788 242379
rect 553876 242323 553878 242379
rect 561874 242323 561876 242379
rect 561964 242344 561966 242379
rect 17922 242024 17923 242064
rect 18324 242024 18407 242064
rect 27919 242032 28903 242118
rect 566247 242034 567231 242120
rect 17922 242023 18407 242024
rect 28002 242024 28003 242032
rect 28820 242024 28903 242032
rect 566330 242025 566331 242034
rect 567148 242025 567231 242034
rect 566330 242024 567231 242025
rect 576826 242066 577228 253056
rect 576826 242025 576827 242066
rect 577228 242025 577311 242066
rect 576826 242024 577311 242025
rect 28002 242023 28903 242024
rect 46792 241322 49192 241802
rect 545958 241322 548358 241802
rect 46792 241314 46852 241322
rect 49132 241314 49224 241322
rect 545958 241314 546018 241322
rect 548298 241314 548390 241322
rect 46792 240754 49192 241314
rect 545958 240754 548358 241314
rect 46792 233806 49192 234366
rect 545958 233806 548358 234366
rect 46792 233798 46852 233806
rect 49132 233798 49224 233806
rect 545958 233798 546018 233806
rect 548298 233798 548390 233806
rect 46792 233318 49192 233798
rect 545958 233318 548358 233798
rect 17839 233096 18410 233182
rect 27916 233096 28903 233182
rect 566247 233097 567234 233183
rect 576740 233097 577311 233183
rect 17922 233054 17923 233096
rect 18324 233054 18407 233096
rect 28002 233086 28903 233096
rect 566330 233088 567231 233097
rect 576826 233056 576827 233097
rect 577228 233056 577311 233097
rect 17922 231028 18324 233054
rect 576826 231028 577228 233056
rect 17922 222064 18324 224000
rect 17922 222024 17923 222064
rect 18324 222024 18407 222064
rect 27919 222032 28903 222092
rect 566247 222034 567231 222092
rect 17922 222023 18407 222024
rect 28002 222024 28003 222032
rect 28820 222024 28903 222032
rect 566330 222025 566331 222034
rect 567148 222025 567231 222034
rect 566330 222024 567231 222025
rect 576826 222066 577228 224092
rect 576826 222025 576827 222066
rect 577228 222025 577311 222066
rect 576826 222024 577311 222025
rect 28002 222023 28903 222024
rect 46792 221322 49192 221802
rect 545958 221322 548358 221802
rect 46792 221314 46852 221322
rect 49132 221314 49224 221322
rect 545958 221314 546018 221322
rect 548298 221314 548390 221322
rect 46792 220754 49192 221314
rect 545958 220754 548358 221314
rect 46792 213806 49192 214366
rect 46792 213798 46852 213806
rect 49132 213798 49224 213806
rect 46792 213318 49192 213798
rect 17839 213096 18410 213182
rect 27916 213096 28903 213182
rect 17922 213054 17923 213096
rect 18324 213054 18407 213096
rect 28002 213086 28903 213096
rect 17922 202064 18324 213054
rect 33184 212741 33186 212776
rect 33274 212741 33276 212797
rect 41272 212741 41274 212797
rect 41362 212741 41364 212776
rect 33184 212565 33186 212601
rect 33274 212475 33276 212601
rect 41272 212475 41274 212601
rect 41362 212565 41364 212601
rect 33184 211357 33186 211390
rect 33274 211357 33276 211480
rect 41272 211357 41274 211480
rect 41362 211357 41364 211390
rect 47518 211276 49130 211328
rect 33184 211179 33186 211217
rect 33274 211161 33276 211217
rect 41272 211161 41274 211217
rect 41362 211179 41364 211217
rect 33184 210973 33186 211004
rect 33274 210973 33276 211029
rect 41272 210973 41274 211029
rect 41362 210973 41364 211004
rect 33184 210793 33186 210833
rect 33274 210703 33276 210833
rect 41272 210703 41274 210833
rect 41362 210793 41364 210833
rect 47518 210800 49130 210852
rect 57402 210509 59558 210592
rect 62776 210509 66032 210592
rect 57485 210141 57486 210509
rect 59475 210141 59558 210509
rect 62859 210141 62860 210509
rect 65949 210141 66032 210509
rect 57402 210120 57961 210141
rect 58999 210120 59558 210141
rect 57402 210119 59558 210120
rect 57402 210055 57961 210119
rect 58999 210055 59558 210119
rect 62776 210120 63335 210141
rect 65473 210120 66032 210141
rect 62776 210119 66032 210120
rect 62776 210055 63335 210119
rect 65473 210055 66032 210119
rect 33184 209589 33186 209630
rect 33274 209589 33276 209720
rect 41272 209589 41274 209720
rect 41362 209589 41364 209630
rect 33184 209419 33186 209449
rect 33274 209393 33276 209449
rect 41272 209393 41274 209449
rect 41362 209419 41364 209449
rect 33184 209205 33186 209239
rect 33274 209205 33276 209261
rect 41272 209205 41274 209261
rect 41362 209205 41364 209239
rect 33184 209028 33186 209065
rect 33274 208938 33276 209065
rect 41272 208938 41274 209065
rect 41362 209028 41364 209065
rect 46792 208330 49192 208810
rect 46792 208322 46852 208330
rect 49132 208322 49224 208330
rect 33184 207821 33186 207858
rect 33274 207821 33276 207948
rect 41272 207821 41274 207948
rect 41362 207821 41364 207858
rect 46792 207762 49192 208322
rect 33184 207647 33186 207681
rect 33274 207625 33276 207681
rect 41272 207625 41274 207681
rect 41362 207647 41364 207681
rect 33184 207437 33186 207470
rect 33274 207437 33276 207493
rect 41272 207437 41274 207493
rect 41362 207437 41364 207470
rect 33184 207259 33186 207297
rect 33274 207169 33276 207297
rect 41272 207169 41274 207297
rect 41362 207259 41364 207297
rect 46792 206798 49192 207358
rect 46792 206790 46852 206798
rect 49132 206790 49224 206798
rect 46792 206310 49192 206790
rect 33184 206053 33186 206088
rect 33274 206053 33276 206178
rect 41272 206053 41274 206178
rect 41362 206053 41364 206088
rect 33184 205877 33186 205913
rect 33274 205857 33276 205913
rect 41272 205857 41274 205913
rect 41362 205877 41364 205913
rect 33184 205669 33186 205701
rect 33274 205669 33276 205725
rect 41272 205669 41274 205725
rect 41362 205669 41364 205701
rect 33184 205490 33186 205529
rect 33274 205400 33276 205529
rect 41272 205400 41274 205529
rect 41362 205490 41364 205529
rect 57485 205087 57486 210055
rect 57875 205087 57961 210055
rect 59085 205087 59086 210055
rect 59475 205087 59558 210055
rect 60188 205165 60278 209955
rect 60370 209882 61964 209972
rect 60370 209728 61024 209818
rect 60342 205447 60432 209673
rect 60968 205447 61058 209673
rect 60370 205302 61024 205392
rect 61122 205306 61212 209814
rect 61304 209728 61958 209818
rect 61276 205447 61366 209673
rect 61902 205447 61992 209673
rect 61304 205302 61958 205392
rect 60370 205148 61964 205238
rect 62056 205165 62146 209955
rect 62859 205087 62860 210055
rect 63249 210036 63335 210055
rect 63249 205087 63332 210036
rect 65559 205087 65560 210055
rect 65949 205087 66032 210055
rect 69038 205697 69184 205749
rect 57402 205001 59558 205087
rect 62776 205084 63332 205087
rect 65476 205084 66032 205087
rect 62776 205001 66032 205084
rect 57485 204612 57486 205001
rect 59475 204612 59558 205001
rect 57485 204611 59558 204612
rect 62859 204612 62860 205001
rect 65949 204612 66032 205001
rect 69094 204851 69184 204880
rect 62859 204611 66032 204612
rect 33184 204285 33186 204322
rect 33274 204285 33276 204412
rect 41272 204285 41274 204412
rect 41362 204285 41364 204322
rect 47518 204268 49130 204320
rect 33184 204111 33186 204145
rect 33274 204089 33276 204145
rect 41272 204089 41274 204145
rect 41362 204111 41364 204145
rect 66692 204138 66838 204162
rect 33184 203901 33186 203935
rect 33274 203901 33276 203957
rect 41272 203901 41274 203957
rect 41362 203901 41364 203935
rect 47518 203792 49130 203844
rect 33184 203724 33186 203761
rect 33274 203634 33276 203761
rect 41272 203634 41274 203761
rect 41362 203724 41364 203761
rect 57555 202949 57701 202988
rect 59943 202949 60089 202988
rect 33184 202517 33186 202549
rect 33274 202517 33276 202639
rect 41272 202517 41274 202639
rect 41362 202517 41364 202549
rect 33184 202338 33186 202377
rect 33274 202321 33276 202377
rect 41272 202321 41274 202377
rect 41362 202338 41364 202377
rect 17922 202024 17923 202064
rect 18324 202024 18407 202064
rect 27919 202032 28903 202118
rect 17922 202023 18407 202024
rect 28002 202024 28003 202032
rect 28820 202024 28903 202032
rect 28002 202023 28903 202024
rect 46792 201322 49192 201802
rect 46792 201314 46852 201322
rect 49132 201314 49224 201322
rect 46792 200754 49192 201314
rect 46792 193806 49192 194366
rect 46792 193798 46852 193806
rect 49132 193798 49224 193806
rect 46792 193318 49192 193798
rect 17839 193096 18410 193182
rect 27916 193096 28903 193182
rect 17922 193054 17923 193096
rect 18324 193054 18407 193096
rect 28002 193086 28903 193096
rect 17922 191028 18324 193054
rect 17922 182064 18324 184092
rect 17922 182024 17923 182064
rect 18324 182024 18407 182064
rect 27919 182032 28903 182092
rect 17922 182023 18407 182024
rect 28002 182024 28003 182032
rect 28820 182024 28903 182032
rect 28002 182023 28903 182024
rect 46792 181322 49192 181802
rect 46792 181314 46852 181322
rect 49132 181314 49224 181322
rect 46792 180754 49192 181314
rect 545958 133806 548358 134366
rect 545958 133798 546018 133806
rect 548298 133798 548390 133806
rect 545958 133318 548358 133798
rect 566247 133097 567234 133183
rect 576740 133097 577311 133183
rect 566330 133088 567231 133097
rect 576826 133056 576827 133097
rect 577228 133056 577311 133097
rect 576826 131028 577228 133056
rect 566247 122034 567231 122092
rect 566330 122025 566331 122034
rect 567148 122025 567231 122034
rect 566330 122024 567231 122025
rect 576826 122066 577228 124092
rect 576826 122025 576827 122066
rect 577228 122025 577311 122066
rect 576826 122024 577311 122025
rect 545958 121322 548358 121802
rect 545958 121314 546018 121322
rect 548298 121314 548390 121322
rect 545958 120754 548358 121314
rect 545958 113806 548358 114366
rect 545958 113798 546018 113806
rect 548298 113798 548390 113806
rect 545958 113318 548358 113798
rect 566247 113097 567234 113183
rect 576740 113097 577311 113183
rect 566330 113088 567231 113097
rect 576826 113056 576827 113097
rect 577228 113056 577311 113097
rect 553786 112743 553788 112782
rect 553876 112743 553878 112799
rect 561874 112743 561876 112799
rect 561964 112743 561966 112782
rect 553786 112571 553788 112603
rect 553876 112481 553878 112603
rect 561874 112481 561876 112603
rect 561964 112571 561966 112603
rect 535061 112188 535151 112227
rect 537505 112188 537595 112227
rect 553786 111359 553788 111396
rect 553876 111359 553878 111486
rect 561874 111359 561876 111486
rect 561964 111359 561966 111396
rect 546020 111276 547632 111328
rect 553786 111185 553788 111219
rect 553876 111163 553878 111219
rect 561874 111163 561876 111219
rect 561964 111185 561966 111219
rect 528368 111014 528458 111038
rect 553786 110975 553788 111009
rect 553876 110975 553878 111031
rect 561874 110975 561876 111031
rect 561964 110975 561966 111009
rect 546020 110800 547632 110852
rect 553786 110798 553788 110835
rect 553876 110708 553878 110835
rect 561874 110708 561876 110835
rect 561964 110798 561966 110835
rect 530544 110592 531740 110595
rect 529118 110509 532374 110592
rect 535592 110509 537748 110592
rect 525966 110296 526112 110325
rect 529201 110141 529202 110509
rect 532291 110141 532374 110509
rect 535675 110141 535676 110509
rect 537665 110141 537748 110509
rect 529118 110120 529677 110141
rect 531815 110120 532374 110141
rect 529118 110119 532374 110120
rect 529118 110055 529677 110119
rect 531815 110055 532374 110119
rect 535592 110120 536151 110141
rect 537189 110120 537748 110141
rect 535592 110119 537748 110120
rect 535592 110055 536151 110119
rect 537189 110055 537748 110119
rect 525966 109427 526056 109479
rect 529201 105087 529202 110055
rect 529591 110036 529677 110055
rect 529591 105087 529674 110036
rect 531901 105087 531902 110055
rect 532291 105087 532374 110055
rect 533004 105165 533094 109955
rect 533186 109882 534780 109972
rect 533192 109728 533846 109818
rect 533158 105447 533248 109673
rect 533784 105447 533874 109673
rect 533192 105302 533846 105392
rect 533938 105306 534028 109814
rect 534126 109728 534780 109818
rect 534092 105447 534182 109673
rect 534718 105447 534808 109673
rect 534126 105302 534780 105392
rect 533186 105148 534780 105238
rect 534872 105165 534962 109955
rect 535675 105087 535676 110055
rect 536065 105087 536151 110055
rect 537275 105087 537276 110055
rect 537665 105087 537748 110055
rect 553786 109591 553788 109630
rect 553876 109591 553878 109720
rect 561874 109591 561876 109720
rect 561964 109591 561966 109630
rect 553786 109419 553788 109451
rect 553876 109395 553878 109451
rect 561874 109395 561876 109451
rect 561964 109419 561966 109451
rect 553786 109207 553788 109243
rect 553876 109207 553878 109263
rect 561874 109207 561876 109263
rect 561964 109207 561966 109243
rect 553786 109032 553788 109067
rect 553876 108942 553878 109067
rect 561874 108942 561876 109067
rect 561964 109032 561966 109067
rect 545958 108330 548358 108810
rect 545958 108322 546018 108330
rect 548298 108322 548390 108330
rect 545958 107762 548358 108322
rect 553786 107823 553788 107861
rect 553876 107823 553878 107951
rect 561874 107823 561876 107951
rect 561964 107823 561966 107861
rect 553786 107650 553788 107683
rect 553876 107627 553878 107683
rect 561874 107627 561876 107683
rect 561964 107650 561966 107683
rect 553786 107439 553788 107473
rect 553876 107439 553878 107495
rect 561874 107439 561876 107495
rect 561964 107439 561966 107473
rect 545958 106798 548358 107358
rect 553786 107262 553788 107299
rect 553876 107172 553878 107299
rect 561874 107172 561876 107299
rect 561964 107262 561966 107299
rect 545958 106790 546018 106798
rect 548298 106790 548390 106798
rect 545958 106310 548358 106790
rect 553786 106055 553788 106092
rect 553876 106055 553878 106182
rect 561874 106055 561876 106182
rect 561964 106055 561966 106092
rect 553786 105881 553788 105915
rect 553876 105859 553878 105915
rect 561874 105859 561876 105915
rect 561964 105881 561966 105915
rect 553786 105671 553788 105701
rect 553876 105671 553878 105727
rect 561874 105671 561876 105727
rect 561964 105671 561966 105701
rect 553786 105490 553788 105531
rect 553876 105400 553878 105531
rect 561874 105400 561876 105531
rect 561964 105490 561966 105531
rect 529118 105084 529674 105087
rect 531818 105084 532374 105087
rect 529118 105001 532374 105084
rect 535592 105001 537748 105087
rect 529201 104612 529202 105001
rect 532291 104612 532374 105001
rect 529201 104611 532374 104612
rect 535675 104612 535676 105001
rect 537665 104612 537748 105001
rect 535675 104611 537748 104612
rect 546020 104268 547632 104320
rect 553786 104287 553788 104327
rect 553876 104287 553878 104417
rect 561874 104287 561876 104417
rect 561964 104287 561966 104327
rect 553786 104116 553788 104147
rect 553876 104091 553878 104147
rect 561874 104091 561876 104147
rect 561964 104116 561966 104147
rect 553786 103903 553788 103941
rect 553876 103903 553878 103959
rect 561874 103903 561876 103959
rect 561964 103903 561966 103941
rect 546020 103792 547632 103844
rect 553786 103730 553788 103763
rect 553876 103640 553878 103763
rect 561874 103640 561876 103763
rect 561964 103730 561966 103763
rect 553786 102519 553788 102555
rect 553876 102519 553878 102645
rect 561874 102519 561876 102645
rect 561964 102519 561966 102555
rect 553786 102344 553788 102379
rect 553876 102323 553878 102379
rect 561874 102323 561876 102379
rect 561964 102344 561966 102379
rect 566247 102034 567231 102120
rect 566330 102025 566331 102034
rect 567148 102025 567231 102034
rect 566330 102024 567231 102025
rect 576826 102066 577228 113056
rect 576826 102025 576827 102066
rect 577228 102025 577311 102066
rect 576826 102024 577311 102025
rect 545958 101322 548358 101802
rect 545958 101314 546018 101322
rect 548298 101314 548390 101322
rect 545958 100754 548358 101314
rect 545958 93806 548358 94366
rect 545958 93798 546018 93806
rect 548298 93798 548390 93806
rect 545958 93318 548358 93798
rect 566247 93097 567234 93183
rect 576740 93097 577311 93183
rect 566330 93088 567231 93097
rect 576826 93056 576827 93097
rect 577228 93056 577311 93097
rect 553786 92743 553788 92782
rect 553876 92743 553878 92799
rect 561874 92743 561876 92799
rect 561964 92743 561966 92782
rect 553786 92571 553788 92603
rect 553876 92481 553878 92603
rect 561874 92481 561876 92603
rect 561964 92571 561966 92603
rect 535061 92188 535151 92227
rect 537505 92188 537595 92227
rect 553786 91359 553788 91396
rect 553876 91359 553878 91486
rect 561874 91359 561876 91486
rect 561964 91359 561966 91396
rect 546020 91276 547632 91328
rect 553786 91185 553788 91219
rect 553876 91163 553878 91219
rect 561874 91163 561876 91219
rect 561964 91185 561966 91219
rect 528368 91014 528458 91038
rect 553786 90975 553788 91009
rect 553876 90975 553878 91031
rect 561874 90975 561876 91031
rect 561964 90975 561966 91009
rect 546020 90800 547632 90852
rect 553786 90798 553788 90835
rect 553876 90708 553878 90835
rect 561874 90708 561876 90835
rect 561964 90798 561966 90835
rect 530544 90592 531740 90595
rect 529118 90509 532374 90592
rect 535592 90509 537748 90592
rect 525966 90296 526112 90325
rect 529201 90141 529202 90509
rect 532291 90141 532374 90509
rect 535675 90141 535676 90509
rect 537665 90141 537748 90509
rect 529118 90120 529677 90141
rect 531815 90120 532374 90141
rect 529118 90119 532374 90120
rect 529118 90055 529677 90119
rect 531815 90055 532374 90119
rect 535592 90120 536151 90141
rect 537189 90120 537748 90141
rect 535592 90119 537748 90120
rect 535592 90055 536151 90119
rect 537189 90055 537748 90119
rect 525966 89427 526056 89479
rect 529201 85087 529202 90055
rect 529591 90036 529677 90055
rect 529591 85087 529674 90036
rect 531901 85087 531902 90055
rect 532291 85087 532374 90055
rect 533004 85165 533094 89955
rect 533186 89882 534780 89972
rect 533192 89728 533846 89818
rect 533158 85447 533248 89673
rect 533784 85447 533874 89673
rect 533192 85302 533846 85392
rect 533938 85306 534028 89814
rect 534126 89728 534780 89818
rect 534092 85447 534182 89673
rect 534718 85447 534808 89673
rect 534126 85302 534780 85392
rect 533186 85148 534780 85238
rect 534872 85165 534962 89955
rect 535675 85087 535676 90055
rect 536065 85087 536151 90055
rect 537275 85087 537276 90055
rect 537665 85087 537748 90055
rect 553786 89591 553788 89630
rect 553876 89591 553878 89720
rect 561874 89591 561876 89720
rect 561964 89591 561966 89630
rect 553786 89419 553788 89451
rect 553876 89395 553878 89451
rect 561874 89395 561876 89451
rect 561964 89419 561966 89451
rect 553786 89207 553788 89243
rect 553876 89207 553878 89263
rect 561874 89207 561876 89263
rect 561964 89207 561966 89243
rect 553786 89032 553788 89067
rect 553876 88942 553878 89067
rect 561874 88942 561876 89067
rect 561964 89032 561966 89067
rect 545958 88330 548358 88810
rect 545958 88322 546018 88330
rect 548298 88322 548390 88330
rect 545958 87762 548358 88322
rect 553786 87823 553788 87861
rect 553876 87823 553878 87951
rect 561874 87823 561876 87951
rect 561964 87823 561966 87861
rect 553786 87650 553788 87683
rect 553876 87627 553878 87683
rect 561874 87627 561876 87683
rect 561964 87650 561966 87683
rect 553786 87439 553788 87473
rect 553876 87439 553878 87495
rect 561874 87439 561876 87495
rect 561964 87439 561966 87473
rect 545958 86798 548358 87358
rect 553786 87262 553788 87299
rect 553876 87172 553878 87299
rect 561874 87172 561876 87299
rect 561964 87262 561966 87299
rect 545958 86790 546018 86798
rect 548298 86790 548390 86798
rect 545958 86310 548358 86790
rect 553786 86055 553788 86092
rect 553876 86055 553878 86182
rect 561874 86055 561876 86182
rect 561964 86055 561966 86092
rect 553786 85881 553788 85915
rect 553876 85859 553878 85915
rect 561874 85859 561876 85915
rect 561964 85881 561966 85915
rect 553786 85671 553788 85701
rect 553876 85671 553878 85727
rect 561874 85671 561876 85727
rect 561964 85671 561966 85701
rect 553786 85490 553788 85531
rect 553876 85400 553878 85531
rect 561874 85400 561876 85531
rect 561964 85490 561966 85531
rect 529118 85084 529674 85087
rect 531818 85084 532374 85087
rect 529118 85001 532374 85084
rect 535592 85001 537748 85087
rect 529201 84612 529202 85001
rect 532291 84612 532374 85001
rect 529201 84611 532374 84612
rect 535675 84612 535676 85001
rect 537665 84612 537748 85001
rect 535675 84611 537748 84612
rect 546020 84268 547632 84320
rect 553786 84287 553788 84327
rect 553876 84287 553878 84417
rect 561874 84287 561876 84417
rect 561964 84287 561966 84327
rect 553786 84116 553788 84147
rect 553876 84091 553878 84147
rect 561874 84091 561876 84147
rect 561964 84116 561966 84147
rect 553786 83903 553788 83941
rect 553876 83903 553878 83959
rect 561874 83903 561876 83959
rect 561964 83903 561966 83941
rect 546020 83792 547632 83844
rect 553786 83730 553788 83763
rect 553876 83640 553878 83763
rect 561874 83640 561876 83763
rect 561964 83730 561966 83763
rect 553786 82519 553788 82555
rect 553876 82519 553878 82645
rect 561874 82519 561876 82645
rect 561964 82519 561966 82555
rect 553786 82344 553788 82379
rect 553876 82323 553878 82379
rect 561874 82323 561876 82379
rect 561964 82344 561966 82379
rect 566247 82034 567231 82120
rect 566330 82025 566331 82034
rect 567148 82025 567231 82034
rect 566330 82024 567231 82025
rect 576826 82066 577228 93056
rect 576826 82025 576827 82066
rect 577228 82025 577311 82066
rect 576826 82024 577311 82025
rect 545958 81322 548358 81802
rect 545958 81314 546018 81322
rect 548298 81314 548390 81322
rect 545958 80754 548358 81314
rect 17157 75060 73873 75113
rect 521418 75060 577624 75112
rect 75060 17496 75112 73702
rect 209427 69064 209479 69154
rect 210296 69064 210325 69154
rect 249427 69064 249479 69154
rect 250296 69064 250325 69154
rect 269427 69064 269479 69154
rect 270296 69064 270325 69154
rect 309427 69064 309479 69154
rect 310296 69064 310325 69154
rect 329427 69064 329479 69154
rect 330296 69064 330325 69154
rect 369427 69064 369479 69154
rect 370296 69064 370325 69154
rect 409427 69064 409479 69154
rect 410296 69064 410325 69154
rect 429427 69064 429479 69154
rect 430296 69064 430325 69154
rect 469427 69064 469479 69154
rect 470296 69064 470325 69154
rect 210958 66752 210982 66808
rect 250958 66752 250982 66808
rect 270958 66752 270982 66808
rect 310958 66752 310982 66808
rect 330958 66752 330982 66808
rect 370958 66752 370982 66808
rect 410958 66752 410982 66808
rect 430958 66752 430982 66808
rect 470958 66752 470982 66808
rect 211014 66662 211038 66752
rect 251014 66662 251038 66752
rect 271014 66662 271038 66752
rect 311014 66662 311038 66752
rect 331014 66662 331038 66752
rect 371014 66662 371038 66752
rect 411014 66662 411038 66752
rect 431014 66662 431038 66752
rect 471014 66662 471038 66752
rect 204528 65919 210592 66002
rect 244528 65919 250592 66002
rect 264528 65919 270592 66002
rect 304528 65919 310592 66002
rect 324528 65919 330592 66002
rect 364528 65919 370592 66002
rect 404528 65919 410592 66002
rect 424528 65919 430592 66002
rect 464528 65919 470592 66002
rect 204611 62830 204612 65919
rect 205001 65530 205087 65919
rect 210055 65530 210141 65919
rect 205001 65529 210141 65530
rect 205001 65446 205087 65529
rect 205001 63305 205084 65446
rect 210119 63305 210120 65529
rect 210509 64576 210592 65919
rect 210509 63380 210595 64576
rect 204979 63302 205084 63305
rect 210036 63302 210141 63305
rect 204979 63219 210141 63302
rect 205001 62830 205087 63219
rect 210055 62830 210141 63219
rect 210509 62830 210592 63380
rect 204611 62829 210592 62830
rect 244611 62830 244612 65919
rect 245001 65530 245087 65919
rect 250055 65530 250141 65919
rect 245001 65529 250141 65530
rect 245001 65446 245087 65529
rect 245001 63305 245084 65446
rect 250119 63305 250120 65529
rect 250509 64576 250592 65919
rect 250509 63380 250595 64576
rect 244979 63302 245084 63305
rect 250036 63302 250141 63305
rect 244979 63219 250141 63302
rect 245001 62830 245087 63219
rect 250055 62830 250141 63219
rect 250509 62830 250592 63380
rect 244611 62829 250592 62830
rect 264611 62830 264612 65919
rect 265001 65530 265087 65919
rect 270055 65530 270141 65919
rect 265001 65529 270141 65530
rect 265001 65446 265087 65529
rect 265001 63305 265084 65446
rect 270119 63305 270120 65529
rect 270509 64576 270592 65919
rect 270509 63380 270595 64576
rect 264979 63302 265084 63305
rect 270036 63302 270141 63305
rect 264979 63219 270141 63302
rect 265001 62830 265087 63219
rect 270055 62830 270141 63219
rect 270509 62830 270592 63380
rect 264611 62829 270592 62830
rect 304611 62830 304612 65919
rect 305001 65530 305087 65919
rect 310055 65530 310141 65919
rect 305001 65529 310141 65530
rect 305001 65446 305087 65529
rect 305001 63305 305084 65446
rect 310119 63305 310120 65529
rect 310509 64576 310592 65919
rect 310509 63380 310595 64576
rect 304979 63302 305084 63305
rect 310036 63302 310141 63305
rect 304979 63219 310141 63302
rect 305001 62830 305087 63219
rect 310055 62830 310141 63219
rect 310509 62830 310592 63380
rect 304611 62829 310592 62830
rect 324611 62830 324612 65919
rect 325001 65530 325087 65919
rect 330055 65530 330141 65919
rect 325001 65529 330141 65530
rect 325001 65446 325087 65529
rect 325001 63305 325084 65446
rect 330119 63305 330120 65529
rect 330509 64576 330592 65919
rect 330509 63380 330595 64576
rect 324979 63302 325084 63305
rect 330036 63302 330141 63305
rect 324979 63219 330141 63302
rect 325001 62830 325087 63219
rect 330055 62830 330141 63219
rect 330509 62830 330592 63380
rect 324611 62829 330592 62830
rect 364611 62830 364612 65919
rect 365001 65530 365087 65919
rect 370055 65530 370141 65919
rect 365001 65529 370141 65530
rect 365001 65446 365087 65529
rect 365001 63305 365084 65446
rect 370119 63305 370120 65529
rect 370509 64576 370592 65919
rect 370509 63380 370595 64576
rect 364979 63302 365084 63305
rect 370036 63302 370141 63305
rect 364979 63219 370141 63302
rect 365001 62830 365087 63219
rect 370055 62830 370141 63219
rect 370509 62830 370592 63380
rect 364611 62829 370592 62830
rect 404611 62830 404612 65919
rect 405001 65530 405087 65919
rect 410055 65530 410141 65919
rect 405001 65529 410141 65530
rect 405001 65446 405087 65529
rect 405001 63305 405084 65446
rect 410119 63305 410120 65529
rect 410509 64576 410592 65919
rect 410509 63380 410595 64576
rect 404979 63302 405084 63305
rect 410036 63302 410141 63305
rect 404979 63219 410141 63302
rect 405001 62830 405087 63219
rect 410055 62830 410141 63219
rect 410509 62830 410592 63380
rect 404611 62829 410592 62830
rect 424611 62830 424612 65919
rect 425001 65530 425087 65919
rect 430055 65530 430141 65919
rect 425001 65529 430141 65530
rect 425001 65446 425087 65529
rect 425001 63305 425084 65446
rect 430119 63305 430120 65529
rect 430509 64576 430592 65919
rect 430509 63380 430595 64576
rect 424979 63302 425084 63305
rect 430036 63302 430141 63305
rect 424979 63219 430141 63302
rect 425001 62830 425087 63219
rect 430055 62830 430141 63219
rect 430509 62830 430592 63380
rect 424611 62829 430592 62830
rect 464611 62830 464612 65919
rect 465001 65530 465087 65919
rect 470055 65530 470141 65919
rect 465001 65529 470141 65530
rect 465001 65446 465087 65529
rect 465001 63305 465084 65446
rect 470119 63305 470120 65529
rect 470509 64576 470592 65919
rect 470509 63380 470595 64576
rect 464979 63302 465084 63305
rect 470036 63302 470141 63305
rect 464979 63219 470141 63302
rect 465001 62830 465087 63219
rect 470055 62830 470141 63219
rect 470509 62830 470592 63380
rect 464611 62829 470592 62830
rect 205165 62026 209955 62116
rect 245165 62026 249955 62116
rect 265165 62026 269955 62116
rect 305165 62026 309955 62116
rect 325165 62026 329955 62116
rect 365165 62026 369955 62116
rect 405165 62026 409955 62116
rect 425165 62026 429955 62116
rect 465165 62026 469955 62116
rect 205148 60340 205238 61934
rect 205302 61274 205392 61928
rect 205447 61872 209673 61962
rect 205447 61246 209673 61336
rect 209728 61274 209818 61928
rect 205306 61092 209814 61182
rect 205302 60340 205392 60994
rect 205447 60938 209673 61028
rect 205447 60312 209673 60402
rect 209728 60340 209818 60994
rect 209882 60340 209972 61934
rect 245148 60340 245238 61934
rect 245302 61274 245392 61928
rect 245447 61872 249673 61962
rect 245447 61246 249673 61336
rect 249728 61274 249818 61928
rect 245306 61092 249814 61182
rect 245302 60340 245392 60994
rect 245447 60938 249673 61028
rect 245447 60312 249673 60402
rect 249728 60340 249818 60994
rect 249882 60340 249972 61934
rect 265148 60340 265238 61934
rect 265302 61274 265392 61928
rect 265447 61872 269673 61962
rect 265447 61246 269673 61336
rect 269728 61274 269818 61928
rect 265306 61092 269814 61182
rect 265302 60340 265392 60994
rect 265447 60938 269673 61028
rect 265447 60312 269673 60402
rect 269728 60340 269818 60994
rect 269882 60340 269972 61934
rect 305148 60340 305238 61934
rect 305302 61274 305392 61928
rect 305447 61872 309673 61962
rect 305447 61246 309673 61336
rect 309728 61274 309818 61928
rect 305306 61092 309814 61182
rect 305302 60340 305392 60994
rect 305447 60938 309673 61028
rect 305447 60312 309673 60402
rect 309728 60340 309818 60994
rect 309882 60340 309972 61934
rect 325148 60340 325238 61934
rect 325302 61274 325392 61928
rect 325447 61872 329673 61962
rect 325447 61246 329673 61336
rect 329728 61274 329818 61928
rect 325306 61092 329814 61182
rect 325302 60340 325392 60994
rect 325447 60938 329673 61028
rect 325447 60312 329673 60402
rect 329728 60340 329818 60994
rect 329882 60340 329972 61934
rect 365148 60340 365238 61934
rect 365302 61274 365392 61928
rect 365447 61872 369673 61962
rect 365447 61246 369673 61336
rect 369728 61274 369818 61928
rect 365306 61092 369814 61182
rect 365302 60340 365392 60994
rect 365447 60938 369673 61028
rect 365447 60312 369673 60402
rect 369728 60340 369818 60994
rect 369882 60340 369972 61934
rect 405148 60340 405238 61934
rect 405302 61274 405392 61928
rect 405447 61872 409673 61962
rect 405447 61246 409673 61336
rect 409728 61274 409818 61928
rect 405306 61092 409814 61182
rect 405302 60340 405392 60994
rect 405447 60938 409673 61028
rect 405447 60312 409673 60402
rect 409728 60340 409818 60994
rect 409882 60340 409972 61934
rect 425148 60340 425238 61934
rect 425302 61274 425392 61928
rect 425447 61872 429673 61962
rect 425447 61246 429673 61336
rect 429728 61274 429818 61928
rect 425306 61092 429814 61182
rect 425302 60340 425392 60994
rect 425447 60938 429673 61028
rect 425447 60312 429673 60402
rect 429728 60340 429818 60994
rect 429882 60340 429972 61934
rect 465148 60340 465238 61934
rect 465302 61274 465392 61928
rect 465447 61872 469673 61962
rect 465447 61246 469673 61336
rect 469728 61274 469818 61928
rect 465306 61092 469814 61182
rect 465302 60340 465392 60994
rect 465447 60938 469673 61028
rect 465447 60312 469673 60402
rect 469728 60340 469818 60994
rect 469882 60340 469972 61934
rect 205165 60158 209955 60248
rect 245165 60158 249955 60248
rect 265165 60158 269955 60248
rect 305165 60158 309955 60248
rect 325165 60158 329955 60248
rect 365165 60158 369955 60248
rect 405165 60158 409955 60248
rect 425165 60158 429955 60248
rect 465165 60158 469955 60248
rect 212188 59969 212227 60059
rect 252188 59969 252227 60059
rect 272188 59969 272227 60059
rect 312188 59969 312227 60059
rect 332188 59969 332227 60059
rect 372188 59969 372227 60059
rect 412188 59969 412227 60059
rect 432188 59969 432227 60059
rect 472188 59969 472227 60059
rect 204528 59445 210592 59528
rect 244528 59445 250592 59528
rect 264528 59445 270592 59528
rect 304528 59445 310592 59528
rect 324528 59445 330592 59528
rect 364528 59445 370592 59528
rect 404528 59445 410592 59528
rect 424528 59445 430592 59528
rect 464528 59445 470592 59528
rect 204611 57456 204612 59445
rect 205001 59056 205087 59445
rect 210055 59056 210141 59445
rect 205001 59055 210141 59056
rect 205001 57931 205087 59055
rect 210119 57931 210120 59055
rect 204979 57845 210141 57931
rect 205001 57456 205087 57845
rect 210055 57456 210141 57845
rect 210509 57456 210592 59445
rect 212132 57615 212171 57671
rect 212188 57525 212227 57615
rect 204611 57455 210592 57456
rect 244611 57456 244612 59445
rect 245001 59056 245087 59445
rect 250055 59056 250141 59445
rect 245001 59055 250141 59056
rect 245001 57931 245087 59055
rect 250119 57931 250120 59055
rect 244979 57845 250141 57931
rect 245001 57456 245087 57845
rect 250055 57456 250141 57845
rect 250509 57456 250592 59445
rect 252132 57615 252171 57671
rect 252188 57525 252227 57615
rect 244611 57455 250592 57456
rect 264611 57456 264612 59445
rect 265001 59056 265087 59445
rect 270055 59056 270141 59445
rect 265001 59055 270141 59056
rect 265001 57931 265087 59055
rect 270119 57931 270120 59055
rect 264979 57845 270141 57931
rect 265001 57456 265087 57845
rect 270055 57456 270141 57845
rect 270509 57456 270592 59445
rect 272132 57615 272171 57671
rect 272188 57525 272227 57615
rect 264611 57455 270592 57456
rect 304611 57456 304612 59445
rect 305001 59056 305087 59445
rect 310055 59056 310141 59445
rect 305001 59055 310141 59056
rect 305001 57931 305087 59055
rect 310119 57931 310120 59055
rect 304979 57845 310141 57931
rect 305001 57456 305087 57845
rect 310055 57456 310141 57845
rect 310509 57456 310592 59445
rect 312132 57615 312171 57671
rect 312188 57525 312227 57615
rect 304611 57455 310592 57456
rect 324611 57456 324612 59445
rect 325001 59056 325087 59445
rect 330055 59056 330141 59445
rect 325001 59055 330141 59056
rect 325001 57931 325087 59055
rect 330119 57931 330120 59055
rect 324979 57845 330141 57931
rect 325001 57456 325087 57845
rect 330055 57456 330141 57845
rect 330509 57456 330592 59445
rect 332132 57615 332171 57671
rect 332188 57525 332227 57615
rect 324611 57455 330592 57456
rect 364611 57456 364612 59445
rect 365001 59056 365087 59445
rect 370055 59056 370141 59445
rect 365001 59055 370141 59056
rect 365001 57931 365087 59055
rect 370119 57931 370120 59055
rect 364979 57845 370141 57931
rect 365001 57456 365087 57845
rect 370055 57456 370141 57845
rect 370509 57456 370592 59445
rect 372132 57615 372171 57671
rect 372188 57525 372227 57615
rect 364611 57455 370592 57456
rect 404611 57456 404612 59445
rect 405001 59056 405087 59445
rect 410055 59056 410141 59445
rect 405001 59055 410141 59056
rect 405001 57931 405087 59055
rect 410119 57931 410120 59055
rect 404979 57845 410141 57931
rect 405001 57456 405087 57845
rect 410055 57456 410141 57845
rect 410509 57456 410592 59445
rect 412132 57615 412171 57671
rect 412188 57525 412227 57615
rect 404611 57455 410592 57456
rect 424611 57456 424612 59445
rect 425001 59056 425087 59445
rect 430055 59056 430141 59445
rect 425001 59055 430141 59056
rect 425001 57931 425087 59055
rect 430119 57931 430120 59055
rect 424979 57845 430141 57931
rect 425001 57456 425087 57845
rect 430055 57456 430141 57845
rect 430509 57456 430592 59445
rect 432132 57615 432171 57671
rect 432188 57525 432227 57615
rect 424611 57455 430592 57456
rect 464611 57456 464612 59445
rect 465001 59056 465087 59445
rect 470055 59056 470141 59445
rect 465001 59055 470141 59056
rect 465001 57931 465087 59055
rect 470119 57931 470120 59055
rect 464979 57845 470141 57931
rect 465001 57456 465087 57845
rect 470055 57456 470141 57845
rect 470509 57456 470592 59445
rect 472132 57615 472171 57671
rect 472188 57525 472227 57615
rect 464611 57455 470592 57456
rect 201314 49162 201322 49194
rect 206790 49162 206798 49194
rect 208322 49162 208330 49194
rect 213798 49162 213806 49194
rect 221314 49162 221322 49194
rect 233798 49162 233806 49194
rect 241314 49162 241322 49194
rect 246790 49162 246798 49194
rect 248322 49162 248330 49194
rect 253798 49162 253806 49194
rect 261314 49162 261322 49194
rect 266790 49162 266798 49194
rect 268322 49162 268330 49194
rect 273798 49162 273806 49194
rect 301314 49162 301322 49194
rect 306790 49162 306798 49194
rect 308322 49162 308330 49194
rect 313798 49162 313806 49194
rect 321314 49162 321322 49194
rect 326790 49162 326798 49194
rect 328322 49162 328330 49194
rect 333798 49162 333806 49194
rect 341314 49162 341322 49194
rect 353798 49162 353806 49194
rect 361314 49162 361322 49194
rect 366790 49162 366798 49194
rect 368322 49162 368330 49194
rect 373798 49162 373806 49194
rect 401314 49162 401322 49194
rect 406790 49162 406798 49194
rect 408322 49162 408330 49194
rect 413798 49162 413806 49194
rect 421314 49162 421322 49194
rect 426790 49162 426798 49194
rect 428322 49162 428330 49194
rect 433798 49162 433806 49194
rect 441314 49162 441322 49194
rect 453798 49162 453806 49194
rect 461314 49162 461322 49194
rect 466790 49162 466798 49194
rect 468322 49162 468330 49194
rect 473798 49162 473806 49194
rect 501314 49162 501322 49194
rect 513798 49162 513806 49194
rect 200754 49102 201802 49162
rect 200754 46822 201314 49102
rect 201322 46822 201802 49102
rect 206310 49102 207358 49162
rect 203792 47488 203844 49100
rect 204268 47488 204320 49100
rect 200754 46762 201802 46822
rect 206310 46822 206790 49102
rect 206798 46822 207358 49102
rect 206310 46762 207358 46822
rect 207762 49102 208810 49162
rect 207762 46822 208322 49102
rect 208330 46822 208810 49102
rect 213318 49102 214366 49162
rect 210800 47488 210852 49100
rect 211276 47488 211328 49100
rect 207762 46762 208810 46822
rect 213318 46822 213798 49102
rect 213806 46822 214366 49102
rect 213318 46762 214366 46822
rect 220754 49102 221802 49162
rect 220754 46822 221314 49102
rect 221322 46822 221802 49102
rect 220754 46762 221802 46822
rect 233318 49102 234366 49162
rect 233318 46822 233798 49102
rect 233806 46822 234366 49102
rect 233318 46762 234366 46822
rect 240754 49102 241802 49162
rect 240754 46822 241314 49102
rect 241322 46822 241802 49102
rect 246310 49102 247358 49162
rect 243792 47488 243844 49100
rect 244268 47488 244320 49100
rect 240754 46762 241802 46822
rect 246310 46822 246790 49102
rect 246798 46822 247358 49102
rect 246310 46762 247358 46822
rect 247762 49102 248810 49162
rect 247762 46822 248322 49102
rect 248330 46822 248810 49102
rect 253318 49102 254366 49162
rect 250800 47488 250852 49100
rect 251276 47488 251328 49100
rect 247762 46762 248810 46822
rect 253318 46822 253798 49102
rect 253806 46822 254366 49102
rect 253318 46762 254366 46822
rect 260754 49102 261802 49162
rect 260754 46822 261314 49102
rect 261322 46822 261802 49102
rect 266310 49102 267358 49162
rect 263792 47488 263844 49100
rect 264268 47488 264320 49100
rect 260754 46762 261802 46822
rect 266310 46822 266790 49102
rect 266798 46822 267358 49102
rect 266310 46762 267358 46822
rect 267762 49102 268810 49162
rect 267762 46822 268322 49102
rect 268330 46822 268810 49102
rect 273318 49102 274366 49162
rect 270800 47488 270852 49100
rect 271276 47488 271328 49100
rect 267762 46762 268810 46822
rect 273318 46822 273798 49102
rect 273806 46822 274366 49102
rect 273318 46762 274366 46822
rect 300754 49102 301802 49162
rect 300754 46822 301314 49102
rect 301322 46822 301802 49102
rect 306310 49102 307358 49162
rect 303792 47488 303844 49100
rect 304268 47488 304320 49100
rect 300754 46762 301802 46822
rect 306310 46822 306790 49102
rect 306798 46822 307358 49102
rect 306310 46762 307358 46822
rect 307762 49102 308810 49162
rect 307762 46822 308322 49102
rect 308330 46822 308810 49102
rect 313318 49102 314366 49162
rect 310800 47488 310852 49100
rect 311276 47488 311328 49100
rect 307762 46762 308810 46822
rect 313318 46822 313798 49102
rect 313806 46822 314366 49102
rect 313318 46762 314366 46822
rect 320754 49102 321802 49162
rect 320754 46822 321314 49102
rect 321322 46822 321802 49102
rect 326310 49102 327358 49162
rect 323792 47488 323844 49100
rect 324268 47488 324320 49100
rect 320754 46762 321802 46822
rect 326310 46822 326790 49102
rect 326798 46822 327358 49102
rect 326310 46762 327358 46822
rect 327762 49102 328810 49162
rect 327762 46822 328322 49102
rect 328330 46822 328810 49102
rect 333318 49102 334366 49162
rect 330800 47488 330852 49100
rect 331276 47488 331328 49100
rect 327762 46762 328810 46822
rect 333318 46822 333798 49102
rect 333806 46822 334366 49102
rect 333318 46762 334366 46822
rect 340754 49102 341802 49162
rect 340754 46822 341314 49102
rect 341322 46822 341802 49102
rect 340754 46762 341802 46822
rect 353318 49102 354366 49162
rect 353318 46822 353798 49102
rect 353806 46822 354366 49102
rect 353318 46762 354366 46822
rect 360754 49102 361802 49162
rect 360754 46822 361314 49102
rect 361322 46822 361802 49102
rect 366310 49102 367358 49162
rect 363792 47488 363844 49100
rect 364268 47488 364320 49100
rect 360754 46762 361802 46822
rect 366310 46822 366790 49102
rect 366798 46822 367358 49102
rect 366310 46762 367358 46822
rect 367762 49102 368810 49162
rect 367762 46822 368322 49102
rect 368330 46822 368810 49102
rect 373318 49102 374366 49162
rect 370800 47488 370852 49100
rect 371276 47488 371328 49100
rect 367762 46762 368810 46822
rect 373318 46822 373798 49102
rect 373806 46822 374366 49102
rect 373318 46762 374366 46822
rect 400754 49102 401802 49162
rect 400754 46822 401314 49102
rect 401322 46822 401802 49102
rect 406310 49102 407358 49162
rect 403792 47488 403844 49100
rect 404268 47488 404320 49100
rect 400754 46762 401802 46822
rect 406310 46822 406790 49102
rect 406798 46822 407358 49102
rect 406310 46762 407358 46822
rect 407762 49102 408810 49162
rect 407762 46822 408322 49102
rect 408330 46822 408810 49102
rect 413318 49102 414366 49162
rect 410800 47488 410852 49100
rect 411276 47488 411328 49100
rect 407762 46762 408810 46822
rect 413318 46822 413798 49102
rect 413806 46822 414366 49102
rect 413318 46762 414366 46822
rect 420754 49102 421802 49162
rect 420754 46822 421314 49102
rect 421322 46822 421802 49102
rect 426310 49102 427358 49162
rect 423792 47488 423844 49100
rect 424268 47488 424320 49100
rect 420754 46762 421802 46822
rect 426310 46822 426790 49102
rect 426798 46822 427358 49102
rect 426310 46762 427358 46822
rect 427762 49102 428810 49162
rect 427762 46822 428322 49102
rect 428330 46822 428810 49102
rect 433318 49102 434366 49162
rect 430800 47488 430852 49100
rect 431276 47488 431328 49100
rect 427762 46762 428810 46822
rect 433318 46822 433798 49102
rect 433806 46822 434366 49102
rect 433318 46762 434366 46822
rect 440754 49102 441802 49162
rect 440754 46822 441314 49102
rect 441322 46822 441802 49102
rect 440754 46762 441802 46822
rect 453318 49102 454366 49162
rect 453318 46822 453798 49102
rect 453806 46822 454366 49102
rect 453318 46762 454366 46822
rect 460754 49102 461802 49162
rect 460754 46822 461314 49102
rect 461322 46822 461802 49102
rect 466310 49102 467358 49162
rect 463792 47488 463844 49100
rect 464268 47488 464320 49100
rect 460754 46762 461802 46822
rect 466310 46822 466790 49102
rect 466798 46822 467358 49102
rect 466310 46762 467358 46822
rect 467762 49102 468810 49162
rect 467762 46822 468322 49102
rect 468330 46822 468810 49102
rect 473318 49102 474366 49162
rect 470800 47488 470852 49100
rect 471276 47488 471328 49100
rect 467762 46762 468810 46822
rect 473318 46822 473798 49102
rect 473806 46822 474366 49102
rect 473318 46762 474366 46822
rect 500754 49102 501802 49162
rect 500754 46822 501314 49102
rect 501322 46822 501802 49102
rect 500754 46762 501802 46822
rect 513318 49102 514366 49162
rect 513318 46822 513798 49102
rect 513806 46822 514366 49102
rect 513318 46762 514366 46822
rect 202344 41332 202379 41334
rect 202519 41332 202555 41334
rect 203730 41332 203763 41334
rect 203903 41332 203941 41334
rect 204116 41332 204147 41334
rect 204287 41332 204327 41334
rect 205490 41332 205531 41334
rect 205671 41332 205701 41334
rect 205881 41332 205915 41334
rect 206055 41332 206092 41334
rect 207262 41332 207299 41334
rect 207439 41332 207473 41334
rect 207650 41332 207683 41334
rect 207823 41332 207861 41334
rect 209032 41332 209067 41334
rect 209207 41332 209243 41334
rect 209419 41332 209451 41334
rect 209591 41332 209630 41334
rect 210798 41332 210835 41334
rect 210975 41332 211009 41334
rect 211185 41332 211219 41334
rect 211359 41332 211396 41334
rect 212571 41332 212603 41334
rect 212743 41332 212782 41334
rect 242344 41332 242379 41334
rect 242519 41332 242555 41334
rect 243730 41332 243763 41334
rect 243903 41332 243941 41334
rect 244116 41332 244147 41334
rect 244287 41332 244327 41334
rect 245490 41332 245531 41334
rect 245671 41332 245701 41334
rect 245881 41332 245915 41334
rect 246055 41332 246092 41334
rect 247262 41332 247299 41334
rect 247439 41332 247473 41334
rect 247650 41332 247683 41334
rect 247823 41332 247861 41334
rect 249032 41332 249067 41334
rect 249207 41332 249243 41334
rect 249419 41332 249451 41334
rect 249591 41332 249630 41334
rect 250798 41332 250835 41334
rect 250975 41332 251009 41334
rect 251185 41332 251219 41334
rect 251359 41332 251396 41334
rect 252571 41332 252603 41334
rect 252743 41332 252782 41334
rect 262344 41332 262379 41334
rect 262519 41332 262555 41334
rect 263730 41332 263763 41334
rect 263903 41332 263941 41334
rect 264116 41332 264147 41334
rect 264287 41332 264327 41334
rect 265490 41332 265531 41334
rect 265671 41332 265701 41334
rect 265881 41332 265915 41334
rect 266055 41332 266092 41334
rect 267262 41332 267299 41334
rect 267439 41332 267473 41334
rect 267650 41332 267683 41334
rect 267823 41332 267861 41334
rect 269032 41332 269067 41334
rect 269207 41332 269243 41334
rect 269419 41332 269451 41334
rect 269591 41332 269630 41334
rect 270798 41332 270835 41334
rect 270975 41332 271009 41334
rect 271185 41332 271219 41334
rect 271359 41332 271396 41334
rect 272571 41332 272603 41334
rect 272743 41332 272782 41334
rect 302344 41332 302379 41334
rect 302519 41332 302555 41334
rect 303730 41332 303763 41334
rect 303903 41332 303941 41334
rect 304116 41332 304147 41334
rect 304287 41332 304327 41334
rect 305490 41332 305531 41334
rect 305671 41332 305701 41334
rect 305881 41332 305915 41334
rect 306055 41332 306092 41334
rect 307262 41332 307299 41334
rect 307439 41332 307473 41334
rect 307650 41332 307683 41334
rect 307823 41332 307861 41334
rect 309032 41332 309067 41334
rect 309207 41332 309243 41334
rect 309419 41332 309451 41334
rect 309591 41332 309630 41334
rect 310798 41332 310835 41334
rect 310975 41332 311009 41334
rect 311185 41332 311219 41334
rect 311359 41332 311396 41334
rect 312571 41332 312603 41334
rect 312743 41332 312782 41334
rect 322344 41332 322379 41334
rect 322519 41332 322555 41334
rect 323730 41332 323763 41334
rect 323903 41332 323941 41334
rect 324116 41332 324147 41334
rect 324287 41332 324327 41334
rect 325490 41332 325531 41334
rect 325671 41332 325701 41334
rect 325881 41332 325915 41334
rect 326055 41332 326092 41334
rect 327262 41332 327299 41334
rect 327439 41332 327473 41334
rect 327650 41332 327683 41334
rect 327823 41332 327861 41334
rect 329032 41332 329067 41334
rect 329207 41332 329243 41334
rect 329419 41332 329451 41334
rect 329591 41332 329630 41334
rect 330798 41332 330835 41334
rect 330975 41332 331009 41334
rect 331185 41332 331219 41334
rect 331359 41332 331396 41334
rect 332571 41332 332603 41334
rect 332743 41332 332782 41334
rect 362344 41332 362379 41334
rect 362519 41332 362555 41334
rect 363730 41332 363763 41334
rect 363903 41332 363941 41334
rect 364116 41332 364147 41334
rect 364287 41332 364327 41334
rect 365490 41332 365531 41334
rect 365671 41332 365701 41334
rect 365881 41332 365915 41334
rect 366055 41332 366092 41334
rect 367262 41332 367299 41334
rect 367439 41332 367473 41334
rect 367650 41332 367683 41334
rect 367823 41332 367861 41334
rect 369032 41332 369067 41334
rect 369207 41332 369243 41334
rect 369419 41332 369451 41334
rect 369591 41332 369630 41334
rect 370798 41332 370835 41334
rect 370975 41332 371009 41334
rect 371185 41332 371219 41334
rect 371359 41332 371396 41334
rect 372571 41332 372603 41334
rect 372743 41332 372782 41334
rect 402344 41332 402379 41334
rect 402519 41332 402555 41334
rect 403730 41332 403763 41334
rect 403903 41332 403941 41334
rect 404116 41332 404147 41334
rect 404287 41332 404327 41334
rect 405490 41332 405531 41334
rect 405671 41332 405701 41334
rect 405881 41332 405915 41334
rect 406055 41332 406092 41334
rect 407262 41332 407299 41334
rect 407439 41332 407473 41334
rect 407650 41332 407683 41334
rect 407823 41332 407861 41334
rect 409032 41332 409067 41334
rect 409207 41332 409243 41334
rect 409419 41332 409451 41334
rect 409591 41332 409630 41334
rect 410798 41332 410835 41334
rect 410975 41332 411009 41334
rect 411185 41332 411219 41334
rect 411359 41332 411396 41334
rect 412571 41332 412603 41334
rect 412743 41332 412782 41334
rect 422344 41332 422379 41334
rect 422519 41332 422555 41334
rect 423730 41332 423763 41334
rect 423903 41332 423941 41334
rect 424116 41332 424147 41334
rect 424287 41332 424327 41334
rect 425490 41332 425531 41334
rect 425671 41332 425701 41334
rect 425881 41332 425915 41334
rect 426055 41332 426092 41334
rect 427262 41332 427299 41334
rect 427439 41332 427473 41334
rect 427650 41332 427683 41334
rect 427823 41332 427861 41334
rect 429032 41332 429067 41334
rect 429207 41332 429243 41334
rect 429419 41332 429451 41334
rect 429591 41332 429630 41334
rect 430798 41332 430835 41334
rect 430975 41332 431009 41334
rect 431185 41332 431219 41334
rect 431359 41332 431396 41334
rect 432571 41332 432603 41334
rect 432743 41332 432782 41334
rect 462344 41332 462379 41334
rect 462519 41332 462555 41334
rect 463730 41332 463763 41334
rect 463903 41332 463941 41334
rect 464116 41332 464147 41334
rect 464287 41332 464327 41334
rect 465490 41332 465531 41334
rect 465671 41332 465701 41334
rect 465881 41332 465915 41334
rect 466055 41332 466092 41334
rect 467262 41332 467299 41334
rect 467439 41332 467473 41334
rect 467650 41332 467683 41334
rect 467823 41332 467861 41334
rect 469032 41332 469067 41334
rect 469207 41332 469243 41334
rect 469419 41332 469451 41334
rect 469591 41332 469630 41334
rect 470798 41332 470835 41334
rect 470975 41332 471009 41334
rect 471185 41332 471219 41334
rect 471359 41332 471396 41334
rect 472571 41332 472603 41334
rect 472743 41332 472782 41334
rect 202323 41242 202379 41244
rect 202519 41242 202645 41244
rect 203640 41242 203763 41244
rect 203903 41242 203959 41244
rect 204091 41242 204147 41244
rect 204287 41242 204417 41244
rect 205400 41242 205531 41244
rect 205671 41242 205727 41244
rect 205859 41242 205915 41244
rect 206055 41242 206182 41244
rect 207172 41242 207299 41244
rect 207439 41242 207495 41244
rect 207627 41242 207683 41244
rect 207823 41242 207951 41244
rect 208942 41242 209067 41244
rect 209207 41242 209263 41244
rect 209395 41242 209451 41244
rect 209591 41242 209720 41244
rect 210708 41242 210835 41244
rect 210975 41242 211031 41244
rect 211163 41242 211219 41244
rect 211359 41242 211486 41244
rect 212481 41242 212603 41244
rect 212743 41242 212799 41244
rect 242323 41242 242379 41244
rect 242519 41242 242645 41244
rect 243640 41242 243763 41244
rect 243903 41242 243959 41244
rect 244091 41242 244147 41244
rect 244287 41242 244417 41244
rect 245400 41242 245531 41244
rect 245671 41242 245727 41244
rect 245859 41242 245915 41244
rect 246055 41242 246182 41244
rect 247172 41242 247299 41244
rect 247439 41242 247495 41244
rect 247627 41242 247683 41244
rect 247823 41242 247951 41244
rect 248942 41242 249067 41244
rect 249207 41242 249263 41244
rect 249395 41242 249451 41244
rect 249591 41242 249720 41244
rect 250708 41242 250835 41244
rect 250975 41242 251031 41244
rect 251163 41242 251219 41244
rect 251359 41242 251486 41244
rect 252481 41242 252603 41244
rect 252743 41242 252799 41244
rect 262323 41242 262379 41244
rect 262519 41242 262645 41244
rect 263640 41242 263763 41244
rect 263903 41242 263959 41244
rect 264091 41242 264147 41244
rect 264287 41242 264417 41244
rect 265400 41242 265531 41244
rect 265671 41242 265727 41244
rect 265859 41242 265915 41244
rect 266055 41242 266182 41244
rect 267172 41242 267299 41244
rect 267439 41242 267495 41244
rect 267627 41242 267683 41244
rect 267823 41242 267951 41244
rect 268942 41242 269067 41244
rect 269207 41242 269263 41244
rect 269395 41242 269451 41244
rect 269591 41242 269720 41244
rect 270708 41242 270835 41244
rect 270975 41242 271031 41244
rect 271163 41242 271219 41244
rect 271359 41242 271486 41244
rect 272481 41242 272603 41244
rect 272743 41242 272799 41244
rect 302323 41242 302379 41244
rect 302519 41242 302645 41244
rect 303640 41242 303763 41244
rect 303903 41242 303959 41244
rect 304091 41242 304147 41244
rect 304287 41242 304417 41244
rect 305400 41242 305531 41244
rect 305671 41242 305727 41244
rect 305859 41242 305915 41244
rect 306055 41242 306182 41244
rect 307172 41242 307299 41244
rect 307439 41242 307495 41244
rect 307627 41242 307683 41244
rect 307823 41242 307951 41244
rect 308942 41242 309067 41244
rect 309207 41242 309263 41244
rect 309395 41242 309451 41244
rect 309591 41242 309720 41244
rect 310708 41242 310835 41244
rect 310975 41242 311031 41244
rect 311163 41242 311219 41244
rect 311359 41242 311486 41244
rect 312481 41242 312603 41244
rect 312743 41242 312799 41244
rect 322323 41242 322379 41244
rect 322519 41242 322645 41244
rect 323640 41242 323763 41244
rect 323903 41242 323959 41244
rect 324091 41242 324147 41244
rect 324287 41242 324417 41244
rect 325400 41242 325531 41244
rect 325671 41242 325727 41244
rect 325859 41242 325915 41244
rect 326055 41242 326182 41244
rect 327172 41242 327299 41244
rect 327439 41242 327495 41244
rect 327627 41242 327683 41244
rect 327823 41242 327951 41244
rect 328942 41242 329067 41244
rect 329207 41242 329263 41244
rect 329395 41242 329451 41244
rect 329591 41242 329720 41244
rect 330708 41242 330835 41244
rect 330975 41242 331031 41244
rect 331163 41242 331219 41244
rect 331359 41242 331486 41244
rect 332481 41242 332603 41244
rect 332743 41242 332799 41244
rect 362323 41242 362379 41244
rect 362519 41242 362645 41244
rect 363640 41242 363763 41244
rect 363903 41242 363959 41244
rect 364091 41242 364147 41244
rect 364287 41242 364417 41244
rect 365400 41242 365531 41244
rect 365671 41242 365727 41244
rect 365859 41242 365915 41244
rect 366055 41242 366182 41244
rect 367172 41242 367299 41244
rect 367439 41242 367495 41244
rect 367627 41242 367683 41244
rect 367823 41242 367951 41244
rect 368942 41242 369067 41244
rect 369207 41242 369263 41244
rect 369395 41242 369451 41244
rect 369591 41242 369720 41244
rect 370708 41242 370835 41244
rect 370975 41242 371031 41244
rect 371163 41242 371219 41244
rect 371359 41242 371486 41244
rect 372481 41242 372603 41244
rect 372743 41242 372799 41244
rect 402323 41242 402379 41244
rect 402519 41242 402645 41244
rect 403640 41242 403763 41244
rect 403903 41242 403959 41244
rect 404091 41242 404147 41244
rect 404287 41242 404417 41244
rect 405400 41242 405531 41244
rect 405671 41242 405727 41244
rect 405859 41242 405915 41244
rect 406055 41242 406182 41244
rect 407172 41242 407299 41244
rect 407439 41242 407495 41244
rect 407627 41242 407683 41244
rect 407823 41242 407951 41244
rect 408942 41242 409067 41244
rect 409207 41242 409263 41244
rect 409395 41242 409451 41244
rect 409591 41242 409720 41244
rect 410708 41242 410835 41244
rect 410975 41242 411031 41244
rect 411163 41242 411219 41244
rect 411359 41242 411486 41244
rect 412481 41242 412603 41244
rect 412743 41242 412799 41244
rect 422323 41242 422379 41244
rect 422519 41242 422645 41244
rect 423640 41242 423763 41244
rect 423903 41242 423959 41244
rect 424091 41242 424147 41244
rect 424287 41242 424417 41244
rect 425400 41242 425531 41244
rect 425671 41242 425727 41244
rect 425859 41242 425915 41244
rect 426055 41242 426182 41244
rect 427172 41242 427299 41244
rect 427439 41242 427495 41244
rect 427627 41242 427683 41244
rect 427823 41242 427951 41244
rect 428942 41242 429067 41244
rect 429207 41242 429263 41244
rect 429395 41242 429451 41244
rect 429591 41242 429720 41244
rect 430708 41242 430835 41244
rect 430975 41242 431031 41244
rect 431163 41242 431219 41244
rect 431359 41242 431486 41244
rect 432481 41242 432603 41244
rect 432743 41242 432799 41244
rect 462323 41242 462379 41244
rect 462519 41242 462645 41244
rect 463640 41242 463763 41244
rect 463903 41242 463959 41244
rect 464091 41242 464147 41244
rect 464287 41242 464417 41244
rect 465400 41242 465531 41244
rect 465671 41242 465727 41244
rect 465859 41242 465915 41244
rect 466055 41242 466182 41244
rect 467172 41242 467299 41244
rect 467439 41242 467495 41244
rect 467627 41242 467683 41244
rect 467823 41242 467951 41244
rect 468942 41242 469067 41244
rect 469207 41242 469263 41244
rect 469395 41242 469451 41244
rect 469591 41242 469720 41244
rect 470708 41242 470835 41244
rect 470975 41242 471031 41244
rect 471163 41242 471219 41244
rect 471359 41242 471486 41244
rect 472481 41242 472603 41244
rect 472743 41242 472799 41244
rect 202323 33244 202379 33246
rect 202519 33244 202645 33246
rect 203640 33244 203763 33246
rect 203903 33244 203959 33246
rect 204091 33244 204147 33246
rect 204287 33244 204417 33246
rect 205400 33244 205531 33246
rect 205671 33244 205727 33246
rect 205859 33244 205915 33246
rect 206055 33244 206182 33246
rect 207172 33244 207299 33246
rect 207439 33244 207495 33246
rect 207627 33244 207683 33246
rect 207823 33244 207951 33246
rect 208942 33244 209067 33246
rect 209207 33244 209263 33246
rect 209395 33244 209451 33246
rect 209591 33244 209720 33246
rect 210708 33244 210835 33246
rect 210975 33244 211031 33246
rect 211163 33244 211219 33246
rect 211359 33244 211486 33246
rect 212481 33244 212603 33246
rect 212743 33244 212799 33246
rect 242323 33244 242379 33246
rect 242519 33244 242645 33246
rect 243640 33244 243763 33246
rect 243903 33244 243959 33246
rect 244091 33244 244147 33246
rect 244287 33244 244417 33246
rect 245400 33244 245531 33246
rect 245671 33244 245727 33246
rect 245859 33244 245915 33246
rect 246055 33244 246182 33246
rect 247172 33244 247299 33246
rect 247439 33244 247495 33246
rect 247627 33244 247683 33246
rect 247823 33244 247951 33246
rect 248942 33244 249067 33246
rect 249207 33244 249263 33246
rect 249395 33244 249451 33246
rect 249591 33244 249720 33246
rect 250708 33244 250835 33246
rect 250975 33244 251031 33246
rect 251163 33244 251219 33246
rect 251359 33244 251486 33246
rect 252481 33244 252603 33246
rect 252743 33244 252799 33246
rect 262323 33244 262379 33246
rect 262519 33244 262645 33246
rect 263640 33244 263763 33246
rect 263903 33244 263959 33246
rect 264091 33244 264147 33246
rect 264287 33244 264417 33246
rect 265400 33244 265531 33246
rect 265671 33244 265727 33246
rect 265859 33244 265915 33246
rect 266055 33244 266182 33246
rect 267172 33244 267299 33246
rect 267439 33244 267495 33246
rect 267627 33244 267683 33246
rect 267823 33244 267951 33246
rect 268942 33244 269067 33246
rect 269207 33244 269263 33246
rect 269395 33244 269451 33246
rect 269591 33244 269720 33246
rect 270708 33244 270835 33246
rect 270975 33244 271031 33246
rect 271163 33244 271219 33246
rect 271359 33244 271486 33246
rect 272481 33244 272603 33246
rect 272743 33244 272799 33246
rect 302323 33244 302379 33246
rect 302519 33244 302645 33246
rect 303640 33244 303763 33246
rect 303903 33244 303959 33246
rect 304091 33244 304147 33246
rect 304287 33244 304417 33246
rect 305400 33244 305531 33246
rect 305671 33244 305727 33246
rect 305859 33244 305915 33246
rect 306055 33244 306182 33246
rect 307172 33244 307299 33246
rect 307439 33244 307495 33246
rect 307627 33244 307683 33246
rect 307823 33244 307951 33246
rect 308942 33244 309067 33246
rect 309207 33244 309263 33246
rect 309395 33244 309451 33246
rect 309591 33244 309720 33246
rect 310708 33244 310835 33246
rect 310975 33244 311031 33246
rect 311163 33244 311219 33246
rect 311359 33244 311486 33246
rect 312481 33244 312603 33246
rect 312743 33244 312799 33246
rect 322323 33244 322379 33246
rect 322519 33244 322645 33246
rect 323640 33244 323763 33246
rect 323903 33244 323959 33246
rect 324091 33244 324147 33246
rect 324287 33244 324417 33246
rect 325400 33244 325531 33246
rect 325671 33244 325727 33246
rect 325859 33244 325915 33246
rect 326055 33244 326182 33246
rect 327172 33244 327299 33246
rect 327439 33244 327495 33246
rect 327627 33244 327683 33246
rect 327823 33244 327951 33246
rect 328942 33244 329067 33246
rect 329207 33244 329263 33246
rect 329395 33244 329451 33246
rect 329591 33244 329720 33246
rect 330708 33244 330835 33246
rect 330975 33244 331031 33246
rect 331163 33244 331219 33246
rect 331359 33244 331486 33246
rect 332481 33244 332603 33246
rect 332743 33244 332799 33246
rect 362323 33244 362379 33246
rect 362519 33244 362645 33246
rect 363640 33244 363763 33246
rect 363903 33244 363959 33246
rect 364091 33244 364147 33246
rect 364287 33244 364417 33246
rect 365400 33244 365531 33246
rect 365671 33244 365727 33246
rect 365859 33244 365915 33246
rect 366055 33244 366182 33246
rect 367172 33244 367299 33246
rect 367439 33244 367495 33246
rect 367627 33244 367683 33246
rect 367823 33244 367951 33246
rect 368942 33244 369067 33246
rect 369207 33244 369263 33246
rect 369395 33244 369451 33246
rect 369591 33244 369720 33246
rect 370708 33244 370835 33246
rect 370975 33244 371031 33246
rect 371163 33244 371219 33246
rect 371359 33244 371486 33246
rect 372481 33244 372603 33246
rect 372743 33244 372799 33246
rect 402323 33244 402379 33246
rect 402519 33244 402645 33246
rect 403640 33244 403763 33246
rect 403903 33244 403959 33246
rect 404091 33244 404147 33246
rect 404287 33244 404417 33246
rect 405400 33244 405531 33246
rect 405671 33244 405727 33246
rect 405859 33244 405915 33246
rect 406055 33244 406182 33246
rect 407172 33244 407299 33246
rect 407439 33244 407495 33246
rect 407627 33244 407683 33246
rect 407823 33244 407951 33246
rect 408942 33244 409067 33246
rect 409207 33244 409263 33246
rect 409395 33244 409451 33246
rect 409591 33244 409720 33246
rect 410708 33244 410835 33246
rect 410975 33244 411031 33246
rect 411163 33244 411219 33246
rect 411359 33244 411486 33246
rect 412481 33244 412603 33246
rect 412743 33244 412799 33246
rect 422323 33244 422379 33246
rect 422519 33244 422645 33246
rect 423640 33244 423763 33246
rect 423903 33244 423959 33246
rect 424091 33244 424147 33246
rect 424287 33244 424417 33246
rect 425400 33244 425531 33246
rect 425671 33244 425727 33246
rect 425859 33244 425915 33246
rect 426055 33244 426182 33246
rect 427172 33244 427299 33246
rect 427439 33244 427495 33246
rect 427627 33244 427683 33246
rect 427823 33244 427951 33246
rect 428942 33244 429067 33246
rect 429207 33244 429263 33246
rect 429395 33244 429451 33246
rect 429591 33244 429720 33246
rect 430708 33244 430835 33246
rect 430975 33244 431031 33246
rect 431163 33244 431219 33246
rect 431359 33244 431486 33246
rect 432481 33244 432603 33246
rect 432743 33244 432799 33246
rect 462323 33244 462379 33246
rect 462519 33244 462645 33246
rect 463640 33244 463763 33246
rect 463903 33244 463959 33246
rect 464091 33244 464147 33246
rect 464287 33244 464417 33246
rect 465400 33244 465531 33246
rect 465671 33244 465727 33246
rect 465859 33244 465915 33246
rect 466055 33244 466182 33246
rect 467172 33244 467299 33246
rect 467439 33244 467495 33246
rect 467627 33244 467683 33246
rect 467823 33244 467951 33246
rect 468942 33244 469067 33246
rect 469207 33244 469263 33246
rect 469395 33244 469451 33246
rect 469591 33244 469720 33246
rect 470708 33244 470835 33246
rect 470975 33244 471031 33246
rect 471163 33244 471219 33246
rect 471359 33244 471486 33246
rect 472481 33244 472603 33246
rect 472743 33244 472799 33246
rect 202344 33154 202379 33156
rect 202519 33154 202555 33156
rect 203730 33154 203763 33156
rect 203903 33154 203941 33156
rect 204116 33154 204147 33156
rect 204287 33154 204327 33156
rect 205490 33154 205531 33156
rect 205671 33154 205701 33156
rect 205881 33154 205915 33156
rect 206055 33154 206092 33156
rect 207262 33154 207299 33156
rect 207439 33154 207473 33156
rect 207650 33154 207683 33156
rect 207823 33154 207861 33156
rect 209032 33154 209067 33156
rect 209207 33154 209243 33156
rect 209419 33154 209451 33156
rect 209591 33154 209630 33156
rect 210798 33154 210835 33156
rect 210975 33154 211009 33156
rect 211185 33154 211219 33156
rect 211359 33154 211396 33156
rect 212571 33154 212603 33156
rect 212743 33154 212782 33156
rect 242344 33154 242379 33156
rect 242519 33154 242555 33156
rect 243730 33154 243763 33156
rect 243903 33154 243941 33156
rect 244116 33154 244147 33156
rect 244287 33154 244327 33156
rect 245490 33154 245531 33156
rect 245671 33154 245701 33156
rect 245881 33154 245915 33156
rect 246055 33154 246092 33156
rect 247262 33154 247299 33156
rect 247439 33154 247473 33156
rect 247650 33154 247683 33156
rect 247823 33154 247861 33156
rect 249032 33154 249067 33156
rect 249207 33154 249243 33156
rect 249419 33154 249451 33156
rect 249591 33154 249630 33156
rect 250798 33154 250835 33156
rect 250975 33154 251009 33156
rect 251185 33154 251219 33156
rect 251359 33154 251396 33156
rect 252571 33154 252603 33156
rect 252743 33154 252782 33156
rect 262344 33154 262379 33156
rect 262519 33154 262555 33156
rect 263730 33154 263763 33156
rect 263903 33154 263941 33156
rect 264116 33154 264147 33156
rect 264287 33154 264327 33156
rect 265490 33154 265531 33156
rect 265671 33154 265701 33156
rect 265881 33154 265915 33156
rect 266055 33154 266092 33156
rect 267262 33154 267299 33156
rect 267439 33154 267473 33156
rect 267650 33154 267683 33156
rect 267823 33154 267861 33156
rect 269032 33154 269067 33156
rect 269207 33154 269243 33156
rect 269419 33154 269451 33156
rect 269591 33154 269630 33156
rect 270798 33154 270835 33156
rect 270975 33154 271009 33156
rect 271185 33154 271219 33156
rect 271359 33154 271396 33156
rect 272571 33154 272603 33156
rect 272743 33154 272782 33156
rect 302344 33154 302379 33156
rect 302519 33154 302555 33156
rect 303730 33154 303763 33156
rect 303903 33154 303941 33156
rect 304116 33154 304147 33156
rect 304287 33154 304327 33156
rect 305490 33154 305531 33156
rect 305671 33154 305701 33156
rect 305881 33154 305915 33156
rect 306055 33154 306092 33156
rect 307262 33154 307299 33156
rect 307439 33154 307473 33156
rect 307650 33154 307683 33156
rect 307823 33154 307861 33156
rect 309032 33154 309067 33156
rect 309207 33154 309243 33156
rect 309419 33154 309451 33156
rect 309591 33154 309630 33156
rect 310798 33154 310835 33156
rect 310975 33154 311009 33156
rect 311185 33154 311219 33156
rect 311359 33154 311396 33156
rect 312571 33154 312603 33156
rect 312743 33154 312782 33156
rect 322344 33154 322379 33156
rect 322519 33154 322555 33156
rect 323730 33154 323763 33156
rect 323903 33154 323941 33156
rect 324116 33154 324147 33156
rect 324287 33154 324327 33156
rect 325490 33154 325531 33156
rect 325671 33154 325701 33156
rect 325881 33154 325915 33156
rect 326055 33154 326092 33156
rect 327262 33154 327299 33156
rect 327439 33154 327473 33156
rect 327650 33154 327683 33156
rect 327823 33154 327861 33156
rect 329032 33154 329067 33156
rect 329207 33154 329243 33156
rect 329419 33154 329451 33156
rect 329591 33154 329630 33156
rect 330798 33154 330835 33156
rect 330975 33154 331009 33156
rect 331185 33154 331219 33156
rect 331359 33154 331396 33156
rect 332571 33154 332603 33156
rect 332743 33154 332782 33156
rect 362344 33154 362379 33156
rect 362519 33154 362555 33156
rect 363730 33154 363763 33156
rect 363903 33154 363941 33156
rect 364116 33154 364147 33156
rect 364287 33154 364327 33156
rect 365490 33154 365531 33156
rect 365671 33154 365701 33156
rect 365881 33154 365915 33156
rect 366055 33154 366092 33156
rect 367262 33154 367299 33156
rect 367439 33154 367473 33156
rect 367650 33154 367683 33156
rect 367823 33154 367861 33156
rect 369032 33154 369067 33156
rect 369207 33154 369243 33156
rect 369419 33154 369451 33156
rect 369591 33154 369630 33156
rect 370798 33154 370835 33156
rect 370975 33154 371009 33156
rect 371185 33154 371219 33156
rect 371359 33154 371396 33156
rect 372571 33154 372603 33156
rect 372743 33154 372782 33156
rect 402344 33154 402379 33156
rect 402519 33154 402555 33156
rect 403730 33154 403763 33156
rect 403903 33154 403941 33156
rect 404116 33154 404147 33156
rect 404287 33154 404327 33156
rect 405490 33154 405531 33156
rect 405671 33154 405701 33156
rect 405881 33154 405915 33156
rect 406055 33154 406092 33156
rect 407262 33154 407299 33156
rect 407439 33154 407473 33156
rect 407650 33154 407683 33156
rect 407823 33154 407861 33156
rect 409032 33154 409067 33156
rect 409207 33154 409243 33156
rect 409419 33154 409451 33156
rect 409591 33154 409630 33156
rect 410798 33154 410835 33156
rect 410975 33154 411009 33156
rect 411185 33154 411219 33156
rect 411359 33154 411396 33156
rect 412571 33154 412603 33156
rect 412743 33154 412782 33156
rect 422344 33154 422379 33156
rect 422519 33154 422555 33156
rect 423730 33154 423763 33156
rect 423903 33154 423941 33156
rect 424116 33154 424147 33156
rect 424287 33154 424327 33156
rect 425490 33154 425531 33156
rect 425671 33154 425701 33156
rect 425881 33154 425915 33156
rect 426055 33154 426092 33156
rect 427262 33154 427299 33156
rect 427439 33154 427473 33156
rect 427650 33154 427683 33156
rect 427823 33154 427861 33156
rect 429032 33154 429067 33156
rect 429207 33154 429243 33156
rect 429419 33154 429451 33156
rect 429591 33154 429630 33156
rect 430798 33154 430835 33156
rect 430975 33154 431009 33156
rect 431185 33154 431219 33156
rect 431359 33154 431396 33156
rect 432571 33154 432603 33156
rect 432743 33154 432782 33156
rect 462344 33154 462379 33156
rect 462519 33154 462555 33156
rect 463730 33154 463763 33156
rect 463903 33154 463941 33156
rect 464116 33154 464147 33156
rect 464287 33154 464327 33156
rect 465490 33154 465531 33156
rect 465671 33154 465701 33156
rect 465881 33154 465915 33156
rect 466055 33154 466092 33156
rect 467262 33154 467299 33156
rect 467439 33154 467473 33156
rect 467650 33154 467683 33156
rect 467823 33154 467861 33156
rect 469032 33154 469067 33156
rect 469207 33154 469243 33156
rect 469419 33154 469451 33156
rect 469591 33154 469630 33156
rect 470798 33154 470835 33156
rect 470975 33154 471009 33156
rect 471185 33154 471219 33156
rect 471359 33154 471396 33156
rect 472571 33154 472603 33156
rect 472743 33154 472782 33156
rect 201938 28790 202120 28873
rect 213002 28790 213183 28873
rect 221938 28790 222092 28873
rect 233028 28790 233183 28873
rect 241938 28790 242120 28873
rect 253002 28790 253183 28873
rect 261938 28790 262120 28873
rect 273002 28790 273183 28873
rect 301938 28790 302120 28873
rect 313002 28790 313183 28873
rect 321938 28790 322120 28873
rect 333002 28790 333183 28873
rect 341938 28790 342092 28873
rect 353028 28790 353183 28873
rect 361938 28790 362120 28873
rect 373002 28790 373183 28873
rect 401938 28790 402120 28873
rect 413002 28790 413183 28873
rect 421938 28790 422120 28873
rect 433002 28790 433183 28873
rect 441938 28790 442092 28873
rect 453028 28790 453183 28873
rect 461938 28790 462120 28873
rect 473002 28790 473183 28873
rect 501938 28790 502092 28873
rect 513028 28790 513183 28873
rect 202024 27973 202025 28790
rect 202034 27973 202120 28790
rect 202024 27972 202120 27973
rect 213088 27972 213183 28790
rect 222024 27973 222025 28790
rect 222034 27973 222092 28790
rect 222024 27972 222092 27973
rect 233088 27972 233183 28790
rect 242024 27973 242025 28790
rect 242034 27973 242120 28790
rect 242024 27972 242120 27973
rect 253088 27972 253183 28790
rect 262024 27973 262025 28790
rect 262034 27973 262120 28790
rect 262024 27972 262120 27973
rect 273088 27972 273183 28790
rect 302024 27973 302025 28790
rect 302034 27973 302120 28790
rect 302024 27972 302120 27973
rect 313088 27972 313183 28790
rect 322024 27973 322025 28790
rect 322034 27973 322120 28790
rect 322024 27972 322120 27973
rect 333088 27972 333183 28790
rect 342024 27973 342025 28790
rect 342034 27973 342092 28790
rect 342024 27972 342092 27973
rect 353088 27972 353183 28790
rect 362024 27973 362025 28790
rect 362034 27973 362120 28790
rect 362024 27972 362120 27973
rect 373088 27972 373183 28790
rect 402024 27973 402025 28790
rect 402034 27973 402120 28790
rect 402024 27972 402120 27973
rect 413088 27972 413183 28790
rect 422024 27973 422025 28790
rect 422034 27973 422120 28790
rect 422024 27972 422120 27973
rect 433088 27972 433183 28790
rect 442024 27973 442025 28790
rect 442034 27973 442092 28790
rect 442024 27972 442092 27973
rect 453088 27972 453183 28790
rect 462024 27973 462025 28790
rect 462034 27973 462120 28790
rect 462024 27972 462120 27973
rect 473088 27972 473183 28790
rect 502024 27973 502025 28790
rect 502034 27973 502092 28790
rect 502024 27972 502092 27973
rect 513088 27972 513183 28790
rect 201938 18377 202024 18380
rect 213097 18377 213183 18380
rect 201938 18294 202066 18377
rect 213056 18294 213183 18377
rect 221938 18377 222024 18380
rect 233097 18377 233183 18380
rect 221938 18294 222066 18377
rect 233056 18294 233183 18377
rect 241938 18377 242024 18380
rect 253097 18377 253183 18380
rect 241938 18294 242066 18377
rect 253056 18294 253183 18377
rect 261938 18377 262024 18380
rect 273097 18377 273183 18380
rect 261938 18294 262066 18377
rect 273056 18294 273183 18377
rect 301938 18377 302024 18380
rect 313097 18377 313183 18380
rect 301938 18294 302066 18377
rect 313056 18294 313183 18377
rect 321938 18377 322024 18380
rect 333097 18377 333183 18380
rect 321938 18294 322066 18377
rect 333056 18294 333183 18377
rect 341938 18377 342024 18380
rect 353097 18377 353183 18380
rect 341938 18294 342066 18377
rect 353056 18294 353183 18377
rect 361938 18377 362024 18380
rect 373097 18377 373183 18380
rect 361938 18294 362066 18377
rect 373056 18294 373183 18377
rect 401938 18377 402024 18380
rect 413097 18377 413183 18380
rect 401938 18294 402066 18377
rect 413056 18294 413183 18377
rect 421938 18377 422024 18380
rect 433097 18377 433183 18380
rect 421938 18294 422066 18377
rect 433056 18294 433183 18377
rect 441938 18377 442024 18380
rect 453097 18377 453183 18380
rect 441938 18294 442066 18377
rect 453056 18294 453183 18377
rect 461938 18377 462024 18380
rect 473097 18377 473183 18380
rect 461938 18294 462066 18377
rect 473056 18294 473183 18377
rect 501938 18377 502024 18380
rect 513097 18377 513183 18380
rect 501938 18294 502066 18377
rect 513056 18294 513183 18377
rect 202024 17893 202025 18294
rect 202066 17893 213056 18294
rect 213097 17893 213183 18294
rect 202024 17892 213183 17893
rect 222024 17893 222025 18294
rect 222066 17893 224000 18294
rect 222024 17892 224000 17893
rect 231028 17893 233056 18294
rect 233097 17893 233183 18294
rect 231028 17892 233183 17893
rect 242024 17893 242025 18294
rect 242066 17893 253056 18294
rect 253097 17893 253183 18294
rect 242024 17892 253183 17893
rect 262024 17893 262025 18294
rect 262066 17893 273056 18294
rect 273097 17893 273183 18294
rect 262024 17892 273183 17893
rect 302024 17893 302025 18294
rect 302066 17893 313056 18294
rect 313097 17893 313183 18294
rect 302024 17892 313183 17893
rect 322024 17893 322025 18294
rect 322066 17893 333056 18294
rect 333097 17893 333183 18294
rect 322024 17892 333183 17893
rect 342024 17893 342025 18294
rect 342066 17893 344092 18294
rect 342024 17892 344092 17893
rect 351028 17893 353056 18294
rect 353097 17893 353183 18294
rect 351028 17892 353183 17893
rect 362024 17893 362025 18294
rect 362066 17893 373056 18294
rect 373097 17893 373183 18294
rect 362024 17892 373183 17893
rect 402024 17893 402025 18294
rect 402066 17893 413056 18294
rect 413097 17893 413183 18294
rect 402024 17892 413183 17893
rect 422024 17893 422025 18294
rect 422066 17893 433056 18294
rect 433097 17893 433183 18294
rect 422024 17892 433183 17893
rect 442024 17893 442025 18294
rect 442066 17893 444092 18294
rect 442024 17892 444092 17893
rect 451028 17893 453056 18294
rect 453097 17893 453183 18294
rect 451028 17892 453183 17893
rect 462024 17893 462025 18294
rect 462066 17893 473056 18294
rect 473097 17893 473183 18294
rect 462024 17892 473183 17893
rect 502024 17893 502025 18294
rect 502066 17893 504092 18294
rect 502024 17892 504092 17893
rect 511028 17893 513056 18294
rect 513097 17893 513183 18294
rect 511028 17892 513183 17893
rect 520063 17415 520116 73873
rect 520007 17351 520060 17407
rect 520063 17157 520116 17351
<< metal1 >>
rect 74569 440932 148250 441191
rect 74569 440906 75058 440932
rect 74569 440888 74846 440906
rect 74569 440812 74676 440888
rect 74752 440830 74846 440888
rect 74922 440856 75058 440906
rect 75134 440856 148250 440932
rect 74922 440830 148250 440856
rect 74752 440812 148250 440830
rect 74569 440782 148250 440812
rect 74569 440706 75037 440782
rect 75113 440706 148250 440782
rect 74569 440632 148250 440706
rect 74569 440625 75036 440632
rect 74569 440619 74825 440625
rect 74569 440543 74655 440619
rect 74731 440549 74825 440619
rect 74901 440556 75036 440625
rect 75112 440556 148250 440632
rect 74901 440549 148250 440556
rect 74731 440543 148250 440549
rect 74569 440510 148250 440543
rect 74574 440509 148250 440510
rect 74339 420662 74977 420665
rect 74339 420581 146967 420662
rect 74339 420555 74830 420581
rect 74339 420537 74618 420555
rect 74339 420461 74448 420537
rect 74524 420479 74618 420537
rect 74694 420505 74830 420555
rect 74906 420505 146967 420581
rect 74694 420479 146967 420505
rect 74524 420461 146967 420479
rect 74339 420431 146967 420461
rect 74339 420355 74809 420431
rect 74885 420355 146967 420431
rect 74339 420281 146967 420355
rect 74339 420274 74808 420281
rect 74339 420268 74597 420274
rect 74339 420192 74427 420268
rect 74503 420198 74597 420268
rect 74673 420205 74808 420274
rect 74884 420205 146967 420281
rect 74673 420198 146967 420205
rect 74503 420192 146967 420198
rect 74339 420136 146967 420192
rect 74306 400767 75158 400768
rect 74306 400684 150157 400767
rect 74306 400658 74797 400684
rect 74306 400640 74585 400658
rect 74306 400564 74415 400640
rect 74491 400582 74585 400640
rect 74661 400608 74797 400658
rect 74873 400608 150157 400684
rect 74661 400582 150157 400608
rect 74491 400564 150157 400582
rect 74306 400534 150157 400564
rect 74306 400458 74776 400534
rect 74852 400458 150157 400534
rect 74306 400384 150157 400458
rect 74306 400377 74775 400384
rect 74306 400371 74564 400377
rect 74306 400295 74394 400371
rect 74470 400301 74564 400371
rect 74640 400308 74775 400377
rect 74851 400308 150157 400384
rect 74640 400301 150157 400308
rect 74470 400295 150157 400301
rect 74306 400239 150157 400295
rect 74131 380767 74983 380768
rect 149400 380767 149928 382857
rect 74131 380684 149928 380767
rect 74131 380658 74622 380684
rect 74131 380640 74410 380658
rect 74131 380564 74240 380640
rect 74316 380582 74410 380640
rect 74486 380608 74622 380658
rect 74698 380608 149928 380684
rect 74486 380582 149928 380608
rect 74316 380564 149928 380582
rect 74131 380534 149928 380564
rect 74131 380458 74601 380534
rect 74677 380458 149928 380534
rect 74131 380384 149928 380458
rect 74131 380377 74600 380384
rect 74131 380371 74389 380377
rect 74131 380295 74219 380371
rect 74295 380301 74389 380371
rect 74465 380308 74600 380377
rect 74676 380308 149928 380384
rect 74465 380301 149928 380308
rect 74295 380295 149928 380301
rect 74131 380239 149928 380295
rect 74194 340743 75046 340744
rect 74194 340660 143989 340743
rect 74194 340634 74685 340660
rect 74194 340616 74473 340634
rect 74194 340540 74303 340616
rect 74379 340558 74473 340616
rect 74549 340584 74685 340634
rect 74761 340584 143989 340660
rect 74549 340558 143989 340584
rect 74379 340540 143989 340558
rect 74194 340510 143989 340540
rect 74194 340434 74664 340510
rect 74740 340434 143989 340510
rect 74194 340360 143989 340434
rect 74194 340353 74663 340360
rect 74194 340347 74452 340353
rect 74194 340271 74282 340347
rect 74358 340277 74452 340347
rect 74528 340284 74663 340353
rect 74739 340284 143989 340360
rect 74528 340277 143989 340284
rect 74358 340271 143989 340277
rect 74194 340215 143989 340271
rect 74144 320736 74818 320888
rect 74144 320735 75032 320736
rect 143492 320735 144020 322602
rect 74144 320652 144020 320735
rect 74144 320626 74671 320652
rect 74144 320608 74459 320626
rect 74144 320532 74289 320608
rect 74365 320550 74459 320608
rect 74535 320576 74671 320626
rect 74747 320576 144020 320652
rect 74535 320550 144020 320576
rect 74365 320532 144020 320550
rect 74144 320502 144020 320532
rect 74144 320426 74650 320502
rect 74726 320426 144020 320502
rect 74144 320352 144020 320426
rect 74144 320345 74649 320352
rect 74144 320339 74438 320345
rect 74144 320263 74268 320339
rect 74344 320269 74438 320339
rect 74514 320276 74649 320345
rect 74725 320276 144020 320352
rect 74514 320269 144020 320276
rect 74344 320263 144020 320269
rect 74144 320207 144020 320263
<< via1 >>
rect 74676 440812 74752 440888
rect 74846 440830 74922 440906
rect 75058 440856 75134 440932
rect 75037 440706 75113 440782
rect 74655 440543 74731 440619
rect 74825 440549 74901 440625
rect 75036 440556 75112 440632
rect 74448 420461 74524 420537
rect 74618 420479 74694 420555
rect 74830 420505 74906 420581
rect 74809 420355 74885 420431
rect 74427 420192 74503 420268
rect 74597 420198 74673 420274
rect 74808 420205 74884 420281
rect 74415 400564 74491 400640
rect 74585 400582 74661 400658
rect 74797 400608 74873 400684
rect 74776 400458 74852 400534
rect 74394 400295 74470 400371
rect 74564 400301 74640 400377
rect 74775 400308 74851 400384
rect 74240 380564 74316 380640
rect 74410 380582 74486 380658
rect 74622 380608 74698 380684
rect 74601 380458 74677 380534
rect 74219 380295 74295 380371
rect 74389 380301 74465 380377
rect 74600 380308 74676 380384
rect 74303 340540 74379 340616
rect 74473 340558 74549 340634
rect 74685 340584 74761 340660
rect 74664 340434 74740 340510
rect 74282 340271 74358 340347
rect 74452 340277 74528 340353
rect 74663 340284 74739 340360
rect 74289 320532 74365 320608
rect 74459 320550 74535 320626
rect 74671 320576 74747 320652
rect 74650 320426 74726 320502
rect 74268 320263 74344 320339
rect 74438 320269 74514 320345
rect 74649 320276 74725 320352
<< metal2 >>
rect 90963 467581 97688 468097
rect 90963 467431 91879 467581
rect 92029 467431 92147 467581
rect 92297 467431 92415 467581
rect 92565 467431 92683 467581
rect 92833 467431 92951 467581
rect 93101 467431 93219 467581
rect 93369 467431 93487 467581
rect 93637 467431 93755 467581
rect 93905 467431 94023 467581
rect 94173 467431 94291 467581
rect 94441 467431 97688 467581
rect 90963 467343 97688 467431
rect 90963 467232 91879 467343
rect 72010 467193 91879 467232
rect 92029 467193 92147 467343
rect 92297 467193 92415 467343
rect 92565 467193 92683 467343
rect 92833 467193 92951 467343
rect 93101 467193 93219 467343
rect 93369 467193 93487 467343
rect 93637 467193 93755 467343
rect 93905 467193 94023 467343
rect 94173 467193 94291 467343
rect 94441 467193 97688 467343
rect 72010 467105 97688 467193
rect 72010 466955 91879 467105
rect 92029 466955 92147 467105
rect 92297 466955 92415 467105
rect 92565 466955 92683 467105
rect 92833 466955 92951 467105
rect 93101 466955 93219 467105
rect 93369 466955 93487 467105
rect 93637 466955 93755 467105
rect 93905 466955 94023 467105
rect 94173 466955 94291 467105
rect 94441 466955 97688 467105
rect 72010 466867 97688 466955
rect 72010 466717 91879 466867
rect 92029 466717 92147 466867
rect 92297 466717 92415 466867
rect 92565 466717 92683 466867
rect 92833 466717 92951 466867
rect 93101 466717 93219 466867
rect 93369 466717 93487 466867
rect 93637 466717 93755 466867
rect 93905 466717 94023 466867
rect 94173 466717 94291 466867
rect 94441 466717 97688 466867
rect 72010 466629 97688 466717
rect 72010 466479 91879 466629
rect 92029 466479 92147 466629
rect 92297 466479 92415 466629
rect 92565 466479 92683 466629
rect 92833 466479 92951 466629
rect 93101 466479 93219 466629
rect 93369 466479 93487 466629
rect 93637 466479 93755 466629
rect 93905 466479 94023 466629
rect 94173 466479 94291 466629
rect 94441 466479 97688 466629
rect 72010 466391 97688 466479
rect 72010 466241 91879 466391
rect 92029 466241 92147 466391
rect 92297 466241 92415 466391
rect 92565 466241 92683 466391
rect 92833 466241 92951 466391
rect 93101 466241 93219 466391
rect 93369 466241 93487 466391
rect 93637 466241 93755 466391
rect 93905 466241 94023 466391
rect 94173 466241 94291 466391
rect 94441 466241 97688 466391
rect 72010 466153 97688 466241
rect 72010 466003 91879 466153
rect 92029 466003 92147 466153
rect 92297 466003 92415 466153
rect 92565 466003 92683 466153
rect 92833 466003 92951 466153
rect 93101 466003 93219 466153
rect 93369 466003 93487 466153
rect 93637 466003 93755 466153
rect 93905 466003 94023 466153
rect 94173 466003 94291 466153
rect 94441 466003 97688 466153
rect 72010 465915 97688 466003
rect 72010 465765 91879 465915
rect 92029 465765 92147 465915
rect 92297 465765 92415 465915
rect 92565 465765 92683 465915
rect 92833 465765 92951 465915
rect 93101 465765 93219 465915
rect 93369 465765 93487 465915
rect 93637 465765 93755 465915
rect 93905 465765 94023 465915
rect 94173 465765 94291 465915
rect 94441 465765 97688 465915
rect 72010 465677 97688 465765
rect 72010 465527 91879 465677
rect 92029 465527 92147 465677
rect 92297 465527 92415 465677
rect 92565 465527 92683 465677
rect 92833 465527 92951 465677
rect 93101 465527 93219 465677
rect 93369 465527 93487 465677
rect 93637 465527 93755 465677
rect 93905 465527 94023 465677
rect 94173 465527 94291 465677
rect 94441 465527 97688 465677
rect 72010 465439 97688 465527
rect 72010 465289 91879 465439
rect 92029 465289 92147 465439
rect 92297 465289 92415 465439
rect 92565 465289 92683 465439
rect 92833 465289 92951 465439
rect 93101 465289 93219 465439
rect 93369 465289 93487 465439
rect 93637 465289 93755 465439
rect 93905 465289 94023 465439
rect 94173 465289 94291 465439
rect 94441 465289 97688 465439
rect 72010 465182 97688 465289
rect 90963 464614 97688 465182
rect 121375 458462 126869 459116
rect 121375 457241 123379 458462
rect 124600 457241 126869 458462
rect 121375 456782 126869 457241
rect 121375 456620 125479 456782
rect 121375 455399 123282 456620
rect 124503 455561 125479 456620
rect 126700 455561 126869 456782
rect 124503 455399 126869 455561
rect 82014 454512 83235 454961
rect 74330 454436 83235 454512
rect 74330 454388 74499 454436
rect 73984 454314 74499 454388
rect 73984 454312 74406 454314
rect 79501 454114 79577 454436
rect 82014 454114 83235 454436
rect 79501 454038 83235 454114
rect 73984 453791 74625 453867
rect 73984 453562 74348 453638
rect 74272 453559 74348 453562
rect 74549 453559 74625 453791
rect 77796 453559 77872 453561
rect 74272 453496 77872 453559
rect 73984 453483 77872 453496
rect 73984 453420 74349 453483
rect 74554 452994 74630 453483
rect 73984 452918 74630 452994
rect 77739 453273 77872 453483
rect 79501 453385 79577 454038
rect 82014 453385 83235 454038
rect 79501 453309 83235 453385
rect 77739 453140 77981 453273
rect 78114 453140 78123 453273
rect 77739 452783 77872 453140
rect 73734 452708 77872 452783
rect 73734 452707 77815 452708
rect 79501 442873 79577 453309
rect 74283 442797 79577 442873
rect 82014 447194 83235 453309
rect 121375 454423 126869 455399
rect 121375 453202 123056 454423
rect 124277 453369 126869 454423
rect 124277 453202 125729 453369
rect 121375 452148 125729 453202
rect 126950 452148 126959 453369
rect 121375 452129 126869 452148
rect 121375 450908 122862 452129
rect 124083 450908 126869 452129
rect 121375 449649 126869 450908
rect 121375 449640 126950 449649
rect 121375 449576 125729 449640
rect 121375 448355 122765 449576
rect 123986 448419 125729 449576
rect 126950 448419 126959 449640
rect 123986 448410 126950 448419
rect 123986 448355 126869 448410
rect 121375 447249 126869 448355
rect 121375 447194 122603 447249
rect 82014 446028 122603 447194
rect 123824 447194 126869 447249
rect 123824 446028 125729 447194
rect 82014 445973 125729 446028
rect 126950 445973 126959 447194
rect 74283 441329 74359 442797
rect 74004 441253 74359 441329
rect 74283 441034 74359 441253
rect 73984 440958 74359 441034
rect 74569 440989 75124 440990
rect 74569 440932 75201 440989
rect 74569 440906 75058 440932
rect 74569 440888 74846 440906
rect 73984 440812 74676 440888
rect 74752 440830 74846 440888
rect 74922 440856 75058 440906
rect 75134 440856 75201 440932
rect 74922 440830 75201 440856
rect 74752 440812 75201 440830
rect 74569 440782 75201 440812
rect 74569 440706 75037 440782
rect 75113 440706 75201 440782
rect 74569 440632 75201 440706
rect 74569 440625 75036 440632
rect 74569 440619 74825 440625
rect 74569 440543 74655 440619
rect 74731 440549 74825 440619
rect 74901 440556 75036 440625
rect 75112 440556 75201 440632
rect 74901 440549 75201 440556
rect 74731 440543 75201 440549
rect 74569 440510 75201 440543
rect 82014 434388 83235 445973
rect 121375 445963 126869 445973
rect 73984 434312 83235 434388
rect 74027 433867 75955 433884
rect 73984 433791 75955 433867
rect 74027 433754 75955 433791
rect 74027 433654 74642 433754
rect 74742 433654 74810 433754
rect 74910 433654 74978 433754
rect 75078 433654 75146 433754
rect 75246 433654 75314 433754
rect 75414 433654 75482 433754
rect 75582 433654 75650 433754
rect 75750 433654 75818 433754
rect 75918 433654 75954 433754
rect 74027 433638 75954 433654
rect 73984 433596 75954 433638
rect 73984 433562 74642 433596
rect 74027 433496 74642 433562
rect 74742 433496 74810 433596
rect 74910 433496 74978 433596
rect 75078 433496 75146 433596
rect 75246 433496 75314 433596
rect 75414 433496 75482 433596
rect 75582 433496 75650 433596
rect 75750 433496 75818 433596
rect 75918 433496 75954 433596
rect 73984 433438 75954 433496
rect 73984 433420 74642 433438
rect 74027 433338 74642 433420
rect 74742 433338 74810 433438
rect 74910 433338 74978 433438
rect 75078 433338 75146 433438
rect 75246 433338 75314 433438
rect 75414 433338 75482 433438
rect 75582 433338 75650 433438
rect 75750 433338 75818 433438
rect 75918 433338 75954 433438
rect 74027 433280 75954 433338
rect 74027 433180 74642 433280
rect 74742 433180 74810 433280
rect 74910 433180 74978 433280
rect 75078 433180 75146 433280
rect 75246 433180 75314 433280
rect 75414 433180 75482 433280
rect 75582 433180 75650 433280
rect 75750 433180 75818 433280
rect 75918 433180 75954 433280
rect 74027 433122 75954 433180
rect 74027 433022 74642 433122
rect 74742 433022 74810 433122
rect 74910 433022 74978 433122
rect 75078 433022 75146 433122
rect 75246 433022 75314 433122
rect 75414 433022 75482 433122
rect 75582 433022 75650 433122
rect 75750 433022 75818 433122
rect 75918 433022 75954 433122
rect 74027 432994 75954 433022
rect 73984 432964 75954 432994
rect 73984 432918 74642 432964
rect 74027 432864 74642 432918
rect 74742 432864 74810 432964
rect 74910 432864 74978 432964
rect 75078 432864 75146 432964
rect 75246 432864 75314 432964
rect 75414 432864 75482 432964
rect 75582 432864 75650 432964
rect 75750 432864 75818 432964
rect 75918 432864 75954 432964
rect 74027 432806 75954 432864
rect 74027 432783 74642 432806
rect 73984 432707 74642 432783
rect 74576 432706 74642 432707
rect 74742 432706 74810 432806
rect 74910 432706 74978 432806
rect 75078 432706 75146 432806
rect 75246 432706 75314 432806
rect 75414 432706 75482 432806
rect 75582 432706 75650 432806
rect 75750 432706 75818 432806
rect 75918 432706 75954 432806
rect 74576 432648 75954 432706
rect 74576 432548 74642 432648
rect 74742 432548 74810 432648
rect 74910 432548 74978 432648
rect 75078 432548 75146 432648
rect 75246 432548 75314 432648
rect 75414 432548 75482 432648
rect 75582 432548 75650 432648
rect 75750 432548 75818 432648
rect 75918 432548 75954 432648
rect 74576 432520 75954 432548
rect 74576 432511 75797 432520
rect 82014 421326 83235 434312
rect 73984 421250 83235 421326
rect 74901 421034 83235 421250
rect 73984 420958 83235 421034
rect 74339 420888 74977 420889
rect 73984 420812 74977 420888
rect 74339 420581 74977 420812
rect 74339 420555 74830 420581
rect 74339 420537 74618 420555
rect 74339 420461 74448 420537
rect 74524 420479 74618 420537
rect 74694 420505 74830 420555
rect 74906 420505 74977 420581
rect 74694 420479 74977 420505
rect 74524 420461 74977 420479
rect 74339 420431 74977 420461
rect 74339 420355 74809 420431
rect 74885 420355 74977 420431
rect 74339 420281 74977 420355
rect 74339 420274 74808 420281
rect 74339 420268 74597 420274
rect 74339 420192 74427 420268
rect 74503 420198 74597 420268
rect 74673 420205 74808 420274
rect 74884 420205 74977 420281
rect 74673 420198 74977 420205
rect 74503 420192 74977 420198
rect 74339 420136 74977 420192
rect 82014 414388 83235 420958
rect 73784 414312 83235 414388
rect 74676 413867 76190 413905
rect 74052 413817 76190 413867
rect 74052 413717 74761 413817
rect 74861 413717 74929 413817
rect 75029 413717 75097 413817
rect 75197 413717 75265 413817
rect 75365 413717 75433 413817
rect 75533 413717 75601 413817
rect 75701 413717 75769 413817
rect 75869 413717 75937 413817
rect 76037 413717 76190 413817
rect 74052 413659 76190 413717
rect 74052 413559 74761 413659
rect 74861 413559 74929 413659
rect 75029 413559 75097 413659
rect 75197 413559 75265 413659
rect 75365 413559 75433 413659
rect 75533 413559 75601 413659
rect 75701 413559 75769 413659
rect 75869 413559 75937 413659
rect 76037 413559 76190 413659
rect 74052 413501 76190 413559
rect 74052 413401 74761 413501
rect 74861 413401 74929 413501
rect 75029 413401 75097 413501
rect 75197 413401 75265 413501
rect 75365 413401 75433 413501
rect 75533 413401 75601 413501
rect 75701 413401 75769 413501
rect 75869 413401 75937 413501
rect 76037 413401 76190 413501
rect 74052 413343 76190 413401
rect 74052 413243 74761 413343
rect 74861 413243 74929 413343
rect 75029 413243 75097 413343
rect 75197 413243 75265 413343
rect 75365 413243 75433 413343
rect 75533 413243 75601 413343
rect 75701 413243 75769 413343
rect 75869 413243 75937 413343
rect 76037 413243 76190 413343
rect 74052 413185 76190 413243
rect 74052 413085 74761 413185
rect 74861 413085 74929 413185
rect 75029 413085 75097 413185
rect 75197 413085 75265 413185
rect 75365 413085 75433 413185
rect 75533 413085 75601 413185
rect 75701 413085 75769 413185
rect 75869 413085 75937 413185
rect 76037 413085 76190 413185
rect 74052 413027 76190 413085
rect 74052 412927 74761 413027
rect 74861 412927 74929 413027
rect 75029 412927 75097 413027
rect 75197 412927 75265 413027
rect 75365 412927 75433 413027
rect 75533 412927 75601 413027
rect 75701 412927 75769 413027
rect 75869 412927 75937 413027
rect 76037 412927 76190 413027
rect 74052 412869 76190 412927
rect 74052 412769 74761 412869
rect 74861 412769 74929 412869
rect 75029 412769 75097 412869
rect 75197 412769 75265 412869
rect 75365 412769 75433 412869
rect 75533 412769 75601 412869
rect 75701 412769 75769 412869
rect 75869 412769 75937 412869
rect 76037 412769 76190 412869
rect 74052 412711 76190 412769
rect 74052 412707 74761 412711
rect 74676 412611 74761 412707
rect 74861 412611 74929 412711
rect 75029 412611 75097 412711
rect 75197 412611 75265 412711
rect 75365 412611 75433 412711
rect 75533 412611 75601 412711
rect 75701 412611 75769 412711
rect 75869 412611 75937 412711
rect 76037 412611 76190 412711
rect 74676 412310 76190 412611
rect 82014 401326 83235 414312
rect 73768 401250 83235 401326
rect 74854 401034 83235 401250
rect 73984 400958 83235 401034
rect 73984 400812 74944 400888
rect 74306 400684 74944 400812
rect 74306 400658 74797 400684
rect 74306 400640 74585 400658
rect 74306 400564 74415 400640
rect 74491 400582 74585 400640
rect 74661 400608 74797 400658
rect 74873 400608 74944 400684
rect 74661 400582 74944 400608
rect 74491 400564 74944 400582
rect 74306 400534 74944 400564
rect 74306 400458 74776 400534
rect 74852 400458 74944 400534
rect 74306 400384 74944 400458
rect 74306 400377 74775 400384
rect 74306 400371 74564 400377
rect 74306 400295 74394 400371
rect 74470 400301 74564 400371
rect 74640 400308 74775 400377
rect 74851 400308 74944 400384
rect 74640 400301 74944 400308
rect 74470 400295 74944 400301
rect 74306 400239 74944 400295
rect 82014 394388 83235 400958
rect 73984 394312 83235 394388
rect 74713 393951 76091 394003
rect 74713 393867 74779 393951
rect 74053 393851 74779 393867
rect 74879 393851 74947 393951
rect 75047 393851 75115 393951
rect 75215 393851 75283 393951
rect 75383 393851 75451 393951
rect 75551 393851 75619 393951
rect 75719 393851 75787 393951
rect 75887 393851 75955 393951
rect 76055 393851 76091 393951
rect 74053 393793 76091 393851
rect 74053 393693 74779 393793
rect 74879 393693 74947 393793
rect 75047 393693 75115 393793
rect 75215 393693 75283 393793
rect 75383 393693 75451 393793
rect 75551 393693 75619 393793
rect 75719 393693 75787 393793
rect 75887 393693 75955 393793
rect 76055 393693 76091 393793
rect 74053 393635 76091 393693
rect 74053 393535 74779 393635
rect 74879 393535 74947 393635
rect 75047 393535 75115 393635
rect 75215 393535 75283 393635
rect 75383 393535 75451 393635
rect 75551 393535 75619 393635
rect 75719 393535 75787 393635
rect 75887 393535 75955 393635
rect 76055 393535 76091 393635
rect 74053 393477 76091 393535
rect 74053 393377 74779 393477
rect 74879 393377 74947 393477
rect 75047 393377 75115 393477
rect 75215 393377 75283 393477
rect 75383 393377 75451 393477
rect 75551 393377 75619 393477
rect 75719 393377 75787 393477
rect 75887 393377 75955 393477
rect 76055 393377 76091 393477
rect 74053 393319 76091 393377
rect 74053 393219 74779 393319
rect 74879 393219 74947 393319
rect 75047 393219 75115 393319
rect 75215 393219 75283 393319
rect 75383 393219 75451 393319
rect 75551 393219 75619 393319
rect 75719 393219 75787 393319
rect 75887 393219 75955 393319
rect 76055 393219 76091 393319
rect 74053 393161 76091 393219
rect 74053 393061 74779 393161
rect 74879 393061 74947 393161
rect 75047 393061 75115 393161
rect 75215 393061 75283 393161
rect 75383 393061 75451 393161
rect 75551 393061 75619 393161
rect 75719 393061 75787 393161
rect 75887 393061 75955 393161
rect 76055 393061 76091 393161
rect 74053 393003 76091 393061
rect 74053 392903 74779 393003
rect 74879 392903 74947 393003
rect 75047 392903 75115 393003
rect 75215 392903 75283 393003
rect 75383 392903 75451 393003
rect 75551 392903 75619 393003
rect 75719 392903 75787 393003
rect 75887 392903 75955 393003
rect 76055 392903 76091 393003
rect 74053 392845 76091 392903
rect 74053 392745 74779 392845
rect 74879 392745 74947 392845
rect 75047 392745 75115 392845
rect 75215 392745 75283 392845
rect 75383 392745 75451 392845
rect 75551 392745 75619 392845
rect 75719 392745 75787 392845
rect 75887 392745 75955 392845
rect 76055 392745 76091 392845
rect 74053 392708 75210 392745
rect 75288 392717 76091 392745
rect 75288 392708 75934 392717
rect 74053 392707 74882 392708
rect 82014 381327 83235 394312
rect 74693 381326 83235 381327
rect 73984 381250 83235 381326
rect 74693 381034 83235 381250
rect 73984 380958 83235 381034
rect 73984 380812 74770 380888
rect 74131 380735 74770 380812
rect 74131 380684 74769 380735
rect 74131 380658 74622 380684
rect 74131 380640 74410 380658
rect 74131 380564 74240 380640
rect 74316 380582 74410 380640
rect 74486 380608 74622 380658
rect 74698 380608 74769 380684
rect 74486 380582 74769 380608
rect 74316 380564 74769 380582
rect 74131 380534 74769 380564
rect 74131 380458 74601 380534
rect 74677 380458 74769 380534
rect 74131 380384 74769 380458
rect 74131 380377 74600 380384
rect 74131 380371 74389 380377
rect 74131 380295 74219 380371
rect 74295 380301 74389 380371
rect 74465 380308 74600 380377
rect 74676 380308 74769 380384
rect 74465 380301 74769 380308
rect 74295 380295 74769 380301
rect 74131 380239 74769 380295
rect 82014 367232 83235 380958
rect 121127 367465 127852 367981
rect 121127 367315 122043 367465
rect 122193 367315 122311 367465
rect 122461 367315 122579 367465
rect 122729 367315 122847 367465
rect 122997 367315 123115 367465
rect 123265 367315 123383 367465
rect 123533 367315 123651 367465
rect 123801 367315 123919 367465
rect 124069 367315 124187 367465
rect 124337 367315 124455 367465
rect 124605 367315 127852 367465
rect 121127 367232 127852 367315
rect 72010 367227 127852 367232
rect 72010 367077 122043 367227
rect 122193 367077 122311 367227
rect 122461 367077 122579 367227
rect 122729 367077 122847 367227
rect 122997 367077 123115 367227
rect 123265 367077 123383 367227
rect 123533 367077 123651 367227
rect 123801 367077 123919 367227
rect 124069 367077 124187 367227
rect 124337 367077 124455 367227
rect 124605 367077 127852 367227
rect 72010 366989 127852 367077
rect 72010 366839 122043 366989
rect 122193 366839 122311 366989
rect 122461 366839 122579 366989
rect 122729 366839 122847 366989
rect 122997 366839 123115 366989
rect 123265 366839 123383 366989
rect 123533 366839 123651 366989
rect 123801 366839 123919 366989
rect 124069 366839 124187 366989
rect 124337 366839 124455 366989
rect 124605 366839 127852 366989
rect 72010 366751 127852 366839
rect 72010 366601 122043 366751
rect 122193 366601 122311 366751
rect 122461 366601 122579 366751
rect 122729 366601 122847 366751
rect 122997 366601 123115 366751
rect 123265 366601 123383 366751
rect 123533 366601 123651 366751
rect 123801 366601 123919 366751
rect 124069 366601 124187 366751
rect 124337 366601 124455 366751
rect 124605 366601 127852 366751
rect 72010 366513 127852 366601
rect 72010 366363 122043 366513
rect 122193 366363 122311 366513
rect 122461 366363 122579 366513
rect 122729 366363 122847 366513
rect 122997 366363 123115 366513
rect 123265 366363 123383 366513
rect 123533 366363 123651 366513
rect 123801 366363 123919 366513
rect 124069 366363 124187 366513
rect 124337 366363 124455 366513
rect 124605 366363 127852 366513
rect 72010 366275 127852 366363
rect 72010 366125 122043 366275
rect 122193 366125 122311 366275
rect 122461 366125 122579 366275
rect 122729 366125 122847 366275
rect 122997 366125 123115 366275
rect 123265 366125 123383 366275
rect 123533 366125 123651 366275
rect 123801 366125 123919 366275
rect 124069 366125 124187 366275
rect 124337 366125 124455 366275
rect 124605 366125 127852 366275
rect 72010 366037 127852 366125
rect 72010 365887 122043 366037
rect 122193 365887 122311 366037
rect 122461 365887 122579 366037
rect 122729 365887 122847 366037
rect 122997 365887 123115 366037
rect 123265 365887 123383 366037
rect 123533 365887 123651 366037
rect 123801 365887 123919 366037
rect 124069 365887 124187 366037
rect 124337 365887 124455 366037
rect 124605 365887 127852 366037
rect 72010 365799 127852 365887
rect 72010 365649 122043 365799
rect 122193 365649 122311 365799
rect 122461 365649 122579 365799
rect 122729 365649 122847 365799
rect 122997 365649 123115 365799
rect 123265 365649 123383 365799
rect 123533 365649 123651 365799
rect 123801 365649 123919 365799
rect 124069 365649 124187 365799
rect 124337 365649 124455 365799
rect 124605 365649 127852 365799
rect 72010 365561 127852 365649
rect 72010 365411 122043 365561
rect 122193 365411 122311 365561
rect 122461 365411 122579 365561
rect 122729 365411 122847 365561
rect 122997 365411 123115 365561
rect 123265 365411 123383 365561
rect 123533 365411 123651 365561
rect 123801 365411 123919 365561
rect 124069 365411 124187 365561
rect 124337 365411 124455 365561
rect 124605 365411 127852 365561
rect 72010 365323 127852 365411
rect 72010 365182 122043 365323
rect 81074 354454 83124 365182
rect 121077 365173 122043 365182
rect 122193 365173 122311 365323
rect 122461 365173 122579 365323
rect 122729 365173 122847 365323
rect 122997 365173 123115 365323
rect 123265 365173 123383 365323
rect 123533 365173 123651 365323
rect 123801 365173 123919 365323
rect 124069 365173 124187 365323
rect 124337 365173 124455 365323
rect 124605 365173 127852 365323
rect 121077 365066 127852 365173
rect 121127 364498 127852 365066
rect 73745 354247 83124 354454
rect 73983 353842 75995 353868
rect 73983 353790 75996 353842
rect 74028 353690 74684 353790
rect 74784 353690 74852 353790
rect 74952 353690 75020 353790
rect 75120 353690 75188 353790
rect 75288 353690 75356 353790
rect 75456 353690 75524 353790
rect 75624 353690 75692 353790
rect 75792 353690 75860 353790
rect 75960 353690 75996 353790
rect 74028 353632 75996 353690
rect 74028 353532 74684 353632
rect 74784 353532 74852 353632
rect 74952 353532 75020 353632
rect 75120 353532 75188 353632
rect 75288 353532 75356 353632
rect 75456 353532 75524 353632
rect 75624 353532 75692 353632
rect 75792 353532 75860 353632
rect 75960 353532 75996 353632
rect 74028 353474 75996 353532
rect 74028 353374 74684 353474
rect 74784 353374 74852 353474
rect 74952 353374 75020 353474
rect 75120 353374 75188 353474
rect 75288 353374 75356 353474
rect 75456 353374 75524 353474
rect 75624 353374 75692 353474
rect 75792 353374 75860 353474
rect 75960 353374 75996 353474
rect 74028 353316 75996 353374
rect 74028 353216 74684 353316
rect 74784 353216 74852 353316
rect 74952 353216 75020 353316
rect 75120 353216 75188 353316
rect 75288 353216 75356 353316
rect 75456 353216 75524 353316
rect 75624 353216 75692 353316
rect 75792 353216 75860 353316
rect 75960 353216 75996 353316
rect 74028 353158 75996 353216
rect 74028 353058 74684 353158
rect 74784 353058 74852 353158
rect 74952 353058 75020 353158
rect 75120 353058 75188 353158
rect 75288 353058 75356 353158
rect 75456 353058 75524 353158
rect 75624 353058 75692 353158
rect 75792 353058 75860 353158
rect 75960 353058 75996 353158
rect 74028 353000 75996 353058
rect 74028 352900 74684 353000
rect 74784 352900 74852 353000
rect 74952 352900 75020 353000
rect 75120 352900 75188 353000
rect 75288 352900 75356 353000
rect 75456 352900 75524 353000
rect 75624 352900 75692 353000
rect 75792 352900 75860 353000
rect 75960 352900 75996 353000
rect 74028 352842 75996 352900
rect 74028 352783 74684 352842
rect 73984 352742 74684 352783
rect 74784 352742 74852 352842
rect 74952 352742 75020 352842
rect 75120 352742 75188 352842
rect 75288 352742 75356 352842
rect 75456 352742 75524 352842
rect 75624 352742 75692 352842
rect 75792 352742 75860 352842
rect 75960 352742 75996 352842
rect 73984 352707 75996 352742
rect 74618 352684 75996 352707
rect 74618 352584 74684 352684
rect 74784 352584 74852 352684
rect 74952 352584 75020 352684
rect 75120 352584 75188 352684
rect 75288 352584 75356 352684
rect 75456 352584 75524 352684
rect 75624 352584 75692 352684
rect 75792 352584 75860 352684
rect 75960 352584 75996 352684
rect 74618 352547 75210 352584
rect 75288 352556 75996 352584
rect 75288 352547 75839 352556
rect 81074 341326 83124 354247
rect 73984 341250 83124 341326
rect 74351 341034 83124 341250
rect 73984 340958 83124 341034
rect 73984 340812 74833 340888
rect 74194 340687 74833 340812
rect 74194 340660 74832 340687
rect 74194 340634 74685 340660
rect 74194 340616 74473 340634
rect 74194 340540 74303 340616
rect 74379 340558 74473 340616
rect 74549 340584 74685 340634
rect 74761 340584 74832 340660
rect 74549 340558 74832 340584
rect 74379 340540 74832 340558
rect 74194 340510 74832 340540
rect 74194 340434 74664 340510
rect 74740 340434 74832 340510
rect 74194 340360 74832 340434
rect 74194 340353 74663 340360
rect 74194 340347 74452 340353
rect 74194 340271 74282 340347
rect 74358 340277 74452 340347
rect 74528 340284 74663 340353
rect 74739 340284 74832 340360
rect 74528 340277 74832 340284
rect 74358 340271 74832 340277
rect 74194 340215 74832 340271
rect 81074 334459 83124 340958
rect 73755 334393 83124 334459
rect 73749 334307 83124 334393
rect 73755 334242 83124 334307
rect 74053 333805 75938 333867
rect 74053 333705 74626 333805
rect 74726 333705 74794 333805
rect 74894 333705 74962 333805
rect 75062 333705 75130 333805
rect 75230 333705 75298 333805
rect 75398 333705 75466 333805
rect 75566 333705 75634 333805
rect 75734 333705 75802 333805
rect 75902 333705 75938 333805
rect 74053 333647 75938 333705
rect 74053 333547 74626 333647
rect 74726 333547 74794 333647
rect 74894 333547 74962 333647
rect 75062 333547 75130 333647
rect 75230 333547 75298 333647
rect 75398 333547 75466 333647
rect 75566 333547 75634 333647
rect 75734 333547 75802 333647
rect 75902 333547 75938 333647
rect 74053 333489 75938 333547
rect 74053 333389 74626 333489
rect 74726 333389 74794 333489
rect 74894 333389 74962 333489
rect 75062 333389 75130 333489
rect 75230 333389 75298 333489
rect 75398 333389 75466 333489
rect 75566 333389 75634 333489
rect 75734 333389 75802 333489
rect 75902 333389 75938 333489
rect 74053 333331 75938 333389
rect 74053 333231 74626 333331
rect 74726 333231 74794 333331
rect 74894 333231 74962 333331
rect 75062 333231 75130 333331
rect 75230 333231 75298 333331
rect 75398 333231 75466 333331
rect 75566 333231 75634 333331
rect 75734 333231 75802 333331
rect 75902 333231 75938 333331
rect 74053 333173 75938 333231
rect 74053 333073 74626 333173
rect 74726 333073 74794 333173
rect 74894 333073 74962 333173
rect 75062 333073 75130 333173
rect 75230 333073 75298 333173
rect 75398 333073 75466 333173
rect 75566 333073 75634 333173
rect 75734 333073 75802 333173
rect 75902 333073 75938 333173
rect 74053 333015 75938 333073
rect 74053 332915 74626 333015
rect 74726 332915 74794 333015
rect 74894 332915 74962 333015
rect 75062 332915 75130 333015
rect 75230 332915 75298 333015
rect 75398 332915 75466 333015
rect 75566 332915 75634 333015
rect 75734 332915 75802 333015
rect 75902 332915 75938 333015
rect 74053 332857 75938 332915
rect 74053 332757 74626 332857
rect 74726 332757 74794 332857
rect 74894 332757 74962 332857
rect 75062 332757 75130 332857
rect 75230 332757 75298 332857
rect 75398 332757 75466 332857
rect 75566 332757 75634 332857
rect 75734 332757 75802 332857
rect 75902 332757 75938 332857
rect 74053 332707 75938 332757
rect 74560 332699 75938 332707
rect 74560 332599 74626 332699
rect 74726 332599 74794 332699
rect 74894 332599 74962 332699
rect 75062 332599 75130 332699
rect 75230 332599 75298 332699
rect 75398 332599 75466 332699
rect 75566 332599 75634 332699
rect 75734 332599 75802 332699
rect 75902 332599 75938 332699
rect 74560 332571 75938 332599
rect 74560 332562 75781 332571
rect 81074 321326 83124 334242
rect 73984 321250 83125 321326
rect 74424 321034 83125 321250
rect 73984 320958 83125 321034
rect 73984 320812 74818 320888
rect 74144 320652 74818 320812
rect 74144 320626 74671 320652
rect 74144 320608 74459 320626
rect 74144 320532 74289 320608
rect 74365 320550 74459 320608
rect 74535 320576 74671 320626
rect 74747 320576 74818 320652
rect 74535 320550 74818 320576
rect 74365 320532 74818 320550
rect 74144 320502 74818 320532
rect 74144 320426 74650 320502
rect 74726 320426 74818 320502
rect 74144 320352 74818 320426
rect 74144 320345 74649 320352
rect 74144 320339 74438 320345
rect 74144 320263 74268 320339
rect 74344 320269 74438 320339
rect 74514 320276 74649 320345
rect 74725 320276 74818 320352
rect 74514 320269 74818 320276
rect 74344 320263 74818 320269
rect 74144 320207 74818 320263
<< via2 >>
rect 91879 467431 92029 467581
rect 92147 467431 92297 467581
rect 92415 467431 92565 467581
rect 92683 467431 92833 467581
rect 92951 467431 93101 467581
rect 93219 467431 93369 467581
rect 93487 467431 93637 467581
rect 93755 467431 93905 467581
rect 94023 467431 94173 467581
rect 94291 467431 94441 467581
rect 91879 467193 92029 467343
rect 92147 467193 92297 467343
rect 92415 467193 92565 467343
rect 92683 467193 92833 467343
rect 92951 467193 93101 467343
rect 93219 467193 93369 467343
rect 93487 467193 93637 467343
rect 93755 467193 93905 467343
rect 94023 467193 94173 467343
rect 94291 467193 94441 467343
rect 91879 466955 92029 467105
rect 92147 466955 92297 467105
rect 92415 466955 92565 467105
rect 92683 466955 92833 467105
rect 92951 466955 93101 467105
rect 93219 466955 93369 467105
rect 93487 466955 93637 467105
rect 93755 466955 93905 467105
rect 94023 466955 94173 467105
rect 94291 466955 94441 467105
rect 91879 466717 92029 466867
rect 92147 466717 92297 466867
rect 92415 466717 92565 466867
rect 92683 466717 92833 466867
rect 92951 466717 93101 466867
rect 93219 466717 93369 466867
rect 93487 466717 93637 466867
rect 93755 466717 93905 466867
rect 94023 466717 94173 466867
rect 94291 466717 94441 466867
rect 91879 466479 92029 466629
rect 92147 466479 92297 466629
rect 92415 466479 92565 466629
rect 92683 466479 92833 466629
rect 92951 466479 93101 466629
rect 93219 466479 93369 466629
rect 93487 466479 93637 466629
rect 93755 466479 93905 466629
rect 94023 466479 94173 466629
rect 94291 466479 94441 466629
rect 91879 466241 92029 466391
rect 92147 466241 92297 466391
rect 92415 466241 92565 466391
rect 92683 466241 92833 466391
rect 92951 466241 93101 466391
rect 93219 466241 93369 466391
rect 93487 466241 93637 466391
rect 93755 466241 93905 466391
rect 94023 466241 94173 466391
rect 94291 466241 94441 466391
rect 91879 466003 92029 466153
rect 92147 466003 92297 466153
rect 92415 466003 92565 466153
rect 92683 466003 92833 466153
rect 92951 466003 93101 466153
rect 93219 466003 93369 466153
rect 93487 466003 93637 466153
rect 93755 466003 93905 466153
rect 94023 466003 94173 466153
rect 94291 466003 94441 466153
rect 91879 465765 92029 465915
rect 92147 465765 92297 465915
rect 92415 465765 92565 465915
rect 92683 465765 92833 465915
rect 92951 465765 93101 465915
rect 93219 465765 93369 465915
rect 93487 465765 93637 465915
rect 93755 465765 93905 465915
rect 94023 465765 94173 465915
rect 94291 465765 94441 465915
rect 91879 465527 92029 465677
rect 92147 465527 92297 465677
rect 92415 465527 92565 465677
rect 92683 465527 92833 465677
rect 92951 465527 93101 465677
rect 93219 465527 93369 465677
rect 93487 465527 93637 465677
rect 93755 465527 93905 465677
rect 94023 465527 94173 465677
rect 94291 465527 94441 465677
rect 91879 465289 92029 465439
rect 92147 465289 92297 465439
rect 92415 465289 92565 465439
rect 92683 465289 92833 465439
rect 92951 465289 93101 465439
rect 93219 465289 93369 465439
rect 93487 465289 93637 465439
rect 93755 465289 93905 465439
rect 94023 465289 94173 465439
rect 94291 465289 94441 465439
rect 123379 457241 124600 458462
rect 123282 455399 124503 456620
rect 125479 455561 126700 456782
rect 77983 453392 78116 453525
rect 77981 453140 78114 453273
rect 77991 452749 78124 452882
rect 123056 453202 124277 454423
rect 125729 452148 126950 453369
rect 122862 450908 124083 452129
rect 122765 448355 123986 449576
rect 125729 448419 126950 449640
rect 122603 446028 123824 447249
rect 125729 445973 126950 447194
rect 74642 433654 74742 433754
rect 74810 433654 74910 433754
rect 74978 433654 75078 433754
rect 75146 433654 75246 433754
rect 75314 433654 75414 433754
rect 75482 433654 75582 433754
rect 75650 433654 75750 433754
rect 75818 433654 75918 433754
rect 74642 433496 74742 433596
rect 74810 433496 74910 433596
rect 74978 433496 75078 433596
rect 75146 433496 75246 433596
rect 75314 433496 75414 433596
rect 75482 433496 75582 433596
rect 75650 433496 75750 433596
rect 75818 433496 75918 433596
rect 74642 433338 74742 433438
rect 74810 433338 74910 433438
rect 74978 433338 75078 433438
rect 75146 433338 75246 433438
rect 75314 433338 75414 433438
rect 75482 433338 75582 433438
rect 75650 433338 75750 433438
rect 75818 433338 75918 433438
rect 74642 433180 74742 433280
rect 74810 433180 74910 433280
rect 74978 433180 75078 433280
rect 75146 433180 75246 433280
rect 75314 433180 75414 433280
rect 75482 433180 75582 433280
rect 75650 433180 75750 433280
rect 75818 433180 75918 433280
rect 74642 433022 74742 433122
rect 74810 433022 74910 433122
rect 74978 433022 75078 433122
rect 75146 433022 75246 433122
rect 75314 433022 75414 433122
rect 75482 433022 75582 433122
rect 75650 433022 75750 433122
rect 75818 433022 75918 433122
rect 74642 432864 74742 432964
rect 74810 432864 74910 432964
rect 74978 432864 75078 432964
rect 75146 432864 75246 432964
rect 75314 432864 75414 432964
rect 75482 432864 75582 432964
rect 75650 432864 75750 432964
rect 75818 432864 75918 432964
rect 74642 432706 74742 432806
rect 74810 432706 74910 432806
rect 74978 432706 75078 432806
rect 75146 432706 75246 432806
rect 75314 432706 75414 432806
rect 75482 432706 75582 432806
rect 75650 432706 75750 432806
rect 75818 432706 75918 432806
rect 74642 432548 74742 432648
rect 74810 432548 74910 432648
rect 74978 432548 75078 432648
rect 75146 432548 75246 432648
rect 75314 432548 75414 432648
rect 75482 432548 75582 432648
rect 75650 432548 75750 432648
rect 75818 432548 75918 432648
rect 74761 413717 74861 413817
rect 74929 413717 75029 413817
rect 75097 413717 75197 413817
rect 75265 413717 75365 413817
rect 75433 413717 75533 413817
rect 75601 413717 75701 413817
rect 75769 413717 75869 413817
rect 75937 413717 76037 413817
rect 74761 413559 74861 413659
rect 74929 413559 75029 413659
rect 75097 413559 75197 413659
rect 75265 413559 75365 413659
rect 75433 413559 75533 413659
rect 75601 413559 75701 413659
rect 75769 413559 75869 413659
rect 75937 413559 76037 413659
rect 74761 413401 74861 413501
rect 74929 413401 75029 413501
rect 75097 413401 75197 413501
rect 75265 413401 75365 413501
rect 75433 413401 75533 413501
rect 75601 413401 75701 413501
rect 75769 413401 75869 413501
rect 75937 413401 76037 413501
rect 74761 413243 74861 413343
rect 74929 413243 75029 413343
rect 75097 413243 75197 413343
rect 75265 413243 75365 413343
rect 75433 413243 75533 413343
rect 75601 413243 75701 413343
rect 75769 413243 75869 413343
rect 75937 413243 76037 413343
rect 74761 413085 74861 413185
rect 74929 413085 75029 413185
rect 75097 413085 75197 413185
rect 75265 413085 75365 413185
rect 75433 413085 75533 413185
rect 75601 413085 75701 413185
rect 75769 413085 75869 413185
rect 75937 413085 76037 413185
rect 74761 412927 74861 413027
rect 74929 412927 75029 413027
rect 75097 412927 75197 413027
rect 75265 412927 75365 413027
rect 75433 412927 75533 413027
rect 75601 412927 75701 413027
rect 75769 412927 75869 413027
rect 75937 412927 76037 413027
rect 74761 412769 74861 412869
rect 74929 412769 75029 412869
rect 75097 412769 75197 412869
rect 75265 412769 75365 412869
rect 75433 412769 75533 412869
rect 75601 412769 75701 412869
rect 75769 412769 75869 412869
rect 75937 412769 76037 412869
rect 74761 412611 74861 412711
rect 74929 412611 75029 412711
rect 75097 412611 75197 412711
rect 75265 412611 75365 412711
rect 75433 412611 75533 412711
rect 75601 412611 75701 412711
rect 75769 412611 75869 412711
rect 75937 412611 76037 412711
rect 74779 393851 74879 393951
rect 74947 393851 75047 393951
rect 75115 393851 75215 393951
rect 75283 393851 75383 393951
rect 75451 393851 75551 393951
rect 75619 393851 75719 393951
rect 75787 393851 75887 393951
rect 75955 393851 76055 393951
rect 74779 393693 74879 393793
rect 74947 393693 75047 393793
rect 75115 393693 75215 393793
rect 75283 393693 75383 393793
rect 75451 393693 75551 393793
rect 75619 393693 75719 393793
rect 75787 393693 75887 393793
rect 75955 393693 76055 393793
rect 74779 393535 74879 393635
rect 74947 393535 75047 393635
rect 75115 393535 75215 393635
rect 75283 393535 75383 393635
rect 75451 393535 75551 393635
rect 75619 393535 75719 393635
rect 75787 393535 75887 393635
rect 75955 393535 76055 393635
rect 74779 393377 74879 393477
rect 74947 393377 75047 393477
rect 75115 393377 75215 393477
rect 75283 393377 75383 393477
rect 75451 393377 75551 393477
rect 75619 393377 75719 393477
rect 75787 393377 75887 393477
rect 75955 393377 76055 393477
rect 74779 393219 74879 393319
rect 74947 393219 75047 393319
rect 75115 393219 75215 393319
rect 75283 393219 75383 393319
rect 75451 393219 75551 393319
rect 75619 393219 75719 393319
rect 75787 393219 75887 393319
rect 75955 393219 76055 393319
rect 74779 393061 74879 393161
rect 74947 393061 75047 393161
rect 75115 393061 75215 393161
rect 75283 393061 75383 393161
rect 75451 393061 75551 393161
rect 75619 393061 75719 393161
rect 75787 393061 75887 393161
rect 75955 393061 76055 393161
rect 74779 392903 74879 393003
rect 74947 392903 75047 393003
rect 75115 392903 75215 393003
rect 75283 392903 75383 393003
rect 75451 392903 75551 393003
rect 75619 392903 75719 393003
rect 75787 392903 75887 393003
rect 75955 392903 76055 393003
rect 74779 392745 74879 392845
rect 74947 392745 75047 392845
rect 75115 392745 75215 392845
rect 75283 392745 75383 392845
rect 75451 392745 75551 392845
rect 75619 392745 75719 392845
rect 75787 392745 75887 392845
rect 75955 392745 76055 392845
rect 122043 367315 122193 367465
rect 122311 367315 122461 367465
rect 122579 367315 122729 367465
rect 122847 367315 122997 367465
rect 123115 367315 123265 367465
rect 123383 367315 123533 367465
rect 123651 367315 123801 367465
rect 123919 367315 124069 367465
rect 124187 367315 124337 367465
rect 124455 367315 124605 367465
rect 122043 367077 122193 367227
rect 122311 367077 122461 367227
rect 122579 367077 122729 367227
rect 122847 367077 122997 367227
rect 123115 367077 123265 367227
rect 123383 367077 123533 367227
rect 123651 367077 123801 367227
rect 123919 367077 124069 367227
rect 124187 367077 124337 367227
rect 124455 367077 124605 367227
rect 122043 366839 122193 366989
rect 122311 366839 122461 366989
rect 122579 366839 122729 366989
rect 122847 366839 122997 366989
rect 123115 366839 123265 366989
rect 123383 366839 123533 366989
rect 123651 366839 123801 366989
rect 123919 366839 124069 366989
rect 124187 366839 124337 366989
rect 124455 366839 124605 366989
rect 122043 366601 122193 366751
rect 122311 366601 122461 366751
rect 122579 366601 122729 366751
rect 122847 366601 122997 366751
rect 123115 366601 123265 366751
rect 123383 366601 123533 366751
rect 123651 366601 123801 366751
rect 123919 366601 124069 366751
rect 124187 366601 124337 366751
rect 124455 366601 124605 366751
rect 122043 366363 122193 366513
rect 122311 366363 122461 366513
rect 122579 366363 122729 366513
rect 122847 366363 122997 366513
rect 123115 366363 123265 366513
rect 123383 366363 123533 366513
rect 123651 366363 123801 366513
rect 123919 366363 124069 366513
rect 124187 366363 124337 366513
rect 124455 366363 124605 366513
rect 122043 366125 122193 366275
rect 122311 366125 122461 366275
rect 122579 366125 122729 366275
rect 122847 366125 122997 366275
rect 123115 366125 123265 366275
rect 123383 366125 123533 366275
rect 123651 366125 123801 366275
rect 123919 366125 124069 366275
rect 124187 366125 124337 366275
rect 124455 366125 124605 366275
rect 122043 365887 122193 366037
rect 122311 365887 122461 366037
rect 122579 365887 122729 366037
rect 122847 365887 122997 366037
rect 123115 365887 123265 366037
rect 123383 365887 123533 366037
rect 123651 365887 123801 366037
rect 123919 365887 124069 366037
rect 124187 365887 124337 366037
rect 124455 365887 124605 366037
rect 122043 365649 122193 365799
rect 122311 365649 122461 365799
rect 122579 365649 122729 365799
rect 122847 365649 122997 365799
rect 123115 365649 123265 365799
rect 123383 365649 123533 365799
rect 123651 365649 123801 365799
rect 123919 365649 124069 365799
rect 124187 365649 124337 365799
rect 124455 365649 124605 365799
rect 122043 365411 122193 365561
rect 122311 365411 122461 365561
rect 122579 365411 122729 365561
rect 122847 365411 122997 365561
rect 123115 365411 123265 365561
rect 123383 365411 123533 365561
rect 123651 365411 123801 365561
rect 123919 365411 124069 365561
rect 124187 365411 124337 365561
rect 124455 365411 124605 365561
rect 122043 365173 122193 365323
rect 122311 365173 122461 365323
rect 122579 365173 122729 365323
rect 122847 365173 122997 365323
rect 123115 365173 123265 365323
rect 123383 365173 123533 365323
rect 123651 365173 123801 365323
rect 123919 365173 124069 365323
rect 124187 365173 124337 365323
rect 124455 365173 124605 365323
rect 74684 353690 74784 353790
rect 74852 353690 74952 353790
rect 75020 353690 75120 353790
rect 75188 353690 75288 353790
rect 75356 353690 75456 353790
rect 75524 353690 75624 353790
rect 75692 353690 75792 353790
rect 75860 353690 75960 353790
rect 74684 353532 74784 353632
rect 74852 353532 74952 353632
rect 75020 353532 75120 353632
rect 75188 353532 75288 353632
rect 75356 353532 75456 353632
rect 75524 353532 75624 353632
rect 75692 353532 75792 353632
rect 75860 353532 75960 353632
rect 74684 353374 74784 353474
rect 74852 353374 74952 353474
rect 75020 353374 75120 353474
rect 75188 353374 75288 353474
rect 75356 353374 75456 353474
rect 75524 353374 75624 353474
rect 75692 353374 75792 353474
rect 75860 353374 75960 353474
rect 74684 353216 74784 353316
rect 74852 353216 74952 353316
rect 75020 353216 75120 353316
rect 75188 353216 75288 353316
rect 75356 353216 75456 353316
rect 75524 353216 75624 353316
rect 75692 353216 75792 353316
rect 75860 353216 75960 353316
rect 74684 353058 74784 353158
rect 74852 353058 74952 353158
rect 75020 353058 75120 353158
rect 75188 353058 75288 353158
rect 75356 353058 75456 353158
rect 75524 353058 75624 353158
rect 75692 353058 75792 353158
rect 75860 353058 75960 353158
rect 74684 352900 74784 353000
rect 74852 352900 74952 353000
rect 75020 352900 75120 353000
rect 75188 352900 75288 353000
rect 75356 352900 75456 353000
rect 75524 352900 75624 353000
rect 75692 352900 75792 353000
rect 75860 352900 75960 353000
rect 74684 352742 74784 352842
rect 74852 352742 74952 352842
rect 75020 352742 75120 352842
rect 75188 352742 75288 352842
rect 75356 352742 75456 352842
rect 75524 352742 75624 352842
rect 75692 352742 75792 352842
rect 75860 352742 75960 352842
rect 74684 352584 74784 352684
rect 74852 352584 74952 352684
rect 75020 352584 75120 352684
rect 75188 352584 75288 352684
rect 75356 352584 75456 352684
rect 75524 352584 75624 352684
rect 75692 352584 75792 352684
rect 75860 352584 75960 352684
rect 74626 333705 74726 333805
rect 74794 333705 74894 333805
rect 74962 333705 75062 333805
rect 75130 333705 75230 333805
rect 75298 333705 75398 333805
rect 75466 333705 75566 333805
rect 75634 333705 75734 333805
rect 75802 333705 75902 333805
rect 74626 333547 74726 333647
rect 74794 333547 74894 333647
rect 74962 333547 75062 333647
rect 75130 333547 75230 333647
rect 75298 333547 75398 333647
rect 75466 333547 75566 333647
rect 75634 333547 75734 333647
rect 75802 333547 75902 333647
rect 74626 333389 74726 333489
rect 74794 333389 74894 333489
rect 74962 333389 75062 333489
rect 75130 333389 75230 333489
rect 75298 333389 75398 333489
rect 75466 333389 75566 333489
rect 75634 333389 75734 333489
rect 75802 333389 75902 333489
rect 74626 333231 74726 333331
rect 74794 333231 74894 333331
rect 74962 333231 75062 333331
rect 75130 333231 75230 333331
rect 75298 333231 75398 333331
rect 75466 333231 75566 333331
rect 75634 333231 75734 333331
rect 75802 333231 75902 333331
rect 74626 333073 74726 333173
rect 74794 333073 74894 333173
rect 74962 333073 75062 333173
rect 75130 333073 75230 333173
rect 75298 333073 75398 333173
rect 75466 333073 75566 333173
rect 75634 333073 75734 333173
rect 75802 333073 75902 333173
rect 74626 332915 74726 333015
rect 74794 332915 74894 333015
rect 74962 332915 75062 333015
rect 75130 332915 75230 333015
rect 75298 332915 75398 333015
rect 75466 332915 75566 333015
rect 75634 332915 75734 333015
rect 75802 332915 75902 333015
rect 74626 332757 74726 332857
rect 74794 332757 74894 332857
rect 74962 332757 75062 332857
rect 75130 332757 75230 332857
rect 75298 332757 75398 332857
rect 75466 332757 75566 332857
rect 75634 332757 75734 332857
rect 75802 332757 75902 332857
rect 74626 332599 74726 332699
rect 74794 332599 74894 332699
rect 74962 332599 75062 332699
rect 75130 332599 75230 332699
rect 75298 332599 75398 332699
rect 75466 332599 75566 332699
rect 75634 332599 75734 332699
rect 75802 332599 75902 332699
<< metal3 >>
rect 87832 510796 112357 510951
rect 87832 510096 87948 510796
rect 88648 510096 88929 510796
rect 89629 510096 89910 510796
rect 90610 510096 90891 510796
rect 91591 510096 91872 510796
rect 92572 510096 92853 510796
rect 93553 510096 93834 510796
rect 94534 510096 94815 510796
rect 95515 510096 95796 510796
rect 96496 510096 96777 510796
rect 97477 510096 97758 510796
rect 98458 510096 98739 510796
rect 99439 510096 99720 510796
rect 100420 510096 100701 510796
rect 101401 510096 101682 510796
rect 102382 510096 102663 510796
rect 103363 510096 103644 510796
rect 104344 510096 104625 510796
rect 105325 510096 105606 510796
rect 106306 510096 106587 510796
rect 107287 510096 107568 510796
rect 108268 510096 108549 510796
rect 109249 510096 109530 510796
rect 110230 510096 110511 510796
rect 111211 510096 111492 510796
rect 112192 510096 112357 510796
rect 87832 509776 112357 510096
rect 87832 509076 87948 509776
rect 88648 509076 88929 509776
rect 89629 509076 89910 509776
rect 90610 509076 90891 509776
rect 91591 509076 91872 509776
rect 92572 509076 92853 509776
rect 93553 509076 93834 509776
rect 94534 509076 94815 509776
rect 95515 509076 95796 509776
rect 96496 509076 96777 509776
rect 97477 509076 97758 509776
rect 98458 509076 98739 509776
rect 99439 509076 99720 509776
rect 100420 509076 100701 509776
rect 101401 509076 101682 509776
rect 102382 509076 102663 509776
rect 103363 509076 103644 509776
rect 104344 509076 104625 509776
rect 105325 509076 105606 509776
rect 106306 509076 106587 509776
rect 107287 509076 107568 509776
rect 108268 509076 108549 509776
rect 109249 509076 109530 509776
rect 110230 509076 110511 509776
rect 111211 509076 111492 509776
rect 112192 509076 112357 509776
rect 87832 508756 112357 509076
rect 87832 508056 87948 508756
rect 88648 508056 88929 508756
rect 89629 508056 89910 508756
rect 90610 508056 90891 508756
rect 91591 508056 91872 508756
rect 92572 508056 92853 508756
rect 93553 508056 93834 508756
rect 94534 508056 94815 508756
rect 95515 508056 95796 508756
rect 96496 508056 96777 508756
rect 97477 508056 97758 508756
rect 98458 508056 98739 508756
rect 99439 508056 99720 508756
rect 100420 508056 100701 508756
rect 101401 508056 101682 508756
rect 102382 508056 102663 508756
rect 103363 508056 103644 508756
rect 104344 508056 104625 508756
rect 105325 508056 105606 508756
rect 106306 508056 106587 508756
rect 107287 508056 107568 508756
rect 108268 508056 108549 508756
rect 109249 508056 109530 508756
rect 110230 508056 110511 508756
rect 111211 508056 111492 508756
rect 112192 508056 112357 508756
rect 87832 507736 112357 508056
rect 87832 507715 87948 507736
rect 87777 507036 87948 507715
rect 88648 507036 88929 507736
rect 89629 507036 89910 507736
rect 90610 507036 90891 507736
rect 91591 507036 91872 507736
rect 92572 507036 92853 507736
rect 93553 507036 93834 507736
rect 94534 507036 94815 507736
rect 95515 507036 95796 507736
rect 96496 507036 96777 507736
rect 97477 507036 97758 507736
rect 98458 507036 98739 507736
rect 99439 507036 99720 507736
rect 100420 507036 100701 507736
rect 101401 507036 101682 507736
rect 102382 507036 102663 507736
rect 103363 507036 103644 507736
rect 104344 507036 104625 507736
rect 105325 507036 105606 507736
rect 106306 507036 106587 507736
rect 107287 507036 107568 507736
rect 108268 507036 108549 507736
rect 109249 507036 109530 507736
rect 110230 507036 110511 507736
rect 111211 507036 111492 507736
rect 112192 507036 112357 507736
rect 482253 508075 507466 508386
rect 482253 507551 482569 508075
rect 87777 506716 112357 507036
rect 87777 506016 87948 506716
rect 88648 506016 88929 506716
rect 89629 506016 89910 506716
rect 90610 506016 90891 506716
rect 91591 506016 91872 506716
rect 92572 506016 92853 506716
rect 93553 506016 93834 506716
rect 94534 506016 94815 506716
rect 95515 506016 95796 506716
rect 96496 506016 96777 506716
rect 97477 506016 97758 506716
rect 98458 506016 98739 506716
rect 99439 506016 99720 506716
rect 100420 506016 100701 506716
rect 101401 506016 101682 506716
rect 102382 506016 102663 506716
rect 103363 506016 103644 506716
rect 104344 506016 104625 506716
rect 105325 506016 105606 506716
rect 106306 506016 106587 506716
rect 107287 506016 107568 506716
rect 108268 506016 108549 506716
rect 109249 506016 109530 506716
rect 110230 506016 110511 506716
rect 111211 506016 111492 506716
rect 112192 506030 112357 506716
rect 481938 507375 482569 507551
rect 483269 507375 483896 508075
rect 484596 507375 485223 508075
rect 485923 507375 486550 508075
rect 487250 507375 487877 508075
rect 488577 507375 489204 508075
rect 489904 507375 490531 508075
rect 491231 507375 491858 508075
rect 492558 507375 493185 508075
rect 493885 507375 494512 508075
rect 495212 507375 495839 508075
rect 496539 507375 497166 508075
rect 497866 507375 498493 508075
rect 499193 507375 499820 508075
rect 500520 507375 501147 508075
rect 501847 507375 502474 508075
rect 503174 507375 503801 508075
rect 504501 507375 505128 508075
rect 505828 507375 506455 508075
rect 507155 507375 507466 508075
rect 481938 506748 507466 507375
rect 481938 506048 482569 506748
rect 483269 506048 483896 506748
rect 484596 506048 485223 506748
rect 485923 506048 486550 506748
rect 487250 506048 487877 506748
rect 488577 506048 489204 506748
rect 489904 506048 490531 506748
rect 491231 506048 491858 506748
rect 492558 506048 493185 506748
rect 493885 506048 494512 506748
rect 495212 506048 495839 506748
rect 496539 506048 497166 506748
rect 497866 506048 498493 506748
rect 499193 506048 499820 506748
rect 500520 506048 501147 506748
rect 501847 506048 502474 506748
rect 503174 506048 503801 506748
rect 504501 506048 505128 506748
rect 505828 506048 506455 506748
rect 507155 506048 507466 506748
rect 481938 506030 507466 506048
rect 112192 506016 507466 506030
rect 87777 505696 507466 506016
rect 87777 504996 87948 505696
rect 88648 504996 88929 505696
rect 89629 504996 89910 505696
rect 90610 504996 90891 505696
rect 91591 504996 91872 505696
rect 92572 504996 92853 505696
rect 93553 504996 93834 505696
rect 94534 504996 94815 505696
rect 95515 504996 95796 505696
rect 96496 504996 96777 505696
rect 97477 504996 97758 505696
rect 98458 504996 98739 505696
rect 99439 504996 99720 505696
rect 100420 504996 100701 505696
rect 101401 504996 101682 505696
rect 102382 504996 102663 505696
rect 103363 504996 103644 505696
rect 104344 504996 104625 505696
rect 105325 504996 105606 505696
rect 106306 504996 106587 505696
rect 107287 504996 107568 505696
rect 108268 504996 108549 505696
rect 109249 504996 109530 505696
rect 110230 504996 110511 505696
rect 111211 504996 111492 505696
rect 112192 505421 507466 505696
rect 112192 504996 482569 505421
rect 87777 504721 482569 504996
rect 483269 504721 483896 505421
rect 484596 504721 485223 505421
rect 485923 504721 486550 505421
rect 487250 504721 487877 505421
rect 488577 504721 489204 505421
rect 489904 504721 490531 505421
rect 491231 504721 491858 505421
rect 492558 504721 493185 505421
rect 493885 504721 494512 505421
rect 495212 504721 495839 505421
rect 496539 504721 497166 505421
rect 497866 504721 498493 505421
rect 499193 504721 499820 505421
rect 500520 504721 501147 505421
rect 501847 504721 502474 505421
rect 503174 504721 503801 505421
rect 504501 504721 505128 505421
rect 505828 504721 506455 505421
rect 507155 504721 507466 505421
rect 87777 504676 507466 504721
rect 87777 503976 87948 504676
rect 88648 503976 88929 504676
rect 89629 503976 89910 504676
rect 90610 503976 90891 504676
rect 91591 503976 91872 504676
rect 92572 503976 92853 504676
rect 93553 503976 93834 504676
rect 94534 503976 94815 504676
rect 95515 503976 95796 504676
rect 96496 503976 96777 504676
rect 97477 503976 97758 504676
rect 98458 503976 98739 504676
rect 99439 503976 99720 504676
rect 100420 503976 100701 504676
rect 101401 503976 101682 504676
rect 102382 503976 102663 504676
rect 103363 503976 103644 504676
rect 104344 503976 104625 504676
rect 105325 503976 105606 504676
rect 106306 503976 106587 504676
rect 107287 503976 107568 504676
rect 108268 503976 108549 504676
rect 109249 503976 109530 504676
rect 110230 503976 110511 504676
rect 111211 503976 111492 504676
rect 112192 504094 507466 504676
rect 112192 503976 482569 504094
rect 87777 503656 482569 503976
rect 87777 502956 87948 503656
rect 88648 502956 88929 503656
rect 89629 502956 89910 503656
rect 90610 502956 90891 503656
rect 91591 502956 91872 503656
rect 92572 502956 92853 503656
rect 93553 502956 93834 503656
rect 94534 502956 94815 503656
rect 95515 502956 95796 503656
rect 96496 502956 96777 503656
rect 97477 502956 97758 503656
rect 98458 502956 98739 503656
rect 99439 502956 99720 503656
rect 100420 502956 100701 503656
rect 101401 502956 101682 503656
rect 102382 502956 102663 503656
rect 103363 502956 103644 503656
rect 104344 502956 104625 503656
rect 105325 502956 105606 503656
rect 106306 502956 106587 503656
rect 107287 502956 107568 503656
rect 108268 502956 108549 503656
rect 109249 502956 109530 503656
rect 110230 502956 110511 503656
rect 111211 502956 111492 503656
rect 112192 503394 482569 503656
rect 483269 503394 483896 504094
rect 484596 503394 485223 504094
rect 485923 503394 486550 504094
rect 487250 503394 487877 504094
rect 488577 503394 489204 504094
rect 489904 503394 490531 504094
rect 491231 503394 491858 504094
rect 492558 503394 493185 504094
rect 493885 503394 494512 504094
rect 495212 503394 495839 504094
rect 496539 503394 497166 504094
rect 497866 503394 498493 504094
rect 499193 503394 499820 504094
rect 500520 503394 501147 504094
rect 501847 503394 502474 504094
rect 503174 503394 503801 504094
rect 504501 503394 505128 504094
rect 505828 503394 506455 504094
rect 507155 503394 507466 504094
rect 112192 502956 507466 503394
rect 87777 502767 507466 502956
rect 87777 502636 482569 502767
rect 87777 501936 87948 502636
rect 88648 501936 88929 502636
rect 89629 501936 89910 502636
rect 90610 501936 90891 502636
rect 91591 501936 91872 502636
rect 92572 501936 92853 502636
rect 93553 501936 93834 502636
rect 94534 501936 94815 502636
rect 95515 501936 95796 502636
rect 96496 501936 96777 502636
rect 97477 501936 97758 502636
rect 98458 501936 98739 502636
rect 99439 501936 99720 502636
rect 100420 501936 100701 502636
rect 101401 501936 101682 502636
rect 102382 501936 102663 502636
rect 103363 501936 103644 502636
rect 104344 501936 104625 502636
rect 105325 501936 105606 502636
rect 106306 501936 106587 502636
rect 107287 501936 107568 502636
rect 108268 501936 108549 502636
rect 109249 501936 109530 502636
rect 110230 501936 110511 502636
rect 111211 501936 111492 502636
rect 112192 502067 482569 502636
rect 483269 502067 483896 502767
rect 484596 502067 485223 502767
rect 485923 502067 486550 502767
rect 487250 502067 487877 502767
rect 488577 502067 489204 502767
rect 489904 502067 490531 502767
rect 491231 502067 491858 502767
rect 492558 502067 493185 502767
rect 493885 502067 494512 502767
rect 495212 502067 495839 502767
rect 496539 502067 497166 502767
rect 497866 502067 498493 502767
rect 499193 502067 499820 502767
rect 500520 502067 501147 502767
rect 501847 502067 502474 502767
rect 503174 502067 503801 502767
rect 504501 502067 505128 502767
rect 505828 502067 506455 502767
rect 507155 502067 507466 502767
rect 112192 501936 507466 502067
rect 87777 501616 507466 501936
rect 87777 500916 87948 501616
rect 88648 500916 88929 501616
rect 89629 500916 89910 501616
rect 90610 500916 90891 501616
rect 91591 500916 91872 501616
rect 92572 500916 92853 501616
rect 93553 500916 93834 501616
rect 94534 500916 94815 501616
rect 95515 500916 95796 501616
rect 96496 500916 96777 501616
rect 97477 500916 97758 501616
rect 98458 500916 98739 501616
rect 99439 500916 99720 501616
rect 100420 500916 100701 501616
rect 101401 500916 101682 501616
rect 102382 500916 102663 501616
rect 103363 500916 103644 501616
rect 104344 500916 104625 501616
rect 105325 500916 105606 501616
rect 106306 500916 106587 501616
rect 107287 500916 107568 501616
rect 108268 500916 108549 501616
rect 109249 500916 109530 501616
rect 110230 500916 110511 501616
rect 111211 500916 111492 501616
rect 112192 501440 507466 501616
rect 112192 500916 482569 501440
rect 87777 500740 482569 500916
rect 483269 500740 483896 501440
rect 484596 500740 485223 501440
rect 485923 500740 486550 501440
rect 487250 500740 487877 501440
rect 488577 500740 489204 501440
rect 489904 500740 490531 501440
rect 491231 500740 491858 501440
rect 492558 500740 493185 501440
rect 493885 500740 494512 501440
rect 495212 500740 495839 501440
rect 496539 500740 497166 501440
rect 497866 500740 498493 501440
rect 499193 500740 499820 501440
rect 500520 500740 501147 501440
rect 501847 500740 502474 501440
rect 503174 500740 503801 501440
rect 504501 500740 505128 501440
rect 505828 500740 506455 501440
rect 507155 500740 507466 501440
rect 87777 500596 507466 500740
rect 87777 499896 87948 500596
rect 88648 499896 88929 500596
rect 89629 499896 89910 500596
rect 90610 499896 90891 500596
rect 91591 499896 91872 500596
rect 92572 499896 92853 500596
rect 93553 499896 93834 500596
rect 94534 499896 94815 500596
rect 95515 499896 95796 500596
rect 96496 499896 96777 500596
rect 97477 499896 97758 500596
rect 98458 499896 98739 500596
rect 99439 499896 99720 500596
rect 100420 499896 100701 500596
rect 101401 499896 101682 500596
rect 102382 499896 102663 500596
rect 103363 499896 103644 500596
rect 104344 499896 104625 500596
rect 105325 499896 105606 500596
rect 106306 499896 106587 500596
rect 107287 499896 107568 500596
rect 108268 499896 108549 500596
rect 109249 499896 109530 500596
rect 110230 499896 110511 500596
rect 111211 499896 111492 500596
rect 112192 500113 507466 500596
rect 112192 499896 482569 500113
rect 87777 499576 482569 499896
rect 87777 498876 87948 499576
rect 88648 498876 88929 499576
rect 89629 498876 89910 499576
rect 90610 498876 90891 499576
rect 91591 498876 91872 499576
rect 92572 498876 92853 499576
rect 93553 498876 93834 499576
rect 94534 498876 94815 499576
rect 95515 498876 95796 499576
rect 96496 498876 96777 499576
rect 97477 498876 97758 499576
rect 98458 498876 98739 499576
rect 99439 498876 99720 499576
rect 100420 498876 100701 499576
rect 101401 498876 101682 499576
rect 102382 498876 102663 499576
rect 103363 498876 103644 499576
rect 104344 498876 104625 499576
rect 105325 498876 105606 499576
rect 106306 498876 106587 499576
rect 107287 498876 107568 499576
rect 108268 498876 108549 499576
rect 109249 498876 109530 499576
rect 110230 498876 110511 499576
rect 111211 498876 111492 499576
rect 112192 499413 482569 499576
rect 483269 499413 483896 500113
rect 484596 499413 485223 500113
rect 485923 499413 486550 500113
rect 487250 499413 487877 500113
rect 488577 499413 489204 500113
rect 489904 499413 490531 500113
rect 491231 499413 491858 500113
rect 492558 499413 493185 500113
rect 493885 499413 494512 500113
rect 495212 499413 495839 500113
rect 496539 499413 497166 500113
rect 497866 499413 498493 500113
rect 499193 499413 499820 500113
rect 500520 499413 501147 500113
rect 501847 499413 502474 500113
rect 503174 499413 503801 500113
rect 504501 499413 505128 500113
rect 505828 499413 506455 500113
rect 507155 499413 507466 500113
rect 112192 498876 507466 499413
rect 87777 498786 507466 498876
rect 87777 498556 482569 498786
rect 87777 497856 87948 498556
rect 88648 497856 88929 498556
rect 89629 497856 89910 498556
rect 90610 497856 90891 498556
rect 91591 497856 91872 498556
rect 92572 497856 92853 498556
rect 93553 497856 93834 498556
rect 94534 497856 94815 498556
rect 95515 497856 95796 498556
rect 96496 497856 96777 498556
rect 97477 497856 97758 498556
rect 98458 497856 98739 498556
rect 99439 497856 99720 498556
rect 100420 497856 100701 498556
rect 101401 497856 101682 498556
rect 102382 497856 102663 498556
rect 103363 497856 103644 498556
rect 104344 497856 104625 498556
rect 105325 497856 105606 498556
rect 106306 497856 106587 498556
rect 107287 497856 107568 498556
rect 108268 497856 108549 498556
rect 109249 497856 109530 498556
rect 110230 497856 110511 498556
rect 111211 497856 111492 498556
rect 112192 498086 482569 498556
rect 483269 498086 483896 498786
rect 484596 498086 485223 498786
rect 485923 498086 486550 498786
rect 487250 498086 487877 498786
rect 488577 498086 489204 498786
rect 489904 498086 490531 498786
rect 491231 498086 491858 498786
rect 492558 498086 493185 498786
rect 493885 498086 494512 498786
rect 495212 498086 495839 498786
rect 496539 498086 497166 498786
rect 497866 498086 498493 498786
rect 499193 498086 499820 498786
rect 500520 498086 501147 498786
rect 501847 498086 502474 498786
rect 503174 498086 503801 498786
rect 504501 498086 505128 498786
rect 505828 498086 506455 498786
rect 507155 498086 507466 498786
rect 112192 497856 507466 498086
rect 87777 497536 507466 497856
rect 87777 496836 87948 497536
rect 88648 496836 88929 497536
rect 89629 496836 89910 497536
rect 90610 496836 90891 497536
rect 91591 496836 91872 497536
rect 92572 496836 92853 497536
rect 93553 496836 93834 497536
rect 94534 496836 94815 497536
rect 95515 496836 95796 497536
rect 96496 496836 96777 497536
rect 97477 496836 97758 497536
rect 98458 496836 98739 497536
rect 99439 496836 99720 497536
rect 100420 496836 100701 497536
rect 101401 496836 101682 497536
rect 102382 496836 102663 497536
rect 103363 496836 103644 497536
rect 104344 496836 104625 497536
rect 105325 496836 105606 497536
rect 106306 496836 106587 497536
rect 107287 496836 107568 497536
rect 108268 496836 108549 497536
rect 109249 496836 109530 497536
rect 110230 496836 110511 497536
rect 111211 496836 111492 497536
rect 112192 497459 507466 497536
rect 112192 496836 482569 497459
rect 87777 496759 482569 496836
rect 483269 496759 483896 497459
rect 484596 496759 485223 497459
rect 485923 496759 486550 497459
rect 487250 496759 487877 497459
rect 488577 496759 489204 497459
rect 489904 496759 490531 497459
rect 491231 496759 491858 497459
rect 492558 496759 493185 497459
rect 493885 496759 494512 497459
rect 495212 496759 495839 497459
rect 496539 496759 497166 497459
rect 497866 496759 498493 497459
rect 499193 496759 499820 497459
rect 500520 496759 501147 497459
rect 501847 496759 502474 497459
rect 503174 496759 503801 497459
rect 504501 496759 505128 497459
rect 505828 496759 506455 497459
rect 507155 496759 507466 497459
rect 87777 496516 507466 496759
rect 87777 495816 87948 496516
rect 88648 495816 88929 496516
rect 89629 495816 89910 496516
rect 90610 495816 90891 496516
rect 91591 495816 91872 496516
rect 92572 495816 92853 496516
rect 93553 495816 93834 496516
rect 94534 495816 94815 496516
rect 95515 495816 95796 496516
rect 96496 495816 96777 496516
rect 97477 495816 97758 496516
rect 98458 495816 98739 496516
rect 99439 495816 99720 496516
rect 100420 495816 100701 496516
rect 101401 495816 101682 496516
rect 102382 495816 102663 496516
rect 103363 495816 103644 496516
rect 104344 495816 104625 496516
rect 105325 495816 105606 496516
rect 106306 495816 106587 496516
rect 107287 495816 107568 496516
rect 108268 495816 108549 496516
rect 109249 495816 109530 496516
rect 110230 495816 110511 496516
rect 111211 495816 111492 496516
rect 112192 496132 507466 496516
rect 112192 495816 482569 496132
rect 87777 495496 482569 495816
rect 87777 494796 87948 495496
rect 88648 494796 88929 495496
rect 89629 494796 89910 495496
rect 90610 494796 90891 495496
rect 91591 494796 91872 495496
rect 92572 494796 92853 495496
rect 93553 494796 93834 495496
rect 94534 494796 94815 495496
rect 95515 494796 95796 495496
rect 96496 494796 96777 495496
rect 97477 494796 97758 495496
rect 98458 494796 98739 495496
rect 99439 494796 99720 495496
rect 100420 494796 100701 495496
rect 101401 494796 101682 495496
rect 102382 494796 102663 495496
rect 103363 494796 103644 495496
rect 104344 494796 104625 495496
rect 105325 494796 105606 495496
rect 106306 494796 106587 495496
rect 107287 494796 107568 495496
rect 108268 494796 108549 495496
rect 109249 494796 109530 495496
rect 110230 494796 110511 495496
rect 111211 494796 111492 495496
rect 112192 495432 482569 495496
rect 483269 495432 483896 496132
rect 484596 495432 485223 496132
rect 485923 495432 486550 496132
rect 487250 495432 487877 496132
rect 488577 495432 489204 496132
rect 489904 495432 490531 496132
rect 491231 495432 491858 496132
rect 492558 495432 493185 496132
rect 493885 495432 494512 496132
rect 495212 495432 495839 496132
rect 496539 495432 497166 496132
rect 497866 495432 498493 496132
rect 499193 495432 499820 496132
rect 500520 495432 501147 496132
rect 501847 495432 502474 496132
rect 503174 495432 503801 496132
rect 504501 495432 505128 496132
rect 505828 495432 506455 496132
rect 507155 495432 507466 496132
rect 112192 494805 507466 495432
rect 112192 494796 482569 494805
rect 87777 494476 482569 494796
rect 87777 493776 87948 494476
rect 88648 493776 88929 494476
rect 89629 493776 89910 494476
rect 90610 493776 90891 494476
rect 91591 493776 91872 494476
rect 92572 493776 92853 494476
rect 93553 493776 93834 494476
rect 94534 493776 94815 494476
rect 95515 493776 95796 494476
rect 96496 493776 96777 494476
rect 97477 493776 97758 494476
rect 98458 493776 98739 494476
rect 99439 493776 99720 494476
rect 100420 493776 100701 494476
rect 101401 493776 101682 494476
rect 102382 493776 102663 494476
rect 103363 493776 103644 494476
rect 104344 493776 104625 494476
rect 105325 493776 105606 494476
rect 106306 493776 106587 494476
rect 107287 493776 107568 494476
rect 108268 493776 108549 494476
rect 109249 493776 109530 494476
rect 110230 493776 110511 494476
rect 111211 493776 111492 494476
rect 112192 494105 482569 494476
rect 483269 494105 483896 494805
rect 484596 494105 485223 494805
rect 485923 494105 486550 494805
rect 487250 494105 487877 494805
rect 488577 494105 489204 494805
rect 489904 494105 490531 494805
rect 491231 494105 491858 494805
rect 492558 494105 493185 494805
rect 493885 494105 494512 494805
rect 495212 494105 495839 494805
rect 496539 494105 497166 494805
rect 497866 494105 498493 494805
rect 499193 494105 499820 494805
rect 500520 494105 501147 494805
rect 501847 494105 502474 494805
rect 503174 494105 503801 494805
rect 504501 494105 505128 494805
rect 505828 494105 506455 494805
rect 507155 494105 507466 494805
rect 112192 493776 507466 494105
rect 87777 493478 507466 493776
rect 87777 493456 482569 493478
rect 87777 492756 87948 493456
rect 88648 492756 88929 493456
rect 89629 492756 89910 493456
rect 90610 492756 90891 493456
rect 91591 492756 91872 493456
rect 92572 492756 92853 493456
rect 93553 492756 93834 493456
rect 94534 492756 94815 493456
rect 95515 492756 95796 493456
rect 96496 492756 96777 493456
rect 97477 492756 97758 493456
rect 98458 492756 98739 493456
rect 99439 492756 99720 493456
rect 100420 492756 100701 493456
rect 101401 492756 101682 493456
rect 102382 492756 102663 493456
rect 103363 492756 103644 493456
rect 104344 492756 104625 493456
rect 105325 492756 105606 493456
rect 106306 492756 106587 493456
rect 107287 492756 107568 493456
rect 108268 492756 108549 493456
rect 109249 492756 109530 493456
rect 110230 492756 110511 493456
rect 111211 492756 111492 493456
rect 112192 492778 482569 493456
rect 483269 492778 483896 493478
rect 484596 492778 485223 493478
rect 485923 492778 486550 493478
rect 487250 492778 487877 493478
rect 488577 492778 489204 493478
rect 489904 492778 490531 493478
rect 491231 492778 491858 493478
rect 492558 492778 493185 493478
rect 493885 492778 494512 493478
rect 495212 492778 495839 493478
rect 496539 492778 497166 493478
rect 497866 492778 498493 493478
rect 499193 492778 499820 493478
rect 500520 492778 501147 493478
rect 501847 492778 502474 493478
rect 503174 492778 503801 493478
rect 504501 492778 505128 493478
rect 505828 492778 506455 493478
rect 507155 492778 507466 493478
rect 112192 492756 507466 492778
rect 87777 492436 507466 492756
rect 87777 491736 87948 492436
rect 88648 491736 88929 492436
rect 89629 491736 89910 492436
rect 90610 491736 90891 492436
rect 91591 491736 91872 492436
rect 92572 491736 92853 492436
rect 93553 491736 93834 492436
rect 94534 491736 94815 492436
rect 95515 491736 95796 492436
rect 96496 491736 96777 492436
rect 97477 491736 97758 492436
rect 98458 491736 98739 492436
rect 99439 491736 99720 492436
rect 100420 491736 100701 492436
rect 101401 491736 101682 492436
rect 102382 491736 102663 492436
rect 103363 491736 103644 492436
rect 104344 491736 104625 492436
rect 105325 491736 105606 492436
rect 106306 491736 106587 492436
rect 107287 491736 107568 492436
rect 108268 491736 108549 492436
rect 109249 491736 109530 492436
rect 110230 491736 110511 492436
rect 111211 491736 111492 492436
rect 112192 492151 507466 492436
rect 112192 491736 482569 492151
rect 87777 491451 482569 491736
rect 483269 491451 483896 492151
rect 484596 491451 485223 492151
rect 485923 491451 486550 492151
rect 487250 491451 487877 492151
rect 488577 491451 489204 492151
rect 489904 491451 490531 492151
rect 491231 491451 491858 492151
rect 492558 491451 493185 492151
rect 493885 491451 494512 492151
rect 495212 491451 495839 492151
rect 496539 491451 497166 492151
rect 497866 491451 498493 492151
rect 499193 491451 499820 492151
rect 500520 491451 501147 492151
rect 501847 491451 502474 492151
rect 503174 491451 503801 492151
rect 504501 491451 505128 492151
rect 505828 491451 506455 492151
rect 507155 491451 507466 492151
rect 87777 491416 507466 491451
rect 87777 490716 87948 491416
rect 88648 490716 88929 491416
rect 89629 490716 89910 491416
rect 90610 490716 90891 491416
rect 91591 490716 91872 491416
rect 92572 490716 92853 491416
rect 93553 490716 93834 491416
rect 94534 490716 94815 491416
rect 95515 490716 95796 491416
rect 96496 490716 96777 491416
rect 97477 490716 97758 491416
rect 98458 490716 98739 491416
rect 99439 490716 99720 491416
rect 100420 490716 100701 491416
rect 101401 490716 101682 491416
rect 102382 490716 102663 491416
rect 103363 490716 103644 491416
rect 104344 490716 104625 491416
rect 105325 490716 105606 491416
rect 106306 490716 106587 491416
rect 107287 490716 107568 491416
rect 108268 490716 108549 491416
rect 109249 490716 109530 491416
rect 110230 490716 110511 491416
rect 111211 490716 111492 491416
rect 112192 490824 507466 491416
rect 112192 490716 482569 490824
rect 87777 490396 482569 490716
rect 87777 489696 87948 490396
rect 88648 489696 88929 490396
rect 89629 489696 89910 490396
rect 90610 489696 90891 490396
rect 91591 489696 91872 490396
rect 92572 489696 92853 490396
rect 93553 489696 93834 490396
rect 94534 489696 94815 490396
rect 95515 489696 95796 490396
rect 96496 489696 96777 490396
rect 97477 489696 97758 490396
rect 98458 489696 98739 490396
rect 99439 489696 99720 490396
rect 100420 489696 100701 490396
rect 101401 489696 101682 490396
rect 102382 489696 102663 490396
rect 103363 489696 103644 490396
rect 104344 489696 104625 490396
rect 105325 489696 105606 490396
rect 106306 489696 106587 490396
rect 107287 489696 107568 490396
rect 108268 489696 108549 490396
rect 109249 489696 109530 490396
rect 110230 489696 110511 490396
rect 111211 489696 111492 490396
rect 112192 490124 482569 490396
rect 483269 490124 483896 490824
rect 484596 490124 485223 490824
rect 485923 490124 486550 490824
rect 487250 490124 487877 490824
rect 488577 490124 489204 490824
rect 489904 490124 490531 490824
rect 491231 490124 491858 490824
rect 492558 490124 493185 490824
rect 493885 490124 494512 490824
rect 495212 490124 495839 490824
rect 496539 490124 497166 490824
rect 497866 490124 498493 490824
rect 499193 490124 499820 490824
rect 500520 490124 501147 490824
rect 501847 490124 502474 490824
rect 503174 490124 503801 490824
rect 504501 490124 505128 490824
rect 505828 490124 506455 490824
rect 507155 490124 507466 490824
rect 112192 489696 507466 490124
rect 87777 489497 507466 489696
rect 87777 489376 482569 489497
rect 87777 488676 87948 489376
rect 88648 488676 88929 489376
rect 89629 488676 89910 489376
rect 90610 488676 90891 489376
rect 91591 488676 91872 489376
rect 92572 488676 92853 489376
rect 93553 488676 93834 489376
rect 94534 488676 94815 489376
rect 95515 488676 95796 489376
rect 96496 488676 96777 489376
rect 97477 488676 97758 489376
rect 98458 488676 98739 489376
rect 99439 488676 99720 489376
rect 100420 488676 100701 489376
rect 101401 488676 101682 489376
rect 102382 488676 102663 489376
rect 103363 488676 103644 489376
rect 104344 488676 104625 489376
rect 105325 488676 105606 489376
rect 106306 488676 106587 489376
rect 107287 488676 107568 489376
rect 108268 488676 108549 489376
rect 109249 488676 109530 489376
rect 110230 488676 110511 489376
rect 111211 488676 111492 489376
rect 112192 488797 482569 489376
rect 483269 488797 483896 489497
rect 484596 488797 485223 489497
rect 485923 488797 486550 489497
rect 487250 488797 487877 489497
rect 488577 488797 489204 489497
rect 489904 488797 490531 489497
rect 491231 488797 491858 489497
rect 492558 488797 493185 489497
rect 493885 488797 494512 489497
rect 495212 488797 495839 489497
rect 496539 488797 497166 489497
rect 497866 488797 498493 489497
rect 499193 488797 499820 489497
rect 500520 488797 501147 489497
rect 501847 488797 502474 489497
rect 503174 488797 503801 489497
rect 504501 488797 505128 489497
rect 505828 488797 506455 489497
rect 507155 488797 507466 489497
rect 112192 488676 507466 488797
rect 87777 488356 507466 488676
rect 87777 487656 87948 488356
rect 88648 487656 88929 488356
rect 89629 487656 89910 488356
rect 90610 487656 90891 488356
rect 91591 487656 91872 488356
rect 92572 487656 92853 488356
rect 93553 487656 93834 488356
rect 94534 487656 94815 488356
rect 95515 487656 95796 488356
rect 96496 487656 96777 488356
rect 97477 487656 97758 488356
rect 98458 487656 98739 488356
rect 99439 487656 99720 488356
rect 100420 487656 100701 488356
rect 101401 487656 101682 488356
rect 102382 487656 102663 488356
rect 103363 487656 103644 488356
rect 104344 487656 104625 488356
rect 105325 487656 105606 488356
rect 106306 487656 106587 488356
rect 107287 487656 107568 488356
rect 108268 487656 108549 488356
rect 109249 487656 109530 488356
rect 110230 487656 110511 488356
rect 111211 487656 111492 488356
rect 112192 488170 507466 488356
rect 112192 487656 482569 488170
rect 87777 487470 482569 487656
rect 483269 487470 483896 488170
rect 484596 487470 485223 488170
rect 485923 487470 486550 488170
rect 487250 487470 487877 488170
rect 488577 487470 489204 488170
rect 489904 487470 490531 488170
rect 491231 487470 491858 488170
rect 492558 487470 493185 488170
rect 493885 487470 494512 488170
rect 495212 487470 495839 488170
rect 496539 487470 497166 488170
rect 497866 487470 498493 488170
rect 499193 487470 499820 488170
rect 500520 487470 501147 488170
rect 501847 487470 502474 488170
rect 503174 487470 503801 488170
rect 504501 487470 505128 488170
rect 505828 487470 506455 488170
rect 507155 487470 507466 488170
rect 87777 487336 507466 487470
rect 87777 486636 87948 487336
rect 88648 486636 88929 487336
rect 89629 486636 89910 487336
rect 90610 486636 90891 487336
rect 91591 486636 91872 487336
rect 92572 486636 92853 487336
rect 93553 486636 93834 487336
rect 94534 486636 94815 487336
rect 95515 486636 95796 487336
rect 96496 486636 96777 487336
rect 97477 486636 97758 487336
rect 98458 486636 98739 487336
rect 99439 486636 99720 487336
rect 100420 486636 100701 487336
rect 101401 486636 101682 487336
rect 102382 486636 102663 487336
rect 103363 486636 103644 487336
rect 104344 486636 104625 487336
rect 105325 486636 105606 487336
rect 106306 486636 106587 487336
rect 107287 486636 107568 487336
rect 108268 486636 108549 487336
rect 109249 486636 109530 487336
rect 110230 486636 110511 487336
rect 111211 486636 111492 487336
rect 112192 487085 507466 487336
rect 112192 486636 112357 487085
rect 87777 486316 112357 486636
rect 87777 485616 87948 486316
rect 88648 485616 88929 486316
rect 89629 485616 89910 486316
rect 90610 485616 90891 486316
rect 91591 485616 91872 486316
rect 92572 485616 92853 486316
rect 93553 485616 93834 486316
rect 94534 485616 94815 486316
rect 95515 485616 95796 486316
rect 96496 485616 96777 486316
rect 97477 485616 97758 486316
rect 98458 485616 98739 486316
rect 99439 485616 99720 486316
rect 100420 485616 100701 486316
rect 101401 485616 101682 486316
rect 102382 485616 102663 486316
rect 103363 485616 103644 486316
rect 104344 485616 104625 486316
rect 105325 485616 105606 486316
rect 106306 485616 106587 486316
rect 107287 485616 107568 486316
rect 108268 485616 108549 486316
rect 109249 485616 109530 486316
rect 110230 485616 110511 486316
rect 111211 485616 111492 486316
rect 112192 485616 112357 486316
rect 87777 485451 112357 485616
rect 481938 486843 507466 487085
rect 481938 486143 482569 486843
rect 483269 486143 483896 486843
rect 484596 486143 485223 486843
rect 485923 486143 486550 486843
rect 487250 486143 487877 486843
rect 488577 486143 489204 486843
rect 489904 486143 490531 486843
rect 491231 486143 491858 486843
rect 492558 486143 493185 486843
rect 493885 486143 494512 486843
rect 495212 486143 495839 486843
rect 496539 486143 497166 486843
rect 497866 486143 498493 486843
rect 499193 486143 499820 486843
rect 500520 486143 501147 486843
rect 501847 486143 502474 486843
rect 503174 486143 503801 486843
rect 504501 486143 505128 486843
rect 505828 486143 506455 486843
rect 507155 486143 507466 486843
rect 481938 485516 507466 486143
rect 87777 485163 110934 485451
rect 481938 484816 482569 485516
rect 483269 484816 483896 485516
rect 484596 484816 485223 485516
rect 485923 484816 486550 485516
rect 487250 484816 487877 485516
rect 488577 484816 489204 485516
rect 489904 484816 490531 485516
rect 491231 484816 491858 485516
rect 492558 484816 493185 485516
rect 493885 484816 494512 485516
rect 495212 484816 495839 485516
rect 496539 484816 497166 485516
rect 497866 484816 498493 485516
rect 499193 484816 499820 485516
rect 500520 484816 501147 485516
rect 501847 484816 502474 485516
rect 503174 484816 503801 485516
rect 504501 484816 505128 485516
rect 505828 484816 506455 485516
rect 507155 484816 507466 485516
rect 481938 484189 507466 484816
rect 481938 483489 482569 484189
rect 483269 483489 483896 484189
rect 484596 483489 485223 484189
rect 485923 483489 486550 484189
rect 487250 483489 487877 484189
rect 488577 483489 489204 484189
rect 489904 483489 490531 484189
rect 491231 483489 491858 484189
rect 492558 483489 493185 484189
rect 493885 483489 494512 484189
rect 495212 483489 495839 484189
rect 496539 483489 497166 484189
rect 497866 483489 498493 484189
rect 499193 483489 499820 484189
rect 500520 483489 501147 484189
rect 501847 483489 502474 484189
rect 503174 483489 503801 484189
rect 504501 483489 505128 484189
rect 505828 483489 506455 484189
rect 507155 483489 507466 484189
rect 481938 483173 507466 483489
rect 481938 482808 506681 483173
rect 444162 480913 468473 481095
rect 444162 480840 444322 480913
rect 118930 480340 144555 480560
rect 444052 480340 444322 480840
rect 118930 480296 444322 480340
rect 118930 479596 119166 480296
rect 119866 479596 120188 480296
rect 120888 479596 121210 480296
rect 121910 479596 122232 480296
rect 122932 479596 123254 480296
rect 123954 479596 124276 480296
rect 124976 479596 125298 480296
rect 125998 479596 126320 480296
rect 127020 479596 127342 480296
rect 128042 479596 128364 480296
rect 129064 479596 129386 480296
rect 130086 479596 130408 480296
rect 131108 479596 131430 480296
rect 132130 479596 132452 480296
rect 133152 479596 133474 480296
rect 134174 479596 134496 480296
rect 135196 479596 135518 480296
rect 136218 479596 136540 480296
rect 137240 479596 137562 480296
rect 138262 479596 138584 480296
rect 139284 479596 139606 480296
rect 140306 479596 140628 480296
rect 141328 479596 141650 480296
rect 142350 479596 142672 480296
rect 143372 479596 143694 480296
rect 144394 480213 444322 480296
rect 445022 480213 445379 480913
rect 446079 480213 446436 480913
rect 447136 480213 447493 480913
rect 448193 480213 448550 480913
rect 449250 480213 449607 480913
rect 450307 480213 450664 480913
rect 451364 480213 451721 480913
rect 452421 480213 452778 480913
rect 453478 480213 453835 480913
rect 454535 480213 454892 480913
rect 455592 480213 455949 480913
rect 456649 480213 457006 480913
rect 457706 480213 458063 480913
rect 458763 480213 459120 480913
rect 459820 480213 460177 480913
rect 460877 480213 461234 480913
rect 461934 480213 462291 480913
rect 462991 480213 463348 480913
rect 464048 480213 464405 480913
rect 465105 480213 465462 480913
rect 466162 480213 466519 480913
rect 467219 480213 467576 480913
rect 468276 480840 468473 480913
rect 468276 480213 468505 480840
rect 144394 479841 468505 480213
rect 144394 479596 444322 479841
rect 118930 479224 444322 479596
rect 118930 478524 119166 479224
rect 119866 478524 120188 479224
rect 120888 478524 121210 479224
rect 121910 478524 122232 479224
rect 122932 478524 123254 479224
rect 123954 478524 124276 479224
rect 124976 478524 125298 479224
rect 125998 478524 126320 479224
rect 127020 478524 127342 479224
rect 128042 478524 128364 479224
rect 129064 478524 129386 479224
rect 130086 478524 130408 479224
rect 131108 478524 131430 479224
rect 132130 478524 132452 479224
rect 133152 478524 133474 479224
rect 134174 478524 134496 479224
rect 135196 478524 135518 479224
rect 136218 478524 136540 479224
rect 137240 478524 137562 479224
rect 138262 478524 138584 479224
rect 139284 478524 139606 479224
rect 140306 478524 140628 479224
rect 141328 478524 141650 479224
rect 142350 478524 142672 479224
rect 143372 478524 143694 479224
rect 144394 479141 444322 479224
rect 445022 479141 445379 479841
rect 446079 479141 446436 479841
rect 447136 479141 447493 479841
rect 448193 479141 448550 479841
rect 449250 479141 449607 479841
rect 450307 479141 450664 479841
rect 451364 479141 451721 479841
rect 452421 479141 452778 479841
rect 453478 479141 453835 479841
rect 454535 479141 454892 479841
rect 455592 479141 455949 479841
rect 456649 479141 457006 479841
rect 457706 479141 458063 479841
rect 458763 479141 459120 479841
rect 459820 479141 460177 479841
rect 460877 479141 461234 479841
rect 461934 479141 462291 479841
rect 462991 479141 463348 479841
rect 464048 479141 464405 479841
rect 465105 479141 465462 479841
rect 466162 479141 466519 479841
rect 467219 479141 467576 479841
rect 468276 479141 468505 479841
rect 144394 478769 468505 479141
rect 144394 478524 444322 478769
rect 118930 478152 444322 478524
rect 118930 477452 119166 478152
rect 119866 477452 120188 478152
rect 120888 477452 121210 478152
rect 121910 477452 122232 478152
rect 122932 477452 123254 478152
rect 123954 477452 124276 478152
rect 124976 477452 125298 478152
rect 125998 477452 126320 478152
rect 127020 477452 127342 478152
rect 128042 477452 128364 478152
rect 129064 477452 129386 478152
rect 130086 477452 130408 478152
rect 131108 477452 131430 478152
rect 132130 477452 132452 478152
rect 133152 477452 133474 478152
rect 134174 477452 134496 478152
rect 135196 477452 135518 478152
rect 136218 477452 136540 478152
rect 137240 477452 137562 478152
rect 138262 477452 138584 478152
rect 139284 477452 139606 478152
rect 140306 477452 140628 478152
rect 141328 477452 141650 478152
rect 142350 477452 142672 478152
rect 143372 477452 143694 478152
rect 144394 478069 444322 478152
rect 445022 478069 445379 478769
rect 446079 478069 446436 478769
rect 447136 478069 447493 478769
rect 448193 478069 448550 478769
rect 449250 478069 449607 478769
rect 450307 478069 450664 478769
rect 451364 478069 451721 478769
rect 452421 478069 452778 478769
rect 453478 478069 453835 478769
rect 454535 478069 454892 478769
rect 455592 478069 455949 478769
rect 456649 478069 457006 478769
rect 457706 478069 458063 478769
rect 458763 478069 459120 478769
rect 459820 478069 460177 478769
rect 460877 478069 461234 478769
rect 461934 478069 462291 478769
rect 462991 478069 463348 478769
rect 464048 478069 464405 478769
rect 465105 478069 465462 478769
rect 466162 478069 466519 478769
rect 467219 478069 467576 478769
rect 468276 478069 468505 478769
rect 144394 477697 468505 478069
rect 144394 477452 444322 477697
rect 118930 477080 444322 477452
rect 118930 476380 119166 477080
rect 119866 476380 120188 477080
rect 120888 476380 121210 477080
rect 121910 476380 122232 477080
rect 122932 476380 123254 477080
rect 123954 476380 124276 477080
rect 124976 476380 125298 477080
rect 125998 476380 126320 477080
rect 127020 476380 127342 477080
rect 128042 476380 128364 477080
rect 129064 476380 129386 477080
rect 130086 476380 130408 477080
rect 131108 476380 131430 477080
rect 132130 476380 132452 477080
rect 133152 476380 133474 477080
rect 134174 476380 134496 477080
rect 135196 476380 135518 477080
rect 136218 476380 136540 477080
rect 137240 476380 137562 477080
rect 138262 476380 138584 477080
rect 139284 476380 139606 477080
rect 140306 476380 140628 477080
rect 141328 476380 141650 477080
rect 142350 476380 142672 477080
rect 143372 476380 143694 477080
rect 144394 476997 444322 477080
rect 445022 476997 445379 477697
rect 446079 476997 446436 477697
rect 447136 476997 447493 477697
rect 448193 476997 448550 477697
rect 449250 476997 449607 477697
rect 450307 476997 450664 477697
rect 451364 476997 451721 477697
rect 452421 476997 452778 477697
rect 453478 476997 453835 477697
rect 454535 476997 454892 477697
rect 455592 476997 455949 477697
rect 456649 476997 457006 477697
rect 457706 476997 458063 477697
rect 458763 476997 459120 477697
rect 459820 476997 460177 477697
rect 460877 476997 461234 477697
rect 461934 476997 462291 477697
rect 462991 476997 463348 477697
rect 464048 476997 464405 477697
rect 465105 476997 465462 477697
rect 466162 476997 466519 477697
rect 467219 476997 467576 477697
rect 468276 476997 468505 477697
rect 144394 476625 468505 476997
rect 144394 476380 444322 476625
rect 118930 476008 444322 476380
rect 118930 475308 119166 476008
rect 119866 475308 120188 476008
rect 120888 475308 121210 476008
rect 121910 475308 122232 476008
rect 122932 475308 123254 476008
rect 123954 475308 124276 476008
rect 124976 475308 125298 476008
rect 125998 475308 126320 476008
rect 127020 475308 127342 476008
rect 128042 475308 128364 476008
rect 129064 475308 129386 476008
rect 130086 475308 130408 476008
rect 131108 475308 131430 476008
rect 132130 475308 132452 476008
rect 133152 475308 133474 476008
rect 134174 475308 134496 476008
rect 135196 475308 135518 476008
rect 136218 475308 136540 476008
rect 137240 475308 137562 476008
rect 138262 475308 138584 476008
rect 139284 475308 139606 476008
rect 140306 475308 140628 476008
rect 141328 475308 141650 476008
rect 142350 475308 142672 476008
rect 143372 475308 143694 476008
rect 144394 475925 444322 476008
rect 445022 475925 445379 476625
rect 446079 475925 446436 476625
rect 447136 475925 447493 476625
rect 448193 475925 448550 476625
rect 449250 475925 449607 476625
rect 450307 475925 450664 476625
rect 451364 475925 451721 476625
rect 452421 475925 452778 476625
rect 453478 475925 453835 476625
rect 454535 475925 454892 476625
rect 455592 475925 455949 476625
rect 456649 475925 457006 476625
rect 457706 475925 458063 476625
rect 458763 475925 459120 476625
rect 459820 475925 460177 476625
rect 460877 475925 461234 476625
rect 461934 475925 462291 476625
rect 462991 475925 463348 476625
rect 464048 475925 464405 476625
rect 465105 475925 465462 476625
rect 466162 475925 466519 476625
rect 467219 475925 467576 476625
rect 468276 475925 468505 476625
rect 144394 475553 468505 475925
rect 144394 475308 444322 475553
rect 118930 474936 444322 475308
rect 118930 474236 119166 474936
rect 119866 474236 120188 474936
rect 120888 474236 121210 474936
rect 121910 474236 122232 474936
rect 122932 474236 123254 474936
rect 123954 474236 124276 474936
rect 124976 474236 125298 474936
rect 125998 474236 126320 474936
rect 127020 474236 127342 474936
rect 128042 474236 128364 474936
rect 129064 474236 129386 474936
rect 130086 474236 130408 474936
rect 131108 474236 131430 474936
rect 132130 474236 132452 474936
rect 133152 474236 133474 474936
rect 134174 474236 134496 474936
rect 135196 474236 135518 474936
rect 136218 474236 136540 474936
rect 137240 474236 137562 474936
rect 138262 474236 138584 474936
rect 139284 474236 139606 474936
rect 140306 474236 140628 474936
rect 141328 474236 141650 474936
rect 142350 474236 142672 474936
rect 143372 474236 143694 474936
rect 144394 474853 444322 474936
rect 445022 474853 445379 475553
rect 446079 474853 446436 475553
rect 447136 474853 447493 475553
rect 448193 474853 448550 475553
rect 449250 474853 449607 475553
rect 450307 474853 450664 475553
rect 451364 474853 451721 475553
rect 452421 474853 452778 475553
rect 453478 474853 453835 475553
rect 454535 474853 454892 475553
rect 455592 474853 455949 475553
rect 456649 474853 457006 475553
rect 457706 474853 458063 475553
rect 458763 474853 459120 475553
rect 459820 474853 460177 475553
rect 460877 474853 461234 475553
rect 461934 474853 462291 475553
rect 462991 474853 463348 475553
rect 464048 474853 464405 475553
rect 465105 474853 465462 475553
rect 466162 474853 466519 475553
rect 467219 474853 467576 475553
rect 468276 474853 468505 475553
rect 144394 474481 468505 474853
rect 144394 474236 444322 474481
rect 118930 473864 444322 474236
rect 118930 473164 119166 473864
rect 119866 473164 120188 473864
rect 120888 473164 121210 473864
rect 121910 473164 122232 473864
rect 122932 473164 123254 473864
rect 123954 473164 124276 473864
rect 124976 473164 125298 473864
rect 125998 473164 126320 473864
rect 127020 473164 127342 473864
rect 128042 473164 128364 473864
rect 129064 473164 129386 473864
rect 130086 473164 130408 473864
rect 131108 473164 131430 473864
rect 132130 473164 132452 473864
rect 133152 473164 133474 473864
rect 134174 473164 134496 473864
rect 135196 473164 135518 473864
rect 136218 473164 136540 473864
rect 137240 473164 137562 473864
rect 138262 473164 138584 473864
rect 139284 473164 139606 473864
rect 140306 473164 140628 473864
rect 141328 473164 141650 473864
rect 142350 473164 142672 473864
rect 143372 473164 143694 473864
rect 144394 473781 444322 473864
rect 445022 473781 445379 474481
rect 446079 473781 446436 474481
rect 447136 473781 447493 474481
rect 448193 473781 448550 474481
rect 449250 473781 449607 474481
rect 450307 473781 450664 474481
rect 451364 473781 451721 474481
rect 452421 473781 452778 474481
rect 453478 473781 453835 474481
rect 454535 473781 454892 474481
rect 455592 473781 455949 474481
rect 456649 473781 457006 474481
rect 457706 473781 458063 474481
rect 458763 473781 459120 474481
rect 459820 473781 460177 474481
rect 460877 473781 461234 474481
rect 461934 473781 462291 474481
rect 462991 473781 463348 474481
rect 464048 473781 464405 474481
rect 465105 473781 465462 474481
rect 466162 473781 466519 474481
rect 467219 473781 467576 474481
rect 468276 473781 468505 474481
rect 144394 473409 468505 473781
rect 144394 473164 444322 473409
rect 118930 472792 444322 473164
rect 118930 472092 119166 472792
rect 119866 472092 120188 472792
rect 120888 472092 121210 472792
rect 121910 472092 122232 472792
rect 122932 472092 123254 472792
rect 123954 472092 124276 472792
rect 124976 472092 125298 472792
rect 125998 472092 126320 472792
rect 127020 472092 127342 472792
rect 128042 472092 128364 472792
rect 129064 472092 129386 472792
rect 130086 472092 130408 472792
rect 131108 472092 131430 472792
rect 132130 472092 132452 472792
rect 133152 472092 133474 472792
rect 134174 472092 134496 472792
rect 135196 472092 135518 472792
rect 136218 472092 136540 472792
rect 137240 472092 137562 472792
rect 138262 472092 138584 472792
rect 139284 472092 139606 472792
rect 140306 472092 140628 472792
rect 141328 472092 141650 472792
rect 142350 472092 142672 472792
rect 143372 472092 143694 472792
rect 144394 472709 444322 472792
rect 445022 472709 445379 473409
rect 446079 472709 446436 473409
rect 447136 472709 447493 473409
rect 448193 472709 448550 473409
rect 449250 472709 449607 473409
rect 450307 472709 450664 473409
rect 451364 472709 451721 473409
rect 452421 472709 452778 473409
rect 453478 472709 453835 473409
rect 454535 472709 454892 473409
rect 455592 472709 455949 473409
rect 456649 472709 457006 473409
rect 457706 472709 458063 473409
rect 458763 472709 459120 473409
rect 459820 472709 460177 473409
rect 460877 472709 461234 473409
rect 461934 472709 462291 473409
rect 462991 472709 463348 473409
rect 464048 472709 464405 473409
rect 465105 472709 465462 473409
rect 466162 472709 466519 473409
rect 467219 472709 467576 473409
rect 468276 472709 468505 473409
rect 144394 472337 468505 472709
rect 144394 472092 444322 472337
rect 118930 471720 444322 472092
rect 118930 471020 119166 471720
rect 119866 471020 120188 471720
rect 120888 471020 121210 471720
rect 121910 471020 122232 471720
rect 122932 471020 123254 471720
rect 123954 471020 124276 471720
rect 124976 471020 125298 471720
rect 125998 471020 126320 471720
rect 127020 471020 127342 471720
rect 128042 471020 128364 471720
rect 129064 471020 129386 471720
rect 130086 471020 130408 471720
rect 131108 471020 131430 471720
rect 132130 471020 132452 471720
rect 133152 471020 133474 471720
rect 134174 471020 134496 471720
rect 135196 471020 135518 471720
rect 136218 471020 136540 471720
rect 137240 471020 137562 471720
rect 138262 471020 138584 471720
rect 139284 471020 139606 471720
rect 140306 471020 140628 471720
rect 141328 471020 141650 471720
rect 142350 471020 142672 471720
rect 143372 471020 143694 471720
rect 144394 471637 444322 471720
rect 445022 471637 445379 472337
rect 446079 471637 446436 472337
rect 447136 471637 447493 472337
rect 448193 471637 448550 472337
rect 449250 471637 449607 472337
rect 450307 471637 450664 472337
rect 451364 471637 451721 472337
rect 452421 471637 452778 472337
rect 453478 471637 453835 472337
rect 454535 471637 454892 472337
rect 455592 471637 455949 472337
rect 456649 471637 457006 472337
rect 457706 471637 458063 472337
rect 458763 471637 459120 472337
rect 459820 471637 460177 472337
rect 460877 471637 461234 472337
rect 461934 471637 462291 472337
rect 462991 471637 463348 472337
rect 464048 471637 464405 472337
rect 465105 471637 465462 472337
rect 466162 471637 466519 472337
rect 467219 471637 467576 472337
rect 468276 471637 468505 472337
rect 144394 471265 468505 471637
rect 144394 471020 444322 471265
rect 118930 470648 444322 471020
rect 118930 469948 119166 470648
rect 119866 469948 120188 470648
rect 120888 469948 121210 470648
rect 121910 469948 122232 470648
rect 122932 469948 123254 470648
rect 123954 469948 124276 470648
rect 124976 469948 125298 470648
rect 125998 469948 126320 470648
rect 127020 469948 127342 470648
rect 128042 469948 128364 470648
rect 129064 469948 129386 470648
rect 130086 469948 130408 470648
rect 131108 469948 131430 470648
rect 132130 469948 132452 470648
rect 133152 469948 133474 470648
rect 134174 469948 134496 470648
rect 135196 469948 135518 470648
rect 136218 469948 136540 470648
rect 137240 469948 137562 470648
rect 138262 469948 138584 470648
rect 139284 469948 139606 470648
rect 140306 469948 140628 470648
rect 141328 469948 141650 470648
rect 142350 469948 142672 470648
rect 143372 469948 143694 470648
rect 144394 470565 444322 470648
rect 445022 470565 445379 471265
rect 446079 470565 446436 471265
rect 447136 470565 447493 471265
rect 448193 470565 448550 471265
rect 449250 470565 449607 471265
rect 450307 470565 450664 471265
rect 451364 470565 451721 471265
rect 452421 470565 452778 471265
rect 453478 470565 453835 471265
rect 454535 470565 454892 471265
rect 455592 470565 455949 471265
rect 456649 470565 457006 471265
rect 457706 470565 458063 471265
rect 458763 470565 459120 471265
rect 459820 470565 460177 471265
rect 460877 470565 461234 471265
rect 461934 470565 462291 471265
rect 462991 470565 463348 471265
rect 464048 470565 464405 471265
rect 465105 470565 465462 471265
rect 466162 470565 466519 471265
rect 467219 470565 467576 471265
rect 468276 470565 468505 471265
rect 144394 470193 468505 470565
rect 144394 469948 444322 470193
rect 118930 469576 444322 469948
rect 118930 468876 119166 469576
rect 119866 468876 120188 469576
rect 120888 468876 121210 469576
rect 121910 468876 122232 469576
rect 122932 468876 123254 469576
rect 123954 468876 124276 469576
rect 124976 468876 125298 469576
rect 125998 468876 126320 469576
rect 127020 468876 127342 469576
rect 128042 468876 128364 469576
rect 129064 468876 129386 469576
rect 130086 468876 130408 469576
rect 131108 468876 131430 469576
rect 132130 468876 132452 469576
rect 133152 468876 133474 469576
rect 134174 468876 134496 469576
rect 135196 468876 135518 469576
rect 136218 468876 136540 469576
rect 137240 468876 137562 469576
rect 138262 468876 138584 469576
rect 139284 468876 139606 469576
rect 140306 468876 140628 469576
rect 141328 468876 141650 469576
rect 142350 468876 142672 469576
rect 143372 468876 143694 469576
rect 144394 469493 444322 469576
rect 445022 469493 445379 470193
rect 446079 469493 446436 470193
rect 447136 469493 447493 470193
rect 448193 469493 448550 470193
rect 449250 469493 449607 470193
rect 450307 469493 450664 470193
rect 451364 469493 451721 470193
rect 452421 469493 452778 470193
rect 453478 469493 453835 470193
rect 454535 469493 454892 470193
rect 455592 469493 455949 470193
rect 456649 469493 457006 470193
rect 457706 469493 458063 470193
rect 458763 469493 459120 470193
rect 459820 469493 460177 470193
rect 460877 469493 461234 470193
rect 461934 469493 462291 470193
rect 462991 469493 463348 470193
rect 464048 469493 464405 470193
rect 465105 469493 465462 470193
rect 466162 469493 466519 470193
rect 467219 469493 467576 470193
rect 468276 469493 468505 470193
rect 144394 469121 468505 469493
rect 144394 468876 444322 469121
rect 118930 468504 444322 468876
rect 90963 467581 97688 468097
rect 90963 467431 91879 467581
rect 92029 467431 92147 467581
rect 92297 467431 92415 467581
rect 92565 467431 92683 467581
rect 92833 467431 92951 467581
rect 93101 467431 93219 467581
rect 93369 467431 93487 467581
rect 93637 467431 93755 467581
rect 93905 467431 94023 467581
rect 94173 467431 94291 467581
rect 94441 467431 97688 467581
rect 90963 467343 97688 467431
rect 90963 467193 91879 467343
rect 92029 467193 92147 467343
rect 92297 467193 92415 467343
rect 92565 467193 92683 467343
rect 92833 467193 92951 467343
rect 93101 467193 93219 467343
rect 93369 467193 93487 467343
rect 93637 467193 93755 467343
rect 93905 467193 94023 467343
rect 94173 467193 94291 467343
rect 94441 467193 97688 467343
rect 90963 467105 97688 467193
rect 90963 466955 91879 467105
rect 92029 466955 92147 467105
rect 92297 466955 92415 467105
rect 92565 466955 92683 467105
rect 92833 466955 92951 467105
rect 93101 466955 93219 467105
rect 93369 466955 93487 467105
rect 93637 466955 93755 467105
rect 93905 466955 94023 467105
rect 94173 466955 94291 467105
rect 94441 466955 97688 467105
rect 90963 466867 97688 466955
rect 90963 466717 91879 466867
rect 92029 466717 92147 466867
rect 92297 466717 92415 466867
rect 92565 466717 92683 466867
rect 92833 466717 92951 466867
rect 93101 466717 93219 466867
rect 93369 466717 93487 466867
rect 93637 466717 93755 466867
rect 93905 466717 94023 466867
rect 94173 466717 94291 466867
rect 94441 466717 97688 466867
rect 90963 466632 97688 466717
rect 85125 466629 97688 466632
rect 85125 466479 91879 466629
rect 92029 466479 92147 466629
rect 92297 466479 92415 466629
rect 92565 466479 92683 466629
rect 92833 466479 92951 466629
rect 93101 466479 93219 466629
rect 93369 466479 93487 466629
rect 93637 466479 93755 466629
rect 93905 466479 94023 466629
rect 94173 466479 94291 466629
rect 94441 466479 97688 466629
rect 85125 466391 97688 466479
rect 85125 466241 91879 466391
rect 92029 466241 92147 466391
rect 92297 466241 92415 466391
rect 92565 466241 92683 466391
rect 92833 466241 92951 466391
rect 93101 466241 93219 466391
rect 93369 466241 93487 466391
rect 93637 466241 93755 466391
rect 93905 466241 94023 466391
rect 94173 466241 94291 466391
rect 94441 466241 97688 466391
rect 85125 466153 97688 466241
rect 85125 466003 91879 466153
rect 92029 466003 92147 466153
rect 92297 466003 92415 466153
rect 92565 466003 92683 466153
rect 92833 466003 92951 466153
rect 93101 466003 93219 466153
rect 93369 466003 93487 466153
rect 93637 466003 93755 466153
rect 93905 466003 94023 466153
rect 94173 466003 94291 466153
rect 94441 466003 97688 466153
rect 85125 465915 97688 466003
rect 85125 465765 91879 465915
rect 92029 465765 92147 465915
rect 92297 465765 92415 465915
rect 92565 465765 92683 465915
rect 92833 465765 92951 465915
rect 93101 465765 93219 465915
rect 93369 465765 93487 465915
rect 93637 465765 93755 465915
rect 93905 465765 94023 465915
rect 94173 465765 94291 465915
rect 94441 465765 97688 465915
rect 85125 465677 97688 465765
rect 85125 465527 91879 465677
rect 92029 465527 92147 465677
rect 92297 465527 92415 465677
rect 92565 465527 92683 465677
rect 92833 465527 92951 465677
rect 93101 465527 93219 465677
rect 93369 465527 93487 465677
rect 93637 465527 93755 465677
rect 93905 465527 94023 465677
rect 94173 465527 94291 465677
rect 94441 465527 97688 465677
rect 85125 465439 97688 465527
rect 85125 465411 91879 465439
rect 77870 453525 78295 453564
rect 77870 453392 77983 453525
rect 78116 453392 78295 453525
rect 77870 453288 78295 453392
rect 85125 453288 86346 465411
rect 90963 465289 91879 465411
rect 92029 465289 92147 465439
rect 92297 465289 92415 465439
rect 92565 465289 92683 465439
rect 92833 465289 92951 465439
rect 93101 465289 93219 465439
rect 93369 465289 93487 465439
rect 93637 465289 93755 465439
rect 93905 465289 94023 465439
rect 94173 465289 94291 465439
rect 94441 465289 97688 465439
rect 90963 464614 97688 465289
rect 118930 467804 119166 468504
rect 119866 467804 120188 468504
rect 120888 467804 121210 468504
rect 121910 467804 122232 468504
rect 122932 467804 123254 468504
rect 123954 467804 124276 468504
rect 124976 467804 125298 468504
rect 125998 467804 126320 468504
rect 127020 467804 127342 468504
rect 128042 467804 128364 468504
rect 129064 467804 129386 468504
rect 130086 467804 130408 468504
rect 131108 467804 131430 468504
rect 132130 467804 132452 468504
rect 133152 467804 133474 468504
rect 134174 467804 134496 468504
rect 135196 467804 135518 468504
rect 136218 467804 136540 468504
rect 137240 467804 137562 468504
rect 138262 467804 138584 468504
rect 139284 467804 139606 468504
rect 140306 467804 140628 468504
rect 141328 467804 141650 468504
rect 142350 467804 142672 468504
rect 143372 467804 143694 468504
rect 144394 468421 444322 468504
rect 445022 468421 445379 469121
rect 446079 468421 446436 469121
rect 447136 468421 447493 469121
rect 448193 468421 448550 469121
rect 449250 468421 449607 469121
rect 450307 468421 450664 469121
rect 451364 468421 451721 469121
rect 452421 468421 452778 469121
rect 453478 468421 453835 469121
rect 454535 468421 454892 469121
rect 455592 468421 455949 469121
rect 456649 468421 457006 469121
rect 457706 468421 458063 469121
rect 458763 468421 459120 469121
rect 459820 468421 460177 469121
rect 460877 468421 461234 469121
rect 461934 468421 462291 469121
rect 462991 468421 463348 469121
rect 464048 468421 464405 469121
rect 465105 468421 465462 469121
rect 466162 468421 466519 469121
rect 467219 468421 467576 469121
rect 468276 468421 468505 469121
rect 144394 468049 468505 468421
rect 144394 467804 444322 468049
rect 118930 467432 444322 467804
rect 118930 466732 119166 467432
rect 119866 466732 120188 467432
rect 120888 466732 121210 467432
rect 121910 466732 122232 467432
rect 122932 466732 123254 467432
rect 123954 466732 124276 467432
rect 124976 466732 125298 467432
rect 125998 466732 126320 467432
rect 127020 466732 127342 467432
rect 128042 466732 128364 467432
rect 129064 466732 129386 467432
rect 130086 466732 130408 467432
rect 131108 466732 131430 467432
rect 132130 466732 132452 467432
rect 133152 466732 133474 467432
rect 134174 466732 134496 467432
rect 135196 466732 135518 467432
rect 136218 466732 136540 467432
rect 137240 466732 137562 467432
rect 138262 466732 138584 467432
rect 139284 466732 139606 467432
rect 140306 466732 140628 467432
rect 141328 466732 141650 467432
rect 142350 466732 142672 467432
rect 143372 466732 143694 467432
rect 144394 467349 444322 467432
rect 445022 467349 445379 468049
rect 446079 467349 446436 468049
rect 447136 467349 447493 468049
rect 448193 467349 448550 468049
rect 449250 467349 449607 468049
rect 450307 467349 450664 468049
rect 451364 467349 451721 468049
rect 452421 467349 452778 468049
rect 453478 467349 453835 468049
rect 454535 467349 454892 468049
rect 455592 467349 455949 468049
rect 456649 467349 457006 468049
rect 457706 467349 458063 468049
rect 458763 467349 459120 468049
rect 459820 467349 460177 468049
rect 460877 467349 461234 468049
rect 461934 467349 462291 468049
rect 462991 467349 463348 468049
rect 464048 467349 464405 468049
rect 465105 467349 465462 468049
rect 466162 467349 466519 468049
rect 467219 467349 467576 468049
rect 468276 467349 468505 468049
rect 144394 466977 468505 467349
rect 144394 466732 444322 466977
rect 118930 466360 444322 466732
rect 118930 465660 119166 466360
rect 119866 465660 120188 466360
rect 120888 465660 121210 466360
rect 121910 465660 122232 466360
rect 122932 465660 123254 466360
rect 123954 465660 124276 466360
rect 124976 465660 125298 466360
rect 125998 465660 126320 466360
rect 127020 465660 127342 466360
rect 128042 465660 128364 466360
rect 129064 465660 129386 466360
rect 130086 465660 130408 466360
rect 131108 465660 131430 466360
rect 132130 465660 132452 466360
rect 133152 465660 133474 466360
rect 134174 465660 134496 466360
rect 135196 465660 135518 466360
rect 136218 465660 136540 466360
rect 137240 465660 137562 466360
rect 138262 465660 138584 466360
rect 139284 465660 139606 466360
rect 140306 465660 140628 466360
rect 141328 465660 141650 466360
rect 142350 465660 142672 466360
rect 143372 465660 143694 466360
rect 144394 466277 444322 466360
rect 445022 466277 445379 466977
rect 446079 466277 446436 466977
rect 447136 466277 447493 466977
rect 448193 466277 448550 466977
rect 449250 466277 449607 466977
rect 450307 466277 450664 466977
rect 451364 466277 451721 466977
rect 452421 466277 452778 466977
rect 453478 466277 453835 466977
rect 454535 466277 454892 466977
rect 455592 466277 455949 466977
rect 456649 466277 457006 466977
rect 457706 466277 458063 466977
rect 458763 466277 459120 466977
rect 459820 466277 460177 466977
rect 460877 466277 461234 466977
rect 461934 466277 462291 466977
rect 462991 466277 463348 466977
rect 464048 466277 464405 466977
rect 465105 466277 465462 466977
rect 466162 466277 466519 466977
rect 467219 466277 467576 466977
rect 468276 466277 468505 466977
rect 144394 465905 468505 466277
rect 144394 465660 444322 465905
rect 118930 465288 444322 465660
rect 118930 464588 119166 465288
rect 119866 464588 120188 465288
rect 120888 464588 121210 465288
rect 121910 464588 122232 465288
rect 122932 464588 123254 465288
rect 123954 464588 124276 465288
rect 124976 464588 125298 465288
rect 125998 464588 126320 465288
rect 127020 464588 127342 465288
rect 128042 464588 128364 465288
rect 129064 464588 129386 465288
rect 130086 464588 130408 465288
rect 131108 464588 131430 465288
rect 132130 464588 132452 465288
rect 133152 464588 133474 465288
rect 134174 464588 134496 465288
rect 135196 464588 135518 465288
rect 136218 464588 136540 465288
rect 137240 464588 137562 465288
rect 138262 464588 138584 465288
rect 139284 464588 139606 465288
rect 140306 464588 140628 465288
rect 141328 464588 141650 465288
rect 142350 464588 142672 465288
rect 143372 464588 143694 465288
rect 144394 465205 444322 465288
rect 445022 465205 445379 465905
rect 446079 465205 446436 465905
rect 447136 465205 447493 465905
rect 448193 465205 448550 465905
rect 449250 465205 449607 465905
rect 450307 465205 450664 465905
rect 451364 465205 451721 465905
rect 452421 465205 452778 465905
rect 453478 465205 453835 465905
rect 454535 465205 454892 465905
rect 455592 465205 455949 465905
rect 456649 465205 457006 465905
rect 457706 465205 458063 465905
rect 458763 465205 459120 465905
rect 459820 465205 460177 465905
rect 460877 465205 461234 465905
rect 461934 465205 462291 465905
rect 462991 465205 463348 465905
rect 464048 465205 464405 465905
rect 465105 465205 465462 465905
rect 466162 465205 466519 465905
rect 467219 465205 467576 465905
rect 468276 465205 468505 465905
rect 144394 464833 468505 465205
rect 144394 464588 444322 464833
rect 118930 464216 444322 464588
rect 118930 463516 119166 464216
rect 119866 463516 120188 464216
rect 120888 463516 121210 464216
rect 121910 463516 122232 464216
rect 122932 463516 123254 464216
rect 123954 463516 124276 464216
rect 124976 463516 125298 464216
rect 125998 463516 126320 464216
rect 127020 463516 127342 464216
rect 128042 463516 128364 464216
rect 129064 463516 129386 464216
rect 130086 463516 130408 464216
rect 131108 463516 131430 464216
rect 132130 463516 132452 464216
rect 133152 463516 133474 464216
rect 134174 463516 134496 464216
rect 135196 463516 135518 464216
rect 136218 463516 136540 464216
rect 137240 463516 137562 464216
rect 138262 463516 138584 464216
rect 139284 463516 139606 464216
rect 140306 463516 140628 464216
rect 141328 463516 141650 464216
rect 142350 463516 142672 464216
rect 143372 463516 143694 464216
rect 144394 464133 444322 464216
rect 445022 464133 445379 464833
rect 446079 464133 446436 464833
rect 447136 464133 447493 464833
rect 448193 464133 448550 464833
rect 449250 464133 449607 464833
rect 450307 464133 450664 464833
rect 451364 464133 451721 464833
rect 452421 464133 452778 464833
rect 453478 464133 453835 464833
rect 454535 464133 454892 464833
rect 455592 464133 455949 464833
rect 456649 464133 457006 464833
rect 457706 464133 458063 464833
rect 458763 464133 459120 464833
rect 459820 464133 460177 464833
rect 460877 464133 461234 464833
rect 461934 464133 462291 464833
rect 462991 464133 463348 464833
rect 464048 464133 464405 464833
rect 465105 464133 465462 464833
rect 466162 464133 466519 464833
rect 467219 464133 467576 464833
rect 468276 464133 468505 464833
rect 144394 463761 468505 464133
rect 144394 463516 444322 463761
rect 118930 463399 444322 463516
rect 118930 463144 144555 463399
rect 118930 462444 119166 463144
rect 119866 462444 120188 463144
rect 120888 462444 121210 463144
rect 121910 462444 122232 463144
rect 122932 462444 123254 463144
rect 123954 462444 124276 463144
rect 124976 462444 125298 463144
rect 125998 462444 126320 463144
rect 127020 462444 127342 463144
rect 128042 462444 128364 463144
rect 129064 462444 129386 463144
rect 130086 462444 130408 463144
rect 131108 462444 131430 463144
rect 132130 462444 132452 463144
rect 133152 462444 133474 463144
rect 134174 462444 134496 463144
rect 135196 462444 135518 463144
rect 136218 462444 136540 463144
rect 137240 462444 137562 463144
rect 138262 462444 138584 463144
rect 139284 462444 139606 463144
rect 140306 462444 140628 463144
rect 141328 462444 141650 463144
rect 142350 462444 142672 463144
rect 143372 462444 143694 463144
rect 144394 462444 144555 463144
rect 118930 462072 144555 462444
rect 118930 461372 119166 462072
rect 119866 461372 120188 462072
rect 120888 461372 121210 462072
rect 121910 461372 122232 462072
rect 122932 461372 123254 462072
rect 123954 461372 124276 462072
rect 124976 461372 125298 462072
rect 125998 461372 126320 462072
rect 127020 461372 127342 462072
rect 128042 461372 128364 462072
rect 129064 461372 129386 462072
rect 130086 461372 130408 462072
rect 131108 461372 131430 462072
rect 132130 461372 132452 462072
rect 133152 461372 133474 462072
rect 134174 461372 134496 462072
rect 135196 461372 135518 462072
rect 136218 461372 136540 462072
rect 137240 461372 137562 462072
rect 138262 461372 138584 462072
rect 139284 461372 139606 462072
rect 140306 461372 140628 462072
rect 141328 461372 141650 462072
rect 142350 461372 142672 462072
rect 143372 461372 143694 462072
rect 144394 461372 144555 462072
rect 118930 461000 144555 461372
rect 118930 460300 119166 461000
rect 119866 460300 120188 461000
rect 120888 460300 121210 461000
rect 121910 460300 122232 461000
rect 122932 460300 123254 461000
rect 123954 460300 124276 461000
rect 124976 460300 125298 461000
rect 125998 460300 126320 461000
rect 127020 460300 127342 461000
rect 128042 460300 128364 461000
rect 129064 460300 129386 461000
rect 130086 460300 130408 461000
rect 131108 460300 131430 461000
rect 132130 460300 132452 461000
rect 133152 460300 133474 461000
rect 134174 460300 134496 461000
rect 135196 460300 135518 461000
rect 136218 460300 136540 461000
rect 137240 460300 137562 461000
rect 138262 460300 138584 461000
rect 139284 460300 139606 461000
rect 140306 460300 140628 461000
rect 141328 460300 141650 461000
rect 142350 460300 142672 461000
rect 143372 460300 143694 461000
rect 144394 460300 144555 461000
rect 118930 459928 144555 460300
rect 118930 459228 119166 459928
rect 119866 459228 120188 459928
rect 120888 459228 121210 459928
rect 121910 459228 122232 459928
rect 122932 459228 123254 459928
rect 123954 459228 124276 459928
rect 124976 459228 125298 459928
rect 125998 459228 126320 459928
rect 127020 459228 127342 459928
rect 128042 459228 128364 459928
rect 129064 459228 129386 459928
rect 130086 459228 130408 459928
rect 131108 459228 131430 459928
rect 132130 459228 132452 459928
rect 133152 459228 133474 459928
rect 134174 459228 134496 459928
rect 135196 459228 135518 459928
rect 136218 459228 136540 459928
rect 137240 459228 137562 459928
rect 138262 459228 138584 459928
rect 139284 459228 139606 459928
rect 140306 459228 140628 459928
rect 141328 459228 141650 459928
rect 142350 459228 142672 459928
rect 143372 459228 143694 459928
rect 144394 459228 144555 459928
rect 118930 459077 144555 459228
rect 444052 463061 444322 463399
rect 445022 463061 445379 463761
rect 446079 463061 446436 463761
rect 447136 463061 447493 463761
rect 448193 463061 448550 463761
rect 449250 463061 449607 463761
rect 450307 463061 450664 463761
rect 451364 463061 451721 463761
rect 452421 463061 452778 463761
rect 453478 463061 453835 463761
rect 454535 463061 454892 463761
rect 455592 463061 455949 463761
rect 456649 463061 457006 463761
rect 457706 463061 458063 463761
rect 458763 463061 459120 463761
rect 459820 463061 460177 463761
rect 460877 463061 461234 463761
rect 461934 463061 462291 463761
rect 462991 463061 463348 463761
rect 464048 463061 464405 463761
rect 465105 463061 465462 463761
rect 466162 463061 466519 463761
rect 467219 463061 467576 463761
rect 468276 463061 468505 463761
rect 444052 462689 468505 463061
rect 444052 461989 444322 462689
rect 445022 461989 445379 462689
rect 446079 461989 446436 462689
rect 447136 461989 447493 462689
rect 448193 461989 448550 462689
rect 449250 461989 449607 462689
rect 450307 461989 450664 462689
rect 451364 461989 451721 462689
rect 452421 461989 452778 462689
rect 453478 461989 453835 462689
rect 454535 461989 454892 462689
rect 455592 461989 455949 462689
rect 456649 461989 457006 462689
rect 457706 461989 458063 462689
rect 458763 461989 459120 462689
rect 459820 461989 460177 462689
rect 460877 461989 461234 462689
rect 461934 461989 462291 462689
rect 462991 461989 463348 462689
rect 464048 461989 464405 462689
rect 465105 461989 465462 462689
rect 466162 461989 466519 462689
rect 467219 461989 467576 462689
rect 468276 461989 468505 462689
rect 444052 461617 468505 461989
rect 444052 460917 444322 461617
rect 445022 460917 445379 461617
rect 446079 460917 446436 461617
rect 447136 460917 447493 461617
rect 448193 460917 448550 461617
rect 449250 460917 449607 461617
rect 450307 460917 450664 461617
rect 451364 460917 451721 461617
rect 452421 460917 452778 461617
rect 453478 460917 453835 461617
rect 454535 460917 454892 461617
rect 455592 460917 455949 461617
rect 456649 460917 457006 461617
rect 457706 460917 458063 461617
rect 458763 460917 459120 461617
rect 459820 460917 460177 461617
rect 460877 460917 461234 461617
rect 461934 460917 462291 461617
rect 462991 460917 463348 461617
rect 464048 460917 464405 461617
rect 465105 460917 465462 461617
rect 466162 460917 466519 461617
rect 467219 460917 467576 461617
rect 468276 460917 468505 461617
rect 444052 460545 468505 460917
rect 444052 459845 444322 460545
rect 445022 459845 445379 460545
rect 446079 459845 446436 460545
rect 447136 459845 447493 460545
rect 448193 459845 448550 460545
rect 449250 459845 449607 460545
rect 450307 459845 450664 460545
rect 451364 459845 451721 460545
rect 452421 459845 452778 460545
rect 453478 459845 453835 460545
rect 454535 459845 454892 460545
rect 455592 459845 455949 460545
rect 456649 459845 457006 460545
rect 457706 459845 458063 460545
rect 458763 459845 459120 460545
rect 459820 459845 460177 460545
rect 460877 459845 461234 460545
rect 461934 459845 462291 460545
rect 462991 459845 463348 460545
rect 464048 459845 464405 460545
rect 465105 459845 465462 460545
rect 466162 459845 466519 460545
rect 467219 459845 467576 460545
rect 468276 459845 468505 460545
rect 444052 459473 468505 459845
rect 118930 458967 143881 459077
rect 77870 453273 86346 453288
rect 77870 453140 77981 453273
rect 78114 453140 86346 453273
rect 77870 453124 86346 453140
rect 77870 452882 78295 453124
rect 77870 452749 77991 452882
rect 78124 452749 78295 452882
rect 77870 452710 78295 452749
rect 74576 433754 75955 433884
rect 74576 433654 74642 433754
rect 74742 433654 74810 433754
rect 74910 433654 74978 433754
rect 75078 433654 75146 433754
rect 75246 433654 75314 433754
rect 75414 433654 75482 433754
rect 75582 433654 75650 433754
rect 75750 433654 75818 433754
rect 75918 433732 75954 433754
rect 85125 433732 86346 453124
rect 121375 458462 126950 458967
rect 121375 457241 123379 458462
rect 124600 457241 126950 458462
rect 444052 458773 444322 459473
rect 445022 458773 445379 459473
rect 446079 458773 446436 459473
rect 447136 458773 447493 459473
rect 448193 458773 448550 459473
rect 449250 458773 449607 459473
rect 450307 458773 450664 459473
rect 451364 458773 451721 459473
rect 452421 458773 452778 459473
rect 453478 458773 453835 459473
rect 454535 458773 454892 459473
rect 455592 458773 455949 459473
rect 456649 458773 457006 459473
rect 457706 458773 458063 459473
rect 458763 458773 459120 459473
rect 459820 458773 460177 459473
rect 460877 458773 461234 459473
rect 461934 458773 462291 459473
rect 462991 458773 463348 459473
rect 464048 458773 464405 459473
rect 465105 458773 465462 459473
rect 466162 458773 466519 459473
rect 467219 458773 467576 459473
rect 468276 458773 468505 459473
rect 444052 458401 468505 458773
rect 444052 457701 444322 458401
rect 445022 457701 445379 458401
rect 446079 457701 446436 458401
rect 447136 457701 447493 458401
rect 448193 457701 448550 458401
rect 449250 457701 449607 458401
rect 450307 457701 450664 458401
rect 451364 457701 451721 458401
rect 452421 457701 452778 458401
rect 453478 457701 453835 458401
rect 454535 457701 454892 458401
rect 455592 457701 455949 458401
rect 456649 457701 457006 458401
rect 457706 457701 458063 458401
rect 458763 457701 459120 458401
rect 459820 457701 460177 458401
rect 460877 457701 461234 458401
rect 461934 457701 462291 458401
rect 462991 457701 463348 458401
rect 464048 457701 464405 458401
rect 465105 457701 465462 458401
rect 466162 457701 466519 458401
rect 467219 457701 467576 458401
rect 468276 457701 468505 458401
rect 444052 457364 468505 457701
rect 121375 456782 126950 457241
rect 121375 456620 125479 456782
rect 121375 455399 123282 456620
rect 124503 455561 125479 456620
rect 126700 455561 126950 456782
rect 124503 455399 126950 455561
rect 121375 454423 126950 455399
rect 121375 453202 123056 454423
rect 124277 453369 126950 454423
rect 124277 453202 125729 453369
rect 121375 452148 125729 453202
rect 121375 452129 126950 452148
rect 121375 450908 122862 452129
rect 124083 450908 126950 452129
rect 121375 449640 126950 450908
rect 121375 449576 125729 449640
rect 121375 448355 122765 449576
rect 123986 448419 125729 449576
rect 126950 448419 126959 449640
rect 123986 448355 126950 448419
rect 121375 447249 126950 448355
rect 121375 446028 122603 447249
rect 123824 447194 126950 447249
rect 123824 446028 125729 447194
rect 121375 445973 125729 446028
rect 121375 445964 126950 445973
rect 121375 445963 126869 445964
rect 75918 433654 86346 433732
rect 74576 433596 86346 433654
rect 74576 433496 74642 433596
rect 74742 433496 74810 433596
rect 74910 433496 74978 433596
rect 75078 433496 75146 433596
rect 75246 433496 75314 433596
rect 75414 433496 75482 433596
rect 75582 433496 75650 433596
rect 75750 433496 75818 433596
rect 75918 433496 86346 433596
rect 74576 433438 86346 433496
rect 74576 433338 74642 433438
rect 74742 433338 74810 433438
rect 74910 433338 74978 433438
rect 75078 433338 75146 433438
rect 75246 433338 75314 433438
rect 75414 433338 75482 433438
rect 75582 433338 75650 433438
rect 75750 433338 75818 433438
rect 75918 433338 86346 433438
rect 74576 433280 86346 433338
rect 74576 433180 74642 433280
rect 74742 433180 74810 433280
rect 74910 433180 74978 433280
rect 75078 433180 75146 433280
rect 75246 433180 75314 433280
rect 75414 433180 75482 433280
rect 75582 433180 75650 433280
rect 75750 433180 75818 433280
rect 75918 433180 86346 433280
rect 74576 433122 86346 433180
rect 74576 433022 74642 433122
rect 74742 433022 74810 433122
rect 74910 433022 74978 433122
rect 75078 433022 75146 433122
rect 75246 433022 75314 433122
rect 75414 433022 75482 433122
rect 75582 433022 75650 433122
rect 75750 433022 75818 433122
rect 75918 433022 86346 433122
rect 74576 432964 86346 433022
rect 74576 432864 74642 432964
rect 74742 432864 74810 432964
rect 74910 432864 74978 432964
rect 75078 432864 75146 432964
rect 75246 432864 75314 432964
rect 75414 432864 75482 432964
rect 75582 432864 75650 432964
rect 75750 432864 75818 432964
rect 75918 432864 86346 432964
rect 74576 432806 86346 432864
rect 74576 432706 74642 432806
rect 74742 432706 74810 432806
rect 74910 432706 74978 432806
rect 75078 432706 75146 432806
rect 75246 432706 75314 432806
rect 75414 432706 75482 432806
rect 75582 432706 75650 432806
rect 75750 432706 75818 432806
rect 75918 432706 86346 432806
rect 74576 432648 86346 432706
rect 74576 432548 74642 432648
rect 74742 432548 74810 432648
rect 74910 432548 74978 432648
rect 75078 432548 75146 432648
rect 75246 432548 75314 432648
rect 75414 432548 75482 432648
rect 75582 432548 75650 432648
rect 75750 432548 75818 432648
rect 75918 432548 86346 432648
rect 74576 432511 86346 432548
rect 74676 413817 76190 413905
rect 74676 413717 74761 413817
rect 74861 413717 74929 413817
rect 75029 413717 75097 413817
rect 75197 413717 75265 413817
rect 75365 413717 75433 413817
rect 75533 413717 75601 413817
rect 75701 413717 75769 413817
rect 75869 413717 75937 413817
rect 76037 413717 76190 413817
rect 74676 413659 76190 413717
rect 74676 413559 74761 413659
rect 74861 413559 74929 413659
rect 75029 413559 75097 413659
rect 75197 413559 75265 413659
rect 75365 413559 75433 413659
rect 75533 413559 75601 413659
rect 75701 413559 75769 413659
rect 75869 413559 75937 413659
rect 76037 413559 76190 413659
rect 74676 413542 76190 413559
rect 85125 413542 86346 432511
rect 74676 413501 86346 413542
rect 74676 413401 74761 413501
rect 74861 413401 74929 413501
rect 75029 413401 75097 413501
rect 75197 413401 75265 413501
rect 75365 413401 75433 413501
rect 75533 413401 75601 413501
rect 75701 413401 75769 413501
rect 75869 413401 75937 413501
rect 76037 413401 86346 413501
rect 74676 413343 86346 413401
rect 74676 413243 74761 413343
rect 74861 413243 74929 413343
rect 75029 413243 75097 413343
rect 75197 413243 75265 413343
rect 75365 413243 75433 413343
rect 75533 413243 75601 413343
rect 75701 413243 75769 413343
rect 75869 413243 75937 413343
rect 76037 413243 86346 413343
rect 74676 413185 86346 413243
rect 74676 413085 74761 413185
rect 74861 413085 74929 413185
rect 75029 413085 75097 413185
rect 75197 413085 75265 413185
rect 75365 413085 75433 413185
rect 75533 413085 75601 413185
rect 75701 413085 75769 413185
rect 75869 413085 75937 413185
rect 76037 413085 86346 413185
rect 74676 413027 86346 413085
rect 74676 412927 74761 413027
rect 74861 412927 74929 413027
rect 75029 412927 75097 413027
rect 75197 412927 75265 413027
rect 75365 412927 75433 413027
rect 75533 412927 75601 413027
rect 75701 412927 75769 413027
rect 75869 412927 75937 413027
rect 76037 412927 86346 413027
rect 74676 412869 86346 412927
rect 74676 412769 74761 412869
rect 74861 412769 74929 412869
rect 75029 412769 75097 412869
rect 75197 412769 75265 412869
rect 75365 412769 75433 412869
rect 75533 412769 75601 412869
rect 75701 412769 75769 412869
rect 75869 412769 75937 412869
rect 76037 412769 86346 412869
rect 74676 412711 86346 412769
rect 74676 412611 74761 412711
rect 74861 412611 74929 412711
rect 75029 412611 75097 412711
rect 75197 412611 75265 412711
rect 75365 412611 75433 412711
rect 75533 412611 75601 412711
rect 75701 412611 75769 412711
rect 75869 412611 75937 412711
rect 76037 412611 86346 412711
rect 74676 412321 86346 412611
rect 74676 412310 76190 412321
rect 74713 393959 76091 394003
rect 85125 393959 86346 412321
rect 74713 393951 86346 393959
rect 74713 393851 74779 393951
rect 74879 393851 74947 393951
rect 75047 393851 75115 393951
rect 75215 393851 75283 393951
rect 75383 393851 75451 393951
rect 75551 393851 75619 393951
rect 75719 393851 75787 393951
rect 75887 393851 75955 393951
rect 76055 393851 86346 393951
rect 74713 393793 86346 393851
rect 74713 393693 74779 393793
rect 74879 393693 74947 393793
rect 75047 393693 75115 393793
rect 75215 393693 75283 393793
rect 75383 393693 75451 393793
rect 75551 393693 75619 393793
rect 75719 393693 75787 393793
rect 75887 393693 75955 393793
rect 76055 393693 86346 393793
rect 74713 393635 86346 393693
rect 74713 393535 74779 393635
rect 74879 393535 74947 393635
rect 75047 393535 75115 393635
rect 75215 393535 75283 393635
rect 75383 393535 75451 393635
rect 75551 393535 75619 393635
rect 75719 393535 75787 393635
rect 75887 393535 75955 393635
rect 76055 393535 86346 393635
rect 74713 393477 86346 393535
rect 74713 393377 74779 393477
rect 74879 393377 74947 393477
rect 75047 393377 75115 393477
rect 75215 393377 75283 393477
rect 75383 393377 75451 393477
rect 75551 393377 75619 393477
rect 75719 393377 75787 393477
rect 75887 393377 75955 393477
rect 76055 393377 86346 393477
rect 74713 393319 86346 393377
rect 74713 393219 74779 393319
rect 74879 393219 74947 393319
rect 75047 393219 75115 393319
rect 75215 393219 75283 393319
rect 75383 393219 75451 393319
rect 75551 393219 75619 393319
rect 75719 393219 75787 393319
rect 75887 393219 75955 393319
rect 76055 393219 86346 393319
rect 74713 393161 86346 393219
rect 74713 393061 74779 393161
rect 74879 393061 74947 393161
rect 75047 393061 75115 393161
rect 75215 393061 75283 393161
rect 75383 393061 75451 393161
rect 75551 393061 75619 393161
rect 75719 393061 75787 393161
rect 75887 393061 75955 393161
rect 76055 393061 86346 393161
rect 74713 393003 86346 393061
rect 74713 392903 74779 393003
rect 74879 392903 74947 393003
rect 75047 392903 75115 393003
rect 75215 392903 75283 393003
rect 75383 392903 75451 393003
rect 75551 392903 75619 393003
rect 75719 392903 75787 393003
rect 75887 392903 75955 393003
rect 76055 392903 86346 393003
rect 74713 392845 86346 392903
rect 74713 392745 74779 392845
rect 74879 392745 74947 392845
rect 75047 392745 75115 392845
rect 75215 392745 75283 392845
rect 75383 392745 75451 392845
rect 75551 392745 75619 392845
rect 75719 392745 75787 392845
rect 75887 392745 75955 392845
rect 76055 392745 86346 392845
rect 74713 392738 86346 392745
rect 74713 392708 76091 392738
rect 74618 353816 75996 353868
rect 85125 353816 86346 392738
rect 121127 367465 127852 367981
rect 121127 367315 122043 367465
rect 122193 367315 122311 367465
rect 122461 367315 122579 367465
rect 122729 367315 122847 367465
rect 122997 367315 123115 367465
rect 123265 367315 123383 367465
rect 123533 367315 123651 367465
rect 123801 367315 123919 367465
rect 124069 367315 124187 367465
rect 124337 367315 124455 367465
rect 124605 367315 127852 367465
rect 121127 367227 127852 367315
rect 121127 367077 122043 367227
rect 122193 367077 122311 367227
rect 122461 367077 122579 367227
rect 122729 367077 122847 367227
rect 122997 367077 123115 367227
rect 123265 367077 123383 367227
rect 123533 367077 123651 367227
rect 123801 367077 123919 367227
rect 124069 367077 124187 367227
rect 124337 367077 124455 367227
rect 124605 367077 127852 367227
rect 121127 366989 127852 367077
rect 121127 366839 122043 366989
rect 122193 366839 122311 366989
rect 122461 366839 122579 366989
rect 122729 366839 122847 366989
rect 122997 366839 123115 366989
rect 123265 366839 123383 366989
rect 123533 366839 123651 366989
rect 123801 366839 123919 366989
rect 124069 366839 124187 366989
rect 124337 366839 124455 366989
rect 124605 366839 127852 366989
rect 121127 366751 127852 366839
rect 121127 366601 122043 366751
rect 122193 366601 122311 366751
rect 122461 366601 122579 366751
rect 122729 366601 122847 366751
rect 122997 366601 123115 366751
rect 123265 366601 123383 366751
rect 123533 366601 123651 366751
rect 123801 366601 123919 366751
rect 124069 366601 124187 366751
rect 124337 366601 124455 366751
rect 124605 366601 127852 366751
rect 121127 366513 127852 366601
rect 121127 366363 122043 366513
rect 122193 366363 122311 366513
rect 122461 366363 122579 366513
rect 122729 366363 122847 366513
rect 122997 366363 123115 366513
rect 123265 366363 123383 366513
rect 123533 366363 123651 366513
rect 123801 366363 123919 366513
rect 124069 366363 124187 366513
rect 124337 366363 124455 366513
rect 124605 366363 127852 366513
rect 121127 366275 127852 366363
rect 121127 366125 122043 366275
rect 122193 366125 122311 366275
rect 122461 366125 122579 366275
rect 122729 366125 122847 366275
rect 122997 366125 123115 366275
rect 123265 366125 123383 366275
rect 123533 366125 123651 366275
rect 123801 366125 123919 366275
rect 124069 366125 124187 366275
rect 124337 366125 124455 366275
rect 124605 366125 127852 366275
rect 121127 366037 127852 366125
rect 121127 365887 122043 366037
rect 122193 365887 122311 366037
rect 122461 365887 122579 366037
rect 122729 365887 122847 366037
rect 122997 365887 123115 366037
rect 123265 365887 123383 366037
rect 123533 365887 123651 366037
rect 123801 365887 123919 366037
rect 124069 365887 124187 366037
rect 124337 365887 124455 366037
rect 124605 365887 127852 366037
rect 121127 365799 127852 365887
rect 121127 365649 122043 365799
rect 122193 365649 122311 365799
rect 122461 365649 122579 365799
rect 122729 365649 122847 365799
rect 122997 365649 123115 365799
rect 123265 365649 123383 365799
rect 123533 365649 123651 365799
rect 123801 365649 123919 365799
rect 124069 365649 124187 365799
rect 124337 365649 124455 365799
rect 124605 365649 127852 365799
rect 121127 365561 127852 365649
rect 121127 365411 122043 365561
rect 122193 365411 122311 365561
rect 122461 365411 122579 365561
rect 122729 365411 122847 365561
rect 122997 365411 123115 365561
rect 123265 365411 123383 365561
rect 123533 365411 123651 365561
rect 123801 365411 123919 365561
rect 124069 365411 124187 365561
rect 124337 365411 124455 365561
rect 124605 365411 127852 365561
rect 121127 365323 127852 365411
rect 121127 365173 122043 365323
rect 122193 365173 122311 365323
rect 122461 365173 122579 365323
rect 122729 365173 122847 365323
rect 122997 365173 123115 365323
rect 123265 365173 123383 365323
rect 123533 365173 123651 365323
rect 123801 365173 123919 365323
rect 124069 365173 124187 365323
rect 124337 365173 124455 365323
rect 124605 365173 127852 365323
rect 121127 364498 127852 365173
rect 74618 353790 86346 353816
rect 74618 353690 74684 353790
rect 74784 353690 74852 353790
rect 74952 353690 75020 353790
rect 75120 353690 75188 353790
rect 75288 353690 75356 353790
rect 75456 353690 75524 353790
rect 75624 353690 75692 353790
rect 75792 353690 75860 353790
rect 75960 353690 86346 353790
rect 74618 353632 86346 353690
rect 74618 353532 74684 353632
rect 74784 353532 74852 353632
rect 74952 353532 75020 353632
rect 75120 353532 75188 353632
rect 75288 353532 75356 353632
rect 75456 353532 75524 353632
rect 75624 353532 75692 353632
rect 75792 353532 75860 353632
rect 75960 353532 86346 353632
rect 74618 353474 86346 353532
rect 74618 353374 74684 353474
rect 74784 353374 74852 353474
rect 74952 353374 75020 353474
rect 75120 353374 75188 353474
rect 75288 353374 75356 353474
rect 75456 353374 75524 353474
rect 75624 353374 75692 353474
rect 75792 353374 75860 353474
rect 75960 353374 86346 353474
rect 74618 353316 86346 353374
rect 74618 353216 74684 353316
rect 74784 353216 74852 353316
rect 74952 353216 75020 353316
rect 75120 353216 75188 353316
rect 75288 353216 75356 353316
rect 75456 353216 75524 353316
rect 75624 353216 75692 353316
rect 75792 353216 75860 353316
rect 75960 353216 86346 353316
rect 74618 353158 86346 353216
rect 74618 353058 74684 353158
rect 74784 353058 74852 353158
rect 74952 353058 75020 353158
rect 75120 353058 75188 353158
rect 75288 353058 75356 353158
rect 75456 353058 75524 353158
rect 75624 353058 75692 353158
rect 75792 353058 75860 353158
rect 75960 353058 86346 353158
rect 74618 353000 86346 353058
rect 74618 352900 74684 353000
rect 74784 352900 74852 353000
rect 74952 352900 75020 353000
rect 75120 352900 75188 353000
rect 75288 352900 75356 353000
rect 75456 352900 75524 353000
rect 75624 352900 75692 353000
rect 75792 352900 75860 353000
rect 75960 352900 86346 353000
rect 74618 352842 86346 352900
rect 74618 352742 74684 352842
rect 74784 352742 74852 352842
rect 74952 352742 75020 352842
rect 75120 352742 75188 352842
rect 75288 352742 75356 352842
rect 75456 352742 75524 352842
rect 75624 352742 75692 352842
rect 75792 352742 75860 352842
rect 75960 352742 86346 352842
rect 74618 352684 86346 352742
rect 74618 352584 74684 352684
rect 74784 352584 74852 352684
rect 74952 352584 75020 352684
rect 75120 352584 75188 352684
rect 75288 352584 75356 352684
rect 75456 352584 75524 352684
rect 75624 352584 75692 352684
rect 75792 352584 75860 352684
rect 75960 352595 86346 352684
rect 75960 352584 75996 352595
rect 74618 352547 75996 352584
rect 85125 333888 86346 352595
rect 74558 333805 86346 333888
rect 74558 333705 74626 333805
rect 74726 333705 74794 333805
rect 74894 333705 74962 333805
rect 75062 333705 75130 333805
rect 75230 333705 75298 333805
rect 75398 333705 75466 333805
rect 75566 333705 75634 333805
rect 75734 333705 75802 333805
rect 75902 333705 86346 333805
rect 74558 333647 86346 333705
rect 74558 333547 74626 333647
rect 74726 333547 74794 333647
rect 74894 333547 74962 333647
rect 75062 333547 75130 333647
rect 75230 333547 75298 333647
rect 75398 333547 75466 333647
rect 75566 333547 75634 333647
rect 75734 333547 75802 333647
rect 75902 333547 86346 333647
rect 74558 333489 86346 333547
rect 74558 333389 74626 333489
rect 74726 333389 74794 333489
rect 74894 333389 74962 333489
rect 75062 333389 75130 333489
rect 75230 333389 75298 333489
rect 75398 333389 75466 333489
rect 75566 333389 75634 333489
rect 75734 333389 75802 333489
rect 75902 333389 86346 333489
rect 74558 333331 86346 333389
rect 74558 333231 74626 333331
rect 74726 333231 74794 333331
rect 74894 333231 74962 333331
rect 75062 333231 75130 333331
rect 75230 333231 75298 333331
rect 75398 333231 75466 333331
rect 75566 333231 75634 333331
rect 75734 333231 75802 333331
rect 75902 333231 86346 333331
rect 74558 333173 86346 333231
rect 74558 333073 74626 333173
rect 74726 333073 74794 333173
rect 74894 333073 74962 333173
rect 75062 333073 75130 333173
rect 75230 333073 75298 333173
rect 75398 333073 75466 333173
rect 75566 333073 75634 333173
rect 75734 333073 75802 333173
rect 75902 333073 86346 333173
rect 74558 333015 86346 333073
rect 74558 332915 74626 333015
rect 74726 332915 74794 333015
rect 74894 332915 74962 333015
rect 75062 332915 75130 333015
rect 75230 332915 75298 333015
rect 75398 332915 75466 333015
rect 75566 332915 75634 333015
rect 75734 332915 75802 333015
rect 75902 332915 86346 333015
rect 74558 332857 86346 332915
rect 74558 332757 74626 332857
rect 74726 332757 74794 332857
rect 74894 332757 74962 332857
rect 75062 332757 75130 332857
rect 75230 332757 75298 332857
rect 75398 332757 75466 332857
rect 75566 332757 75634 332857
rect 75734 332757 75802 332857
rect 75902 332757 86346 332857
rect 74558 332699 86346 332757
rect 74558 332667 74626 332699
rect 74560 332599 74626 332667
rect 74726 332599 74794 332699
rect 74894 332599 74962 332699
rect 75062 332599 75130 332699
rect 75230 332599 75298 332699
rect 75398 332599 75466 332699
rect 75566 332599 75634 332699
rect 75734 332599 75802 332699
rect 75902 332667 86346 332699
rect 75902 332599 75938 332667
rect 74560 332562 75938 332599
rect 85125 321317 86346 332667
rect 443499 149850 468321 150276
rect 443499 149665 468566 149850
rect 443499 148965 443943 149665
rect 444643 148965 445021 149665
rect 445721 148965 446099 149665
rect 446799 148965 447177 149665
rect 447877 148965 448255 149665
rect 448955 148965 449333 149665
rect 450033 148965 450411 149665
rect 451111 148965 451489 149665
rect 452189 148965 452567 149665
rect 453267 148965 453645 149665
rect 454345 148965 454723 149665
rect 455423 148965 455801 149665
rect 456501 148965 456879 149665
rect 457579 148965 457957 149665
rect 458657 148965 459035 149665
rect 459735 148965 460113 149665
rect 460813 148965 461191 149665
rect 461891 148965 462269 149665
rect 462969 148965 463347 149665
rect 464047 148965 464425 149665
rect 465125 148965 465503 149665
rect 466203 148965 466581 149665
rect 467281 148965 467659 149665
rect 468359 148965 468566 149665
rect 443499 148644 468566 148965
rect 443499 147944 443943 148644
rect 444643 147944 445021 148644
rect 445721 147944 446099 148644
rect 446799 147944 447177 148644
rect 447877 147944 448255 148644
rect 448955 147944 449333 148644
rect 450033 147944 450411 148644
rect 451111 147944 451489 148644
rect 452189 147944 452567 148644
rect 453267 147944 453645 148644
rect 454345 147944 454723 148644
rect 455423 147944 455801 148644
rect 456501 147944 456879 148644
rect 457579 147944 457957 148644
rect 458657 147944 459035 148644
rect 459735 147944 460113 148644
rect 460813 147944 461191 148644
rect 461891 147944 462269 148644
rect 462969 147944 463347 148644
rect 464047 147944 464425 148644
rect 465125 147944 465503 148644
rect 466203 147944 466581 148644
rect 467281 147944 467659 148644
rect 468359 147944 468566 148644
rect 443499 147623 468566 147944
rect 443499 146923 443943 147623
rect 444643 146923 445021 147623
rect 445721 146923 446099 147623
rect 446799 146923 447177 147623
rect 447877 146923 448255 147623
rect 448955 146923 449333 147623
rect 450033 146923 450411 147623
rect 451111 146923 451489 147623
rect 452189 146923 452567 147623
rect 453267 146923 453645 147623
rect 454345 146923 454723 147623
rect 455423 146923 455801 147623
rect 456501 146923 456879 147623
rect 457579 146923 457957 147623
rect 458657 146923 459035 147623
rect 459735 146923 460113 147623
rect 460813 146923 461191 147623
rect 461891 146923 462269 147623
rect 462969 146923 463347 147623
rect 464047 146923 464425 147623
rect 465125 146923 465503 147623
rect 466203 146923 466581 147623
rect 467281 146923 467659 147623
rect 468359 146923 468566 147623
rect 443499 146602 468566 146923
rect 121369 145939 142442 146041
rect 443499 145939 443943 146602
rect 121363 145902 443943 145939
rect 444643 145902 445021 146602
rect 445721 145902 446099 146602
rect 446799 145902 447177 146602
rect 447877 145902 448255 146602
rect 448955 145902 449333 146602
rect 450033 145902 450411 146602
rect 451111 145902 451489 146602
rect 452189 145902 452567 146602
rect 453267 145902 453645 146602
rect 454345 145902 454723 146602
rect 455423 145902 455801 146602
rect 456501 145902 456879 146602
rect 457579 145902 457957 146602
rect 458657 145902 459035 146602
rect 459735 145902 460113 146602
rect 460813 145902 461191 146602
rect 461891 145902 462269 146602
rect 462969 145902 463347 146602
rect 464047 145902 464425 146602
rect 465125 145902 465503 146602
rect 466203 145902 466581 146602
rect 467281 145902 467659 146602
rect 468359 145902 468566 146602
rect 121363 145581 468566 145902
rect 121363 145196 443943 145581
rect 121363 144196 121694 145196
rect 122694 144196 123035 145196
rect 124035 144196 124376 145196
rect 125376 144196 125717 145196
rect 126717 144196 127058 145196
rect 128058 144196 128399 145196
rect 129399 144196 129740 145196
rect 130740 144196 131081 145196
rect 132081 144196 132422 145196
rect 133422 144196 133763 145196
rect 134763 144196 135104 145196
rect 136104 144196 136445 145196
rect 137445 144196 137786 145196
rect 138786 144196 139127 145196
rect 140127 144196 140468 145196
rect 141468 144881 443943 145196
rect 444643 144881 445021 145581
rect 445721 144881 446099 145581
rect 446799 144881 447177 145581
rect 447877 144881 448255 145581
rect 448955 144881 449333 145581
rect 450033 144881 450411 145581
rect 451111 144881 451489 145581
rect 452189 144881 452567 145581
rect 453267 144881 453645 145581
rect 454345 144881 454723 145581
rect 455423 144881 455801 145581
rect 456501 144881 456879 145581
rect 457579 144881 457957 145581
rect 458657 144881 459035 145581
rect 459735 144881 460113 145581
rect 460813 144881 461191 145581
rect 461891 144881 462269 145581
rect 462969 144881 463347 145581
rect 464047 144881 464425 145581
rect 465125 144881 465503 145581
rect 466203 144881 466581 145581
rect 467281 144881 467659 145581
rect 468359 144881 468566 145581
rect 141468 144560 468566 144881
rect 141468 144196 443943 144560
rect 121363 143860 443943 144196
rect 444643 143860 445021 144560
rect 445721 143860 446099 144560
rect 446799 143860 447177 144560
rect 447877 143860 448255 144560
rect 448955 143860 449333 144560
rect 450033 143860 450411 144560
rect 451111 143860 451489 144560
rect 452189 143860 452567 144560
rect 453267 143860 453645 144560
rect 454345 143860 454723 144560
rect 455423 143860 455801 144560
rect 456501 143860 456879 144560
rect 457579 143860 457957 144560
rect 458657 143860 459035 144560
rect 459735 143860 460113 144560
rect 460813 143860 461191 144560
rect 461891 143860 462269 144560
rect 462969 143860 463347 144560
rect 464047 143860 464425 144560
rect 465125 143860 465503 144560
rect 466203 143860 466581 144560
rect 467281 143860 467659 144560
rect 468359 143860 468566 144560
rect 121363 143855 468566 143860
rect 121363 142855 121694 143855
rect 122694 142855 123035 143855
rect 124035 142855 124376 143855
rect 125376 142855 125717 143855
rect 126717 142855 127058 143855
rect 128058 142855 128399 143855
rect 129399 142855 129740 143855
rect 130740 142855 131081 143855
rect 132081 142855 132422 143855
rect 133422 142855 133763 143855
rect 134763 142855 135104 143855
rect 136104 142855 136445 143855
rect 137445 142855 137786 143855
rect 138786 142855 139127 143855
rect 140127 142855 140468 143855
rect 141468 143539 468566 143855
rect 141468 142855 443943 143539
rect 121363 142839 443943 142855
rect 444643 142839 445021 143539
rect 445721 142839 446099 143539
rect 446799 142839 447177 143539
rect 447877 142839 448255 143539
rect 448955 142839 449333 143539
rect 450033 142839 450411 143539
rect 451111 142839 451489 143539
rect 452189 142839 452567 143539
rect 453267 142839 453645 143539
rect 454345 142839 454723 143539
rect 455423 142839 455801 143539
rect 456501 142839 456879 143539
rect 457579 142839 457957 143539
rect 458657 142839 459035 143539
rect 459735 142839 460113 143539
rect 460813 142839 461191 143539
rect 461891 142839 462269 143539
rect 462969 142839 463347 143539
rect 464047 142839 464425 143539
rect 465125 142839 465503 143539
rect 466203 142839 466581 143539
rect 467281 142839 467659 143539
rect 468359 142839 468566 143539
rect 121363 142518 468566 142839
rect 121363 142514 443943 142518
rect 121363 141514 121694 142514
rect 122694 141514 123035 142514
rect 124035 141514 124376 142514
rect 125376 141514 125717 142514
rect 126717 141514 127058 142514
rect 128058 141514 128399 142514
rect 129399 141514 129740 142514
rect 130740 141514 131081 142514
rect 132081 141514 132422 142514
rect 133422 141514 133763 142514
rect 134763 141514 135104 142514
rect 136104 141514 136445 142514
rect 137445 141514 137786 142514
rect 138786 141514 139127 142514
rect 140127 141514 140468 142514
rect 141468 141818 443943 142514
rect 444643 141818 445021 142518
rect 445721 141818 446099 142518
rect 446799 141818 447177 142518
rect 447877 141818 448255 142518
rect 448955 141818 449333 142518
rect 450033 141818 450411 142518
rect 451111 141818 451489 142518
rect 452189 141818 452567 142518
rect 453267 141818 453645 142518
rect 454345 141818 454723 142518
rect 455423 141818 455801 142518
rect 456501 141818 456879 142518
rect 457579 141818 457957 142518
rect 458657 141818 459035 142518
rect 459735 141818 460113 142518
rect 460813 141818 461191 142518
rect 461891 141818 462269 142518
rect 462969 141818 463347 142518
rect 464047 141818 464425 142518
rect 465125 141818 465503 142518
rect 466203 141818 466581 142518
rect 467281 141818 467659 142518
rect 468359 141818 468566 142518
rect 141468 141514 468566 141818
rect 121363 141497 468566 141514
rect 121363 141173 443943 141497
rect 121363 140173 121694 141173
rect 122694 140173 123035 141173
rect 124035 140173 124376 141173
rect 125376 140173 125717 141173
rect 126717 140173 127058 141173
rect 128058 140173 128399 141173
rect 129399 140173 129740 141173
rect 130740 140173 131081 141173
rect 132081 140173 132422 141173
rect 133422 140173 133763 141173
rect 134763 140173 135104 141173
rect 136104 140173 136445 141173
rect 137445 140173 137786 141173
rect 138786 140173 139127 141173
rect 140127 140173 140468 141173
rect 141468 140797 443943 141173
rect 444643 140797 445021 141497
rect 445721 140797 446099 141497
rect 446799 140797 447177 141497
rect 447877 140797 448255 141497
rect 448955 140797 449333 141497
rect 450033 140797 450411 141497
rect 451111 140797 451489 141497
rect 452189 140797 452567 141497
rect 453267 140797 453645 141497
rect 454345 140797 454723 141497
rect 455423 140797 455801 141497
rect 456501 140797 456879 141497
rect 457579 140797 457957 141497
rect 458657 140797 459035 141497
rect 459735 140797 460113 141497
rect 460813 140797 461191 141497
rect 461891 140797 462269 141497
rect 462969 140797 463347 141497
rect 464047 140797 464425 141497
rect 465125 140797 465503 141497
rect 466203 140797 466581 141497
rect 467281 140797 467659 141497
rect 468359 140797 468566 141497
rect 141468 140476 468566 140797
rect 141468 140173 443943 140476
rect 121363 139832 443943 140173
rect 121363 138832 121694 139832
rect 122694 138832 123035 139832
rect 124035 138832 124376 139832
rect 125376 138832 125717 139832
rect 126717 138832 127058 139832
rect 128058 138832 128399 139832
rect 129399 138832 129740 139832
rect 130740 138832 131081 139832
rect 132081 138832 132422 139832
rect 133422 138832 133763 139832
rect 134763 138832 135104 139832
rect 136104 138832 136445 139832
rect 137445 138832 137786 139832
rect 138786 138832 139127 139832
rect 140127 138832 140468 139832
rect 141468 139776 443943 139832
rect 444643 139776 445021 140476
rect 445721 139776 446099 140476
rect 446799 139776 447177 140476
rect 447877 139776 448255 140476
rect 448955 139776 449333 140476
rect 450033 139776 450411 140476
rect 451111 139776 451489 140476
rect 452189 139776 452567 140476
rect 453267 139776 453645 140476
rect 454345 139776 454723 140476
rect 455423 139776 455801 140476
rect 456501 139776 456879 140476
rect 457579 139776 457957 140476
rect 458657 139776 459035 140476
rect 459735 139776 460113 140476
rect 460813 139776 461191 140476
rect 461891 139776 462269 140476
rect 462969 139776 463347 140476
rect 464047 139776 464425 140476
rect 465125 139776 465503 140476
rect 466203 139776 466581 140476
rect 467281 139776 467659 140476
rect 468359 139776 468566 140476
rect 141468 139455 468566 139776
rect 141468 138832 443943 139455
rect 121363 138755 443943 138832
rect 444643 138755 445021 139455
rect 445721 138755 446099 139455
rect 446799 138755 447177 139455
rect 447877 138755 448255 139455
rect 448955 138755 449333 139455
rect 450033 138755 450411 139455
rect 451111 138755 451489 139455
rect 452189 138755 452567 139455
rect 453267 138755 453645 139455
rect 454345 138755 454723 139455
rect 455423 138755 455801 139455
rect 456501 138755 456879 139455
rect 457579 138755 457957 139455
rect 458657 138755 459035 139455
rect 459735 138755 460113 139455
rect 460813 138755 461191 139455
rect 461891 138755 462269 139455
rect 462969 138755 463347 139455
rect 464047 138755 464425 139455
rect 465125 138755 465503 139455
rect 466203 138755 466581 139455
rect 467281 138755 467659 139455
rect 468359 138755 468566 139455
rect 121363 138491 468566 138755
rect 121363 137491 121694 138491
rect 122694 137491 123035 138491
rect 124035 137491 124376 138491
rect 125376 137491 125717 138491
rect 126717 137491 127058 138491
rect 128058 137491 128399 138491
rect 129399 137491 129740 138491
rect 130740 137491 131081 138491
rect 132081 137491 132422 138491
rect 133422 137491 133763 138491
rect 134763 137491 135104 138491
rect 136104 137491 136445 138491
rect 137445 137491 137786 138491
rect 138786 137491 139127 138491
rect 140127 137491 140468 138491
rect 141468 138434 468566 138491
rect 141468 137734 443943 138434
rect 444643 137734 445021 138434
rect 445721 137734 446099 138434
rect 446799 137734 447177 138434
rect 447877 137734 448255 138434
rect 448955 137734 449333 138434
rect 450033 137734 450411 138434
rect 451111 137734 451489 138434
rect 452189 137734 452567 138434
rect 453267 137734 453645 138434
rect 454345 137734 454723 138434
rect 455423 137734 455801 138434
rect 456501 137734 456879 138434
rect 457579 137734 457957 138434
rect 458657 137734 459035 138434
rect 459735 137734 460113 138434
rect 460813 137734 461191 138434
rect 461891 137734 462269 138434
rect 462969 137734 463347 138434
rect 464047 137734 464425 138434
rect 465125 137734 465503 138434
rect 466203 137734 466581 138434
rect 467281 137734 467659 138434
rect 468359 137734 468566 138434
rect 141468 137491 468566 137734
rect 121363 137413 468566 137491
rect 121363 137150 443943 137413
rect 121363 136150 121694 137150
rect 122694 136150 123035 137150
rect 124035 136150 124376 137150
rect 125376 136150 125717 137150
rect 126717 136150 127058 137150
rect 128058 136150 128399 137150
rect 129399 136150 129740 137150
rect 130740 136150 131081 137150
rect 132081 136150 132422 137150
rect 133422 136150 133763 137150
rect 134763 136150 135104 137150
rect 136104 136150 136445 137150
rect 137445 136150 137786 137150
rect 138786 136150 139127 137150
rect 140127 136150 140468 137150
rect 141468 136713 443943 137150
rect 444643 136713 445021 137413
rect 445721 136713 446099 137413
rect 446799 136713 447177 137413
rect 447877 136713 448255 137413
rect 448955 136713 449333 137413
rect 450033 136713 450411 137413
rect 451111 136713 451489 137413
rect 452189 136713 452567 137413
rect 453267 136713 453645 137413
rect 454345 136713 454723 137413
rect 455423 136713 455801 137413
rect 456501 136713 456879 137413
rect 457579 136713 457957 137413
rect 458657 136713 459035 137413
rect 459735 136713 460113 137413
rect 460813 136713 461191 137413
rect 461891 136713 462269 137413
rect 462969 136713 463347 137413
rect 464047 136713 464425 137413
rect 465125 136713 465503 137413
rect 466203 136713 466581 137413
rect 467281 136713 467659 137413
rect 468359 136713 468566 137413
rect 141468 136392 468566 136713
rect 141468 136150 443943 136392
rect 121363 135809 443943 136150
rect 121363 134809 121694 135809
rect 122694 134809 123035 135809
rect 124035 134809 124376 135809
rect 125376 134809 125717 135809
rect 126717 134809 127058 135809
rect 128058 134809 128399 135809
rect 129399 134809 129740 135809
rect 130740 134809 131081 135809
rect 132081 134809 132422 135809
rect 133422 134809 133763 135809
rect 134763 134809 135104 135809
rect 136104 134809 136445 135809
rect 137445 134809 137786 135809
rect 138786 134809 139127 135809
rect 140127 134809 140468 135809
rect 141468 135692 443943 135809
rect 444643 135692 445021 136392
rect 445721 135692 446099 136392
rect 446799 135692 447177 136392
rect 447877 135692 448255 136392
rect 448955 135692 449333 136392
rect 450033 135692 450411 136392
rect 451111 135692 451489 136392
rect 452189 135692 452567 136392
rect 453267 135692 453645 136392
rect 454345 135692 454723 136392
rect 455423 135692 455801 136392
rect 456501 135692 456879 136392
rect 457579 135692 457957 136392
rect 458657 135692 459035 136392
rect 459735 135692 460113 136392
rect 460813 135692 461191 136392
rect 461891 135692 462269 136392
rect 462969 135692 463347 136392
rect 464047 135692 464425 136392
rect 465125 135692 465503 136392
rect 466203 135692 466581 136392
rect 467281 135692 467659 136392
rect 468359 135692 468566 136392
rect 141468 135371 468566 135692
rect 141468 134809 443943 135371
rect 121363 134671 443943 134809
rect 444643 134671 445021 135371
rect 445721 134671 446099 135371
rect 446799 134671 447177 135371
rect 447877 134671 448255 135371
rect 448955 134671 449333 135371
rect 450033 134671 450411 135371
rect 451111 134671 451489 135371
rect 452189 134671 452567 135371
rect 453267 134671 453645 135371
rect 454345 134671 454723 135371
rect 455423 134671 455801 135371
rect 456501 134671 456879 135371
rect 457579 134671 457957 135371
rect 458657 134671 459035 135371
rect 459735 134671 460113 135371
rect 460813 134671 461191 135371
rect 461891 134671 462269 135371
rect 462969 134671 463347 135371
rect 464047 134671 464425 135371
rect 465125 134671 465503 135371
rect 466203 134671 466581 135371
rect 467281 134671 467659 135371
rect 468359 134671 468566 135371
rect 121363 134468 468566 134671
rect 121363 133468 121694 134468
rect 122694 133468 123035 134468
rect 124035 133468 124376 134468
rect 125376 133468 125717 134468
rect 126717 133468 127058 134468
rect 128058 133468 128399 134468
rect 129399 133468 129740 134468
rect 130740 133468 131081 134468
rect 132081 133468 132422 134468
rect 133422 133468 133763 134468
rect 134763 133468 135104 134468
rect 136104 133468 136445 134468
rect 137445 133468 137786 134468
rect 138786 133468 139127 134468
rect 140127 133468 140468 134468
rect 141468 134350 468566 134468
rect 141468 133650 443943 134350
rect 444643 133650 445021 134350
rect 445721 133650 446099 134350
rect 446799 133650 447177 134350
rect 447877 133650 448255 134350
rect 448955 133650 449333 134350
rect 450033 133650 450411 134350
rect 451111 133650 451489 134350
rect 452189 133650 452567 134350
rect 453267 133650 453645 134350
rect 454345 133650 454723 134350
rect 455423 133650 455801 134350
rect 456501 133650 456879 134350
rect 457579 133650 457957 134350
rect 458657 133650 459035 134350
rect 459735 133650 460113 134350
rect 460813 133650 461191 134350
rect 461891 133650 462269 134350
rect 462969 133650 463347 134350
rect 464047 133650 464425 134350
rect 465125 133650 465503 134350
rect 466203 133650 466581 134350
rect 467281 133650 467659 134350
rect 468359 133650 468566 134350
rect 141468 133468 468566 133650
rect 121363 133329 468566 133468
rect 121363 133127 443943 133329
rect 121363 132127 121694 133127
rect 122694 132127 123035 133127
rect 124035 132127 124376 133127
rect 125376 132127 125717 133127
rect 126717 132127 127058 133127
rect 128058 132127 128399 133127
rect 129399 132127 129740 133127
rect 130740 132127 131081 133127
rect 132081 132127 132422 133127
rect 133422 132127 133763 133127
rect 134763 132127 135104 133127
rect 136104 132127 136445 133127
rect 137445 132127 137786 133127
rect 138786 132127 139127 133127
rect 140127 132127 140468 133127
rect 141468 132629 443943 133127
rect 444643 132629 445021 133329
rect 445721 132629 446099 133329
rect 446799 132629 447177 133329
rect 447877 132629 448255 133329
rect 448955 132629 449333 133329
rect 450033 132629 450411 133329
rect 451111 132629 451489 133329
rect 452189 132629 452567 133329
rect 453267 132629 453645 133329
rect 454345 132629 454723 133329
rect 455423 132629 455801 133329
rect 456501 132629 456879 133329
rect 457579 132629 457957 133329
rect 458657 132629 459035 133329
rect 459735 132629 460113 133329
rect 460813 132629 461191 133329
rect 461891 132629 462269 133329
rect 462969 132629 463347 133329
rect 464047 132629 464425 133329
rect 465125 132629 465503 133329
rect 466203 132629 466581 133329
rect 467281 132629 467659 133329
rect 468359 132629 468566 133329
rect 141468 132308 468566 132629
rect 141468 132127 443943 132308
rect 121363 131786 443943 132127
rect 121363 130786 121694 131786
rect 122694 130786 123035 131786
rect 124035 130786 124376 131786
rect 125376 130786 125717 131786
rect 126717 130786 127058 131786
rect 128058 130786 128399 131786
rect 129399 130786 129740 131786
rect 130740 130786 131081 131786
rect 132081 130786 132422 131786
rect 133422 130786 133763 131786
rect 134763 130786 135104 131786
rect 136104 130786 136445 131786
rect 137445 130786 137786 131786
rect 138786 130786 139127 131786
rect 140127 130786 140468 131786
rect 141468 131608 443943 131786
rect 444643 131608 445021 132308
rect 445721 131608 446099 132308
rect 446799 131608 447177 132308
rect 447877 131608 448255 132308
rect 448955 131608 449333 132308
rect 450033 131608 450411 132308
rect 451111 131608 451489 132308
rect 452189 131608 452567 132308
rect 453267 131608 453645 132308
rect 454345 131608 454723 132308
rect 455423 131608 455801 132308
rect 456501 131608 456879 132308
rect 457579 131608 457957 132308
rect 458657 131608 459035 132308
rect 459735 131608 460113 132308
rect 460813 131608 461191 132308
rect 461891 131608 462269 132308
rect 462969 131608 463347 132308
rect 464047 131608 464425 132308
rect 465125 131608 465503 132308
rect 466203 131608 466581 132308
rect 467281 131608 467659 132308
rect 468359 131608 468566 132308
rect 141468 131287 468566 131608
rect 141468 130786 443943 131287
rect 121363 130587 443943 130786
rect 444643 130587 445021 131287
rect 445721 130587 446099 131287
rect 446799 130587 447177 131287
rect 447877 130587 448255 131287
rect 448955 130587 449333 131287
rect 450033 130587 450411 131287
rect 451111 130587 451489 131287
rect 452189 130587 452567 131287
rect 453267 130587 453645 131287
rect 454345 130587 454723 131287
rect 455423 130587 455801 131287
rect 456501 130587 456879 131287
rect 457579 130587 457957 131287
rect 458657 130587 459035 131287
rect 459735 130587 460113 131287
rect 460813 130587 461191 131287
rect 461891 130587 462269 131287
rect 462969 130587 463347 131287
rect 464047 130587 464425 131287
rect 465125 130587 465503 131287
rect 466203 130587 466581 131287
rect 467281 130587 467659 131287
rect 468359 130587 468566 131287
rect 121363 130445 468566 130587
rect 121363 129445 121694 130445
rect 122694 129445 123035 130445
rect 124035 129445 124376 130445
rect 125376 129445 125717 130445
rect 126717 129445 127058 130445
rect 128058 129445 128399 130445
rect 129399 129445 129740 130445
rect 130740 129445 131081 130445
rect 132081 129445 132422 130445
rect 133422 129445 133763 130445
rect 134763 129445 135104 130445
rect 136104 129445 136445 130445
rect 137445 129445 137786 130445
rect 138786 129445 139127 130445
rect 140127 129445 140468 130445
rect 141468 130266 468566 130445
rect 141468 129566 443943 130266
rect 444643 129566 445021 130266
rect 445721 129566 446099 130266
rect 446799 129566 447177 130266
rect 447877 129566 448255 130266
rect 448955 129566 449333 130266
rect 450033 129566 450411 130266
rect 451111 129566 451489 130266
rect 452189 129566 452567 130266
rect 453267 129566 453645 130266
rect 454345 129566 454723 130266
rect 455423 129566 455801 130266
rect 456501 129566 456879 130266
rect 457579 129566 457957 130266
rect 458657 129566 459035 130266
rect 459735 129566 460113 130266
rect 460813 129566 461191 130266
rect 461891 129566 462269 130266
rect 462969 129566 463347 130266
rect 464047 129566 464425 130266
rect 465125 129566 465503 130266
rect 466203 129566 466581 130266
rect 467281 129566 467659 130266
rect 468359 129566 468566 130266
rect 141468 129445 468566 129566
rect 121363 129245 468566 129445
rect 121363 129104 443943 129245
rect 121363 128104 121694 129104
rect 122694 128104 123035 129104
rect 124035 128104 124376 129104
rect 125376 128104 125717 129104
rect 126717 128104 127058 129104
rect 128058 128104 128399 129104
rect 129399 128104 129740 129104
rect 130740 128104 131081 129104
rect 132081 128104 132422 129104
rect 133422 128104 133763 129104
rect 134763 128104 135104 129104
rect 136104 128104 136445 129104
rect 137445 128104 137786 129104
rect 138786 128104 139127 129104
rect 140127 128104 140468 129104
rect 141468 128545 443943 129104
rect 444643 128545 445021 129245
rect 445721 128545 446099 129245
rect 446799 128545 447177 129245
rect 447877 128545 448255 129245
rect 448955 128545 449333 129245
rect 450033 128545 450411 129245
rect 451111 128545 451489 129245
rect 452189 128545 452567 129245
rect 453267 128545 453645 129245
rect 454345 128545 454723 129245
rect 455423 128545 455801 129245
rect 456501 128545 456879 129245
rect 457579 128545 457957 129245
rect 458657 128545 459035 129245
rect 459735 128545 460113 129245
rect 460813 128545 461191 129245
rect 461891 128545 462269 129245
rect 462969 128545 463347 129245
rect 464047 128545 464425 129245
rect 465125 128545 465503 129245
rect 466203 128545 466581 129245
rect 467281 128545 467659 129245
rect 468359 128545 468566 129245
rect 141468 128224 468566 128545
rect 141468 128104 443943 128224
rect 121363 127763 443943 128104
rect 121363 126763 121694 127763
rect 122694 126763 123035 127763
rect 124035 126763 124376 127763
rect 125376 126763 125717 127763
rect 126717 126763 127058 127763
rect 128058 126763 128399 127763
rect 129399 126763 129740 127763
rect 130740 126763 131081 127763
rect 132081 126763 132422 127763
rect 133422 126763 133763 127763
rect 134763 126763 135104 127763
rect 136104 126763 136445 127763
rect 137445 126763 137786 127763
rect 138786 126763 139127 127763
rect 140127 126763 140468 127763
rect 141468 127524 443943 127763
rect 444643 127524 445021 128224
rect 445721 127524 446099 128224
rect 446799 127524 447177 128224
rect 447877 127524 448255 128224
rect 448955 127524 449333 128224
rect 450033 127524 450411 128224
rect 451111 127524 451489 128224
rect 452189 127524 452567 128224
rect 453267 127524 453645 128224
rect 454345 127524 454723 128224
rect 455423 127524 455801 128224
rect 456501 127524 456879 128224
rect 457579 127524 457957 128224
rect 458657 127524 459035 128224
rect 459735 127524 460113 128224
rect 460813 127524 461191 128224
rect 461891 127524 462269 128224
rect 462969 127524 463347 128224
rect 464047 127524 464425 128224
rect 465125 127524 465503 128224
rect 466203 127524 466581 128224
rect 467281 127524 467659 128224
rect 468359 127524 468566 128224
rect 141468 127203 468566 127524
rect 141468 126763 443943 127203
rect 121363 126503 443943 126763
rect 444643 126503 445021 127203
rect 445721 126503 446099 127203
rect 446799 126503 447177 127203
rect 447877 126503 448255 127203
rect 448955 126503 449333 127203
rect 450033 126503 450411 127203
rect 451111 126503 451489 127203
rect 452189 126503 452567 127203
rect 453267 126503 453645 127203
rect 454345 126503 454723 127203
rect 455423 126503 455801 127203
rect 456501 126503 456879 127203
rect 457579 126503 457957 127203
rect 458657 126503 459035 127203
rect 459735 126503 460113 127203
rect 460813 126503 461191 127203
rect 461891 126503 462269 127203
rect 462969 126503 463347 127203
rect 464047 126503 464425 127203
rect 465125 126503 465503 127203
rect 466203 126503 466581 127203
rect 467281 126503 467659 127203
rect 468359 126503 468566 127203
rect 121363 126422 468566 126503
rect 121363 125422 121694 126422
rect 122694 125422 123035 126422
rect 124035 125422 124376 126422
rect 125376 125422 125717 126422
rect 126717 125422 127058 126422
rect 128058 125422 128399 126422
rect 129399 125422 129740 126422
rect 130740 125422 131081 126422
rect 132081 125422 132422 126422
rect 133422 125422 133763 126422
rect 134763 125422 135104 126422
rect 136104 125422 136445 126422
rect 137445 125422 137786 126422
rect 138786 125422 139127 126422
rect 140127 125422 140468 126422
rect 141468 126182 468566 126422
rect 141468 125482 443943 126182
rect 444643 125482 445021 126182
rect 445721 125482 446099 126182
rect 446799 125482 447177 126182
rect 447877 125482 448255 126182
rect 448955 125482 449333 126182
rect 450033 125482 450411 126182
rect 451111 125482 451489 126182
rect 452189 125482 452567 126182
rect 453267 125482 453645 126182
rect 454345 125482 454723 126182
rect 455423 125482 455801 126182
rect 456501 125482 456879 126182
rect 457579 125482 457957 126182
rect 458657 125482 459035 126182
rect 459735 125482 460113 126182
rect 460813 125482 461191 126182
rect 461891 125482 462269 126182
rect 462969 125482 463347 126182
rect 464047 125482 464425 126182
rect 465125 125482 465503 126182
rect 466203 125482 466581 126182
rect 467281 125482 467659 126182
rect 468359 125482 468566 126182
rect 141468 125422 468566 125482
rect 121363 125346 468566 125422
rect 121363 125186 468321 125346
rect 121369 124678 142442 125186
rect 443499 125098 468321 125186
rect 481895 124824 508199 125045
rect 481895 124124 482072 124824
rect 482772 124124 483168 124824
rect 483868 124124 484264 124824
rect 484964 124124 485360 124824
rect 486060 124124 486456 124824
rect 487156 124124 487552 124824
rect 488252 124124 488648 124824
rect 489348 124124 489744 124824
rect 490444 124124 490840 124824
rect 491540 124124 491936 124824
rect 492636 124124 493032 124824
rect 493732 124124 494128 124824
rect 494828 124124 495224 124824
rect 495924 124124 496320 124824
rect 497020 124124 497416 124824
rect 498116 124124 498512 124824
rect 499212 124124 499608 124824
rect 500308 124124 500704 124824
rect 501404 124124 501800 124824
rect 502500 124124 502896 124824
rect 503596 124124 503992 124824
rect 504692 124124 505088 124824
rect 505788 124124 506184 124824
rect 506884 124124 507280 124824
rect 507980 124124 508199 124824
rect 481895 123677 508199 124124
rect 481670 123673 508199 123677
rect 481670 122973 482072 123673
rect 482772 122973 483168 123673
rect 483868 122973 484264 123673
rect 484964 122973 485360 123673
rect 486060 122973 486456 123673
rect 487156 122973 487552 123673
rect 488252 122973 488648 123673
rect 489348 122973 489744 123673
rect 490444 122973 490840 123673
rect 491540 122973 491936 123673
rect 492636 122973 493032 123673
rect 493732 122973 494128 123673
rect 494828 122973 495224 123673
rect 495924 122973 496320 123673
rect 497020 122973 497416 123673
rect 498116 122973 498512 123673
rect 499212 122973 499608 123673
rect 500308 122973 500704 123673
rect 501404 122973 501800 123673
rect 502500 122973 502896 123673
rect 503596 122973 503992 123673
rect 504692 122973 505088 123673
rect 505788 122973 506184 123673
rect 506884 122973 507280 123673
rect 507980 122973 508199 123673
rect 481670 122522 508199 122973
rect 481670 121822 482072 122522
rect 482772 121822 483168 122522
rect 483868 121822 484264 122522
rect 484964 121822 485360 122522
rect 486060 121822 486456 122522
rect 487156 121822 487552 122522
rect 488252 121822 488648 122522
rect 489348 121822 489744 122522
rect 490444 121822 490840 122522
rect 491540 121822 491936 122522
rect 492636 121822 493032 122522
rect 493732 121822 494128 122522
rect 494828 121822 495224 122522
rect 495924 121822 496320 122522
rect 497020 121822 497416 122522
rect 498116 121822 498512 122522
rect 499212 121822 499608 122522
rect 500308 121822 500704 122522
rect 501404 121822 501800 122522
rect 502500 121822 502896 122522
rect 503596 121822 503992 122522
rect 504692 121822 505088 122522
rect 505788 121822 506184 122522
rect 506884 121822 507280 122522
rect 507980 121822 508199 122522
rect 481670 121371 508199 121822
rect 481670 120671 482072 121371
rect 482772 120671 483168 121371
rect 483868 120671 484264 121371
rect 484964 120671 485360 121371
rect 486060 120671 486456 121371
rect 487156 120671 487552 121371
rect 488252 120671 488648 121371
rect 489348 120671 489744 121371
rect 490444 120671 490840 121371
rect 491540 120671 491936 121371
rect 492636 120671 493032 121371
rect 493732 120671 494128 121371
rect 494828 120671 495224 121371
rect 495924 120671 496320 121371
rect 497020 120671 497416 121371
rect 498116 120671 498512 121371
rect 499212 120671 499608 121371
rect 500308 120671 500704 121371
rect 501404 120671 501800 121371
rect 502500 120671 502896 121371
rect 503596 120671 503992 121371
rect 504692 120671 505088 121371
rect 505788 120671 506184 121371
rect 506884 120671 507280 121371
rect 507980 120671 508199 121371
rect 88384 119846 111541 120594
rect 88384 119146 89225 119846
rect 89925 119146 90134 119846
rect 90834 119146 91043 119846
rect 91743 119146 91952 119846
rect 92652 119146 92861 119846
rect 93561 119146 93770 119846
rect 94470 119146 94679 119846
rect 95379 119146 95588 119846
rect 96288 119146 96497 119846
rect 97197 119146 97406 119846
rect 98106 119146 98315 119846
rect 99015 119146 99224 119846
rect 99924 119146 100133 119846
rect 100833 119146 101042 119846
rect 101742 119146 101951 119846
rect 102651 119146 102860 119846
rect 103560 119146 103769 119846
rect 104469 119146 104678 119846
rect 105378 119146 105587 119846
rect 106287 119146 106496 119846
rect 107196 119146 107405 119846
rect 108105 119146 108314 119846
rect 109014 119146 109223 119846
rect 109923 119146 110132 119846
rect 110832 119146 111541 119846
rect 88384 118958 111541 119146
rect 88384 118258 89225 118958
rect 89925 118258 90134 118958
rect 90834 118258 91043 118958
rect 91743 118258 91952 118958
rect 92652 118258 92861 118958
rect 93561 118258 93770 118958
rect 94470 118258 94679 118958
rect 95379 118258 95588 118958
rect 96288 118258 96497 118958
rect 97197 118258 97406 118958
rect 98106 118258 98315 118958
rect 99015 118258 99224 118958
rect 99924 118258 100133 118958
rect 100833 118258 101042 118958
rect 101742 118258 101951 118958
rect 102651 118258 102860 118958
rect 103560 118258 103769 118958
rect 104469 118258 104678 118958
rect 105378 118258 105587 118958
rect 106287 118258 106496 118958
rect 107196 118258 107405 118958
rect 108105 118258 108314 118958
rect 109014 118258 109223 118958
rect 109923 118258 110132 118958
rect 110832 118512 111541 118958
rect 481670 120220 508199 120671
rect 481670 119520 482072 120220
rect 482772 119520 483168 120220
rect 483868 119520 484264 120220
rect 484964 119520 485360 120220
rect 486060 119520 486456 120220
rect 487156 119520 487552 120220
rect 488252 119520 488648 120220
rect 489348 119520 489744 120220
rect 490444 119520 490840 120220
rect 491540 119520 491936 120220
rect 492636 119520 493032 120220
rect 493732 119520 494128 120220
rect 494828 119520 495224 120220
rect 495924 119520 496320 120220
rect 497020 119520 497416 120220
rect 498116 119520 498512 120220
rect 499212 119520 499608 120220
rect 500308 119520 500704 120220
rect 501404 119520 501800 120220
rect 502500 119520 502896 120220
rect 503596 119520 503992 120220
rect 504692 119520 505088 120220
rect 505788 119520 506184 120220
rect 506884 119520 507280 120220
rect 507980 119520 508199 120220
rect 481670 119069 508199 119520
rect 481670 118512 482072 119069
rect 110832 118369 482072 118512
rect 482772 118369 483168 119069
rect 483868 118369 484264 119069
rect 484964 118369 485360 119069
rect 486060 118369 486456 119069
rect 487156 118369 487552 119069
rect 488252 118369 488648 119069
rect 489348 118369 489744 119069
rect 490444 118369 490840 119069
rect 491540 118369 491936 119069
rect 492636 118369 493032 119069
rect 493732 118369 494128 119069
rect 494828 118369 495224 119069
rect 495924 118369 496320 119069
rect 497020 118369 497416 119069
rect 498116 118369 498512 119069
rect 499212 118369 499608 119069
rect 500308 118369 500704 119069
rect 501404 118369 501800 119069
rect 502500 118369 502896 119069
rect 503596 118369 503992 119069
rect 504692 118369 505088 119069
rect 505788 118369 506184 119069
rect 506884 118369 507280 119069
rect 507980 118369 508199 119069
rect 110832 118258 508199 118369
rect 88384 118070 508199 118258
rect 88384 117370 89225 118070
rect 89925 117370 90134 118070
rect 90834 117370 91043 118070
rect 91743 117370 91952 118070
rect 92652 117370 92861 118070
rect 93561 117370 93770 118070
rect 94470 117370 94679 118070
rect 95379 117370 95588 118070
rect 96288 117370 96497 118070
rect 97197 117370 97406 118070
rect 98106 117370 98315 118070
rect 99015 117370 99224 118070
rect 99924 117370 100133 118070
rect 100833 117370 101042 118070
rect 101742 117370 101951 118070
rect 102651 117370 102860 118070
rect 103560 117370 103769 118070
rect 104469 117370 104678 118070
rect 105378 117370 105587 118070
rect 106287 117370 106496 118070
rect 107196 117370 107405 118070
rect 108105 117370 108314 118070
rect 109014 117370 109223 118070
rect 109923 117370 110132 118070
rect 110832 117918 508199 118070
rect 110832 117370 482072 117918
rect 88384 117218 482072 117370
rect 482772 117218 483168 117918
rect 483868 117218 484264 117918
rect 484964 117218 485360 117918
rect 486060 117218 486456 117918
rect 487156 117218 487552 117918
rect 488252 117218 488648 117918
rect 489348 117218 489744 117918
rect 490444 117218 490840 117918
rect 491540 117218 491936 117918
rect 492636 117218 493032 117918
rect 493732 117218 494128 117918
rect 494828 117218 495224 117918
rect 495924 117218 496320 117918
rect 497020 117218 497416 117918
rect 498116 117218 498512 117918
rect 499212 117218 499608 117918
rect 500308 117218 500704 117918
rect 501404 117218 501800 117918
rect 502500 117218 502896 117918
rect 503596 117218 503992 117918
rect 504692 117218 505088 117918
rect 505788 117218 506184 117918
rect 506884 117218 507280 117918
rect 507980 117218 508199 117918
rect 88384 117182 508199 117218
rect 88384 116482 89225 117182
rect 89925 116482 90134 117182
rect 90834 116482 91043 117182
rect 91743 116482 91952 117182
rect 92652 116482 92861 117182
rect 93561 116482 93770 117182
rect 94470 116482 94679 117182
rect 95379 116482 95588 117182
rect 96288 116482 96497 117182
rect 97197 116482 97406 117182
rect 98106 116482 98315 117182
rect 99015 116482 99224 117182
rect 99924 116482 100133 117182
rect 100833 116482 101042 117182
rect 101742 116482 101951 117182
rect 102651 116482 102860 117182
rect 103560 116482 103769 117182
rect 104469 116482 104678 117182
rect 105378 116482 105587 117182
rect 106287 116482 106496 117182
rect 107196 116482 107405 117182
rect 108105 116482 108314 117182
rect 109014 116482 109223 117182
rect 109923 116482 110132 117182
rect 110832 116767 508199 117182
rect 110832 116482 482072 116767
rect 88384 116294 482072 116482
rect 88384 115594 89225 116294
rect 89925 115594 90134 116294
rect 90834 115594 91043 116294
rect 91743 115594 91952 116294
rect 92652 115594 92861 116294
rect 93561 115594 93770 116294
rect 94470 115594 94679 116294
rect 95379 115594 95588 116294
rect 96288 115594 96497 116294
rect 97197 115594 97406 116294
rect 98106 115594 98315 116294
rect 99015 115594 99224 116294
rect 99924 115594 100133 116294
rect 100833 115594 101042 116294
rect 101742 115594 101951 116294
rect 102651 115594 102860 116294
rect 103560 115594 103769 116294
rect 104469 115594 104678 116294
rect 105378 115594 105587 116294
rect 106287 115594 106496 116294
rect 107196 115594 107405 116294
rect 108105 115594 108314 116294
rect 109014 115594 109223 116294
rect 109923 115594 110132 116294
rect 110832 116067 482072 116294
rect 482772 116067 483168 116767
rect 483868 116067 484264 116767
rect 484964 116067 485360 116767
rect 486060 116067 486456 116767
rect 487156 116067 487552 116767
rect 488252 116067 488648 116767
rect 489348 116067 489744 116767
rect 490444 116067 490840 116767
rect 491540 116067 491936 116767
rect 492636 116067 493032 116767
rect 493732 116067 494128 116767
rect 494828 116067 495224 116767
rect 495924 116067 496320 116767
rect 497020 116067 497416 116767
rect 498116 116067 498512 116767
rect 499212 116067 499608 116767
rect 500308 116067 500704 116767
rect 501404 116067 501800 116767
rect 502500 116067 502896 116767
rect 503596 116067 503992 116767
rect 504692 116067 505088 116767
rect 505788 116067 506184 116767
rect 506884 116067 507280 116767
rect 507980 116067 508199 116767
rect 110832 115616 508199 116067
rect 110832 115594 482072 115616
rect 88384 115406 482072 115594
rect 88384 114706 89225 115406
rect 89925 114706 90134 115406
rect 90834 114706 91043 115406
rect 91743 114706 91952 115406
rect 92652 114706 92861 115406
rect 93561 114706 93770 115406
rect 94470 114706 94679 115406
rect 95379 114706 95588 115406
rect 96288 114706 96497 115406
rect 97197 114706 97406 115406
rect 98106 114706 98315 115406
rect 99015 114706 99224 115406
rect 99924 114706 100133 115406
rect 100833 114706 101042 115406
rect 101742 114706 101951 115406
rect 102651 114706 102860 115406
rect 103560 114706 103769 115406
rect 104469 114706 104678 115406
rect 105378 114706 105587 115406
rect 106287 114706 106496 115406
rect 107196 114706 107405 115406
rect 108105 114706 108314 115406
rect 109014 114706 109223 115406
rect 109923 114706 110132 115406
rect 110832 114916 482072 115406
rect 482772 114916 483168 115616
rect 483868 114916 484264 115616
rect 484964 114916 485360 115616
rect 486060 114916 486456 115616
rect 487156 114916 487552 115616
rect 488252 114916 488648 115616
rect 489348 114916 489744 115616
rect 490444 114916 490840 115616
rect 491540 114916 491936 115616
rect 492636 114916 493032 115616
rect 493732 114916 494128 115616
rect 494828 114916 495224 115616
rect 495924 114916 496320 115616
rect 497020 114916 497416 115616
rect 498116 114916 498512 115616
rect 499212 114916 499608 115616
rect 500308 114916 500704 115616
rect 501404 114916 501800 115616
rect 502500 114916 502896 115616
rect 503596 114916 503992 115616
rect 504692 114916 505088 115616
rect 505788 114916 506184 115616
rect 506884 114916 507280 115616
rect 507980 114916 508199 115616
rect 110832 114706 508199 114916
rect 88384 114518 508199 114706
rect 88384 113818 89225 114518
rect 89925 113818 90134 114518
rect 90834 113818 91043 114518
rect 91743 113818 91952 114518
rect 92652 113818 92861 114518
rect 93561 113818 93770 114518
rect 94470 113818 94679 114518
rect 95379 113818 95588 114518
rect 96288 113818 96497 114518
rect 97197 113818 97406 114518
rect 98106 113818 98315 114518
rect 99015 113818 99224 114518
rect 99924 113818 100133 114518
rect 100833 113818 101042 114518
rect 101742 113818 101951 114518
rect 102651 113818 102860 114518
rect 103560 113818 103769 114518
rect 104469 113818 104678 114518
rect 105378 113818 105587 114518
rect 106287 113818 106496 114518
rect 107196 113818 107405 114518
rect 108105 113818 108314 114518
rect 109014 113818 109223 114518
rect 109923 113818 110132 114518
rect 110832 114465 508199 114518
rect 110832 113818 482072 114465
rect 88384 113765 482072 113818
rect 482772 113765 483168 114465
rect 483868 113765 484264 114465
rect 484964 113765 485360 114465
rect 486060 113765 486456 114465
rect 487156 113765 487552 114465
rect 488252 113765 488648 114465
rect 489348 113765 489744 114465
rect 490444 113765 490840 114465
rect 491540 113765 491936 114465
rect 492636 113765 493032 114465
rect 493732 113765 494128 114465
rect 494828 113765 495224 114465
rect 495924 113765 496320 114465
rect 497020 113765 497416 114465
rect 498116 113765 498512 114465
rect 499212 113765 499608 114465
rect 500308 113765 500704 114465
rect 501404 113765 501800 114465
rect 502500 113765 502896 114465
rect 503596 113765 503992 114465
rect 504692 113765 505088 114465
rect 505788 113765 506184 114465
rect 506884 113765 507280 114465
rect 507980 113765 508199 114465
rect 88384 113630 508199 113765
rect 88384 112930 89225 113630
rect 89925 112930 90134 113630
rect 90834 112930 91043 113630
rect 91743 112930 91952 113630
rect 92652 112930 92861 113630
rect 93561 112930 93770 113630
rect 94470 112930 94679 113630
rect 95379 112930 95588 113630
rect 96288 112930 96497 113630
rect 97197 112930 97406 113630
rect 98106 112930 98315 113630
rect 99015 112930 99224 113630
rect 99924 112930 100133 113630
rect 100833 112930 101042 113630
rect 101742 112930 101951 113630
rect 102651 112930 102860 113630
rect 103560 112930 103769 113630
rect 104469 112930 104678 113630
rect 105378 112930 105587 113630
rect 106287 112930 106496 113630
rect 107196 112930 107405 113630
rect 108105 112930 108314 113630
rect 109014 112930 109223 113630
rect 109923 112930 110132 113630
rect 110832 113314 508199 113630
rect 110832 112930 482072 113314
rect 88384 112742 482072 112930
rect 88384 112042 89225 112742
rect 89925 112042 90134 112742
rect 90834 112042 91043 112742
rect 91743 112042 91952 112742
rect 92652 112042 92861 112742
rect 93561 112042 93770 112742
rect 94470 112042 94679 112742
rect 95379 112042 95588 112742
rect 96288 112042 96497 112742
rect 97197 112042 97406 112742
rect 98106 112042 98315 112742
rect 99015 112042 99224 112742
rect 99924 112042 100133 112742
rect 100833 112042 101042 112742
rect 101742 112042 101951 112742
rect 102651 112042 102860 112742
rect 103560 112042 103769 112742
rect 104469 112042 104678 112742
rect 105378 112042 105587 112742
rect 106287 112042 106496 112742
rect 107196 112042 107405 112742
rect 108105 112042 108314 112742
rect 109014 112042 109223 112742
rect 109923 112042 110132 112742
rect 110832 112614 482072 112742
rect 482772 112614 483168 113314
rect 483868 112614 484264 113314
rect 484964 112614 485360 113314
rect 486060 112614 486456 113314
rect 487156 112614 487552 113314
rect 488252 112614 488648 113314
rect 489348 112614 489744 113314
rect 490444 112614 490840 113314
rect 491540 112614 491936 113314
rect 492636 112614 493032 113314
rect 493732 112614 494128 113314
rect 494828 112614 495224 113314
rect 495924 112614 496320 113314
rect 497020 112614 497416 113314
rect 498116 112614 498512 113314
rect 499212 112614 499608 113314
rect 500308 112614 500704 113314
rect 501404 112614 501800 113314
rect 502500 112614 502896 113314
rect 503596 112614 503992 113314
rect 504692 112614 505088 113314
rect 505788 112614 506184 113314
rect 506884 112614 507280 113314
rect 507980 112614 508199 113314
rect 110832 112163 508199 112614
rect 110832 112042 482072 112163
rect 88384 111854 482072 112042
rect 88384 111154 89225 111854
rect 89925 111154 90134 111854
rect 90834 111154 91043 111854
rect 91743 111154 91952 111854
rect 92652 111154 92861 111854
rect 93561 111154 93770 111854
rect 94470 111154 94679 111854
rect 95379 111154 95588 111854
rect 96288 111154 96497 111854
rect 97197 111154 97406 111854
rect 98106 111154 98315 111854
rect 99015 111154 99224 111854
rect 99924 111154 100133 111854
rect 100833 111154 101042 111854
rect 101742 111154 101951 111854
rect 102651 111154 102860 111854
rect 103560 111154 103769 111854
rect 104469 111154 104678 111854
rect 105378 111154 105587 111854
rect 106287 111154 106496 111854
rect 107196 111154 107405 111854
rect 108105 111154 108314 111854
rect 109014 111154 109223 111854
rect 109923 111154 110132 111854
rect 110832 111463 482072 111854
rect 482772 111463 483168 112163
rect 483868 111463 484264 112163
rect 484964 111463 485360 112163
rect 486060 111463 486456 112163
rect 487156 111463 487552 112163
rect 488252 111463 488648 112163
rect 489348 111463 489744 112163
rect 490444 111463 490840 112163
rect 491540 111463 491936 112163
rect 492636 111463 493032 112163
rect 493732 111463 494128 112163
rect 494828 111463 495224 112163
rect 495924 111463 496320 112163
rect 497020 111463 497416 112163
rect 498116 111463 498512 112163
rect 499212 111463 499608 112163
rect 500308 111463 500704 112163
rect 501404 111463 501800 112163
rect 502500 111463 502896 112163
rect 503596 111463 503992 112163
rect 504692 111463 505088 112163
rect 505788 111463 506184 112163
rect 506884 111463 507280 112163
rect 507980 111463 508199 112163
rect 110832 111154 508199 111463
rect 88384 111012 508199 111154
rect 88384 110966 482072 111012
rect 88384 110266 89225 110966
rect 89925 110266 90134 110966
rect 90834 110266 91043 110966
rect 91743 110266 91952 110966
rect 92652 110266 92861 110966
rect 93561 110266 93770 110966
rect 94470 110266 94679 110966
rect 95379 110266 95588 110966
rect 96288 110266 96497 110966
rect 97197 110266 97406 110966
rect 98106 110266 98315 110966
rect 99015 110266 99224 110966
rect 99924 110266 100133 110966
rect 100833 110266 101042 110966
rect 101742 110266 101951 110966
rect 102651 110266 102860 110966
rect 103560 110266 103769 110966
rect 104469 110266 104678 110966
rect 105378 110266 105587 110966
rect 106287 110266 106496 110966
rect 107196 110266 107405 110966
rect 108105 110266 108314 110966
rect 109014 110266 109223 110966
rect 109923 110266 110132 110966
rect 110832 110312 482072 110966
rect 482772 110312 483168 111012
rect 483868 110312 484264 111012
rect 484964 110312 485360 111012
rect 486060 110312 486456 111012
rect 487156 110312 487552 111012
rect 488252 110312 488648 111012
rect 489348 110312 489744 111012
rect 490444 110312 490840 111012
rect 491540 110312 491936 111012
rect 492636 110312 493032 111012
rect 493732 110312 494128 111012
rect 494828 110312 495224 111012
rect 495924 110312 496320 111012
rect 497020 110312 497416 111012
rect 498116 110312 498512 111012
rect 499212 110312 499608 111012
rect 500308 110312 500704 111012
rect 501404 110312 501800 111012
rect 502500 110312 502896 111012
rect 503596 110312 503992 111012
rect 504692 110312 505088 111012
rect 505788 110312 506184 111012
rect 506884 110312 507280 111012
rect 507980 110312 508199 111012
rect 110832 110266 508199 110312
rect 88384 110078 508199 110266
rect 88384 109378 89225 110078
rect 89925 109378 90134 110078
rect 90834 109378 91043 110078
rect 91743 109378 91952 110078
rect 92652 109378 92861 110078
rect 93561 109378 93770 110078
rect 94470 109378 94679 110078
rect 95379 109378 95588 110078
rect 96288 109378 96497 110078
rect 97197 109378 97406 110078
rect 98106 109378 98315 110078
rect 99015 109378 99224 110078
rect 99924 109378 100133 110078
rect 100833 109378 101042 110078
rect 101742 109378 101951 110078
rect 102651 109378 102860 110078
rect 103560 109378 103769 110078
rect 104469 109378 104678 110078
rect 105378 109378 105587 110078
rect 106287 109378 106496 110078
rect 107196 109378 107405 110078
rect 108105 109378 108314 110078
rect 109014 109378 109223 110078
rect 109923 109378 110132 110078
rect 110832 109861 508199 110078
rect 110832 109378 482072 109861
rect 88384 109190 482072 109378
rect 88384 108490 89225 109190
rect 89925 108490 90134 109190
rect 90834 108490 91043 109190
rect 91743 108490 91952 109190
rect 92652 108490 92861 109190
rect 93561 108490 93770 109190
rect 94470 108490 94679 109190
rect 95379 108490 95588 109190
rect 96288 108490 96497 109190
rect 97197 108490 97406 109190
rect 98106 108490 98315 109190
rect 99015 108490 99224 109190
rect 99924 108490 100133 109190
rect 100833 108490 101042 109190
rect 101742 108490 101951 109190
rect 102651 108490 102860 109190
rect 103560 108490 103769 109190
rect 104469 108490 104678 109190
rect 105378 108490 105587 109190
rect 106287 108490 106496 109190
rect 107196 108490 107405 109190
rect 108105 108490 108314 109190
rect 109014 108490 109223 109190
rect 109923 108490 110132 109190
rect 110832 109161 482072 109190
rect 482772 109161 483168 109861
rect 483868 109161 484264 109861
rect 484964 109161 485360 109861
rect 486060 109161 486456 109861
rect 487156 109161 487552 109861
rect 488252 109161 488648 109861
rect 489348 109161 489744 109861
rect 490444 109161 490840 109861
rect 491540 109161 491936 109861
rect 492636 109161 493032 109861
rect 493732 109161 494128 109861
rect 494828 109161 495224 109861
rect 495924 109161 496320 109861
rect 497020 109161 497416 109861
rect 498116 109161 498512 109861
rect 499212 109161 499608 109861
rect 500308 109161 500704 109861
rect 501404 109161 501800 109861
rect 502500 109161 502896 109861
rect 503596 109161 503992 109861
rect 504692 109161 505088 109861
rect 505788 109161 506184 109861
rect 506884 109161 507280 109861
rect 507980 109161 508199 109861
rect 110832 108710 508199 109161
rect 110832 108490 482072 108710
rect 88384 108302 482072 108490
rect 88384 107602 89225 108302
rect 89925 107602 90134 108302
rect 90834 107602 91043 108302
rect 91743 107602 91952 108302
rect 92652 107602 92861 108302
rect 93561 107602 93770 108302
rect 94470 107602 94679 108302
rect 95379 107602 95588 108302
rect 96288 107602 96497 108302
rect 97197 107602 97406 108302
rect 98106 107602 98315 108302
rect 99015 107602 99224 108302
rect 99924 107602 100133 108302
rect 100833 107602 101042 108302
rect 101742 107602 101951 108302
rect 102651 107602 102860 108302
rect 103560 107602 103769 108302
rect 104469 107602 104678 108302
rect 105378 107602 105587 108302
rect 106287 107602 106496 108302
rect 107196 107602 107405 108302
rect 108105 107602 108314 108302
rect 109014 107602 109223 108302
rect 109923 107602 110132 108302
rect 110832 108010 482072 108302
rect 482772 108010 483168 108710
rect 483868 108010 484264 108710
rect 484964 108010 485360 108710
rect 486060 108010 486456 108710
rect 487156 108010 487552 108710
rect 488252 108010 488648 108710
rect 489348 108010 489744 108710
rect 490444 108010 490840 108710
rect 491540 108010 491936 108710
rect 492636 108010 493032 108710
rect 493732 108010 494128 108710
rect 494828 108010 495224 108710
rect 495924 108010 496320 108710
rect 497020 108010 497416 108710
rect 498116 108010 498512 108710
rect 499212 108010 499608 108710
rect 500308 108010 500704 108710
rect 501404 108010 501800 108710
rect 502500 108010 502896 108710
rect 503596 108010 503992 108710
rect 504692 108010 505088 108710
rect 505788 108010 506184 108710
rect 506884 108010 507280 108710
rect 507980 108010 508199 108710
rect 110832 107602 508199 108010
rect 88384 107559 508199 107602
rect 88384 107414 482072 107559
rect 88384 106714 89225 107414
rect 89925 106714 90134 107414
rect 90834 106714 91043 107414
rect 91743 106714 91952 107414
rect 92652 106714 92861 107414
rect 93561 106714 93770 107414
rect 94470 106714 94679 107414
rect 95379 106714 95588 107414
rect 96288 106714 96497 107414
rect 97197 106714 97406 107414
rect 98106 106714 98315 107414
rect 99015 106714 99224 107414
rect 99924 106714 100133 107414
rect 100833 106714 101042 107414
rect 101742 106714 101951 107414
rect 102651 106714 102860 107414
rect 103560 106714 103769 107414
rect 104469 106714 104678 107414
rect 105378 106714 105587 107414
rect 106287 106714 106496 107414
rect 107196 106714 107405 107414
rect 108105 106714 108314 107414
rect 109014 106714 109223 107414
rect 109923 106714 110132 107414
rect 110832 106859 482072 107414
rect 482772 106859 483168 107559
rect 483868 106859 484264 107559
rect 484964 106859 485360 107559
rect 486060 106859 486456 107559
rect 487156 106859 487552 107559
rect 488252 106859 488648 107559
rect 489348 106859 489744 107559
rect 490444 106859 490840 107559
rect 491540 106859 491936 107559
rect 492636 106859 493032 107559
rect 493732 106859 494128 107559
rect 494828 106859 495224 107559
rect 495924 106859 496320 107559
rect 497020 106859 497416 107559
rect 498116 106859 498512 107559
rect 499212 106859 499608 107559
rect 500308 106859 500704 107559
rect 501404 106859 501800 107559
rect 502500 106859 502896 107559
rect 503596 106859 503992 107559
rect 504692 106859 505088 107559
rect 505788 106859 506184 107559
rect 506884 106859 507280 107559
rect 507980 106859 508199 107559
rect 110832 106714 508199 106859
rect 88384 106526 508199 106714
rect 88384 105826 89225 106526
rect 89925 105826 90134 106526
rect 90834 105826 91043 106526
rect 91743 105826 91952 106526
rect 92652 105826 92861 106526
rect 93561 105826 93770 106526
rect 94470 105826 94679 106526
rect 95379 105826 95588 106526
rect 96288 105826 96497 106526
rect 97197 105826 97406 106526
rect 98106 105826 98315 106526
rect 99015 105826 99224 106526
rect 99924 105826 100133 106526
rect 100833 105826 101042 106526
rect 101742 105826 101951 106526
rect 102651 105826 102860 106526
rect 103560 105826 103769 106526
rect 104469 105826 104678 106526
rect 105378 105826 105587 106526
rect 106287 105826 106496 106526
rect 107196 105826 107405 106526
rect 108105 105826 108314 106526
rect 109014 105826 109223 106526
rect 109923 105826 110132 106526
rect 110832 106408 508199 106526
rect 110832 105826 482072 106408
rect 88384 105708 482072 105826
rect 482772 105708 483168 106408
rect 483868 105708 484264 106408
rect 484964 105708 485360 106408
rect 486060 105708 486456 106408
rect 487156 105708 487552 106408
rect 488252 105708 488648 106408
rect 489348 105708 489744 106408
rect 490444 105708 490840 106408
rect 491540 105708 491936 106408
rect 492636 105708 493032 106408
rect 493732 105708 494128 106408
rect 494828 105708 495224 106408
rect 495924 105708 496320 106408
rect 497020 105708 497416 106408
rect 498116 105708 498512 106408
rect 499212 105708 499608 106408
rect 500308 105708 500704 106408
rect 501404 105708 501800 106408
rect 502500 105708 502896 106408
rect 503596 105708 503992 106408
rect 504692 105708 505088 106408
rect 505788 105708 506184 106408
rect 506884 105708 507280 106408
rect 507980 105708 508199 106408
rect 88384 105638 508199 105708
rect 88384 104938 89225 105638
rect 89925 104938 90134 105638
rect 90834 104938 91043 105638
rect 91743 104938 91952 105638
rect 92652 104938 92861 105638
rect 93561 104938 93770 105638
rect 94470 104938 94679 105638
rect 95379 104938 95588 105638
rect 96288 104938 96497 105638
rect 97197 104938 97406 105638
rect 98106 104938 98315 105638
rect 99015 104938 99224 105638
rect 99924 104938 100133 105638
rect 100833 104938 101042 105638
rect 101742 104938 101951 105638
rect 102651 104938 102860 105638
rect 103560 104938 103769 105638
rect 104469 104938 104678 105638
rect 105378 104938 105587 105638
rect 106287 104938 106496 105638
rect 107196 104938 107405 105638
rect 108105 104938 108314 105638
rect 109014 104938 109223 105638
rect 109923 104938 110132 105638
rect 110832 105257 508199 105638
rect 110832 104938 482072 105257
rect 88384 104750 482072 104938
rect 88384 104050 89225 104750
rect 89925 104050 90134 104750
rect 90834 104050 91043 104750
rect 91743 104050 91952 104750
rect 92652 104050 92861 104750
rect 93561 104050 93770 104750
rect 94470 104050 94679 104750
rect 95379 104050 95588 104750
rect 96288 104050 96497 104750
rect 97197 104050 97406 104750
rect 98106 104050 98315 104750
rect 99015 104050 99224 104750
rect 99924 104050 100133 104750
rect 100833 104050 101042 104750
rect 101742 104050 101951 104750
rect 102651 104050 102860 104750
rect 103560 104050 103769 104750
rect 104469 104050 104678 104750
rect 105378 104050 105587 104750
rect 106287 104050 106496 104750
rect 107196 104050 107405 104750
rect 108105 104050 108314 104750
rect 109014 104050 109223 104750
rect 109923 104050 110132 104750
rect 110832 104557 482072 104750
rect 482772 104557 483168 105257
rect 483868 104557 484264 105257
rect 484964 104557 485360 105257
rect 486060 104557 486456 105257
rect 487156 104557 487552 105257
rect 488252 104557 488648 105257
rect 489348 104557 489744 105257
rect 490444 104557 490840 105257
rect 491540 104557 491936 105257
rect 492636 104557 493032 105257
rect 493732 104557 494128 105257
rect 494828 104557 495224 105257
rect 495924 104557 496320 105257
rect 497020 104557 497416 105257
rect 498116 104557 498512 105257
rect 499212 104557 499608 105257
rect 500308 104557 500704 105257
rect 501404 104557 501800 105257
rect 502500 104557 502896 105257
rect 503596 104557 503992 105257
rect 504692 104557 505088 105257
rect 505788 104557 506184 105257
rect 506884 104557 507280 105257
rect 507980 104557 508199 105257
rect 110832 104106 508199 104557
rect 110832 104050 482072 104106
rect 88384 103862 482072 104050
rect 88384 103162 89225 103862
rect 89925 103162 90134 103862
rect 90834 103162 91043 103862
rect 91743 103162 91952 103862
rect 92652 103162 92861 103862
rect 93561 103162 93770 103862
rect 94470 103162 94679 103862
rect 95379 103162 95588 103862
rect 96288 103162 96497 103862
rect 97197 103162 97406 103862
rect 98106 103162 98315 103862
rect 99015 103162 99224 103862
rect 99924 103162 100133 103862
rect 100833 103162 101042 103862
rect 101742 103162 101951 103862
rect 102651 103162 102860 103862
rect 103560 103162 103769 103862
rect 104469 103162 104678 103862
rect 105378 103162 105587 103862
rect 106287 103162 106496 103862
rect 107196 103162 107405 103862
rect 108105 103162 108314 103862
rect 109014 103162 109223 103862
rect 109923 103162 110132 103862
rect 110832 103406 482072 103862
rect 482772 103406 483168 104106
rect 483868 103406 484264 104106
rect 484964 103406 485360 104106
rect 486060 103406 486456 104106
rect 487156 103406 487552 104106
rect 488252 103406 488648 104106
rect 489348 103406 489744 104106
rect 490444 103406 490840 104106
rect 491540 103406 491936 104106
rect 492636 103406 493032 104106
rect 493732 103406 494128 104106
rect 494828 103406 495224 104106
rect 495924 103406 496320 104106
rect 497020 103406 497416 104106
rect 498116 103406 498512 104106
rect 499212 103406 499608 104106
rect 500308 103406 500704 104106
rect 501404 103406 501800 104106
rect 502500 103406 502896 104106
rect 503596 103406 503992 104106
rect 504692 103406 505088 104106
rect 505788 103406 506184 104106
rect 506884 103406 507280 104106
rect 507980 103406 508199 104106
rect 110832 103162 508199 103406
rect 88384 102974 508199 103162
rect 88384 102274 89225 102974
rect 89925 102274 90134 102974
rect 90834 102274 91043 102974
rect 91743 102274 91952 102974
rect 92652 102274 92861 102974
rect 93561 102274 93770 102974
rect 94470 102274 94679 102974
rect 95379 102274 95588 102974
rect 96288 102274 96497 102974
rect 97197 102274 97406 102974
rect 98106 102274 98315 102974
rect 99015 102274 99224 102974
rect 99924 102274 100133 102974
rect 100833 102274 101042 102974
rect 101742 102274 101951 102974
rect 102651 102274 102860 102974
rect 103560 102274 103769 102974
rect 104469 102274 104678 102974
rect 105378 102274 105587 102974
rect 106287 102274 106496 102974
rect 107196 102274 107405 102974
rect 108105 102274 108314 102974
rect 109014 102274 109223 102974
rect 109923 102274 110132 102974
rect 110832 102955 508199 102974
rect 110832 102596 482072 102955
rect 110832 102274 111541 102596
rect 88384 102086 111541 102274
rect 88384 101386 89225 102086
rect 89925 101386 90134 102086
rect 90834 101386 91043 102086
rect 91743 101386 91952 102086
rect 92652 101386 92861 102086
rect 93561 101386 93770 102086
rect 94470 101386 94679 102086
rect 95379 101386 95588 102086
rect 96288 101386 96497 102086
rect 97197 101386 97406 102086
rect 98106 101386 98315 102086
rect 99015 101386 99224 102086
rect 99924 101386 100133 102086
rect 100833 101386 101042 102086
rect 101742 101386 101951 102086
rect 102651 101386 102860 102086
rect 103560 101386 103769 102086
rect 104469 101386 104678 102086
rect 105378 101386 105587 102086
rect 106287 101386 106496 102086
rect 107196 101386 107405 102086
rect 108105 101386 108314 102086
rect 109014 101386 109223 102086
rect 109923 101386 110132 102086
rect 110832 101386 111541 102086
rect 88384 101198 111541 101386
rect 88384 100498 89225 101198
rect 89925 100498 90134 101198
rect 90834 100498 91043 101198
rect 91743 100498 91952 101198
rect 92652 100498 92861 101198
rect 93561 100498 93770 101198
rect 94470 100498 94679 101198
rect 95379 100498 95588 101198
rect 96288 100498 96497 101198
rect 97197 100498 97406 101198
rect 98106 100498 98315 101198
rect 99015 100498 99224 101198
rect 99924 100498 100133 101198
rect 100833 100498 101042 101198
rect 101742 100498 101951 101198
rect 102651 100498 102860 101198
rect 103560 100498 103769 101198
rect 104469 100498 104678 101198
rect 105378 100498 105587 101198
rect 106287 100498 106496 101198
rect 107196 100498 107405 101198
rect 108105 100498 108314 101198
rect 109014 100498 109223 101198
rect 109923 100498 110132 101198
rect 110832 100498 111541 101198
rect 88384 100310 111541 100498
rect 88384 99610 89225 100310
rect 89925 99610 90134 100310
rect 90834 99610 91043 100310
rect 91743 99610 91952 100310
rect 92652 99610 92861 100310
rect 93561 99610 93770 100310
rect 94470 99610 94679 100310
rect 95379 99610 95588 100310
rect 96288 99610 96497 100310
rect 97197 99610 97406 100310
rect 98106 99610 98315 100310
rect 99015 99610 99224 100310
rect 99924 99610 100133 100310
rect 100833 99610 101042 100310
rect 101742 99610 101951 100310
rect 102651 99610 102860 100310
rect 103560 99610 103769 100310
rect 104469 99610 104678 100310
rect 105378 99610 105587 100310
rect 106287 99610 106496 100310
rect 107196 99610 107405 100310
rect 108105 99610 108314 100310
rect 109014 99610 109223 100310
rect 109923 99610 110132 100310
rect 110832 99610 111541 100310
rect 88384 99422 111541 99610
rect 481670 102255 482072 102596
rect 482772 102255 483168 102955
rect 483868 102255 484264 102955
rect 484964 102255 485360 102955
rect 486060 102255 486456 102955
rect 487156 102255 487552 102955
rect 488252 102255 488648 102955
rect 489348 102255 489744 102955
rect 490444 102255 490840 102955
rect 491540 102255 491936 102955
rect 492636 102255 493032 102955
rect 493732 102255 494128 102955
rect 494828 102255 495224 102955
rect 495924 102255 496320 102955
rect 497020 102255 497416 102955
rect 498116 102255 498512 102955
rect 499212 102255 499608 102955
rect 500308 102255 500704 102955
rect 501404 102255 501800 102955
rect 502500 102255 502896 102955
rect 503596 102255 503992 102955
rect 504692 102255 505088 102955
rect 505788 102255 506184 102955
rect 506884 102255 507280 102955
rect 507980 102255 508199 102955
rect 481670 101804 508199 102255
rect 481670 101104 482072 101804
rect 482772 101104 483168 101804
rect 483868 101104 484264 101804
rect 484964 101104 485360 101804
rect 486060 101104 486456 101804
rect 487156 101104 487552 101804
rect 488252 101104 488648 101804
rect 489348 101104 489744 101804
rect 490444 101104 490840 101804
rect 491540 101104 491936 101804
rect 492636 101104 493032 101804
rect 493732 101104 494128 101804
rect 494828 101104 495224 101804
rect 495924 101104 496320 101804
rect 497020 101104 497416 101804
rect 498116 101104 498512 101804
rect 499212 101104 499608 101804
rect 500308 101104 500704 101804
rect 501404 101104 501800 101804
rect 502500 101104 502896 101804
rect 503596 101104 503992 101804
rect 504692 101104 505088 101804
rect 505788 101104 506184 101804
rect 506884 101104 507280 101804
rect 507980 101104 508199 101804
rect 481670 100653 508199 101104
rect 481670 99953 482072 100653
rect 482772 99953 483168 100653
rect 483868 99953 484264 100653
rect 484964 99953 485360 100653
rect 486060 99953 486456 100653
rect 487156 99953 487552 100653
rect 488252 99953 488648 100653
rect 489348 99953 489744 100653
rect 490444 99953 490840 100653
rect 491540 99953 491936 100653
rect 492636 99953 493032 100653
rect 493732 99953 494128 100653
rect 494828 99953 495224 100653
rect 495924 99953 496320 100653
rect 497020 99953 497416 100653
rect 498116 99953 498512 100653
rect 499212 99953 499608 100653
rect 500308 99953 500704 100653
rect 501404 99953 501800 100653
rect 502500 99953 502896 100653
rect 503596 99953 503992 100653
rect 504692 99953 505088 100653
rect 505788 99953 506184 100653
rect 506884 99953 507280 100653
rect 507980 99953 508199 100653
rect 481670 99723 508199 99953
rect 481670 99532 507195 99723
rect 88384 98722 89225 99422
rect 89925 98722 90134 99422
rect 90834 98722 91043 99422
rect 91743 98722 91952 99422
rect 92652 98722 92861 99422
rect 93561 98722 93770 99422
rect 94470 98722 94679 99422
rect 95379 98722 95588 99422
rect 96288 98722 96497 99422
rect 97197 98722 97406 99422
rect 98106 98722 98315 99422
rect 99015 98722 99224 99422
rect 99924 98722 100133 99422
rect 100833 98722 101042 99422
rect 101742 98722 101951 99422
rect 102651 98722 102860 99422
rect 103560 98722 103769 99422
rect 104469 98722 104678 99422
rect 105378 98722 105587 99422
rect 106287 98722 106496 99422
rect 107196 98722 107405 99422
rect 108105 98722 108314 99422
rect 109014 98722 109223 99422
rect 109923 98722 110132 99422
rect 110832 98722 111541 99422
rect 88384 98042 111541 98722
<< via3 >>
rect 87948 510096 88648 510796
rect 88929 510096 89629 510796
rect 89910 510096 90610 510796
rect 90891 510096 91591 510796
rect 91872 510096 92572 510796
rect 92853 510096 93553 510796
rect 93834 510096 94534 510796
rect 94815 510096 95515 510796
rect 95796 510096 96496 510796
rect 96777 510096 97477 510796
rect 97758 510096 98458 510796
rect 98739 510096 99439 510796
rect 99720 510096 100420 510796
rect 100701 510096 101401 510796
rect 101682 510096 102382 510796
rect 102663 510096 103363 510796
rect 103644 510096 104344 510796
rect 104625 510096 105325 510796
rect 105606 510096 106306 510796
rect 106587 510096 107287 510796
rect 107568 510096 108268 510796
rect 108549 510096 109249 510796
rect 109530 510096 110230 510796
rect 110511 510096 111211 510796
rect 111492 510096 112192 510796
rect 87948 509076 88648 509776
rect 88929 509076 89629 509776
rect 89910 509076 90610 509776
rect 90891 509076 91591 509776
rect 91872 509076 92572 509776
rect 92853 509076 93553 509776
rect 93834 509076 94534 509776
rect 94815 509076 95515 509776
rect 95796 509076 96496 509776
rect 96777 509076 97477 509776
rect 97758 509076 98458 509776
rect 98739 509076 99439 509776
rect 99720 509076 100420 509776
rect 100701 509076 101401 509776
rect 101682 509076 102382 509776
rect 102663 509076 103363 509776
rect 103644 509076 104344 509776
rect 104625 509076 105325 509776
rect 105606 509076 106306 509776
rect 106587 509076 107287 509776
rect 107568 509076 108268 509776
rect 108549 509076 109249 509776
rect 109530 509076 110230 509776
rect 110511 509076 111211 509776
rect 111492 509076 112192 509776
rect 87948 508056 88648 508756
rect 88929 508056 89629 508756
rect 89910 508056 90610 508756
rect 90891 508056 91591 508756
rect 91872 508056 92572 508756
rect 92853 508056 93553 508756
rect 93834 508056 94534 508756
rect 94815 508056 95515 508756
rect 95796 508056 96496 508756
rect 96777 508056 97477 508756
rect 97758 508056 98458 508756
rect 98739 508056 99439 508756
rect 99720 508056 100420 508756
rect 100701 508056 101401 508756
rect 101682 508056 102382 508756
rect 102663 508056 103363 508756
rect 103644 508056 104344 508756
rect 104625 508056 105325 508756
rect 105606 508056 106306 508756
rect 106587 508056 107287 508756
rect 107568 508056 108268 508756
rect 108549 508056 109249 508756
rect 109530 508056 110230 508756
rect 110511 508056 111211 508756
rect 111492 508056 112192 508756
rect 87948 507036 88648 507736
rect 88929 507036 89629 507736
rect 89910 507036 90610 507736
rect 90891 507036 91591 507736
rect 91872 507036 92572 507736
rect 92853 507036 93553 507736
rect 93834 507036 94534 507736
rect 94815 507036 95515 507736
rect 95796 507036 96496 507736
rect 96777 507036 97477 507736
rect 97758 507036 98458 507736
rect 98739 507036 99439 507736
rect 99720 507036 100420 507736
rect 100701 507036 101401 507736
rect 101682 507036 102382 507736
rect 102663 507036 103363 507736
rect 103644 507036 104344 507736
rect 104625 507036 105325 507736
rect 105606 507036 106306 507736
rect 106587 507036 107287 507736
rect 107568 507036 108268 507736
rect 108549 507036 109249 507736
rect 109530 507036 110230 507736
rect 110511 507036 111211 507736
rect 111492 507036 112192 507736
rect 87948 506016 88648 506716
rect 88929 506016 89629 506716
rect 89910 506016 90610 506716
rect 90891 506016 91591 506716
rect 91872 506016 92572 506716
rect 92853 506016 93553 506716
rect 93834 506016 94534 506716
rect 94815 506016 95515 506716
rect 95796 506016 96496 506716
rect 96777 506016 97477 506716
rect 97758 506016 98458 506716
rect 98739 506016 99439 506716
rect 99720 506016 100420 506716
rect 100701 506016 101401 506716
rect 101682 506016 102382 506716
rect 102663 506016 103363 506716
rect 103644 506016 104344 506716
rect 104625 506016 105325 506716
rect 105606 506016 106306 506716
rect 106587 506016 107287 506716
rect 107568 506016 108268 506716
rect 108549 506016 109249 506716
rect 109530 506016 110230 506716
rect 110511 506016 111211 506716
rect 111492 506016 112192 506716
rect 482569 507375 483269 508075
rect 483896 507375 484596 508075
rect 485223 507375 485923 508075
rect 486550 507375 487250 508075
rect 487877 507375 488577 508075
rect 489204 507375 489904 508075
rect 490531 507375 491231 508075
rect 491858 507375 492558 508075
rect 493185 507375 493885 508075
rect 494512 507375 495212 508075
rect 495839 507375 496539 508075
rect 497166 507375 497866 508075
rect 498493 507375 499193 508075
rect 499820 507375 500520 508075
rect 501147 507375 501847 508075
rect 502474 507375 503174 508075
rect 503801 507375 504501 508075
rect 505128 507375 505828 508075
rect 506455 507375 507155 508075
rect 482569 506048 483269 506748
rect 483896 506048 484596 506748
rect 485223 506048 485923 506748
rect 486550 506048 487250 506748
rect 487877 506048 488577 506748
rect 489204 506048 489904 506748
rect 490531 506048 491231 506748
rect 491858 506048 492558 506748
rect 493185 506048 493885 506748
rect 494512 506048 495212 506748
rect 495839 506048 496539 506748
rect 497166 506048 497866 506748
rect 498493 506048 499193 506748
rect 499820 506048 500520 506748
rect 501147 506048 501847 506748
rect 502474 506048 503174 506748
rect 503801 506048 504501 506748
rect 505128 506048 505828 506748
rect 506455 506048 507155 506748
rect 87948 504996 88648 505696
rect 88929 504996 89629 505696
rect 89910 504996 90610 505696
rect 90891 504996 91591 505696
rect 91872 504996 92572 505696
rect 92853 504996 93553 505696
rect 93834 504996 94534 505696
rect 94815 504996 95515 505696
rect 95796 504996 96496 505696
rect 96777 504996 97477 505696
rect 97758 504996 98458 505696
rect 98739 504996 99439 505696
rect 99720 504996 100420 505696
rect 100701 504996 101401 505696
rect 101682 504996 102382 505696
rect 102663 504996 103363 505696
rect 103644 504996 104344 505696
rect 104625 504996 105325 505696
rect 105606 504996 106306 505696
rect 106587 504996 107287 505696
rect 107568 504996 108268 505696
rect 108549 504996 109249 505696
rect 109530 504996 110230 505696
rect 110511 504996 111211 505696
rect 111492 504996 112192 505696
rect 482569 504721 483269 505421
rect 483896 504721 484596 505421
rect 485223 504721 485923 505421
rect 486550 504721 487250 505421
rect 487877 504721 488577 505421
rect 489204 504721 489904 505421
rect 490531 504721 491231 505421
rect 491858 504721 492558 505421
rect 493185 504721 493885 505421
rect 494512 504721 495212 505421
rect 495839 504721 496539 505421
rect 497166 504721 497866 505421
rect 498493 504721 499193 505421
rect 499820 504721 500520 505421
rect 501147 504721 501847 505421
rect 502474 504721 503174 505421
rect 503801 504721 504501 505421
rect 505128 504721 505828 505421
rect 506455 504721 507155 505421
rect 87948 503976 88648 504676
rect 88929 503976 89629 504676
rect 89910 503976 90610 504676
rect 90891 503976 91591 504676
rect 91872 503976 92572 504676
rect 92853 503976 93553 504676
rect 93834 503976 94534 504676
rect 94815 503976 95515 504676
rect 95796 503976 96496 504676
rect 96777 503976 97477 504676
rect 97758 503976 98458 504676
rect 98739 503976 99439 504676
rect 99720 503976 100420 504676
rect 100701 503976 101401 504676
rect 101682 503976 102382 504676
rect 102663 503976 103363 504676
rect 103644 503976 104344 504676
rect 104625 503976 105325 504676
rect 105606 503976 106306 504676
rect 106587 503976 107287 504676
rect 107568 503976 108268 504676
rect 108549 503976 109249 504676
rect 109530 503976 110230 504676
rect 110511 503976 111211 504676
rect 111492 503976 112192 504676
rect 87948 502956 88648 503656
rect 88929 502956 89629 503656
rect 89910 502956 90610 503656
rect 90891 502956 91591 503656
rect 91872 502956 92572 503656
rect 92853 502956 93553 503656
rect 93834 502956 94534 503656
rect 94815 502956 95515 503656
rect 95796 502956 96496 503656
rect 96777 502956 97477 503656
rect 97758 502956 98458 503656
rect 98739 502956 99439 503656
rect 99720 502956 100420 503656
rect 100701 502956 101401 503656
rect 101682 502956 102382 503656
rect 102663 502956 103363 503656
rect 103644 502956 104344 503656
rect 104625 502956 105325 503656
rect 105606 502956 106306 503656
rect 106587 502956 107287 503656
rect 107568 502956 108268 503656
rect 108549 502956 109249 503656
rect 109530 502956 110230 503656
rect 110511 502956 111211 503656
rect 111492 502956 112192 503656
rect 482569 503394 483269 504094
rect 483896 503394 484596 504094
rect 485223 503394 485923 504094
rect 486550 503394 487250 504094
rect 487877 503394 488577 504094
rect 489204 503394 489904 504094
rect 490531 503394 491231 504094
rect 491858 503394 492558 504094
rect 493185 503394 493885 504094
rect 494512 503394 495212 504094
rect 495839 503394 496539 504094
rect 497166 503394 497866 504094
rect 498493 503394 499193 504094
rect 499820 503394 500520 504094
rect 501147 503394 501847 504094
rect 502474 503394 503174 504094
rect 503801 503394 504501 504094
rect 505128 503394 505828 504094
rect 506455 503394 507155 504094
rect 87948 501936 88648 502636
rect 88929 501936 89629 502636
rect 89910 501936 90610 502636
rect 90891 501936 91591 502636
rect 91872 501936 92572 502636
rect 92853 501936 93553 502636
rect 93834 501936 94534 502636
rect 94815 501936 95515 502636
rect 95796 501936 96496 502636
rect 96777 501936 97477 502636
rect 97758 501936 98458 502636
rect 98739 501936 99439 502636
rect 99720 501936 100420 502636
rect 100701 501936 101401 502636
rect 101682 501936 102382 502636
rect 102663 501936 103363 502636
rect 103644 501936 104344 502636
rect 104625 501936 105325 502636
rect 105606 501936 106306 502636
rect 106587 501936 107287 502636
rect 107568 501936 108268 502636
rect 108549 501936 109249 502636
rect 109530 501936 110230 502636
rect 110511 501936 111211 502636
rect 111492 501936 112192 502636
rect 482569 502067 483269 502767
rect 483896 502067 484596 502767
rect 485223 502067 485923 502767
rect 486550 502067 487250 502767
rect 487877 502067 488577 502767
rect 489204 502067 489904 502767
rect 490531 502067 491231 502767
rect 491858 502067 492558 502767
rect 493185 502067 493885 502767
rect 494512 502067 495212 502767
rect 495839 502067 496539 502767
rect 497166 502067 497866 502767
rect 498493 502067 499193 502767
rect 499820 502067 500520 502767
rect 501147 502067 501847 502767
rect 502474 502067 503174 502767
rect 503801 502067 504501 502767
rect 505128 502067 505828 502767
rect 506455 502067 507155 502767
rect 87948 500916 88648 501616
rect 88929 500916 89629 501616
rect 89910 500916 90610 501616
rect 90891 500916 91591 501616
rect 91872 500916 92572 501616
rect 92853 500916 93553 501616
rect 93834 500916 94534 501616
rect 94815 500916 95515 501616
rect 95796 500916 96496 501616
rect 96777 500916 97477 501616
rect 97758 500916 98458 501616
rect 98739 500916 99439 501616
rect 99720 500916 100420 501616
rect 100701 500916 101401 501616
rect 101682 500916 102382 501616
rect 102663 500916 103363 501616
rect 103644 500916 104344 501616
rect 104625 500916 105325 501616
rect 105606 500916 106306 501616
rect 106587 500916 107287 501616
rect 107568 500916 108268 501616
rect 108549 500916 109249 501616
rect 109530 500916 110230 501616
rect 110511 500916 111211 501616
rect 111492 500916 112192 501616
rect 482569 500740 483269 501440
rect 483896 500740 484596 501440
rect 485223 500740 485923 501440
rect 486550 500740 487250 501440
rect 487877 500740 488577 501440
rect 489204 500740 489904 501440
rect 490531 500740 491231 501440
rect 491858 500740 492558 501440
rect 493185 500740 493885 501440
rect 494512 500740 495212 501440
rect 495839 500740 496539 501440
rect 497166 500740 497866 501440
rect 498493 500740 499193 501440
rect 499820 500740 500520 501440
rect 501147 500740 501847 501440
rect 502474 500740 503174 501440
rect 503801 500740 504501 501440
rect 505128 500740 505828 501440
rect 506455 500740 507155 501440
rect 87948 499896 88648 500596
rect 88929 499896 89629 500596
rect 89910 499896 90610 500596
rect 90891 499896 91591 500596
rect 91872 499896 92572 500596
rect 92853 499896 93553 500596
rect 93834 499896 94534 500596
rect 94815 499896 95515 500596
rect 95796 499896 96496 500596
rect 96777 499896 97477 500596
rect 97758 499896 98458 500596
rect 98739 499896 99439 500596
rect 99720 499896 100420 500596
rect 100701 499896 101401 500596
rect 101682 499896 102382 500596
rect 102663 499896 103363 500596
rect 103644 499896 104344 500596
rect 104625 499896 105325 500596
rect 105606 499896 106306 500596
rect 106587 499896 107287 500596
rect 107568 499896 108268 500596
rect 108549 499896 109249 500596
rect 109530 499896 110230 500596
rect 110511 499896 111211 500596
rect 111492 499896 112192 500596
rect 87948 498876 88648 499576
rect 88929 498876 89629 499576
rect 89910 498876 90610 499576
rect 90891 498876 91591 499576
rect 91872 498876 92572 499576
rect 92853 498876 93553 499576
rect 93834 498876 94534 499576
rect 94815 498876 95515 499576
rect 95796 498876 96496 499576
rect 96777 498876 97477 499576
rect 97758 498876 98458 499576
rect 98739 498876 99439 499576
rect 99720 498876 100420 499576
rect 100701 498876 101401 499576
rect 101682 498876 102382 499576
rect 102663 498876 103363 499576
rect 103644 498876 104344 499576
rect 104625 498876 105325 499576
rect 105606 498876 106306 499576
rect 106587 498876 107287 499576
rect 107568 498876 108268 499576
rect 108549 498876 109249 499576
rect 109530 498876 110230 499576
rect 110511 498876 111211 499576
rect 111492 498876 112192 499576
rect 482569 499413 483269 500113
rect 483896 499413 484596 500113
rect 485223 499413 485923 500113
rect 486550 499413 487250 500113
rect 487877 499413 488577 500113
rect 489204 499413 489904 500113
rect 490531 499413 491231 500113
rect 491858 499413 492558 500113
rect 493185 499413 493885 500113
rect 494512 499413 495212 500113
rect 495839 499413 496539 500113
rect 497166 499413 497866 500113
rect 498493 499413 499193 500113
rect 499820 499413 500520 500113
rect 501147 499413 501847 500113
rect 502474 499413 503174 500113
rect 503801 499413 504501 500113
rect 505128 499413 505828 500113
rect 506455 499413 507155 500113
rect 87948 497856 88648 498556
rect 88929 497856 89629 498556
rect 89910 497856 90610 498556
rect 90891 497856 91591 498556
rect 91872 497856 92572 498556
rect 92853 497856 93553 498556
rect 93834 497856 94534 498556
rect 94815 497856 95515 498556
rect 95796 497856 96496 498556
rect 96777 497856 97477 498556
rect 97758 497856 98458 498556
rect 98739 497856 99439 498556
rect 99720 497856 100420 498556
rect 100701 497856 101401 498556
rect 101682 497856 102382 498556
rect 102663 497856 103363 498556
rect 103644 497856 104344 498556
rect 104625 497856 105325 498556
rect 105606 497856 106306 498556
rect 106587 497856 107287 498556
rect 107568 497856 108268 498556
rect 108549 497856 109249 498556
rect 109530 497856 110230 498556
rect 110511 497856 111211 498556
rect 111492 497856 112192 498556
rect 482569 498086 483269 498786
rect 483896 498086 484596 498786
rect 485223 498086 485923 498786
rect 486550 498086 487250 498786
rect 487877 498086 488577 498786
rect 489204 498086 489904 498786
rect 490531 498086 491231 498786
rect 491858 498086 492558 498786
rect 493185 498086 493885 498786
rect 494512 498086 495212 498786
rect 495839 498086 496539 498786
rect 497166 498086 497866 498786
rect 498493 498086 499193 498786
rect 499820 498086 500520 498786
rect 501147 498086 501847 498786
rect 502474 498086 503174 498786
rect 503801 498086 504501 498786
rect 505128 498086 505828 498786
rect 506455 498086 507155 498786
rect 87948 496836 88648 497536
rect 88929 496836 89629 497536
rect 89910 496836 90610 497536
rect 90891 496836 91591 497536
rect 91872 496836 92572 497536
rect 92853 496836 93553 497536
rect 93834 496836 94534 497536
rect 94815 496836 95515 497536
rect 95796 496836 96496 497536
rect 96777 496836 97477 497536
rect 97758 496836 98458 497536
rect 98739 496836 99439 497536
rect 99720 496836 100420 497536
rect 100701 496836 101401 497536
rect 101682 496836 102382 497536
rect 102663 496836 103363 497536
rect 103644 496836 104344 497536
rect 104625 496836 105325 497536
rect 105606 496836 106306 497536
rect 106587 496836 107287 497536
rect 107568 496836 108268 497536
rect 108549 496836 109249 497536
rect 109530 496836 110230 497536
rect 110511 496836 111211 497536
rect 111492 496836 112192 497536
rect 482569 496759 483269 497459
rect 483896 496759 484596 497459
rect 485223 496759 485923 497459
rect 486550 496759 487250 497459
rect 487877 496759 488577 497459
rect 489204 496759 489904 497459
rect 490531 496759 491231 497459
rect 491858 496759 492558 497459
rect 493185 496759 493885 497459
rect 494512 496759 495212 497459
rect 495839 496759 496539 497459
rect 497166 496759 497866 497459
rect 498493 496759 499193 497459
rect 499820 496759 500520 497459
rect 501147 496759 501847 497459
rect 502474 496759 503174 497459
rect 503801 496759 504501 497459
rect 505128 496759 505828 497459
rect 506455 496759 507155 497459
rect 87948 495816 88648 496516
rect 88929 495816 89629 496516
rect 89910 495816 90610 496516
rect 90891 495816 91591 496516
rect 91872 495816 92572 496516
rect 92853 495816 93553 496516
rect 93834 495816 94534 496516
rect 94815 495816 95515 496516
rect 95796 495816 96496 496516
rect 96777 495816 97477 496516
rect 97758 495816 98458 496516
rect 98739 495816 99439 496516
rect 99720 495816 100420 496516
rect 100701 495816 101401 496516
rect 101682 495816 102382 496516
rect 102663 495816 103363 496516
rect 103644 495816 104344 496516
rect 104625 495816 105325 496516
rect 105606 495816 106306 496516
rect 106587 495816 107287 496516
rect 107568 495816 108268 496516
rect 108549 495816 109249 496516
rect 109530 495816 110230 496516
rect 110511 495816 111211 496516
rect 111492 495816 112192 496516
rect 87948 494796 88648 495496
rect 88929 494796 89629 495496
rect 89910 494796 90610 495496
rect 90891 494796 91591 495496
rect 91872 494796 92572 495496
rect 92853 494796 93553 495496
rect 93834 494796 94534 495496
rect 94815 494796 95515 495496
rect 95796 494796 96496 495496
rect 96777 494796 97477 495496
rect 97758 494796 98458 495496
rect 98739 494796 99439 495496
rect 99720 494796 100420 495496
rect 100701 494796 101401 495496
rect 101682 494796 102382 495496
rect 102663 494796 103363 495496
rect 103644 494796 104344 495496
rect 104625 494796 105325 495496
rect 105606 494796 106306 495496
rect 106587 494796 107287 495496
rect 107568 494796 108268 495496
rect 108549 494796 109249 495496
rect 109530 494796 110230 495496
rect 110511 494796 111211 495496
rect 111492 494796 112192 495496
rect 482569 495432 483269 496132
rect 483896 495432 484596 496132
rect 485223 495432 485923 496132
rect 486550 495432 487250 496132
rect 487877 495432 488577 496132
rect 489204 495432 489904 496132
rect 490531 495432 491231 496132
rect 491858 495432 492558 496132
rect 493185 495432 493885 496132
rect 494512 495432 495212 496132
rect 495839 495432 496539 496132
rect 497166 495432 497866 496132
rect 498493 495432 499193 496132
rect 499820 495432 500520 496132
rect 501147 495432 501847 496132
rect 502474 495432 503174 496132
rect 503801 495432 504501 496132
rect 505128 495432 505828 496132
rect 506455 495432 507155 496132
rect 87948 493776 88648 494476
rect 88929 493776 89629 494476
rect 89910 493776 90610 494476
rect 90891 493776 91591 494476
rect 91872 493776 92572 494476
rect 92853 493776 93553 494476
rect 93834 493776 94534 494476
rect 94815 493776 95515 494476
rect 95796 493776 96496 494476
rect 96777 493776 97477 494476
rect 97758 493776 98458 494476
rect 98739 493776 99439 494476
rect 99720 493776 100420 494476
rect 100701 493776 101401 494476
rect 101682 493776 102382 494476
rect 102663 493776 103363 494476
rect 103644 493776 104344 494476
rect 104625 493776 105325 494476
rect 105606 493776 106306 494476
rect 106587 493776 107287 494476
rect 107568 493776 108268 494476
rect 108549 493776 109249 494476
rect 109530 493776 110230 494476
rect 110511 493776 111211 494476
rect 111492 493776 112192 494476
rect 482569 494105 483269 494805
rect 483896 494105 484596 494805
rect 485223 494105 485923 494805
rect 486550 494105 487250 494805
rect 487877 494105 488577 494805
rect 489204 494105 489904 494805
rect 490531 494105 491231 494805
rect 491858 494105 492558 494805
rect 493185 494105 493885 494805
rect 494512 494105 495212 494805
rect 495839 494105 496539 494805
rect 497166 494105 497866 494805
rect 498493 494105 499193 494805
rect 499820 494105 500520 494805
rect 501147 494105 501847 494805
rect 502474 494105 503174 494805
rect 503801 494105 504501 494805
rect 505128 494105 505828 494805
rect 506455 494105 507155 494805
rect 87948 492756 88648 493456
rect 88929 492756 89629 493456
rect 89910 492756 90610 493456
rect 90891 492756 91591 493456
rect 91872 492756 92572 493456
rect 92853 492756 93553 493456
rect 93834 492756 94534 493456
rect 94815 492756 95515 493456
rect 95796 492756 96496 493456
rect 96777 492756 97477 493456
rect 97758 492756 98458 493456
rect 98739 492756 99439 493456
rect 99720 492756 100420 493456
rect 100701 492756 101401 493456
rect 101682 492756 102382 493456
rect 102663 492756 103363 493456
rect 103644 492756 104344 493456
rect 104625 492756 105325 493456
rect 105606 492756 106306 493456
rect 106587 492756 107287 493456
rect 107568 492756 108268 493456
rect 108549 492756 109249 493456
rect 109530 492756 110230 493456
rect 110511 492756 111211 493456
rect 111492 492756 112192 493456
rect 482569 492778 483269 493478
rect 483896 492778 484596 493478
rect 485223 492778 485923 493478
rect 486550 492778 487250 493478
rect 487877 492778 488577 493478
rect 489204 492778 489904 493478
rect 490531 492778 491231 493478
rect 491858 492778 492558 493478
rect 493185 492778 493885 493478
rect 494512 492778 495212 493478
rect 495839 492778 496539 493478
rect 497166 492778 497866 493478
rect 498493 492778 499193 493478
rect 499820 492778 500520 493478
rect 501147 492778 501847 493478
rect 502474 492778 503174 493478
rect 503801 492778 504501 493478
rect 505128 492778 505828 493478
rect 506455 492778 507155 493478
rect 87948 491736 88648 492436
rect 88929 491736 89629 492436
rect 89910 491736 90610 492436
rect 90891 491736 91591 492436
rect 91872 491736 92572 492436
rect 92853 491736 93553 492436
rect 93834 491736 94534 492436
rect 94815 491736 95515 492436
rect 95796 491736 96496 492436
rect 96777 491736 97477 492436
rect 97758 491736 98458 492436
rect 98739 491736 99439 492436
rect 99720 491736 100420 492436
rect 100701 491736 101401 492436
rect 101682 491736 102382 492436
rect 102663 491736 103363 492436
rect 103644 491736 104344 492436
rect 104625 491736 105325 492436
rect 105606 491736 106306 492436
rect 106587 491736 107287 492436
rect 107568 491736 108268 492436
rect 108549 491736 109249 492436
rect 109530 491736 110230 492436
rect 110511 491736 111211 492436
rect 111492 491736 112192 492436
rect 482569 491451 483269 492151
rect 483896 491451 484596 492151
rect 485223 491451 485923 492151
rect 486550 491451 487250 492151
rect 487877 491451 488577 492151
rect 489204 491451 489904 492151
rect 490531 491451 491231 492151
rect 491858 491451 492558 492151
rect 493185 491451 493885 492151
rect 494512 491451 495212 492151
rect 495839 491451 496539 492151
rect 497166 491451 497866 492151
rect 498493 491451 499193 492151
rect 499820 491451 500520 492151
rect 501147 491451 501847 492151
rect 502474 491451 503174 492151
rect 503801 491451 504501 492151
rect 505128 491451 505828 492151
rect 506455 491451 507155 492151
rect 87948 490716 88648 491416
rect 88929 490716 89629 491416
rect 89910 490716 90610 491416
rect 90891 490716 91591 491416
rect 91872 490716 92572 491416
rect 92853 490716 93553 491416
rect 93834 490716 94534 491416
rect 94815 490716 95515 491416
rect 95796 490716 96496 491416
rect 96777 490716 97477 491416
rect 97758 490716 98458 491416
rect 98739 490716 99439 491416
rect 99720 490716 100420 491416
rect 100701 490716 101401 491416
rect 101682 490716 102382 491416
rect 102663 490716 103363 491416
rect 103644 490716 104344 491416
rect 104625 490716 105325 491416
rect 105606 490716 106306 491416
rect 106587 490716 107287 491416
rect 107568 490716 108268 491416
rect 108549 490716 109249 491416
rect 109530 490716 110230 491416
rect 110511 490716 111211 491416
rect 111492 490716 112192 491416
rect 87948 489696 88648 490396
rect 88929 489696 89629 490396
rect 89910 489696 90610 490396
rect 90891 489696 91591 490396
rect 91872 489696 92572 490396
rect 92853 489696 93553 490396
rect 93834 489696 94534 490396
rect 94815 489696 95515 490396
rect 95796 489696 96496 490396
rect 96777 489696 97477 490396
rect 97758 489696 98458 490396
rect 98739 489696 99439 490396
rect 99720 489696 100420 490396
rect 100701 489696 101401 490396
rect 101682 489696 102382 490396
rect 102663 489696 103363 490396
rect 103644 489696 104344 490396
rect 104625 489696 105325 490396
rect 105606 489696 106306 490396
rect 106587 489696 107287 490396
rect 107568 489696 108268 490396
rect 108549 489696 109249 490396
rect 109530 489696 110230 490396
rect 110511 489696 111211 490396
rect 111492 489696 112192 490396
rect 482569 490124 483269 490824
rect 483896 490124 484596 490824
rect 485223 490124 485923 490824
rect 486550 490124 487250 490824
rect 487877 490124 488577 490824
rect 489204 490124 489904 490824
rect 490531 490124 491231 490824
rect 491858 490124 492558 490824
rect 493185 490124 493885 490824
rect 494512 490124 495212 490824
rect 495839 490124 496539 490824
rect 497166 490124 497866 490824
rect 498493 490124 499193 490824
rect 499820 490124 500520 490824
rect 501147 490124 501847 490824
rect 502474 490124 503174 490824
rect 503801 490124 504501 490824
rect 505128 490124 505828 490824
rect 506455 490124 507155 490824
rect 87948 488676 88648 489376
rect 88929 488676 89629 489376
rect 89910 488676 90610 489376
rect 90891 488676 91591 489376
rect 91872 488676 92572 489376
rect 92853 488676 93553 489376
rect 93834 488676 94534 489376
rect 94815 488676 95515 489376
rect 95796 488676 96496 489376
rect 96777 488676 97477 489376
rect 97758 488676 98458 489376
rect 98739 488676 99439 489376
rect 99720 488676 100420 489376
rect 100701 488676 101401 489376
rect 101682 488676 102382 489376
rect 102663 488676 103363 489376
rect 103644 488676 104344 489376
rect 104625 488676 105325 489376
rect 105606 488676 106306 489376
rect 106587 488676 107287 489376
rect 107568 488676 108268 489376
rect 108549 488676 109249 489376
rect 109530 488676 110230 489376
rect 110511 488676 111211 489376
rect 111492 488676 112192 489376
rect 482569 488797 483269 489497
rect 483896 488797 484596 489497
rect 485223 488797 485923 489497
rect 486550 488797 487250 489497
rect 487877 488797 488577 489497
rect 489204 488797 489904 489497
rect 490531 488797 491231 489497
rect 491858 488797 492558 489497
rect 493185 488797 493885 489497
rect 494512 488797 495212 489497
rect 495839 488797 496539 489497
rect 497166 488797 497866 489497
rect 498493 488797 499193 489497
rect 499820 488797 500520 489497
rect 501147 488797 501847 489497
rect 502474 488797 503174 489497
rect 503801 488797 504501 489497
rect 505128 488797 505828 489497
rect 506455 488797 507155 489497
rect 87948 487656 88648 488356
rect 88929 487656 89629 488356
rect 89910 487656 90610 488356
rect 90891 487656 91591 488356
rect 91872 487656 92572 488356
rect 92853 487656 93553 488356
rect 93834 487656 94534 488356
rect 94815 487656 95515 488356
rect 95796 487656 96496 488356
rect 96777 487656 97477 488356
rect 97758 487656 98458 488356
rect 98739 487656 99439 488356
rect 99720 487656 100420 488356
rect 100701 487656 101401 488356
rect 101682 487656 102382 488356
rect 102663 487656 103363 488356
rect 103644 487656 104344 488356
rect 104625 487656 105325 488356
rect 105606 487656 106306 488356
rect 106587 487656 107287 488356
rect 107568 487656 108268 488356
rect 108549 487656 109249 488356
rect 109530 487656 110230 488356
rect 110511 487656 111211 488356
rect 111492 487656 112192 488356
rect 482569 487470 483269 488170
rect 483896 487470 484596 488170
rect 485223 487470 485923 488170
rect 486550 487470 487250 488170
rect 487877 487470 488577 488170
rect 489204 487470 489904 488170
rect 490531 487470 491231 488170
rect 491858 487470 492558 488170
rect 493185 487470 493885 488170
rect 494512 487470 495212 488170
rect 495839 487470 496539 488170
rect 497166 487470 497866 488170
rect 498493 487470 499193 488170
rect 499820 487470 500520 488170
rect 501147 487470 501847 488170
rect 502474 487470 503174 488170
rect 503801 487470 504501 488170
rect 505128 487470 505828 488170
rect 506455 487470 507155 488170
rect 87948 486636 88648 487336
rect 88929 486636 89629 487336
rect 89910 486636 90610 487336
rect 90891 486636 91591 487336
rect 91872 486636 92572 487336
rect 92853 486636 93553 487336
rect 93834 486636 94534 487336
rect 94815 486636 95515 487336
rect 95796 486636 96496 487336
rect 96777 486636 97477 487336
rect 97758 486636 98458 487336
rect 98739 486636 99439 487336
rect 99720 486636 100420 487336
rect 100701 486636 101401 487336
rect 101682 486636 102382 487336
rect 102663 486636 103363 487336
rect 103644 486636 104344 487336
rect 104625 486636 105325 487336
rect 105606 486636 106306 487336
rect 106587 486636 107287 487336
rect 107568 486636 108268 487336
rect 108549 486636 109249 487336
rect 109530 486636 110230 487336
rect 110511 486636 111211 487336
rect 111492 486636 112192 487336
rect 87948 485616 88648 486316
rect 88929 485616 89629 486316
rect 89910 485616 90610 486316
rect 90891 485616 91591 486316
rect 91872 485616 92572 486316
rect 92853 485616 93553 486316
rect 93834 485616 94534 486316
rect 94815 485616 95515 486316
rect 95796 485616 96496 486316
rect 96777 485616 97477 486316
rect 97758 485616 98458 486316
rect 98739 485616 99439 486316
rect 99720 485616 100420 486316
rect 100701 485616 101401 486316
rect 101682 485616 102382 486316
rect 102663 485616 103363 486316
rect 103644 485616 104344 486316
rect 104625 485616 105325 486316
rect 105606 485616 106306 486316
rect 106587 485616 107287 486316
rect 107568 485616 108268 486316
rect 108549 485616 109249 486316
rect 109530 485616 110230 486316
rect 110511 485616 111211 486316
rect 111492 485616 112192 486316
rect 482569 486143 483269 486843
rect 483896 486143 484596 486843
rect 485223 486143 485923 486843
rect 486550 486143 487250 486843
rect 487877 486143 488577 486843
rect 489204 486143 489904 486843
rect 490531 486143 491231 486843
rect 491858 486143 492558 486843
rect 493185 486143 493885 486843
rect 494512 486143 495212 486843
rect 495839 486143 496539 486843
rect 497166 486143 497866 486843
rect 498493 486143 499193 486843
rect 499820 486143 500520 486843
rect 501147 486143 501847 486843
rect 502474 486143 503174 486843
rect 503801 486143 504501 486843
rect 505128 486143 505828 486843
rect 506455 486143 507155 486843
rect 482569 484816 483269 485516
rect 483896 484816 484596 485516
rect 485223 484816 485923 485516
rect 486550 484816 487250 485516
rect 487877 484816 488577 485516
rect 489204 484816 489904 485516
rect 490531 484816 491231 485516
rect 491858 484816 492558 485516
rect 493185 484816 493885 485516
rect 494512 484816 495212 485516
rect 495839 484816 496539 485516
rect 497166 484816 497866 485516
rect 498493 484816 499193 485516
rect 499820 484816 500520 485516
rect 501147 484816 501847 485516
rect 502474 484816 503174 485516
rect 503801 484816 504501 485516
rect 505128 484816 505828 485516
rect 506455 484816 507155 485516
rect 482569 483489 483269 484189
rect 483896 483489 484596 484189
rect 485223 483489 485923 484189
rect 486550 483489 487250 484189
rect 487877 483489 488577 484189
rect 489204 483489 489904 484189
rect 490531 483489 491231 484189
rect 491858 483489 492558 484189
rect 493185 483489 493885 484189
rect 494512 483489 495212 484189
rect 495839 483489 496539 484189
rect 497166 483489 497866 484189
rect 498493 483489 499193 484189
rect 499820 483489 500520 484189
rect 501147 483489 501847 484189
rect 502474 483489 503174 484189
rect 503801 483489 504501 484189
rect 505128 483489 505828 484189
rect 506455 483489 507155 484189
rect 119166 479596 119866 480296
rect 120188 479596 120888 480296
rect 121210 479596 121910 480296
rect 122232 479596 122932 480296
rect 123254 479596 123954 480296
rect 124276 479596 124976 480296
rect 125298 479596 125998 480296
rect 126320 479596 127020 480296
rect 127342 479596 128042 480296
rect 128364 479596 129064 480296
rect 129386 479596 130086 480296
rect 130408 479596 131108 480296
rect 131430 479596 132130 480296
rect 132452 479596 133152 480296
rect 133474 479596 134174 480296
rect 134496 479596 135196 480296
rect 135518 479596 136218 480296
rect 136540 479596 137240 480296
rect 137562 479596 138262 480296
rect 138584 479596 139284 480296
rect 139606 479596 140306 480296
rect 140628 479596 141328 480296
rect 141650 479596 142350 480296
rect 142672 479596 143372 480296
rect 143694 479596 144394 480296
rect 444322 480213 445022 480913
rect 445379 480213 446079 480913
rect 446436 480213 447136 480913
rect 447493 480213 448193 480913
rect 448550 480213 449250 480913
rect 449607 480213 450307 480913
rect 450664 480213 451364 480913
rect 451721 480213 452421 480913
rect 452778 480213 453478 480913
rect 453835 480213 454535 480913
rect 454892 480213 455592 480913
rect 455949 480213 456649 480913
rect 457006 480213 457706 480913
rect 458063 480213 458763 480913
rect 459120 480213 459820 480913
rect 460177 480213 460877 480913
rect 461234 480213 461934 480913
rect 462291 480213 462991 480913
rect 463348 480213 464048 480913
rect 464405 480213 465105 480913
rect 465462 480213 466162 480913
rect 466519 480213 467219 480913
rect 467576 480213 468276 480913
rect 119166 478524 119866 479224
rect 120188 478524 120888 479224
rect 121210 478524 121910 479224
rect 122232 478524 122932 479224
rect 123254 478524 123954 479224
rect 124276 478524 124976 479224
rect 125298 478524 125998 479224
rect 126320 478524 127020 479224
rect 127342 478524 128042 479224
rect 128364 478524 129064 479224
rect 129386 478524 130086 479224
rect 130408 478524 131108 479224
rect 131430 478524 132130 479224
rect 132452 478524 133152 479224
rect 133474 478524 134174 479224
rect 134496 478524 135196 479224
rect 135518 478524 136218 479224
rect 136540 478524 137240 479224
rect 137562 478524 138262 479224
rect 138584 478524 139284 479224
rect 139606 478524 140306 479224
rect 140628 478524 141328 479224
rect 141650 478524 142350 479224
rect 142672 478524 143372 479224
rect 143694 478524 144394 479224
rect 444322 479141 445022 479841
rect 445379 479141 446079 479841
rect 446436 479141 447136 479841
rect 447493 479141 448193 479841
rect 448550 479141 449250 479841
rect 449607 479141 450307 479841
rect 450664 479141 451364 479841
rect 451721 479141 452421 479841
rect 452778 479141 453478 479841
rect 453835 479141 454535 479841
rect 454892 479141 455592 479841
rect 455949 479141 456649 479841
rect 457006 479141 457706 479841
rect 458063 479141 458763 479841
rect 459120 479141 459820 479841
rect 460177 479141 460877 479841
rect 461234 479141 461934 479841
rect 462291 479141 462991 479841
rect 463348 479141 464048 479841
rect 464405 479141 465105 479841
rect 465462 479141 466162 479841
rect 466519 479141 467219 479841
rect 467576 479141 468276 479841
rect 119166 477452 119866 478152
rect 120188 477452 120888 478152
rect 121210 477452 121910 478152
rect 122232 477452 122932 478152
rect 123254 477452 123954 478152
rect 124276 477452 124976 478152
rect 125298 477452 125998 478152
rect 126320 477452 127020 478152
rect 127342 477452 128042 478152
rect 128364 477452 129064 478152
rect 129386 477452 130086 478152
rect 130408 477452 131108 478152
rect 131430 477452 132130 478152
rect 132452 477452 133152 478152
rect 133474 477452 134174 478152
rect 134496 477452 135196 478152
rect 135518 477452 136218 478152
rect 136540 477452 137240 478152
rect 137562 477452 138262 478152
rect 138584 477452 139284 478152
rect 139606 477452 140306 478152
rect 140628 477452 141328 478152
rect 141650 477452 142350 478152
rect 142672 477452 143372 478152
rect 143694 477452 144394 478152
rect 444322 478069 445022 478769
rect 445379 478069 446079 478769
rect 446436 478069 447136 478769
rect 447493 478069 448193 478769
rect 448550 478069 449250 478769
rect 449607 478069 450307 478769
rect 450664 478069 451364 478769
rect 451721 478069 452421 478769
rect 452778 478069 453478 478769
rect 453835 478069 454535 478769
rect 454892 478069 455592 478769
rect 455949 478069 456649 478769
rect 457006 478069 457706 478769
rect 458063 478069 458763 478769
rect 459120 478069 459820 478769
rect 460177 478069 460877 478769
rect 461234 478069 461934 478769
rect 462291 478069 462991 478769
rect 463348 478069 464048 478769
rect 464405 478069 465105 478769
rect 465462 478069 466162 478769
rect 466519 478069 467219 478769
rect 467576 478069 468276 478769
rect 119166 476380 119866 477080
rect 120188 476380 120888 477080
rect 121210 476380 121910 477080
rect 122232 476380 122932 477080
rect 123254 476380 123954 477080
rect 124276 476380 124976 477080
rect 125298 476380 125998 477080
rect 126320 476380 127020 477080
rect 127342 476380 128042 477080
rect 128364 476380 129064 477080
rect 129386 476380 130086 477080
rect 130408 476380 131108 477080
rect 131430 476380 132130 477080
rect 132452 476380 133152 477080
rect 133474 476380 134174 477080
rect 134496 476380 135196 477080
rect 135518 476380 136218 477080
rect 136540 476380 137240 477080
rect 137562 476380 138262 477080
rect 138584 476380 139284 477080
rect 139606 476380 140306 477080
rect 140628 476380 141328 477080
rect 141650 476380 142350 477080
rect 142672 476380 143372 477080
rect 143694 476380 144394 477080
rect 444322 476997 445022 477697
rect 445379 476997 446079 477697
rect 446436 476997 447136 477697
rect 447493 476997 448193 477697
rect 448550 476997 449250 477697
rect 449607 476997 450307 477697
rect 450664 476997 451364 477697
rect 451721 476997 452421 477697
rect 452778 476997 453478 477697
rect 453835 476997 454535 477697
rect 454892 476997 455592 477697
rect 455949 476997 456649 477697
rect 457006 476997 457706 477697
rect 458063 476997 458763 477697
rect 459120 476997 459820 477697
rect 460177 476997 460877 477697
rect 461234 476997 461934 477697
rect 462291 476997 462991 477697
rect 463348 476997 464048 477697
rect 464405 476997 465105 477697
rect 465462 476997 466162 477697
rect 466519 476997 467219 477697
rect 467576 476997 468276 477697
rect 119166 475308 119866 476008
rect 120188 475308 120888 476008
rect 121210 475308 121910 476008
rect 122232 475308 122932 476008
rect 123254 475308 123954 476008
rect 124276 475308 124976 476008
rect 125298 475308 125998 476008
rect 126320 475308 127020 476008
rect 127342 475308 128042 476008
rect 128364 475308 129064 476008
rect 129386 475308 130086 476008
rect 130408 475308 131108 476008
rect 131430 475308 132130 476008
rect 132452 475308 133152 476008
rect 133474 475308 134174 476008
rect 134496 475308 135196 476008
rect 135518 475308 136218 476008
rect 136540 475308 137240 476008
rect 137562 475308 138262 476008
rect 138584 475308 139284 476008
rect 139606 475308 140306 476008
rect 140628 475308 141328 476008
rect 141650 475308 142350 476008
rect 142672 475308 143372 476008
rect 143694 475308 144394 476008
rect 444322 475925 445022 476625
rect 445379 475925 446079 476625
rect 446436 475925 447136 476625
rect 447493 475925 448193 476625
rect 448550 475925 449250 476625
rect 449607 475925 450307 476625
rect 450664 475925 451364 476625
rect 451721 475925 452421 476625
rect 452778 475925 453478 476625
rect 453835 475925 454535 476625
rect 454892 475925 455592 476625
rect 455949 475925 456649 476625
rect 457006 475925 457706 476625
rect 458063 475925 458763 476625
rect 459120 475925 459820 476625
rect 460177 475925 460877 476625
rect 461234 475925 461934 476625
rect 462291 475925 462991 476625
rect 463348 475925 464048 476625
rect 464405 475925 465105 476625
rect 465462 475925 466162 476625
rect 466519 475925 467219 476625
rect 467576 475925 468276 476625
rect 119166 474236 119866 474936
rect 120188 474236 120888 474936
rect 121210 474236 121910 474936
rect 122232 474236 122932 474936
rect 123254 474236 123954 474936
rect 124276 474236 124976 474936
rect 125298 474236 125998 474936
rect 126320 474236 127020 474936
rect 127342 474236 128042 474936
rect 128364 474236 129064 474936
rect 129386 474236 130086 474936
rect 130408 474236 131108 474936
rect 131430 474236 132130 474936
rect 132452 474236 133152 474936
rect 133474 474236 134174 474936
rect 134496 474236 135196 474936
rect 135518 474236 136218 474936
rect 136540 474236 137240 474936
rect 137562 474236 138262 474936
rect 138584 474236 139284 474936
rect 139606 474236 140306 474936
rect 140628 474236 141328 474936
rect 141650 474236 142350 474936
rect 142672 474236 143372 474936
rect 143694 474236 144394 474936
rect 444322 474853 445022 475553
rect 445379 474853 446079 475553
rect 446436 474853 447136 475553
rect 447493 474853 448193 475553
rect 448550 474853 449250 475553
rect 449607 474853 450307 475553
rect 450664 474853 451364 475553
rect 451721 474853 452421 475553
rect 452778 474853 453478 475553
rect 453835 474853 454535 475553
rect 454892 474853 455592 475553
rect 455949 474853 456649 475553
rect 457006 474853 457706 475553
rect 458063 474853 458763 475553
rect 459120 474853 459820 475553
rect 460177 474853 460877 475553
rect 461234 474853 461934 475553
rect 462291 474853 462991 475553
rect 463348 474853 464048 475553
rect 464405 474853 465105 475553
rect 465462 474853 466162 475553
rect 466519 474853 467219 475553
rect 467576 474853 468276 475553
rect 119166 473164 119866 473864
rect 120188 473164 120888 473864
rect 121210 473164 121910 473864
rect 122232 473164 122932 473864
rect 123254 473164 123954 473864
rect 124276 473164 124976 473864
rect 125298 473164 125998 473864
rect 126320 473164 127020 473864
rect 127342 473164 128042 473864
rect 128364 473164 129064 473864
rect 129386 473164 130086 473864
rect 130408 473164 131108 473864
rect 131430 473164 132130 473864
rect 132452 473164 133152 473864
rect 133474 473164 134174 473864
rect 134496 473164 135196 473864
rect 135518 473164 136218 473864
rect 136540 473164 137240 473864
rect 137562 473164 138262 473864
rect 138584 473164 139284 473864
rect 139606 473164 140306 473864
rect 140628 473164 141328 473864
rect 141650 473164 142350 473864
rect 142672 473164 143372 473864
rect 143694 473164 144394 473864
rect 444322 473781 445022 474481
rect 445379 473781 446079 474481
rect 446436 473781 447136 474481
rect 447493 473781 448193 474481
rect 448550 473781 449250 474481
rect 449607 473781 450307 474481
rect 450664 473781 451364 474481
rect 451721 473781 452421 474481
rect 452778 473781 453478 474481
rect 453835 473781 454535 474481
rect 454892 473781 455592 474481
rect 455949 473781 456649 474481
rect 457006 473781 457706 474481
rect 458063 473781 458763 474481
rect 459120 473781 459820 474481
rect 460177 473781 460877 474481
rect 461234 473781 461934 474481
rect 462291 473781 462991 474481
rect 463348 473781 464048 474481
rect 464405 473781 465105 474481
rect 465462 473781 466162 474481
rect 466519 473781 467219 474481
rect 467576 473781 468276 474481
rect 119166 472092 119866 472792
rect 120188 472092 120888 472792
rect 121210 472092 121910 472792
rect 122232 472092 122932 472792
rect 123254 472092 123954 472792
rect 124276 472092 124976 472792
rect 125298 472092 125998 472792
rect 126320 472092 127020 472792
rect 127342 472092 128042 472792
rect 128364 472092 129064 472792
rect 129386 472092 130086 472792
rect 130408 472092 131108 472792
rect 131430 472092 132130 472792
rect 132452 472092 133152 472792
rect 133474 472092 134174 472792
rect 134496 472092 135196 472792
rect 135518 472092 136218 472792
rect 136540 472092 137240 472792
rect 137562 472092 138262 472792
rect 138584 472092 139284 472792
rect 139606 472092 140306 472792
rect 140628 472092 141328 472792
rect 141650 472092 142350 472792
rect 142672 472092 143372 472792
rect 143694 472092 144394 472792
rect 444322 472709 445022 473409
rect 445379 472709 446079 473409
rect 446436 472709 447136 473409
rect 447493 472709 448193 473409
rect 448550 472709 449250 473409
rect 449607 472709 450307 473409
rect 450664 472709 451364 473409
rect 451721 472709 452421 473409
rect 452778 472709 453478 473409
rect 453835 472709 454535 473409
rect 454892 472709 455592 473409
rect 455949 472709 456649 473409
rect 457006 472709 457706 473409
rect 458063 472709 458763 473409
rect 459120 472709 459820 473409
rect 460177 472709 460877 473409
rect 461234 472709 461934 473409
rect 462291 472709 462991 473409
rect 463348 472709 464048 473409
rect 464405 472709 465105 473409
rect 465462 472709 466162 473409
rect 466519 472709 467219 473409
rect 467576 472709 468276 473409
rect 119166 471020 119866 471720
rect 120188 471020 120888 471720
rect 121210 471020 121910 471720
rect 122232 471020 122932 471720
rect 123254 471020 123954 471720
rect 124276 471020 124976 471720
rect 125298 471020 125998 471720
rect 126320 471020 127020 471720
rect 127342 471020 128042 471720
rect 128364 471020 129064 471720
rect 129386 471020 130086 471720
rect 130408 471020 131108 471720
rect 131430 471020 132130 471720
rect 132452 471020 133152 471720
rect 133474 471020 134174 471720
rect 134496 471020 135196 471720
rect 135518 471020 136218 471720
rect 136540 471020 137240 471720
rect 137562 471020 138262 471720
rect 138584 471020 139284 471720
rect 139606 471020 140306 471720
rect 140628 471020 141328 471720
rect 141650 471020 142350 471720
rect 142672 471020 143372 471720
rect 143694 471020 144394 471720
rect 444322 471637 445022 472337
rect 445379 471637 446079 472337
rect 446436 471637 447136 472337
rect 447493 471637 448193 472337
rect 448550 471637 449250 472337
rect 449607 471637 450307 472337
rect 450664 471637 451364 472337
rect 451721 471637 452421 472337
rect 452778 471637 453478 472337
rect 453835 471637 454535 472337
rect 454892 471637 455592 472337
rect 455949 471637 456649 472337
rect 457006 471637 457706 472337
rect 458063 471637 458763 472337
rect 459120 471637 459820 472337
rect 460177 471637 460877 472337
rect 461234 471637 461934 472337
rect 462291 471637 462991 472337
rect 463348 471637 464048 472337
rect 464405 471637 465105 472337
rect 465462 471637 466162 472337
rect 466519 471637 467219 472337
rect 467576 471637 468276 472337
rect 119166 469948 119866 470648
rect 120188 469948 120888 470648
rect 121210 469948 121910 470648
rect 122232 469948 122932 470648
rect 123254 469948 123954 470648
rect 124276 469948 124976 470648
rect 125298 469948 125998 470648
rect 126320 469948 127020 470648
rect 127342 469948 128042 470648
rect 128364 469948 129064 470648
rect 129386 469948 130086 470648
rect 130408 469948 131108 470648
rect 131430 469948 132130 470648
rect 132452 469948 133152 470648
rect 133474 469948 134174 470648
rect 134496 469948 135196 470648
rect 135518 469948 136218 470648
rect 136540 469948 137240 470648
rect 137562 469948 138262 470648
rect 138584 469948 139284 470648
rect 139606 469948 140306 470648
rect 140628 469948 141328 470648
rect 141650 469948 142350 470648
rect 142672 469948 143372 470648
rect 143694 469948 144394 470648
rect 444322 470565 445022 471265
rect 445379 470565 446079 471265
rect 446436 470565 447136 471265
rect 447493 470565 448193 471265
rect 448550 470565 449250 471265
rect 449607 470565 450307 471265
rect 450664 470565 451364 471265
rect 451721 470565 452421 471265
rect 452778 470565 453478 471265
rect 453835 470565 454535 471265
rect 454892 470565 455592 471265
rect 455949 470565 456649 471265
rect 457006 470565 457706 471265
rect 458063 470565 458763 471265
rect 459120 470565 459820 471265
rect 460177 470565 460877 471265
rect 461234 470565 461934 471265
rect 462291 470565 462991 471265
rect 463348 470565 464048 471265
rect 464405 470565 465105 471265
rect 465462 470565 466162 471265
rect 466519 470565 467219 471265
rect 467576 470565 468276 471265
rect 119166 468876 119866 469576
rect 120188 468876 120888 469576
rect 121210 468876 121910 469576
rect 122232 468876 122932 469576
rect 123254 468876 123954 469576
rect 124276 468876 124976 469576
rect 125298 468876 125998 469576
rect 126320 468876 127020 469576
rect 127342 468876 128042 469576
rect 128364 468876 129064 469576
rect 129386 468876 130086 469576
rect 130408 468876 131108 469576
rect 131430 468876 132130 469576
rect 132452 468876 133152 469576
rect 133474 468876 134174 469576
rect 134496 468876 135196 469576
rect 135518 468876 136218 469576
rect 136540 468876 137240 469576
rect 137562 468876 138262 469576
rect 138584 468876 139284 469576
rect 139606 468876 140306 469576
rect 140628 468876 141328 469576
rect 141650 468876 142350 469576
rect 142672 468876 143372 469576
rect 143694 468876 144394 469576
rect 444322 469493 445022 470193
rect 445379 469493 446079 470193
rect 446436 469493 447136 470193
rect 447493 469493 448193 470193
rect 448550 469493 449250 470193
rect 449607 469493 450307 470193
rect 450664 469493 451364 470193
rect 451721 469493 452421 470193
rect 452778 469493 453478 470193
rect 453835 469493 454535 470193
rect 454892 469493 455592 470193
rect 455949 469493 456649 470193
rect 457006 469493 457706 470193
rect 458063 469493 458763 470193
rect 459120 469493 459820 470193
rect 460177 469493 460877 470193
rect 461234 469493 461934 470193
rect 462291 469493 462991 470193
rect 463348 469493 464048 470193
rect 464405 469493 465105 470193
rect 465462 469493 466162 470193
rect 466519 469493 467219 470193
rect 467576 469493 468276 470193
rect 91879 467431 92029 467581
rect 92147 467431 92297 467581
rect 92415 467431 92565 467581
rect 92683 467431 92833 467581
rect 92951 467431 93101 467581
rect 93219 467431 93369 467581
rect 93487 467431 93637 467581
rect 93755 467431 93905 467581
rect 94023 467431 94173 467581
rect 94291 467431 94441 467581
rect 91879 467193 92029 467343
rect 92147 467193 92297 467343
rect 92415 467193 92565 467343
rect 92683 467193 92833 467343
rect 92951 467193 93101 467343
rect 93219 467193 93369 467343
rect 93487 467193 93637 467343
rect 93755 467193 93905 467343
rect 94023 467193 94173 467343
rect 94291 467193 94441 467343
rect 91879 466955 92029 467105
rect 92147 466955 92297 467105
rect 92415 466955 92565 467105
rect 92683 466955 92833 467105
rect 92951 466955 93101 467105
rect 93219 466955 93369 467105
rect 93487 466955 93637 467105
rect 93755 466955 93905 467105
rect 94023 466955 94173 467105
rect 94291 466955 94441 467105
rect 91879 466717 92029 466867
rect 92147 466717 92297 466867
rect 92415 466717 92565 466867
rect 92683 466717 92833 466867
rect 92951 466717 93101 466867
rect 93219 466717 93369 466867
rect 93487 466717 93637 466867
rect 93755 466717 93905 466867
rect 94023 466717 94173 466867
rect 94291 466717 94441 466867
rect 91879 466479 92029 466629
rect 92147 466479 92297 466629
rect 92415 466479 92565 466629
rect 92683 466479 92833 466629
rect 92951 466479 93101 466629
rect 93219 466479 93369 466629
rect 93487 466479 93637 466629
rect 93755 466479 93905 466629
rect 94023 466479 94173 466629
rect 94291 466479 94441 466629
rect 91879 466241 92029 466391
rect 92147 466241 92297 466391
rect 92415 466241 92565 466391
rect 92683 466241 92833 466391
rect 92951 466241 93101 466391
rect 93219 466241 93369 466391
rect 93487 466241 93637 466391
rect 93755 466241 93905 466391
rect 94023 466241 94173 466391
rect 94291 466241 94441 466391
rect 91879 466003 92029 466153
rect 92147 466003 92297 466153
rect 92415 466003 92565 466153
rect 92683 466003 92833 466153
rect 92951 466003 93101 466153
rect 93219 466003 93369 466153
rect 93487 466003 93637 466153
rect 93755 466003 93905 466153
rect 94023 466003 94173 466153
rect 94291 466003 94441 466153
rect 91879 465765 92029 465915
rect 92147 465765 92297 465915
rect 92415 465765 92565 465915
rect 92683 465765 92833 465915
rect 92951 465765 93101 465915
rect 93219 465765 93369 465915
rect 93487 465765 93637 465915
rect 93755 465765 93905 465915
rect 94023 465765 94173 465915
rect 94291 465765 94441 465915
rect 91879 465527 92029 465677
rect 92147 465527 92297 465677
rect 92415 465527 92565 465677
rect 92683 465527 92833 465677
rect 92951 465527 93101 465677
rect 93219 465527 93369 465677
rect 93487 465527 93637 465677
rect 93755 465527 93905 465677
rect 94023 465527 94173 465677
rect 94291 465527 94441 465677
rect 91879 465289 92029 465439
rect 92147 465289 92297 465439
rect 92415 465289 92565 465439
rect 92683 465289 92833 465439
rect 92951 465289 93101 465439
rect 93219 465289 93369 465439
rect 93487 465289 93637 465439
rect 93755 465289 93905 465439
rect 94023 465289 94173 465439
rect 94291 465289 94441 465439
rect 119166 467804 119866 468504
rect 120188 467804 120888 468504
rect 121210 467804 121910 468504
rect 122232 467804 122932 468504
rect 123254 467804 123954 468504
rect 124276 467804 124976 468504
rect 125298 467804 125998 468504
rect 126320 467804 127020 468504
rect 127342 467804 128042 468504
rect 128364 467804 129064 468504
rect 129386 467804 130086 468504
rect 130408 467804 131108 468504
rect 131430 467804 132130 468504
rect 132452 467804 133152 468504
rect 133474 467804 134174 468504
rect 134496 467804 135196 468504
rect 135518 467804 136218 468504
rect 136540 467804 137240 468504
rect 137562 467804 138262 468504
rect 138584 467804 139284 468504
rect 139606 467804 140306 468504
rect 140628 467804 141328 468504
rect 141650 467804 142350 468504
rect 142672 467804 143372 468504
rect 143694 467804 144394 468504
rect 444322 468421 445022 469121
rect 445379 468421 446079 469121
rect 446436 468421 447136 469121
rect 447493 468421 448193 469121
rect 448550 468421 449250 469121
rect 449607 468421 450307 469121
rect 450664 468421 451364 469121
rect 451721 468421 452421 469121
rect 452778 468421 453478 469121
rect 453835 468421 454535 469121
rect 454892 468421 455592 469121
rect 455949 468421 456649 469121
rect 457006 468421 457706 469121
rect 458063 468421 458763 469121
rect 459120 468421 459820 469121
rect 460177 468421 460877 469121
rect 461234 468421 461934 469121
rect 462291 468421 462991 469121
rect 463348 468421 464048 469121
rect 464405 468421 465105 469121
rect 465462 468421 466162 469121
rect 466519 468421 467219 469121
rect 467576 468421 468276 469121
rect 119166 466732 119866 467432
rect 120188 466732 120888 467432
rect 121210 466732 121910 467432
rect 122232 466732 122932 467432
rect 123254 466732 123954 467432
rect 124276 466732 124976 467432
rect 125298 466732 125998 467432
rect 126320 466732 127020 467432
rect 127342 466732 128042 467432
rect 128364 466732 129064 467432
rect 129386 466732 130086 467432
rect 130408 466732 131108 467432
rect 131430 466732 132130 467432
rect 132452 466732 133152 467432
rect 133474 466732 134174 467432
rect 134496 466732 135196 467432
rect 135518 466732 136218 467432
rect 136540 466732 137240 467432
rect 137562 466732 138262 467432
rect 138584 466732 139284 467432
rect 139606 466732 140306 467432
rect 140628 466732 141328 467432
rect 141650 466732 142350 467432
rect 142672 466732 143372 467432
rect 143694 466732 144394 467432
rect 444322 467349 445022 468049
rect 445379 467349 446079 468049
rect 446436 467349 447136 468049
rect 447493 467349 448193 468049
rect 448550 467349 449250 468049
rect 449607 467349 450307 468049
rect 450664 467349 451364 468049
rect 451721 467349 452421 468049
rect 452778 467349 453478 468049
rect 453835 467349 454535 468049
rect 454892 467349 455592 468049
rect 455949 467349 456649 468049
rect 457006 467349 457706 468049
rect 458063 467349 458763 468049
rect 459120 467349 459820 468049
rect 460177 467349 460877 468049
rect 461234 467349 461934 468049
rect 462291 467349 462991 468049
rect 463348 467349 464048 468049
rect 464405 467349 465105 468049
rect 465462 467349 466162 468049
rect 466519 467349 467219 468049
rect 467576 467349 468276 468049
rect 119166 465660 119866 466360
rect 120188 465660 120888 466360
rect 121210 465660 121910 466360
rect 122232 465660 122932 466360
rect 123254 465660 123954 466360
rect 124276 465660 124976 466360
rect 125298 465660 125998 466360
rect 126320 465660 127020 466360
rect 127342 465660 128042 466360
rect 128364 465660 129064 466360
rect 129386 465660 130086 466360
rect 130408 465660 131108 466360
rect 131430 465660 132130 466360
rect 132452 465660 133152 466360
rect 133474 465660 134174 466360
rect 134496 465660 135196 466360
rect 135518 465660 136218 466360
rect 136540 465660 137240 466360
rect 137562 465660 138262 466360
rect 138584 465660 139284 466360
rect 139606 465660 140306 466360
rect 140628 465660 141328 466360
rect 141650 465660 142350 466360
rect 142672 465660 143372 466360
rect 143694 465660 144394 466360
rect 444322 466277 445022 466977
rect 445379 466277 446079 466977
rect 446436 466277 447136 466977
rect 447493 466277 448193 466977
rect 448550 466277 449250 466977
rect 449607 466277 450307 466977
rect 450664 466277 451364 466977
rect 451721 466277 452421 466977
rect 452778 466277 453478 466977
rect 453835 466277 454535 466977
rect 454892 466277 455592 466977
rect 455949 466277 456649 466977
rect 457006 466277 457706 466977
rect 458063 466277 458763 466977
rect 459120 466277 459820 466977
rect 460177 466277 460877 466977
rect 461234 466277 461934 466977
rect 462291 466277 462991 466977
rect 463348 466277 464048 466977
rect 464405 466277 465105 466977
rect 465462 466277 466162 466977
rect 466519 466277 467219 466977
rect 467576 466277 468276 466977
rect 119166 464588 119866 465288
rect 120188 464588 120888 465288
rect 121210 464588 121910 465288
rect 122232 464588 122932 465288
rect 123254 464588 123954 465288
rect 124276 464588 124976 465288
rect 125298 464588 125998 465288
rect 126320 464588 127020 465288
rect 127342 464588 128042 465288
rect 128364 464588 129064 465288
rect 129386 464588 130086 465288
rect 130408 464588 131108 465288
rect 131430 464588 132130 465288
rect 132452 464588 133152 465288
rect 133474 464588 134174 465288
rect 134496 464588 135196 465288
rect 135518 464588 136218 465288
rect 136540 464588 137240 465288
rect 137562 464588 138262 465288
rect 138584 464588 139284 465288
rect 139606 464588 140306 465288
rect 140628 464588 141328 465288
rect 141650 464588 142350 465288
rect 142672 464588 143372 465288
rect 143694 464588 144394 465288
rect 444322 465205 445022 465905
rect 445379 465205 446079 465905
rect 446436 465205 447136 465905
rect 447493 465205 448193 465905
rect 448550 465205 449250 465905
rect 449607 465205 450307 465905
rect 450664 465205 451364 465905
rect 451721 465205 452421 465905
rect 452778 465205 453478 465905
rect 453835 465205 454535 465905
rect 454892 465205 455592 465905
rect 455949 465205 456649 465905
rect 457006 465205 457706 465905
rect 458063 465205 458763 465905
rect 459120 465205 459820 465905
rect 460177 465205 460877 465905
rect 461234 465205 461934 465905
rect 462291 465205 462991 465905
rect 463348 465205 464048 465905
rect 464405 465205 465105 465905
rect 465462 465205 466162 465905
rect 466519 465205 467219 465905
rect 467576 465205 468276 465905
rect 119166 463516 119866 464216
rect 120188 463516 120888 464216
rect 121210 463516 121910 464216
rect 122232 463516 122932 464216
rect 123254 463516 123954 464216
rect 124276 463516 124976 464216
rect 125298 463516 125998 464216
rect 126320 463516 127020 464216
rect 127342 463516 128042 464216
rect 128364 463516 129064 464216
rect 129386 463516 130086 464216
rect 130408 463516 131108 464216
rect 131430 463516 132130 464216
rect 132452 463516 133152 464216
rect 133474 463516 134174 464216
rect 134496 463516 135196 464216
rect 135518 463516 136218 464216
rect 136540 463516 137240 464216
rect 137562 463516 138262 464216
rect 138584 463516 139284 464216
rect 139606 463516 140306 464216
rect 140628 463516 141328 464216
rect 141650 463516 142350 464216
rect 142672 463516 143372 464216
rect 143694 463516 144394 464216
rect 444322 464133 445022 464833
rect 445379 464133 446079 464833
rect 446436 464133 447136 464833
rect 447493 464133 448193 464833
rect 448550 464133 449250 464833
rect 449607 464133 450307 464833
rect 450664 464133 451364 464833
rect 451721 464133 452421 464833
rect 452778 464133 453478 464833
rect 453835 464133 454535 464833
rect 454892 464133 455592 464833
rect 455949 464133 456649 464833
rect 457006 464133 457706 464833
rect 458063 464133 458763 464833
rect 459120 464133 459820 464833
rect 460177 464133 460877 464833
rect 461234 464133 461934 464833
rect 462291 464133 462991 464833
rect 463348 464133 464048 464833
rect 464405 464133 465105 464833
rect 465462 464133 466162 464833
rect 466519 464133 467219 464833
rect 467576 464133 468276 464833
rect 119166 462444 119866 463144
rect 120188 462444 120888 463144
rect 121210 462444 121910 463144
rect 122232 462444 122932 463144
rect 123254 462444 123954 463144
rect 124276 462444 124976 463144
rect 125298 462444 125998 463144
rect 126320 462444 127020 463144
rect 127342 462444 128042 463144
rect 128364 462444 129064 463144
rect 129386 462444 130086 463144
rect 130408 462444 131108 463144
rect 131430 462444 132130 463144
rect 132452 462444 133152 463144
rect 133474 462444 134174 463144
rect 134496 462444 135196 463144
rect 135518 462444 136218 463144
rect 136540 462444 137240 463144
rect 137562 462444 138262 463144
rect 138584 462444 139284 463144
rect 139606 462444 140306 463144
rect 140628 462444 141328 463144
rect 141650 462444 142350 463144
rect 142672 462444 143372 463144
rect 143694 462444 144394 463144
rect 119166 461372 119866 462072
rect 120188 461372 120888 462072
rect 121210 461372 121910 462072
rect 122232 461372 122932 462072
rect 123254 461372 123954 462072
rect 124276 461372 124976 462072
rect 125298 461372 125998 462072
rect 126320 461372 127020 462072
rect 127342 461372 128042 462072
rect 128364 461372 129064 462072
rect 129386 461372 130086 462072
rect 130408 461372 131108 462072
rect 131430 461372 132130 462072
rect 132452 461372 133152 462072
rect 133474 461372 134174 462072
rect 134496 461372 135196 462072
rect 135518 461372 136218 462072
rect 136540 461372 137240 462072
rect 137562 461372 138262 462072
rect 138584 461372 139284 462072
rect 139606 461372 140306 462072
rect 140628 461372 141328 462072
rect 141650 461372 142350 462072
rect 142672 461372 143372 462072
rect 143694 461372 144394 462072
rect 119166 460300 119866 461000
rect 120188 460300 120888 461000
rect 121210 460300 121910 461000
rect 122232 460300 122932 461000
rect 123254 460300 123954 461000
rect 124276 460300 124976 461000
rect 125298 460300 125998 461000
rect 126320 460300 127020 461000
rect 127342 460300 128042 461000
rect 128364 460300 129064 461000
rect 129386 460300 130086 461000
rect 130408 460300 131108 461000
rect 131430 460300 132130 461000
rect 132452 460300 133152 461000
rect 133474 460300 134174 461000
rect 134496 460300 135196 461000
rect 135518 460300 136218 461000
rect 136540 460300 137240 461000
rect 137562 460300 138262 461000
rect 138584 460300 139284 461000
rect 139606 460300 140306 461000
rect 140628 460300 141328 461000
rect 141650 460300 142350 461000
rect 142672 460300 143372 461000
rect 143694 460300 144394 461000
rect 119166 459228 119866 459928
rect 120188 459228 120888 459928
rect 121210 459228 121910 459928
rect 122232 459228 122932 459928
rect 123254 459228 123954 459928
rect 124276 459228 124976 459928
rect 125298 459228 125998 459928
rect 126320 459228 127020 459928
rect 127342 459228 128042 459928
rect 128364 459228 129064 459928
rect 129386 459228 130086 459928
rect 130408 459228 131108 459928
rect 131430 459228 132130 459928
rect 132452 459228 133152 459928
rect 133474 459228 134174 459928
rect 134496 459228 135196 459928
rect 135518 459228 136218 459928
rect 136540 459228 137240 459928
rect 137562 459228 138262 459928
rect 138584 459228 139284 459928
rect 139606 459228 140306 459928
rect 140628 459228 141328 459928
rect 141650 459228 142350 459928
rect 142672 459228 143372 459928
rect 143694 459228 144394 459928
rect 444322 463061 445022 463761
rect 445379 463061 446079 463761
rect 446436 463061 447136 463761
rect 447493 463061 448193 463761
rect 448550 463061 449250 463761
rect 449607 463061 450307 463761
rect 450664 463061 451364 463761
rect 451721 463061 452421 463761
rect 452778 463061 453478 463761
rect 453835 463061 454535 463761
rect 454892 463061 455592 463761
rect 455949 463061 456649 463761
rect 457006 463061 457706 463761
rect 458063 463061 458763 463761
rect 459120 463061 459820 463761
rect 460177 463061 460877 463761
rect 461234 463061 461934 463761
rect 462291 463061 462991 463761
rect 463348 463061 464048 463761
rect 464405 463061 465105 463761
rect 465462 463061 466162 463761
rect 466519 463061 467219 463761
rect 467576 463061 468276 463761
rect 444322 461989 445022 462689
rect 445379 461989 446079 462689
rect 446436 461989 447136 462689
rect 447493 461989 448193 462689
rect 448550 461989 449250 462689
rect 449607 461989 450307 462689
rect 450664 461989 451364 462689
rect 451721 461989 452421 462689
rect 452778 461989 453478 462689
rect 453835 461989 454535 462689
rect 454892 461989 455592 462689
rect 455949 461989 456649 462689
rect 457006 461989 457706 462689
rect 458063 461989 458763 462689
rect 459120 461989 459820 462689
rect 460177 461989 460877 462689
rect 461234 461989 461934 462689
rect 462291 461989 462991 462689
rect 463348 461989 464048 462689
rect 464405 461989 465105 462689
rect 465462 461989 466162 462689
rect 466519 461989 467219 462689
rect 467576 461989 468276 462689
rect 444322 460917 445022 461617
rect 445379 460917 446079 461617
rect 446436 460917 447136 461617
rect 447493 460917 448193 461617
rect 448550 460917 449250 461617
rect 449607 460917 450307 461617
rect 450664 460917 451364 461617
rect 451721 460917 452421 461617
rect 452778 460917 453478 461617
rect 453835 460917 454535 461617
rect 454892 460917 455592 461617
rect 455949 460917 456649 461617
rect 457006 460917 457706 461617
rect 458063 460917 458763 461617
rect 459120 460917 459820 461617
rect 460177 460917 460877 461617
rect 461234 460917 461934 461617
rect 462291 460917 462991 461617
rect 463348 460917 464048 461617
rect 464405 460917 465105 461617
rect 465462 460917 466162 461617
rect 466519 460917 467219 461617
rect 467576 460917 468276 461617
rect 444322 459845 445022 460545
rect 445379 459845 446079 460545
rect 446436 459845 447136 460545
rect 447493 459845 448193 460545
rect 448550 459845 449250 460545
rect 449607 459845 450307 460545
rect 450664 459845 451364 460545
rect 451721 459845 452421 460545
rect 452778 459845 453478 460545
rect 453835 459845 454535 460545
rect 454892 459845 455592 460545
rect 455949 459845 456649 460545
rect 457006 459845 457706 460545
rect 458063 459845 458763 460545
rect 459120 459845 459820 460545
rect 460177 459845 460877 460545
rect 461234 459845 461934 460545
rect 462291 459845 462991 460545
rect 463348 459845 464048 460545
rect 464405 459845 465105 460545
rect 465462 459845 466162 460545
rect 466519 459845 467219 460545
rect 467576 459845 468276 460545
rect 444322 458773 445022 459473
rect 445379 458773 446079 459473
rect 446436 458773 447136 459473
rect 447493 458773 448193 459473
rect 448550 458773 449250 459473
rect 449607 458773 450307 459473
rect 450664 458773 451364 459473
rect 451721 458773 452421 459473
rect 452778 458773 453478 459473
rect 453835 458773 454535 459473
rect 454892 458773 455592 459473
rect 455949 458773 456649 459473
rect 457006 458773 457706 459473
rect 458063 458773 458763 459473
rect 459120 458773 459820 459473
rect 460177 458773 460877 459473
rect 461234 458773 461934 459473
rect 462291 458773 462991 459473
rect 463348 458773 464048 459473
rect 464405 458773 465105 459473
rect 465462 458773 466162 459473
rect 466519 458773 467219 459473
rect 467576 458773 468276 459473
rect 444322 457701 445022 458401
rect 445379 457701 446079 458401
rect 446436 457701 447136 458401
rect 447493 457701 448193 458401
rect 448550 457701 449250 458401
rect 449607 457701 450307 458401
rect 450664 457701 451364 458401
rect 451721 457701 452421 458401
rect 452778 457701 453478 458401
rect 453835 457701 454535 458401
rect 454892 457701 455592 458401
rect 455949 457701 456649 458401
rect 457006 457701 457706 458401
rect 458063 457701 458763 458401
rect 459120 457701 459820 458401
rect 460177 457701 460877 458401
rect 461234 457701 461934 458401
rect 462291 457701 462991 458401
rect 463348 457701 464048 458401
rect 464405 457701 465105 458401
rect 465462 457701 466162 458401
rect 466519 457701 467219 458401
rect 467576 457701 468276 458401
rect 122043 367315 122193 367465
rect 122311 367315 122461 367465
rect 122579 367315 122729 367465
rect 122847 367315 122997 367465
rect 123115 367315 123265 367465
rect 123383 367315 123533 367465
rect 123651 367315 123801 367465
rect 123919 367315 124069 367465
rect 124187 367315 124337 367465
rect 124455 367315 124605 367465
rect 122043 367077 122193 367227
rect 122311 367077 122461 367227
rect 122579 367077 122729 367227
rect 122847 367077 122997 367227
rect 123115 367077 123265 367227
rect 123383 367077 123533 367227
rect 123651 367077 123801 367227
rect 123919 367077 124069 367227
rect 124187 367077 124337 367227
rect 124455 367077 124605 367227
rect 122043 366839 122193 366989
rect 122311 366839 122461 366989
rect 122579 366839 122729 366989
rect 122847 366839 122997 366989
rect 123115 366839 123265 366989
rect 123383 366839 123533 366989
rect 123651 366839 123801 366989
rect 123919 366839 124069 366989
rect 124187 366839 124337 366989
rect 124455 366839 124605 366989
rect 122043 366601 122193 366751
rect 122311 366601 122461 366751
rect 122579 366601 122729 366751
rect 122847 366601 122997 366751
rect 123115 366601 123265 366751
rect 123383 366601 123533 366751
rect 123651 366601 123801 366751
rect 123919 366601 124069 366751
rect 124187 366601 124337 366751
rect 124455 366601 124605 366751
rect 122043 366363 122193 366513
rect 122311 366363 122461 366513
rect 122579 366363 122729 366513
rect 122847 366363 122997 366513
rect 123115 366363 123265 366513
rect 123383 366363 123533 366513
rect 123651 366363 123801 366513
rect 123919 366363 124069 366513
rect 124187 366363 124337 366513
rect 124455 366363 124605 366513
rect 122043 366125 122193 366275
rect 122311 366125 122461 366275
rect 122579 366125 122729 366275
rect 122847 366125 122997 366275
rect 123115 366125 123265 366275
rect 123383 366125 123533 366275
rect 123651 366125 123801 366275
rect 123919 366125 124069 366275
rect 124187 366125 124337 366275
rect 124455 366125 124605 366275
rect 122043 365887 122193 366037
rect 122311 365887 122461 366037
rect 122579 365887 122729 366037
rect 122847 365887 122997 366037
rect 123115 365887 123265 366037
rect 123383 365887 123533 366037
rect 123651 365887 123801 366037
rect 123919 365887 124069 366037
rect 124187 365887 124337 366037
rect 124455 365887 124605 366037
rect 122043 365649 122193 365799
rect 122311 365649 122461 365799
rect 122579 365649 122729 365799
rect 122847 365649 122997 365799
rect 123115 365649 123265 365799
rect 123383 365649 123533 365799
rect 123651 365649 123801 365799
rect 123919 365649 124069 365799
rect 124187 365649 124337 365799
rect 124455 365649 124605 365799
rect 122043 365411 122193 365561
rect 122311 365411 122461 365561
rect 122579 365411 122729 365561
rect 122847 365411 122997 365561
rect 123115 365411 123265 365561
rect 123383 365411 123533 365561
rect 123651 365411 123801 365561
rect 123919 365411 124069 365561
rect 124187 365411 124337 365561
rect 124455 365411 124605 365561
rect 122043 365173 122193 365323
rect 122311 365173 122461 365323
rect 122579 365173 122729 365323
rect 122847 365173 122997 365323
rect 123115 365173 123265 365323
rect 123383 365173 123533 365323
rect 123651 365173 123801 365323
rect 123919 365173 124069 365323
rect 124187 365173 124337 365323
rect 124455 365173 124605 365323
rect 443943 148965 444643 149665
rect 445021 148965 445721 149665
rect 446099 148965 446799 149665
rect 447177 148965 447877 149665
rect 448255 148965 448955 149665
rect 449333 148965 450033 149665
rect 450411 148965 451111 149665
rect 451489 148965 452189 149665
rect 452567 148965 453267 149665
rect 453645 148965 454345 149665
rect 454723 148965 455423 149665
rect 455801 148965 456501 149665
rect 456879 148965 457579 149665
rect 457957 148965 458657 149665
rect 459035 148965 459735 149665
rect 460113 148965 460813 149665
rect 461191 148965 461891 149665
rect 462269 148965 462969 149665
rect 463347 148965 464047 149665
rect 464425 148965 465125 149665
rect 465503 148965 466203 149665
rect 466581 148965 467281 149665
rect 467659 148965 468359 149665
rect 443943 147944 444643 148644
rect 445021 147944 445721 148644
rect 446099 147944 446799 148644
rect 447177 147944 447877 148644
rect 448255 147944 448955 148644
rect 449333 147944 450033 148644
rect 450411 147944 451111 148644
rect 451489 147944 452189 148644
rect 452567 147944 453267 148644
rect 453645 147944 454345 148644
rect 454723 147944 455423 148644
rect 455801 147944 456501 148644
rect 456879 147944 457579 148644
rect 457957 147944 458657 148644
rect 459035 147944 459735 148644
rect 460113 147944 460813 148644
rect 461191 147944 461891 148644
rect 462269 147944 462969 148644
rect 463347 147944 464047 148644
rect 464425 147944 465125 148644
rect 465503 147944 466203 148644
rect 466581 147944 467281 148644
rect 467659 147944 468359 148644
rect 443943 146923 444643 147623
rect 445021 146923 445721 147623
rect 446099 146923 446799 147623
rect 447177 146923 447877 147623
rect 448255 146923 448955 147623
rect 449333 146923 450033 147623
rect 450411 146923 451111 147623
rect 451489 146923 452189 147623
rect 452567 146923 453267 147623
rect 453645 146923 454345 147623
rect 454723 146923 455423 147623
rect 455801 146923 456501 147623
rect 456879 146923 457579 147623
rect 457957 146923 458657 147623
rect 459035 146923 459735 147623
rect 460113 146923 460813 147623
rect 461191 146923 461891 147623
rect 462269 146923 462969 147623
rect 463347 146923 464047 147623
rect 464425 146923 465125 147623
rect 465503 146923 466203 147623
rect 466581 146923 467281 147623
rect 467659 146923 468359 147623
rect 443943 145902 444643 146602
rect 445021 145902 445721 146602
rect 446099 145902 446799 146602
rect 447177 145902 447877 146602
rect 448255 145902 448955 146602
rect 449333 145902 450033 146602
rect 450411 145902 451111 146602
rect 451489 145902 452189 146602
rect 452567 145902 453267 146602
rect 453645 145902 454345 146602
rect 454723 145902 455423 146602
rect 455801 145902 456501 146602
rect 456879 145902 457579 146602
rect 457957 145902 458657 146602
rect 459035 145902 459735 146602
rect 460113 145902 460813 146602
rect 461191 145902 461891 146602
rect 462269 145902 462969 146602
rect 463347 145902 464047 146602
rect 464425 145902 465125 146602
rect 465503 145902 466203 146602
rect 466581 145902 467281 146602
rect 467659 145902 468359 146602
rect 121694 144196 122694 145196
rect 123035 144196 124035 145196
rect 124376 144196 125376 145196
rect 125717 144196 126717 145196
rect 127058 144196 128058 145196
rect 128399 144196 129399 145196
rect 129740 144196 130740 145196
rect 131081 144196 132081 145196
rect 132422 144196 133422 145196
rect 133763 144196 134763 145196
rect 135104 144196 136104 145196
rect 136445 144196 137445 145196
rect 137786 144196 138786 145196
rect 139127 144196 140127 145196
rect 140468 144196 141468 145196
rect 443943 144881 444643 145581
rect 445021 144881 445721 145581
rect 446099 144881 446799 145581
rect 447177 144881 447877 145581
rect 448255 144881 448955 145581
rect 449333 144881 450033 145581
rect 450411 144881 451111 145581
rect 451489 144881 452189 145581
rect 452567 144881 453267 145581
rect 453645 144881 454345 145581
rect 454723 144881 455423 145581
rect 455801 144881 456501 145581
rect 456879 144881 457579 145581
rect 457957 144881 458657 145581
rect 459035 144881 459735 145581
rect 460113 144881 460813 145581
rect 461191 144881 461891 145581
rect 462269 144881 462969 145581
rect 463347 144881 464047 145581
rect 464425 144881 465125 145581
rect 465503 144881 466203 145581
rect 466581 144881 467281 145581
rect 467659 144881 468359 145581
rect 443943 143860 444643 144560
rect 445021 143860 445721 144560
rect 446099 143860 446799 144560
rect 447177 143860 447877 144560
rect 448255 143860 448955 144560
rect 449333 143860 450033 144560
rect 450411 143860 451111 144560
rect 451489 143860 452189 144560
rect 452567 143860 453267 144560
rect 453645 143860 454345 144560
rect 454723 143860 455423 144560
rect 455801 143860 456501 144560
rect 456879 143860 457579 144560
rect 457957 143860 458657 144560
rect 459035 143860 459735 144560
rect 460113 143860 460813 144560
rect 461191 143860 461891 144560
rect 462269 143860 462969 144560
rect 463347 143860 464047 144560
rect 464425 143860 465125 144560
rect 465503 143860 466203 144560
rect 466581 143860 467281 144560
rect 467659 143860 468359 144560
rect 121694 142855 122694 143855
rect 123035 142855 124035 143855
rect 124376 142855 125376 143855
rect 125717 142855 126717 143855
rect 127058 142855 128058 143855
rect 128399 142855 129399 143855
rect 129740 142855 130740 143855
rect 131081 142855 132081 143855
rect 132422 142855 133422 143855
rect 133763 142855 134763 143855
rect 135104 142855 136104 143855
rect 136445 142855 137445 143855
rect 137786 142855 138786 143855
rect 139127 142855 140127 143855
rect 140468 142855 141468 143855
rect 443943 142839 444643 143539
rect 445021 142839 445721 143539
rect 446099 142839 446799 143539
rect 447177 142839 447877 143539
rect 448255 142839 448955 143539
rect 449333 142839 450033 143539
rect 450411 142839 451111 143539
rect 451489 142839 452189 143539
rect 452567 142839 453267 143539
rect 453645 142839 454345 143539
rect 454723 142839 455423 143539
rect 455801 142839 456501 143539
rect 456879 142839 457579 143539
rect 457957 142839 458657 143539
rect 459035 142839 459735 143539
rect 460113 142839 460813 143539
rect 461191 142839 461891 143539
rect 462269 142839 462969 143539
rect 463347 142839 464047 143539
rect 464425 142839 465125 143539
rect 465503 142839 466203 143539
rect 466581 142839 467281 143539
rect 467659 142839 468359 143539
rect 121694 141514 122694 142514
rect 123035 141514 124035 142514
rect 124376 141514 125376 142514
rect 125717 141514 126717 142514
rect 127058 141514 128058 142514
rect 128399 141514 129399 142514
rect 129740 141514 130740 142514
rect 131081 141514 132081 142514
rect 132422 141514 133422 142514
rect 133763 141514 134763 142514
rect 135104 141514 136104 142514
rect 136445 141514 137445 142514
rect 137786 141514 138786 142514
rect 139127 141514 140127 142514
rect 140468 141514 141468 142514
rect 443943 141818 444643 142518
rect 445021 141818 445721 142518
rect 446099 141818 446799 142518
rect 447177 141818 447877 142518
rect 448255 141818 448955 142518
rect 449333 141818 450033 142518
rect 450411 141818 451111 142518
rect 451489 141818 452189 142518
rect 452567 141818 453267 142518
rect 453645 141818 454345 142518
rect 454723 141818 455423 142518
rect 455801 141818 456501 142518
rect 456879 141818 457579 142518
rect 457957 141818 458657 142518
rect 459035 141818 459735 142518
rect 460113 141818 460813 142518
rect 461191 141818 461891 142518
rect 462269 141818 462969 142518
rect 463347 141818 464047 142518
rect 464425 141818 465125 142518
rect 465503 141818 466203 142518
rect 466581 141818 467281 142518
rect 467659 141818 468359 142518
rect 121694 140173 122694 141173
rect 123035 140173 124035 141173
rect 124376 140173 125376 141173
rect 125717 140173 126717 141173
rect 127058 140173 128058 141173
rect 128399 140173 129399 141173
rect 129740 140173 130740 141173
rect 131081 140173 132081 141173
rect 132422 140173 133422 141173
rect 133763 140173 134763 141173
rect 135104 140173 136104 141173
rect 136445 140173 137445 141173
rect 137786 140173 138786 141173
rect 139127 140173 140127 141173
rect 140468 140173 141468 141173
rect 443943 140797 444643 141497
rect 445021 140797 445721 141497
rect 446099 140797 446799 141497
rect 447177 140797 447877 141497
rect 448255 140797 448955 141497
rect 449333 140797 450033 141497
rect 450411 140797 451111 141497
rect 451489 140797 452189 141497
rect 452567 140797 453267 141497
rect 453645 140797 454345 141497
rect 454723 140797 455423 141497
rect 455801 140797 456501 141497
rect 456879 140797 457579 141497
rect 457957 140797 458657 141497
rect 459035 140797 459735 141497
rect 460113 140797 460813 141497
rect 461191 140797 461891 141497
rect 462269 140797 462969 141497
rect 463347 140797 464047 141497
rect 464425 140797 465125 141497
rect 465503 140797 466203 141497
rect 466581 140797 467281 141497
rect 467659 140797 468359 141497
rect 121694 138832 122694 139832
rect 123035 138832 124035 139832
rect 124376 138832 125376 139832
rect 125717 138832 126717 139832
rect 127058 138832 128058 139832
rect 128399 138832 129399 139832
rect 129740 138832 130740 139832
rect 131081 138832 132081 139832
rect 132422 138832 133422 139832
rect 133763 138832 134763 139832
rect 135104 138832 136104 139832
rect 136445 138832 137445 139832
rect 137786 138832 138786 139832
rect 139127 138832 140127 139832
rect 140468 138832 141468 139832
rect 443943 139776 444643 140476
rect 445021 139776 445721 140476
rect 446099 139776 446799 140476
rect 447177 139776 447877 140476
rect 448255 139776 448955 140476
rect 449333 139776 450033 140476
rect 450411 139776 451111 140476
rect 451489 139776 452189 140476
rect 452567 139776 453267 140476
rect 453645 139776 454345 140476
rect 454723 139776 455423 140476
rect 455801 139776 456501 140476
rect 456879 139776 457579 140476
rect 457957 139776 458657 140476
rect 459035 139776 459735 140476
rect 460113 139776 460813 140476
rect 461191 139776 461891 140476
rect 462269 139776 462969 140476
rect 463347 139776 464047 140476
rect 464425 139776 465125 140476
rect 465503 139776 466203 140476
rect 466581 139776 467281 140476
rect 467659 139776 468359 140476
rect 443943 138755 444643 139455
rect 445021 138755 445721 139455
rect 446099 138755 446799 139455
rect 447177 138755 447877 139455
rect 448255 138755 448955 139455
rect 449333 138755 450033 139455
rect 450411 138755 451111 139455
rect 451489 138755 452189 139455
rect 452567 138755 453267 139455
rect 453645 138755 454345 139455
rect 454723 138755 455423 139455
rect 455801 138755 456501 139455
rect 456879 138755 457579 139455
rect 457957 138755 458657 139455
rect 459035 138755 459735 139455
rect 460113 138755 460813 139455
rect 461191 138755 461891 139455
rect 462269 138755 462969 139455
rect 463347 138755 464047 139455
rect 464425 138755 465125 139455
rect 465503 138755 466203 139455
rect 466581 138755 467281 139455
rect 467659 138755 468359 139455
rect 121694 137491 122694 138491
rect 123035 137491 124035 138491
rect 124376 137491 125376 138491
rect 125717 137491 126717 138491
rect 127058 137491 128058 138491
rect 128399 137491 129399 138491
rect 129740 137491 130740 138491
rect 131081 137491 132081 138491
rect 132422 137491 133422 138491
rect 133763 137491 134763 138491
rect 135104 137491 136104 138491
rect 136445 137491 137445 138491
rect 137786 137491 138786 138491
rect 139127 137491 140127 138491
rect 140468 137491 141468 138491
rect 443943 137734 444643 138434
rect 445021 137734 445721 138434
rect 446099 137734 446799 138434
rect 447177 137734 447877 138434
rect 448255 137734 448955 138434
rect 449333 137734 450033 138434
rect 450411 137734 451111 138434
rect 451489 137734 452189 138434
rect 452567 137734 453267 138434
rect 453645 137734 454345 138434
rect 454723 137734 455423 138434
rect 455801 137734 456501 138434
rect 456879 137734 457579 138434
rect 457957 137734 458657 138434
rect 459035 137734 459735 138434
rect 460113 137734 460813 138434
rect 461191 137734 461891 138434
rect 462269 137734 462969 138434
rect 463347 137734 464047 138434
rect 464425 137734 465125 138434
rect 465503 137734 466203 138434
rect 466581 137734 467281 138434
rect 467659 137734 468359 138434
rect 121694 136150 122694 137150
rect 123035 136150 124035 137150
rect 124376 136150 125376 137150
rect 125717 136150 126717 137150
rect 127058 136150 128058 137150
rect 128399 136150 129399 137150
rect 129740 136150 130740 137150
rect 131081 136150 132081 137150
rect 132422 136150 133422 137150
rect 133763 136150 134763 137150
rect 135104 136150 136104 137150
rect 136445 136150 137445 137150
rect 137786 136150 138786 137150
rect 139127 136150 140127 137150
rect 140468 136150 141468 137150
rect 443943 136713 444643 137413
rect 445021 136713 445721 137413
rect 446099 136713 446799 137413
rect 447177 136713 447877 137413
rect 448255 136713 448955 137413
rect 449333 136713 450033 137413
rect 450411 136713 451111 137413
rect 451489 136713 452189 137413
rect 452567 136713 453267 137413
rect 453645 136713 454345 137413
rect 454723 136713 455423 137413
rect 455801 136713 456501 137413
rect 456879 136713 457579 137413
rect 457957 136713 458657 137413
rect 459035 136713 459735 137413
rect 460113 136713 460813 137413
rect 461191 136713 461891 137413
rect 462269 136713 462969 137413
rect 463347 136713 464047 137413
rect 464425 136713 465125 137413
rect 465503 136713 466203 137413
rect 466581 136713 467281 137413
rect 467659 136713 468359 137413
rect 121694 134809 122694 135809
rect 123035 134809 124035 135809
rect 124376 134809 125376 135809
rect 125717 134809 126717 135809
rect 127058 134809 128058 135809
rect 128399 134809 129399 135809
rect 129740 134809 130740 135809
rect 131081 134809 132081 135809
rect 132422 134809 133422 135809
rect 133763 134809 134763 135809
rect 135104 134809 136104 135809
rect 136445 134809 137445 135809
rect 137786 134809 138786 135809
rect 139127 134809 140127 135809
rect 140468 134809 141468 135809
rect 443943 135692 444643 136392
rect 445021 135692 445721 136392
rect 446099 135692 446799 136392
rect 447177 135692 447877 136392
rect 448255 135692 448955 136392
rect 449333 135692 450033 136392
rect 450411 135692 451111 136392
rect 451489 135692 452189 136392
rect 452567 135692 453267 136392
rect 453645 135692 454345 136392
rect 454723 135692 455423 136392
rect 455801 135692 456501 136392
rect 456879 135692 457579 136392
rect 457957 135692 458657 136392
rect 459035 135692 459735 136392
rect 460113 135692 460813 136392
rect 461191 135692 461891 136392
rect 462269 135692 462969 136392
rect 463347 135692 464047 136392
rect 464425 135692 465125 136392
rect 465503 135692 466203 136392
rect 466581 135692 467281 136392
rect 467659 135692 468359 136392
rect 443943 134671 444643 135371
rect 445021 134671 445721 135371
rect 446099 134671 446799 135371
rect 447177 134671 447877 135371
rect 448255 134671 448955 135371
rect 449333 134671 450033 135371
rect 450411 134671 451111 135371
rect 451489 134671 452189 135371
rect 452567 134671 453267 135371
rect 453645 134671 454345 135371
rect 454723 134671 455423 135371
rect 455801 134671 456501 135371
rect 456879 134671 457579 135371
rect 457957 134671 458657 135371
rect 459035 134671 459735 135371
rect 460113 134671 460813 135371
rect 461191 134671 461891 135371
rect 462269 134671 462969 135371
rect 463347 134671 464047 135371
rect 464425 134671 465125 135371
rect 465503 134671 466203 135371
rect 466581 134671 467281 135371
rect 467659 134671 468359 135371
rect 121694 133468 122694 134468
rect 123035 133468 124035 134468
rect 124376 133468 125376 134468
rect 125717 133468 126717 134468
rect 127058 133468 128058 134468
rect 128399 133468 129399 134468
rect 129740 133468 130740 134468
rect 131081 133468 132081 134468
rect 132422 133468 133422 134468
rect 133763 133468 134763 134468
rect 135104 133468 136104 134468
rect 136445 133468 137445 134468
rect 137786 133468 138786 134468
rect 139127 133468 140127 134468
rect 140468 133468 141468 134468
rect 443943 133650 444643 134350
rect 445021 133650 445721 134350
rect 446099 133650 446799 134350
rect 447177 133650 447877 134350
rect 448255 133650 448955 134350
rect 449333 133650 450033 134350
rect 450411 133650 451111 134350
rect 451489 133650 452189 134350
rect 452567 133650 453267 134350
rect 453645 133650 454345 134350
rect 454723 133650 455423 134350
rect 455801 133650 456501 134350
rect 456879 133650 457579 134350
rect 457957 133650 458657 134350
rect 459035 133650 459735 134350
rect 460113 133650 460813 134350
rect 461191 133650 461891 134350
rect 462269 133650 462969 134350
rect 463347 133650 464047 134350
rect 464425 133650 465125 134350
rect 465503 133650 466203 134350
rect 466581 133650 467281 134350
rect 467659 133650 468359 134350
rect 121694 132127 122694 133127
rect 123035 132127 124035 133127
rect 124376 132127 125376 133127
rect 125717 132127 126717 133127
rect 127058 132127 128058 133127
rect 128399 132127 129399 133127
rect 129740 132127 130740 133127
rect 131081 132127 132081 133127
rect 132422 132127 133422 133127
rect 133763 132127 134763 133127
rect 135104 132127 136104 133127
rect 136445 132127 137445 133127
rect 137786 132127 138786 133127
rect 139127 132127 140127 133127
rect 140468 132127 141468 133127
rect 443943 132629 444643 133329
rect 445021 132629 445721 133329
rect 446099 132629 446799 133329
rect 447177 132629 447877 133329
rect 448255 132629 448955 133329
rect 449333 132629 450033 133329
rect 450411 132629 451111 133329
rect 451489 132629 452189 133329
rect 452567 132629 453267 133329
rect 453645 132629 454345 133329
rect 454723 132629 455423 133329
rect 455801 132629 456501 133329
rect 456879 132629 457579 133329
rect 457957 132629 458657 133329
rect 459035 132629 459735 133329
rect 460113 132629 460813 133329
rect 461191 132629 461891 133329
rect 462269 132629 462969 133329
rect 463347 132629 464047 133329
rect 464425 132629 465125 133329
rect 465503 132629 466203 133329
rect 466581 132629 467281 133329
rect 467659 132629 468359 133329
rect 121694 130786 122694 131786
rect 123035 130786 124035 131786
rect 124376 130786 125376 131786
rect 125717 130786 126717 131786
rect 127058 130786 128058 131786
rect 128399 130786 129399 131786
rect 129740 130786 130740 131786
rect 131081 130786 132081 131786
rect 132422 130786 133422 131786
rect 133763 130786 134763 131786
rect 135104 130786 136104 131786
rect 136445 130786 137445 131786
rect 137786 130786 138786 131786
rect 139127 130786 140127 131786
rect 140468 130786 141468 131786
rect 443943 131608 444643 132308
rect 445021 131608 445721 132308
rect 446099 131608 446799 132308
rect 447177 131608 447877 132308
rect 448255 131608 448955 132308
rect 449333 131608 450033 132308
rect 450411 131608 451111 132308
rect 451489 131608 452189 132308
rect 452567 131608 453267 132308
rect 453645 131608 454345 132308
rect 454723 131608 455423 132308
rect 455801 131608 456501 132308
rect 456879 131608 457579 132308
rect 457957 131608 458657 132308
rect 459035 131608 459735 132308
rect 460113 131608 460813 132308
rect 461191 131608 461891 132308
rect 462269 131608 462969 132308
rect 463347 131608 464047 132308
rect 464425 131608 465125 132308
rect 465503 131608 466203 132308
rect 466581 131608 467281 132308
rect 467659 131608 468359 132308
rect 443943 130587 444643 131287
rect 445021 130587 445721 131287
rect 446099 130587 446799 131287
rect 447177 130587 447877 131287
rect 448255 130587 448955 131287
rect 449333 130587 450033 131287
rect 450411 130587 451111 131287
rect 451489 130587 452189 131287
rect 452567 130587 453267 131287
rect 453645 130587 454345 131287
rect 454723 130587 455423 131287
rect 455801 130587 456501 131287
rect 456879 130587 457579 131287
rect 457957 130587 458657 131287
rect 459035 130587 459735 131287
rect 460113 130587 460813 131287
rect 461191 130587 461891 131287
rect 462269 130587 462969 131287
rect 463347 130587 464047 131287
rect 464425 130587 465125 131287
rect 465503 130587 466203 131287
rect 466581 130587 467281 131287
rect 467659 130587 468359 131287
rect 121694 129445 122694 130445
rect 123035 129445 124035 130445
rect 124376 129445 125376 130445
rect 125717 129445 126717 130445
rect 127058 129445 128058 130445
rect 128399 129445 129399 130445
rect 129740 129445 130740 130445
rect 131081 129445 132081 130445
rect 132422 129445 133422 130445
rect 133763 129445 134763 130445
rect 135104 129445 136104 130445
rect 136445 129445 137445 130445
rect 137786 129445 138786 130445
rect 139127 129445 140127 130445
rect 140468 129445 141468 130445
rect 443943 129566 444643 130266
rect 445021 129566 445721 130266
rect 446099 129566 446799 130266
rect 447177 129566 447877 130266
rect 448255 129566 448955 130266
rect 449333 129566 450033 130266
rect 450411 129566 451111 130266
rect 451489 129566 452189 130266
rect 452567 129566 453267 130266
rect 453645 129566 454345 130266
rect 454723 129566 455423 130266
rect 455801 129566 456501 130266
rect 456879 129566 457579 130266
rect 457957 129566 458657 130266
rect 459035 129566 459735 130266
rect 460113 129566 460813 130266
rect 461191 129566 461891 130266
rect 462269 129566 462969 130266
rect 463347 129566 464047 130266
rect 464425 129566 465125 130266
rect 465503 129566 466203 130266
rect 466581 129566 467281 130266
rect 467659 129566 468359 130266
rect 121694 128104 122694 129104
rect 123035 128104 124035 129104
rect 124376 128104 125376 129104
rect 125717 128104 126717 129104
rect 127058 128104 128058 129104
rect 128399 128104 129399 129104
rect 129740 128104 130740 129104
rect 131081 128104 132081 129104
rect 132422 128104 133422 129104
rect 133763 128104 134763 129104
rect 135104 128104 136104 129104
rect 136445 128104 137445 129104
rect 137786 128104 138786 129104
rect 139127 128104 140127 129104
rect 140468 128104 141468 129104
rect 443943 128545 444643 129245
rect 445021 128545 445721 129245
rect 446099 128545 446799 129245
rect 447177 128545 447877 129245
rect 448255 128545 448955 129245
rect 449333 128545 450033 129245
rect 450411 128545 451111 129245
rect 451489 128545 452189 129245
rect 452567 128545 453267 129245
rect 453645 128545 454345 129245
rect 454723 128545 455423 129245
rect 455801 128545 456501 129245
rect 456879 128545 457579 129245
rect 457957 128545 458657 129245
rect 459035 128545 459735 129245
rect 460113 128545 460813 129245
rect 461191 128545 461891 129245
rect 462269 128545 462969 129245
rect 463347 128545 464047 129245
rect 464425 128545 465125 129245
rect 465503 128545 466203 129245
rect 466581 128545 467281 129245
rect 467659 128545 468359 129245
rect 121694 126763 122694 127763
rect 123035 126763 124035 127763
rect 124376 126763 125376 127763
rect 125717 126763 126717 127763
rect 127058 126763 128058 127763
rect 128399 126763 129399 127763
rect 129740 126763 130740 127763
rect 131081 126763 132081 127763
rect 132422 126763 133422 127763
rect 133763 126763 134763 127763
rect 135104 126763 136104 127763
rect 136445 126763 137445 127763
rect 137786 126763 138786 127763
rect 139127 126763 140127 127763
rect 140468 126763 141468 127763
rect 443943 127524 444643 128224
rect 445021 127524 445721 128224
rect 446099 127524 446799 128224
rect 447177 127524 447877 128224
rect 448255 127524 448955 128224
rect 449333 127524 450033 128224
rect 450411 127524 451111 128224
rect 451489 127524 452189 128224
rect 452567 127524 453267 128224
rect 453645 127524 454345 128224
rect 454723 127524 455423 128224
rect 455801 127524 456501 128224
rect 456879 127524 457579 128224
rect 457957 127524 458657 128224
rect 459035 127524 459735 128224
rect 460113 127524 460813 128224
rect 461191 127524 461891 128224
rect 462269 127524 462969 128224
rect 463347 127524 464047 128224
rect 464425 127524 465125 128224
rect 465503 127524 466203 128224
rect 466581 127524 467281 128224
rect 467659 127524 468359 128224
rect 443943 126503 444643 127203
rect 445021 126503 445721 127203
rect 446099 126503 446799 127203
rect 447177 126503 447877 127203
rect 448255 126503 448955 127203
rect 449333 126503 450033 127203
rect 450411 126503 451111 127203
rect 451489 126503 452189 127203
rect 452567 126503 453267 127203
rect 453645 126503 454345 127203
rect 454723 126503 455423 127203
rect 455801 126503 456501 127203
rect 456879 126503 457579 127203
rect 457957 126503 458657 127203
rect 459035 126503 459735 127203
rect 460113 126503 460813 127203
rect 461191 126503 461891 127203
rect 462269 126503 462969 127203
rect 463347 126503 464047 127203
rect 464425 126503 465125 127203
rect 465503 126503 466203 127203
rect 466581 126503 467281 127203
rect 467659 126503 468359 127203
rect 121694 125422 122694 126422
rect 123035 125422 124035 126422
rect 124376 125422 125376 126422
rect 125717 125422 126717 126422
rect 127058 125422 128058 126422
rect 128399 125422 129399 126422
rect 129740 125422 130740 126422
rect 131081 125422 132081 126422
rect 132422 125422 133422 126422
rect 133763 125422 134763 126422
rect 135104 125422 136104 126422
rect 136445 125422 137445 126422
rect 137786 125422 138786 126422
rect 139127 125422 140127 126422
rect 140468 125422 141468 126422
rect 443943 125482 444643 126182
rect 445021 125482 445721 126182
rect 446099 125482 446799 126182
rect 447177 125482 447877 126182
rect 448255 125482 448955 126182
rect 449333 125482 450033 126182
rect 450411 125482 451111 126182
rect 451489 125482 452189 126182
rect 452567 125482 453267 126182
rect 453645 125482 454345 126182
rect 454723 125482 455423 126182
rect 455801 125482 456501 126182
rect 456879 125482 457579 126182
rect 457957 125482 458657 126182
rect 459035 125482 459735 126182
rect 460113 125482 460813 126182
rect 461191 125482 461891 126182
rect 462269 125482 462969 126182
rect 463347 125482 464047 126182
rect 464425 125482 465125 126182
rect 465503 125482 466203 126182
rect 466581 125482 467281 126182
rect 467659 125482 468359 126182
rect 482072 124124 482772 124824
rect 483168 124124 483868 124824
rect 484264 124124 484964 124824
rect 485360 124124 486060 124824
rect 486456 124124 487156 124824
rect 487552 124124 488252 124824
rect 488648 124124 489348 124824
rect 489744 124124 490444 124824
rect 490840 124124 491540 124824
rect 491936 124124 492636 124824
rect 493032 124124 493732 124824
rect 494128 124124 494828 124824
rect 495224 124124 495924 124824
rect 496320 124124 497020 124824
rect 497416 124124 498116 124824
rect 498512 124124 499212 124824
rect 499608 124124 500308 124824
rect 500704 124124 501404 124824
rect 501800 124124 502500 124824
rect 502896 124124 503596 124824
rect 503992 124124 504692 124824
rect 505088 124124 505788 124824
rect 506184 124124 506884 124824
rect 507280 124124 507980 124824
rect 482072 122973 482772 123673
rect 483168 122973 483868 123673
rect 484264 122973 484964 123673
rect 485360 122973 486060 123673
rect 486456 122973 487156 123673
rect 487552 122973 488252 123673
rect 488648 122973 489348 123673
rect 489744 122973 490444 123673
rect 490840 122973 491540 123673
rect 491936 122973 492636 123673
rect 493032 122973 493732 123673
rect 494128 122973 494828 123673
rect 495224 122973 495924 123673
rect 496320 122973 497020 123673
rect 497416 122973 498116 123673
rect 498512 122973 499212 123673
rect 499608 122973 500308 123673
rect 500704 122973 501404 123673
rect 501800 122973 502500 123673
rect 502896 122973 503596 123673
rect 503992 122973 504692 123673
rect 505088 122973 505788 123673
rect 506184 122973 506884 123673
rect 507280 122973 507980 123673
rect 482072 121822 482772 122522
rect 483168 121822 483868 122522
rect 484264 121822 484964 122522
rect 485360 121822 486060 122522
rect 486456 121822 487156 122522
rect 487552 121822 488252 122522
rect 488648 121822 489348 122522
rect 489744 121822 490444 122522
rect 490840 121822 491540 122522
rect 491936 121822 492636 122522
rect 493032 121822 493732 122522
rect 494128 121822 494828 122522
rect 495224 121822 495924 122522
rect 496320 121822 497020 122522
rect 497416 121822 498116 122522
rect 498512 121822 499212 122522
rect 499608 121822 500308 122522
rect 500704 121822 501404 122522
rect 501800 121822 502500 122522
rect 502896 121822 503596 122522
rect 503992 121822 504692 122522
rect 505088 121822 505788 122522
rect 506184 121822 506884 122522
rect 507280 121822 507980 122522
rect 482072 120671 482772 121371
rect 483168 120671 483868 121371
rect 484264 120671 484964 121371
rect 485360 120671 486060 121371
rect 486456 120671 487156 121371
rect 487552 120671 488252 121371
rect 488648 120671 489348 121371
rect 489744 120671 490444 121371
rect 490840 120671 491540 121371
rect 491936 120671 492636 121371
rect 493032 120671 493732 121371
rect 494128 120671 494828 121371
rect 495224 120671 495924 121371
rect 496320 120671 497020 121371
rect 497416 120671 498116 121371
rect 498512 120671 499212 121371
rect 499608 120671 500308 121371
rect 500704 120671 501404 121371
rect 501800 120671 502500 121371
rect 502896 120671 503596 121371
rect 503992 120671 504692 121371
rect 505088 120671 505788 121371
rect 506184 120671 506884 121371
rect 507280 120671 507980 121371
rect 89225 119146 89925 119846
rect 90134 119146 90834 119846
rect 91043 119146 91743 119846
rect 91952 119146 92652 119846
rect 92861 119146 93561 119846
rect 93770 119146 94470 119846
rect 94679 119146 95379 119846
rect 95588 119146 96288 119846
rect 96497 119146 97197 119846
rect 97406 119146 98106 119846
rect 98315 119146 99015 119846
rect 99224 119146 99924 119846
rect 100133 119146 100833 119846
rect 101042 119146 101742 119846
rect 101951 119146 102651 119846
rect 102860 119146 103560 119846
rect 103769 119146 104469 119846
rect 104678 119146 105378 119846
rect 105587 119146 106287 119846
rect 106496 119146 107196 119846
rect 107405 119146 108105 119846
rect 108314 119146 109014 119846
rect 109223 119146 109923 119846
rect 110132 119146 110832 119846
rect 89225 118258 89925 118958
rect 90134 118258 90834 118958
rect 91043 118258 91743 118958
rect 91952 118258 92652 118958
rect 92861 118258 93561 118958
rect 93770 118258 94470 118958
rect 94679 118258 95379 118958
rect 95588 118258 96288 118958
rect 96497 118258 97197 118958
rect 97406 118258 98106 118958
rect 98315 118258 99015 118958
rect 99224 118258 99924 118958
rect 100133 118258 100833 118958
rect 101042 118258 101742 118958
rect 101951 118258 102651 118958
rect 102860 118258 103560 118958
rect 103769 118258 104469 118958
rect 104678 118258 105378 118958
rect 105587 118258 106287 118958
rect 106496 118258 107196 118958
rect 107405 118258 108105 118958
rect 108314 118258 109014 118958
rect 109223 118258 109923 118958
rect 110132 118258 110832 118958
rect 482072 119520 482772 120220
rect 483168 119520 483868 120220
rect 484264 119520 484964 120220
rect 485360 119520 486060 120220
rect 486456 119520 487156 120220
rect 487552 119520 488252 120220
rect 488648 119520 489348 120220
rect 489744 119520 490444 120220
rect 490840 119520 491540 120220
rect 491936 119520 492636 120220
rect 493032 119520 493732 120220
rect 494128 119520 494828 120220
rect 495224 119520 495924 120220
rect 496320 119520 497020 120220
rect 497416 119520 498116 120220
rect 498512 119520 499212 120220
rect 499608 119520 500308 120220
rect 500704 119520 501404 120220
rect 501800 119520 502500 120220
rect 502896 119520 503596 120220
rect 503992 119520 504692 120220
rect 505088 119520 505788 120220
rect 506184 119520 506884 120220
rect 507280 119520 507980 120220
rect 482072 118369 482772 119069
rect 483168 118369 483868 119069
rect 484264 118369 484964 119069
rect 485360 118369 486060 119069
rect 486456 118369 487156 119069
rect 487552 118369 488252 119069
rect 488648 118369 489348 119069
rect 489744 118369 490444 119069
rect 490840 118369 491540 119069
rect 491936 118369 492636 119069
rect 493032 118369 493732 119069
rect 494128 118369 494828 119069
rect 495224 118369 495924 119069
rect 496320 118369 497020 119069
rect 497416 118369 498116 119069
rect 498512 118369 499212 119069
rect 499608 118369 500308 119069
rect 500704 118369 501404 119069
rect 501800 118369 502500 119069
rect 502896 118369 503596 119069
rect 503992 118369 504692 119069
rect 505088 118369 505788 119069
rect 506184 118369 506884 119069
rect 507280 118369 507980 119069
rect 89225 117370 89925 118070
rect 90134 117370 90834 118070
rect 91043 117370 91743 118070
rect 91952 117370 92652 118070
rect 92861 117370 93561 118070
rect 93770 117370 94470 118070
rect 94679 117370 95379 118070
rect 95588 117370 96288 118070
rect 96497 117370 97197 118070
rect 97406 117370 98106 118070
rect 98315 117370 99015 118070
rect 99224 117370 99924 118070
rect 100133 117370 100833 118070
rect 101042 117370 101742 118070
rect 101951 117370 102651 118070
rect 102860 117370 103560 118070
rect 103769 117370 104469 118070
rect 104678 117370 105378 118070
rect 105587 117370 106287 118070
rect 106496 117370 107196 118070
rect 107405 117370 108105 118070
rect 108314 117370 109014 118070
rect 109223 117370 109923 118070
rect 110132 117370 110832 118070
rect 482072 117218 482772 117918
rect 483168 117218 483868 117918
rect 484264 117218 484964 117918
rect 485360 117218 486060 117918
rect 486456 117218 487156 117918
rect 487552 117218 488252 117918
rect 488648 117218 489348 117918
rect 489744 117218 490444 117918
rect 490840 117218 491540 117918
rect 491936 117218 492636 117918
rect 493032 117218 493732 117918
rect 494128 117218 494828 117918
rect 495224 117218 495924 117918
rect 496320 117218 497020 117918
rect 497416 117218 498116 117918
rect 498512 117218 499212 117918
rect 499608 117218 500308 117918
rect 500704 117218 501404 117918
rect 501800 117218 502500 117918
rect 502896 117218 503596 117918
rect 503992 117218 504692 117918
rect 505088 117218 505788 117918
rect 506184 117218 506884 117918
rect 507280 117218 507980 117918
rect 89225 116482 89925 117182
rect 90134 116482 90834 117182
rect 91043 116482 91743 117182
rect 91952 116482 92652 117182
rect 92861 116482 93561 117182
rect 93770 116482 94470 117182
rect 94679 116482 95379 117182
rect 95588 116482 96288 117182
rect 96497 116482 97197 117182
rect 97406 116482 98106 117182
rect 98315 116482 99015 117182
rect 99224 116482 99924 117182
rect 100133 116482 100833 117182
rect 101042 116482 101742 117182
rect 101951 116482 102651 117182
rect 102860 116482 103560 117182
rect 103769 116482 104469 117182
rect 104678 116482 105378 117182
rect 105587 116482 106287 117182
rect 106496 116482 107196 117182
rect 107405 116482 108105 117182
rect 108314 116482 109014 117182
rect 109223 116482 109923 117182
rect 110132 116482 110832 117182
rect 89225 115594 89925 116294
rect 90134 115594 90834 116294
rect 91043 115594 91743 116294
rect 91952 115594 92652 116294
rect 92861 115594 93561 116294
rect 93770 115594 94470 116294
rect 94679 115594 95379 116294
rect 95588 115594 96288 116294
rect 96497 115594 97197 116294
rect 97406 115594 98106 116294
rect 98315 115594 99015 116294
rect 99224 115594 99924 116294
rect 100133 115594 100833 116294
rect 101042 115594 101742 116294
rect 101951 115594 102651 116294
rect 102860 115594 103560 116294
rect 103769 115594 104469 116294
rect 104678 115594 105378 116294
rect 105587 115594 106287 116294
rect 106496 115594 107196 116294
rect 107405 115594 108105 116294
rect 108314 115594 109014 116294
rect 109223 115594 109923 116294
rect 110132 115594 110832 116294
rect 482072 116067 482772 116767
rect 483168 116067 483868 116767
rect 484264 116067 484964 116767
rect 485360 116067 486060 116767
rect 486456 116067 487156 116767
rect 487552 116067 488252 116767
rect 488648 116067 489348 116767
rect 489744 116067 490444 116767
rect 490840 116067 491540 116767
rect 491936 116067 492636 116767
rect 493032 116067 493732 116767
rect 494128 116067 494828 116767
rect 495224 116067 495924 116767
rect 496320 116067 497020 116767
rect 497416 116067 498116 116767
rect 498512 116067 499212 116767
rect 499608 116067 500308 116767
rect 500704 116067 501404 116767
rect 501800 116067 502500 116767
rect 502896 116067 503596 116767
rect 503992 116067 504692 116767
rect 505088 116067 505788 116767
rect 506184 116067 506884 116767
rect 507280 116067 507980 116767
rect 89225 114706 89925 115406
rect 90134 114706 90834 115406
rect 91043 114706 91743 115406
rect 91952 114706 92652 115406
rect 92861 114706 93561 115406
rect 93770 114706 94470 115406
rect 94679 114706 95379 115406
rect 95588 114706 96288 115406
rect 96497 114706 97197 115406
rect 97406 114706 98106 115406
rect 98315 114706 99015 115406
rect 99224 114706 99924 115406
rect 100133 114706 100833 115406
rect 101042 114706 101742 115406
rect 101951 114706 102651 115406
rect 102860 114706 103560 115406
rect 103769 114706 104469 115406
rect 104678 114706 105378 115406
rect 105587 114706 106287 115406
rect 106496 114706 107196 115406
rect 107405 114706 108105 115406
rect 108314 114706 109014 115406
rect 109223 114706 109923 115406
rect 110132 114706 110832 115406
rect 482072 114916 482772 115616
rect 483168 114916 483868 115616
rect 484264 114916 484964 115616
rect 485360 114916 486060 115616
rect 486456 114916 487156 115616
rect 487552 114916 488252 115616
rect 488648 114916 489348 115616
rect 489744 114916 490444 115616
rect 490840 114916 491540 115616
rect 491936 114916 492636 115616
rect 493032 114916 493732 115616
rect 494128 114916 494828 115616
rect 495224 114916 495924 115616
rect 496320 114916 497020 115616
rect 497416 114916 498116 115616
rect 498512 114916 499212 115616
rect 499608 114916 500308 115616
rect 500704 114916 501404 115616
rect 501800 114916 502500 115616
rect 502896 114916 503596 115616
rect 503992 114916 504692 115616
rect 505088 114916 505788 115616
rect 506184 114916 506884 115616
rect 507280 114916 507980 115616
rect 89225 113818 89925 114518
rect 90134 113818 90834 114518
rect 91043 113818 91743 114518
rect 91952 113818 92652 114518
rect 92861 113818 93561 114518
rect 93770 113818 94470 114518
rect 94679 113818 95379 114518
rect 95588 113818 96288 114518
rect 96497 113818 97197 114518
rect 97406 113818 98106 114518
rect 98315 113818 99015 114518
rect 99224 113818 99924 114518
rect 100133 113818 100833 114518
rect 101042 113818 101742 114518
rect 101951 113818 102651 114518
rect 102860 113818 103560 114518
rect 103769 113818 104469 114518
rect 104678 113818 105378 114518
rect 105587 113818 106287 114518
rect 106496 113818 107196 114518
rect 107405 113818 108105 114518
rect 108314 113818 109014 114518
rect 109223 113818 109923 114518
rect 110132 113818 110832 114518
rect 482072 113765 482772 114465
rect 483168 113765 483868 114465
rect 484264 113765 484964 114465
rect 485360 113765 486060 114465
rect 486456 113765 487156 114465
rect 487552 113765 488252 114465
rect 488648 113765 489348 114465
rect 489744 113765 490444 114465
rect 490840 113765 491540 114465
rect 491936 113765 492636 114465
rect 493032 113765 493732 114465
rect 494128 113765 494828 114465
rect 495224 113765 495924 114465
rect 496320 113765 497020 114465
rect 497416 113765 498116 114465
rect 498512 113765 499212 114465
rect 499608 113765 500308 114465
rect 500704 113765 501404 114465
rect 501800 113765 502500 114465
rect 502896 113765 503596 114465
rect 503992 113765 504692 114465
rect 505088 113765 505788 114465
rect 506184 113765 506884 114465
rect 507280 113765 507980 114465
rect 89225 112930 89925 113630
rect 90134 112930 90834 113630
rect 91043 112930 91743 113630
rect 91952 112930 92652 113630
rect 92861 112930 93561 113630
rect 93770 112930 94470 113630
rect 94679 112930 95379 113630
rect 95588 112930 96288 113630
rect 96497 112930 97197 113630
rect 97406 112930 98106 113630
rect 98315 112930 99015 113630
rect 99224 112930 99924 113630
rect 100133 112930 100833 113630
rect 101042 112930 101742 113630
rect 101951 112930 102651 113630
rect 102860 112930 103560 113630
rect 103769 112930 104469 113630
rect 104678 112930 105378 113630
rect 105587 112930 106287 113630
rect 106496 112930 107196 113630
rect 107405 112930 108105 113630
rect 108314 112930 109014 113630
rect 109223 112930 109923 113630
rect 110132 112930 110832 113630
rect 89225 112042 89925 112742
rect 90134 112042 90834 112742
rect 91043 112042 91743 112742
rect 91952 112042 92652 112742
rect 92861 112042 93561 112742
rect 93770 112042 94470 112742
rect 94679 112042 95379 112742
rect 95588 112042 96288 112742
rect 96497 112042 97197 112742
rect 97406 112042 98106 112742
rect 98315 112042 99015 112742
rect 99224 112042 99924 112742
rect 100133 112042 100833 112742
rect 101042 112042 101742 112742
rect 101951 112042 102651 112742
rect 102860 112042 103560 112742
rect 103769 112042 104469 112742
rect 104678 112042 105378 112742
rect 105587 112042 106287 112742
rect 106496 112042 107196 112742
rect 107405 112042 108105 112742
rect 108314 112042 109014 112742
rect 109223 112042 109923 112742
rect 110132 112042 110832 112742
rect 482072 112614 482772 113314
rect 483168 112614 483868 113314
rect 484264 112614 484964 113314
rect 485360 112614 486060 113314
rect 486456 112614 487156 113314
rect 487552 112614 488252 113314
rect 488648 112614 489348 113314
rect 489744 112614 490444 113314
rect 490840 112614 491540 113314
rect 491936 112614 492636 113314
rect 493032 112614 493732 113314
rect 494128 112614 494828 113314
rect 495224 112614 495924 113314
rect 496320 112614 497020 113314
rect 497416 112614 498116 113314
rect 498512 112614 499212 113314
rect 499608 112614 500308 113314
rect 500704 112614 501404 113314
rect 501800 112614 502500 113314
rect 502896 112614 503596 113314
rect 503992 112614 504692 113314
rect 505088 112614 505788 113314
rect 506184 112614 506884 113314
rect 507280 112614 507980 113314
rect 89225 111154 89925 111854
rect 90134 111154 90834 111854
rect 91043 111154 91743 111854
rect 91952 111154 92652 111854
rect 92861 111154 93561 111854
rect 93770 111154 94470 111854
rect 94679 111154 95379 111854
rect 95588 111154 96288 111854
rect 96497 111154 97197 111854
rect 97406 111154 98106 111854
rect 98315 111154 99015 111854
rect 99224 111154 99924 111854
rect 100133 111154 100833 111854
rect 101042 111154 101742 111854
rect 101951 111154 102651 111854
rect 102860 111154 103560 111854
rect 103769 111154 104469 111854
rect 104678 111154 105378 111854
rect 105587 111154 106287 111854
rect 106496 111154 107196 111854
rect 107405 111154 108105 111854
rect 108314 111154 109014 111854
rect 109223 111154 109923 111854
rect 110132 111154 110832 111854
rect 482072 111463 482772 112163
rect 483168 111463 483868 112163
rect 484264 111463 484964 112163
rect 485360 111463 486060 112163
rect 486456 111463 487156 112163
rect 487552 111463 488252 112163
rect 488648 111463 489348 112163
rect 489744 111463 490444 112163
rect 490840 111463 491540 112163
rect 491936 111463 492636 112163
rect 493032 111463 493732 112163
rect 494128 111463 494828 112163
rect 495224 111463 495924 112163
rect 496320 111463 497020 112163
rect 497416 111463 498116 112163
rect 498512 111463 499212 112163
rect 499608 111463 500308 112163
rect 500704 111463 501404 112163
rect 501800 111463 502500 112163
rect 502896 111463 503596 112163
rect 503992 111463 504692 112163
rect 505088 111463 505788 112163
rect 506184 111463 506884 112163
rect 507280 111463 507980 112163
rect 89225 110266 89925 110966
rect 90134 110266 90834 110966
rect 91043 110266 91743 110966
rect 91952 110266 92652 110966
rect 92861 110266 93561 110966
rect 93770 110266 94470 110966
rect 94679 110266 95379 110966
rect 95588 110266 96288 110966
rect 96497 110266 97197 110966
rect 97406 110266 98106 110966
rect 98315 110266 99015 110966
rect 99224 110266 99924 110966
rect 100133 110266 100833 110966
rect 101042 110266 101742 110966
rect 101951 110266 102651 110966
rect 102860 110266 103560 110966
rect 103769 110266 104469 110966
rect 104678 110266 105378 110966
rect 105587 110266 106287 110966
rect 106496 110266 107196 110966
rect 107405 110266 108105 110966
rect 108314 110266 109014 110966
rect 109223 110266 109923 110966
rect 110132 110266 110832 110966
rect 482072 110312 482772 111012
rect 483168 110312 483868 111012
rect 484264 110312 484964 111012
rect 485360 110312 486060 111012
rect 486456 110312 487156 111012
rect 487552 110312 488252 111012
rect 488648 110312 489348 111012
rect 489744 110312 490444 111012
rect 490840 110312 491540 111012
rect 491936 110312 492636 111012
rect 493032 110312 493732 111012
rect 494128 110312 494828 111012
rect 495224 110312 495924 111012
rect 496320 110312 497020 111012
rect 497416 110312 498116 111012
rect 498512 110312 499212 111012
rect 499608 110312 500308 111012
rect 500704 110312 501404 111012
rect 501800 110312 502500 111012
rect 502896 110312 503596 111012
rect 503992 110312 504692 111012
rect 505088 110312 505788 111012
rect 506184 110312 506884 111012
rect 507280 110312 507980 111012
rect 89225 109378 89925 110078
rect 90134 109378 90834 110078
rect 91043 109378 91743 110078
rect 91952 109378 92652 110078
rect 92861 109378 93561 110078
rect 93770 109378 94470 110078
rect 94679 109378 95379 110078
rect 95588 109378 96288 110078
rect 96497 109378 97197 110078
rect 97406 109378 98106 110078
rect 98315 109378 99015 110078
rect 99224 109378 99924 110078
rect 100133 109378 100833 110078
rect 101042 109378 101742 110078
rect 101951 109378 102651 110078
rect 102860 109378 103560 110078
rect 103769 109378 104469 110078
rect 104678 109378 105378 110078
rect 105587 109378 106287 110078
rect 106496 109378 107196 110078
rect 107405 109378 108105 110078
rect 108314 109378 109014 110078
rect 109223 109378 109923 110078
rect 110132 109378 110832 110078
rect 89225 108490 89925 109190
rect 90134 108490 90834 109190
rect 91043 108490 91743 109190
rect 91952 108490 92652 109190
rect 92861 108490 93561 109190
rect 93770 108490 94470 109190
rect 94679 108490 95379 109190
rect 95588 108490 96288 109190
rect 96497 108490 97197 109190
rect 97406 108490 98106 109190
rect 98315 108490 99015 109190
rect 99224 108490 99924 109190
rect 100133 108490 100833 109190
rect 101042 108490 101742 109190
rect 101951 108490 102651 109190
rect 102860 108490 103560 109190
rect 103769 108490 104469 109190
rect 104678 108490 105378 109190
rect 105587 108490 106287 109190
rect 106496 108490 107196 109190
rect 107405 108490 108105 109190
rect 108314 108490 109014 109190
rect 109223 108490 109923 109190
rect 110132 108490 110832 109190
rect 482072 109161 482772 109861
rect 483168 109161 483868 109861
rect 484264 109161 484964 109861
rect 485360 109161 486060 109861
rect 486456 109161 487156 109861
rect 487552 109161 488252 109861
rect 488648 109161 489348 109861
rect 489744 109161 490444 109861
rect 490840 109161 491540 109861
rect 491936 109161 492636 109861
rect 493032 109161 493732 109861
rect 494128 109161 494828 109861
rect 495224 109161 495924 109861
rect 496320 109161 497020 109861
rect 497416 109161 498116 109861
rect 498512 109161 499212 109861
rect 499608 109161 500308 109861
rect 500704 109161 501404 109861
rect 501800 109161 502500 109861
rect 502896 109161 503596 109861
rect 503992 109161 504692 109861
rect 505088 109161 505788 109861
rect 506184 109161 506884 109861
rect 507280 109161 507980 109861
rect 89225 107602 89925 108302
rect 90134 107602 90834 108302
rect 91043 107602 91743 108302
rect 91952 107602 92652 108302
rect 92861 107602 93561 108302
rect 93770 107602 94470 108302
rect 94679 107602 95379 108302
rect 95588 107602 96288 108302
rect 96497 107602 97197 108302
rect 97406 107602 98106 108302
rect 98315 107602 99015 108302
rect 99224 107602 99924 108302
rect 100133 107602 100833 108302
rect 101042 107602 101742 108302
rect 101951 107602 102651 108302
rect 102860 107602 103560 108302
rect 103769 107602 104469 108302
rect 104678 107602 105378 108302
rect 105587 107602 106287 108302
rect 106496 107602 107196 108302
rect 107405 107602 108105 108302
rect 108314 107602 109014 108302
rect 109223 107602 109923 108302
rect 110132 107602 110832 108302
rect 482072 108010 482772 108710
rect 483168 108010 483868 108710
rect 484264 108010 484964 108710
rect 485360 108010 486060 108710
rect 486456 108010 487156 108710
rect 487552 108010 488252 108710
rect 488648 108010 489348 108710
rect 489744 108010 490444 108710
rect 490840 108010 491540 108710
rect 491936 108010 492636 108710
rect 493032 108010 493732 108710
rect 494128 108010 494828 108710
rect 495224 108010 495924 108710
rect 496320 108010 497020 108710
rect 497416 108010 498116 108710
rect 498512 108010 499212 108710
rect 499608 108010 500308 108710
rect 500704 108010 501404 108710
rect 501800 108010 502500 108710
rect 502896 108010 503596 108710
rect 503992 108010 504692 108710
rect 505088 108010 505788 108710
rect 506184 108010 506884 108710
rect 507280 108010 507980 108710
rect 89225 106714 89925 107414
rect 90134 106714 90834 107414
rect 91043 106714 91743 107414
rect 91952 106714 92652 107414
rect 92861 106714 93561 107414
rect 93770 106714 94470 107414
rect 94679 106714 95379 107414
rect 95588 106714 96288 107414
rect 96497 106714 97197 107414
rect 97406 106714 98106 107414
rect 98315 106714 99015 107414
rect 99224 106714 99924 107414
rect 100133 106714 100833 107414
rect 101042 106714 101742 107414
rect 101951 106714 102651 107414
rect 102860 106714 103560 107414
rect 103769 106714 104469 107414
rect 104678 106714 105378 107414
rect 105587 106714 106287 107414
rect 106496 106714 107196 107414
rect 107405 106714 108105 107414
rect 108314 106714 109014 107414
rect 109223 106714 109923 107414
rect 110132 106714 110832 107414
rect 482072 106859 482772 107559
rect 483168 106859 483868 107559
rect 484264 106859 484964 107559
rect 485360 106859 486060 107559
rect 486456 106859 487156 107559
rect 487552 106859 488252 107559
rect 488648 106859 489348 107559
rect 489744 106859 490444 107559
rect 490840 106859 491540 107559
rect 491936 106859 492636 107559
rect 493032 106859 493732 107559
rect 494128 106859 494828 107559
rect 495224 106859 495924 107559
rect 496320 106859 497020 107559
rect 497416 106859 498116 107559
rect 498512 106859 499212 107559
rect 499608 106859 500308 107559
rect 500704 106859 501404 107559
rect 501800 106859 502500 107559
rect 502896 106859 503596 107559
rect 503992 106859 504692 107559
rect 505088 106859 505788 107559
rect 506184 106859 506884 107559
rect 507280 106859 507980 107559
rect 89225 105826 89925 106526
rect 90134 105826 90834 106526
rect 91043 105826 91743 106526
rect 91952 105826 92652 106526
rect 92861 105826 93561 106526
rect 93770 105826 94470 106526
rect 94679 105826 95379 106526
rect 95588 105826 96288 106526
rect 96497 105826 97197 106526
rect 97406 105826 98106 106526
rect 98315 105826 99015 106526
rect 99224 105826 99924 106526
rect 100133 105826 100833 106526
rect 101042 105826 101742 106526
rect 101951 105826 102651 106526
rect 102860 105826 103560 106526
rect 103769 105826 104469 106526
rect 104678 105826 105378 106526
rect 105587 105826 106287 106526
rect 106496 105826 107196 106526
rect 107405 105826 108105 106526
rect 108314 105826 109014 106526
rect 109223 105826 109923 106526
rect 110132 105826 110832 106526
rect 482072 105708 482772 106408
rect 483168 105708 483868 106408
rect 484264 105708 484964 106408
rect 485360 105708 486060 106408
rect 486456 105708 487156 106408
rect 487552 105708 488252 106408
rect 488648 105708 489348 106408
rect 489744 105708 490444 106408
rect 490840 105708 491540 106408
rect 491936 105708 492636 106408
rect 493032 105708 493732 106408
rect 494128 105708 494828 106408
rect 495224 105708 495924 106408
rect 496320 105708 497020 106408
rect 497416 105708 498116 106408
rect 498512 105708 499212 106408
rect 499608 105708 500308 106408
rect 500704 105708 501404 106408
rect 501800 105708 502500 106408
rect 502896 105708 503596 106408
rect 503992 105708 504692 106408
rect 505088 105708 505788 106408
rect 506184 105708 506884 106408
rect 507280 105708 507980 106408
rect 89225 104938 89925 105638
rect 90134 104938 90834 105638
rect 91043 104938 91743 105638
rect 91952 104938 92652 105638
rect 92861 104938 93561 105638
rect 93770 104938 94470 105638
rect 94679 104938 95379 105638
rect 95588 104938 96288 105638
rect 96497 104938 97197 105638
rect 97406 104938 98106 105638
rect 98315 104938 99015 105638
rect 99224 104938 99924 105638
rect 100133 104938 100833 105638
rect 101042 104938 101742 105638
rect 101951 104938 102651 105638
rect 102860 104938 103560 105638
rect 103769 104938 104469 105638
rect 104678 104938 105378 105638
rect 105587 104938 106287 105638
rect 106496 104938 107196 105638
rect 107405 104938 108105 105638
rect 108314 104938 109014 105638
rect 109223 104938 109923 105638
rect 110132 104938 110832 105638
rect 89225 104050 89925 104750
rect 90134 104050 90834 104750
rect 91043 104050 91743 104750
rect 91952 104050 92652 104750
rect 92861 104050 93561 104750
rect 93770 104050 94470 104750
rect 94679 104050 95379 104750
rect 95588 104050 96288 104750
rect 96497 104050 97197 104750
rect 97406 104050 98106 104750
rect 98315 104050 99015 104750
rect 99224 104050 99924 104750
rect 100133 104050 100833 104750
rect 101042 104050 101742 104750
rect 101951 104050 102651 104750
rect 102860 104050 103560 104750
rect 103769 104050 104469 104750
rect 104678 104050 105378 104750
rect 105587 104050 106287 104750
rect 106496 104050 107196 104750
rect 107405 104050 108105 104750
rect 108314 104050 109014 104750
rect 109223 104050 109923 104750
rect 110132 104050 110832 104750
rect 482072 104557 482772 105257
rect 483168 104557 483868 105257
rect 484264 104557 484964 105257
rect 485360 104557 486060 105257
rect 486456 104557 487156 105257
rect 487552 104557 488252 105257
rect 488648 104557 489348 105257
rect 489744 104557 490444 105257
rect 490840 104557 491540 105257
rect 491936 104557 492636 105257
rect 493032 104557 493732 105257
rect 494128 104557 494828 105257
rect 495224 104557 495924 105257
rect 496320 104557 497020 105257
rect 497416 104557 498116 105257
rect 498512 104557 499212 105257
rect 499608 104557 500308 105257
rect 500704 104557 501404 105257
rect 501800 104557 502500 105257
rect 502896 104557 503596 105257
rect 503992 104557 504692 105257
rect 505088 104557 505788 105257
rect 506184 104557 506884 105257
rect 507280 104557 507980 105257
rect 89225 103162 89925 103862
rect 90134 103162 90834 103862
rect 91043 103162 91743 103862
rect 91952 103162 92652 103862
rect 92861 103162 93561 103862
rect 93770 103162 94470 103862
rect 94679 103162 95379 103862
rect 95588 103162 96288 103862
rect 96497 103162 97197 103862
rect 97406 103162 98106 103862
rect 98315 103162 99015 103862
rect 99224 103162 99924 103862
rect 100133 103162 100833 103862
rect 101042 103162 101742 103862
rect 101951 103162 102651 103862
rect 102860 103162 103560 103862
rect 103769 103162 104469 103862
rect 104678 103162 105378 103862
rect 105587 103162 106287 103862
rect 106496 103162 107196 103862
rect 107405 103162 108105 103862
rect 108314 103162 109014 103862
rect 109223 103162 109923 103862
rect 110132 103162 110832 103862
rect 482072 103406 482772 104106
rect 483168 103406 483868 104106
rect 484264 103406 484964 104106
rect 485360 103406 486060 104106
rect 486456 103406 487156 104106
rect 487552 103406 488252 104106
rect 488648 103406 489348 104106
rect 489744 103406 490444 104106
rect 490840 103406 491540 104106
rect 491936 103406 492636 104106
rect 493032 103406 493732 104106
rect 494128 103406 494828 104106
rect 495224 103406 495924 104106
rect 496320 103406 497020 104106
rect 497416 103406 498116 104106
rect 498512 103406 499212 104106
rect 499608 103406 500308 104106
rect 500704 103406 501404 104106
rect 501800 103406 502500 104106
rect 502896 103406 503596 104106
rect 503992 103406 504692 104106
rect 505088 103406 505788 104106
rect 506184 103406 506884 104106
rect 507280 103406 507980 104106
rect 89225 102274 89925 102974
rect 90134 102274 90834 102974
rect 91043 102274 91743 102974
rect 91952 102274 92652 102974
rect 92861 102274 93561 102974
rect 93770 102274 94470 102974
rect 94679 102274 95379 102974
rect 95588 102274 96288 102974
rect 96497 102274 97197 102974
rect 97406 102274 98106 102974
rect 98315 102274 99015 102974
rect 99224 102274 99924 102974
rect 100133 102274 100833 102974
rect 101042 102274 101742 102974
rect 101951 102274 102651 102974
rect 102860 102274 103560 102974
rect 103769 102274 104469 102974
rect 104678 102274 105378 102974
rect 105587 102274 106287 102974
rect 106496 102274 107196 102974
rect 107405 102274 108105 102974
rect 108314 102274 109014 102974
rect 109223 102274 109923 102974
rect 110132 102274 110832 102974
rect 89225 101386 89925 102086
rect 90134 101386 90834 102086
rect 91043 101386 91743 102086
rect 91952 101386 92652 102086
rect 92861 101386 93561 102086
rect 93770 101386 94470 102086
rect 94679 101386 95379 102086
rect 95588 101386 96288 102086
rect 96497 101386 97197 102086
rect 97406 101386 98106 102086
rect 98315 101386 99015 102086
rect 99224 101386 99924 102086
rect 100133 101386 100833 102086
rect 101042 101386 101742 102086
rect 101951 101386 102651 102086
rect 102860 101386 103560 102086
rect 103769 101386 104469 102086
rect 104678 101386 105378 102086
rect 105587 101386 106287 102086
rect 106496 101386 107196 102086
rect 107405 101386 108105 102086
rect 108314 101386 109014 102086
rect 109223 101386 109923 102086
rect 110132 101386 110832 102086
rect 89225 100498 89925 101198
rect 90134 100498 90834 101198
rect 91043 100498 91743 101198
rect 91952 100498 92652 101198
rect 92861 100498 93561 101198
rect 93770 100498 94470 101198
rect 94679 100498 95379 101198
rect 95588 100498 96288 101198
rect 96497 100498 97197 101198
rect 97406 100498 98106 101198
rect 98315 100498 99015 101198
rect 99224 100498 99924 101198
rect 100133 100498 100833 101198
rect 101042 100498 101742 101198
rect 101951 100498 102651 101198
rect 102860 100498 103560 101198
rect 103769 100498 104469 101198
rect 104678 100498 105378 101198
rect 105587 100498 106287 101198
rect 106496 100498 107196 101198
rect 107405 100498 108105 101198
rect 108314 100498 109014 101198
rect 109223 100498 109923 101198
rect 110132 100498 110832 101198
rect 89225 99610 89925 100310
rect 90134 99610 90834 100310
rect 91043 99610 91743 100310
rect 91952 99610 92652 100310
rect 92861 99610 93561 100310
rect 93770 99610 94470 100310
rect 94679 99610 95379 100310
rect 95588 99610 96288 100310
rect 96497 99610 97197 100310
rect 97406 99610 98106 100310
rect 98315 99610 99015 100310
rect 99224 99610 99924 100310
rect 100133 99610 100833 100310
rect 101042 99610 101742 100310
rect 101951 99610 102651 100310
rect 102860 99610 103560 100310
rect 103769 99610 104469 100310
rect 104678 99610 105378 100310
rect 105587 99610 106287 100310
rect 106496 99610 107196 100310
rect 107405 99610 108105 100310
rect 108314 99610 109014 100310
rect 109223 99610 109923 100310
rect 110132 99610 110832 100310
rect 482072 102255 482772 102955
rect 483168 102255 483868 102955
rect 484264 102255 484964 102955
rect 485360 102255 486060 102955
rect 486456 102255 487156 102955
rect 487552 102255 488252 102955
rect 488648 102255 489348 102955
rect 489744 102255 490444 102955
rect 490840 102255 491540 102955
rect 491936 102255 492636 102955
rect 493032 102255 493732 102955
rect 494128 102255 494828 102955
rect 495224 102255 495924 102955
rect 496320 102255 497020 102955
rect 497416 102255 498116 102955
rect 498512 102255 499212 102955
rect 499608 102255 500308 102955
rect 500704 102255 501404 102955
rect 501800 102255 502500 102955
rect 502896 102255 503596 102955
rect 503992 102255 504692 102955
rect 505088 102255 505788 102955
rect 506184 102255 506884 102955
rect 507280 102255 507980 102955
rect 482072 101104 482772 101804
rect 483168 101104 483868 101804
rect 484264 101104 484964 101804
rect 485360 101104 486060 101804
rect 486456 101104 487156 101804
rect 487552 101104 488252 101804
rect 488648 101104 489348 101804
rect 489744 101104 490444 101804
rect 490840 101104 491540 101804
rect 491936 101104 492636 101804
rect 493032 101104 493732 101804
rect 494128 101104 494828 101804
rect 495224 101104 495924 101804
rect 496320 101104 497020 101804
rect 497416 101104 498116 101804
rect 498512 101104 499212 101804
rect 499608 101104 500308 101804
rect 500704 101104 501404 101804
rect 501800 101104 502500 101804
rect 502896 101104 503596 101804
rect 503992 101104 504692 101804
rect 505088 101104 505788 101804
rect 506184 101104 506884 101804
rect 507280 101104 507980 101804
rect 482072 99953 482772 100653
rect 483168 99953 483868 100653
rect 484264 99953 484964 100653
rect 485360 99953 486060 100653
rect 486456 99953 487156 100653
rect 487552 99953 488252 100653
rect 488648 99953 489348 100653
rect 489744 99953 490444 100653
rect 490840 99953 491540 100653
rect 491936 99953 492636 100653
rect 493032 99953 493732 100653
rect 494128 99953 494828 100653
rect 495224 99953 495924 100653
rect 496320 99953 497020 100653
rect 497416 99953 498116 100653
rect 498512 99953 499212 100653
rect 499608 99953 500308 100653
rect 500704 99953 501404 100653
rect 501800 99953 502500 100653
rect 502896 99953 503596 100653
rect 503992 99953 504692 100653
rect 505088 99953 505788 100653
rect 506184 99953 506884 100653
rect 507280 99953 507980 100653
rect 89225 98722 89925 99422
rect 90134 98722 90834 99422
rect 91043 98722 91743 99422
rect 91952 98722 92652 99422
rect 92861 98722 93561 99422
rect 93770 98722 94470 99422
rect 94679 98722 95379 99422
rect 95588 98722 96288 99422
rect 96497 98722 97197 99422
rect 97406 98722 98106 99422
rect 98315 98722 99015 99422
rect 99224 98722 99924 99422
rect 100133 98722 100833 99422
rect 101042 98722 101742 99422
rect 101951 98722 102651 99422
rect 102860 98722 103560 99422
rect 103769 98722 104469 99422
rect 104678 98722 105378 99422
rect 105587 98722 106287 99422
rect 106496 98722 107196 99422
rect 107405 98722 108105 99422
rect 108314 98722 109014 99422
rect 109223 98722 109923 99422
rect 110132 98722 110832 99422
<< metal4 >>
rect 87832 510796 112357 510951
rect 87832 510096 87948 510796
rect 88648 510096 88929 510796
rect 89629 510096 89910 510796
rect 90610 510096 90891 510796
rect 91591 510096 91872 510796
rect 92572 510096 92853 510796
rect 93553 510096 93834 510796
rect 94534 510096 94815 510796
rect 95515 510096 95796 510796
rect 96496 510096 96777 510796
rect 97477 510096 97758 510796
rect 98458 510096 98739 510796
rect 99439 510096 99720 510796
rect 100420 510096 100701 510796
rect 101401 510096 101682 510796
rect 102382 510096 102663 510796
rect 103363 510096 103644 510796
rect 104344 510096 104625 510796
rect 105325 510096 105606 510796
rect 106306 510096 106587 510796
rect 107287 510096 107568 510796
rect 108268 510096 108549 510796
rect 109249 510096 109530 510796
rect 110230 510096 110511 510796
rect 111211 510096 111492 510796
rect 112192 510096 112357 510796
rect 87832 509776 112357 510096
rect 87832 509076 87948 509776
rect 88648 509076 88929 509776
rect 89629 509076 89910 509776
rect 90610 509076 90891 509776
rect 91591 509076 91872 509776
rect 92572 509076 92853 509776
rect 93553 509076 93834 509776
rect 94534 509076 94815 509776
rect 95515 509076 95796 509776
rect 96496 509076 96777 509776
rect 97477 509076 97758 509776
rect 98458 509076 98739 509776
rect 99439 509076 99720 509776
rect 100420 509076 100701 509776
rect 101401 509076 101682 509776
rect 102382 509076 102663 509776
rect 103363 509076 103644 509776
rect 104344 509076 104625 509776
rect 105325 509076 105606 509776
rect 106306 509076 106587 509776
rect 107287 509076 107568 509776
rect 108268 509076 108549 509776
rect 109249 509076 109530 509776
rect 110230 509076 110511 509776
rect 111211 509076 111492 509776
rect 112192 509076 112357 509776
rect 87832 508756 112357 509076
rect 87832 508056 87948 508756
rect 88648 508056 88929 508756
rect 89629 508056 89910 508756
rect 90610 508056 90891 508756
rect 91591 508056 91872 508756
rect 92572 508056 92853 508756
rect 93553 508056 93834 508756
rect 94534 508056 94815 508756
rect 95515 508056 95796 508756
rect 96496 508056 96777 508756
rect 97477 508056 97758 508756
rect 98458 508056 98739 508756
rect 99439 508056 99720 508756
rect 100420 508056 100701 508756
rect 101401 508056 101682 508756
rect 102382 508056 102663 508756
rect 103363 508056 103644 508756
rect 104344 508056 104625 508756
rect 105325 508056 105606 508756
rect 106306 508056 106587 508756
rect 107287 508056 107568 508756
rect 108268 508056 108549 508756
rect 109249 508056 109530 508756
rect 110230 508056 110511 508756
rect 111211 508056 111492 508756
rect 112192 508056 112357 508756
rect 87832 507736 112357 508056
rect 87832 507715 87948 507736
rect 87777 507036 87948 507715
rect 88648 507036 88929 507736
rect 89629 507036 89910 507736
rect 90610 507036 90891 507736
rect 91591 507036 91872 507736
rect 92572 507036 92853 507736
rect 93553 507036 93834 507736
rect 94534 507036 94815 507736
rect 95515 507036 95796 507736
rect 96496 507036 96777 507736
rect 97477 507036 97758 507736
rect 98458 507036 98739 507736
rect 99439 507036 99720 507736
rect 100420 507036 100701 507736
rect 101401 507036 101682 507736
rect 102382 507036 102663 507736
rect 103363 507036 103644 507736
rect 104344 507036 104625 507736
rect 105325 507036 105606 507736
rect 106306 507036 106587 507736
rect 107287 507036 107568 507736
rect 108268 507036 108549 507736
rect 109249 507036 109530 507736
rect 110230 507036 110511 507736
rect 111211 507036 111492 507736
rect 112192 507036 112357 507736
rect 482253 508075 507466 508386
rect 482253 507551 482569 508075
rect 87777 506716 112357 507036
rect 87777 506016 87948 506716
rect 88648 506016 88929 506716
rect 89629 506016 89910 506716
rect 90610 506016 90891 506716
rect 91591 506016 91872 506716
rect 92572 506016 92853 506716
rect 93553 506016 93834 506716
rect 94534 506016 94815 506716
rect 95515 506016 95796 506716
rect 96496 506016 96777 506716
rect 97477 506016 97758 506716
rect 98458 506016 98739 506716
rect 99439 506016 99720 506716
rect 100420 506016 100701 506716
rect 101401 506016 101682 506716
rect 102382 506016 102663 506716
rect 103363 506016 103644 506716
rect 104344 506016 104625 506716
rect 105325 506016 105606 506716
rect 106306 506016 106587 506716
rect 107287 506016 107568 506716
rect 108268 506016 108549 506716
rect 109249 506016 109530 506716
rect 110230 506016 110511 506716
rect 111211 506016 111492 506716
rect 112192 506016 112357 506716
rect 87777 505696 112357 506016
rect 87777 504996 87948 505696
rect 88648 504996 88929 505696
rect 89629 504996 89910 505696
rect 90610 504996 90891 505696
rect 91591 504996 91872 505696
rect 92572 504996 92853 505696
rect 93553 504996 93834 505696
rect 94534 504996 94815 505696
rect 95515 504996 95796 505696
rect 96496 504996 96777 505696
rect 97477 504996 97758 505696
rect 98458 504996 98739 505696
rect 99439 504996 99720 505696
rect 100420 504996 100701 505696
rect 101401 504996 101682 505696
rect 102382 504996 102663 505696
rect 103363 504996 103644 505696
rect 104344 504996 104625 505696
rect 105325 504996 105606 505696
rect 106306 504996 106587 505696
rect 107287 504996 107568 505696
rect 108268 504996 108549 505696
rect 109249 504996 109530 505696
rect 110230 504996 110511 505696
rect 111211 504996 111492 505696
rect 112192 504996 112357 505696
rect 87777 504676 112357 504996
rect 87777 503976 87948 504676
rect 88648 503976 88929 504676
rect 89629 503976 89910 504676
rect 90610 503976 90891 504676
rect 91591 503976 91872 504676
rect 92572 503976 92853 504676
rect 93553 503976 93834 504676
rect 94534 503976 94815 504676
rect 95515 503976 95796 504676
rect 96496 503976 96777 504676
rect 97477 503976 97758 504676
rect 98458 503976 98739 504676
rect 99439 503976 99720 504676
rect 100420 503976 100701 504676
rect 101401 503976 101682 504676
rect 102382 503976 102663 504676
rect 103363 503976 103644 504676
rect 104344 503976 104625 504676
rect 105325 503976 105606 504676
rect 106306 503976 106587 504676
rect 107287 503976 107568 504676
rect 108268 503976 108549 504676
rect 109249 503976 109530 504676
rect 110230 503976 110511 504676
rect 111211 503976 111492 504676
rect 112192 503976 112357 504676
rect 87777 503656 112357 503976
rect 87777 502956 87948 503656
rect 88648 502956 88929 503656
rect 89629 502956 89910 503656
rect 90610 502956 90891 503656
rect 91591 502956 91872 503656
rect 92572 502956 92853 503656
rect 93553 502956 93834 503656
rect 94534 502956 94815 503656
rect 95515 502956 95796 503656
rect 96496 502956 96777 503656
rect 97477 502956 97758 503656
rect 98458 502956 98739 503656
rect 99439 502956 99720 503656
rect 100420 502956 100701 503656
rect 101401 502956 101682 503656
rect 102382 502956 102663 503656
rect 103363 502956 103644 503656
rect 104344 502956 104625 503656
rect 105325 502956 105606 503656
rect 106306 502956 106587 503656
rect 107287 502956 107568 503656
rect 108268 502956 108549 503656
rect 109249 502956 109530 503656
rect 110230 502956 110511 503656
rect 111211 502956 111492 503656
rect 112192 502956 112357 503656
rect 87777 502636 112357 502956
rect 87777 501936 87948 502636
rect 88648 501936 88929 502636
rect 89629 501936 89910 502636
rect 90610 501936 90891 502636
rect 91591 501936 91872 502636
rect 92572 501936 92853 502636
rect 93553 501936 93834 502636
rect 94534 501936 94815 502636
rect 95515 501936 95796 502636
rect 96496 501936 96777 502636
rect 97477 501936 97758 502636
rect 98458 501936 98739 502636
rect 99439 501936 99720 502636
rect 100420 501936 100701 502636
rect 101401 501936 101682 502636
rect 102382 501936 102663 502636
rect 103363 501936 103644 502636
rect 104344 501936 104625 502636
rect 105325 501936 105606 502636
rect 106306 501936 106587 502636
rect 107287 501936 107568 502636
rect 108268 501936 108549 502636
rect 109249 501936 109530 502636
rect 110230 501936 110511 502636
rect 111211 501936 111492 502636
rect 112192 501936 112357 502636
rect 87777 501616 112357 501936
rect 87777 500916 87948 501616
rect 88648 500916 88929 501616
rect 89629 500916 89910 501616
rect 90610 500916 90891 501616
rect 91591 500916 91872 501616
rect 92572 500916 92853 501616
rect 93553 500916 93834 501616
rect 94534 500916 94815 501616
rect 95515 500916 95796 501616
rect 96496 500916 96777 501616
rect 97477 500916 97758 501616
rect 98458 500916 98739 501616
rect 99439 500916 99720 501616
rect 100420 500916 100701 501616
rect 101401 500916 101682 501616
rect 102382 500916 102663 501616
rect 103363 500916 103644 501616
rect 104344 500916 104625 501616
rect 105325 500916 105606 501616
rect 106306 500916 106587 501616
rect 107287 500916 107568 501616
rect 108268 500916 108549 501616
rect 109249 500916 109530 501616
rect 110230 500916 110511 501616
rect 111211 500916 111492 501616
rect 112192 500916 112357 501616
rect 87777 500596 112357 500916
rect 87777 499896 87948 500596
rect 88648 499896 88929 500596
rect 89629 499896 89910 500596
rect 90610 499896 90891 500596
rect 91591 499896 91872 500596
rect 92572 499896 92853 500596
rect 93553 499896 93834 500596
rect 94534 499896 94815 500596
rect 95515 499896 95796 500596
rect 96496 499896 96777 500596
rect 97477 499896 97758 500596
rect 98458 499896 98739 500596
rect 99439 499896 99720 500596
rect 100420 499896 100701 500596
rect 101401 499896 101682 500596
rect 102382 499896 102663 500596
rect 103363 499896 103644 500596
rect 104344 499896 104625 500596
rect 105325 499896 105606 500596
rect 106306 499896 106587 500596
rect 107287 499896 107568 500596
rect 108268 499896 108549 500596
rect 109249 499896 109530 500596
rect 110230 499896 110511 500596
rect 111211 499896 111492 500596
rect 112192 499896 112357 500596
rect 87777 499576 112357 499896
rect 87777 498876 87948 499576
rect 88648 498876 88929 499576
rect 89629 498876 89910 499576
rect 90610 498876 90891 499576
rect 91591 498876 91872 499576
rect 92572 498876 92853 499576
rect 93553 498876 93834 499576
rect 94534 498876 94815 499576
rect 95515 498876 95796 499576
rect 96496 498876 96777 499576
rect 97477 498876 97758 499576
rect 98458 498876 98739 499576
rect 99439 498876 99720 499576
rect 100420 498876 100701 499576
rect 101401 498876 101682 499576
rect 102382 498876 102663 499576
rect 103363 498876 103644 499576
rect 104344 498876 104625 499576
rect 105325 498876 105606 499576
rect 106306 498876 106587 499576
rect 107287 498876 107568 499576
rect 108268 498876 108549 499576
rect 109249 498876 109530 499576
rect 110230 498876 110511 499576
rect 111211 498876 111492 499576
rect 112192 498876 112357 499576
rect 87777 498556 112357 498876
rect 87777 497856 87948 498556
rect 88648 497856 88929 498556
rect 89629 497856 89910 498556
rect 90610 497856 90891 498556
rect 91591 497856 91872 498556
rect 92572 497856 92853 498556
rect 93553 497856 93834 498556
rect 94534 497856 94815 498556
rect 95515 497856 95796 498556
rect 96496 497856 96777 498556
rect 97477 497856 97758 498556
rect 98458 497856 98739 498556
rect 99439 497856 99720 498556
rect 100420 497856 100701 498556
rect 101401 497856 101682 498556
rect 102382 497856 102663 498556
rect 103363 497856 103644 498556
rect 104344 497856 104625 498556
rect 105325 497856 105606 498556
rect 106306 497856 106587 498556
rect 107287 497856 107568 498556
rect 108268 497856 108549 498556
rect 109249 497856 109530 498556
rect 110230 497856 110511 498556
rect 111211 497856 111492 498556
rect 112192 497856 112357 498556
rect 87777 497536 112357 497856
rect 87777 496836 87948 497536
rect 88648 496836 88929 497536
rect 89629 496836 89910 497536
rect 90610 496836 90891 497536
rect 91591 496836 91872 497536
rect 92572 496836 92853 497536
rect 93553 496836 93834 497536
rect 94534 496836 94815 497536
rect 95515 496836 95796 497536
rect 96496 496836 96777 497536
rect 97477 496836 97758 497536
rect 98458 496836 98739 497536
rect 99439 496836 99720 497536
rect 100420 496836 100701 497536
rect 101401 496836 101682 497536
rect 102382 496836 102663 497536
rect 103363 496836 103644 497536
rect 104344 496836 104625 497536
rect 105325 496836 105606 497536
rect 106306 496836 106587 497536
rect 107287 496836 107568 497536
rect 108268 496836 108549 497536
rect 109249 496836 109530 497536
rect 110230 496836 110511 497536
rect 111211 496836 111492 497536
rect 112192 496836 112357 497536
rect 87777 496516 112357 496836
rect 87777 495816 87948 496516
rect 88648 495816 88929 496516
rect 89629 495816 89910 496516
rect 90610 495816 90891 496516
rect 91591 495816 91872 496516
rect 92572 495816 92853 496516
rect 93553 495816 93834 496516
rect 94534 495816 94815 496516
rect 95515 495816 95796 496516
rect 96496 495816 96777 496516
rect 97477 495816 97758 496516
rect 98458 495816 98739 496516
rect 99439 495816 99720 496516
rect 100420 495816 100701 496516
rect 101401 495816 101682 496516
rect 102382 495816 102663 496516
rect 103363 495816 103644 496516
rect 104344 495816 104625 496516
rect 105325 495816 105606 496516
rect 106306 495816 106587 496516
rect 107287 495816 107568 496516
rect 108268 495816 108549 496516
rect 109249 495816 109530 496516
rect 110230 495816 110511 496516
rect 111211 495816 111492 496516
rect 112192 495816 112357 496516
rect 87777 495496 112357 495816
rect 87777 494796 87948 495496
rect 88648 494796 88929 495496
rect 89629 494796 89910 495496
rect 90610 494796 90891 495496
rect 91591 494796 91872 495496
rect 92572 494796 92853 495496
rect 93553 494796 93834 495496
rect 94534 494796 94815 495496
rect 95515 494796 95796 495496
rect 96496 494796 96777 495496
rect 97477 494796 97758 495496
rect 98458 494796 98739 495496
rect 99439 494796 99720 495496
rect 100420 494796 100701 495496
rect 101401 494796 101682 495496
rect 102382 494796 102663 495496
rect 103363 494796 103644 495496
rect 104344 494796 104625 495496
rect 105325 494796 105606 495496
rect 106306 494796 106587 495496
rect 107287 494796 107568 495496
rect 108268 494796 108549 495496
rect 109249 494796 109530 495496
rect 110230 494796 110511 495496
rect 111211 494796 111492 495496
rect 112192 494796 112357 495496
rect 87777 494476 112357 494796
rect 87777 493776 87948 494476
rect 88648 493776 88929 494476
rect 89629 493776 89910 494476
rect 90610 493776 90891 494476
rect 91591 493776 91872 494476
rect 92572 493776 92853 494476
rect 93553 493776 93834 494476
rect 94534 493776 94815 494476
rect 95515 493776 95796 494476
rect 96496 493776 96777 494476
rect 97477 493776 97758 494476
rect 98458 493776 98739 494476
rect 99439 493776 99720 494476
rect 100420 493776 100701 494476
rect 101401 493776 101682 494476
rect 102382 493776 102663 494476
rect 103363 493776 103644 494476
rect 104344 493776 104625 494476
rect 105325 493776 105606 494476
rect 106306 493776 106587 494476
rect 107287 493776 107568 494476
rect 108268 493776 108549 494476
rect 109249 493776 109530 494476
rect 110230 493776 110511 494476
rect 111211 493776 111492 494476
rect 112192 493776 112357 494476
rect 87777 493456 112357 493776
rect 87777 492756 87948 493456
rect 88648 492756 88929 493456
rect 89629 492756 89910 493456
rect 90610 492756 90891 493456
rect 91591 492756 91872 493456
rect 92572 492756 92853 493456
rect 93553 492756 93834 493456
rect 94534 492756 94815 493456
rect 95515 492756 95796 493456
rect 96496 492756 96777 493456
rect 97477 492756 97758 493456
rect 98458 492756 98739 493456
rect 99439 492756 99720 493456
rect 100420 492756 100701 493456
rect 101401 492756 101682 493456
rect 102382 492756 102663 493456
rect 103363 492756 103644 493456
rect 104344 492756 104625 493456
rect 105325 492756 105606 493456
rect 106306 492756 106587 493456
rect 107287 492756 107568 493456
rect 108268 492756 108549 493456
rect 109249 492756 109530 493456
rect 110230 492756 110511 493456
rect 111211 492756 111492 493456
rect 112192 492756 112357 493456
rect 87777 492436 112357 492756
rect 87777 491736 87948 492436
rect 88648 491736 88929 492436
rect 89629 491736 89910 492436
rect 90610 491736 90891 492436
rect 91591 491736 91872 492436
rect 92572 491736 92853 492436
rect 93553 491736 93834 492436
rect 94534 491736 94815 492436
rect 95515 491736 95796 492436
rect 96496 491736 96777 492436
rect 97477 491736 97758 492436
rect 98458 491736 98739 492436
rect 99439 491736 99720 492436
rect 100420 491736 100701 492436
rect 101401 491736 101682 492436
rect 102382 491736 102663 492436
rect 103363 491736 103644 492436
rect 104344 491736 104625 492436
rect 105325 491736 105606 492436
rect 106306 491736 106587 492436
rect 107287 491736 107568 492436
rect 108268 491736 108549 492436
rect 109249 491736 109530 492436
rect 110230 491736 110511 492436
rect 111211 491736 111492 492436
rect 112192 491736 112357 492436
rect 87777 491416 112357 491736
rect 87777 490716 87948 491416
rect 88648 490716 88929 491416
rect 89629 490716 89910 491416
rect 90610 490716 90891 491416
rect 91591 490716 91872 491416
rect 92572 490716 92853 491416
rect 93553 490716 93834 491416
rect 94534 490716 94815 491416
rect 95515 490716 95796 491416
rect 96496 490716 96777 491416
rect 97477 490716 97758 491416
rect 98458 490716 98739 491416
rect 99439 490716 99720 491416
rect 100420 490716 100701 491416
rect 101401 490716 101682 491416
rect 102382 490716 102663 491416
rect 103363 490716 103644 491416
rect 104344 490716 104625 491416
rect 105325 490716 105606 491416
rect 106306 490716 106587 491416
rect 107287 490716 107568 491416
rect 108268 490716 108549 491416
rect 109249 490716 109530 491416
rect 110230 490716 110511 491416
rect 111211 490716 111492 491416
rect 112192 490716 112357 491416
rect 87777 490396 112357 490716
rect 87777 489696 87948 490396
rect 88648 489696 88929 490396
rect 89629 489696 89910 490396
rect 90610 489696 90891 490396
rect 91591 489696 91872 490396
rect 92572 489696 92853 490396
rect 93553 489696 93834 490396
rect 94534 489696 94815 490396
rect 95515 489696 95796 490396
rect 96496 489696 96777 490396
rect 97477 489696 97758 490396
rect 98458 489696 98739 490396
rect 99439 489696 99720 490396
rect 100420 489696 100701 490396
rect 101401 489696 101682 490396
rect 102382 489696 102663 490396
rect 103363 489696 103644 490396
rect 104344 489696 104625 490396
rect 105325 489696 105606 490396
rect 106306 489696 106587 490396
rect 107287 489696 107568 490396
rect 108268 489696 108549 490396
rect 109249 489696 109530 490396
rect 110230 489696 110511 490396
rect 111211 489696 111492 490396
rect 112192 489696 112357 490396
rect 87777 489376 112357 489696
rect 87777 488676 87948 489376
rect 88648 488676 88929 489376
rect 89629 488676 89910 489376
rect 90610 488676 90891 489376
rect 91591 488676 91872 489376
rect 92572 488676 92853 489376
rect 93553 488676 93834 489376
rect 94534 488676 94815 489376
rect 95515 488676 95796 489376
rect 96496 488676 96777 489376
rect 97477 488676 97758 489376
rect 98458 488676 98739 489376
rect 99439 488676 99720 489376
rect 100420 488676 100701 489376
rect 101401 488676 101682 489376
rect 102382 488676 102663 489376
rect 103363 488676 103644 489376
rect 104344 488676 104625 489376
rect 105325 488676 105606 489376
rect 106306 488676 106587 489376
rect 107287 488676 107568 489376
rect 108268 488676 108549 489376
rect 109249 488676 109530 489376
rect 110230 488676 110511 489376
rect 111211 488676 111492 489376
rect 112192 488676 112357 489376
rect 87777 488356 112357 488676
rect 87777 487656 87948 488356
rect 88648 487656 88929 488356
rect 89629 487656 89910 488356
rect 90610 487656 90891 488356
rect 91591 487656 91872 488356
rect 92572 487656 92853 488356
rect 93553 487656 93834 488356
rect 94534 487656 94815 488356
rect 95515 487656 95796 488356
rect 96496 487656 96777 488356
rect 97477 487656 97758 488356
rect 98458 487656 98739 488356
rect 99439 487656 99720 488356
rect 100420 487656 100701 488356
rect 101401 487656 101682 488356
rect 102382 487656 102663 488356
rect 103363 487656 103644 488356
rect 104344 487656 104625 488356
rect 105325 487656 105606 488356
rect 106306 487656 106587 488356
rect 107287 487656 107568 488356
rect 108268 487656 108549 488356
rect 109249 487656 109530 488356
rect 110230 487656 110511 488356
rect 111211 487656 111492 488356
rect 112192 487656 112357 488356
rect 87777 487336 112357 487656
rect 87777 486636 87948 487336
rect 88648 486636 88929 487336
rect 89629 486636 89910 487336
rect 90610 486636 90891 487336
rect 91591 486636 91872 487336
rect 92572 486636 92853 487336
rect 93553 486636 93834 487336
rect 94534 486636 94815 487336
rect 95515 486636 95796 487336
rect 96496 486636 96777 487336
rect 97477 486636 97758 487336
rect 98458 486636 98739 487336
rect 99439 486636 99720 487336
rect 100420 486636 100701 487336
rect 101401 486636 101682 487336
rect 102382 486636 102663 487336
rect 103363 486636 103644 487336
rect 104344 486636 104625 487336
rect 105325 486636 105606 487336
rect 106306 486636 106587 487336
rect 107287 486636 107568 487336
rect 108268 486636 108549 487336
rect 109249 486636 109530 487336
rect 110230 486636 110511 487336
rect 111211 486636 111492 487336
rect 112192 486636 112357 487336
rect 87777 486316 112357 486636
rect 87777 485616 87948 486316
rect 88648 485616 88929 486316
rect 89629 485616 89910 486316
rect 90610 485616 90891 486316
rect 91591 485616 91872 486316
rect 92572 485616 92853 486316
rect 93553 485616 93834 486316
rect 94534 485616 94815 486316
rect 95515 485616 95796 486316
rect 96496 485616 96777 486316
rect 97477 485616 97758 486316
rect 98458 485616 98739 486316
rect 99439 485616 99720 486316
rect 100420 485616 100701 486316
rect 101401 485616 101682 486316
rect 102382 485616 102663 486316
rect 103363 485616 103644 486316
rect 104344 485616 104625 486316
rect 105325 485616 105606 486316
rect 106306 485616 106587 486316
rect 107287 485616 107568 486316
rect 108268 485616 108549 486316
rect 109249 485616 109530 486316
rect 110230 485616 110511 486316
rect 111211 485616 111492 486316
rect 112192 485616 112357 486316
rect 87777 485451 112357 485616
rect 481938 507375 482569 507551
rect 483269 507375 483896 508075
rect 484596 507375 485223 508075
rect 485923 507375 486550 508075
rect 487250 507375 487877 508075
rect 488577 507375 489204 508075
rect 489904 507375 490531 508075
rect 491231 507375 491858 508075
rect 492558 507375 493185 508075
rect 493885 507375 494512 508075
rect 495212 507375 495839 508075
rect 496539 507375 497166 508075
rect 497866 507375 498493 508075
rect 499193 507375 499820 508075
rect 500520 507375 501147 508075
rect 501847 507375 502474 508075
rect 503174 507375 503801 508075
rect 504501 507375 505128 508075
rect 505828 507375 506455 508075
rect 507155 507375 507466 508075
rect 481938 506748 507466 507375
rect 481938 506048 482569 506748
rect 483269 506048 483896 506748
rect 484596 506048 485223 506748
rect 485923 506048 486550 506748
rect 487250 506048 487877 506748
rect 488577 506048 489204 506748
rect 489904 506048 490531 506748
rect 491231 506048 491858 506748
rect 492558 506048 493185 506748
rect 493885 506048 494512 506748
rect 495212 506048 495839 506748
rect 496539 506048 497166 506748
rect 497866 506048 498493 506748
rect 499193 506048 499820 506748
rect 500520 506048 501147 506748
rect 501847 506048 502474 506748
rect 503174 506048 503801 506748
rect 504501 506048 505128 506748
rect 505828 506048 506455 506748
rect 507155 506048 507466 506748
rect 481938 505421 507466 506048
rect 481938 504721 482569 505421
rect 483269 504721 483896 505421
rect 484596 504721 485223 505421
rect 485923 504721 486550 505421
rect 487250 504721 487877 505421
rect 488577 504721 489204 505421
rect 489904 504721 490531 505421
rect 491231 504721 491858 505421
rect 492558 504721 493185 505421
rect 493885 504721 494512 505421
rect 495212 504721 495839 505421
rect 496539 504721 497166 505421
rect 497866 504721 498493 505421
rect 499193 504721 499820 505421
rect 500520 504721 501147 505421
rect 501847 504721 502474 505421
rect 503174 504721 503801 505421
rect 504501 504721 505128 505421
rect 505828 504721 506455 505421
rect 507155 504721 507466 505421
rect 481938 504094 507466 504721
rect 481938 503394 482569 504094
rect 483269 503394 483896 504094
rect 484596 503394 485223 504094
rect 485923 503394 486550 504094
rect 487250 503394 487877 504094
rect 488577 503394 489204 504094
rect 489904 503394 490531 504094
rect 491231 503394 491858 504094
rect 492558 503394 493185 504094
rect 493885 503394 494512 504094
rect 495212 503394 495839 504094
rect 496539 503394 497166 504094
rect 497866 503394 498493 504094
rect 499193 503394 499820 504094
rect 500520 503394 501147 504094
rect 501847 503394 502474 504094
rect 503174 503394 503801 504094
rect 504501 503394 505128 504094
rect 505828 503394 506455 504094
rect 507155 503394 507466 504094
rect 481938 502767 507466 503394
rect 481938 502067 482569 502767
rect 483269 502067 483896 502767
rect 484596 502067 485223 502767
rect 485923 502067 486550 502767
rect 487250 502067 487877 502767
rect 488577 502067 489204 502767
rect 489904 502067 490531 502767
rect 491231 502067 491858 502767
rect 492558 502067 493185 502767
rect 493885 502067 494512 502767
rect 495212 502067 495839 502767
rect 496539 502067 497166 502767
rect 497866 502067 498493 502767
rect 499193 502067 499820 502767
rect 500520 502067 501147 502767
rect 501847 502067 502474 502767
rect 503174 502067 503801 502767
rect 504501 502067 505128 502767
rect 505828 502067 506455 502767
rect 507155 502067 507466 502767
rect 481938 501440 507466 502067
rect 481938 500740 482569 501440
rect 483269 500740 483896 501440
rect 484596 500740 485223 501440
rect 485923 500740 486550 501440
rect 487250 500740 487877 501440
rect 488577 500740 489204 501440
rect 489904 500740 490531 501440
rect 491231 500740 491858 501440
rect 492558 500740 493185 501440
rect 493885 500740 494512 501440
rect 495212 500740 495839 501440
rect 496539 500740 497166 501440
rect 497866 500740 498493 501440
rect 499193 500740 499820 501440
rect 500520 500740 501147 501440
rect 501847 500740 502474 501440
rect 503174 500740 503801 501440
rect 504501 500740 505128 501440
rect 505828 500740 506455 501440
rect 507155 500740 507466 501440
rect 481938 500113 507466 500740
rect 481938 499413 482569 500113
rect 483269 499413 483896 500113
rect 484596 499413 485223 500113
rect 485923 499413 486550 500113
rect 487250 499413 487877 500113
rect 488577 499413 489204 500113
rect 489904 499413 490531 500113
rect 491231 499413 491858 500113
rect 492558 499413 493185 500113
rect 493885 499413 494512 500113
rect 495212 499413 495839 500113
rect 496539 499413 497166 500113
rect 497866 499413 498493 500113
rect 499193 499413 499820 500113
rect 500520 499413 501147 500113
rect 501847 499413 502474 500113
rect 503174 499413 503801 500113
rect 504501 499413 505128 500113
rect 505828 499413 506455 500113
rect 507155 499413 507466 500113
rect 481938 498786 507466 499413
rect 481938 498086 482569 498786
rect 483269 498086 483896 498786
rect 484596 498086 485223 498786
rect 485923 498086 486550 498786
rect 487250 498086 487877 498786
rect 488577 498086 489204 498786
rect 489904 498086 490531 498786
rect 491231 498086 491858 498786
rect 492558 498086 493185 498786
rect 493885 498086 494512 498786
rect 495212 498086 495839 498786
rect 496539 498086 497166 498786
rect 497866 498086 498493 498786
rect 499193 498086 499820 498786
rect 500520 498086 501147 498786
rect 501847 498086 502474 498786
rect 503174 498086 503801 498786
rect 504501 498086 505128 498786
rect 505828 498086 506455 498786
rect 507155 498086 507466 498786
rect 481938 497459 507466 498086
rect 481938 496759 482569 497459
rect 483269 496759 483896 497459
rect 484596 496759 485223 497459
rect 485923 496759 486550 497459
rect 487250 496759 487877 497459
rect 488577 496759 489204 497459
rect 489904 496759 490531 497459
rect 491231 496759 491858 497459
rect 492558 496759 493185 497459
rect 493885 496759 494512 497459
rect 495212 496759 495839 497459
rect 496539 496759 497166 497459
rect 497866 496759 498493 497459
rect 499193 496759 499820 497459
rect 500520 496759 501147 497459
rect 501847 496759 502474 497459
rect 503174 496759 503801 497459
rect 504501 496759 505128 497459
rect 505828 496759 506455 497459
rect 507155 496759 507466 497459
rect 481938 496132 507466 496759
rect 481938 495432 482569 496132
rect 483269 495432 483896 496132
rect 484596 495432 485223 496132
rect 485923 495432 486550 496132
rect 487250 495432 487877 496132
rect 488577 495432 489204 496132
rect 489904 495432 490531 496132
rect 491231 495432 491858 496132
rect 492558 495432 493185 496132
rect 493885 495432 494512 496132
rect 495212 495432 495839 496132
rect 496539 495432 497166 496132
rect 497866 495432 498493 496132
rect 499193 495432 499820 496132
rect 500520 495432 501147 496132
rect 501847 495432 502474 496132
rect 503174 495432 503801 496132
rect 504501 495432 505128 496132
rect 505828 495432 506455 496132
rect 507155 495432 507466 496132
rect 481938 494805 507466 495432
rect 481938 494105 482569 494805
rect 483269 494105 483896 494805
rect 484596 494105 485223 494805
rect 485923 494105 486550 494805
rect 487250 494105 487877 494805
rect 488577 494105 489204 494805
rect 489904 494105 490531 494805
rect 491231 494105 491858 494805
rect 492558 494105 493185 494805
rect 493885 494105 494512 494805
rect 495212 494105 495839 494805
rect 496539 494105 497166 494805
rect 497866 494105 498493 494805
rect 499193 494105 499820 494805
rect 500520 494105 501147 494805
rect 501847 494105 502474 494805
rect 503174 494105 503801 494805
rect 504501 494105 505128 494805
rect 505828 494105 506455 494805
rect 507155 494105 507466 494805
rect 481938 493478 507466 494105
rect 481938 492778 482569 493478
rect 483269 492778 483896 493478
rect 484596 492778 485223 493478
rect 485923 492778 486550 493478
rect 487250 492778 487877 493478
rect 488577 492778 489204 493478
rect 489904 492778 490531 493478
rect 491231 492778 491858 493478
rect 492558 492778 493185 493478
rect 493885 492778 494512 493478
rect 495212 492778 495839 493478
rect 496539 492778 497166 493478
rect 497866 492778 498493 493478
rect 499193 492778 499820 493478
rect 500520 492778 501147 493478
rect 501847 492778 502474 493478
rect 503174 492778 503801 493478
rect 504501 492778 505128 493478
rect 505828 492778 506455 493478
rect 507155 492778 507466 493478
rect 481938 492151 507466 492778
rect 481938 491451 482569 492151
rect 483269 491451 483896 492151
rect 484596 491451 485223 492151
rect 485923 491451 486550 492151
rect 487250 491451 487877 492151
rect 488577 491451 489204 492151
rect 489904 491451 490531 492151
rect 491231 491451 491858 492151
rect 492558 491451 493185 492151
rect 493885 491451 494512 492151
rect 495212 491451 495839 492151
rect 496539 491451 497166 492151
rect 497866 491451 498493 492151
rect 499193 491451 499820 492151
rect 500520 491451 501147 492151
rect 501847 491451 502474 492151
rect 503174 491451 503801 492151
rect 504501 491451 505128 492151
rect 505828 491451 506455 492151
rect 507155 491451 507466 492151
rect 481938 490824 507466 491451
rect 481938 490124 482569 490824
rect 483269 490124 483896 490824
rect 484596 490124 485223 490824
rect 485923 490124 486550 490824
rect 487250 490124 487877 490824
rect 488577 490124 489204 490824
rect 489904 490124 490531 490824
rect 491231 490124 491858 490824
rect 492558 490124 493185 490824
rect 493885 490124 494512 490824
rect 495212 490124 495839 490824
rect 496539 490124 497166 490824
rect 497866 490124 498493 490824
rect 499193 490124 499820 490824
rect 500520 490124 501147 490824
rect 501847 490124 502474 490824
rect 503174 490124 503801 490824
rect 504501 490124 505128 490824
rect 505828 490124 506455 490824
rect 507155 490124 507466 490824
rect 481938 489497 507466 490124
rect 481938 488797 482569 489497
rect 483269 488797 483896 489497
rect 484596 488797 485223 489497
rect 485923 488797 486550 489497
rect 487250 488797 487877 489497
rect 488577 488797 489204 489497
rect 489904 488797 490531 489497
rect 491231 488797 491858 489497
rect 492558 488797 493185 489497
rect 493885 488797 494512 489497
rect 495212 488797 495839 489497
rect 496539 488797 497166 489497
rect 497866 488797 498493 489497
rect 499193 488797 499820 489497
rect 500520 488797 501147 489497
rect 501847 488797 502474 489497
rect 503174 488797 503801 489497
rect 504501 488797 505128 489497
rect 505828 488797 506455 489497
rect 507155 488797 507466 489497
rect 481938 488170 507466 488797
rect 481938 487470 482569 488170
rect 483269 487470 483896 488170
rect 484596 487470 485223 488170
rect 485923 487470 486550 488170
rect 487250 487470 487877 488170
rect 488577 487470 489204 488170
rect 489904 487470 490531 488170
rect 491231 487470 491858 488170
rect 492558 487470 493185 488170
rect 493885 487470 494512 488170
rect 495212 487470 495839 488170
rect 496539 487470 497166 488170
rect 497866 487470 498493 488170
rect 499193 487470 499820 488170
rect 500520 487470 501147 488170
rect 501847 487470 502474 488170
rect 503174 487470 503801 488170
rect 504501 487470 505128 488170
rect 505828 487470 506455 488170
rect 507155 487470 507466 488170
rect 481938 486843 507466 487470
rect 481938 486143 482569 486843
rect 483269 486143 483896 486843
rect 484596 486143 485223 486843
rect 485923 486143 486550 486843
rect 487250 486143 487877 486843
rect 488577 486143 489204 486843
rect 489904 486143 490531 486843
rect 491231 486143 491858 486843
rect 492558 486143 493185 486843
rect 493885 486143 494512 486843
rect 495212 486143 495839 486843
rect 496539 486143 497166 486843
rect 497866 486143 498493 486843
rect 499193 486143 499820 486843
rect 500520 486143 501147 486843
rect 501847 486143 502474 486843
rect 503174 486143 503801 486843
rect 504501 486143 505128 486843
rect 505828 486143 506455 486843
rect 507155 486143 507466 486843
rect 481938 485516 507466 486143
rect 87777 485163 110934 485451
rect 91770 468097 108327 485163
rect 481938 484816 482569 485516
rect 483269 484816 483896 485516
rect 484596 484816 485223 485516
rect 485923 484816 486550 485516
rect 487250 484816 487877 485516
rect 488577 484816 489204 485516
rect 489904 484816 490531 485516
rect 491231 484816 491858 485516
rect 492558 484816 493185 485516
rect 493885 484816 494512 485516
rect 495212 484816 495839 485516
rect 496539 484816 497166 485516
rect 497866 484816 498493 485516
rect 499193 484816 499820 485516
rect 500520 484816 501147 485516
rect 501847 484816 502474 485516
rect 503174 484816 503801 485516
rect 504501 484816 505128 485516
rect 505828 484816 506455 485516
rect 507155 484816 507466 485516
rect 481938 484189 507466 484816
rect 481938 483489 482569 484189
rect 483269 483489 483896 484189
rect 484596 483489 485223 484189
rect 485923 483489 486550 484189
rect 487250 483489 487877 484189
rect 488577 483489 489204 484189
rect 489904 483489 490531 484189
rect 491231 483489 491858 484189
rect 492558 483489 493185 484189
rect 493885 483489 494512 484189
rect 495212 483489 495839 484189
rect 496539 483489 497166 484189
rect 497866 483489 498493 484189
rect 499193 483489 499820 484189
rect 500520 483489 501147 484189
rect 501847 483489 502474 484189
rect 503174 483489 503801 484189
rect 504501 483489 505128 484189
rect 505828 483489 506455 484189
rect 507155 483489 507466 484189
rect 481938 483173 507466 483489
rect 481938 482808 506681 483173
rect 444162 480913 468473 481095
rect 444162 480840 444322 480913
rect 90963 467581 108327 468097
rect 90963 467431 91879 467581
rect 92029 467431 92147 467581
rect 92297 467431 92415 467581
rect 92565 467431 92683 467581
rect 92833 467431 92951 467581
rect 93101 467431 93219 467581
rect 93369 467431 93487 467581
rect 93637 467431 93755 467581
rect 93905 467431 94023 467581
rect 94173 467431 94291 467581
rect 94441 467431 108327 467581
rect 90963 467343 108327 467431
rect 90963 467193 91879 467343
rect 92029 467193 92147 467343
rect 92297 467193 92415 467343
rect 92565 467193 92683 467343
rect 92833 467193 92951 467343
rect 93101 467193 93219 467343
rect 93369 467193 93487 467343
rect 93637 467193 93755 467343
rect 93905 467193 94023 467343
rect 94173 467193 94291 467343
rect 94441 467193 108327 467343
rect 90963 467105 108327 467193
rect 90963 466955 91879 467105
rect 92029 466955 92147 467105
rect 92297 466955 92415 467105
rect 92565 466955 92683 467105
rect 92833 466955 92951 467105
rect 93101 466955 93219 467105
rect 93369 466955 93487 467105
rect 93637 466955 93755 467105
rect 93905 466955 94023 467105
rect 94173 466955 94291 467105
rect 94441 466955 108327 467105
rect 90963 466867 108327 466955
rect 90963 466717 91879 466867
rect 92029 466717 92147 466867
rect 92297 466717 92415 466867
rect 92565 466717 92683 466867
rect 92833 466717 92951 466867
rect 93101 466717 93219 466867
rect 93369 466717 93487 466867
rect 93637 466717 93755 466867
rect 93905 466717 94023 466867
rect 94173 466717 94291 466867
rect 94441 466717 108327 466867
rect 90963 466629 108327 466717
rect 90963 466479 91879 466629
rect 92029 466479 92147 466629
rect 92297 466479 92415 466629
rect 92565 466479 92683 466629
rect 92833 466479 92951 466629
rect 93101 466479 93219 466629
rect 93369 466479 93487 466629
rect 93637 466479 93755 466629
rect 93905 466479 94023 466629
rect 94173 466479 94291 466629
rect 94441 466479 108327 466629
rect 90963 466391 108327 466479
rect 90963 466241 91879 466391
rect 92029 466241 92147 466391
rect 92297 466241 92415 466391
rect 92565 466241 92683 466391
rect 92833 466241 92951 466391
rect 93101 466241 93219 466391
rect 93369 466241 93487 466391
rect 93637 466241 93755 466391
rect 93905 466241 94023 466391
rect 94173 466241 94291 466391
rect 94441 466241 108327 466391
rect 90963 466153 108327 466241
rect 90963 466003 91879 466153
rect 92029 466003 92147 466153
rect 92297 466003 92415 466153
rect 92565 466003 92683 466153
rect 92833 466003 92951 466153
rect 93101 466003 93219 466153
rect 93369 466003 93487 466153
rect 93637 466003 93755 466153
rect 93905 466003 94023 466153
rect 94173 466003 94291 466153
rect 94441 466003 108327 466153
rect 90963 465915 108327 466003
rect 90963 465765 91879 465915
rect 92029 465765 92147 465915
rect 92297 465765 92415 465915
rect 92565 465765 92683 465915
rect 92833 465765 92951 465915
rect 93101 465765 93219 465915
rect 93369 465765 93487 465915
rect 93637 465765 93755 465915
rect 93905 465765 94023 465915
rect 94173 465765 94291 465915
rect 94441 465765 108327 465915
rect 90963 465677 108327 465765
rect 90963 465527 91879 465677
rect 92029 465527 92147 465677
rect 92297 465527 92415 465677
rect 92565 465527 92683 465677
rect 92833 465527 92951 465677
rect 93101 465527 93219 465677
rect 93369 465527 93487 465677
rect 93637 465527 93755 465677
rect 93905 465527 94023 465677
rect 94173 465527 94291 465677
rect 94441 465527 108327 465677
rect 90963 465439 108327 465527
rect 90963 465289 91879 465439
rect 92029 465289 92147 465439
rect 92297 465289 92415 465439
rect 92565 465289 92683 465439
rect 92833 465289 92951 465439
rect 93101 465289 93219 465439
rect 93369 465289 93487 465439
rect 93637 465289 93755 465439
rect 93905 465289 94023 465439
rect 94173 465289 94291 465439
rect 94441 465289 108327 465439
rect 90963 464614 108327 465289
rect 91770 120594 108327 464614
rect 118930 480296 144555 480560
rect 118930 479596 119166 480296
rect 119866 479596 120188 480296
rect 120888 479596 121210 480296
rect 121910 479596 122232 480296
rect 122932 479596 123254 480296
rect 123954 479596 124276 480296
rect 124976 479596 125298 480296
rect 125998 479596 126320 480296
rect 127020 479596 127342 480296
rect 128042 479596 128364 480296
rect 129064 479596 129386 480296
rect 130086 479596 130408 480296
rect 131108 479596 131430 480296
rect 132130 479596 132452 480296
rect 133152 479596 133474 480296
rect 134174 479596 134496 480296
rect 135196 479596 135518 480296
rect 136218 479596 136540 480296
rect 137240 479596 137562 480296
rect 138262 479596 138584 480296
rect 139284 479596 139606 480296
rect 140306 479596 140628 480296
rect 141328 479596 141650 480296
rect 142350 479596 142672 480296
rect 143372 479596 143694 480296
rect 144394 479596 144555 480296
rect 118930 479224 144555 479596
rect 118930 478524 119166 479224
rect 119866 478524 120188 479224
rect 120888 478524 121210 479224
rect 121910 478524 122232 479224
rect 122932 478524 123254 479224
rect 123954 478524 124276 479224
rect 124976 478524 125298 479224
rect 125998 478524 126320 479224
rect 127020 478524 127342 479224
rect 128042 478524 128364 479224
rect 129064 478524 129386 479224
rect 130086 478524 130408 479224
rect 131108 478524 131430 479224
rect 132130 478524 132452 479224
rect 133152 478524 133474 479224
rect 134174 478524 134496 479224
rect 135196 478524 135518 479224
rect 136218 478524 136540 479224
rect 137240 478524 137562 479224
rect 138262 478524 138584 479224
rect 139284 478524 139606 479224
rect 140306 478524 140628 479224
rect 141328 478524 141650 479224
rect 142350 478524 142672 479224
rect 143372 478524 143694 479224
rect 144394 478524 144555 479224
rect 118930 478152 144555 478524
rect 118930 477452 119166 478152
rect 119866 477452 120188 478152
rect 120888 477452 121210 478152
rect 121910 477452 122232 478152
rect 122932 477452 123254 478152
rect 123954 477452 124276 478152
rect 124976 477452 125298 478152
rect 125998 477452 126320 478152
rect 127020 477452 127342 478152
rect 128042 477452 128364 478152
rect 129064 477452 129386 478152
rect 130086 477452 130408 478152
rect 131108 477452 131430 478152
rect 132130 477452 132452 478152
rect 133152 477452 133474 478152
rect 134174 477452 134496 478152
rect 135196 477452 135518 478152
rect 136218 477452 136540 478152
rect 137240 477452 137562 478152
rect 138262 477452 138584 478152
rect 139284 477452 139606 478152
rect 140306 477452 140628 478152
rect 141328 477452 141650 478152
rect 142350 477452 142672 478152
rect 143372 477452 143694 478152
rect 144394 477452 144555 478152
rect 118930 477080 144555 477452
rect 118930 476380 119166 477080
rect 119866 476380 120188 477080
rect 120888 476380 121210 477080
rect 121910 476380 122232 477080
rect 122932 476380 123254 477080
rect 123954 476380 124276 477080
rect 124976 476380 125298 477080
rect 125998 476380 126320 477080
rect 127020 476380 127342 477080
rect 128042 476380 128364 477080
rect 129064 476380 129386 477080
rect 130086 476380 130408 477080
rect 131108 476380 131430 477080
rect 132130 476380 132452 477080
rect 133152 476380 133474 477080
rect 134174 476380 134496 477080
rect 135196 476380 135518 477080
rect 136218 476380 136540 477080
rect 137240 476380 137562 477080
rect 138262 476380 138584 477080
rect 139284 476380 139606 477080
rect 140306 476380 140628 477080
rect 141328 476380 141650 477080
rect 142350 476380 142672 477080
rect 143372 476380 143694 477080
rect 144394 476380 144555 477080
rect 118930 476008 144555 476380
rect 118930 475308 119166 476008
rect 119866 475308 120188 476008
rect 120888 475308 121210 476008
rect 121910 475308 122232 476008
rect 122932 475308 123254 476008
rect 123954 475308 124276 476008
rect 124976 475308 125298 476008
rect 125998 475308 126320 476008
rect 127020 475308 127342 476008
rect 128042 475308 128364 476008
rect 129064 475308 129386 476008
rect 130086 475308 130408 476008
rect 131108 475308 131430 476008
rect 132130 475308 132452 476008
rect 133152 475308 133474 476008
rect 134174 475308 134496 476008
rect 135196 475308 135518 476008
rect 136218 475308 136540 476008
rect 137240 475308 137562 476008
rect 138262 475308 138584 476008
rect 139284 475308 139606 476008
rect 140306 475308 140628 476008
rect 141328 475308 141650 476008
rect 142350 475308 142672 476008
rect 143372 475308 143694 476008
rect 144394 475308 144555 476008
rect 118930 474936 144555 475308
rect 118930 474236 119166 474936
rect 119866 474236 120188 474936
rect 120888 474236 121210 474936
rect 121910 474236 122232 474936
rect 122932 474236 123254 474936
rect 123954 474236 124276 474936
rect 124976 474236 125298 474936
rect 125998 474236 126320 474936
rect 127020 474236 127342 474936
rect 128042 474236 128364 474936
rect 129064 474236 129386 474936
rect 130086 474236 130408 474936
rect 131108 474236 131430 474936
rect 132130 474236 132452 474936
rect 133152 474236 133474 474936
rect 134174 474236 134496 474936
rect 135196 474236 135518 474936
rect 136218 474236 136540 474936
rect 137240 474236 137562 474936
rect 138262 474236 138584 474936
rect 139284 474236 139606 474936
rect 140306 474236 140628 474936
rect 141328 474236 141650 474936
rect 142350 474236 142672 474936
rect 143372 474236 143694 474936
rect 144394 474236 144555 474936
rect 118930 473864 144555 474236
rect 118930 473164 119166 473864
rect 119866 473164 120188 473864
rect 120888 473164 121210 473864
rect 121910 473164 122232 473864
rect 122932 473164 123254 473864
rect 123954 473164 124276 473864
rect 124976 473164 125298 473864
rect 125998 473164 126320 473864
rect 127020 473164 127342 473864
rect 128042 473164 128364 473864
rect 129064 473164 129386 473864
rect 130086 473164 130408 473864
rect 131108 473164 131430 473864
rect 132130 473164 132452 473864
rect 133152 473164 133474 473864
rect 134174 473164 134496 473864
rect 135196 473164 135518 473864
rect 136218 473164 136540 473864
rect 137240 473164 137562 473864
rect 138262 473164 138584 473864
rect 139284 473164 139606 473864
rect 140306 473164 140628 473864
rect 141328 473164 141650 473864
rect 142350 473164 142672 473864
rect 143372 473164 143694 473864
rect 144394 473164 144555 473864
rect 118930 472792 144555 473164
rect 118930 472092 119166 472792
rect 119866 472092 120188 472792
rect 120888 472092 121210 472792
rect 121910 472092 122232 472792
rect 122932 472092 123254 472792
rect 123954 472092 124276 472792
rect 124976 472092 125298 472792
rect 125998 472092 126320 472792
rect 127020 472092 127342 472792
rect 128042 472092 128364 472792
rect 129064 472092 129386 472792
rect 130086 472092 130408 472792
rect 131108 472092 131430 472792
rect 132130 472092 132452 472792
rect 133152 472092 133474 472792
rect 134174 472092 134496 472792
rect 135196 472092 135518 472792
rect 136218 472092 136540 472792
rect 137240 472092 137562 472792
rect 138262 472092 138584 472792
rect 139284 472092 139606 472792
rect 140306 472092 140628 472792
rect 141328 472092 141650 472792
rect 142350 472092 142672 472792
rect 143372 472092 143694 472792
rect 144394 472092 144555 472792
rect 118930 471720 144555 472092
rect 118930 471020 119166 471720
rect 119866 471020 120188 471720
rect 120888 471020 121210 471720
rect 121910 471020 122232 471720
rect 122932 471020 123254 471720
rect 123954 471020 124276 471720
rect 124976 471020 125298 471720
rect 125998 471020 126320 471720
rect 127020 471020 127342 471720
rect 128042 471020 128364 471720
rect 129064 471020 129386 471720
rect 130086 471020 130408 471720
rect 131108 471020 131430 471720
rect 132130 471020 132452 471720
rect 133152 471020 133474 471720
rect 134174 471020 134496 471720
rect 135196 471020 135518 471720
rect 136218 471020 136540 471720
rect 137240 471020 137562 471720
rect 138262 471020 138584 471720
rect 139284 471020 139606 471720
rect 140306 471020 140628 471720
rect 141328 471020 141650 471720
rect 142350 471020 142672 471720
rect 143372 471020 143694 471720
rect 144394 471020 144555 471720
rect 118930 470648 144555 471020
rect 118930 469948 119166 470648
rect 119866 469948 120188 470648
rect 120888 469948 121210 470648
rect 121910 469948 122232 470648
rect 122932 469948 123254 470648
rect 123954 469948 124276 470648
rect 124976 469948 125298 470648
rect 125998 469948 126320 470648
rect 127020 469948 127342 470648
rect 128042 469948 128364 470648
rect 129064 469948 129386 470648
rect 130086 469948 130408 470648
rect 131108 469948 131430 470648
rect 132130 469948 132452 470648
rect 133152 469948 133474 470648
rect 134174 469948 134496 470648
rect 135196 469948 135518 470648
rect 136218 469948 136540 470648
rect 137240 469948 137562 470648
rect 138262 469948 138584 470648
rect 139284 469948 139606 470648
rect 140306 469948 140628 470648
rect 141328 469948 141650 470648
rect 142350 469948 142672 470648
rect 143372 469948 143694 470648
rect 144394 469948 144555 470648
rect 118930 469576 144555 469948
rect 118930 468876 119166 469576
rect 119866 468876 120188 469576
rect 120888 468876 121210 469576
rect 121910 468876 122232 469576
rect 122932 468876 123254 469576
rect 123954 468876 124276 469576
rect 124976 468876 125298 469576
rect 125998 468876 126320 469576
rect 127020 468876 127342 469576
rect 128042 468876 128364 469576
rect 129064 468876 129386 469576
rect 130086 468876 130408 469576
rect 131108 468876 131430 469576
rect 132130 468876 132452 469576
rect 133152 468876 133474 469576
rect 134174 468876 134496 469576
rect 135196 468876 135518 469576
rect 136218 468876 136540 469576
rect 137240 468876 137562 469576
rect 138262 468876 138584 469576
rect 139284 468876 139606 469576
rect 140306 468876 140628 469576
rect 141328 468876 141650 469576
rect 142350 468876 142672 469576
rect 143372 468876 143694 469576
rect 144394 468876 144555 469576
rect 118930 468504 144555 468876
rect 118930 467804 119166 468504
rect 119866 467804 120188 468504
rect 120888 467804 121210 468504
rect 121910 467804 122232 468504
rect 122932 467804 123254 468504
rect 123954 467804 124276 468504
rect 124976 467804 125298 468504
rect 125998 467804 126320 468504
rect 127020 467804 127342 468504
rect 128042 467804 128364 468504
rect 129064 467804 129386 468504
rect 130086 467804 130408 468504
rect 131108 467804 131430 468504
rect 132130 467804 132452 468504
rect 133152 467804 133474 468504
rect 134174 467804 134496 468504
rect 135196 467804 135518 468504
rect 136218 467804 136540 468504
rect 137240 467804 137562 468504
rect 138262 467804 138584 468504
rect 139284 467804 139606 468504
rect 140306 467804 140628 468504
rect 141328 467804 141650 468504
rect 142350 467804 142672 468504
rect 143372 467804 143694 468504
rect 144394 467804 144555 468504
rect 118930 467432 144555 467804
rect 118930 466732 119166 467432
rect 119866 466732 120188 467432
rect 120888 466732 121210 467432
rect 121910 466732 122232 467432
rect 122932 466732 123254 467432
rect 123954 466732 124276 467432
rect 124976 466732 125298 467432
rect 125998 466732 126320 467432
rect 127020 466732 127342 467432
rect 128042 466732 128364 467432
rect 129064 466732 129386 467432
rect 130086 466732 130408 467432
rect 131108 466732 131430 467432
rect 132130 466732 132452 467432
rect 133152 466732 133474 467432
rect 134174 466732 134496 467432
rect 135196 466732 135518 467432
rect 136218 466732 136540 467432
rect 137240 466732 137562 467432
rect 138262 466732 138584 467432
rect 139284 466732 139606 467432
rect 140306 466732 140628 467432
rect 141328 466732 141650 467432
rect 142350 466732 142672 467432
rect 143372 466732 143694 467432
rect 144394 466732 144555 467432
rect 118930 466360 144555 466732
rect 118930 465660 119166 466360
rect 119866 465660 120188 466360
rect 120888 465660 121210 466360
rect 121910 465660 122232 466360
rect 122932 465660 123254 466360
rect 123954 465660 124276 466360
rect 124976 465660 125298 466360
rect 125998 465660 126320 466360
rect 127020 465660 127342 466360
rect 128042 465660 128364 466360
rect 129064 465660 129386 466360
rect 130086 465660 130408 466360
rect 131108 465660 131430 466360
rect 132130 465660 132452 466360
rect 133152 465660 133474 466360
rect 134174 465660 134496 466360
rect 135196 465660 135518 466360
rect 136218 465660 136540 466360
rect 137240 465660 137562 466360
rect 138262 465660 138584 466360
rect 139284 465660 139606 466360
rect 140306 465660 140628 466360
rect 141328 465660 141650 466360
rect 142350 465660 142672 466360
rect 143372 465660 143694 466360
rect 144394 465660 144555 466360
rect 118930 465288 144555 465660
rect 118930 464588 119166 465288
rect 119866 464588 120188 465288
rect 120888 464588 121210 465288
rect 121910 464588 122232 465288
rect 122932 464588 123254 465288
rect 123954 464588 124276 465288
rect 124976 464588 125298 465288
rect 125998 464588 126320 465288
rect 127020 464588 127342 465288
rect 128042 464588 128364 465288
rect 129064 464588 129386 465288
rect 130086 464588 130408 465288
rect 131108 464588 131430 465288
rect 132130 464588 132452 465288
rect 133152 464588 133474 465288
rect 134174 464588 134496 465288
rect 135196 464588 135518 465288
rect 136218 464588 136540 465288
rect 137240 464588 137562 465288
rect 138262 464588 138584 465288
rect 139284 464588 139606 465288
rect 140306 464588 140628 465288
rect 141328 464588 141650 465288
rect 142350 464588 142672 465288
rect 143372 464588 143694 465288
rect 144394 464588 144555 465288
rect 118930 464216 144555 464588
rect 118930 463516 119166 464216
rect 119866 463516 120188 464216
rect 120888 463516 121210 464216
rect 121910 463516 122232 464216
rect 122932 463516 123254 464216
rect 123954 463516 124276 464216
rect 124976 463516 125298 464216
rect 125998 463516 126320 464216
rect 127020 463516 127342 464216
rect 128042 463516 128364 464216
rect 129064 463516 129386 464216
rect 130086 463516 130408 464216
rect 131108 463516 131430 464216
rect 132130 463516 132452 464216
rect 133152 463516 133474 464216
rect 134174 463516 134496 464216
rect 135196 463516 135518 464216
rect 136218 463516 136540 464216
rect 137240 463516 137562 464216
rect 138262 463516 138584 464216
rect 139284 463516 139606 464216
rect 140306 463516 140628 464216
rect 141328 463516 141650 464216
rect 142350 463516 142672 464216
rect 143372 463516 143694 464216
rect 144394 463516 144555 464216
rect 118930 463144 144555 463516
rect 118930 462444 119166 463144
rect 119866 462444 120188 463144
rect 120888 462444 121210 463144
rect 121910 462444 122232 463144
rect 122932 462444 123254 463144
rect 123954 462444 124276 463144
rect 124976 462444 125298 463144
rect 125998 462444 126320 463144
rect 127020 462444 127342 463144
rect 128042 462444 128364 463144
rect 129064 462444 129386 463144
rect 130086 462444 130408 463144
rect 131108 462444 131430 463144
rect 132130 462444 132452 463144
rect 133152 462444 133474 463144
rect 134174 462444 134496 463144
rect 135196 462444 135518 463144
rect 136218 462444 136540 463144
rect 137240 462444 137562 463144
rect 138262 462444 138584 463144
rect 139284 462444 139606 463144
rect 140306 462444 140628 463144
rect 141328 462444 141650 463144
rect 142350 462444 142672 463144
rect 143372 462444 143694 463144
rect 144394 462444 144555 463144
rect 118930 462072 144555 462444
rect 118930 461372 119166 462072
rect 119866 461372 120188 462072
rect 120888 461372 121210 462072
rect 121910 461372 122232 462072
rect 122932 461372 123254 462072
rect 123954 461372 124276 462072
rect 124976 461372 125298 462072
rect 125998 461372 126320 462072
rect 127020 461372 127342 462072
rect 128042 461372 128364 462072
rect 129064 461372 129386 462072
rect 130086 461372 130408 462072
rect 131108 461372 131430 462072
rect 132130 461372 132452 462072
rect 133152 461372 133474 462072
rect 134174 461372 134496 462072
rect 135196 461372 135518 462072
rect 136218 461372 136540 462072
rect 137240 461372 137562 462072
rect 138262 461372 138584 462072
rect 139284 461372 139606 462072
rect 140306 461372 140628 462072
rect 141328 461372 141650 462072
rect 142350 461372 142672 462072
rect 143372 461372 143694 462072
rect 144394 461372 144555 462072
rect 118930 461000 144555 461372
rect 118930 460300 119166 461000
rect 119866 460300 120188 461000
rect 120888 460300 121210 461000
rect 121910 460300 122232 461000
rect 122932 460300 123254 461000
rect 123954 460300 124276 461000
rect 124976 460300 125298 461000
rect 125998 460300 126320 461000
rect 127020 460300 127342 461000
rect 128042 460300 128364 461000
rect 129064 460300 129386 461000
rect 130086 460300 130408 461000
rect 131108 460300 131430 461000
rect 132130 460300 132452 461000
rect 133152 460300 133474 461000
rect 134174 460300 134496 461000
rect 135196 460300 135518 461000
rect 136218 460300 136540 461000
rect 137240 460300 137562 461000
rect 138262 460300 138584 461000
rect 139284 460300 139606 461000
rect 140306 460300 140628 461000
rect 141328 460300 141650 461000
rect 142350 460300 142672 461000
rect 143372 460300 143694 461000
rect 144394 460300 144555 461000
rect 118930 459928 144555 460300
rect 118930 459228 119166 459928
rect 119866 459228 120188 459928
rect 120888 459228 121210 459928
rect 121910 459228 122232 459928
rect 122932 459228 123254 459928
rect 123954 459228 124276 459928
rect 124976 459228 125298 459928
rect 125998 459228 126320 459928
rect 127020 459228 127342 459928
rect 128042 459228 128364 459928
rect 129064 459228 129386 459928
rect 130086 459228 130408 459928
rect 131108 459228 131430 459928
rect 132130 459228 132452 459928
rect 133152 459228 133474 459928
rect 134174 459228 134496 459928
rect 135196 459228 135518 459928
rect 136218 459228 136540 459928
rect 137240 459228 137562 459928
rect 138262 459228 138584 459928
rect 139284 459228 139606 459928
rect 140306 459228 140628 459928
rect 141328 459228 141650 459928
rect 142350 459228 142672 459928
rect 143372 459228 143694 459928
rect 144394 459228 144555 459928
rect 118930 459077 144555 459228
rect 444052 480213 444322 480840
rect 445022 480213 445379 480913
rect 446079 480213 446436 480913
rect 447136 480213 447493 480913
rect 448193 480213 448550 480913
rect 449250 480213 449607 480913
rect 450307 480213 450664 480913
rect 451364 480213 451721 480913
rect 452421 480213 452778 480913
rect 453478 480213 453835 480913
rect 454535 480213 454892 480913
rect 455592 480213 455949 480913
rect 456649 480213 457006 480913
rect 457706 480213 458063 480913
rect 458763 480213 459120 480913
rect 459820 480213 460177 480913
rect 460877 480213 461234 480913
rect 461934 480213 462291 480913
rect 462991 480213 463348 480913
rect 464048 480213 464405 480913
rect 465105 480213 465462 480913
rect 466162 480213 466519 480913
rect 467219 480213 467576 480913
rect 468276 480840 468473 480913
rect 468276 480213 468505 480840
rect 444052 479841 468505 480213
rect 444052 479141 444322 479841
rect 445022 479141 445379 479841
rect 446079 479141 446436 479841
rect 447136 479141 447493 479841
rect 448193 479141 448550 479841
rect 449250 479141 449607 479841
rect 450307 479141 450664 479841
rect 451364 479141 451721 479841
rect 452421 479141 452778 479841
rect 453478 479141 453835 479841
rect 454535 479141 454892 479841
rect 455592 479141 455949 479841
rect 456649 479141 457006 479841
rect 457706 479141 458063 479841
rect 458763 479141 459120 479841
rect 459820 479141 460177 479841
rect 460877 479141 461234 479841
rect 461934 479141 462291 479841
rect 462991 479141 463348 479841
rect 464048 479141 464405 479841
rect 465105 479141 465462 479841
rect 466162 479141 466519 479841
rect 467219 479141 467576 479841
rect 468276 479141 468505 479841
rect 444052 478769 468505 479141
rect 444052 478069 444322 478769
rect 445022 478069 445379 478769
rect 446079 478069 446436 478769
rect 447136 478069 447493 478769
rect 448193 478069 448550 478769
rect 449250 478069 449607 478769
rect 450307 478069 450664 478769
rect 451364 478069 451721 478769
rect 452421 478069 452778 478769
rect 453478 478069 453835 478769
rect 454535 478069 454892 478769
rect 455592 478069 455949 478769
rect 456649 478069 457006 478769
rect 457706 478069 458063 478769
rect 458763 478069 459120 478769
rect 459820 478069 460177 478769
rect 460877 478069 461234 478769
rect 461934 478069 462291 478769
rect 462991 478069 463348 478769
rect 464048 478069 464405 478769
rect 465105 478069 465462 478769
rect 466162 478069 466519 478769
rect 467219 478069 467576 478769
rect 468276 478069 468505 478769
rect 444052 477697 468505 478069
rect 444052 476997 444322 477697
rect 445022 476997 445379 477697
rect 446079 476997 446436 477697
rect 447136 476997 447493 477697
rect 448193 476997 448550 477697
rect 449250 476997 449607 477697
rect 450307 476997 450664 477697
rect 451364 476997 451721 477697
rect 452421 476997 452778 477697
rect 453478 476997 453835 477697
rect 454535 476997 454892 477697
rect 455592 476997 455949 477697
rect 456649 476997 457006 477697
rect 457706 476997 458063 477697
rect 458763 476997 459120 477697
rect 459820 476997 460177 477697
rect 460877 476997 461234 477697
rect 461934 476997 462291 477697
rect 462991 476997 463348 477697
rect 464048 476997 464405 477697
rect 465105 476997 465462 477697
rect 466162 476997 466519 477697
rect 467219 476997 467576 477697
rect 468276 476997 468505 477697
rect 444052 476625 468505 476997
rect 444052 475925 444322 476625
rect 445022 475925 445379 476625
rect 446079 475925 446436 476625
rect 447136 475925 447493 476625
rect 448193 475925 448550 476625
rect 449250 475925 449607 476625
rect 450307 475925 450664 476625
rect 451364 475925 451721 476625
rect 452421 475925 452778 476625
rect 453478 475925 453835 476625
rect 454535 475925 454892 476625
rect 455592 475925 455949 476625
rect 456649 475925 457006 476625
rect 457706 475925 458063 476625
rect 458763 475925 459120 476625
rect 459820 475925 460177 476625
rect 460877 475925 461234 476625
rect 461934 475925 462291 476625
rect 462991 475925 463348 476625
rect 464048 475925 464405 476625
rect 465105 475925 465462 476625
rect 466162 475925 466519 476625
rect 467219 475925 467576 476625
rect 468276 475925 468505 476625
rect 444052 475553 468505 475925
rect 444052 474853 444322 475553
rect 445022 474853 445379 475553
rect 446079 474853 446436 475553
rect 447136 474853 447493 475553
rect 448193 474853 448550 475553
rect 449250 474853 449607 475553
rect 450307 474853 450664 475553
rect 451364 474853 451721 475553
rect 452421 474853 452778 475553
rect 453478 474853 453835 475553
rect 454535 474853 454892 475553
rect 455592 474853 455949 475553
rect 456649 474853 457006 475553
rect 457706 474853 458063 475553
rect 458763 474853 459120 475553
rect 459820 474853 460177 475553
rect 460877 474853 461234 475553
rect 461934 474853 462291 475553
rect 462991 474853 463348 475553
rect 464048 474853 464405 475553
rect 465105 474853 465462 475553
rect 466162 474853 466519 475553
rect 467219 474853 467576 475553
rect 468276 474853 468505 475553
rect 444052 474481 468505 474853
rect 444052 473781 444322 474481
rect 445022 473781 445379 474481
rect 446079 473781 446436 474481
rect 447136 473781 447493 474481
rect 448193 473781 448550 474481
rect 449250 473781 449607 474481
rect 450307 473781 450664 474481
rect 451364 473781 451721 474481
rect 452421 473781 452778 474481
rect 453478 473781 453835 474481
rect 454535 473781 454892 474481
rect 455592 473781 455949 474481
rect 456649 473781 457006 474481
rect 457706 473781 458063 474481
rect 458763 473781 459120 474481
rect 459820 473781 460177 474481
rect 460877 473781 461234 474481
rect 461934 473781 462291 474481
rect 462991 473781 463348 474481
rect 464048 473781 464405 474481
rect 465105 473781 465462 474481
rect 466162 473781 466519 474481
rect 467219 473781 467576 474481
rect 468276 473781 468505 474481
rect 444052 473409 468505 473781
rect 444052 472709 444322 473409
rect 445022 472709 445379 473409
rect 446079 472709 446436 473409
rect 447136 472709 447493 473409
rect 448193 472709 448550 473409
rect 449250 472709 449607 473409
rect 450307 472709 450664 473409
rect 451364 472709 451721 473409
rect 452421 472709 452778 473409
rect 453478 472709 453835 473409
rect 454535 472709 454892 473409
rect 455592 472709 455949 473409
rect 456649 472709 457006 473409
rect 457706 472709 458063 473409
rect 458763 472709 459120 473409
rect 459820 472709 460177 473409
rect 460877 472709 461234 473409
rect 461934 472709 462291 473409
rect 462991 472709 463348 473409
rect 464048 472709 464405 473409
rect 465105 472709 465462 473409
rect 466162 472709 466519 473409
rect 467219 472709 467576 473409
rect 468276 472709 468505 473409
rect 444052 472337 468505 472709
rect 444052 471637 444322 472337
rect 445022 471637 445379 472337
rect 446079 471637 446436 472337
rect 447136 471637 447493 472337
rect 448193 471637 448550 472337
rect 449250 471637 449607 472337
rect 450307 471637 450664 472337
rect 451364 471637 451721 472337
rect 452421 471637 452778 472337
rect 453478 471637 453835 472337
rect 454535 471637 454892 472337
rect 455592 471637 455949 472337
rect 456649 471637 457006 472337
rect 457706 471637 458063 472337
rect 458763 471637 459120 472337
rect 459820 471637 460177 472337
rect 460877 471637 461234 472337
rect 461934 471637 462291 472337
rect 462991 471637 463348 472337
rect 464048 471637 464405 472337
rect 465105 471637 465462 472337
rect 466162 471637 466519 472337
rect 467219 471637 467576 472337
rect 468276 471637 468505 472337
rect 444052 471265 468505 471637
rect 444052 470565 444322 471265
rect 445022 470565 445379 471265
rect 446079 470565 446436 471265
rect 447136 470565 447493 471265
rect 448193 470565 448550 471265
rect 449250 470565 449607 471265
rect 450307 470565 450664 471265
rect 451364 470565 451721 471265
rect 452421 470565 452778 471265
rect 453478 470565 453835 471265
rect 454535 470565 454892 471265
rect 455592 470565 455949 471265
rect 456649 470565 457006 471265
rect 457706 470565 458063 471265
rect 458763 470565 459120 471265
rect 459820 470565 460177 471265
rect 460877 470565 461234 471265
rect 461934 470565 462291 471265
rect 462991 470565 463348 471265
rect 464048 470565 464405 471265
rect 465105 470565 465462 471265
rect 466162 470565 466519 471265
rect 467219 470565 467576 471265
rect 468276 470565 468505 471265
rect 444052 470193 468505 470565
rect 444052 469493 444322 470193
rect 445022 469493 445379 470193
rect 446079 469493 446436 470193
rect 447136 469493 447493 470193
rect 448193 469493 448550 470193
rect 449250 469493 449607 470193
rect 450307 469493 450664 470193
rect 451364 469493 451721 470193
rect 452421 469493 452778 470193
rect 453478 469493 453835 470193
rect 454535 469493 454892 470193
rect 455592 469493 455949 470193
rect 456649 469493 457006 470193
rect 457706 469493 458063 470193
rect 458763 469493 459120 470193
rect 459820 469493 460177 470193
rect 460877 469493 461234 470193
rect 461934 469493 462291 470193
rect 462991 469493 463348 470193
rect 464048 469493 464405 470193
rect 465105 469493 465462 470193
rect 466162 469493 466519 470193
rect 467219 469493 467576 470193
rect 468276 469493 468505 470193
rect 444052 469121 468505 469493
rect 444052 468421 444322 469121
rect 445022 468421 445379 469121
rect 446079 468421 446436 469121
rect 447136 468421 447493 469121
rect 448193 468421 448550 469121
rect 449250 468421 449607 469121
rect 450307 468421 450664 469121
rect 451364 468421 451721 469121
rect 452421 468421 452778 469121
rect 453478 468421 453835 469121
rect 454535 468421 454892 469121
rect 455592 468421 455949 469121
rect 456649 468421 457006 469121
rect 457706 468421 458063 469121
rect 458763 468421 459120 469121
rect 459820 468421 460177 469121
rect 460877 468421 461234 469121
rect 461934 468421 462291 469121
rect 462991 468421 463348 469121
rect 464048 468421 464405 469121
rect 465105 468421 465462 469121
rect 466162 468421 466519 469121
rect 467219 468421 467576 469121
rect 468276 468421 468505 469121
rect 444052 468049 468505 468421
rect 444052 467349 444322 468049
rect 445022 467349 445379 468049
rect 446079 467349 446436 468049
rect 447136 467349 447493 468049
rect 448193 467349 448550 468049
rect 449250 467349 449607 468049
rect 450307 467349 450664 468049
rect 451364 467349 451721 468049
rect 452421 467349 452778 468049
rect 453478 467349 453835 468049
rect 454535 467349 454892 468049
rect 455592 467349 455949 468049
rect 456649 467349 457006 468049
rect 457706 467349 458063 468049
rect 458763 467349 459120 468049
rect 459820 467349 460177 468049
rect 460877 467349 461234 468049
rect 461934 467349 462291 468049
rect 462991 467349 463348 468049
rect 464048 467349 464405 468049
rect 465105 467349 465462 468049
rect 466162 467349 466519 468049
rect 467219 467349 467576 468049
rect 468276 467349 468505 468049
rect 444052 466977 468505 467349
rect 444052 466277 444322 466977
rect 445022 466277 445379 466977
rect 446079 466277 446436 466977
rect 447136 466277 447493 466977
rect 448193 466277 448550 466977
rect 449250 466277 449607 466977
rect 450307 466277 450664 466977
rect 451364 466277 451721 466977
rect 452421 466277 452778 466977
rect 453478 466277 453835 466977
rect 454535 466277 454892 466977
rect 455592 466277 455949 466977
rect 456649 466277 457006 466977
rect 457706 466277 458063 466977
rect 458763 466277 459120 466977
rect 459820 466277 460177 466977
rect 460877 466277 461234 466977
rect 461934 466277 462291 466977
rect 462991 466277 463348 466977
rect 464048 466277 464405 466977
rect 465105 466277 465462 466977
rect 466162 466277 466519 466977
rect 467219 466277 467576 466977
rect 468276 466277 468505 466977
rect 444052 465905 468505 466277
rect 444052 465205 444322 465905
rect 445022 465205 445379 465905
rect 446079 465205 446436 465905
rect 447136 465205 447493 465905
rect 448193 465205 448550 465905
rect 449250 465205 449607 465905
rect 450307 465205 450664 465905
rect 451364 465205 451721 465905
rect 452421 465205 452778 465905
rect 453478 465205 453835 465905
rect 454535 465205 454892 465905
rect 455592 465205 455949 465905
rect 456649 465205 457006 465905
rect 457706 465205 458063 465905
rect 458763 465205 459120 465905
rect 459820 465205 460177 465905
rect 460877 465205 461234 465905
rect 461934 465205 462291 465905
rect 462991 465205 463348 465905
rect 464048 465205 464405 465905
rect 465105 465205 465462 465905
rect 466162 465205 466519 465905
rect 467219 465205 467576 465905
rect 468276 465205 468505 465905
rect 444052 464833 468505 465205
rect 444052 464133 444322 464833
rect 445022 464133 445379 464833
rect 446079 464133 446436 464833
rect 447136 464133 447493 464833
rect 448193 464133 448550 464833
rect 449250 464133 449607 464833
rect 450307 464133 450664 464833
rect 451364 464133 451721 464833
rect 452421 464133 452778 464833
rect 453478 464133 453835 464833
rect 454535 464133 454892 464833
rect 455592 464133 455949 464833
rect 456649 464133 457006 464833
rect 457706 464133 458063 464833
rect 458763 464133 459120 464833
rect 459820 464133 460177 464833
rect 460877 464133 461234 464833
rect 461934 464133 462291 464833
rect 462991 464133 463348 464833
rect 464048 464133 464405 464833
rect 465105 464133 465462 464833
rect 466162 464133 466519 464833
rect 467219 464133 467576 464833
rect 468276 464133 468505 464833
rect 444052 463761 468505 464133
rect 444052 463061 444322 463761
rect 445022 463061 445379 463761
rect 446079 463061 446436 463761
rect 447136 463061 447493 463761
rect 448193 463061 448550 463761
rect 449250 463061 449607 463761
rect 450307 463061 450664 463761
rect 451364 463061 451721 463761
rect 452421 463061 452778 463761
rect 453478 463061 453835 463761
rect 454535 463061 454892 463761
rect 455592 463061 455949 463761
rect 456649 463061 457006 463761
rect 457706 463061 458063 463761
rect 458763 463061 459120 463761
rect 459820 463061 460177 463761
rect 460877 463061 461234 463761
rect 461934 463061 462291 463761
rect 462991 463061 463348 463761
rect 464048 463061 464405 463761
rect 465105 463061 465462 463761
rect 466162 463061 466519 463761
rect 467219 463061 467576 463761
rect 468276 463061 468505 463761
rect 444052 462689 468505 463061
rect 444052 461989 444322 462689
rect 445022 461989 445379 462689
rect 446079 461989 446436 462689
rect 447136 461989 447493 462689
rect 448193 461989 448550 462689
rect 449250 461989 449607 462689
rect 450307 461989 450664 462689
rect 451364 461989 451721 462689
rect 452421 461989 452778 462689
rect 453478 461989 453835 462689
rect 454535 461989 454892 462689
rect 455592 461989 455949 462689
rect 456649 461989 457006 462689
rect 457706 461989 458063 462689
rect 458763 461989 459120 462689
rect 459820 461989 460177 462689
rect 460877 461989 461234 462689
rect 461934 461989 462291 462689
rect 462991 461989 463348 462689
rect 464048 461989 464405 462689
rect 465105 461989 465462 462689
rect 466162 461989 466519 462689
rect 467219 461989 467576 462689
rect 468276 461989 468505 462689
rect 444052 461617 468505 461989
rect 444052 460917 444322 461617
rect 445022 460917 445379 461617
rect 446079 460917 446436 461617
rect 447136 460917 447493 461617
rect 448193 460917 448550 461617
rect 449250 460917 449607 461617
rect 450307 460917 450664 461617
rect 451364 460917 451721 461617
rect 452421 460917 452778 461617
rect 453478 460917 453835 461617
rect 454535 460917 454892 461617
rect 455592 460917 455949 461617
rect 456649 460917 457006 461617
rect 457706 460917 458063 461617
rect 458763 460917 459120 461617
rect 459820 460917 460177 461617
rect 460877 460917 461234 461617
rect 461934 460917 462291 461617
rect 462991 460917 463348 461617
rect 464048 460917 464405 461617
rect 465105 460917 465462 461617
rect 466162 460917 466519 461617
rect 467219 460917 467576 461617
rect 468276 460917 468505 461617
rect 444052 460545 468505 460917
rect 444052 459845 444322 460545
rect 445022 459845 445379 460545
rect 446079 459845 446436 460545
rect 447136 459845 447493 460545
rect 448193 459845 448550 460545
rect 449250 459845 449607 460545
rect 450307 459845 450664 460545
rect 451364 459845 451721 460545
rect 452421 459845 452778 460545
rect 453478 459845 453835 460545
rect 454535 459845 454892 460545
rect 455592 459845 455949 460545
rect 456649 459845 457006 460545
rect 457706 459845 458063 460545
rect 458763 459845 459120 460545
rect 459820 459845 460177 460545
rect 460877 459845 461234 460545
rect 461934 459845 462291 460545
rect 462991 459845 463348 460545
rect 464048 459845 464405 460545
rect 465105 459845 465462 460545
rect 466162 459845 466519 460545
rect 467219 459845 467576 460545
rect 468276 459845 468505 460545
rect 444052 459473 468505 459845
rect 118930 458967 143881 459077
rect 121375 445963 137991 458967
rect 444052 458773 444322 459473
rect 445022 458773 445379 459473
rect 446079 458773 446436 459473
rect 447136 458773 447493 459473
rect 448193 458773 448550 459473
rect 449250 458773 449607 459473
rect 450307 458773 450664 459473
rect 451364 458773 451721 459473
rect 452421 458773 452778 459473
rect 453478 458773 453835 459473
rect 454535 458773 454892 459473
rect 455592 458773 455949 459473
rect 456649 458773 457006 459473
rect 457706 458773 458063 459473
rect 458763 458773 459120 459473
rect 459820 458773 460177 459473
rect 460877 458773 461234 459473
rect 461934 458773 462291 459473
rect 462991 458773 463348 459473
rect 464048 458773 464405 459473
rect 465105 458773 465462 459473
rect 466162 458773 466519 459473
rect 467219 458773 467576 459473
rect 468276 458773 468505 459473
rect 444052 458401 468505 458773
rect 444052 457701 444322 458401
rect 445022 457701 445379 458401
rect 446079 457701 446436 458401
rect 447136 457701 447493 458401
rect 448193 457701 448550 458401
rect 449250 457701 449607 458401
rect 450307 457701 450664 458401
rect 451364 457701 451721 458401
rect 452421 457701 452778 458401
rect 453478 457701 453835 458401
rect 454535 457701 454892 458401
rect 455592 457701 455949 458401
rect 456649 457701 457006 458401
rect 457706 457701 458063 458401
rect 458763 457701 459120 458401
rect 459820 457701 460177 458401
rect 460877 457701 461234 458401
rect 461934 457701 462291 458401
rect 462991 457701 463348 458401
rect 464048 457701 464405 458401
rect 465105 457701 465462 458401
rect 466162 457701 466519 458401
rect 467219 457701 467576 458401
rect 468276 457701 468505 458401
rect 444052 457364 468505 457701
rect 121434 367981 137991 445963
rect 121127 367465 137991 367981
rect 121127 367315 122043 367465
rect 122193 367315 122311 367465
rect 122461 367315 122579 367465
rect 122729 367315 122847 367465
rect 122997 367315 123115 367465
rect 123265 367315 123383 367465
rect 123533 367315 123651 367465
rect 123801 367315 123919 367465
rect 124069 367315 124187 367465
rect 124337 367315 124455 367465
rect 124605 367315 137991 367465
rect 121127 367227 137991 367315
rect 121127 367077 122043 367227
rect 122193 367077 122311 367227
rect 122461 367077 122579 367227
rect 122729 367077 122847 367227
rect 122997 367077 123115 367227
rect 123265 367077 123383 367227
rect 123533 367077 123651 367227
rect 123801 367077 123919 367227
rect 124069 367077 124187 367227
rect 124337 367077 124455 367227
rect 124605 367077 137991 367227
rect 121127 366989 137991 367077
rect 121127 366839 122043 366989
rect 122193 366839 122311 366989
rect 122461 366839 122579 366989
rect 122729 366839 122847 366989
rect 122997 366839 123115 366989
rect 123265 366839 123383 366989
rect 123533 366839 123651 366989
rect 123801 366839 123919 366989
rect 124069 366839 124187 366989
rect 124337 366839 124455 366989
rect 124605 366839 137991 366989
rect 121127 366751 137991 366839
rect 121127 366601 122043 366751
rect 122193 366601 122311 366751
rect 122461 366601 122579 366751
rect 122729 366601 122847 366751
rect 122997 366601 123115 366751
rect 123265 366601 123383 366751
rect 123533 366601 123651 366751
rect 123801 366601 123919 366751
rect 124069 366601 124187 366751
rect 124337 366601 124455 366751
rect 124605 366601 137991 366751
rect 121127 366513 137991 366601
rect 121127 366363 122043 366513
rect 122193 366363 122311 366513
rect 122461 366363 122579 366513
rect 122729 366363 122847 366513
rect 122997 366363 123115 366513
rect 123265 366363 123383 366513
rect 123533 366363 123651 366513
rect 123801 366363 123919 366513
rect 124069 366363 124187 366513
rect 124337 366363 124455 366513
rect 124605 366363 137991 366513
rect 121127 366275 137991 366363
rect 121127 366125 122043 366275
rect 122193 366125 122311 366275
rect 122461 366125 122579 366275
rect 122729 366125 122847 366275
rect 122997 366125 123115 366275
rect 123265 366125 123383 366275
rect 123533 366125 123651 366275
rect 123801 366125 123919 366275
rect 124069 366125 124187 366275
rect 124337 366125 124455 366275
rect 124605 366125 137991 366275
rect 121127 366037 137991 366125
rect 121127 365887 122043 366037
rect 122193 365887 122311 366037
rect 122461 365887 122579 366037
rect 122729 365887 122847 366037
rect 122997 365887 123115 366037
rect 123265 365887 123383 366037
rect 123533 365887 123651 366037
rect 123801 365887 123919 366037
rect 124069 365887 124187 366037
rect 124337 365887 124455 366037
rect 124605 365887 137991 366037
rect 121127 365799 137991 365887
rect 121127 365649 122043 365799
rect 122193 365649 122311 365799
rect 122461 365649 122579 365799
rect 122729 365649 122847 365799
rect 122997 365649 123115 365799
rect 123265 365649 123383 365799
rect 123533 365649 123651 365799
rect 123801 365649 123919 365799
rect 124069 365649 124187 365799
rect 124337 365649 124455 365799
rect 124605 365649 137991 365799
rect 121127 365561 137991 365649
rect 121127 365411 122043 365561
rect 122193 365411 122311 365561
rect 122461 365411 122579 365561
rect 122729 365411 122847 365561
rect 122997 365411 123115 365561
rect 123265 365411 123383 365561
rect 123533 365411 123651 365561
rect 123801 365411 123919 365561
rect 124069 365411 124187 365561
rect 124337 365411 124455 365561
rect 124605 365411 137991 365561
rect 121127 365323 137991 365411
rect 121127 365173 122043 365323
rect 122193 365173 122311 365323
rect 122461 365173 122579 365323
rect 122729 365173 122847 365323
rect 122997 365173 123115 365323
rect 123265 365173 123383 365323
rect 123533 365173 123651 365323
rect 123801 365173 123919 365323
rect 124069 365173 124187 365323
rect 124337 365173 124455 365323
rect 124605 365173 137991 365323
rect 121127 364498 137991 365173
rect 121434 146041 137991 364498
rect 451564 150276 468121 457364
rect 443499 149850 468321 150276
rect 443499 149665 468566 149850
rect 443499 148965 443943 149665
rect 444643 148965 445021 149665
rect 445721 148965 446099 149665
rect 446799 148965 447177 149665
rect 447877 148965 448255 149665
rect 448955 148965 449333 149665
rect 450033 148965 450411 149665
rect 451111 148965 451489 149665
rect 452189 148965 452567 149665
rect 453267 148965 453645 149665
rect 454345 148965 454723 149665
rect 455423 148965 455801 149665
rect 456501 148965 456879 149665
rect 457579 148965 457957 149665
rect 458657 148965 459035 149665
rect 459735 148965 460113 149665
rect 460813 148965 461191 149665
rect 461891 148965 462269 149665
rect 462969 148965 463347 149665
rect 464047 148965 464425 149665
rect 465125 148965 465503 149665
rect 466203 148965 466581 149665
rect 467281 148965 467659 149665
rect 468359 148965 468566 149665
rect 443499 148644 468566 148965
rect 443499 147944 443943 148644
rect 444643 147944 445021 148644
rect 445721 147944 446099 148644
rect 446799 147944 447177 148644
rect 447877 147944 448255 148644
rect 448955 147944 449333 148644
rect 450033 147944 450411 148644
rect 451111 147944 451489 148644
rect 452189 147944 452567 148644
rect 453267 147944 453645 148644
rect 454345 147944 454723 148644
rect 455423 147944 455801 148644
rect 456501 147944 456879 148644
rect 457579 147944 457957 148644
rect 458657 147944 459035 148644
rect 459735 147944 460113 148644
rect 460813 147944 461191 148644
rect 461891 147944 462269 148644
rect 462969 147944 463347 148644
rect 464047 147944 464425 148644
rect 465125 147944 465503 148644
rect 466203 147944 466581 148644
rect 467281 147944 467659 148644
rect 468359 147944 468566 148644
rect 443499 147623 468566 147944
rect 443499 146923 443943 147623
rect 444643 146923 445021 147623
rect 445721 146923 446099 147623
rect 446799 146923 447177 147623
rect 447877 146923 448255 147623
rect 448955 146923 449333 147623
rect 450033 146923 450411 147623
rect 451111 146923 451489 147623
rect 452189 146923 452567 147623
rect 453267 146923 453645 147623
rect 454345 146923 454723 147623
rect 455423 146923 455801 147623
rect 456501 146923 456879 147623
rect 457579 146923 457957 147623
rect 458657 146923 459035 147623
rect 459735 146923 460113 147623
rect 460813 146923 461191 147623
rect 461891 146923 462269 147623
rect 462969 146923 463347 147623
rect 464047 146923 464425 147623
rect 465125 146923 465503 147623
rect 466203 146923 466581 147623
rect 467281 146923 467659 147623
rect 468359 146923 468566 147623
rect 443499 146602 468566 146923
rect 121369 145196 142442 146041
rect 121369 144196 121694 145196
rect 122694 144196 123035 145196
rect 124035 144196 124376 145196
rect 125376 144196 125717 145196
rect 126717 144196 127058 145196
rect 128058 144196 128399 145196
rect 129399 144196 129740 145196
rect 130740 144196 131081 145196
rect 132081 144196 132422 145196
rect 133422 144196 133763 145196
rect 134763 144196 135104 145196
rect 136104 144196 136445 145196
rect 137445 144196 137786 145196
rect 138786 144196 139127 145196
rect 140127 144196 140468 145196
rect 141468 144196 142442 145196
rect 121369 143855 142442 144196
rect 121369 142855 121694 143855
rect 122694 142855 123035 143855
rect 124035 142855 124376 143855
rect 125376 142855 125717 143855
rect 126717 142855 127058 143855
rect 128058 142855 128399 143855
rect 129399 142855 129740 143855
rect 130740 142855 131081 143855
rect 132081 142855 132422 143855
rect 133422 142855 133763 143855
rect 134763 142855 135104 143855
rect 136104 142855 136445 143855
rect 137445 142855 137786 143855
rect 138786 142855 139127 143855
rect 140127 142855 140468 143855
rect 141468 142855 142442 143855
rect 121369 142514 142442 142855
rect 121369 141514 121694 142514
rect 122694 141514 123035 142514
rect 124035 141514 124376 142514
rect 125376 141514 125717 142514
rect 126717 141514 127058 142514
rect 128058 141514 128399 142514
rect 129399 141514 129740 142514
rect 130740 141514 131081 142514
rect 132081 141514 132422 142514
rect 133422 141514 133763 142514
rect 134763 141514 135104 142514
rect 136104 141514 136445 142514
rect 137445 141514 137786 142514
rect 138786 141514 139127 142514
rect 140127 141514 140468 142514
rect 141468 141514 142442 142514
rect 121369 141173 142442 141514
rect 121369 140173 121694 141173
rect 122694 140173 123035 141173
rect 124035 140173 124376 141173
rect 125376 140173 125717 141173
rect 126717 140173 127058 141173
rect 128058 140173 128399 141173
rect 129399 140173 129740 141173
rect 130740 140173 131081 141173
rect 132081 140173 132422 141173
rect 133422 140173 133763 141173
rect 134763 140173 135104 141173
rect 136104 140173 136445 141173
rect 137445 140173 137786 141173
rect 138786 140173 139127 141173
rect 140127 140173 140468 141173
rect 141468 140173 142442 141173
rect 121369 139832 142442 140173
rect 121369 138832 121694 139832
rect 122694 138832 123035 139832
rect 124035 138832 124376 139832
rect 125376 138832 125717 139832
rect 126717 138832 127058 139832
rect 128058 138832 128399 139832
rect 129399 138832 129740 139832
rect 130740 138832 131081 139832
rect 132081 138832 132422 139832
rect 133422 138832 133763 139832
rect 134763 138832 135104 139832
rect 136104 138832 136445 139832
rect 137445 138832 137786 139832
rect 138786 138832 139127 139832
rect 140127 138832 140468 139832
rect 141468 138832 142442 139832
rect 121369 138491 142442 138832
rect 121369 137491 121694 138491
rect 122694 137491 123035 138491
rect 124035 137491 124376 138491
rect 125376 137491 125717 138491
rect 126717 137491 127058 138491
rect 128058 137491 128399 138491
rect 129399 137491 129740 138491
rect 130740 137491 131081 138491
rect 132081 137491 132422 138491
rect 133422 137491 133763 138491
rect 134763 137491 135104 138491
rect 136104 137491 136445 138491
rect 137445 137491 137786 138491
rect 138786 137491 139127 138491
rect 140127 137491 140468 138491
rect 141468 137491 142442 138491
rect 121369 137150 142442 137491
rect 121369 136150 121694 137150
rect 122694 136150 123035 137150
rect 124035 136150 124376 137150
rect 125376 136150 125717 137150
rect 126717 136150 127058 137150
rect 128058 136150 128399 137150
rect 129399 136150 129740 137150
rect 130740 136150 131081 137150
rect 132081 136150 132422 137150
rect 133422 136150 133763 137150
rect 134763 136150 135104 137150
rect 136104 136150 136445 137150
rect 137445 136150 137786 137150
rect 138786 136150 139127 137150
rect 140127 136150 140468 137150
rect 141468 136150 142442 137150
rect 121369 135809 142442 136150
rect 121369 134809 121694 135809
rect 122694 134809 123035 135809
rect 124035 134809 124376 135809
rect 125376 134809 125717 135809
rect 126717 134809 127058 135809
rect 128058 134809 128399 135809
rect 129399 134809 129740 135809
rect 130740 134809 131081 135809
rect 132081 134809 132422 135809
rect 133422 134809 133763 135809
rect 134763 134809 135104 135809
rect 136104 134809 136445 135809
rect 137445 134809 137786 135809
rect 138786 134809 139127 135809
rect 140127 134809 140468 135809
rect 141468 134809 142442 135809
rect 121369 134468 142442 134809
rect 121369 133468 121694 134468
rect 122694 133468 123035 134468
rect 124035 133468 124376 134468
rect 125376 133468 125717 134468
rect 126717 133468 127058 134468
rect 128058 133468 128399 134468
rect 129399 133468 129740 134468
rect 130740 133468 131081 134468
rect 132081 133468 132422 134468
rect 133422 133468 133763 134468
rect 134763 133468 135104 134468
rect 136104 133468 136445 134468
rect 137445 133468 137786 134468
rect 138786 133468 139127 134468
rect 140127 133468 140468 134468
rect 141468 133468 142442 134468
rect 121369 133127 142442 133468
rect 121369 132127 121694 133127
rect 122694 132127 123035 133127
rect 124035 132127 124376 133127
rect 125376 132127 125717 133127
rect 126717 132127 127058 133127
rect 128058 132127 128399 133127
rect 129399 132127 129740 133127
rect 130740 132127 131081 133127
rect 132081 132127 132422 133127
rect 133422 132127 133763 133127
rect 134763 132127 135104 133127
rect 136104 132127 136445 133127
rect 137445 132127 137786 133127
rect 138786 132127 139127 133127
rect 140127 132127 140468 133127
rect 141468 132127 142442 133127
rect 121369 131786 142442 132127
rect 121369 130786 121694 131786
rect 122694 130786 123035 131786
rect 124035 130786 124376 131786
rect 125376 130786 125717 131786
rect 126717 130786 127058 131786
rect 128058 130786 128399 131786
rect 129399 130786 129740 131786
rect 130740 130786 131081 131786
rect 132081 130786 132422 131786
rect 133422 130786 133763 131786
rect 134763 130786 135104 131786
rect 136104 130786 136445 131786
rect 137445 130786 137786 131786
rect 138786 130786 139127 131786
rect 140127 130786 140468 131786
rect 141468 130786 142442 131786
rect 121369 130445 142442 130786
rect 121369 129445 121694 130445
rect 122694 129445 123035 130445
rect 124035 129445 124376 130445
rect 125376 129445 125717 130445
rect 126717 129445 127058 130445
rect 128058 129445 128399 130445
rect 129399 129445 129740 130445
rect 130740 129445 131081 130445
rect 132081 129445 132422 130445
rect 133422 129445 133763 130445
rect 134763 129445 135104 130445
rect 136104 129445 136445 130445
rect 137445 129445 137786 130445
rect 138786 129445 139127 130445
rect 140127 129445 140468 130445
rect 141468 129445 142442 130445
rect 121369 129104 142442 129445
rect 121369 128104 121694 129104
rect 122694 128104 123035 129104
rect 124035 128104 124376 129104
rect 125376 128104 125717 129104
rect 126717 128104 127058 129104
rect 128058 128104 128399 129104
rect 129399 128104 129740 129104
rect 130740 128104 131081 129104
rect 132081 128104 132422 129104
rect 133422 128104 133763 129104
rect 134763 128104 135104 129104
rect 136104 128104 136445 129104
rect 137445 128104 137786 129104
rect 138786 128104 139127 129104
rect 140127 128104 140468 129104
rect 141468 128104 142442 129104
rect 121369 127763 142442 128104
rect 121369 126763 121694 127763
rect 122694 126763 123035 127763
rect 124035 126763 124376 127763
rect 125376 126763 125717 127763
rect 126717 126763 127058 127763
rect 128058 126763 128399 127763
rect 129399 126763 129740 127763
rect 130740 126763 131081 127763
rect 132081 126763 132422 127763
rect 133422 126763 133763 127763
rect 134763 126763 135104 127763
rect 136104 126763 136445 127763
rect 137445 126763 137786 127763
rect 138786 126763 139127 127763
rect 140127 126763 140468 127763
rect 141468 126763 142442 127763
rect 121369 126422 142442 126763
rect 121369 125422 121694 126422
rect 122694 125422 123035 126422
rect 124035 125422 124376 126422
rect 125376 125422 125717 126422
rect 126717 125422 127058 126422
rect 128058 125422 128399 126422
rect 129399 125422 129740 126422
rect 130740 125422 131081 126422
rect 132081 125422 132422 126422
rect 133422 125422 133763 126422
rect 134763 125422 135104 126422
rect 136104 125422 136445 126422
rect 137445 125422 137786 126422
rect 138786 125422 139127 126422
rect 140127 125422 140468 126422
rect 141468 125422 142442 126422
rect 121369 124678 142442 125422
rect 443499 145902 443943 146602
rect 444643 145902 445021 146602
rect 445721 145902 446099 146602
rect 446799 145902 447177 146602
rect 447877 145902 448255 146602
rect 448955 145902 449333 146602
rect 450033 145902 450411 146602
rect 451111 145902 451489 146602
rect 452189 145902 452567 146602
rect 453267 145902 453645 146602
rect 454345 145902 454723 146602
rect 455423 145902 455801 146602
rect 456501 145902 456879 146602
rect 457579 145902 457957 146602
rect 458657 145902 459035 146602
rect 459735 145902 460113 146602
rect 460813 145902 461191 146602
rect 461891 145902 462269 146602
rect 462969 145902 463347 146602
rect 464047 145902 464425 146602
rect 465125 145902 465503 146602
rect 466203 145902 466581 146602
rect 467281 145902 467659 146602
rect 468359 145902 468566 146602
rect 443499 145581 468566 145902
rect 443499 144881 443943 145581
rect 444643 144881 445021 145581
rect 445721 144881 446099 145581
rect 446799 144881 447177 145581
rect 447877 144881 448255 145581
rect 448955 144881 449333 145581
rect 450033 144881 450411 145581
rect 451111 144881 451489 145581
rect 452189 144881 452567 145581
rect 453267 144881 453645 145581
rect 454345 144881 454723 145581
rect 455423 144881 455801 145581
rect 456501 144881 456879 145581
rect 457579 144881 457957 145581
rect 458657 144881 459035 145581
rect 459735 144881 460113 145581
rect 460813 144881 461191 145581
rect 461891 144881 462269 145581
rect 462969 144881 463347 145581
rect 464047 144881 464425 145581
rect 465125 144881 465503 145581
rect 466203 144881 466581 145581
rect 467281 144881 467659 145581
rect 468359 144881 468566 145581
rect 443499 144560 468566 144881
rect 443499 143860 443943 144560
rect 444643 143860 445021 144560
rect 445721 143860 446099 144560
rect 446799 143860 447177 144560
rect 447877 143860 448255 144560
rect 448955 143860 449333 144560
rect 450033 143860 450411 144560
rect 451111 143860 451489 144560
rect 452189 143860 452567 144560
rect 453267 143860 453645 144560
rect 454345 143860 454723 144560
rect 455423 143860 455801 144560
rect 456501 143860 456879 144560
rect 457579 143860 457957 144560
rect 458657 143860 459035 144560
rect 459735 143860 460113 144560
rect 460813 143860 461191 144560
rect 461891 143860 462269 144560
rect 462969 143860 463347 144560
rect 464047 143860 464425 144560
rect 465125 143860 465503 144560
rect 466203 143860 466581 144560
rect 467281 143860 467659 144560
rect 468359 143860 468566 144560
rect 443499 143539 468566 143860
rect 443499 142839 443943 143539
rect 444643 142839 445021 143539
rect 445721 142839 446099 143539
rect 446799 142839 447177 143539
rect 447877 142839 448255 143539
rect 448955 142839 449333 143539
rect 450033 142839 450411 143539
rect 451111 142839 451489 143539
rect 452189 142839 452567 143539
rect 453267 142839 453645 143539
rect 454345 142839 454723 143539
rect 455423 142839 455801 143539
rect 456501 142839 456879 143539
rect 457579 142839 457957 143539
rect 458657 142839 459035 143539
rect 459735 142839 460113 143539
rect 460813 142839 461191 143539
rect 461891 142839 462269 143539
rect 462969 142839 463347 143539
rect 464047 142839 464425 143539
rect 465125 142839 465503 143539
rect 466203 142839 466581 143539
rect 467281 142839 467659 143539
rect 468359 142839 468566 143539
rect 443499 142518 468566 142839
rect 443499 141818 443943 142518
rect 444643 141818 445021 142518
rect 445721 141818 446099 142518
rect 446799 141818 447177 142518
rect 447877 141818 448255 142518
rect 448955 141818 449333 142518
rect 450033 141818 450411 142518
rect 451111 141818 451489 142518
rect 452189 141818 452567 142518
rect 453267 141818 453645 142518
rect 454345 141818 454723 142518
rect 455423 141818 455801 142518
rect 456501 141818 456879 142518
rect 457579 141818 457957 142518
rect 458657 141818 459035 142518
rect 459735 141818 460113 142518
rect 460813 141818 461191 142518
rect 461891 141818 462269 142518
rect 462969 141818 463347 142518
rect 464047 141818 464425 142518
rect 465125 141818 465503 142518
rect 466203 141818 466581 142518
rect 467281 141818 467659 142518
rect 468359 141818 468566 142518
rect 443499 141497 468566 141818
rect 443499 140797 443943 141497
rect 444643 140797 445021 141497
rect 445721 140797 446099 141497
rect 446799 140797 447177 141497
rect 447877 140797 448255 141497
rect 448955 140797 449333 141497
rect 450033 140797 450411 141497
rect 451111 140797 451489 141497
rect 452189 140797 452567 141497
rect 453267 140797 453645 141497
rect 454345 140797 454723 141497
rect 455423 140797 455801 141497
rect 456501 140797 456879 141497
rect 457579 140797 457957 141497
rect 458657 140797 459035 141497
rect 459735 140797 460113 141497
rect 460813 140797 461191 141497
rect 461891 140797 462269 141497
rect 462969 140797 463347 141497
rect 464047 140797 464425 141497
rect 465125 140797 465503 141497
rect 466203 140797 466581 141497
rect 467281 140797 467659 141497
rect 468359 140797 468566 141497
rect 443499 140476 468566 140797
rect 443499 139776 443943 140476
rect 444643 139776 445021 140476
rect 445721 139776 446099 140476
rect 446799 139776 447177 140476
rect 447877 139776 448255 140476
rect 448955 139776 449333 140476
rect 450033 139776 450411 140476
rect 451111 139776 451489 140476
rect 452189 139776 452567 140476
rect 453267 139776 453645 140476
rect 454345 139776 454723 140476
rect 455423 139776 455801 140476
rect 456501 139776 456879 140476
rect 457579 139776 457957 140476
rect 458657 139776 459035 140476
rect 459735 139776 460113 140476
rect 460813 139776 461191 140476
rect 461891 139776 462269 140476
rect 462969 139776 463347 140476
rect 464047 139776 464425 140476
rect 465125 139776 465503 140476
rect 466203 139776 466581 140476
rect 467281 139776 467659 140476
rect 468359 139776 468566 140476
rect 443499 139455 468566 139776
rect 443499 138755 443943 139455
rect 444643 138755 445021 139455
rect 445721 138755 446099 139455
rect 446799 138755 447177 139455
rect 447877 138755 448255 139455
rect 448955 138755 449333 139455
rect 450033 138755 450411 139455
rect 451111 138755 451489 139455
rect 452189 138755 452567 139455
rect 453267 138755 453645 139455
rect 454345 138755 454723 139455
rect 455423 138755 455801 139455
rect 456501 138755 456879 139455
rect 457579 138755 457957 139455
rect 458657 138755 459035 139455
rect 459735 138755 460113 139455
rect 460813 138755 461191 139455
rect 461891 138755 462269 139455
rect 462969 138755 463347 139455
rect 464047 138755 464425 139455
rect 465125 138755 465503 139455
rect 466203 138755 466581 139455
rect 467281 138755 467659 139455
rect 468359 138755 468566 139455
rect 443499 138434 468566 138755
rect 443499 137734 443943 138434
rect 444643 137734 445021 138434
rect 445721 137734 446099 138434
rect 446799 137734 447177 138434
rect 447877 137734 448255 138434
rect 448955 137734 449333 138434
rect 450033 137734 450411 138434
rect 451111 137734 451489 138434
rect 452189 137734 452567 138434
rect 453267 137734 453645 138434
rect 454345 137734 454723 138434
rect 455423 137734 455801 138434
rect 456501 137734 456879 138434
rect 457579 137734 457957 138434
rect 458657 137734 459035 138434
rect 459735 137734 460113 138434
rect 460813 137734 461191 138434
rect 461891 137734 462269 138434
rect 462969 137734 463347 138434
rect 464047 137734 464425 138434
rect 465125 137734 465503 138434
rect 466203 137734 466581 138434
rect 467281 137734 467659 138434
rect 468359 137734 468566 138434
rect 443499 137413 468566 137734
rect 443499 136713 443943 137413
rect 444643 136713 445021 137413
rect 445721 136713 446099 137413
rect 446799 136713 447177 137413
rect 447877 136713 448255 137413
rect 448955 136713 449333 137413
rect 450033 136713 450411 137413
rect 451111 136713 451489 137413
rect 452189 136713 452567 137413
rect 453267 136713 453645 137413
rect 454345 136713 454723 137413
rect 455423 136713 455801 137413
rect 456501 136713 456879 137413
rect 457579 136713 457957 137413
rect 458657 136713 459035 137413
rect 459735 136713 460113 137413
rect 460813 136713 461191 137413
rect 461891 136713 462269 137413
rect 462969 136713 463347 137413
rect 464047 136713 464425 137413
rect 465125 136713 465503 137413
rect 466203 136713 466581 137413
rect 467281 136713 467659 137413
rect 468359 136713 468566 137413
rect 443499 136392 468566 136713
rect 443499 135692 443943 136392
rect 444643 135692 445021 136392
rect 445721 135692 446099 136392
rect 446799 135692 447177 136392
rect 447877 135692 448255 136392
rect 448955 135692 449333 136392
rect 450033 135692 450411 136392
rect 451111 135692 451489 136392
rect 452189 135692 452567 136392
rect 453267 135692 453645 136392
rect 454345 135692 454723 136392
rect 455423 135692 455801 136392
rect 456501 135692 456879 136392
rect 457579 135692 457957 136392
rect 458657 135692 459035 136392
rect 459735 135692 460113 136392
rect 460813 135692 461191 136392
rect 461891 135692 462269 136392
rect 462969 135692 463347 136392
rect 464047 135692 464425 136392
rect 465125 135692 465503 136392
rect 466203 135692 466581 136392
rect 467281 135692 467659 136392
rect 468359 135692 468566 136392
rect 443499 135371 468566 135692
rect 443499 134671 443943 135371
rect 444643 134671 445021 135371
rect 445721 134671 446099 135371
rect 446799 134671 447177 135371
rect 447877 134671 448255 135371
rect 448955 134671 449333 135371
rect 450033 134671 450411 135371
rect 451111 134671 451489 135371
rect 452189 134671 452567 135371
rect 453267 134671 453645 135371
rect 454345 134671 454723 135371
rect 455423 134671 455801 135371
rect 456501 134671 456879 135371
rect 457579 134671 457957 135371
rect 458657 134671 459035 135371
rect 459735 134671 460113 135371
rect 460813 134671 461191 135371
rect 461891 134671 462269 135371
rect 462969 134671 463347 135371
rect 464047 134671 464425 135371
rect 465125 134671 465503 135371
rect 466203 134671 466581 135371
rect 467281 134671 467659 135371
rect 468359 134671 468566 135371
rect 443499 134350 468566 134671
rect 443499 133650 443943 134350
rect 444643 133650 445021 134350
rect 445721 133650 446099 134350
rect 446799 133650 447177 134350
rect 447877 133650 448255 134350
rect 448955 133650 449333 134350
rect 450033 133650 450411 134350
rect 451111 133650 451489 134350
rect 452189 133650 452567 134350
rect 453267 133650 453645 134350
rect 454345 133650 454723 134350
rect 455423 133650 455801 134350
rect 456501 133650 456879 134350
rect 457579 133650 457957 134350
rect 458657 133650 459035 134350
rect 459735 133650 460113 134350
rect 460813 133650 461191 134350
rect 461891 133650 462269 134350
rect 462969 133650 463347 134350
rect 464047 133650 464425 134350
rect 465125 133650 465503 134350
rect 466203 133650 466581 134350
rect 467281 133650 467659 134350
rect 468359 133650 468566 134350
rect 443499 133329 468566 133650
rect 443499 132629 443943 133329
rect 444643 132629 445021 133329
rect 445721 132629 446099 133329
rect 446799 132629 447177 133329
rect 447877 132629 448255 133329
rect 448955 132629 449333 133329
rect 450033 132629 450411 133329
rect 451111 132629 451489 133329
rect 452189 132629 452567 133329
rect 453267 132629 453645 133329
rect 454345 132629 454723 133329
rect 455423 132629 455801 133329
rect 456501 132629 456879 133329
rect 457579 132629 457957 133329
rect 458657 132629 459035 133329
rect 459735 132629 460113 133329
rect 460813 132629 461191 133329
rect 461891 132629 462269 133329
rect 462969 132629 463347 133329
rect 464047 132629 464425 133329
rect 465125 132629 465503 133329
rect 466203 132629 466581 133329
rect 467281 132629 467659 133329
rect 468359 132629 468566 133329
rect 443499 132308 468566 132629
rect 443499 131608 443943 132308
rect 444643 131608 445021 132308
rect 445721 131608 446099 132308
rect 446799 131608 447177 132308
rect 447877 131608 448255 132308
rect 448955 131608 449333 132308
rect 450033 131608 450411 132308
rect 451111 131608 451489 132308
rect 452189 131608 452567 132308
rect 453267 131608 453645 132308
rect 454345 131608 454723 132308
rect 455423 131608 455801 132308
rect 456501 131608 456879 132308
rect 457579 131608 457957 132308
rect 458657 131608 459035 132308
rect 459735 131608 460113 132308
rect 460813 131608 461191 132308
rect 461891 131608 462269 132308
rect 462969 131608 463347 132308
rect 464047 131608 464425 132308
rect 465125 131608 465503 132308
rect 466203 131608 466581 132308
rect 467281 131608 467659 132308
rect 468359 131608 468566 132308
rect 443499 131287 468566 131608
rect 443499 130587 443943 131287
rect 444643 130587 445021 131287
rect 445721 130587 446099 131287
rect 446799 130587 447177 131287
rect 447877 130587 448255 131287
rect 448955 130587 449333 131287
rect 450033 130587 450411 131287
rect 451111 130587 451489 131287
rect 452189 130587 452567 131287
rect 453267 130587 453645 131287
rect 454345 130587 454723 131287
rect 455423 130587 455801 131287
rect 456501 130587 456879 131287
rect 457579 130587 457957 131287
rect 458657 130587 459035 131287
rect 459735 130587 460113 131287
rect 460813 130587 461191 131287
rect 461891 130587 462269 131287
rect 462969 130587 463347 131287
rect 464047 130587 464425 131287
rect 465125 130587 465503 131287
rect 466203 130587 466581 131287
rect 467281 130587 467659 131287
rect 468359 130587 468566 131287
rect 443499 130266 468566 130587
rect 443499 129566 443943 130266
rect 444643 129566 445021 130266
rect 445721 129566 446099 130266
rect 446799 129566 447177 130266
rect 447877 129566 448255 130266
rect 448955 129566 449333 130266
rect 450033 129566 450411 130266
rect 451111 129566 451489 130266
rect 452189 129566 452567 130266
rect 453267 129566 453645 130266
rect 454345 129566 454723 130266
rect 455423 129566 455801 130266
rect 456501 129566 456879 130266
rect 457579 129566 457957 130266
rect 458657 129566 459035 130266
rect 459735 129566 460113 130266
rect 460813 129566 461191 130266
rect 461891 129566 462269 130266
rect 462969 129566 463347 130266
rect 464047 129566 464425 130266
rect 465125 129566 465503 130266
rect 466203 129566 466581 130266
rect 467281 129566 467659 130266
rect 468359 129566 468566 130266
rect 443499 129245 468566 129566
rect 443499 128545 443943 129245
rect 444643 128545 445021 129245
rect 445721 128545 446099 129245
rect 446799 128545 447177 129245
rect 447877 128545 448255 129245
rect 448955 128545 449333 129245
rect 450033 128545 450411 129245
rect 451111 128545 451489 129245
rect 452189 128545 452567 129245
rect 453267 128545 453645 129245
rect 454345 128545 454723 129245
rect 455423 128545 455801 129245
rect 456501 128545 456879 129245
rect 457579 128545 457957 129245
rect 458657 128545 459035 129245
rect 459735 128545 460113 129245
rect 460813 128545 461191 129245
rect 461891 128545 462269 129245
rect 462969 128545 463347 129245
rect 464047 128545 464425 129245
rect 465125 128545 465503 129245
rect 466203 128545 466581 129245
rect 467281 128545 467659 129245
rect 468359 128545 468566 129245
rect 443499 128224 468566 128545
rect 443499 127524 443943 128224
rect 444643 127524 445021 128224
rect 445721 127524 446099 128224
rect 446799 127524 447177 128224
rect 447877 127524 448255 128224
rect 448955 127524 449333 128224
rect 450033 127524 450411 128224
rect 451111 127524 451489 128224
rect 452189 127524 452567 128224
rect 453267 127524 453645 128224
rect 454345 127524 454723 128224
rect 455423 127524 455801 128224
rect 456501 127524 456879 128224
rect 457579 127524 457957 128224
rect 458657 127524 459035 128224
rect 459735 127524 460113 128224
rect 460813 127524 461191 128224
rect 461891 127524 462269 128224
rect 462969 127524 463347 128224
rect 464047 127524 464425 128224
rect 465125 127524 465503 128224
rect 466203 127524 466581 128224
rect 467281 127524 467659 128224
rect 468359 127524 468566 128224
rect 443499 127203 468566 127524
rect 443499 126503 443943 127203
rect 444643 126503 445021 127203
rect 445721 126503 446099 127203
rect 446799 126503 447177 127203
rect 447877 126503 448255 127203
rect 448955 126503 449333 127203
rect 450033 126503 450411 127203
rect 451111 126503 451489 127203
rect 452189 126503 452567 127203
rect 453267 126503 453645 127203
rect 454345 126503 454723 127203
rect 455423 126503 455801 127203
rect 456501 126503 456879 127203
rect 457579 126503 457957 127203
rect 458657 126503 459035 127203
rect 459735 126503 460113 127203
rect 460813 126503 461191 127203
rect 461891 126503 462269 127203
rect 462969 126503 463347 127203
rect 464047 126503 464425 127203
rect 465125 126503 465503 127203
rect 466203 126503 466581 127203
rect 467281 126503 467659 127203
rect 468359 126503 468566 127203
rect 443499 126182 468566 126503
rect 443499 125482 443943 126182
rect 444643 125482 445021 126182
rect 445721 125482 446099 126182
rect 446799 125482 447177 126182
rect 447877 125482 448255 126182
rect 448955 125482 449333 126182
rect 450033 125482 450411 126182
rect 451111 125482 451489 126182
rect 452189 125482 452567 126182
rect 453267 125482 453645 126182
rect 454345 125482 454723 126182
rect 455423 125482 455801 126182
rect 456501 125482 456879 126182
rect 457579 125482 457957 126182
rect 458657 125482 459035 126182
rect 459735 125482 460113 126182
rect 460813 125482 461191 126182
rect 461891 125482 462269 126182
rect 462969 125482 463347 126182
rect 464047 125482 464425 126182
rect 465125 125482 465503 126182
rect 466203 125482 466581 126182
rect 467281 125482 467659 126182
rect 468359 125482 468566 126182
rect 443499 125346 468566 125482
rect 443499 125098 468321 125346
rect 485637 125045 502194 482808
rect 481895 124824 508199 125045
rect 481895 124124 482072 124824
rect 482772 124124 483168 124824
rect 483868 124124 484264 124824
rect 484964 124124 485360 124824
rect 486060 124124 486456 124824
rect 487156 124124 487552 124824
rect 488252 124124 488648 124824
rect 489348 124124 489744 124824
rect 490444 124124 490840 124824
rect 491540 124124 491936 124824
rect 492636 124124 493032 124824
rect 493732 124124 494128 124824
rect 494828 124124 495224 124824
rect 495924 124124 496320 124824
rect 497020 124124 497416 124824
rect 498116 124124 498512 124824
rect 499212 124124 499608 124824
rect 500308 124124 500704 124824
rect 501404 124124 501800 124824
rect 502500 124124 502896 124824
rect 503596 124124 503992 124824
rect 504692 124124 505088 124824
rect 505788 124124 506184 124824
rect 506884 124124 507280 124824
rect 507980 124124 508199 124824
rect 481895 123677 508199 124124
rect 481670 123673 508199 123677
rect 481670 122973 482072 123673
rect 482772 122973 483168 123673
rect 483868 122973 484264 123673
rect 484964 122973 485360 123673
rect 486060 122973 486456 123673
rect 487156 122973 487552 123673
rect 488252 122973 488648 123673
rect 489348 122973 489744 123673
rect 490444 122973 490840 123673
rect 491540 122973 491936 123673
rect 492636 122973 493032 123673
rect 493732 122973 494128 123673
rect 494828 122973 495224 123673
rect 495924 122973 496320 123673
rect 497020 122973 497416 123673
rect 498116 122973 498512 123673
rect 499212 122973 499608 123673
rect 500308 122973 500704 123673
rect 501404 122973 501800 123673
rect 502500 122973 502896 123673
rect 503596 122973 503992 123673
rect 504692 122973 505088 123673
rect 505788 122973 506184 123673
rect 506884 122973 507280 123673
rect 507980 122973 508199 123673
rect 481670 122522 508199 122973
rect 481670 121822 482072 122522
rect 482772 121822 483168 122522
rect 483868 121822 484264 122522
rect 484964 121822 485360 122522
rect 486060 121822 486456 122522
rect 487156 121822 487552 122522
rect 488252 121822 488648 122522
rect 489348 121822 489744 122522
rect 490444 121822 490840 122522
rect 491540 121822 491936 122522
rect 492636 121822 493032 122522
rect 493732 121822 494128 122522
rect 494828 121822 495224 122522
rect 495924 121822 496320 122522
rect 497020 121822 497416 122522
rect 498116 121822 498512 122522
rect 499212 121822 499608 122522
rect 500308 121822 500704 122522
rect 501404 121822 501800 122522
rect 502500 121822 502896 122522
rect 503596 121822 503992 122522
rect 504692 121822 505088 122522
rect 505788 121822 506184 122522
rect 506884 121822 507280 122522
rect 507980 121822 508199 122522
rect 481670 121371 508199 121822
rect 481670 120671 482072 121371
rect 482772 120671 483168 121371
rect 483868 120671 484264 121371
rect 484964 120671 485360 121371
rect 486060 120671 486456 121371
rect 487156 120671 487552 121371
rect 488252 120671 488648 121371
rect 489348 120671 489744 121371
rect 490444 120671 490840 121371
rect 491540 120671 491936 121371
rect 492636 120671 493032 121371
rect 493732 120671 494128 121371
rect 494828 120671 495224 121371
rect 495924 120671 496320 121371
rect 497020 120671 497416 121371
rect 498116 120671 498512 121371
rect 499212 120671 499608 121371
rect 500308 120671 500704 121371
rect 501404 120671 501800 121371
rect 502500 120671 502896 121371
rect 503596 120671 503992 121371
rect 504692 120671 505088 121371
rect 505788 120671 506184 121371
rect 506884 120671 507280 121371
rect 507980 120671 508199 121371
rect 88384 119846 111541 120594
rect 88384 119146 89225 119846
rect 89925 119146 90134 119846
rect 90834 119146 91043 119846
rect 91743 119146 91952 119846
rect 92652 119146 92861 119846
rect 93561 119146 93770 119846
rect 94470 119146 94679 119846
rect 95379 119146 95588 119846
rect 96288 119146 96497 119846
rect 97197 119146 97406 119846
rect 98106 119146 98315 119846
rect 99015 119146 99224 119846
rect 99924 119146 100133 119846
rect 100833 119146 101042 119846
rect 101742 119146 101951 119846
rect 102651 119146 102860 119846
rect 103560 119146 103769 119846
rect 104469 119146 104678 119846
rect 105378 119146 105587 119846
rect 106287 119146 106496 119846
rect 107196 119146 107405 119846
rect 108105 119146 108314 119846
rect 109014 119146 109223 119846
rect 109923 119146 110132 119846
rect 110832 119146 111541 119846
rect 88384 118958 111541 119146
rect 88384 118258 89225 118958
rect 89925 118258 90134 118958
rect 90834 118258 91043 118958
rect 91743 118258 91952 118958
rect 92652 118258 92861 118958
rect 93561 118258 93770 118958
rect 94470 118258 94679 118958
rect 95379 118258 95588 118958
rect 96288 118258 96497 118958
rect 97197 118258 97406 118958
rect 98106 118258 98315 118958
rect 99015 118258 99224 118958
rect 99924 118258 100133 118958
rect 100833 118258 101042 118958
rect 101742 118258 101951 118958
rect 102651 118258 102860 118958
rect 103560 118258 103769 118958
rect 104469 118258 104678 118958
rect 105378 118258 105587 118958
rect 106287 118258 106496 118958
rect 107196 118258 107405 118958
rect 108105 118258 108314 118958
rect 109014 118258 109223 118958
rect 109923 118258 110132 118958
rect 110832 118258 111541 118958
rect 88384 118070 111541 118258
rect 88384 117370 89225 118070
rect 89925 117370 90134 118070
rect 90834 117370 91043 118070
rect 91743 117370 91952 118070
rect 92652 117370 92861 118070
rect 93561 117370 93770 118070
rect 94470 117370 94679 118070
rect 95379 117370 95588 118070
rect 96288 117370 96497 118070
rect 97197 117370 97406 118070
rect 98106 117370 98315 118070
rect 99015 117370 99224 118070
rect 99924 117370 100133 118070
rect 100833 117370 101042 118070
rect 101742 117370 101951 118070
rect 102651 117370 102860 118070
rect 103560 117370 103769 118070
rect 104469 117370 104678 118070
rect 105378 117370 105587 118070
rect 106287 117370 106496 118070
rect 107196 117370 107405 118070
rect 108105 117370 108314 118070
rect 109014 117370 109223 118070
rect 109923 117370 110132 118070
rect 110832 117370 111541 118070
rect 88384 117182 111541 117370
rect 88384 116482 89225 117182
rect 89925 116482 90134 117182
rect 90834 116482 91043 117182
rect 91743 116482 91952 117182
rect 92652 116482 92861 117182
rect 93561 116482 93770 117182
rect 94470 116482 94679 117182
rect 95379 116482 95588 117182
rect 96288 116482 96497 117182
rect 97197 116482 97406 117182
rect 98106 116482 98315 117182
rect 99015 116482 99224 117182
rect 99924 116482 100133 117182
rect 100833 116482 101042 117182
rect 101742 116482 101951 117182
rect 102651 116482 102860 117182
rect 103560 116482 103769 117182
rect 104469 116482 104678 117182
rect 105378 116482 105587 117182
rect 106287 116482 106496 117182
rect 107196 116482 107405 117182
rect 108105 116482 108314 117182
rect 109014 116482 109223 117182
rect 109923 116482 110132 117182
rect 110832 116482 111541 117182
rect 88384 116294 111541 116482
rect 88384 115594 89225 116294
rect 89925 115594 90134 116294
rect 90834 115594 91043 116294
rect 91743 115594 91952 116294
rect 92652 115594 92861 116294
rect 93561 115594 93770 116294
rect 94470 115594 94679 116294
rect 95379 115594 95588 116294
rect 96288 115594 96497 116294
rect 97197 115594 97406 116294
rect 98106 115594 98315 116294
rect 99015 115594 99224 116294
rect 99924 115594 100133 116294
rect 100833 115594 101042 116294
rect 101742 115594 101951 116294
rect 102651 115594 102860 116294
rect 103560 115594 103769 116294
rect 104469 115594 104678 116294
rect 105378 115594 105587 116294
rect 106287 115594 106496 116294
rect 107196 115594 107405 116294
rect 108105 115594 108314 116294
rect 109014 115594 109223 116294
rect 109923 115594 110132 116294
rect 110832 115594 111541 116294
rect 88384 115406 111541 115594
rect 88384 114706 89225 115406
rect 89925 114706 90134 115406
rect 90834 114706 91043 115406
rect 91743 114706 91952 115406
rect 92652 114706 92861 115406
rect 93561 114706 93770 115406
rect 94470 114706 94679 115406
rect 95379 114706 95588 115406
rect 96288 114706 96497 115406
rect 97197 114706 97406 115406
rect 98106 114706 98315 115406
rect 99015 114706 99224 115406
rect 99924 114706 100133 115406
rect 100833 114706 101042 115406
rect 101742 114706 101951 115406
rect 102651 114706 102860 115406
rect 103560 114706 103769 115406
rect 104469 114706 104678 115406
rect 105378 114706 105587 115406
rect 106287 114706 106496 115406
rect 107196 114706 107405 115406
rect 108105 114706 108314 115406
rect 109014 114706 109223 115406
rect 109923 114706 110132 115406
rect 110832 114706 111541 115406
rect 88384 114518 111541 114706
rect 88384 113818 89225 114518
rect 89925 113818 90134 114518
rect 90834 113818 91043 114518
rect 91743 113818 91952 114518
rect 92652 113818 92861 114518
rect 93561 113818 93770 114518
rect 94470 113818 94679 114518
rect 95379 113818 95588 114518
rect 96288 113818 96497 114518
rect 97197 113818 97406 114518
rect 98106 113818 98315 114518
rect 99015 113818 99224 114518
rect 99924 113818 100133 114518
rect 100833 113818 101042 114518
rect 101742 113818 101951 114518
rect 102651 113818 102860 114518
rect 103560 113818 103769 114518
rect 104469 113818 104678 114518
rect 105378 113818 105587 114518
rect 106287 113818 106496 114518
rect 107196 113818 107405 114518
rect 108105 113818 108314 114518
rect 109014 113818 109223 114518
rect 109923 113818 110132 114518
rect 110832 113818 111541 114518
rect 88384 113630 111541 113818
rect 88384 112930 89225 113630
rect 89925 112930 90134 113630
rect 90834 112930 91043 113630
rect 91743 112930 91952 113630
rect 92652 112930 92861 113630
rect 93561 112930 93770 113630
rect 94470 112930 94679 113630
rect 95379 112930 95588 113630
rect 96288 112930 96497 113630
rect 97197 112930 97406 113630
rect 98106 112930 98315 113630
rect 99015 112930 99224 113630
rect 99924 112930 100133 113630
rect 100833 112930 101042 113630
rect 101742 112930 101951 113630
rect 102651 112930 102860 113630
rect 103560 112930 103769 113630
rect 104469 112930 104678 113630
rect 105378 112930 105587 113630
rect 106287 112930 106496 113630
rect 107196 112930 107405 113630
rect 108105 112930 108314 113630
rect 109014 112930 109223 113630
rect 109923 112930 110132 113630
rect 110832 112930 111541 113630
rect 88384 112742 111541 112930
rect 88384 112042 89225 112742
rect 89925 112042 90134 112742
rect 90834 112042 91043 112742
rect 91743 112042 91952 112742
rect 92652 112042 92861 112742
rect 93561 112042 93770 112742
rect 94470 112042 94679 112742
rect 95379 112042 95588 112742
rect 96288 112042 96497 112742
rect 97197 112042 97406 112742
rect 98106 112042 98315 112742
rect 99015 112042 99224 112742
rect 99924 112042 100133 112742
rect 100833 112042 101042 112742
rect 101742 112042 101951 112742
rect 102651 112042 102860 112742
rect 103560 112042 103769 112742
rect 104469 112042 104678 112742
rect 105378 112042 105587 112742
rect 106287 112042 106496 112742
rect 107196 112042 107405 112742
rect 108105 112042 108314 112742
rect 109014 112042 109223 112742
rect 109923 112042 110132 112742
rect 110832 112042 111541 112742
rect 88384 111854 111541 112042
rect 88384 111154 89225 111854
rect 89925 111154 90134 111854
rect 90834 111154 91043 111854
rect 91743 111154 91952 111854
rect 92652 111154 92861 111854
rect 93561 111154 93770 111854
rect 94470 111154 94679 111854
rect 95379 111154 95588 111854
rect 96288 111154 96497 111854
rect 97197 111154 97406 111854
rect 98106 111154 98315 111854
rect 99015 111154 99224 111854
rect 99924 111154 100133 111854
rect 100833 111154 101042 111854
rect 101742 111154 101951 111854
rect 102651 111154 102860 111854
rect 103560 111154 103769 111854
rect 104469 111154 104678 111854
rect 105378 111154 105587 111854
rect 106287 111154 106496 111854
rect 107196 111154 107405 111854
rect 108105 111154 108314 111854
rect 109014 111154 109223 111854
rect 109923 111154 110132 111854
rect 110832 111154 111541 111854
rect 88384 110966 111541 111154
rect 88384 110266 89225 110966
rect 89925 110266 90134 110966
rect 90834 110266 91043 110966
rect 91743 110266 91952 110966
rect 92652 110266 92861 110966
rect 93561 110266 93770 110966
rect 94470 110266 94679 110966
rect 95379 110266 95588 110966
rect 96288 110266 96497 110966
rect 97197 110266 97406 110966
rect 98106 110266 98315 110966
rect 99015 110266 99224 110966
rect 99924 110266 100133 110966
rect 100833 110266 101042 110966
rect 101742 110266 101951 110966
rect 102651 110266 102860 110966
rect 103560 110266 103769 110966
rect 104469 110266 104678 110966
rect 105378 110266 105587 110966
rect 106287 110266 106496 110966
rect 107196 110266 107405 110966
rect 108105 110266 108314 110966
rect 109014 110266 109223 110966
rect 109923 110266 110132 110966
rect 110832 110266 111541 110966
rect 88384 110078 111541 110266
rect 88384 109378 89225 110078
rect 89925 109378 90134 110078
rect 90834 109378 91043 110078
rect 91743 109378 91952 110078
rect 92652 109378 92861 110078
rect 93561 109378 93770 110078
rect 94470 109378 94679 110078
rect 95379 109378 95588 110078
rect 96288 109378 96497 110078
rect 97197 109378 97406 110078
rect 98106 109378 98315 110078
rect 99015 109378 99224 110078
rect 99924 109378 100133 110078
rect 100833 109378 101042 110078
rect 101742 109378 101951 110078
rect 102651 109378 102860 110078
rect 103560 109378 103769 110078
rect 104469 109378 104678 110078
rect 105378 109378 105587 110078
rect 106287 109378 106496 110078
rect 107196 109378 107405 110078
rect 108105 109378 108314 110078
rect 109014 109378 109223 110078
rect 109923 109378 110132 110078
rect 110832 109378 111541 110078
rect 88384 109190 111541 109378
rect 88384 108490 89225 109190
rect 89925 108490 90134 109190
rect 90834 108490 91043 109190
rect 91743 108490 91952 109190
rect 92652 108490 92861 109190
rect 93561 108490 93770 109190
rect 94470 108490 94679 109190
rect 95379 108490 95588 109190
rect 96288 108490 96497 109190
rect 97197 108490 97406 109190
rect 98106 108490 98315 109190
rect 99015 108490 99224 109190
rect 99924 108490 100133 109190
rect 100833 108490 101042 109190
rect 101742 108490 101951 109190
rect 102651 108490 102860 109190
rect 103560 108490 103769 109190
rect 104469 108490 104678 109190
rect 105378 108490 105587 109190
rect 106287 108490 106496 109190
rect 107196 108490 107405 109190
rect 108105 108490 108314 109190
rect 109014 108490 109223 109190
rect 109923 108490 110132 109190
rect 110832 108490 111541 109190
rect 88384 108302 111541 108490
rect 88384 107602 89225 108302
rect 89925 107602 90134 108302
rect 90834 107602 91043 108302
rect 91743 107602 91952 108302
rect 92652 107602 92861 108302
rect 93561 107602 93770 108302
rect 94470 107602 94679 108302
rect 95379 107602 95588 108302
rect 96288 107602 96497 108302
rect 97197 107602 97406 108302
rect 98106 107602 98315 108302
rect 99015 107602 99224 108302
rect 99924 107602 100133 108302
rect 100833 107602 101042 108302
rect 101742 107602 101951 108302
rect 102651 107602 102860 108302
rect 103560 107602 103769 108302
rect 104469 107602 104678 108302
rect 105378 107602 105587 108302
rect 106287 107602 106496 108302
rect 107196 107602 107405 108302
rect 108105 107602 108314 108302
rect 109014 107602 109223 108302
rect 109923 107602 110132 108302
rect 110832 107602 111541 108302
rect 88384 107414 111541 107602
rect 88384 106714 89225 107414
rect 89925 106714 90134 107414
rect 90834 106714 91043 107414
rect 91743 106714 91952 107414
rect 92652 106714 92861 107414
rect 93561 106714 93770 107414
rect 94470 106714 94679 107414
rect 95379 106714 95588 107414
rect 96288 106714 96497 107414
rect 97197 106714 97406 107414
rect 98106 106714 98315 107414
rect 99015 106714 99224 107414
rect 99924 106714 100133 107414
rect 100833 106714 101042 107414
rect 101742 106714 101951 107414
rect 102651 106714 102860 107414
rect 103560 106714 103769 107414
rect 104469 106714 104678 107414
rect 105378 106714 105587 107414
rect 106287 106714 106496 107414
rect 107196 106714 107405 107414
rect 108105 106714 108314 107414
rect 109014 106714 109223 107414
rect 109923 106714 110132 107414
rect 110832 106714 111541 107414
rect 88384 106526 111541 106714
rect 88384 105826 89225 106526
rect 89925 105826 90134 106526
rect 90834 105826 91043 106526
rect 91743 105826 91952 106526
rect 92652 105826 92861 106526
rect 93561 105826 93770 106526
rect 94470 105826 94679 106526
rect 95379 105826 95588 106526
rect 96288 105826 96497 106526
rect 97197 105826 97406 106526
rect 98106 105826 98315 106526
rect 99015 105826 99224 106526
rect 99924 105826 100133 106526
rect 100833 105826 101042 106526
rect 101742 105826 101951 106526
rect 102651 105826 102860 106526
rect 103560 105826 103769 106526
rect 104469 105826 104678 106526
rect 105378 105826 105587 106526
rect 106287 105826 106496 106526
rect 107196 105826 107405 106526
rect 108105 105826 108314 106526
rect 109014 105826 109223 106526
rect 109923 105826 110132 106526
rect 110832 105826 111541 106526
rect 88384 105638 111541 105826
rect 88384 104938 89225 105638
rect 89925 104938 90134 105638
rect 90834 104938 91043 105638
rect 91743 104938 91952 105638
rect 92652 104938 92861 105638
rect 93561 104938 93770 105638
rect 94470 104938 94679 105638
rect 95379 104938 95588 105638
rect 96288 104938 96497 105638
rect 97197 104938 97406 105638
rect 98106 104938 98315 105638
rect 99015 104938 99224 105638
rect 99924 104938 100133 105638
rect 100833 104938 101042 105638
rect 101742 104938 101951 105638
rect 102651 104938 102860 105638
rect 103560 104938 103769 105638
rect 104469 104938 104678 105638
rect 105378 104938 105587 105638
rect 106287 104938 106496 105638
rect 107196 104938 107405 105638
rect 108105 104938 108314 105638
rect 109014 104938 109223 105638
rect 109923 104938 110132 105638
rect 110832 104938 111541 105638
rect 88384 104750 111541 104938
rect 88384 104050 89225 104750
rect 89925 104050 90134 104750
rect 90834 104050 91043 104750
rect 91743 104050 91952 104750
rect 92652 104050 92861 104750
rect 93561 104050 93770 104750
rect 94470 104050 94679 104750
rect 95379 104050 95588 104750
rect 96288 104050 96497 104750
rect 97197 104050 97406 104750
rect 98106 104050 98315 104750
rect 99015 104050 99224 104750
rect 99924 104050 100133 104750
rect 100833 104050 101042 104750
rect 101742 104050 101951 104750
rect 102651 104050 102860 104750
rect 103560 104050 103769 104750
rect 104469 104050 104678 104750
rect 105378 104050 105587 104750
rect 106287 104050 106496 104750
rect 107196 104050 107405 104750
rect 108105 104050 108314 104750
rect 109014 104050 109223 104750
rect 109923 104050 110132 104750
rect 110832 104050 111541 104750
rect 88384 103862 111541 104050
rect 88384 103162 89225 103862
rect 89925 103162 90134 103862
rect 90834 103162 91043 103862
rect 91743 103162 91952 103862
rect 92652 103162 92861 103862
rect 93561 103162 93770 103862
rect 94470 103162 94679 103862
rect 95379 103162 95588 103862
rect 96288 103162 96497 103862
rect 97197 103162 97406 103862
rect 98106 103162 98315 103862
rect 99015 103162 99224 103862
rect 99924 103162 100133 103862
rect 100833 103162 101042 103862
rect 101742 103162 101951 103862
rect 102651 103162 102860 103862
rect 103560 103162 103769 103862
rect 104469 103162 104678 103862
rect 105378 103162 105587 103862
rect 106287 103162 106496 103862
rect 107196 103162 107405 103862
rect 108105 103162 108314 103862
rect 109014 103162 109223 103862
rect 109923 103162 110132 103862
rect 110832 103162 111541 103862
rect 88384 102974 111541 103162
rect 88384 102274 89225 102974
rect 89925 102274 90134 102974
rect 90834 102274 91043 102974
rect 91743 102274 91952 102974
rect 92652 102274 92861 102974
rect 93561 102274 93770 102974
rect 94470 102274 94679 102974
rect 95379 102274 95588 102974
rect 96288 102274 96497 102974
rect 97197 102274 97406 102974
rect 98106 102274 98315 102974
rect 99015 102274 99224 102974
rect 99924 102274 100133 102974
rect 100833 102274 101042 102974
rect 101742 102274 101951 102974
rect 102651 102274 102860 102974
rect 103560 102274 103769 102974
rect 104469 102274 104678 102974
rect 105378 102274 105587 102974
rect 106287 102274 106496 102974
rect 107196 102274 107405 102974
rect 108105 102274 108314 102974
rect 109014 102274 109223 102974
rect 109923 102274 110132 102974
rect 110832 102274 111541 102974
rect 88384 102086 111541 102274
rect 88384 101386 89225 102086
rect 89925 101386 90134 102086
rect 90834 101386 91043 102086
rect 91743 101386 91952 102086
rect 92652 101386 92861 102086
rect 93561 101386 93770 102086
rect 94470 101386 94679 102086
rect 95379 101386 95588 102086
rect 96288 101386 96497 102086
rect 97197 101386 97406 102086
rect 98106 101386 98315 102086
rect 99015 101386 99224 102086
rect 99924 101386 100133 102086
rect 100833 101386 101042 102086
rect 101742 101386 101951 102086
rect 102651 101386 102860 102086
rect 103560 101386 103769 102086
rect 104469 101386 104678 102086
rect 105378 101386 105587 102086
rect 106287 101386 106496 102086
rect 107196 101386 107405 102086
rect 108105 101386 108314 102086
rect 109014 101386 109223 102086
rect 109923 101386 110132 102086
rect 110832 101386 111541 102086
rect 88384 101198 111541 101386
rect 88384 100498 89225 101198
rect 89925 100498 90134 101198
rect 90834 100498 91043 101198
rect 91743 100498 91952 101198
rect 92652 100498 92861 101198
rect 93561 100498 93770 101198
rect 94470 100498 94679 101198
rect 95379 100498 95588 101198
rect 96288 100498 96497 101198
rect 97197 100498 97406 101198
rect 98106 100498 98315 101198
rect 99015 100498 99224 101198
rect 99924 100498 100133 101198
rect 100833 100498 101042 101198
rect 101742 100498 101951 101198
rect 102651 100498 102860 101198
rect 103560 100498 103769 101198
rect 104469 100498 104678 101198
rect 105378 100498 105587 101198
rect 106287 100498 106496 101198
rect 107196 100498 107405 101198
rect 108105 100498 108314 101198
rect 109014 100498 109223 101198
rect 109923 100498 110132 101198
rect 110832 100498 111541 101198
rect 88384 100310 111541 100498
rect 88384 99610 89225 100310
rect 89925 99610 90134 100310
rect 90834 99610 91043 100310
rect 91743 99610 91952 100310
rect 92652 99610 92861 100310
rect 93561 99610 93770 100310
rect 94470 99610 94679 100310
rect 95379 99610 95588 100310
rect 96288 99610 96497 100310
rect 97197 99610 97406 100310
rect 98106 99610 98315 100310
rect 99015 99610 99224 100310
rect 99924 99610 100133 100310
rect 100833 99610 101042 100310
rect 101742 99610 101951 100310
rect 102651 99610 102860 100310
rect 103560 99610 103769 100310
rect 104469 99610 104678 100310
rect 105378 99610 105587 100310
rect 106287 99610 106496 100310
rect 107196 99610 107405 100310
rect 108105 99610 108314 100310
rect 109014 99610 109223 100310
rect 109923 99610 110132 100310
rect 110832 99610 111541 100310
rect 88384 99422 111541 99610
rect 481670 120220 508199 120671
rect 481670 119520 482072 120220
rect 482772 119520 483168 120220
rect 483868 119520 484264 120220
rect 484964 119520 485360 120220
rect 486060 119520 486456 120220
rect 487156 119520 487552 120220
rect 488252 119520 488648 120220
rect 489348 119520 489744 120220
rect 490444 119520 490840 120220
rect 491540 119520 491936 120220
rect 492636 119520 493032 120220
rect 493732 119520 494128 120220
rect 494828 119520 495224 120220
rect 495924 119520 496320 120220
rect 497020 119520 497416 120220
rect 498116 119520 498512 120220
rect 499212 119520 499608 120220
rect 500308 119520 500704 120220
rect 501404 119520 501800 120220
rect 502500 119520 502896 120220
rect 503596 119520 503992 120220
rect 504692 119520 505088 120220
rect 505788 119520 506184 120220
rect 506884 119520 507280 120220
rect 507980 119520 508199 120220
rect 481670 119069 508199 119520
rect 481670 118369 482072 119069
rect 482772 118369 483168 119069
rect 483868 118369 484264 119069
rect 484964 118369 485360 119069
rect 486060 118369 486456 119069
rect 487156 118369 487552 119069
rect 488252 118369 488648 119069
rect 489348 118369 489744 119069
rect 490444 118369 490840 119069
rect 491540 118369 491936 119069
rect 492636 118369 493032 119069
rect 493732 118369 494128 119069
rect 494828 118369 495224 119069
rect 495924 118369 496320 119069
rect 497020 118369 497416 119069
rect 498116 118369 498512 119069
rect 499212 118369 499608 119069
rect 500308 118369 500704 119069
rect 501404 118369 501800 119069
rect 502500 118369 502896 119069
rect 503596 118369 503992 119069
rect 504692 118369 505088 119069
rect 505788 118369 506184 119069
rect 506884 118369 507280 119069
rect 507980 118369 508199 119069
rect 481670 117918 508199 118369
rect 481670 117218 482072 117918
rect 482772 117218 483168 117918
rect 483868 117218 484264 117918
rect 484964 117218 485360 117918
rect 486060 117218 486456 117918
rect 487156 117218 487552 117918
rect 488252 117218 488648 117918
rect 489348 117218 489744 117918
rect 490444 117218 490840 117918
rect 491540 117218 491936 117918
rect 492636 117218 493032 117918
rect 493732 117218 494128 117918
rect 494828 117218 495224 117918
rect 495924 117218 496320 117918
rect 497020 117218 497416 117918
rect 498116 117218 498512 117918
rect 499212 117218 499608 117918
rect 500308 117218 500704 117918
rect 501404 117218 501800 117918
rect 502500 117218 502896 117918
rect 503596 117218 503992 117918
rect 504692 117218 505088 117918
rect 505788 117218 506184 117918
rect 506884 117218 507280 117918
rect 507980 117218 508199 117918
rect 481670 116767 508199 117218
rect 481670 116067 482072 116767
rect 482772 116067 483168 116767
rect 483868 116067 484264 116767
rect 484964 116067 485360 116767
rect 486060 116067 486456 116767
rect 487156 116067 487552 116767
rect 488252 116067 488648 116767
rect 489348 116067 489744 116767
rect 490444 116067 490840 116767
rect 491540 116067 491936 116767
rect 492636 116067 493032 116767
rect 493732 116067 494128 116767
rect 494828 116067 495224 116767
rect 495924 116067 496320 116767
rect 497020 116067 497416 116767
rect 498116 116067 498512 116767
rect 499212 116067 499608 116767
rect 500308 116067 500704 116767
rect 501404 116067 501800 116767
rect 502500 116067 502896 116767
rect 503596 116067 503992 116767
rect 504692 116067 505088 116767
rect 505788 116067 506184 116767
rect 506884 116067 507280 116767
rect 507980 116067 508199 116767
rect 481670 115616 508199 116067
rect 481670 114916 482072 115616
rect 482772 114916 483168 115616
rect 483868 114916 484264 115616
rect 484964 114916 485360 115616
rect 486060 114916 486456 115616
rect 487156 114916 487552 115616
rect 488252 114916 488648 115616
rect 489348 114916 489744 115616
rect 490444 114916 490840 115616
rect 491540 114916 491936 115616
rect 492636 114916 493032 115616
rect 493732 114916 494128 115616
rect 494828 114916 495224 115616
rect 495924 114916 496320 115616
rect 497020 114916 497416 115616
rect 498116 114916 498512 115616
rect 499212 114916 499608 115616
rect 500308 114916 500704 115616
rect 501404 114916 501800 115616
rect 502500 114916 502896 115616
rect 503596 114916 503992 115616
rect 504692 114916 505088 115616
rect 505788 114916 506184 115616
rect 506884 114916 507280 115616
rect 507980 114916 508199 115616
rect 481670 114465 508199 114916
rect 481670 113765 482072 114465
rect 482772 113765 483168 114465
rect 483868 113765 484264 114465
rect 484964 113765 485360 114465
rect 486060 113765 486456 114465
rect 487156 113765 487552 114465
rect 488252 113765 488648 114465
rect 489348 113765 489744 114465
rect 490444 113765 490840 114465
rect 491540 113765 491936 114465
rect 492636 113765 493032 114465
rect 493732 113765 494128 114465
rect 494828 113765 495224 114465
rect 495924 113765 496320 114465
rect 497020 113765 497416 114465
rect 498116 113765 498512 114465
rect 499212 113765 499608 114465
rect 500308 113765 500704 114465
rect 501404 113765 501800 114465
rect 502500 113765 502896 114465
rect 503596 113765 503992 114465
rect 504692 113765 505088 114465
rect 505788 113765 506184 114465
rect 506884 113765 507280 114465
rect 507980 113765 508199 114465
rect 481670 113314 508199 113765
rect 481670 112614 482072 113314
rect 482772 112614 483168 113314
rect 483868 112614 484264 113314
rect 484964 112614 485360 113314
rect 486060 112614 486456 113314
rect 487156 112614 487552 113314
rect 488252 112614 488648 113314
rect 489348 112614 489744 113314
rect 490444 112614 490840 113314
rect 491540 112614 491936 113314
rect 492636 112614 493032 113314
rect 493732 112614 494128 113314
rect 494828 112614 495224 113314
rect 495924 112614 496320 113314
rect 497020 112614 497416 113314
rect 498116 112614 498512 113314
rect 499212 112614 499608 113314
rect 500308 112614 500704 113314
rect 501404 112614 501800 113314
rect 502500 112614 502896 113314
rect 503596 112614 503992 113314
rect 504692 112614 505088 113314
rect 505788 112614 506184 113314
rect 506884 112614 507280 113314
rect 507980 112614 508199 113314
rect 481670 112163 508199 112614
rect 481670 111463 482072 112163
rect 482772 111463 483168 112163
rect 483868 111463 484264 112163
rect 484964 111463 485360 112163
rect 486060 111463 486456 112163
rect 487156 111463 487552 112163
rect 488252 111463 488648 112163
rect 489348 111463 489744 112163
rect 490444 111463 490840 112163
rect 491540 111463 491936 112163
rect 492636 111463 493032 112163
rect 493732 111463 494128 112163
rect 494828 111463 495224 112163
rect 495924 111463 496320 112163
rect 497020 111463 497416 112163
rect 498116 111463 498512 112163
rect 499212 111463 499608 112163
rect 500308 111463 500704 112163
rect 501404 111463 501800 112163
rect 502500 111463 502896 112163
rect 503596 111463 503992 112163
rect 504692 111463 505088 112163
rect 505788 111463 506184 112163
rect 506884 111463 507280 112163
rect 507980 111463 508199 112163
rect 481670 111012 508199 111463
rect 481670 110312 482072 111012
rect 482772 110312 483168 111012
rect 483868 110312 484264 111012
rect 484964 110312 485360 111012
rect 486060 110312 486456 111012
rect 487156 110312 487552 111012
rect 488252 110312 488648 111012
rect 489348 110312 489744 111012
rect 490444 110312 490840 111012
rect 491540 110312 491936 111012
rect 492636 110312 493032 111012
rect 493732 110312 494128 111012
rect 494828 110312 495224 111012
rect 495924 110312 496320 111012
rect 497020 110312 497416 111012
rect 498116 110312 498512 111012
rect 499212 110312 499608 111012
rect 500308 110312 500704 111012
rect 501404 110312 501800 111012
rect 502500 110312 502896 111012
rect 503596 110312 503992 111012
rect 504692 110312 505088 111012
rect 505788 110312 506184 111012
rect 506884 110312 507280 111012
rect 507980 110312 508199 111012
rect 481670 109861 508199 110312
rect 481670 109161 482072 109861
rect 482772 109161 483168 109861
rect 483868 109161 484264 109861
rect 484964 109161 485360 109861
rect 486060 109161 486456 109861
rect 487156 109161 487552 109861
rect 488252 109161 488648 109861
rect 489348 109161 489744 109861
rect 490444 109161 490840 109861
rect 491540 109161 491936 109861
rect 492636 109161 493032 109861
rect 493732 109161 494128 109861
rect 494828 109161 495224 109861
rect 495924 109161 496320 109861
rect 497020 109161 497416 109861
rect 498116 109161 498512 109861
rect 499212 109161 499608 109861
rect 500308 109161 500704 109861
rect 501404 109161 501800 109861
rect 502500 109161 502896 109861
rect 503596 109161 503992 109861
rect 504692 109161 505088 109861
rect 505788 109161 506184 109861
rect 506884 109161 507280 109861
rect 507980 109161 508199 109861
rect 481670 108710 508199 109161
rect 481670 108010 482072 108710
rect 482772 108010 483168 108710
rect 483868 108010 484264 108710
rect 484964 108010 485360 108710
rect 486060 108010 486456 108710
rect 487156 108010 487552 108710
rect 488252 108010 488648 108710
rect 489348 108010 489744 108710
rect 490444 108010 490840 108710
rect 491540 108010 491936 108710
rect 492636 108010 493032 108710
rect 493732 108010 494128 108710
rect 494828 108010 495224 108710
rect 495924 108010 496320 108710
rect 497020 108010 497416 108710
rect 498116 108010 498512 108710
rect 499212 108010 499608 108710
rect 500308 108010 500704 108710
rect 501404 108010 501800 108710
rect 502500 108010 502896 108710
rect 503596 108010 503992 108710
rect 504692 108010 505088 108710
rect 505788 108010 506184 108710
rect 506884 108010 507280 108710
rect 507980 108010 508199 108710
rect 481670 107559 508199 108010
rect 481670 106859 482072 107559
rect 482772 106859 483168 107559
rect 483868 106859 484264 107559
rect 484964 106859 485360 107559
rect 486060 106859 486456 107559
rect 487156 106859 487552 107559
rect 488252 106859 488648 107559
rect 489348 106859 489744 107559
rect 490444 106859 490840 107559
rect 491540 106859 491936 107559
rect 492636 106859 493032 107559
rect 493732 106859 494128 107559
rect 494828 106859 495224 107559
rect 495924 106859 496320 107559
rect 497020 106859 497416 107559
rect 498116 106859 498512 107559
rect 499212 106859 499608 107559
rect 500308 106859 500704 107559
rect 501404 106859 501800 107559
rect 502500 106859 502896 107559
rect 503596 106859 503992 107559
rect 504692 106859 505088 107559
rect 505788 106859 506184 107559
rect 506884 106859 507280 107559
rect 507980 106859 508199 107559
rect 481670 106408 508199 106859
rect 481670 105708 482072 106408
rect 482772 105708 483168 106408
rect 483868 105708 484264 106408
rect 484964 105708 485360 106408
rect 486060 105708 486456 106408
rect 487156 105708 487552 106408
rect 488252 105708 488648 106408
rect 489348 105708 489744 106408
rect 490444 105708 490840 106408
rect 491540 105708 491936 106408
rect 492636 105708 493032 106408
rect 493732 105708 494128 106408
rect 494828 105708 495224 106408
rect 495924 105708 496320 106408
rect 497020 105708 497416 106408
rect 498116 105708 498512 106408
rect 499212 105708 499608 106408
rect 500308 105708 500704 106408
rect 501404 105708 501800 106408
rect 502500 105708 502896 106408
rect 503596 105708 503992 106408
rect 504692 105708 505088 106408
rect 505788 105708 506184 106408
rect 506884 105708 507280 106408
rect 507980 105708 508199 106408
rect 481670 105257 508199 105708
rect 481670 104557 482072 105257
rect 482772 104557 483168 105257
rect 483868 104557 484264 105257
rect 484964 104557 485360 105257
rect 486060 104557 486456 105257
rect 487156 104557 487552 105257
rect 488252 104557 488648 105257
rect 489348 104557 489744 105257
rect 490444 104557 490840 105257
rect 491540 104557 491936 105257
rect 492636 104557 493032 105257
rect 493732 104557 494128 105257
rect 494828 104557 495224 105257
rect 495924 104557 496320 105257
rect 497020 104557 497416 105257
rect 498116 104557 498512 105257
rect 499212 104557 499608 105257
rect 500308 104557 500704 105257
rect 501404 104557 501800 105257
rect 502500 104557 502896 105257
rect 503596 104557 503992 105257
rect 504692 104557 505088 105257
rect 505788 104557 506184 105257
rect 506884 104557 507280 105257
rect 507980 104557 508199 105257
rect 481670 104106 508199 104557
rect 481670 103406 482072 104106
rect 482772 103406 483168 104106
rect 483868 103406 484264 104106
rect 484964 103406 485360 104106
rect 486060 103406 486456 104106
rect 487156 103406 487552 104106
rect 488252 103406 488648 104106
rect 489348 103406 489744 104106
rect 490444 103406 490840 104106
rect 491540 103406 491936 104106
rect 492636 103406 493032 104106
rect 493732 103406 494128 104106
rect 494828 103406 495224 104106
rect 495924 103406 496320 104106
rect 497020 103406 497416 104106
rect 498116 103406 498512 104106
rect 499212 103406 499608 104106
rect 500308 103406 500704 104106
rect 501404 103406 501800 104106
rect 502500 103406 502896 104106
rect 503596 103406 503992 104106
rect 504692 103406 505088 104106
rect 505788 103406 506184 104106
rect 506884 103406 507280 104106
rect 507980 103406 508199 104106
rect 481670 102955 508199 103406
rect 481670 102255 482072 102955
rect 482772 102255 483168 102955
rect 483868 102255 484264 102955
rect 484964 102255 485360 102955
rect 486060 102255 486456 102955
rect 487156 102255 487552 102955
rect 488252 102255 488648 102955
rect 489348 102255 489744 102955
rect 490444 102255 490840 102955
rect 491540 102255 491936 102955
rect 492636 102255 493032 102955
rect 493732 102255 494128 102955
rect 494828 102255 495224 102955
rect 495924 102255 496320 102955
rect 497020 102255 497416 102955
rect 498116 102255 498512 102955
rect 499212 102255 499608 102955
rect 500308 102255 500704 102955
rect 501404 102255 501800 102955
rect 502500 102255 502896 102955
rect 503596 102255 503992 102955
rect 504692 102255 505088 102955
rect 505788 102255 506184 102955
rect 506884 102255 507280 102955
rect 507980 102255 508199 102955
rect 481670 101804 508199 102255
rect 481670 101104 482072 101804
rect 482772 101104 483168 101804
rect 483868 101104 484264 101804
rect 484964 101104 485360 101804
rect 486060 101104 486456 101804
rect 487156 101104 487552 101804
rect 488252 101104 488648 101804
rect 489348 101104 489744 101804
rect 490444 101104 490840 101804
rect 491540 101104 491936 101804
rect 492636 101104 493032 101804
rect 493732 101104 494128 101804
rect 494828 101104 495224 101804
rect 495924 101104 496320 101804
rect 497020 101104 497416 101804
rect 498116 101104 498512 101804
rect 499212 101104 499608 101804
rect 500308 101104 500704 101804
rect 501404 101104 501800 101804
rect 502500 101104 502896 101804
rect 503596 101104 503992 101804
rect 504692 101104 505088 101804
rect 505788 101104 506184 101804
rect 506884 101104 507280 101804
rect 507980 101104 508199 101804
rect 481670 100653 508199 101104
rect 481670 99953 482072 100653
rect 482772 99953 483168 100653
rect 483868 99953 484264 100653
rect 484964 99953 485360 100653
rect 486060 99953 486456 100653
rect 487156 99953 487552 100653
rect 488252 99953 488648 100653
rect 489348 99953 489744 100653
rect 490444 99953 490840 100653
rect 491540 99953 491936 100653
rect 492636 99953 493032 100653
rect 493732 99953 494128 100653
rect 494828 99953 495224 100653
rect 495924 99953 496320 100653
rect 497020 99953 497416 100653
rect 498116 99953 498512 100653
rect 499212 99953 499608 100653
rect 500308 99953 500704 100653
rect 501404 99953 501800 100653
rect 502500 99953 502896 100653
rect 503596 99953 503992 100653
rect 504692 99953 505088 100653
rect 505788 99953 506184 100653
rect 506884 99953 507280 100653
rect 507980 99953 508199 100653
rect 481670 99723 508199 99953
rect 481670 99532 507195 99723
rect 88384 98722 89225 99422
rect 89925 98722 90134 99422
rect 90834 98722 91043 99422
rect 91743 98722 91952 99422
rect 92652 98722 92861 99422
rect 93561 98722 93770 99422
rect 94470 98722 94679 99422
rect 95379 98722 95588 99422
rect 96288 98722 96497 99422
rect 97197 98722 97406 99422
rect 98106 98722 98315 99422
rect 99015 98722 99224 99422
rect 99924 98722 100133 99422
rect 100833 98722 101042 99422
rect 101742 98722 101951 99422
rect 102651 98722 102860 99422
rect 103560 98722 103769 99422
rect 104469 98722 104678 99422
rect 105378 98722 105587 99422
rect 106287 98722 106496 99422
rect 107196 98722 107405 99422
rect 108105 98722 108314 99422
rect 109014 98722 109223 99422
rect 109923 98722 110132 99422
rect 110832 98722 111541 99422
rect 88384 98042 111541 98722
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_0
timestamp 1713338890
transform 0 1 4060 -1 0 115060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_1
timestamp 1713338890
transform 0 1 4060 -1 0 135060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_2
timestamp 1713338890
transform 1 0 100060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_3
timestamp 1713338890
transform 1 0 80060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_4
timestamp 1713338890
transform 1 0 120060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_5
timestamp 1713338890
transform 1 0 160060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_6
timestamp 1713338890
transform 0 -1 591060 1 0 160060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_7
timestamp 1713338890
transform 0 -1 591060 1 0 180060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_8
timestamp 1713338890
transform 0 -1 591060 1 0 480060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_9
timestamp 1713338890
transform -1 0 215060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_10
timestamp 1713338890
transform -1 0 235060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_11
timestamp 1713338890
transform -1 0 255060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_12
timestamp 1713338890
transform -1 0 275060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_13
timestamp 1713338890
transform -1 0 315060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_14
timestamp 1713338890
transform -1 0 335060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_15
timestamp 1713338890
transform -1 0 375060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_16
timestamp 1713338890
transform -1 0 395060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__asig_5p0  gf180mcu_fd_io__asig_5p0_17
timestamp 1713338890
transform -1 0 435060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_0
timestamp 1713338890
transform 0 1 4060 -1 0 195060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_1
timestamp 1713338890
transform 0 1 4060 -1 0 215060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_2
timestamp 1713338890
transform 0 1 4060 -1 0 235060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_3
timestamp 1713338890
transform 0 1 4060 -1 0 255060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_4
timestamp 1713338890
transform 0 1 4060 -1 0 295060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_5
timestamp 1713338890
transform 0 1 4060 -1 0 315060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_6
timestamp 1713338890
transform 0 1 4060 -1 0 335060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_7
timestamp 1713338890
transform 0 1 4060 -1 0 355060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_8
timestamp 1713338890
transform 0 1 4060 -1 0 395060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_9
timestamp 1713338890
transform 0 1 4060 -1 0 415060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_10
timestamp 1713338890
transform 0 1 4060 -1 0 435060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_11
timestamp 1713338890
transform 0 1 4060 -1 0 455060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_12
timestamp 1713338890
transform 0 1 4060 -1 0 495060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_13
timestamp 1713338890
transform 0 1 4060 -1 0 515060
box -32 0 15032 70000
use gf180mcu_fd_io__bi_t  gf180mcu_fd_io__bi_t_14
timestamp 1713338890
transform -1 0 95060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__brk5_vss_dvdd  gf180mcu_fd_io__brk5_vss_dvdd_0
timestamp 1713338890
transform -1 0 136060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__brk5_vss_dvss  gf180mcu_fd_io__brk5_vss_dvss_0
timestamp 1713338890
transform 1 0 199060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__brk5_vss_dvss  gf180mcu_fd_io__brk5_vss_dvss_1
timestamp 1713338890
transform 0 1 4060 -1 0 176060
box -32 13097 1032 69968
use gf180mcu_fd_io__brk5_vss_dvss  gf180mcu_fd_io__brk5_vss_dvss_2
timestamp 1713338890
transform 0 -1 591060 1 0 219060
box -32 13097 1032 69968
use gf180mcu_fd_io__brk5_vss_vdd  gf180mcu_fd_io__brk5_vss_vdd_0
timestamp 1713338890
transform -1 0 176060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__cor  gf180mcu_fd_io__cor_0
timestamp 1713338890
transform 1 0 4060 0 1 4060
box 13097 13097 71000 71000
use gf180mcu_fd_io__cor  gf180mcu_fd_io__cor_1
timestamp 1713338890
transform 0 -1 591060 1 0 4060
box 13097 13097 71000 71000
use gf180mcu_fd_io__cor  gf180mcu_fd_io__cor_2
timestamp 1713338890
transform 0 1 4060 -1 0 591060
box 13097 13097 71000 71000
use gf180mcu_fd_io__cor  gf180mcu_fd_io__cor_3
timestamp 1713338890
transform -1 0 591060 0 -1 591060
box 13097 13097 71000 71000
use gf180mcu_fd_io__dvdd  gf180mcu_fd_io__dvdd_0
timestamp 1713338890
transform 1 0 280060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  gf180mcu_fd_io__dvdd_1
timestamp 1713338890
transform 1 0 480060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  gf180mcu_fd_io__dvdd_2
timestamp 1713338890
transform 0 1 4060 -1 0 155060
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  gf180mcu_fd_io__dvdd_3
timestamp 1713338890
transform 0 1 4060 -1 0 275060
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  gf180mcu_fd_io__dvdd_4
timestamp 1713338890
transform 0 1 4060 -1 0 475060
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  gf180mcu_fd_io__dvdd_5
timestamp 1713338890
transform -1 0 135060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  gf180mcu_fd_io__dvdd_6
timestamp 1713338890
transform -1 0 195060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__dvdd  gf180mcu_fd_io__dvdd_7
timestamp 1713338890
transform -1 0 495060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_0
timestamp 1713338890
transform 0 1 4060 -1 0 95060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_1
timestamp 1713338890
transform 1 0 140060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_2
timestamp 1713338890
transform 1 0 180060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_3
timestamp 1713338890
transform 1 0 380060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_4
timestamp 1713338890
transform 0 1 4060 -1 0 175060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_5
timestamp 1713338890
transform 0 -1 591060 1 0 140060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_6
timestamp 1713338890
transform 0 -1 591060 1 0 200060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_7
timestamp 1713338890
transform 0 1 4060 -1 0 375060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_8
timestamp 1713338890
transform 0 -1 591060 1 0 460060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_9
timestamp 1713338890
transform 0 -1 591060 1 0 500060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_10
timestamp 1713338890
transform -1 0 115060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_11
timestamp 1713338890
transform -1 0 295060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_12
timestamp 1713338890
transform -1 0 355060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__dvss  gf180mcu_fd_io__dvss_13
timestamp 1713338890
transform -1 0 415060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_0
timestamp 1713338890
transform 1 0 99060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_1
timestamp 1713338890
transform 1 0 79060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_2
timestamp 1713338890
transform 0 1 4060 -1 0 76060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_3
timestamp 1713338890
transform 0 1 4060 -1 0 96060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_4
timestamp 1713338890
transform 0 1 4060 -1 0 116060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_5
timestamp 1713338890
transform 1 0 119060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_6
timestamp 1713338890
transform 1 0 139060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_7
timestamp 1713338890
transform 1 0 159060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_8
timestamp 1713338890
transform 1 0 179060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_9
timestamp 1713338890
transform 1 0 219060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_10
timestamp 1713338890
transform 1 0 239060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_11
timestamp 1713338890
transform 1 0 259060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_12
timestamp 1713338890
transform 1 0 279060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_13
timestamp 1713338890
transform 1 0 299060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_14
timestamp 1713338890
transform 1 0 319060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_15
timestamp 1713338890
transform 1 0 339060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_16
timestamp 1713338890
transform 1 0 359060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_17
timestamp 1713338890
transform 1 0 379060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_18
timestamp 1713338890
transform 1 0 399060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_19
timestamp 1713338890
transform 1 0 419060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_20
timestamp 1713338890
transform 1 0 479060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_21
timestamp 1713338890
transform 1 0 459060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_22
timestamp 1713338890
transform 1 0 439060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_23
timestamp 1713338890
transform 1 0 519060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_24
timestamp 1713338890
transform 1 0 499060 0 1 4060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_25
timestamp 1713338890
transform 0 -1 591060 1 0 79060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_26
timestamp 1713338890
transform 0 -1 591060 1 0 99060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_27
timestamp 1713338890
transform 0 -1 591060 1 0 119060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_28
timestamp 1713338890
transform 0 1 4060 -1 0 136060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_29
timestamp 1713338890
transform 0 1 4060 -1 0 156060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_30
timestamp 1713338890
transform 0 1 4060 -1 0 196060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_31
timestamp 1713338890
transform 0 1 4060 -1 0 216060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_32
timestamp 1713338890
transform 0 1 4060 -1 0 236060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_33
timestamp 1713338890
transform 0 1 4060 -1 0 256060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_34
timestamp 1713338890
transform 0 -1 591060 1 0 139060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_35
timestamp 1713338890
transform 0 -1 591060 1 0 159060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_36
timestamp 1713338890
transform 0 -1 591060 1 0 179060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_37
timestamp 1713338890
transform 0 -1 591060 1 0 199060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_38
timestamp 1713338890
transform 0 -1 591060 1 0 239060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_39
timestamp 1713338890
transform 0 1 4060 -1 0 276060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_40
timestamp 1713338890
transform 0 1 4060 -1 0 296060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_41
timestamp 1713338890
transform 0 1 4060 -1 0 316060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_42
timestamp 1713338890
transform 0 1 4060 -1 0 336060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_43
timestamp 1713338890
transform 0 1 4060 -1 0 356060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_44
timestamp 1713338890
transform 0 1 4060 -1 0 376060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_45
timestamp 1713338890
transform 0 -1 591060 1 0 259060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_46
timestamp 1713338890
transform 0 -1 591060 1 0 279060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_47
timestamp 1713338890
transform 0 -1 591060 1 0 299060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_48
timestamp 1713338890
transform 0 -1 591060 1 0 319060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_49
timestamp 1713338890
transform 0 -1 591060 1 0 339060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_50
timestamp 1713338890
transform 0 -1 591060 1 0 359060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_51
timestamp 1713338890
transform 0 -1 591060 1 0 379060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_52
timestamp 1713338890
transform 0 1 4060 -1 0 396060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_53
timestamp 1713338890
transform 0 1 4060 -1 0 416060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_54
timestamp 1713338890
transform 0 1 4060 -1 0 436060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_55
timestamp 1713338890
transform 0 1 4060 -1 0 456060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_56
timestamp 1713338890
transform 0 1 4060 -1 0 476060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_57
timestamp 1713338890
transform 0 1 4060 -1 0 496060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_58
timestamp 1713338890
transform 0 -1 591060 1 0 399060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_59
timestamp 1713338890
transform 0 -1 591060 1 0 419060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_60
timestamp 1713338890
transform 0 -1 591060 1 0 439060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_61
timestamp 1713338890
transform 0 -1 591060 1 0 459060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_62
timestamp 1713338890
transform 0 -1 591060 1 0 479060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_63
timestamp 1713338890
transform 0 -1 591060 1 0 499060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_64
timestamp 1713338890
transform -1 0 96060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_65
timestamp 1713338890
transform -1 0 76060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_66
timestamp 1713338890
transform 0 1 4060 -1 0 516060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_67
timestamp 1713338890
transform -1 0 116060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_68
timestamp 1713338890
transform -1 0 156060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_69
timestamp 1713338890
transform -1 0 196060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_70
timestamp 1713338890
transform -1 0 216060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_71
timestamp 1713338890
transform -1 0 236060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_72
timestamp 1713338890
transform -1 0 256060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_73
timestamp 1713338890
transform -1 0 276060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_74
timestamp 1713338890
transform -1 0 296060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_75
timestamp 1713338890
transform -1 0 316060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_76
timestamp 1713338890
transform -1 0 336060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_77
timestamp 1713338890
transform -1 0 356060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_78
timestamp 1713338890
transform -1 0 376060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_79
timestamp 1713338890
transform -1 0 396060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_80
timestamp 1713338890
transform -1 0 416060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_81
timestamp 1713338890
transform -1 0 436060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_82
timestamp 1713338890
transform -1 0 456060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_83
timestamp 1713338890
transform -1 0 476060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_84
timestamp 1713338890
transform -1 0 496060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_85
timestamp 1713338890
transform -1 0 516060 0 -1 591060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_86
timestamp 1713338890
transform 0 -1 591060 1 0 519060
box -32 13097 1032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_0
timestamp 1713338890
transform 1 0 95060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_1
timestamp 1713338890
transform 1 0 97060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_2
timestamp 1713338890
transform 1 0 77060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_3
timestamp 1713338890
transform 1 0 75060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_4
timestamp 1713338890
transform 0 1 4060 -1 0 78060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_5
timestamp 1713338890
transform 0 1 4060 -1 0 80060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_6
timestamp 1713338890
transform 0 1 4060 -1 0 98060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_7
timestamp 1713338890
transform 0 1 4060 -1 0 100060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_8
timestamp 1713338890
transform 0 1 4060 -1 0 120060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_9
timestamp 1713338890
transform 0 1 4060 -1 0 118060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_10
timestamp 1713338890
transform 1 0 117060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_11
timestamp 1713338890
transform 1 0 115060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_12
timestamp 1713338890
transform 1 0 137060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_13
timestamp 1713338890
transform 1 0 135060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_14
timestamp 1713338890
transform 1 0 155060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_15
timestamp 1713338890
transform 1 0 157060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_16
timestamp 1713338890
transform 1 0 177060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_17
timestamp 1713338890
transform 1 0 175060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_18
timestamp 1713338890
transform 1 0 195060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_19
timestamp 1713338890
transform 1 0 197060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_20
timestamp 1713338890
transform 1 0 215060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_21
timestamp 1713338890
transform 1 0 217060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_22
timestamp 1713338890
transform 1 0 235060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_23
timestamp 1713338890
transform 1 0 237060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_24
timestamp 1713338890
transform 1 0 255060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_25
timestamp 1713338890
transform 1 0 257060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_26
timestamp 1713338890
transform 1 0 275060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_27
timestamp 1713338890
transform 1 0 277060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_28
timestamp 1713338890
transform 1 0 295060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_29
timestamp 1713338890
transform 1 0 297060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_30
timestamp 1713338890
transform 1 0 315060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_31
timestamp 1713338890
transform 1 0 317060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_32
timestamp 1713338890
transform 1 0 335060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_33
timestamp 1713338890
transform 1 0 337060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_34
timestamp 1713338890
transform 1 0 355060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_35
timestamp 1713338890
transform 1 0 357060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_36
timestamp 1713338890
transform 1 0 375060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_37
timestamp 1713338890
transform 1 0 377060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_38
timestamp 1713338890
transform 1 0 395060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_39
timestamp 1713338890
transform 1 0 397060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_40
timestamp 1713338890
transform 1 0 415060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_41
timestamp 1713338890
transform 1 0 417060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_42
timestamp 1713338890
transform 1 0 477060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_43
timestamp 1713338890
transform 1 0 475060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_44
timestamp 1713338890
transform 1 0 457060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_45
timestamp 1713338890
transform 1 0 455060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_46
timestamp 1713338890
transform 1 0 437060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_47
timestamp 1713338890
transform 1 0 435060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_48
timestamp 1713338890
transform 1 0 515060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_49
timestamp 1713338890
transform 1 0 517060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_50
timestamp 1713338890
transform 1 0 497060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_51
timestamp 1713338890
transform 1 0 495060 0 1 4060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_52
timestamp 1713338890
transform 0 -1 591060 1 0 77060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_53
timestamp 1713338890
transform 0 -1 591060 1 0 75060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_54
timestamp 1713338890
transform 0 -1 591060 1 0 95060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_55
timestamp 1713338890
transform 0 -1 591060 1 0 97060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_56
timestamp 1713338890
transform 0 -1 591060 1 0 117060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_57
timestamp 1713338890
transform 0 -1 591060 1 0 115060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_58
timestamp 1713338890
transform 0 1 4060 -1 0 140060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_59
timestamp 1713338890
transform 0 1 4060 -1 0 138060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_60
timestamp 1713338890
transform 0 1 4060 -1 0 160060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_61
timestamp 1713338890
transform 0 1 4060 -1 0 158060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_62
timestamp 1713338890
transform 0 1 4060 -1 0 180060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_63
timestamp 1713338890
transform 0 1 4060 -1 0 178060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_64
timestamp 1713338890
transform 0 1 4060 -1 0 200060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_65
timestamp 1713338890
transform 0 1 4060 -1 0 198060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_66
timestamp 1713338890
transform 0 1 4060 -1 0 220060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_67
timestamp 1713338890
transform 0 1 4060 -1 0 218060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_68
timestamp 1713338890
transform 0 1 4060 -1 0 240060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_69
timestamp 1713338890
transform 0 1 4060 -1 0 238060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_70
timestamp 1713338890
transform 0 -1 591060 1 0 135060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_71
timestamp 1713338890
transform 0 -1 591060 1 0 137060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_72
timestamp 1713338890
transform 0 -1 591060 1 0 155060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_73
timestamp 1713338890
transform 0 -1 591060 1 0 157060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_74
timestamp 1713338890
transform 0 -1 591060 1 0 175060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_75
timestamp 1713338890
transform 0 -1 591060 1 0 177060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_76
timestamp 1713338890
transform 0 -1 591060 1 0 195060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_77
timestamp 1713338890
transform 0 -1 591060 1 0 197060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_78
timestamp 1713338890
transform 0 -1 591060 1 0 215060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_79
timestamp 1713338890
transform 0 -1 591060 1 0 217060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_80
timestamp 1713338890
transform 0 -1 591060 1 0 235060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_81
timestamp 1713338890
transform 0 -1 591060 1 0 237060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_82
timestamp 1713338890
transform 0 -1 591060 1 0 255060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_83
timestamp 1713338890
transform 0 1 4060 -1 0 260060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_84
timestamp 1713338890
transform 0 1 4060 -1 0 258060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_85
timestamp 1713338890
transform 0 1 4060 -1 0 280060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_86
timestamp 1713338890
transform 0 1 4060 -1 0 278060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_87
timestamp 1713338890
transform 0 1 4060 -1 0 300060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_88
timestamp 1713338890
transform 0 1 4060 -1 0 298060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_89
timestamp 1713338890
transform 0 1 4060 -1 0 320060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_90
timestamp 1713338890
transform 0 1 4060 -1 0 318060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_91
timestamp 1713338890
transform 0 1 4060 -1 0 340060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_92
timestamp 1713338890
transform 0 1 4060 -1 0 338060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_93
timestamp 1713338890
transform 0 1 4060 -1 0 358060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_94
timestamp 1713338890
transform 0 1 4060 -1 0 360060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_95
timestamp 1713338890
transform 0 1 4060 -1 0 378060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_96
timestamp 1713338890
transform 0 1 4060 -1 0 380060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_97
timestamp 1713338890
transform 0 -1 591060 1 0 257060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_98
timestamp 1713338890
transform 0 -1 591060 1 0 277060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_99
timestamp 1713338890
transform 0 -1 591060 1 0 275060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_100
timestamp 1713338890
transform 0 -1 591060 1 0 297060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_101
timestamp 1713338890
transform 0 -1 591060 1 0 295060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_102
timestamp 1713338890
transform 0 -1 591060 1 0 315060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_103
timestamp 1713338890
transform 0 -1 591060 1 0 317060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_104
timestamp 1713338890
transform 0 -1 591060 1 0 337060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_105
timestamp 1713338890
transform 0 -1 591060 1 0 335060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_106
timestamp 1713338890
transform 0 -1 591060 1 0 357060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_107
timestamp 1713338890
transform 0 -1 591060 1 0 355060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_108
timestamp 1713338890
transform 0 -1 591060 1 0 375060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_109
timestamp 1713338890
transform 0 -1 591060 1 0 377060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_110
timestamp 1713338890
transform 0 1 4060 -1 0 398060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_111
timestamp 1713338890
transform 0 1 4060 -1 0 400060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_112
timestamp 1713338890
transform 0 1 4060 -1 0 418060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_113
timestamp 1713338890
transform 0 1 4060 -1 0 420060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_114
timestamp 1713338890
transform 0 1 4060 -1 0 438060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_115
timestamp 1713338890
transform 0 1 4060 -1 0 440060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_116
timestamp 1713338890
transform 0 1 4060 -1 0 458060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_117
timestamp 1713338890
transform 0 1 4060 -1 0 460060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_118
timestamp 1713338890
transform 0 1 4060 -1 0 480060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_119
timestamp 1713338890
transform 0 1 4060 -1 0 478060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_120
timestamp 1713338890
transform 0 1 4060 -1 0 500060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_121
timestamp 1713338890
transform 0 1 4060 -1 0 498060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_122
timestamp 1713338890
transform 0 -1 591060 1 0 395060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_123
timestamp 1713338890
transform 0 -1 591060 1 0 397060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_124
timestamp 1713338890
transform 0 -1 591060 1 0 415060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_125
timestamp 1713338890
transform 0 -1 591060 1 0 417060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_126
timestamp 1713338890
transform 0 -1 591060 1 0 435060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_127
timestamp 1713338890
transform 0 -1 591060 1 0 437060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_128
timestamp 1713338890
transform 0 -1 591060 1 0 455060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_129
timestamp 1713338890
transform 0 -1 591060 1 0 457060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_130
timestamp 1713338890
transform 0 -1 591060 1 0 475060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_131
timestamp 1713338890
transform 0 -1 591060 1 0 477060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_132
timestamp 1713338890
transform 0 -1 591060 1 0 495060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_133
timestamp 1713338890
transform 0 -1 591060 1 0 497060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_134
timestamp 1713338890
transform -1 0 100060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_135
timestamp 1713338890
transform -1 0 98060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_136
timestamp 1713338890
transform -1 0 78060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_137
timestamp 1713338890
transform -1 0 80060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_138
timestamp 1713338890
transform 0 1 4060 -1 0 518060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_139
timestamp 1713338890
transform 0 1 4060 -1 0 520060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_140
timestamp 1713338890
transform -1 0 118060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_141
timestamp 1713338890
transform -1 0 120060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_142
timestamp 1713338890
transform -1 0 138060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_143
timestamp 1713338890
transform -1 0 140060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_144
timestamp 1713338890
transform -1 0 158060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_145
timestamp 1713338890
transform -1 0 160060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_146
timestamp 1713338890
transform -1 0 180060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_147
timestamp 1713338890
transform -1 0 178060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_148
timestamp 1713338890
transform -1 0 200060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_149
timestamp 1713338890
transform -1 0 198060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_150
timestamp 1713338890
transform -1 0 218060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_151
timestamp 1713338890
transform -1 0 220060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_152
timestamp 1713338890
transform -1 0 240060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_153
timestamp 1713338890
transform -1 0 238060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_154
timestamp 1713338890
transform -1 0 260060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_155
timestamp 1713338890
transform -1 0 258060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_156
timestamp 1713338890
transform -1 0 280060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_157
timestamp 1713338890
transform -1 0 278060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_158
timestamp 1713338890
transform -1 0 300060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_159
timestamp 1713338890
transform -1 0 298060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_160
timestamp 1713338890
transform -1 0 320060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_161
timestamp 1713338890
transform -1 0 318060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_162
timestamp 1713338890
transform -1 0 338060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_163
timestamp 1713338890
transform -1 0 340060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_164
timestamp 1713338890
transform -1 0 358060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_165
timestamp 1713338890
transform -1 0 360060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_166
timestamp 1713338890
transform -1 0 378060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_167
timestamp 1713338890
transform -1 0 380060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_168
timestamp 1713338890
transform -1 0 400060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_169
timestamp 1713338890
transform -1 0 398060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_170
timestamp 1713338890
transform -1 0 418060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_171
timestamp 1713338890
transform -1 0 420060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_172
timestamp 1713338890
transform -1 0 440060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_173
timestamp 1713338890
transform -1 0 438060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_174
timestamp 1713338890
transform -1 0 460060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_175
timestamp 1713338890
transform -1 0 458060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_176
timestamp 1713338890
transform -1 0 480060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_177
timestamp 1713338890
transform -1 0 478060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_178
timestamp 1713338890
transform -1 0 500060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_179
timestamp 1713338890
transform -1 0 498060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_180
timestamp 1713338890
transform -1 0 518060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_181
timestamp 1713338890
transform -1 0 520060 0 -1 591060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_182
timestamp 1713338890
transform 0 -1 591060 1 0 517060
box -32 13097 2032 69968
use gf180mcu_fd_io__fill10  gf180mcu_fd_io__fill10_183
timestamp 1713338890
transform 0 -1 591060 1 0 515060
box -32 13097 2032 69968
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_0
timestamp 1713338890
transform 1 0 200060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_1
timestamp 1713338890
transform 1 0 220060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_2
timestamp 1713338890
transform 1 0 240060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_3
timestamp 1713338890
transform 1 0 260060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_4
timestamp 1713338890
transform 1 0 300060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_5
timestamp 1713338890
transform 1 0 320060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_6
timestamp 1713338890
transform 1 0 340060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_7
timestamp 1713338890
transform 1 0 360060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_8
timestamp 1713338890
transform 1 0 400060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_9
timestamp 1713338890
transform 1 0 420060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_10
timestamp 1713338890
transform 0 -1 591060 1 0 80060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_11
timestamp 1713338890
transform 0 -1 591060 1 0 100060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_12
timestamp 1713338890
transform 0 -1 591060 1 0 120060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_13
timestamp 1713338890
transform 1 0 460060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_14
timestamp 1713338890
transform 1 0 440060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_15
timestamp 1713338890
transform 1 0 500060 0 1 4060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_16
timestamp 1713338890
transform -1 0 155060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_17
timestamp 1713338890
transform -1 0 175060 0 -1 591060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_18
timestamp 1713338890
transform 0 -1 591060 1 0 220060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_19
timestamp 1713338890
transform 0 -1 591060 1 0 240060
box -32 0 15032 70000
use gf180mcu_fd_io__in_c  gf180mcu_fd_io__in_c_20
timestamp 1713338890
transform 0 -1 591060 1 0 260060
box -32 0 15032 70000
use pad_fill_75  pad_fill_75_3
timestamp 1713338890
transform 0 -1 591060 1 0 280060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_4
timestamp 1713338890
transform 0 -1 591060 1 0 300060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_5
timestamp 1713338890
transform 0 -1 591060 1 0 320060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_6
timestamp 1713338890
transform 0 -1 591060 1 0 340060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_7
timestamp 1713338890
transform 0 -1 591060 1 0 360060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_8
timestamp 1713338890
transform 0 -1 591060 1 0 380060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_9
timestamp 1713338890
transform 0 -1 591060 1 0 400060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_10
timestamp 1713338890
transform 0 -1 591060 1 0 420060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_11
timestamp 1713338890
transform 0 -1 591060 1 0 440060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_12
timestamp 1713338890
transform -1 0 455060 0 -1 591060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_13
timestamp 1713338890
transform -1 0 475060 0 -1 591060
box -32 13097 15032 69968
use pad_fill_75  pad_fill_75_14
timestamp 1713338890
transform -1 0 515060 0 -1 591060
box -32 13097 15032 69968
<< end >>
