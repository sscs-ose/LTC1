magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect 285 -1968 12576 14320
<< psubdiff >>
rect 2285 12298 2621 12320
rect 2285 12252 2307 12298
rect 2353 12252 2421 12298
rect 2467 12252 2621 12298
rect 2285 12184 2621 12252
rect 2285 12138 2307 12184
rect 2353 12138 2421 12184
rect 2467 12138 2621 12184
rect 2285 12116 2621 12138
rect 10213 12116 10423 12320
rect 2285 12070 2489 12116
rect 2285 12024 2307 12070
rect 2353 12024 2421 12070
rect 2467 12024 2489 12070
rect 2285 11500 2489 12024
rect 2285 11454 2307 11500
rect 2353 11454 2421 11500
rect 2467 11454 2489 11500
rect 2285 11386 2489 11454
rect 2285 11340 2307 11386
rect 2353 11340 2421 11386
rect 2467 11340 2489 11386
rect 2285 11272 2489 11340
rect 2285 11226 2307 11272
rect 2353 11226 2421 11272
rect 2467 11226 2489 11272
rect 2285 11158 2489 11226
rect 2285 11112 2307 11158
rect 2353 11112 2421 11158
rect 2467 11112 2489 11158
rect 2285 11044 2489 11112
rect 2285 10998 2307 11044
rect 2353 10998 2421 11044
rect 2467 10998 2489 11044
rect 2285 10930 2489 10998
rect 2285 10884 2307 10930
rect 2353 10884 2421 10930
rect 2467 10884 2489 10930
rect 2285 10816 2489 10884
rect 2285 10770 2307 10816
rect 2353 10770 2421 10816
rect 2467 10770 2489 10816
rect 2285 10702 2489 10770
rect 2285 10656 2307 10702
rect 2353 10656 2421 10702
rect 2467 10656 2489 10702
rect 2285 10588 2489 10656
rect 2285 10542 2307 10588
rect 2353 10542 2421 10588
rect 2467 10542 2489 10588
rect 2285 10474 2489 10542
rect 2285 10428 2307 10474
rect 2353 10428 2421 10474
rect 2467 10428 2489 10474
rect 2285 10360 2489 10428
rect 2285 10314 2307 10360
rect 2353 10314 2421 10360
rect 2467 10314 2489 10360
rect 2285 10246 2489 10314
rect 2285 10200 2307 10246
rect 2353 10200 2421 10246
rect 2467 10200 2489 10246
rect 2285 10132 2489 10200
rect 2285 10086 2307 10132
rect 2353 10086 2421 10132
rect 2467 10086 2489 10132
rect 2285 10018 2489 10086
rect 2285 9972 2307 10018
rect 2353 9972 2421 10018
rect 2467 9972 2489 10018
rect 2285 9904 2489 9972
rect 2285 9858 2307 9904
rect 2353 9858 2421 9904
rect 2467 9858 2489 9904
rect 2285 9790 2489 9858
rect 2285 9744 2307 9790
rect 2353 9744 2421 9790
rect 2467 9744 2489 9790
rect 2285 9676 2489 9744
rect 2285 9630 2307 9676
rect 2353 9630 2421 9676
rect 2467 9630 2489 9676
rect 2285 9562 2489 9630
rect 2285 9516 2307 9562
rect 2353 9516 2421 9562
rect 2467 9516 2489 9562
rect 2285 9448 2489 9516
rect 2285 9402 2307 9448
rect 2353 9402 2421 9448
rect 2467 9402 2489 9448
rect 2285 9334 2489 9402
rect 2285 9288 2307 9334
rect 2353 9288 2421 9334
rect 2467 9288 2489 9334
rect 2285 9220 2489 9288
rect 2285 9174 2307 9220
rect 2353 9174 2421 9220
rect 2467 9174 2489 9220
rect 2285 9106 2489 9174
rect 2285 9060 2307 9106
rect 2353 9060 2421 9106
rect 2467 9060 2489 9106
rect 2285 8992 2489 9060
rect 2285 8946 2307 8992
rect 2353 8946 2421 8992
rect 2467 8946 2489 8992
rect 2285 8878 2489 8946
rect 2285 8832 2307 8878
rect 2353 8832 2421 8878
rect 2467 8832 2489 8878
rect 2285 8764 2489 8832
rect 2285 8718 2307 8764
rect 2353 8718 2421 8764
rect 2467 8718 2489 8764
rect 2285 8650 2489 8718
rect 2285 8604 2307 8650
rect 2353 8604 2421 8650
rect 2467 8604 2489 8650
rect 2285 8536 2489 8604
rect 2285 8490 2307 8536
rect 2353 8490 2421 8536
rect 2467 8490 2489 8536
rect 2285 8422 2489 8490
rect 2285 8376 2307 8422
rect 2353 8376 2421 8422
rect 2467 8376 2489 8422
rect 2285 8308 2489 8376
rect 2285 8262 2307 8308
rect 2353 8262 2421 8308
rect 2467 8262 2489 8308
rect 2285 8194 2489 8262
rect 2285 8148 2307 8194
rect 2353 8148 2421 8194
rect 2467 8148 2489 8194
rect 2285 8080 2489 8148
rect 2285 8034 2307 8080
rect 2353 8034 2421 8080
rect 2467 8034 2489 8080
rect 2285 7966 2489 8034
rect 2285 7920 2307 7966
rect 2353 7920 2421 7966
rect 2467 7920 2489 7966
rect 2285 7852 2489 7920
rect 2285 7806 2307 7852
rect 2353 7806 2421 7852
rect 2467 7806 2489 7852
rect 2285 7738 2489 7806
rect 2285 7692 2307 7738
rect 2353 7692 2421 7738
rect 2467 7692 2489 7738
rect 2285 7624 2489 7692
rect 2285 7578 2307 7624
rect 2353 7578 2421 7624
rect 2467 7578 2489 7624
rect 2285 7510 2489 7578
rect 2285 7464 2307 7510
rect 2353 7464 2421 7510
rect 2467 7464 2489 7510
rect 2285 7396 2489 7464
rect 2285 7350 2307 7396
rect 2353 7350 2421 7396
rect 2467 7350 2489 7396
rect 2285 7282 2489 7350
rect 2285 7236 2307 7282
rect 2353 7236 2421 7282
rect 2467 7236 2489 7282
rect 2285 7168 2489 7236
rect 2285 7122 2307 7168
rect 2353 7122 2421 7168
rect 2467 7122 2489 7168
rect 2285 7054 2489 7122
rect 2285 7008 2307 7054
rect 2353 7008 2421 7054
rect 2467 7008 2489 7054
rect 2285 6940 2489 7008
rect 2285 6894 2307 6940
rect 2353 6894 2421 6940
rect 2467 6894 2489 6940
rect 2285 6826 2489 6894
rect 2285 6780 2307 6826
rect 2353 6780 2421 6826
rect 2467 6780 2489 6826
rect 2285 6712 2489 6780
rect 2285 6666 2307 6712
rect 2353 6666 2421 6712
rect 2467 6666 2489 6712
rect 2285 6598 2489 6666
rect 2285 6552 2307 6598
rect 2353 6552 2421 6598
rect 2467 6552 2489 6598
rect 2285 6484 2489 6552
rect 2285 6438 2307 6484
rect 2353 6438 2421 6484
rect 2467 6438 2489 6484
rect 2285 6370 2489 6438
rect 2285 6324 2307 6370
rect 2353 6324 2421 6370
rect 2467 6324 2489 6370
rect 2285 6229 2489 6324
rect 2285 6025 2553 6229
rect 7260 32 10423 236
<< psubdiffcont >>
rect 2307 12252 2353 12298
rect 2421 12252 2467 12298
rect 2307 12138 2353 12184
rect 2421 12138 2467 12184
rect 2307 12024 2353 12070
rect 2421 12024 2467 12070
rect 2307 11454 2353 11500
rect 2421 11454 2467 11500
rect 2307 11340 2353 11386
rect 2421 11340 2467 11386
rect 2307 11226 2353 11272
rect 2421 11226 2467 11272
rect 2307 11112 2353 11158
rect 2421 11112 2467 11158
rect 2307 10998 2353 11044
rect 2421 10998 2467 11044
rect 2307 10884 2353 10930
rect 2421 10884 2467 10930
rect 2307 10770 2353 10816
rect 2421 10770 2467 10816
rect 2307 10656 2353 10702
rect 2421 10656 2467 10702
rect 2307 10542 2353 10588
rect 2421 10542 2467 10588
rect 2307 10428 2353 10474
rect 2421 10428 2467 10474
rect 2307 10314 2353 10360
rect 2421 10314 2467 10360
rect 2307 10200 2353 10246
rect 2421 10200 2467 10246
rect 2307 10086 2353 10132
rect 2421 10086 2467 10132
rect 2307 9972 2353 10018
rect 2421 9972 2467 10018
rect 2307 9858 2353 9904
rect 2421 9858 2467 9904
rect 2307 9744 2353 9790
rect 2421 9744 2467 9790
rect 2307 9630 2353 9676
rect 2421 9630 2467 9676
rect 2307 9516 2353 9562
rect 2421 9516 2467 9562
rect 2307 9402 2353 9448
rect 2421 9402 2467 9448
rect 2307 9288 2353 9334
rect 2421 9288 2467 9334
rect 2307 9174 2353 9220
rect 2421 9174 2467 9220
rect 2307 9060 2353 9106
rect 2421 9060 2467 9106
rect 2307 8946 2353 8992
rect 2421 8946 2467 8992
rect 2307 8832 2353 8878
rect 2421 8832 2467 8878
rect 2307 8718 2353 8764
rect 2421 8718 2467 8764
rect 2307 8604 2353 8650
rect 2421 8604 2467 8650
rect 2307 8490 2353 8536
rect 2421 8490 2467 8536
rect 2307 8376 2353 8422
rect 2421 8376 2467 8422
rect 2307 8262 2353 8308
rect 2421 8262 2467 8308
rect 2307 8148 2353 8194
rect 2421 8148 2467 8194
rect 2307 8034 2353 8080
rect 2421 8034 2467 8080
rect 2307 7920 2353 7966
rect 2421 7920 2467 7966
rect 2307 7806 2353 7852
rect 2421 7806 2467 7852
rect 2307 7692 2353 7738
rect 2421 7692 2467 7738
rect 2307 7578 2353 7624
rect 2421 7578 2467 7624
rect 2307 7464 2353 7510
rect 2421 7464 2467 7510
rect 2307 7350 2353 7396
rect 2421 7350 2467 7396
rect 2307 7236 2353 7282
rect 2421 7236 2467 7282
rect 2307 7122 2353 7168
rect 2421 7122 2467 7168
rect 2307 7008 2353 7054
rect 2421 7008 2467 7054
rect 2307 6894 2353 6940
rect 2421 6894 2467 6940
rect 2307 6780 2353 6826
rect 2421 6780 2467 6826
rect 2307 6666 2353 6712
rect 2421 6666 2467 6712
rect 2307 6552 2353 6598
rect 2421 6552 2467 6598
rect 2307 6438 2353 6484
rect 2421 6438 2467 6484
rect 2307 6324 2353 6370
rect 2421 6324 2467 6370
<< metal1 >>
rect 2296 12298 10565 12310
rect 2296 12252 2307 12298
rect 2353 12252 2421 12298
rect 2467 12252 10565 12298
rect 2296 12184 10565 12252
rect 2296 12138 2307 12184
rect 2353 12138 2421 12184
rect 2467 12138 10565 12184
rect 2296 12126 10565 12138
rect 2296 12070 2478 12126
rect 2296 12024 2307 12070
rect 2353 12024 2421 12070
rect 2467 12024 2478 12070
rect 2296 11633 2478 12024
rect 3125 11723 9913 11855
rect 3125 11655 5041 11723
rect 5561 11655 7477 11723
rect 7997 11655 9913 11723
rect 2296 11500 2914 11633
rect 2296 11454 2307 11500
rect 2353 11454 2421 11500
rect 2467 11454 2914 11500
rect 2296 11386 2914 11454
rect 2296 11340 2307 11386
rect 2353 11340 2421 11386
rect 2467 11340 2914 11386
rect 2296 11272 2914 11340
rect 2296 11226 2307 11272
rect 2353 11226 2421 11272
rect 2467 11226 2914 11272
rect 2296 11158 2914 11226
rect 2296 11112 2307 11158
rect 2353 11112 2421 11158
rect 2467 11112 2914 11158
rect 2296 11044 2914 11112
rect 2296 10998 2307 11044
rect 2353 10998 2421 11044
rect 2467 10998 2914 11044
rect 2296 10930 2914 10998
rect 2296 10884 2307 10930
rect 2353 10884 2421 10930
rect 2467 10884 2914 10930
rect 2296 10816 2914 10884
rect 2296 10770 2307 10816
rect 2353 10770 2421 10816
rect 2467 10770 2914 10816
rect 2296 10702 2914 10770
rect 2296 10656 2307 10702
rect 2353 10656 2421 10702
rect 2467 10656 2914 10702
rect 2296 10588 2914 10656
rect 2296 10542 2307 10588
rect 2353 10542 2421 10588
rect 2467 10542 2914 10588
rect 2296 10474 2914 10542
rect 2296 10428 2307 10474
rect 2353 10428 2421 10474
rect 2467 10428 2914 10474
rect 2296 10360 2914 10428
rect 2296 10314 2307 10360
rect 2353 10314 2421 10360
rect 2467 10314 2914 10360
rect 2296 10246 2914 10314
rect 2296 10200 2307 10246
rect 2353 10200 2421 10246
rect 2467 10200 2914 10246
rect 2296 10132 2914 10200
rect 2296 10086 2307 10132
rect 2353 10086 2421 10132
rect 2467 10086 2914 10132
rect 2296 10018 2914 10086
rect 2296 9972 2307 10018
rect 2353 9972 2421 10018
rect 2467 9972 2914 10018
rect 2296 9904 2914 9972
rect 2296 9858 2307 9904
rect 2353 9858 2421 9904
rect 2467 9858 2914 9904
rect 2296 9790 2914 9858
rect 2296 9744 2307 9790
rect 2353 9744 2421 9790
rect 2467 9744 2914 9790
rect 2296 9676 2914 9744
rect 2296 9630 2307 9676
rect 2353 9630 2421 9676
rect 2467 9630 2914 9676
rect 2296 9562 2914 9630
rect 2296 9516 2307 9562
rect 2353 9516 2421 9562
rect 2467 9516 2914 9562
rect 2296 9448 2914 9516
rect 2296 9402 2307 9448
rect 2353 9402 2421 9448
rect 2467 9402 2914 9448
rect 2296 9334 2914 9402
rect 2296 9288 2307 9334
rect 2353 9288 2421 9334
rect 2467 9288 2914 9334
rect 2296 9220 2914 9288
rect 2296 9174 2307 9220
rect 2353 9174 2421 9220
rect 2467 9174 2914 9220
rect 2296 9106 2914 9174
rect 2296 9060 2307 9106
rect 2353 9060 2421 9106
rect 2467 9060 2914 9106
rect 2296 8992 2914 9060
rect 2296 8946 2307 8992
rect 2353 8946 2421 8992
rect 2467 8946 2914 8992
rect 2296 8878 2914 8946
rect 2296 8832 2307 8878
rect 2353 8832 2421 8878
rect 2467 8832 2914 8878
rect 2296 8764 2914 8832
rect 2296 8718 2307 8764
rect 2353 8718 2421 8764
rect 2467 8718 2914 8764
rect 2296 8650 2914 8718
rect 2296 8604 2307 8650
rect 2353 8604 2421 8650
rect 2467 8604 2914 8650
rect 2296 8536 2914 8604
rect 2296 8490 2307 8536
rect 2353 8490 2421 8536
rect 2467 8490 2914 8536
rect 2296 8422 2914 8490
rect 2296 8376 2307 8422
rect 2353 8376 2421 8422
rect 2467 8376 2914 8422
rect 2296 8308 2914 8376
rect 2296 8262 2307 8308
rect 2353 8262 2421 8308
rect 2467 8262 2914 8308
rect 2296 8194 2914 8262
rect 2296 8148 2307 8194
rect 2353 8148 2421 8194
rect 2467 8148 2914 8194
rect 2296 8080 2914 8148
rect 2296 8034 2307 8080
rect 2353 8034 2421 8080
rect 2467 8034 2914 8080
rect 2296 7966 2914 8034
rect 2296 7920 2307 7966
rect 2353 7920 2421 7966
rect 2467 7920 2914 7966
rect 2296 7852 2914 7920
rect 2296 7806 2307 7852
rect 2353 7806 2421 7852
rect 2467 7806 2914 7852
rect 2296 7738 2914 7806
rect 2296 7692 2307 7738
rect 2353 7692 2421 7738
rect 2467 7692 2914 7738
rect 2296 7624 2914 7692
rect 2296 7578 2307 7624
rect 2353 7578 2421 7624
rect 2467 7578 2914 7624
rect 2296 7510 2914 7578
rect 2296 7464 2307 7510
rect 2353 7464 2421 7510
rect 2467 7464 2914 7510
rect 2296 7396 2914 7464
rect 2296 7350 2307 7396
rect 2353 7350 2421 7396
rect 2467 7350 2914 7396
rect 2296 7282 2914 7350
rect 2296 7236 2307 7282
rect 2353 7236 2421 7282
rect 2467 7236 2914 7282
rect 2296 7168 2914 7236
rect 2296 7122 2307 7168
rect 2353 7122 2421 7168
rect 2467 7122 2914 7168
rect 2296 7054 2914 7122
rect 2296 7008 2307 7054
rect 2353 7008 2421 7054
rect 2467 7008 2914 7054
rect 2296 6940 2914 7008
rect 2296 6894 2307 6940
rect 2353 6894 2421 6940
rect 2467 6894 2914 6940
rect 2296 6826 2914 6894
rect 2296 6780 2307 6826
rect 2353 6780 2421 6826
rect 2467 6780 2914 6826
rect 2296 6712 2914 6780
rect 2296 6666 2307 6712
rect 2353 6666 2421 6712
rect 2467 6666 2914 6712
rect 2296 6598 2914 6666
rect 2296 6552 2307 6598
rect 2353 6552 2421 6598
rect 2467 6552 2914 6598
rect 2296 6484 2914 6552
rect 2296 6438 2307 6484
rect 2353 6438 2421 6484
rect 2467 6483 2914 6484
rect 10173 6483 10383 11633
rect 2467 6438 10383 6483
rect 2296 6370 10383 6438
rect 2296 6324 2307 6370
rect 2353 6324 2421 6370
rect 2467 6324 10383 6370
rect 2296 5771 10383 6324
rect 7425 226 7743 5771
rect 10173 621 10383 5771
rect 7997 399 9913 599
rect 7271 42 10565 226
use M1_PSUB_CDNS_69033583165351  M1_PSUB_CDNS_69033583165351_0
timestamp 1713338890
transform 1 0 10474 0 1 6176
box -102 -6144 102 6144
use M1_PSUB_CDNS_69033583165480  M1_PSUB_CDNS_69033583165480_0
timestamp 1713338890
transform 0 -1 6417 1 0 12218
box -102 -3864 102 3864
use M1_PSUB_CDNS_69033583165481  M1_PSUB_CDNS_69033583165481_0
timestamp 1713338890
transform 0 -1 8946 1 0 134
box -102 -1356 102 1356
use M1_PSUB_CDNS_69033583165482  M1_PSUB_CDNS_69033583165482_0
timestamp 1713338890
transform 1 0 7367 0 1 3014
box -107 -2959 107 2959
use M1_PSUB_CDNS_69033583165483  M1_PSUB_CDNS_69033583165483_0
timestamp 1713338890
transform 0 -1 6439 1 0 6127
box -102 -3921 102 3921
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_0
timestamp 1713338890
transform 1 0 3083 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_1
timestamp 1713338890
transform 1 0 5519 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_2
timestamp 1713338890
transform 1 0 7955 0 1 6633
box -218 -350 2218 5092
use nmoscap_6p0_CDNS_406619531454  nmoscap_6p0_CDNS_406619531454_3
timestamp 1713338890
transform 1 0 7955 0 -1 5621
box -218 -350 2218 5092
<< labels >>
rlabel metal1 s 5302 6126 5302 6126 4 VMINUS
port 1 nsew
<< end >>
