magic
tech gf180mcuC
magscale 1 10
timestamp 1695206022
<< metal1 >>
rect 3441 11130 15727 11389
rect 3167 10828 3337 10885
rect 3167 10725 3209 10828
rect 3308 10725 3337 10828
rect 3167 10699 3337 10725
rect 16031 9653 16201 9722
rect 9465 9581 9726 9653
rect 15843 9581 16201 9653
rect 3334 9069 3556 9088
rect 3334 8950 3365 9069
rect 3527 8950 3556 9069
rect 3334 8919 3556 8950
rect 3268 8711 3883 8712
rect 3265 8654 3883 8711
rect 3265 6163 3337 8654
rect 7101 8106 7360 9145
rect 7828 8106 8087 9160
rect 8571 8106 8830 9176
rect 9668 8712 9726 9581
rect 16031 9534 16201 9581
rect 9668 8654 10254 8712
rect 12784 8106 13043 9210
rect 13591 8106 13850 9148
rect 14228 8106 14487 9171
rect 14958 8106 15217 9156
rect 3722 7847 15709 8106
rect 3794 6554 3987 7847
rect 4476 6554 4669 7847
rect 5101 6543 5294 7847
rect 5852 6554 6045 7847
rect 6671 6554 6864 7847
rect 7501 6577 7694 7847
rect 8240 6599 8433 7847
rect 9047 6577 9240 7847
rect 9946 6565 10139 7847
rect 15313 7053 15572 7122
rect 3265 6091 3505 6163
rect 3334 5879 3436 5894
rect 3334 5797 3344 5879
rect 3418 5797 3436 5879
rect 3334 5788 3436 5797
rect 3626 4330 15583 4614
<< via1 >>
rect 3209 10725 3308 10828
rect 3365 8950 3527 9069
rect 3344 5797 3418 5879
<< metal2 >>
rect 3167 10870 3337 10885
rect 3167 10710 3192 10870
rect 3323 10710 3337 10870
rect 3167 10699 3337 10710
rect 3334 9069 3556 9088
rect 3334 8950 3365 9069
rect 3527 9065 3556 9069
rect 3527 8963 3558 9065
rect 3527 8950 3556 8963
rect 3334 8919 3556 8950
rect 3334 5879 3436 8919
rect 3334 5797 3344 5879
rect 3418 5797 3436 5879
rect 3334 5788 3436 5797
<< via2 >>
rect 3192 10828 3323 10870
rect 3192 10725 3209 10828
rect 3209 10725 3308 10828
rect 3308 10725 3323 10828
rect 3192 10710 3323 10725
<< metal3 >>
rect 6461 10966 12885 11009
rect 6460 10909 12885 10966
rect 3167 10870 3337 10885
rect 3167 10710 3192 10870
rect 3323 10802 3337 10870
rect 3323 10725 6443 10802
rect 6461 10745 6518 10909
rect 12828 10745 12885 10909
rect 3323 10710 3337 10725
rect 3167 10699 3337 10710
rect 6366 5054 6443 10725
use CLK_div_3_mag  CLK_div_3_mag_0
timestamp 1695206022
transform -1 0 9601 0 -1 11239
box -34 -1 6461 3249
use CLK_div_3_mag  CLK_div_3_mag_1
timestamp 1695206022
transform -1 0 15970 0 -1 11239
box -34 -1 6461 3249
use CLK_div_10_mag  CLK_div_10_mag_0
timestamp 1695206022
transform 1 0 3386 0 1 4505
box -34 0 12197 3533
<< labels >>
flabel metal1 15535 7087 15535 7087 0 FreeSans 640 0 0 0 Vdiv90
port 0 nsew
flabel metal1 14713 7982 14713 7982 0 FreeSans 640 0 0 0 VDD
port 1 nsew
flabel metal1 12372 4448 12372 4448 0 FreeSans 640 0 0 0 VSS
port 2 nsew
flabel metal1 16073 9616 16073 9616 0 FreeSans 640 0 0 0 CLK
port 3 nsew
flabel via2 3249 10795 3249 10795 0 FreeSans 960 0 0 0 RST
port 4 nsew
<< end >>
