* NGSPICE file created from CLK_div_90_mag_flat.ext - technology: gf180mcuC

.subckt pex_CLK_div_90_mag VSS VDD RST Vdiv90 CLK
X0 a_4437_8231# CLK_div_3_mag_0.Q0.t3 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t54 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X1 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 a_12896_6955# VSS.t268 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_4898_4717# VSS.t43 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t223 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X4 a_4174_4717# CLK_div_10_mag_0.CLK a_4014_4717# VSS.t221 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X5 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.Q0.t3 VDD.t113 VDD.t112 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_10363_9798# VSS.t14 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X7 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VDD.t414 VDD.t413 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 a_11337_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t11 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X9 VDD CLK_div_3_mag_1.Q1.t3 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t456 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X10 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t61 VDD.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 VDD CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t46 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X12 VDD CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.CLK.t0 VDD.t440 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X13 a_11496_4761# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t62 VSS.t61 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X14 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t384 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X15 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t250 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X16 VDD CLK_div_3_mag_1.JK_FF_mag_1.K.t2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t374 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X17 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q2 a_12060_4761# VSS.t267 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X18 a_10363_9798# CLK_div_3_mag_1.JK_FF_mag_1.K.t3 CLK_div_3_mag_1.Q0.t1 VSS.t251 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X19 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_10209_10895# VSS.t293 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X20 VSS CLK_div_3_mag_1.Q1.t4 a_12215_9798# VSS.t296 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X21 VSS CLK.t0 a_11779_8699# VSS.t238 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X22 a_10960_6955# CLK_div_10_mag_0.Q1 VSS.t100 VSS.t99 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X23 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q1 VSS.t98 VSS.t97 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X24 VDD CLK_div_3_mag_0.Q0.t4 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t51 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X25 VDD CLK.t1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t362 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X26 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t11 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X27 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.and2_mag_1.OUT VDD.t184 VDD.t183 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X28 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_7761_5858# VSS.t125 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X29 a_5128_10895# RST.t0 a_4968_10895# VSS.t54 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X30 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1.t3 VDD.t412 VDD.t411 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t439 VDD.t438 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X32 a_12060_4761# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t70 VSS.t69 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X33 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t236 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 VSS CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.CLK.t1 VSS.t288 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X35 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK.t2 VDD.t366 VDD.t365 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X36 a_11779_8699# CLK_div_3_mag_1.Q1.t5 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t238 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X37 a_11906_5858# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t195 VSS.t194 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X38 VDD CLK.t3 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD.t367 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X39 a_7421_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t144 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X40 a_7761_5858# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t205 VSS.t204 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X41 a_11342_5858# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t208 VSS.t207 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X42 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK.t4 VDD.t371 VDD.t370 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X43 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t292 VSS.t291 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X44 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_8325_5858# VSS.t81 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X45 VDD RST.t1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t347 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X46 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.Q1.t6 VDD.t460 VDD.t459 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X47 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB VDD.t387 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X48 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t2 VDD.t351 VDD.t350 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X49 VDD CLK_div_3_mag_1.or_2_mag_0.IN2 a_10806_8231# VDD.t218 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X50 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.QB a_11906_5858# VSS.t270 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X51 a_7011_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1.t1 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X52 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VSS.t28 VSS.t27 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X53 VSS VDD.t469 a_12221_10895# VSS.t185 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X54 VSS CLK_div_3_mag_0.JK_FF_mag_1.K.t3 a_8863_9798# VSS.t84 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X55 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VDD.t119 VDD.t118 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X56 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_7575_9798# VSS.t45 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X57 VDD CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.Q1 VDD.t124 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X58 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4744_5858# VSS.t143 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X59 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t254 VDD.t253 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X60 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t400 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X61 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t308 VDD.t307 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X62 a_13949_4717# RST.t3 a_13789_4717# VSS.t232 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X63 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t134 VDD.t133 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X64 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K.t1 VDD.t289 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X65 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t182 VDD.t181 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t205 VDD.t204 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X67 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t298 VDD.t297 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X68 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_14514_10895# VSS.t209 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X69 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.CLK.t2 VDD.t136 VDD.t135 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X70 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_7011_9798# VSS.t45 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X71 a_8863_9798# CLK_div_3_mag_0.CLK.t3 a_8703_9798# VSS.t84 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X72 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t186 VDD.t185 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X73 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t41 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X74 a_7575_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X75 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t177 VDD.t176 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X76 a_7037_5814# CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VSS.t76 VSS.t75 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X77 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t309 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X78 a_14508_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t259 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X79 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t38 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X80 a_13789_4717# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t163 VSS.t162 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X81 VSS CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS.t72 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X82 a_4738_4717# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t197 VSS.t196 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X83 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB VDD.t35 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X84 a_15232_9798# CLK.t5 a_15072_9798# VSS.t241 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X85 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t427 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X86 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t79 VDD.t78 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X87 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_13949_4717# VSS.t131 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X88 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t286 VDD.t288 VDD.t287 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X89 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t59 VDD.t58 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X90 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t304 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X91 VDD CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_10_mag_0.CLK VDD.t55 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X92 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t178 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X93 a_13225_4717# CLK_div_10_mag_0.Q0 a_13065_4717# VSS.t26 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X94 VDD RST.t4 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t352 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X95 a_10209_10895# CLK_div_3_mag_1.Q0.t4 CLK_div_3_mag_1.JK_FF_mag_1.K VSS.t71 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X96 VDD VDD.t282 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t283 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X97 a_3994_9798# CLK_div_3_mag_0.JK_FF_mag_1.K.t4 CLK_div_3_mag_0.Q0.t2 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X98 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VDD.t34 VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X99 a_7197_5814# CLK_div_10_mag_0.Q0 a_7037_5814# VSS.t25 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X100 a_15078_10895# CLK_div_3_mag_1.Q1.t7 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t299 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X101 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.CLK VDD.t330 VDD.t329 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X102 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t65 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X103 a_10927_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t38 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X104 a_15072_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t30 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X105 VDD CLK_div_3_mag_0.Q1.t4 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t443 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X106 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t279 VDD.t281 VDD.t280 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X107 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VDD.t121 VDD.t120 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X108 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t195 VDD.t194 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X109 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.Q2 VDD.t399 VDD.t398 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X110 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t209 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X111 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB VDD.t84 VDD.t83 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X112 VDD CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.Q0 VDD.t80 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X113 a_13065_4717# VDD.t471 VSS.t184 VSS.t183 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X114 a_10932_4717# RST.t5 a_10772_4717# VSS.t233 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X115 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_8479_4761# VSS.t80 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X116 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t188 VDD.t187 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X117 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_13790_10895# VSS.t256 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X118 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_11491_9798# VSS.t159 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X119 a_12055_9798# CLK_div_3_mag_1.JK_FF_mag_1.K.t4 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t252 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X120 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t109 VDD.t108 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X121 a_9043_4761# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t104 VSS.t103 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X122 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t317 VDD.t316 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X123 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.Q0.t5 VSS.t73 VSS.t72 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X124 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t342 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X125 VDD VDD.t275 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t276 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X126 VSS CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_10_mag_0.CLK VSS.t34 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X127 a_5692_10895# CLK_div_3_mag_0.Q0.t5 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t33 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X128 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q0.t0 VDD.t212 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X129 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t334 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X130 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t426 VDD.t425 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X131 a_4020_5814# VDD.t473 VSS.t182 VSS.t181 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X132 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.K.t6 a_13231_5814# VSS.t77 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X133 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_10927_9798# VSS.t8 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X134 VSS CLK.t6 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t242 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X135 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t75 VDD.t74 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X136 VDD CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t326 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X137 a_10772_4717# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t115 VSS.t114 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X138 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_10_mag_0.Q2 a_10208_4717# VSS.t266 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X139 a_8479_4761# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t124 VSS.t123 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X140 a_6857_10895# CLK_div_3_mag_0.Q1.t5 CLK_div_3_mag_0.JK_FF_mag_1.QB VSS.t154 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X141 a_11491_9798# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t287 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X142 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.QB a_4180_5814# VSS.t50 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X143 a_7985_10895# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t148 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X144 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t408 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X145 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_10932_4717# VSS.t206 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X146 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.Q1 a_9043_4761# VSS.t96 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X147 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t466 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X148 a_12215_9798# CLK.t7 a_12055_9798# VSS.t245 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X149 VDD CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.IN2 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X150 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.Q1.t8 VDD.t462 VDD.t461 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X151 VSS CLK_div_3_mag_0.CLK.t4 a_5410_8699# VSS.t87 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X152 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 a_10960_6955# VSS.t265 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X153 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.QB a_8889_5858# VSS.t79 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X154 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t247 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X155 a_4180_5814# CLK_div_10_mag_0.CLK a_4020_5814# VSS.t220 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X156 a_12221_10895# CLK.t8 a_12061_10895# VSS.t246 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X157 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB VDD.t407 VDD.t406 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X158 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_14513_4761# VSS.t102 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X159 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5462_4761# VSS.t223 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X160 a_8889_5858# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t106 VSS.t105 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X161 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_13226_10895# VSS.t260 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X162 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0.t6 VDD.t50 VDD.t49 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X163 VDD CLK_div_3_mag_0.CLK.t5 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t137 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X164 a_14514_10895# RST.t6 a_14354_10895# VSS.t234 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X165 VDD CLK_div_3_mag_0.Q1.t6 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t299 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X166 VSS CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t2 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X167 a_8325_5858# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t48 VSS.t47 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X168 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_13795_5858# VSS.t109 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X169 Vdiv90 CLK_div_10_mag_0.Q3 VSS.t66 VSS.t65 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X170 a_5462_4761# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t142 VSS.t141 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X171 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB a_10214_5814# VSS.t269 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X172 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST.t7 VDD.t356 VDD.t355 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X173 VSS CLK.t9 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t247 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X174 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_3840_10895# VSS.t188 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X175 a_10806_8231# CLK_div_3_mag_1.Q0.t6 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD.t114 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X176 a_8869_10895# CLK_div_3_mag_0.CLK.t6 a_8709_10895# VSS.t90 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X177 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 VDD.t397 VDD.t396 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X178 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB a_5872_5858# VSS.t49 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X179 a_13795_5858# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t122 VSS.t121 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X180 a_4744_5858# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t68 VSS.t67 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X181 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_8145_10895# VSS.t201 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X182 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK.t10 VDD.t373 VDD.t372 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X183 VDD CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VDD.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X184 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8139_9798# VSS.t45 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X185 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t200 VSS.t199 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X186 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5308_5858# VSS.t222 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X187 a_10773_10895# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t37 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X188 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t206 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X189 a_8703_9798# CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t84 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X190 a_5872_5858# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t278 VSS.t277 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X191 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t165 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X192 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t96 VDD.t95 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X193 a_14964_7257# CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD.t346 VDD.t345 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X194 VSS CLK_div_10_mag_0.and2_mag_0.OUT Vdiv90.t2 VSS.t126 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X195 VSS VDD.t474 a_15238_10895# VSS.t178 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X196 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.CLK.t7 VDD.t141 VDD.t140 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X197 Vdiv90 CLK_div_10_mag_0.Q3 a_15124_7257# VDD.t104 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X198 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VSS.t24 VSS.t23 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X199 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t193 VDD.t192 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X200 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t73 VDD.t72 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X201 VDD CLK_div_3_mag_0.CLK.t8 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t142 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X202 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.CLK VSS.t219 VSS.t218 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X203 VSS CLK_div_3_mag_0.Q1.t7 a_5846_9798# VSS.t84 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X204 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t243 VDD.t242 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X205 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t230 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X206 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_4558_9798# VSS.t45 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X207 VDD RST.t8 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t357 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X208 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4404_10895# VSS.t227 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X209 VSS VDD.t475 a_5852_10895# VSS.t175 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X210 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t9 VDD.t361 VDD.t360 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X211 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X212 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t424 VDD.t423 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X213 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t101 VDD.t100 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X214 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_3994_9798# VSS.t45 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X215 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.CLK.t9 VDD.t146 VDD.t145 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X216 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t30 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X217 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t162 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X218 a_4558_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X219 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.QB VDD.t393 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X220 a_7915_4717# RST.t10 a_7755_4717# VSS.t235 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X221 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t17 VDD.t16 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X222 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_5122_9798# VSS.t45 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X223 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t77 VDD.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X224 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_11497_10895# VSS.t301 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X225 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t203 VDD.t202 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X226 VDD CLK_div_3_mag_0.JK_FF_mag_1.K.t5 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t415 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X227 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t71 VDD.t70 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X228 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t97 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X229 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.K VDD.t434 VDD.t433 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X230 a_13226_10895# CLK_div_3_mag_1.Q1.t9 CLK_div_3_mag_1.JK_FF_mag_1.QB VSS.t300 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X231 a_14354_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t158 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X232 VDD CLK_div_10_mag_0.JK_FF_mag_2.K.t7 CLK_div_10_mag_0.Q3 VDD.t430 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X233 a_10208_4717# CLK_div_10_mag_0.Q1 a_10048_4717# VSS.t95 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X234 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t111 VDD.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X235 a_13231_5814# CLK_div_10_mag_0.Q0 a_13071_5814# VSS.t22 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X236 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t337 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X237 VDD CLK_div_3_mag_0.CLK.t10 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t147 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X238 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t341 VDD.t340 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X239 a_11928_6955# CLK_div_10_mag_0.Q2 VSS.t264 VSS.t263 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X240 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_7915_4717# VSS.t46 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X241 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.and2_mag_1.OUT VSS.t111 VSS.t110 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X242 a_5410_8699# CLK_div_3_mag_0.Q1.t8 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t87 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X243 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X244 a_13071_5814# CLK_div_10_mag_0.JK_FF_mag_0.K VSS.t283 VSS.t282 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X245 a_3840_10895# CLK_div_3_mag_0.Q0.t7 CLK_div_3_mag_0.JK_FF_mag_1.K VSS.t32 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X246 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t239 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X247 VDD VDD.t271 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t272 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X248 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.Q1.t2 VDD.t189 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X249 a_6026_4761# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t83 VSS.t82 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X250 a_8709_10895# CLK_div_3_mag_0.Q1.t9 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t198 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X251 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t15 VDD.t14 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X252 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t62 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X253 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t159 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X254 a_14513_4761# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t108 VSS.t107 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X255 VDD CLK_div_3_mag_1.Q0.t7 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t115 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X256 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 a_11928_6955# VSS.t94 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X257 a_8145_10895# RST.t11 a_7985_10895# VSS.t236 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X258 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X259 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t435 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X260 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q1.t10 VDD.t422 VDD.t421 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X261 VDD CLK_div_3_mag_1.JK_FF_mag_1.K.t5 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t377 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X262 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.Q0 a_6026_4761# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X263 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t244 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X264 VDD CLK_div_3_mag_0.or_2_mag_0.IN2 a_4437_8231# VDD.t5 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X265 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t268 VDD.t270 VDD.t269 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X266 a_10214_5814# CLK_div_10_mag_0.Q1 a_10054_5814# VSS.t93 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X267 a_15238_10895# CLK.t11 a_15078_10895# VSS.t250 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X268 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_14359_5858# VSS.t101 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X269 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11496_4761# VSS.t40 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X270 a_14923_5858# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t276 VSS.t275 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X271 a_4968_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t132 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X272 a_10048_4717# VDD.t477 VSS.t174 VSS.t173 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X273 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.Q0.t0 VDD.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X274 a_4404_10895# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t44 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X275 a_5852_10895# CLK_div_3_mag_0.CLK.t11 a_5692_10895# VSS.t91 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X276 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X277 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q0 VDD.t29 VDD.t28 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X278 a_14359_5858# CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t130 VSS.t129 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X279 a_8139_9798# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X280 VSS CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t5 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X281 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t113 VSS.t112 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X282 a_5308_5858# CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t42 VSS.t41 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X283 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_10778_5858# VSS.t60 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X284 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_6857_10895# VSS.t145 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X285 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_2.K.t8 a_14923_5858# VSS.t281 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X286 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K.t1 VDD.t453 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X287 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VDD.t381 VDD.t380 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X288 a_15124_7257# CLK_div_10_mag_0.and2_mag_0.OUT a_14964_7257# VDD.t201 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X289 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.Q1 VDD.t153 VDD.t152 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X290 a_11497_10895# RST.t12 a_11337_10895# VSS.t237 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X291 VDD CLK_div_3_mag_1.Q1.t10 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t463 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X292 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t59 VSS.t58 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X293 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t265 VDD.t267 VDD.t266 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X294 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t130 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X295 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t262 VDD.t264 VDD.t263 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X296 a_5846_9798# CLK_div_3_mag_0.CLK.t12 a_5686_9798# VSS.t84 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X297 VDD CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t390 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X298 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t175 VDD.t174 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X299 a_10778_5858# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X300 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t447 VDD.t446 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X301 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t94 VDD.t93 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X302 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.Q1 VDD.t158 VDD.t157 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X303 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST.t13 VDD.t89 VDD.t88 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X304 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11342_5858# VSS.t39 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X305 a_13790_10895# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t13 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X306 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t200 VDD.t199 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X307 a_5686_9798# CLK_div_3_mag_0.JK_FF_mag_1.K.t6 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t84 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X308 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0.t8 VSS.t31 VSS.t5 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X309 a_10054_5814# VDD.t478 VSS.t172 VSS.t171 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X310 a_7031_4717# VDD.t479 VSS.t170 VSS.t169 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X311 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t229 VDD.t228 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X312 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_10_mag_0.Q1 a_7191_4717# VSS.t92 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X313 VDD CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.QB VDD.t154 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X314 VDD CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t25 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X315 a_7755_4717# CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t57 VSS.t56 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X316 VSS CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_5128_10895# VSS.t224 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X317 a_5122_9798# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X318 VSS CLK_div_3_mag_0.CLK.t13 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t212 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X319 VDD CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.IN2 VDD.t292 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X320 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q1 VDD.t151 VDD.t150 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X321 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t196 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X322 VSS CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_7421_10895# VSS.t151 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X323 VSS VDD.t480 a_8869_10895# VSS.t166 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X324 a_7191_4717# CLK_div_10_mag_0.Q0 a_7031_4717# VSS.t20 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X325 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t168 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X326 VDD RST.t14 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X327 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_13380_9798# VSS.t116 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X328 a_13944_9798# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t12 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X329 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.Q0 VDD.t24 VDD.t23 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X330 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t259 VDD.t261 VDD.t260 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X331 VDD VDD.t255 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t256 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X332 VDD CLK_div_3_mag_0.JK_FF_mag_1.K.t7 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t418 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X333 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_0.Q3 VDD.t103 VDD.t102 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X334 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t331 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X335 a_12061_10895# CLK_div_3_mag_1.Q0.t8 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t74 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X336 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t233 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X337 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t296 VDD.t295 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X338 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.Q0 VDD.t22 VDD.t21 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X339 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_14508_9798# VSS.t51 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X340 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.QB VDD.t123 VDD.t122 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X341 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t313 VDD.t312 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X342 a_13380_9798# CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.Q1.t1 VSS.t29 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X343 VSS CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.IN2 VSS.t191 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X344 a_12896_6955# CLK_div_10_mag_0.Q0 VSS.t19 VSS.t18 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X345 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.Q3 a_15077_4761# VSS.t64 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X346 a_4898_4717# RST.t15 a_4738_4717# VSS.t55 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X347 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_10773_10895# VSS.t284 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X348 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t318 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X349 VSS CLK_div_3_mag_1.JK_FF_mag_1.K.t7 a_15232_9798# VSS.t253 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X350 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t127 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X351 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t315 VDD.t314 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X352 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t69 VDD.t68 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X353 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1.t0 VDD.t215 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X354 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.CLK.t14 VDD.t322 VDD.t321 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X355 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_10_mag_0.Q3 a_13225_4717# VSS.t63 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X356 a_4014_4717# VDD.t482 VSS.t165 VSS.t164 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X357 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t222 VDD.t221 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X358 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_13944_9798# VSS.t155 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X359 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t227 VDD.t226 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X360 VDD CLK.t12 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t448 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X361 VDD CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t323 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X362 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t383 VDD.t382 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X363 VDD CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.Q2 VDD.t403 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X364 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.QB a_7197_5814# VSS.t78 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X365 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_10_mag_0.Q0 a_4174_4717# VSS.t17 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X366 VSS CLK_div_3_mag_0.CLK.t15 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t215 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X367 a_15077_4761# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t120 VSS.t119 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X368 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK.t13 VDD.t452 VDD.t451 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X369 Vdiv90 CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS.t231 VSS.t230 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
R0 CLK_div_3_mag_0.Q0.n2 CLK_div_3_mag_0.Q0.t5 36.935
R1 CLK_div_3_mag_0.Q0.n3 CLK_div_3_mag_0.Q0.t7 31.4332
R2 CLK_div_3_mag_0.Q0.n5 CLK_div_3_mag_0.Q0.t3 29.8135
R3 CLK_div_3_mag_0.Q0.n5 CLK_div_3_mag_0.Q0.t8 27.8352
R4 CLK_div_3_mag_0.Q0.n2 CLK_div_3_mag_0.Q0.t4 18.1962
R5 CLK_div_3_mag_0.Q0.n3 CLK_div_3_mag_0.Q0.t6 15.3826
R6 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.t2 7.09905
R7 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n3 6.86029
R8 CLK_div_3_mag_0.Q0.n4 CLK_div_3_mag_0.Q0 5.01077
R9 CLK_div_3_mag_0.Q0.n6 CLK_div_3_mag_0.Q0 3.41843
R10 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n1 3.25053
R11 CLK_div_3_mag_0.Q0.n1 CLK_div_3_mag_0.Q0.t0 2.2755
R12 CLK_div_3_mag_0.Q0.n1 CLK_div_3_mag_0.Q0.n0 2.2755
R13 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n6 2.2505
R14 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n2 2.13459
R15 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q0.n5 1.74998
R16 CLK_div_3_mag_0.Q0.n6 CLK_div_3_mag_0.Q0.n4 1.50381
R17 CLK_div_3_mag_0.Q0.n4 CLK_div_3_mag_0.Q0 1.12067
R18 VDD.n160 VDD.n12 11185.2
R19 VDD.n200 VDD.n193 11185.2
R20 VDD.n233 VDD.n225 11185.2
R21 VDD.n140 VDD.t185 1105.93
R22 VDD.t62 VDD.t295 961.905
R23 VDD.t406 VDD.t0 961.905
R24 VDD.t127 VDD.t176 961.905
R25 VDD.t122 VDD.t312 961.905
R26 VDD.t425 VDD.t334 961.905
R27 VDD.t108 VDD.t83 961.905
R28 VDD.t318 VDD.t456 765.152
R29 VDD.t247 VDD.t384 765.152
R30 VDD.t387 VDD.t16 765.152
R31 VDD.t46 VDD.t85 765.152
R32 VDD.t244 VDD.t382 765.152
R33 VDD.t189 VDD.t14 765.152
R34 VDD.t374 VDD.t250 765.152
R35 VDD.t11 VDD.t438 765.152
R36 VDD.t18 VDD.t60 765.152
R37 VDD.t466 VDD.t115 765.152
R38 VDD.t8 VDD.t435 765.152
R39 VDD.t453 VDD.t58 765.152
R40 VDD.t130 VDD.t174 765.152
R41 VDD.t76 VDD.t199 765.152
R42 VDD.t157 VDD.t93 765.152
R43 VDD.t427 VDD.t304 765.152
R44 VDD.t242 VDD.t233 765.152
R45 VDD.t215 VDD.t226 765.152
R46 VDD.t309 VDD.t299 765.152
R47 VDD.t236 VDD.t239 765.152
R48 VDD.t230 VDD.t228 765.152
R49 VDD.t415 VDD.t408 765.152
R50 VDD.t209 VDD.t340 765.152
R51 VDD.t212 VDD.t74 765.152
R52 VDD.t337 VDD.t51 765.152
R53 VDD.t206 VDD.t342 765.152
R54 VDD.t289 VDD.t72 765.152
R55 VDD.t331 VDD.t133 765.152
R56 VDD.t68 VDD.t221 765.152
R57 VDD.t21 VDD.t297 765.152
R58 VDD.t423 VDD.t171 765.152
R59 VDD.t178 VDD.t202 765.152
R60 VDD.t194 VDD.t120 765.152
R61 VDD.t168 VDD.t192 765.152
R62 VDD.t204 VDD.t181 765.152
R63 VDD.t102 VDD.t253 765.152
R64 VDD.t65 VDD.t110 765.152
R65 VDD.t316 VDD.t100 765.152
R66 VDD.t398 VDD.t187 765.152
R67 VDD.n136 VDD.t345 747.159
R68 VDD.t314 VDD.n12 676.191
R69 VDD.n193 VDD.t78 676.191
R70 VDD.n225 VDD.t70 676.191
R71 VDD.t446 VDD.t183 645.307
R72 VDD.n160 VDD.t266 485.714
R73 VDD.n200 VDD.t118 485.714
R74 VDD.t280 VDD.n233 485.714
R75 VDD VDD.n93 429.187
R76 VDD.n151 VDD 427.092
R77 VDD.n146 VDD 427.092
R78 VDD.n439 VDD 426.699
R79 VDD VDD.n504 426.699
R80 VDD VDD.n285 426.699
R81 VDD.n307 VDD 426.699
R82 VDD.t152 VDD.n160 426.44
R83 VDD.t23 VDD.n200 426.44
R84 VDD.n233 VDD.t329 426.44
R85 VDD.n141 VDD 425.019
R86 VDD.n393 VDD 424.618
R87 VDD.n228 VDD 424.618
R88 VDD VDD.n395 418.495
R89 VDD VDD.n208 418.495
R90 VDD.n146 VDD.t28 386.365
R91 VDD.n151 VDD.t396 386.365
R92 VDD.t377 VDD.n439 386.365
R93 VDD.n504 VDD.t463 386.365
R94 VDD.n285 VDD.t418 386.365
R95 VDD.t443 VDD.n307 386.365
R96 VDD.n93 VDD.t433 386.365
R97 VDD.t159 VDD.t406 380.952
R98 VDD.t38 VDD.t122 380.952
R99 VDD.t83 VDD.t326 380.952
R100 VDD.t390 VDD.n141 378.788
R101 VDD.t165 VDD.n146 378.788
R102 VDD.t400 VDD.n151 378.788
R103 VDD.n395 VDD.t459 378.788
R104 VDD.n208 VDD.t421 378.788
R105 VDD.n395 VDD.t218 322.223
R106 VDD.t5 VDD.n208 322.223
R107 VDD.t114 VDD.n393 320.635
R108 VDD.t54 VDD.n228 320.635
R109 VDD.t456 VDD.t372 303.031
R110 VDD.t350 VDD.t247 303.031
R111 VDD.t451 VDD.t46 303.031
R112 VDD.t365 VDD.t374 303.031
R113 VDD.t115 VDD.t370 303.031
R114 VDD.t360 VDD.t8 303.031
R115 VDD.t357 VDD.t76 303.031
R116 VDD.t25 VDD.t157 303.031
R117 VDD.t304 VDD.t321 303.031
R118 VDD.t299 VDD.t135 303.031
R119 VDD.t355 VDD.t236 303.031
R120 VDD.t145 VDD.t415 303.031
R121 VDD.t51 VDD.t140 303.031
R122 VDD.t88 VDD.t206 303.031
R123 VDD.t90 VDD.t68 303.031
R124 VDD.t323 VDD.t21 303.031
R125 VDD.t120 VDD.t30 303.031
R126 VDD.t347 VDD.t204 303.031
R127 VDD.t41 VDD.t102 303.031
R128 VDD.t352 VDD.t316 303.031
R129 VDD.t162 VDD.t398 303.031
R130 VDD.t97 VDD.n12 285.714
R131 VDD.n193 VDD.t196 285.714
R132 VDD.n225 VDD.t223 285.714
R133 VDD.n120 VDD.t403 242.857
R134 VDD.n121 VDD.t62 242.857
R135 VDD.n158 VDD.t97 242.857
R136 VDD.n159 VDD.t159 242.857
R137 VDD.n161 VDD.t124 242.857
R138 VDD.n163 VDD.t127 242.857
R139 VDD.t196 VDD.n166 242.857
R140 VDD.n199 VDD.t38 242.857
R141 VDD.n219 VDD.t80 242.857
R142 VDD.n224 VDD.t334 242.857
R143 VDD.n235 VDD.t223 242.857
R144 VDD.t326 VDD.n234 242.857
R145 VDD.n142 VDD.t390 193.183
R146 VDD.n147 VDD.t165 193.183
R147 VDD.n152 VDD.t400 193.183
R148 VDD.n366 VDD.t154 193.183
R149 VDD.n368 VDD.t130 193.183
R150 VDD.n371 VDD.t357 193.183
R151 VDD.n374 VDD.t25 193.183
R152 VDD.n173 VDD.t35 193.183
R153 VDD.n175 VDD.t331 193.183
R154 VDD.n178 VDD.t90 193.183
R155 VDD.n181 VDD.t323 193.183
R156 VDD.n80 VDD.t430 193.183
R157 VDD.n86 VDD.t171 193.183
R158 VDD.n87 VDD.t178 193.183
R159 VDD.n92 VDD.t30 193.183
R160 VDD.n25 VDD.t105 193.183
R161 VDD.n27 VDD.t168 193.183
R162 VDD.n30 VDD.t347 193.183
R163 VDD.n33 VDD.t41 193.183
R164 VDD.n96 VDD.t393 193.183
R165 VDD.n98 VDD.t65 193.183
R166 VDD.n101 VDD.t352 193.183
R167 VDD.n104 VDD.t162 193.183
R168 VDD.t459 VDD.n4 191.288
R169 VDD.t372 VDD.n420 191.288
R170 VDD.n421 VDD.t350 191.288
R171 VDD.t16 VDD.n429 191.288
R172 VDD.n430 VDD.t461 191.288
R173 VDD.n440 VDD.t451 191.288
R174 VDD.t382 VDD.n447 191.288
R175 VDD.t14 VDD.n452 191.288
R176 VDD.n453 VDD.t44 191.288
R177 VDD.n503 VDD.t365 191.288
R178 VDD.n502 VDD.t438 191.288
R179 VDD.t60 VDD.n468 191.288
R180 VDD.n470 VDD.t380 191.288
R181 VDD.t370 VDD.n481 191.288
R182 VDD.n482 VDD.t360 191.288
R183 VDD.t58 VDD.n490 191.288
R184 VDD.n491 VDD.t112 191.288
R185 VDD.t421 VDD.n206 191.288
R186 VDD.t321 VDD.n294 191.288
R187 VDD.n295 VDD.t242 191.288
R188 VDD.t226 VDD.n301 191.288
R189 VDD.n302 VDD.t302 191.288
R190 VDD.t135 VDD.n269 191.288
R191 VDD.n270 VDD.t355 191.288
R192 VDD.t228 VDD.n278 191.288
R193 VDD.n279 VDD.t411 191.288
R194 VDD.n346 VDD.t145 191.288
R195 VDD.n345 VDD.t340 191.288
R196 VDD.t74 VDD.n311 191.288
R197 VDD.n313 VDD.t413 191.288
R198 VDD.t140 VDD.n324 191.288
R199 VDD.n325 VDD.t88 191.288
R200 VDD.t72 VDD.n333 191.288
R201 VDD.n334 VDD.t49 191.288
R202 VDD.t201 VDD.t104 175.631
R203 VDD.t345 VDD.n135 153.678
R204 VDD.n394 VDD.t114 142.857
R205 VDD.n229 VDD.t54 142.857
R206 VDD.t295 VDD.n120 138.095
R207 VDD.n121 VDD.t314 138.095
R208 VDD.t0 VDD.n158 138.095
R209 VDD.t266 VDD.n159 138.095
R210 VDD.t176 VDD.n161 138.095
R211 VDD.t78 VDD.n163 138.095
R212 VDD.t312 VDD.n166 138.095
R213 VDD.t118 VDD.n199 138.095
R214 VDD.n219 VDD.t425 138.095
R215 VDD.t70 VDD.n224 138.095
R216 VDD.n235 VDD.t108 138.095
R217 VDD.n234 VDD.t280 138.095
R218 VDD.n4 VDD.t367 111.743
R219 VDD.n420 VDD.t283 111.743
R220 VDD.n421 VDD.t318 111.743
R221 VDD.n429 VDD.t384 111.743
R222 VDD.n430 VDD.t387 111.743
R223 VDD.n440 VDD.t377 111.743
R224 VDD.n447 VDD.t85 111.743
R225 VDD.n452 VDD.t244 111.743
R226 VDD.n453 VDD.t189 111.743
R227 VDD.t463 VDD.n503 111.743
R228 VDD.t250 VDD.n502 111.743
R229 VDD.n468 VDD.t11 111.743
R230 VDD.n470 VDD.t18 111.743
R231 VDD.n481 VDD.t256 111.743
R232 VDD.n482 VDD.t466 111.743
R233 VDD.n490 VDD.t435 111.743
R234 VDD.n491 VDD.t453 111.743
R235 VDD.n206 VDD.t137 111.743
R236 VDD.n294 VDD.t418 111.743
R237 VDD.n295 VDD.t427 111.743
R238 VDD.n301 VDD.t233 111.743
R239 VDD.n302 VDD.t215 111.743
R240 VDD.n269 VDD.t272 111.743
R241 VDD.n270 VDD.t309 111.743
R242 VDD.n278 VDD.t239 111.743
R243 VDD.n279 VDD.t230 111.743
R244 VDD.n346 VDD.t443 111.743
R245 VDD.t408 VDD.n345 111.743
R246 VDD.n311 VDD.t209 111.743
R247 VDD.n313 VDD.t212 111.743
R248 VDD.n324 VDD.t276 111.743
R249 VDD.n325 VDD.t337 111.743
R250 VDD.n333 VDD.t342 111.743
R251 VDD.n334 VDD.t289 111.743
R252 VDD.t218 VDD.n394 111.112
R253 VDD.n229 VDD.t5 111.112
R254 VDD.n142 VDD.t28 109.849
R255 VDD.n147 VDD.t396 109.849
R256 VDD.n152 VDD.t150 109.849
R257 VDD.t174 VDD.n366 109.849
R258 VDD.t199 VDD.n368 109.849
R259 VDD.t93 VDD.n371 109.849
R260 VDD.n374 VDD.t263 109.849
R261 VDD.t133 VDD.n173 109.849
R262 VDD.t221 VDD.n175 109.849
R263 VDD.t297 VDD.n178 109.849
R264 VDD.n181 VDD.t260 109.849
R265 VDD.n80 VDD.t423 109.849
R266 VDD.t202 VDD.n86 109.849
R267 VDD.n87 VDD.t194 109.849
R268 VDD.t433 VDD.n92 109.849
R269 VDD.t192 VDD.n25 109.849
R270 VDD.t181 VDD.n27 109.849
R271 VDD.t253 VDD.n30 109.849
R272 VDD.n33 VDD.t287 109.849
R273 VDD.t110 VDD.n96 109.849
R274 VDD.t100 VDD.n98 109.849
R275 VDD.t187 VDD.n101 109.849
R276 VDD.n104 VDD.t269 109.849
R277 VDD.n439 VDD.t448 62.1896
R278 VDD.n504 VDD.t362 62.1896
R279 VDD.n285 VDD.t142 62.1896
R280 VDD.n307 VDD.t147 62.1896
R281 VDD.n393 VDD.t440 61.8817
R282 VDD.n228 VDD.t55 61.8817
R283 VDD.n395 VDD.t292 60.9761
R284 VDD.n208 VDD.t2 60.9761
R285 VDD.n93 VDD.t33 59.702
R286 VDD.n146 VDD.t95 59.4064
R287 VDD.n151 VDD.t307 59.4064
R288 VDD.n141 VDD.t446 59.1138
R289 VDD.t185 VDD.n136 55.0852
R290 VDD.t183 VDD.n140 55.0852
R291 VDD.n407 VDD.t255 30.9379
R292 VDD.n259 VDD.t275 30.9379
R293 VDD.n34 VDD.t286 30.9379
R294 VDD.n36 VDD.t262 30.9379
R295 VDD.n57 VDD.t265 30.721
R296 VDD.n47 VDD.t279 30.7203
R297 VDD.n54 VDD.t268 30.3459
R298 VDD.n410 VDD.t282 30.2877
R299 VDD.n258 VDD.t271 30.2877
R300 VDD.n42 VDD.t259 30.0062
R301 VDD.n54 VDD.t477 24.8618
R302 VDD.n411 VDD.t474 24.5101
R303 VDD.n407 VDD.t469 24.5101
R304 VDD.n257 VDD.t480 24.5101
R305 VDD.n259 VDD.t475 24.5101
R306 VDD.n34 VDD.t471 24.5101
R307 VDD.n36 VDD.t479 24.5101
R308 VDD.n57 VDD.t478 24.4816
R309 VDD.n47 VDD.t473 24.4814
R310 VDD.n44 VDD.t482 24.4392
R311 VDD.n135 VDD.t201 21.9544
R312 VDD VDD.t152 10.5649
R313 VDD.t329 VDD 10.5649
R314 VDD VDD.t23 10.5649
R315 VDD.n261 VDD.n260 8.14231
R316 VDD.n409 VDD.n408 8.14083
R317 VDD.n412 VDD.n411 8.0005
R318 VDD.n257 VDD.n256 8.0005
R319 VDD.n44 VDD.n43 8.0005
R320 VDD.n64 VDD.n63 6.39748
R321 VDD VDD.n219 6.30459
R322 VDD.n420 VDD.n419 6.3005
R323 VDD.n422 VDD.n421 6.3005
R324 VDD.n429 VDD.n428 6.3005
R325 VDD.n431 VDD.n430 6.3005
R326 VDD.n441 VDD.n440 6.3005
R327 VDD.n447 VDD.n446 6.3005
R328 VDD.n452 VDD.n451 6.3005
R329 VDD.n454 VDD.n453 6.3005
R330 VDD.n481 VDD.n480 6.3005
R331 VDD.n483 VDD.n482 6.3005
R332 VDD.n490 VDD.n489 6.3005
R333 VDD.n492 VDD.n491 6.3005
R334 VDD.n502 VDD.n501 6.3005
R335 VDD.n498 VDD.n468 6.3005
R336 VDD.n495 VDD.n470 6.3005
R337 VDD.n503 VDD.n460 6.3005
R338 VDD.n398 VDD.n4 6.3005
R339 VDD.n394 VDD.n8 6.3005
R340 VDD.n375 VDD.n374 6.3005
R341 VDD.n378 VDD.n371 6.3005
R342 VDD.n381 VDD.n368 6.3005
R343 VDD.n384 VDD.n366 6.3005
R344 VDD.n234 VDD.n217 6.3005
R345 VDD.n230 VDD.n229 6.3005
R346 VDD.n236 VDD.n235 6.3005
R347 VDD.n224 VDD.n223 6.3005
R348 VDD.n243 VDD.n206 6.3005
R349 VDD.n294 VDD.n293 6.3005
R350 VDD.n296 VDD.n295 6.3005
R351 VDD.n301 VDD.n300 6.3005
R352 VDD.n303 VDD.n302 6.3005
R353 VDD.n280 VDD.n279 6.3005
R354 VDD.n278 VDD.n277 6.3005
R355 VDD.n271 VDD.n270 6.3005
R356 VDD.n269 VDD.n268 6.3005
R357 VDD.n324 VDD.n323 6.3005
R358 VDD.n326 VDD.n325 6.3005
R359 VDD.n333 VDD.n332 6.3005
R360 VDD.n335 VDD.n334 6.3005
R361 VDD.n345 VDD.n344 6.3005
R362 VDD.n341 VDD.n311 6.3005
R363 VDD.n338 VDD.n313 6.3005
R364 VDD.n347 VDD.n346 6.3005
R365 VDD.n182 VDD.n181 6.3005
R366 VDD.n185 VDD.n178 6.3005
R367 VDD.n188 VDD.n175 6.3005
R368 VDD.n191 VDD.n173 6.3005
R369 VDD.n199 VDD.n198 6.3005
R370 VDD.n355 VDD.n166 6.3005
R371 VDD.n359 VDD.n163 6.3005
R372 VDD.n362 VDD.n161 6.3005
R373 VDD.n159 VDD.n11 6.3005
R374 VDD.n68 VDD.n33 6.3005
R375 VDD.n71 VDD.n30 6.3005
R376 VDD.n74 VDD.n27 6.3005
R377 VDD.n77 VDD.n25 6.3005
R378 VDD.n92 VDD.n91 6.3005
R379 VDD.n88 VDD.n87 6.3005
R380 VDD.n86 VDD.n85 6.3005
R381 VDD.n81 VDD.n80 6.3005
R382 VDD.n105 VDD.n104 6.3005
R383 VDD.n108 VDD.n101 6.3005
R384 VDD.n111 VDD.n98 6.3005
R385 VDD.n114 VDD.n96 6.3005
R386 VDD.n158 VDD.n157 6.3005
R387 VDD.n122 VDD.n121 6.3005
R388 VDD.n120 VDD.n119 6.3005
R389 VDD.n153 VDD.n152 6.3005
R390 VDD.n148 VDD.n147 6.3005
R391 VDD.n143 VDD.n142 6.3005
R392 VDD.n140 VDD.n139 6.3005
R393 VDD.n136 VDD 6.3005
R394 VDD.n135 VDD.n0 6.3005
R395 VDD.n240 VDD.n209 5.85007
R396 VDD.n53 VDD.n52 5.30657
R397 VDD.n480 VDD.n476 5.213
R398 VDD.n375 VDD.t264 5.213
R399 VDD.n323 VDD.n319 5.213
R400 VDD.n182 VDD.t261 5.213
R401 VDD.n105 VDD.t270 5.213
R402 VDD.n232 VDD.t281 5.16878
R403 VDD.n237 VDD.t109 5.16878
R404 VDD.n207 VDD.t71 5.16878
R405 VDD.n354 VDD.t313 5.16878
R406 VDD.n364 VDD.n363 5.16878
R407 VDD VDD.t330 5.16454
R408 VDD VDD.n438 5.16369
R409 VDD VDD.n284 5.16369
R410 VDD.n1 VDD.t383 5.15997
R411 VDD.n297 VDD.t243 5.15997
R412 VDD.n169 VDD.n168 5.15997
R413 VDD.n138 VDD.t184 5.14212
R414 VDD.n459 VDD.n458 5.13287
R415 VDD.n405 VDD.n404 5.13287
R416 VDD.n424 VDD.n401 5.13287
R417 VDD.n427 VDD.t17 5.13287
R418 VDD.n426 VDD.n425 5.13287
R419 VDD.n432 VDD.t462 5.13287
R420 VDD.n437 VDD.n436 5.13287
R421 VDD.n445 VDD.n435 5.13287
R422 VDD.n449 VDD.n448 5.13287
R423 VDD.n450 VDD.t15 5.13287
R424 VDD.n434 VDD.n433 5.13287
R425 VDD.n455 VDD.t45 5.13287
R426 VDD.n466 VDD.n461 5.13287
R427 VDD.n500 VDD.t439 5.13287
R428 VDD.n499 VDD.n467 5.13287
R429 VDD.n497 VDD.t61 5.13287
R430 VDD.n496 VDD.n469 5.13287
R431 VDD.n494 VDD.t381 5.13287
R432 VDD.n475 VDD.n474 5.13287
R433 VDD.n485 VDD.n471 5.13287
R434 VDD.n488 VDD.t59 5.13287
R435 VDD.n487 VDD.n486 5.13287
R436 VDD.n493 VDD.t113 5.13287
R437 VDD.n399 VDD.n3 5.13287
R438 VDD.n397 VDD.t460 5.13287
R439 VDD.n377 VDD.t94 5.13287
R440 VDD.n380 VDD.t200 5.13287
R441 VDD.n382 VDD.n367 5.13287
R442 VDD.n383 VDD.t175 5.13287
R443 VDD.n385 VDD.n365 5.13287
R444 VDD.n244 VDD.n205 5.13287
R445 VDD.n242 VDD.t422 5.13287
R446 VDD.n222 VDD.n218 5.13287
R447 VDD.n221 VDD.t426 5.13287
R448 VDD.n213 VDD.n212 5.13287
R449 VDD.n249 VDD.n248 5.13287
R450 VDD.n286 VDD.n283 5.13287
R451 VDD.n291 VDD.n290 5.13287
R452 VDD.n298 VDD.n282 5.13287
R453 VDD.n299 VDD.t227 5.13287
R454 VDD.n304 VDD.t303 5.13287
R455 VDD.n255 VDD.n254 5.13287
R456 VDD.n273 VDD.n251 5.13287
R457 VDD.n276 VDD.t229 5.13287
R458 VDD.n275 VDD.n274 5.13287
R459 VDD.n281 VDD.t412 5.13287
R460 VDD.n309 VDD.n308 5.13287
R461 VDD.n343 VDD.t341 5.13287
R462 VDD.n342 VDD.n310 5.13287
R463 VDD.n340 VDD.t75 5.13287
R464 VDD.n339 VDD.n312 5.13287
R465 VDD.n337 VDD.t414 5.13287
R466 VDD.n318 VDD.n317 5.13287
R467 VDD.n328 VDD.n314 5.13287
R468 VDD.n331 VDD.t73 5.13287
R469 VDD.n330 VDD.n329 5.13287
R470 VDD.n336 VDD.t50 5.13287
R471 VDD.n203 VDD.n171 5.13287
R472 VDD.n184 VDD.t298 5.13287
R473 VDD.n187 VDD.t222 5.13287
R474 VDD.n189 VDD.n174 5.13287
R475 VDD.n190 VDD.t134 5.13287
R476 VDD.n192 VDD.n172 5.13287
R477 VDD.n197 VDD.t119 5.13287
R478 VDD.n356 VDD.n165 5.13287
R479 VDD.n357 VDD.t79 5.13287
R480 VDD.n360 VDD.n162 5.13287
R481 VDD.n361 VDD.t177 5.13287
R482 VDD.n388 VDD.t267 5.13287
R483 VDD.n17 VDD.t434 5.13287
R484 VDD.n89 VDD.t195 5.13287
R485 VDD.n21 VDD.n20 5.13287
R486 VDD.n84 VDD.t203 5.13287
R487 VDD.n83 VDD.n22 5.13287
R488 VDD.n82 VDD.t424 5.13287
R489 VDD.n79 VDD.n23 5.13287
R490 VDD.n70 VDD.t254 5.13287
R491 VDD.n73 VDD.t182 5.13287
R492 VDD.n75 VDD.n26 5.13287
R493 VDD.n76 VDD.t193 5.13287
R494 VDD.n78 VDD.n24 5.13287
R495 VDD.n107 VDD.t188 5.13287
R496 VDD.n110 VDD.t101 5.13287
R497 VDD.n112 VDD.n97 5.13287
R498 VDD.n113 VDD.t111 5.13287
R499 VDD.n115 VDD.n95 5.13287
R500 VDD.n156 VDD.t1 5.13287
R501 VDD.n124 VDD.n13 5.13287
R502 VDD.n123 VDD.t315 5.13287
R503 VDD.n15 VDD.n14 5.13287
R504 VDD.n118 VDD.t296 5.13287
R505 VDD.n117 VDD.n16 5.13287
R506 VDD.n154 VDD.t151 5.13287
R507 VDD.n129 VDD.n128 5.13287
R508 VDD.n149 VDD.t397 5.13287
R509 VDD.n131 VDD.n130 5.13287
R510 VDD.n144 VDD.t29 5.13287
R511 VDD.n133 VDD.n132 5.13287
R512 VDD.n137 VDD.t186 5.09693
R513 VDD.n505 VDD.n457 5.09407
R514 VDD.n396 VDD.n5 5.09407
R515 VDD.n392 VDD.n9 5.09407
R516 VDD.n387 VDD.t153 5.09407
R517 VDD.n227 VDD.n226 5.09407
R518 VDD.n306 VDD.n250 5.09407
R519 VDD.n201 VDD.t24 5.09407
R520 VDD.n94 VDD.t34 5.09407
R521 VDD.n150 VDD.t308 5.09407
R522 VDD.n145 VDD.t96 5.09407
R523 VDD.n134 VDD.t447 5.09407
R524 VDD.n415 VDD.n414 4.8755
R525 VDD.n264 VDD.n263 4.8755
R526 VDD.n67 VDD.t288 4.8755
R527 VDD.n63 VDD.n53 4.84121
R528 VDD.n45 VDD.n44 4.5005
R529 VDD.n48 VDD.n46 4.5005
R530 VDD.n49 VDD.n46 4.5005
R531 VDD.n37 VDD.n35 4.5005
R532 VDD.n38 VDD.n35 4.5005
R533 VDD.n58 VDD.n56 4.5005
R534 VDD.n59 VDD.n56 4.5005
R535 VDD.n7 VDD.n6 4.12326
R536 VDD.n211 VDD.n210 4.12326
R537 VDD.n511 VDD.t346 3.94862
R538 VDD.n42 VDD.n41 3.61662
R539 VDD.n444 VDD.n443 2.88497
R540 VDD.n292 VDD.n288 2.88497
R541 VDD.n64 VDD.n34 2.88182
R542 VDD.n418 VDD.n417 2.85787
R543 VDD.n423 VDD.n403 2.85787
R544 VDD.n465 VDD.n463 2.85787
R545 VDD.n479 VDD.n478 2.85787
R546 VDD.n484 VDD.n473 2.85787
R547 VDD.n376 VDD.n373 2.85787
R548 VDD.n379 VDD.n370 2.85787
R549 VDD.n216 VDD.n215 2.85787
R550 VDD.n267 VDD.n266 2.85787
R551 VDD.n272 VDD.n253 2.85787
R552 VDD.n247 VDD.n246 2.85787
R553 VDD.n322 VDD.n321 2.85787
R554 VDD.n327 VDD.n316 2.85787
R555 VDD.n183 VDD.n180 2.85787
R556 VDD.n186 VDD.n177 2.85787
R557 VDD.n196 VDD.n195 2.85787
R558 VDD.n90 VDD.n19 2.85787
R559 VDD.n69 VDD.n32 2.85787
R560 VDD.n72 VDD.n29 2.85787
R561 VDD.n106 VDD.n103 2.85787
R562 VDD.n109 VDD.n100 2.85787
R563 VDD.n127 VDD.n126 2.85787
R564 VDD.n417 VDD.t373 2.2755
R565 VDD.n417 VDD.n416 2.2755
R566 VDD.n403 VDD.t351 2.2755
R567 VDD.n403 VDD.n402 2.2755
R568 VDD.n443 VDD.t452 2.2755
R569 VDD.n443 VDD.n442 2.2755
R570 VDD.n463 VDD.t366 2.2755
R571 VDD.n463 VDD.n462 2.2755
R572 VDD.n478 VDD.t371 2.2755
R573 VDD.n478 VDD.n477 2.2755
R574 VDD.n473 VDD.t361 2.2755
R575 VDD.n473 VDD.n472 2.2755
R576 VDD.n373 VDD.t158 2.2755
R577 VDD.n373 VDD.n372 2.2755
R578 VDD.n370 VDD.t77 2.2755
R579 VDD.n370 VDD.n369 2.2755
R580 VDD.n215 VDD.t84 2.2755
R581 VDD.n215 VDD.n214 2.2755
R582 VDD.n288 VDD.t322 2.2755
R583 VDD.n288 VDD.n287 2.2755
R584 VDD.n266 VDD.t136 2.2755
R585 VDD.n266 VDD.n265 2.2755
R586 VDD.n253 VDD.t356 2.2755
R587 VDD.n253 VDD.n252 2.2755
R588 VDD.n246 VDD.t146 2.2755
R589 VDD.n246 VDD.n245 2.2755
R590 VDD.n321 VDD.t141 2.2755
R591 VDD.n321 VDD.n320 2.2755
R592 VDD.n316 VDD.t89 2.2755
R593 VDD.n316 VDD.n315 2.2755
R594 VDD.n180 VDD.t22 2.2755
R595 VDD.n180 VDD.n179 2.2755
R596 VDD.n177 VDD.t69 2.2755
R597 VDD.n177 VDD.n176 2.2755
R598 VDD.n195 VDD.t123 2.2755
R599 VDD.n195 VDD.n194 2.2755
R600 VDD.n19 VDD.t121 2.2755
R601 VDD.n19 VDD.n18 2.2755
R602 VDD.n32 VDD.t103 2.2755
R603 VDD.n32 VDD.n31 2.2755
R604 VDD.n29 VDD.t205 2.2755
R605 VDD.n29 VDD.n28 2.2755
R606 VDD.n103 VDD.t399 2.2755
R607 VDD.n103 VDD.n102 2.2755
R608 VDD.n100 VDD.t317 2.2755
R609 VDD.n100 VDD.n99 2.2755
R610 VDD.n126 VDD.t407 2.2755
R611 VDD.n126 VDD.n125 2.2755
R612 VDD.n51 VDD.n50 2.2439
R613 VDD.n61 VDD.n60 2.2439
R614 VDD.n40 VDD.n39 2.24362
R615 VDD.n37 VDD.n36 2.12257
R616 VDD.n408 VDD.n407 2.11346
R617 VDD.n260 VDD.n259 2.11346
R618 VDD.n261 VDD.n258 1.8236
R619 VDD.n410 VDD.n409 1.82345
R620 VDD VDD.n459 1.81843
R621 VDD VDD.n437 1.81843
R622 VDD VDD.n249 1.81843
R623 VDD.n286 VDD 1.81843
R624 VDD.n55 VDD.n54 1.81789
R625 VDD.n388 VDD 1.77285
R626 VDD VDD.n17 1.77285
R627 VDD VDD.n149 1.77285
R628 VDD VDD.n144 1.77285
R629 VDD VDD.n232 1.70433
R630 VDD.n52 VDD.n51 1.62565
R631 VDD.n62 VDD.n61 1.62565
R632 VDD.n58 VDD.n57 1.39782
R633 VDD.n48 VDD.n47 1.39728
R634 VDD.n79 VDD.n78 1.16167
R635 VDD.n494 VDD.n493 1.16051
R636 VDD.n337 VDD.n336 1.16051
R637 VDD.n52 VDD.n45 1.12171
R638 VDD.n62 VDD.n55 1.12171
R639 VDD.n386 VDD.n385 1.07428
R640 VDD.n202 VDD.n192 1.07428
R641 VDD.n116 VDD.n115 1.07428
R642 VDD.n305 VDD.n281 1.0737
R643 VDD.n456 VDD.n432 1.01824
R644 VDD.n44 VDD.n42 0.840632
R645 VDD.n232 VDD.n231 0.788255
R646 VDD.n231 VDD.n227 0.760634
R647 VDD.n155 VDD.n154 0.715235
R648 VDD.n204 VDD.n203 0.671656
R649 VDD.n264 VDD.n262 0.608132
R650 VDD.n238 VDD.n237 0.593661
R651 VDD.n241 VDD.n207 0.593661
R652 VDD.n351 VDD.n170 0.593661
R653 VDD.n354 VDD.n353 0.593661
R654 VDD.n364 VDD.n10 0.593661
R655 VDD.n358 VDD.n164 0.557288
R656 VDD.n390 VDD.n389 0.557288
R657 VDD.n63 VDD.n62 0.5228
R658 VDD.n53 VDD.n40 0.497812
R659 VDD.n220 VDD.n204 0.488955
R660 VDD.n464 VDD 0.468385
R661 VDD VDD.n348 0.468385
R662 VDD.n231 VDD.n211 0.439524
R663 VDD.n411 VDD.n410 0.404541
R664 VDD.n258 VDD.n257 0.404541
R665 VDD.n444 VDD.n0 0.372824
R666 VDD.n509 VDD.n1 0.369535
R667 VDD.n292 VDD.n289 0.369535
R668 VDD.n297 VDD.n167 0.369535
R669 VDD.n352 VDD.n169 0.369535
R670 VDD.n508 VDD.n2 0.342778
R671 VDD.n507 VDD.n506 0.342778
R672 VDD.n510 VDD 0.338387
R673 VDD.n419 VDD.n415 0.337997
R674 VDD.n268 VDD.n264 0.337997
R675 VDD.n68 VDD.n67 0.337997
R676 VDD.n138 VDD 0.334577
R677 VDD.n67 VDD.n66 0.333658
R678 VDD.n350 VDD.n204 0.329033
R679 VDD.n415 VDD.n413 0.328132
R680 VDD.n139 VDD.n137 0.317357
R681 VDD.n390 VDD.n10 0.312894
R682 VDD.n508 VDD.n507 0.280925
R683 VDD.n239 VDD.n211 0.277085
R684 VDD.n351 VDD.n350 0.274194
R685 VDD.n418 VDD.n405 0.233919
R686 VDD.n424 VDD.n423 0.233919
R687 VDD.n479 VDD.n475 0.233919
R688 VDD.n485 VDD.n484 0.233919
R689 VDD.n380 VDD.n379 0.233919
R690 VDD.n377 VDD.n376 0.233919
R691 VDD.n267 VDD.n255 0.233919
R692 VDD.n273 VDD.n272 0.233919
R693 VDD.n322 VDD.n318 0.233919
R694 VDD.n328 VDD.n327 0.233919
R695 VDD.n187 VDD.n186 0.233919
R696 VDD.n184 VDD.n183 0.233919
R697 VDD.n73 VDD.n72 0.233919
R698 VDD.n70 VDD.n69 0.233919
R699 VDD.n110 VDD.n109 0.233919
R700 VDD.n107 VDD.n106 0.233919
R701 VDD.n507 VDD.n400 0.226218
R702 VDD.n509 VDD.n508 0.221851
R703 VDD.n349 VDD 0.184731
R704 VDD.n150 VDD.n129 0.170231
R705 VDD.n145 VDD.n131 0.170231
R706 VDD.n134 VDD.n133 0.170231
R707 VDD.n391 VDD.n390 0.169866
R708 VDD.n352 VDD.n351 0.161388
R709 VDD.n289 VDD.n10 0.154438
R710 VDD.n137 VDD 0.147133
R711 VDD.n305 VDD.n304 0.143967
R712 VDD.n203 VDD.n202 0.143501
R713 VDD.n117 VDD.n116 0.143501
R714 VDD.n427 VDD.n426 0.141016
R715 VDD.n488 VDD.n487 0.141016
R716 VDD.n500 VDD.n499 0.141016
R717 VDD.n497 VDD.n496 0.141016
R718 VDD.n383 VDD.n382 0.141016
R719 VDD.n222 VDD.n221 0.141016
R720 VDD.n276 VDD.n275 0.141016
R721 VDD.n331 VDD.n330 0.141016
R722 VDD.n343 VDD.n342 0.141016
R723 VDD.n340 VDD.n339 0.141016
R724 VDD.n190 VDD.n189 0.141016
R725 VDD.n357 VDD.n356 0.141016
R726 VDD.n361 VDD.n360 0.141016
R727 VDD.n76 VDD.n75 0.141016
R728 VDD.n83 VDD.n82 0.141016
R729 VDD.n84 VDD.n21 0.141016
R730 VDD.n113 VDD.n112 0.141016
R731 VDD.n118 VDD.n15 0.141016
R732 VDD.n124 VDD.n123 0.141016
R733 VDD.n306 VDD.n305 0.139745
R734 VDD.n387 VDD.n386 0.138896
R735 VDD.n116 VDD.n94 0.138896
R736 VDD.n392 VDD.n391 0.137219
R737 VDD.n167 VDD.n164 0.132199
R738 VDD.n456 VDD.n455 0.130793
R739 VDD.n353 VDD.n352 0.128029
R740 VDD VDD.n201 0.127858
R741 VDD.n289 VDD.n164 0.126986
R742 VDD.n353 VDD.n167 0.125597
R743 VDD.n445 VDD 0.123016
R744 VDD.n466 VDD 0.123016
R745 VDD VDD.n291 0.123016
R746 VDD.n309 VDD 0.123016
R747 VDD VDD.n89 0.122435
R748 VDD VDD.n400 0.122231
R749 VDD.n216 VDD 0.111984
R750 VDD.n196 VDD 0.111984
R751 VDD.n90 VDD 0.111984
R752 VDD VDD.n127 0.111984
R753 VDD VDD.n465 0.111403
R754 VDD VDD.n247 0.111403
R755 VDD.n55 VDD 0.110941
R756 VDD.n408 VDD 0.107393
R757 VDD.n260 VDD 0.107393
R758 VDD.n428 VDD.n427 0.107339
R759 VDD.n432 VDD.n431 0.107339
R760 VDD.n451 VDD.n450 0.107339
R761 VDD.n455 VDD.n454 0.107339
R762 VDD.n489 VDD.n488 0.107339
R763 VDD.n493 VDD.n492 0.107339
R764 VDD.n501 VDD.n500 0.107339
R765 VDD.n498 VDD.n497 0.107339
R766 VDD.n495 VDD.n494 0.107339
R767 VDD.n385 VDD.n384 0.107339
R768 VDD.n382 VDD.n381 0.107339
R769 VDD.n236 VDD.n213 0.107339
R770 VDD.n223 VDD.n222 0.107339
R771 VDD.n300 VDD.n299 0.107339
R772 VDD.n304 VDD.n303 0.107339
R773 VDD.n277 VDD.n276 0.107339
R774 VDD.n281 VDD.n280 0.107339
R775 VDD.n332 VDD.n331 0.107339
R776 VDD.n336 VDD.n335 0.107339
R777 VDD.n344 VDD.n343 0.107339
R778 VDD.n341 VDD.n340 0.107339
R779 VDD.n338 VDD.n337 0.107339
R780 VDD.n192 VDD.n191 0.107339
R781 VDD.n189 VDD.n188 0.107339
R782 VDD.n360 VDD.n359 0.107339
R783 VDD.n356 VDD.n355 0.107339
R784 VDD.n78 VDD.n77 0.107339
R785 VDD.n75 VDD.n74 0.107339
R786 VDD.n81 VDD.n79 0.107339
R787 VDD.n85 VDD.n83 0.107339
R788 VDD.n88 VDD.n21 0.107339
R789 VDD.n115 VDD.n114 0.107339
R790 VDD.n112 VDD.n111 0.107339
R791 VDD.n119 VDD.n117 0.107339
R792 VDD.n122 VDD.n15 0.107339
R793 VDD.n157 VDD.n124 0.107339
R794 VDD.n153 VDD.n129 0.107339
R795 VDD.n148 VDD.n131 0.107339
R796 VDD.n143 VDD.n133 0.107339
R797 VDD VDD.n418 0.106758
R798 VDD.n423 VDD 0.106758
R799 VDD VDD.n479 0.106758
R800 VDD.n484 VDD 0.106758
R801 VDD VDD.n267 0.106758
R802 VDD.n272 VDD 0.106758
R803 VDD VDD.n322 0.106758
R804 VDD.n327 VDD 0.106758
R805 VDD.n379 VDD 0.106177
R806 VDD.n376 VDD 0.106177
R807 VDD VDD.n216 0.106177
R808 VDD.n186 VDD 0.106177
R809 VDD.n183 VDD 0.106177
R810 VDD VDD.n196 0.106177
R811 VDD.n127 VDD 0.106177
R812 VDD.n72 VDD 0.106177
R813 VDD.n69 VDD 0.106177
R814 VDD VDD.n90 0.106177
R815 VDD.n109 VDD 0.106177
R816 VDD.n106 VDD 0.106177
R817 VDD.n391 VDD.n8 0.1004
R818 VDD.n256 VDD 0.100075
R819 VDD.n510 VDD.n509 0.0980478
R820 VDD VDD.n7 0.0975258
R821 VDD.n43 VDD 0.0839415
R822 VDD.n213 VDD.n207 0.0835323
R823 VDD.n155 VDD 0.082371
R824 VDD.n49 VDD 0.0816915
R825 VDD.n422 VDD.n405 0.080629
R826 VDD.n441 VDD.n437 0.080629
R827 VDD.n483 VDD.n475 0.080629
R828 VDD.n378 VDD.n377 0.080629
R829 VDD.n293 VDD.n286 0.080629
R830 VDD.n271 VDD.n255 0.080629
R831 VDD.n326 VDD.n318 0.080629
R832 VDD.n185 VDD.n184 0.080629
R833 VDD.n198 VDD.n197 0.080629
R834 VDD.n71 VDD.n70 0.080629
R835 VDD.n91 VDD.n17 0.080629
R836 VDD.n108 VDD.n107 0.080629
R837 VDD.n59 VDD 0.0805665
R838 VDD.n400 VDD.n399 0.0795385
R839 VDD VDD.n383 0.0794677
R840 VDD VDD.n380 0.0794677
R841 VDD VDD.n190 0.0794677
R842 VDD VDD.n187 0.0794677
R843 VDD VDD.n361 0.0794677
R844 VDD VDD.n76 0.0794677
R845 VDD VDD.n73 0.0794677
R846 VDD.n82 VDD 0.0794677
R847 VDD VDD.n84 0.0794677
R848 VDD.n89 VDD 0.0794677
R849 VDD VDD.n113 0.0794677
R850 VDD VDD.n110 0.0794677
R851 VDD VDD.n118 0.0794677
R852 VDD.n123 VDD 0.0794677
R853 VDD VDD.n156 0.0794677
R854 VDD VDD.n138 0.0794623
R855 VDD VDD.n424 0.0788871
R856 VDD.n426 VDD 0.0788871
R857 VDD VDD.n445 0.0788871
R858 VDD VDD.n449 0.0788871
R859 VDD VDD.n434 0.0788871
R860 VDD VDD.n485 0.0788871
R861 VDD.n487 VDD 0.0788871
R862 VDD VDD.n466 0.0788871
R863 VDD.n499 VDD 0.0788871
R864 VDD.n496 VDD 0.0788871
R865 VDD.n291 VDD 0.0788871
R866 VDD VDD.n298 0.0788871
R867 VDD VDD.n273 0.0788871
R868 VDD.n275 VDD 0.0788871
R869 VDD VDD.n328 0.0788871
R870 VDD.n330 VDD 0.0788871
R871 VDD VDD.n309 0.0788871
R872 VDD.n342 VDD 0.0788871
R873 VDD.n339 VDD 0.0788871
R874 VDD.n154 VDD 0.0759839
R875 VDD.n149 VDD 0.0759839
R876 VDD.n144 VDD 0.0759839
R877 VDD.n434 VDD.n2 0.0754032
R878 VDD.n364 VDD.n362 0.0748226
R879 VDD.n38 VDD 0.0738165
R880 VDD.n297 VDD.n296 0.0730806
R881 VDD.n66 VDD.n64 0.0725
R882 VDD VDD.n170 0.0717592
R883 VDD.n239 VDD.n238 0.071388
R884 VDD VDD.n387 0.0709717
R885 VDD.n201 VDD 0.0709717
R886 VDD.n94 VDD 0.0709717
R887 VDD VDD.n150 0.0709717
R888 VDD VDD.n145 0.0709717
R889 VDD VDD.n134 0.0709717
R890 VDD.n506 VDD.n456 0.0708636
R891 VDD.n397 VDD.n396 0.0704581
R892 VDD VDD.n392 0.0701226
R893 VDD VDD.n227 0.0701226
R894 VDD VDD.n306 0.0701226
R895 VDD.n65 VDD 0.0700455
R896 VDD.n358 VDD.n357 0.0695968
R897 VDD.n406 VDD 0.0690714
R898 VDD.n450 VDD.n2 0.0661129
R899 VDD VDD.n511 0.0659817
R900 VDD.n241 VDD 0.0656
R901 VDD.n386 VDD.n364 0.0639524
R902 VDD VDD.n292 0.0614677
R903 VDD.n240 VDD.n239 0.0611
R904 VDD.n299 VDD.n169 0.0608871
R905 VDD.n237 VDD 0.0603065
R906 VDD.n389 VDD.n388 0.0562419
R907 VDD.n398 VDD.n397 0.0557
R908 VDD.n243 VDD.n242 0.0557
R909 VDD.n464 VDD.n459 0.0556613
R910 VDD.n348 VDD.n249 0.0556613
R911 VDD VDD.n354 0.0556613
R912 VDD.n446 VDD.n1 0.0550806
R913 VDD.n505 VDD 0.0546389
R914 VDD.n221 VDD.n220 0.0515968
R915 VDD.n444 VDD 0.0510161
R916 VDD.n413 VDD.n406 0.0471071
R917 VDD.n66 VDD.n65 0.0455
R918 VDD VDD.n7 0.0437
R919 VDD.n511 VDD 0.0432575
R920 VDD.n506 VDD.n505 0.0430455
R921 VDD.n449 VDD.n1 0.0428871
R922 VDD.n465 VDD.n464 0.0417258
R923 VDD.n348 VDD.n247 0.0417258
R924 VDD.n156 VDD.n155 0.0405645
R925 VDD.n399 VDD 0.0392
R926 VDD.n244 VDD 0.0392
R927 VDD.n412 VDD.n409 0.0387493
R928 VDD.n197 VDD.n170 0.0382419
R929 VDD.n349 VDD.n244 0.038
R930 VDD.n232 VDD.n217 0.0370806
R931 VDD.n413 VDD.n412 0.0358571
R932 VDD.n262 VDD.n261 0.0344878
R933 VDD.n354 VDD 0.0341774
R934 VDD.n242 VDD.n241 0.0311
R935 VDD.n237 VDD 0.0295323
R936 VDD.n50 VDD.n49 0.0275
R937 VDD.n43 VDD.n41 0.0275
R938 VDD.n60 VDD.n59 0.026375
R939 VDD.n51 VDD.n46 0.025705
R940 VDD.n61 VDD.n56 0.025705
R941 VDD VDD.n207 0.0248871
R942 VDD.n298 VDD.n297 0.0248871
R943 VDD.n389 VDD.n11 0.0248871
R944 VDD.n396 VDD 0.0243065
R945 VDD.n220 VDD 0.0242273
R946 VDD.n238 VDD 0.0234344
R947 VDD VDD.n510 0.0211312
R948 VDD.n39 VDD.n38 0.02075
R949 VDD.n464 VDD.n460 0.0206923
R950 VDD.n348 VDD.n347 0.0206923
R951 VDD.n231 VDD.n230 0.017527
R952 VDD.n40 VDD.n35 0.0169383
R953 VDD VDD.n444 0.0167581
R954 VDD.n350 VDD.n349 0.0157185
R955 VDD.n262 VDD.n256 0.0119894
R956 VDD.n202 VDD 0.0115377
R957 VDD VDD.n358 0.010371
R958 VDD.n39 VDD.n37 0.0095
R959 VDD.n406 VDD 0.00907143
R960 VDD VDD.n169 0.00862903
R961 VDD.n292 VDD 0.00630645
R962 VDD VDD.n153 0.00514516
R963 VDD VDD.n148 0.00514516
R964 VDD VDD.n143 0.00514516
R965 VDD.n65 VDD 0.00459091
R966 VDD.n60 VDD.n58 0.003875
R967 VDD VDD.n398 0.0032
R968 VDD VDD.n243 0.0032
R969 VDD.n230 VDD 0.00293243
R970 VDD.n50 VDD.n48 0.00275
R971 VDD.n8 VDD 0.0026
R972 VDD.n428 VDD 0.00224194
R973 VDD.n431 VDD 0.00224194
R974 VDD.n446 VDD 0.00224194
R975 VDD.n451 VDD 0.00224194
R976 VDD.n454 VDD 0.00224194
R977 VDD.n489 VDD 0.00224194
R978 VDD.n492 VDD 0.00224194
R979 VDD.n501 VDD 0.00224194
R980 VDD VDD.n498 0.00224194
R981 VDD VDD.n495 0.00224194
R982 VDD.n296 VDD 0.00224194
R983 VDD.n300 VDD 0.00224194
R984 VDD.n303 VDD 0.00224194
R985 VDD.n277 VDD 0.00224194
R986 VDD.n280 VDD 0.00224194
R987 VDD.n332 VDD 0.00224194
R988 VDD.n335 VDD 0.00224194
R989 VDD.n344 VDD 0.00224194
R990 VDD VDD.n341 0.00224194
R991 VDD VDD.n338 0.00224194
R992 VDD.n139 VDD 0.00219811
R993 VDD.n384 VDD 0.00166129
R994 VDD.n381 VDD 0.00166129
R995 VDD VDD.n378 0.00166129
R996 VDD VDD.n375 0.00166129
R997 VDD.n217 VDD 0.00166129
R998 VDD VDD.n236 0.00166129
R999 VDD.n223 VDD 0.00166129
R1000 VDD.n191 VDD 0.00166129
R1001 VDD.n188 VDD 0.00166129
R1002 VDD VDD.n185 0.00166129
R1003 VDD VDD.n182 0.00166129
R1004 VDD.n198 VDD 0.00166129
R1005 VDD.n359 VDD 0.00166129
R1006 VDD.n355 VDD 0.00166129
R1007 VDD.n362 VDD 0.00166129
R1008 VDD VDD.n11 0.00166129
R1009 VDD.n77 VDD 0.00166129
R1010 VDD.n74 VDD 0.00166129
R1011 VDD VDD.n71 0.00166129
R1012 VDD VDD.n68 0.00166129
R1013 VDD VDD.n81 0.00166129
R1014 VDD.n85 VDD 0.00166129
R1015 VDD VDD.n88 0.00166129
R1016 VDD.n91 VDD 0.00166129
R1017 VDD.n114 VDD 0.00166129
R1018 VDD.n111 VDD 0.00166129
R1019 VDD VDD.n108 0.00166129
R1020 VDD VDD.n105 0.00166129
R1021 VDD.n119 VDD 0.00166129
R1022 VDD VDD.n122 0.00166129
R1023 VDD.n157 VDD 0.00166129
R1024 VDD.n45 VDD.n41 0.001625
R1025 VDD VDD.n240 0.0011
R1026 VDD.n419 VDD 0.00108064
R1027 VDD VDD.n422 0.00108064
R1028 VDD VDD.n441 0.00108064
R1029 VDD.n480 VDD 0.00108064
R1030 VDD VDD.n483 0.00108064
R1031 VDD.n293 VDD 0.00108064
R1032 VDD.n268 VDD 0.00108064
R1033 VDD VDD.n271 0.00108064
R1034 VDD.n323 VDD 0.00108064
R1035 VDD VDD.n326 0.00108064
R1036 VDD.n460 VDD 0.00107692
R1037 VDD.n347 VDD 0.00107692
R1038 VDD VDD.n0 0.000799003
R1039 VSS.n153 VSS.n152 20141.5
R1040 VSS.n279 VSS.n260 18801.2
R1041 VSS.n155 VSS.t242 18488.2
R1042 VSS.n284 VSS.n283 13936
R1043 VSS.n215 VSS.n67 9584.01
R1044 VSS.t32 VSS.n323 7469.08
R1045 VSS.n155 VSS.n154 6872.87
R1046 VSS.n104 VSS.t178 6700.22
R1047 VSS.n241 VSS.t164 6664.41
R1048 VSS.n278 VSS.n277 6129.95
R1049 VSS.n281 VSS.n280 5655.34
R1050 VSS.n198 VSS.t64 5525.09
R1051 VSS.n323 VSS.n32 5466.04
R1052 VSS.n283 VSS.n282 5050.96
R1053 VSS.t65 VSS.n155 4508.16
R1054 VSS.n282 VSS.n65 4367.83
R1055 VSS.n307 VSS.n15 3956.92
R1056 VSS.n198 VSS.n156 3904.35
R1057 VSS.n230 VSS.n66 3893.61
R1058 VSS.n250 VSS.n236 3893.61
R1059 VSS.n214 VSS.n68 3893.61
R1060 VSS.n282 VSS.n279 3791.26
R1061 VSS.n161 VSS.t112 3606.54
R1062 VSS.n282 VSS.n281 3531.55
R1063 VSS.t291 VSS.t110 3055.32
R1064 VSS.n284 VSS.t251 2673.11
R1065 VSS.t199 VSS.t263 2307.56
R1066 VSS.t30 VSS.t51 2307.56
R1067 VSS.t259 VSS.t155 2307.56
R1068 VSS.t247 VSS.t296 2307.56
R1069 VSS.t159 VSS.t252 2307.56
R1070 VSS.t8 VSS.t287 2307.56
R1071 VSS.t14 VSS.t38 2307.56
R1072 VSS.t129 VSS.t109 2307.56
R1073 VSS.t77 VSS.t121 2307.56
R1074 VSS.t282 VSS.t23 2307.56
R1075 VSS.t60 VSS.t207 2307.56
R1076 VSS.t0 VSS.t269 2307.56
R1077 VSS.t97 VSS.t171 2307.56
R1078 VSS.t105 VSS.t81 2307.56
R1079 VSS.t47 VSS.t125 2307.56
R1080 VSS.t204 VSS.t78 2307.56
R1081 VSS.t75 VSS.t27 2307.56
R1082 VSS.t277 VSS.t222 2307.56
R1083 VSS.t41 VSS.t143 2307.56
R1084 VSS.t67 VSS.t50 2307.56
R1085 VSS.n289 VSS.t166 2214.94
R1086 VSS.t71 VSS.n289 2208.57
R1087 VSS.n307 VSS.t154 2042.72
R1088 VSS.t185 VSS.n121 2037.89
R1089 VSS.t175 VSS.n307 2037.89
R1090 VSS.t183 VSS.n68 1969.56
R1091 VSS.t173 VSS.n66 1969.56
R1092 VSS.n236 VSS.t169 1969.56
R1093 VSS.t267 VSS.n68 1964.9
R1094 VSS.n66 VSS.t96 1964.9
R1095 VSS.n236 VSS.t21 1964.9
R1096 VSS.t209 VSS.t299 1950.97
R1097 VSS.t260 VSS.t13 1950.97
R1098 VSS.t301 VSS.t74 1950.97
R1099 VSS.t37 VSS.t293 1950.97
R1100 VSS.t201 VSS.t198 1950.97
R1101 VSS.t224 VSS.t33 1950.97
R1102 VSS.t188 VSS.t44 1950.97
R1103 VSS.t119 VSS.t102 1881.09
R1104 VSS.t63 VSS.t162 1881.09
R1105 VSS.t40 VSS.t69 1881.09
R1106 VSS.t114 VSS.t266 1881.09
R1107 VSS.t80 VSS.t103 1881.09
R1108 VSS.t92 VSS.t56 1881.09
R1109 VSS.t223 VSS.t82 1881.09
R1110 VSS.t17 VSS.t196 1881.09
R1111 VSS.n279 VSS.n278 1724.9
R1112 VSS.n152 VSS.t29 1719.24
R1113 VSS.t270 VSS.n215 1713.53
R1114 VSS.n260 VSS.t79 1713.53
R1115 VSS.n249 VSS.t49 1713.53
R1116 VSS.n152 VSS.n151 1565.03
R1117 VSS.n288 VSS.n284 1565.03
R1118 VSS.n215 VSS.n214 1565.03
R1119 VSS.n260 VSS.n230 1565.03
R1120 VSS.n250 VSS.n249 1565.03
R1121 VSS.n104 VSS.t253 1199.47
R1122 VSS.t181 VSS.n241 1199.47
R1123 VSS.t281 VSS.n198 1153.78
R1124 VSS.t126 VSS.n156 1151.02
R1125 VSS.n323 VSS.t212 1108.08
R1126 VSS.n288 VSS.n287 1073.81
R1127 VSS.t241 VSS.t30 913.885
R1128 VSS.t252 VSS.t245 913.885
R1129 VSS.t22 VSS.t77 913.885
R1130 VSS.t269 VSS.t93 913.885
R1131 VSS.t78 VSS.t25 913.885
R1132 VSS.n173 VSS.t58 838.187
R1133 VSS.n12 VSS.t218 819.106
R1134 VSS.n105 VSS.t242 803.429
R1135 VSS.t299 VSS.t250 772.66
R1136 VSS.t234 VSS.t158 772.66
R1137 VSS.t74 VSS.t246 772.66
R1138 VSS.t237 VSS.t11 772.66
R1139 VSS.t198 VSS.t90 772.66
R1140 VSS.t236 VSS.t148 772.66
R1141 VSS.t33 VSS.t91 772.66
R1142 VSS.t54 VSS.t132 772.66
R1143 VSS.n289 VSS.n288 758.845
R1144 VSS.t232 VSS.t131 744.986
R1145 VSS.t26 VSS.t63 744.986
R1146 VSS.t233 VSS.t206 744.986
R1147 VSS.t266 VSS.t95 744.986
R1148 VSS.t235 VSS.t46 744.986
R1149 VSS.t20 VSS.t92 744.986
R1150 VSS.t55 VSS.t43 744.986
R1151 VSS.t221 VSS.t17 744.986
R1152 VSS.n159 VSS.t126 671.942
R1153 VSS.n154 VSS.n153 619.048
R1154 VSS.n164 VSS.t94 548.331
R1155 VSS.n166 VSS.t265 548.331
R1156 VSS.n163 VSS.t268 548.331
R1157 VSS.n103 VSS.t241 548.331
R1158 VSS.n102 VSS.t259 548.331
R1159 VSS.n101 VSS.t12 548.331
R1160 VSS.n97 VSS.t29 548.331
R1161 VSS.t287 VSS.n137 548.331
R1162 VSS.t38 VSS.n139 548.331
R1163 VSS.n141 VSS.t251 548.331
R1164 VSS.n199 VSS.t281 548.331
R1165 VSS.n202 VSS.t101 548.331
R1166 VSS.n207 VSS.t109 548.331
R1167 VSS.n208 VSS.t22 548.331
R1168 VSS.n216 VSS.t270 548.331
R1169 VSS.n221 VSS.t39 548.331
R1170 VSS.n222 VSS.t60 548.331
R1171 VSS.n227 VSS.t93 548.331
R1172 VSS.t79 VSS.n259 548.331
R1173 VSS.t81 VSS.n258 548.331
R1174 VSS.t125 VSS.n257 548.331
R1175 VSS.t49 VSS.n248 548.331
R1176 VSS.t222 VSS.n247 548.331
R1177 VSS.t143 VSS.n246 548.331
R1178 VSS.n242 VSS.t220 548.331
R1179 VSS.n159 VSS.t230 479.959
R1180 VSS.t250 VSS.n112 463.596
R1181 VSS.n113 VSS.t234 463.596
R1182 VSS.t13 VSS.n117 463.596
R1183 VSS.n118 VSS.t300 463.596
R1184 VSS.t246 VSS.n122 463.596
R1185 VSS.n124 VSS.t237 463.596
R1186 VSS.n126 VSS.t37 463.596
R1187 VSS.n290 VSS.t71 463.596
R1188 VSS.t90 VSS.n298 463.596
R1189 VSS.n299 VSS.t236 463.596
R1190 VSS.n302 VSS.t144 463.596
R1191 VSS.t154 VSS.n306 463.596
R1192 VSS.t91 VSS.n308 463.596
R1193 VSS.n310 VSS.t54 463.596
R1194 VSS.n324 VSS.t32 463.596
R1195 VSS.t64 VSS.n197 446.991
R1196 VSS.t102 VSS.n196 446.991
R1197 VSS.n188 VSS.t232 446.991
R1198 VSS.n189 VSS.t26 446.991
R1199 VSS.n69 VSS.t267 446.991
R1200 VSS.n70 VSS.t40 446.991
R1201 VSS.n72 VSS.t233 446.991
R1202 VSS.t95 VSS.n71 446.991
R1203 VSS.t96 VSS.n2 446.991
R1204 VSS.n3 VSS.t80 446.991
R1205 VSS.n4 VSS.t235 446.991
R1206 VSS.n5 VSS.t20 446.991
R1207 VSS.t21 VSS.n7 446.991
R1208 VSS.n8 VSS.t223 446.991
R1209 VSS.n9 VSS.t55 446.991
R1210 VSS.n10 VSS.t221 446.991
R1211 VSS.t263 VSS.n164 365.555
R1212 VSS.n166 VSS.t99 365.555
R1213 VSS.n163 VSS.t18 365.555
R1214 VSS.t253 VSS.n103 365.555
R1215 VSS.t51 VSS.n102 365.555
R1216 VSS.t155 VSS.n101 365.555
R1217 VSS.n97 VSS.t116 365.555
R1218 VSS.t296 VSS.n149 365.555
R1219 VSS.n137 VSS.t159 365.555
R1220 VSS.n139 VSS.t8 365.555
R1221 VSS.n141 VSS.t14 365.555
R1222 VSS.n199 VSS.t275 365.555
R1223 VSS.n202 VSS.t129 365.555
R1224 VSS.t121 VSS.n207 365.555
R1225 VSS.n208 VSS.t282 365.555
R1226 VSS.n216 VSS.t194 365.555
R1227 VSS.t207 VSS.n221 365.555
R1228 VSS.n222 VSS.t0 365.555
R1229 VSS.t171 VSS.n227 365.555
R1230 VSS.n259 VSS.t105 365.555
R1231 VSS.n258 VSS.t47 365.555
R1232 VSS.n257 VSS.t204 365.555
R1233 VSS.n252 VSS.t75 365.555
R1234 VSS.n248 VSS.t277 365.555
R1235 VSS.n247 VSS.t41 365.555
R1236 VSS.n246 VSS.t67 365.555
R1237 VSS.n242 VSS.t181 365.555
R1238 VSS.t87 VSS.t2 327.675
R1239 VSS.t238 VSS.t191 327.675
R1240 VSS.n112 VSS.t178 309.065
R1241 VSS.n113 VSS.t209 309.065
R1242 VSS.n117 VSS.t256 309.065
R1243 VSS.n118 VSS.t260 309.065
R1244 VSS.n122 VSS.t185 309.065
R1245 VSS.n124 VSS.t301 309.065
R1246 VSS.n126 VSS.t284 309.065
R1247 VSS.n290 VSS.t293 309.065
R1248 VSS.n298 VSS.t166 309.065
R1249 VSS.n299 VSS.t201 309.065
R1250 VSS.n302 VSS.t151 309.065
R1251 VSS.n306 VSS.t145 309.065
R1252 VSS.n308 VSS.t175 309.065
R1253 VSS.n310 VSS.t224 309.065
R1254 VSS.n312 VSS.t227 309.065
R1255 VSS.n324 VSS.t188 309.065
R1256 VSS.n197 VSS.t119 297.995
R1257 VSS.n196 VSS.t107 297.995
R1258 VSS.t162 VSS.n188 297.995
R1259 VSS.n189 VSS.t183 297.995
R1260 VSS.t69 VSS.n69 297.995
R1261 VSS.n70 VSS.t61 297.995
R1262 VSS.n72 VSS.t114 297.995
R1263 VSS.n71 VSS.t173 297.995
R1264 VSS.t103 VSS.n2 297.995
R1265 VSS.n3 VSS.t123 297.995
R1266 VSS.t56 VSS.n4 297.995
R1267 VSS.t169 VSS.n5 297.995
R1268 VSS.t82 VSS.n7 297.995
R1269 VSS.n8 VSS.t141 297.995
R1270 VSS.t196 VSS.n9 297.995
R1271 VSS.t164 VSS.n10 297.995
R1272 VSS.n32 VSS.n31 270.834
R1273 VSS.n277 VSS.n276 270.834
R1274 VSS.n32 VSS.n16 251.548
R1275 VSS.n277 VSS.n261 251.548
R1276 VSS.n30 VSS.t87 190.587
R1277 VSS.n275 VSS.t238 190.587
R1278 VSS.n32 VSS.t5 174.407
R1279 VSS.n277 VSS.t72 174.407
R1280 VSS.t18 VSS.n67 165.642
R1281 VSS.t112 VSS.n160 150.845
R1282 VSS.t110 VSS.n161 150.845
R1283 VSS.n214 VSS.n213 119.948
R1284 VSS.n230 VSS.n229 119.948
R1285 VSS.n251 VSS.n250 119.948
R1286 VSS.n151 VSS.n150 114.236
R1287 VSS.n323 VSS.n15 106.921
R1288 VSS.t5 VSS.t34 93.9117
R1289 VSS.t72 VSS.t288 93.9117
R1290 VSS.t45 VSS.t215 58.5375
R1291 VSS.n165 VSS.t199 34.2711
R1292 VSS.n162 VSS.t291 34.2711
R1293 VSS.n150 VSS.t247 34.2711
R1294 VSS.n287 VSS.t212 34.2711
R1295 VSS.n213 VSS.t23 34.2711
R1296 VSS.n229 VSS.t97 34.2711
R1297 VSS.t27 VSS.n251 34.2711
R1298 VSS.n173 VSS.n67 27.0388
R1299 VSS.n241 VSS.n12 26.4233
R1300 VSS.n322 VSS.t84 20.9066
R1301 VSS.n105 VSS.n104 20.7342
R1302 VSS.n31 VSS.n30 16.7186
R1303 VSS.n276 VSS.n275 16.7186
R1304 VSS.t84 VSS.t45 13.1415
R1305 VSS.n183 VSS.t231 9.37686
R1306 VSS.n235 VSS.t28 9.3736
R1307 VSS.n228 VSS.t98 9.3736
R1308 VSS.n212 VSS.t24 9.3736
R1309 VSS.n321 VSS.n33 9.37275
R1310 VSS.n286 VSS.n285 9.37275
R1311 VSS.n81 VSS.n80 9.37275
R1312 VSS.n106 VSS.n89 9.37275
R1313 VSS.n24 VSS.t31 9.3221
R1314 VSS.n26 VSS.n20 9.3221
R1315 VSS.n269 VSS.t73 9.3221
R1316 VSS.n271 VSS.n265 9.3221
R1317 VSS.n327 VSS.t219 9.30652
R1318 VSS.n28 VSS.n17 9.30652
R1319 VSS.n23 VSS.n21 9.30652
R1320 VSS.n273 VSS.n262 9.30652
R1321 VSS.n268 VSS.n266 9.30652
R1322 VSS.n177 VSS.t292 9.30652
R1323 VSS.n172 VSS.t59 9.30652
R1324 VSS.n168 VSS.t200 9.30652
R1325 VSS.n181 VSS.t113 9.30518
R1326 VSS.n179 VSS.t111 9.25414
R1327 VSS.n327 VSS.n326 7.3796
R1328 VSS VSS.n18 7.30633
R1329 VSS VSS.n263 7.30633
R1330 VSS VSS.t100 7.30633
R1331 VSS.n187 VSS.t120 7.19156
R1332 VSS.n194 VSS.t108 7.19156
R1333 VSS.n77 VSS.t70 7.19156
R1334 VSS.n75 VSS.t62 7.19156
R1335 VSS.n345 VSS.t104 7.19156
R1336 VSS.n343 VSS.t124 7.19156
R1337 VSS.n336 VSS.t83 7.19156
R1338 VSS.n334 VSS.t142 7.19156
R1339 VSS.n232 VSS.t106 7.19156
R1340 VSS.n234 VSS.t48 7.19156
R1341 VSS.n255 VSS.t205 7.19156
R1342 VSS.n218 VSS.t195 7.19156
R1343 VSS.n219 VSS.t208 7.19156
R1344 VSS.n224 VSS.t1 7.19156
R1345 VSS.n201 VSS.t276 7.19156
R1346 VSS.n204 VSS.t130 7.19156
R1347 VSS.n205 VSS.t122 7.19156
R1348 VSS.n14 VSS.n13 7.19156
R1349 VSS.n314 VSS.n311 7.19156
R1350 VSS.n39 VSS.n37 7.19156
R1351 VSS.n41 VSS.n36 7.19156
R1352 VSS.n43 VSS.n35 7.19156
R1353 VSS.n304 VSS.n47 7.19156
R1354 VSS.n301 VSS.n48 7.19156
R1355 VSS.n55 VSS.n53 7.19156
R1356 VSS.n57 VSS.n52 7.19156
R1357 VSS.n59 VSS.n51 7.19156
R1358 VSS.n64 VSS.n63 7.19156
R1359 VSS.n128 VSS.n125 7.19156
R1360 VSS.n143 VSS.n140 7.19156
R1361 VSS.n145 VSS.n138 7.19156
R1362 VSS.n147 VSS.n136 7.19156
R1363 VSS.n84 VSS.n83 7.19156
R1364 VSS.n115 VSS.n85 7.19156
R1365 VSS.n99 VSS.n96 7.19156
R1366 VSS.n95 VSS.n94 7.19156
R1367 VSS.n92 VSS.n91 7.19156
R1368 VSS.n238 VSS.t278 7.19156
R1369 VSS.n240 VSS.t42 7.19156
R1370 VSS.n244 VSS.t68 7.19156
R1371 VSS.n175 VSS.t19 6.88656
R1372 VSS.n170 VSS.t264 6.88656
R1373 VSS.n158 VSS.n157 6.01414
R1374 VSS.n158 VSS.t66 6.01414
R1375 VSS.n192 VSS.t163 5.91399
R1376 VSS.n190 VSS.t184 5.91399
R1377 VSS.n73 VSS.t115 5.91399
R1378 VSS.n348 VSS.t174 5.91399
R1379 VSS.n341 VSS.t57 5.91399
R1380 VSS.n339 VSS.t170 5.91399
R1381 VSS.n332 VSS.t197 5.91399
R1382 VSS.n330 VSS.t165 5.91399
R1383 VSS.n253 VSS.t76 5.91399
R1384 VSS.n225 VSS.t172 5.91399
R1385 VSS.n210 VSS.t283 5.91399
R1386 VSS.n316 VSS.n309 5.91399
R1387 VSS.n318 VSS.n46 5.91399
R1388 VSS.n45 VSS.n34 5.91399
R1389 VSS.n296 VSS.n295 5.91399
R1390 VSS.n294 VSS.n49 5.91399
R1391 VSS.n61 VSS.n50 5.91399
R1392 VSS.n130 VSS.n123 5.91399
R1393 VSS.n132 VSS.n120 5.91399
R1394 VSS.n135 VSS.n82 5.91399
R1395 VSS.n110 VSS.n109 5.91399
R1396 VSS.n108 VSS.n86 5.91399
R1397 VSS.n88 VSS.n87 5.91399
R1398 VSS.n11 VSS.t182 5.91399
R1399 VSS.n30 VSS.n29 5.2005
R1400 VSS.n22 VSS.n16 5.2005
R1401 VSS.n275 VSS.n274 5.2005
R1402 VSS.n267 VSS.n261 5.2005
R1403 VSS.n112 VSS.n111 5.2005
R1404 VSS.n114 VSS.n113 5.2005
R1405 VSS.n117 VSS.n116 5.2005
R1406 VSS.n119 VSS.n118 5.2005
R1407 VSS.n131 VSS.n122 5.2005
R1408 VSS.n129 VSS.n124 5.2005
R1409 VSS.n127 VSS.n126 5.2005
R1410 VSS.n291 VSS.n290 5.2005
R1411 VSS.n106 VSS.n105 5.2005
R1412 VSS.n167 VSS.n166 5.2005
R1413 VSS.n169 VSS.n165 5.2005
R1414 VSS.n171 VSS.n164 5.2005
R1415 VSS.n174 VSS.n173 5.2005
R1416 VSS.n178 VSS.n162 5.2005
R1417 VSS.n176 VSS.n163 5.2005
R1418 VSS.n184 VSS.n159 5.2005
R1419 VSS.n182 VSS.n160 5.2005
R1420 VSS.n180 VSS.n161 5.2005
R1421 VSS.n287 VSS.n286 5.2005
R1422 VSS.n142 VSS.n141 5.2005
R1423 VSS.n144 VSS.n139 5.2005
R1424 VSS.n146 VSS.n137 5.2005
R1425 VSS.n149 VSS.n148 5.2005
R1426 VSS.n150 VSS.n81 5.2005
R1427 VSS.n98 VSS.n97 5.2005
R1428 VSS.n101 VSS.n100 5.2005
R1429 VSS.n102 VSS.n93 5.2005
R1430 VSS.n103 VSS.n90 5.2005
R1431 VSS.n38 VSS.n15 5.2005
R1432 VSS.n40 VSS.n15 5.2005
R1433 VSS.n42 VSS.n15 5.2005
R1434 VSS.n44 VSS.n15 5.2005
R1435 VSS.n322 VSS.n321 5.2005
R1436 VSS.n54 VSS.n15 5.2005
R1437 VSS.n56 VSS.n15 5.2005
R1438 VSS.n58 VSS.n15 5.2005
R1439 VSS.n60 VSS.n15 5.2005
R1440 VSS.n298 VSS.n297 5.2005
R1441 VSS.n300 VSS.n299 5.2005
R1442 VSS.n303 VSS.n302 5.2005
R1443 VSS.n306 VSS.n305 5.2005
R1444 VSS.n317 VSS.n308 5.2005
R1445 VSS.n315 VSS.n310 5.2005
R1446 VSS.n313 VSS.n312 5.2005
R1447 VSS.n325 VSS.n324 5.2005
R1448 VSS.n328 VSS.n12 5.2005
R1449 VSS.n200 VSS.n199 5.2005
R1450 VSS.n203 VSS.n202 5.2005
R1451 VSS.n207 VSS.n206 5.2005
R1452 VSS.n209 VSS.n208 5.2005
R1453 VSS.n213 VSS.n212 5.2005
R1454 VSS.n217 VSS.n216 5.2005
R1455 VSS.n221 VSS.n220 5.2005
R1456 VSS.n223 VSS.n222 5.2005
R1457 VSS.n227 VSS.n226 5.2005
R1458 VSS.n229 VSS.n228 5.2005
R1459 VSS.n259 VSS.n231 5.2005
R1460 VSS.n258 VSS.n233 5.2005
R1461 VSS.n257 VSS.n256 5.2005
R1462 VSS.n254 VSS.n252 5.2005
R1463 VSS.n251 VSS.n235 5.2005
R1464 VSS.n243 VSS.n242 5.2005
R1465 VSS.n246 VSS.n245 5.2005
R1466 VSS.n247 VSS.n239 5.2005
R1467 VSS.n248 VSS.n237 5.2005
R1468 VSS.n331 VSS.n10 5.2005
R1469 VSS.n333 VSS.n9 5.2005
R1470 VSS.n335 VSS.n8 5.2005
R1471 VSS.n337 VSS.n7 5.2005
R1472 VSS.n340 VSS.n5 5.2005
R1473 VSS.n342 VSS.n4 5.2005
R1474 VSS.n344 VSS.n3 5.2005
R1475 VSS.n346 VSS.n2 5.2005
R1476 VSS.n71 VSS.n0 5.2005
R1477 VSS.n74 VSS.n72 5.2005
R1478 VSS.n76 VSS.n70 5.2005
R1479 VSS.n78 VSS.n69 5.2005
R1480 VSS.n191 VSS.n189 5.2005
R1481 VSS.n193 VSS.n188 5.2005
R1482 VSS.n196 VSS.n195 5.2005
R1483 VSS.n197 VSS.n186 5.2005
R1484 VSS.n185 VSS.n158 3.36323
R1485 VSS.n107 VSS 2.84263
R1486 VSS.n323 VSS.n322 2.38977
R1487 VSS.n292 VSS 2.24014
R1488 VSS VSS.n185 2.19933
R1489 VSS.n326 VSS 1.92724
R1490 VSS.n330 VSS.n329 0.917851
R1491 VSS.n108 VSS.n107 0.899322
R1492 VSS.n320 VSS.n319 0.846463
R1493 VSS.n293 VSS.n62 0.846463
R1494 VSS.n134 VSS.n133 0.846463
R1495 VSS.n338 VSS.n6 0.845914
R1496 VSS.n347 VSS.n1 0.845914
R1497 VSS.n211 VSS.n79 0.845914
R1498 VSS.n156 VSS.t65 0.631859
R1499 VSS.n177 VSS.n176 0.396455
R1500 VSS.n168 VSS.n167 0.396455
R1501 VSS.n172 VSS.n171 0.396455
R1502 VSS.n326 VSS 0.392281
R1503 VSS.n183 VSS 0.379596
R1504 VSS VSS.n232 0.343161
R1505 VSS VSS.n234 0.343161
R1506 VSS VSS.n218 0.343161
R1507 VSS.n219 VSS 0.343161
R1508 VSS VSS.n201 0.343161
R1509 VSS VSS.n204 0.343161
R1510 VSS VSS.n41 0.343161
R1511 VSS VSS.n39 0.343161
R1512 VSS VSS.n57 0.343161
R1513 VSS VSS.n55 0.343161
R1514 VSS VSS.n145 0.343161
R1515 VSS VSS.n143 0.343161
R1516 VSS.n95 VSS 0.343161
R1517 VSS VSS.n99 0.343161
R1518 VSS VSS.n238 0.343161
R1519 VSS VSS.n240 0.343161
R1520 VSS.n181 VSS 0.310668
R1521 VSS.n27 VSS.n26 0.310174
R1522 VSS.n272 VSS.n271 0.310174
R1523 VSS VSS.n254 0.289491
R1524 VSS.n226 VSS 0.289491
R1525 VSS.n209 VSS 0.289491
R1526 VSS.n44 VSS 0.289491
R1527 VSS.n60 VSS 0.289491
R1528 VSS.n148 VSS 0.289491
R1529 VSS VSS.n90 0.289491
R1530 VSS VSS.n243 0.289491
R1531 VSS.n170 VSS 0.27984
R1532 VSS.n175 VSS 0.27984
R1533 VSS.n27 VSS.n19 0.254245
R1534 VSS.n272 VSS.n264 0.254245
R1535 VSS.n179 VSS 0.250123
R1536 VSS.n180 VSS.n179 0.247195
R1537 VSS VSS.n175 0.243604
R1538 VSS VSS.n170 0.243604
R1539 VSS.n111 VSS.n110 0.202392
R1540 VSS.n115 VSS.n114 0.202392
R1541 VSS.n131 VSS.n130 0.202392
R1542 VSS.n129 VSS.n128 0.202392
R1543 VSS.n297 VSS.n296 0.202392
R1544 VSS.n301 VSS.n300 0.202392
R1545 VSS.n317 VSS.n316 0.202392
R1546 VSS.n315 VSS.n314 0.202392
R1547 VSS.n347 VSS 0.199831
R1548 VSS.n293 VSS.n292 0.193357
R1549 VSS.n255 VSS 0.191234
R1550 VSS VSS.n224 0.191234
R1551 VSS.n205 VSS 0.191234
R1552 VSS VSS.n43 0.191234
R1553 VSS VSS.n59 0.191234
R1554 VSS VSS.n147 0.191234
R1555 VSS.n92 VSS 0.191234
R1556 VSS.n244 VSS 0.191234
R1557 VSS.n194 VSS.n193 0.18462
R1558 VSS.n192 VSS.n191 0.18462
R1559 VSS.n75 VSS.n74 0.18462
R1560 VSS.n73 VSS.n0 0.18462
R1561 VSS.n343 VSS.n342 0.18462
R1562 VSS.n341 VSS.n340 0.18462
R1563 VSS.n334 VSS.n333 0.18462
R1564 VSS.n332 VSS.n331 0.18462
R1565 VSS.n24 VSS.n23 0.168072
R1566 VSS.n269 VSS.n268 0.168072
R1567 VSS.n182 VSS.n181 0.152211
R1568 VSS VSS.n84 0.144708
R1569 VSS VSS.n64 0.144708
R1570 VSS.n304 VSS 0.144708
R1571 VSS VSS.n14 0.144708
R1572 VSS.n292 VSS 0.142971
R1573 VSS.n28 VSS.n27 0.142796
R1574 VSS.n273 VSS.n272 0.142796
R1575 VSS.n185 VSS.n184 0.138903
R1576 VSS VSS.n6 0.137685
R1577 VSS VSS.n1 0.137685
R1578 VSS VSS.n211 0.137685
R1579 VSS.n329 VSS 0.137685
R1580 VSS.n25 VSS.n24 0.137391
R1581 VSS.n270 VSS.n269 0.137391
R1582 VSS VSS.n320 0.137136
R1583 VSS VSS.n62 0.137136
R1584 VSS.n134 VSS 0.137136
R1585 VSS.n107 VSS.n88 0.136196
R1586 VSS VSS.n187 0.132014
R1587 VSS.n77 VSS 0.132014
R1588 VSS.n345 VSS 0.132014
R1589 VSS.n336 VSS 0.132014
R1590 VSS.n232 VSS.n231 0.118573
R1591 VSS.n234 VSS.n233 0.118573
R1592 VSS.n256 VSS.n255 0.118573
R1593 VSS.n218 VSS.n217 0.118573
R1594 VSS.n220 VSS.n219 0.118573
R1595 VSS.n224 VSS.n223 0.118573
R1596 VSS.n201 VSS.n200 0.118573
R1597 VSS.n204 VSS.n203 0.118573
R1598 VSS.n206 VSS.n205 0.118573
R1599 VSS.n43 VSS.n42 0.118573
R1600 VSS.n41 VSS.n40 0.118573
R1601 VSS.n39 VSS.n38 0.118573
R1602 VSS.n59 VSS.n58 0.118573
R1603 VSS.n57 VSS.n56 0.118573
R1604 VSS.n55 VSS.n54 0.118573
R1605 VSS.n147 VSS.n146 0.118573
R1606 VSS.n145 VSS.n144 0.118573
R1607 VSS.n143 VSS.n142 0.118573
R1608 VSS.n93 VSS.n92 0.118573
R1609 VSS.n100 VSS.n95 0.118573
R1610 VSS.n99 VSS.n98 0.118573
R1611 VSS.n238 VSS.n237 0.118573
R1612 VSS.n240 VSS.n239 0.118573
R1613 VSS.n245 VSS.n244 0.118573
R1614 VSS VSS.n253 0.115271
R1615 VSS VSS.n225 0.115271
R1616 VSS.n210 VSS 0.115271
R1617 VSS.n45 VSS 0.115271
R1618 VSS.n61 VSS 0.115271
R1619 VSS VSS.n135 0.115271
R1620 VSS VSS.n88 0.115271
R1621 VSS VSS.n11 0.115271
R1622 VSS.n26 VSS 0.114702
R1623 VSS.n271 VSS 0.114702
R1624 VSS.n79 VSS 0.114268
R1625 VSS VSS.n183 0.113945
R1626 VSS.n253 VSS.n6 0.10206
R1627 VSS.n225 VSS.n1 0.10206
R1628 VSS.n211 VSS.n210 0.10206
R1629 VSS.n320 VSS.n45 0.10206
R1630 VSS.n62 VSS.n61 0.10206
R1631 VSS.n135 VSS.n134 0.10206
R1632 VSS.n329 VSS.n11 0.10206
R1633 VSS.n338 VSS 0.0835282
R1634 VSS.n133 VSS.n132 0.0790328
R1635 VSS.n294 VSS.n293 0.0790328
R1636 VSS.n319 VSS.n318 0.0790328
R1637 VSS.n133 VSS 0.0779904
R1638 VSS.n319 VSS 0.0779904
R1639 VSS.n190 VSS.n79 0.0724366
R1640 VSS.n348 VSS.n347 0.0724366
R1641 VSS.n339 VSS.n338 0.0724366
R1642 VSS.n328 VSS.n327 0.0675755
R1643 VSS.n178 VSS.n177 0.0675755
R1644 VSS.n169 VSS.n168 0.0675755
R1645 VSS.n174 VSS.n172 0.0675755
R1646 VSS.n29 VSS.n28 0.0667264
R1647 VSS.n274 VSS.n273 0.0667264
R1648 VSS.n23 VSS.n22 0.0557756
R1649 VSS.n268 VSS.n267 0.0557756
R1650 VSS.n116 VSS.n115 0.0501911
R1651 VSS.n119 VSS.n84 0.0501911
R1652 VSS.n128 VSS.n127 0.0501911
R1653 VSS.n291 VSS.n64 0.0501911
R1654 VSS.n303 VSS.n301 0.0501911
R1655 VSS.n305 VSS.n304 0.0501911
R1656 VSS.n314 VSS.n313 0.0501911
R1657 VSS.n325 VSS.n14 0.0501911
R1658 VSS VSS.n108 0.0488012
R1659 VSS.n110 VSS 0.0488012
R1660 VSS.n132 VSS 0.0488012
R1661 VSS.n130 VSS 0.0488012
R1662 VSS VSS.n294 0.0488012
R1663 VSS.n296 VSS 0.0488012
R1664 VSS.n318 VSS 0.0488012
R1665 VSS.n316 VSS 0.0488012
R1666 VSS.n187 VSS.n186 0.0458169
R1667 VSS.n195 VSS.n194 0.0458169
R1668 VSS.n78 VSS.n77 0.0458169
R1669 VSS.n76 VSS.n75 0.0458169
R1670 VSS.n346 VSS.n345 0.0458169
R1671 VSS.n344 VSS.n343 0.0458169
R1672 VSS.n337 VSS.n336 0.0458169
R1673 VSS.n335 VSS.n334 0.0458169
R1674 VSS VSS.n192 0.0445493
R1675 VSS VSS.n190 0.0445493
R1676 VSS VSS.n73 0.0445493
R1677 VSS VSS.n348 0.0445493
R1678 VSS VSS.n341 0.0445493
R1679 VSS VSS.n339 0.0445493
R1680 VSS VSS.n332 0.0445493
R1681 VSS VSS.n330 0.0445493
R1682 VSS.n231 VSS 0.00545413
R1683 VSS.n233 VSS 0.00545413
R1684 VSS.n256 VSS 0.00545413
R1685 VSS.n217 VSS 0.00545413
R1686 VSS.n220 VSS 0.00545413
R1687 VSS.n223 VSS 0.00545413
R1688 VSS.n200 VSS 0.00545413
R1689 VSS.n203 VSS 0.00545413
R1690 VSS.n206 VSS 0.00545413
R1691 VSS.n42 VSS 0.00545413
R1692 VSS.n40 VSS 0.00545413
R1693 VSS.n38 VSS 0.00545413
R1694 VSS.n58 VSS 0.00545413
R1695 VSS.n56 VSS 0.00545413
R1696 VSS.n54 VSS 0.00545413
R1697 VSS.n146 VSS 0.00545413
R1698 VSS.n144 VSS 0.00545413
R1699 VSS.n142 VSS 0.00545413
R1700 VSS VSS.n93 0.00545413
R1701 VSS.n100 VSS 0.00545413
R1702 VSS.n98 VSS 0.00545413
R1703 VSS.n237 VSS 0.00545413
R1704 VSS.n239 VSS 0.00545413
R1705 VSS.n245 VSS 0.00545413
R1706 VSS.n254 VSS 0.00380275
R1707 VSS.n226 VSS 0.00380275
R1708 VSS VSS.n209 0.00380275
R1709 VSS.n19 VSS 0.00380275
R1710 VSS VSS.n44 0.00380275
R1711 VSS VSS.n60 0.00380275
R1712 VSS.n264 VSS 0.00380275
R1713 VSS.n148 VSS 0.00380275
R1714 VSS.n90 VSS 0.00380275
R1715 VSS.n176 VSS 0.00380275
R1716 VSS.n167 VSS 0.00380275
R1717 VSS.n171 VSS 0.00380275
R1718 VSS.n243 VSS 0.00380275
R1719 VSS VSS.n25 0.00352521
R1720 VSS VSS.n270 0.00352521
R1721 VSS.n184 VSS 0.00352521
R1722 VSS.n116 VSS 0.00258494
R1723 VSS VSS.n119 0.00258494
R1724 VSS.n127 VSS 0.00258494
R1725 VSS VSS.n291 0.00258494
R1726 VSS VSS.n303 0.00258494
R1727 VSS.n305 VSS 0.00258494
R1728 VSS.n313 VSS 0.00258494
R1729 VSS VSS.n325 0.00258494
R1730 VSS.n186 VSS 0.00240141
R1731 VSS.n195 VSS 0.00240141
R1732 VSS VSS.n78 0.00240141
R1733 VSS VSS.n76 0.00240141
R1734 VSS VSS.n346 0.00240141
R1735 VSS VSS.n344 0.00240141
R1736 VSS VSS.n337 0.00240141
R1737 VSS VSS.n335 0.00240141
R1738 VSS.n235 VSS 0.00219811
R1739 VSS.n228 VSS 0.00219811
R1740 VSS.n212 VSS 0.00219811
R1741 VSS VSS.n328 0.00219811
R1742 VSS.n29 VSS 0.00219811
R1743 VSS.n321 VSS 0.00219811
R1744 VSS.n286 VSS 0.00219811
R1745 VSS.n274 VSS 0.00219811
R1746 VSS VSS.n81 0.00219811
R1747 VSS VSS.n106 0.00219811
R1748 VSS VSS.n182 0.00219811
R1749 VSS VSS.n180 0.00219811
R1750 VSS VSS.n178 0.00219811
R1751 VSS VSS.n169 0.00219811
R1752 VSS VSS.n174 0.00219811
R1753 VSS.n22 VSS 0.00191732
R1754 VSS.n267 VSS 0.00191732
R1755 VSS.n111 VSS 0.00188996
R1756 VSS.n114 VSS 0.00188996
R1757 VSS VSS.n131 0.00188996
R1758 VSS VSS.n129 0.00188996
R1759 VSS.n297 VSS 0.00188996
R1760 VSS.n300 VSS 0.00188996
R1761 VSS VSS.n317 0.00188996
R1762 VSS VSS.n315 0.00188996
R1763 VSS.n193 VSS 0.00176761
R1764 VSS.n191 VSS 0.00176761
R1765 VSS.n74 VSS 0.00176761
R1766 VSS VSS.n0 0.00176761
R1767 VSS.n342 VSS 0.00176761
R1768 VSS.n340 VSS 0.00176761
R1769 VSS.n333 VSS 0.00176761
R1770 VSS.n331 VSS 0.00176761
R1771 CLK_div_3_mag_1.Q0.n2 CLK_div_3_mag_1.Q0.t8 36.935
R1772 CLK_div_3_mag_1.Q0.n3 CLK_div_3_mag_1.Q0.t4 31.4332
R1773 CLK_div_3_mag_1.Q0.n5 CLK_div_3_mag_1.Q0.t6 29.8135
R1774 CLK_div_3_mag_1.Q0.n5 CLK_div_3_mag_1.Q0.t5 27.8352
R1775 CLK_div_3_mag_1.Q0.n2 CLK_div_3_mag_1.Q0.t7 18.1962
R1776 CLK_div_3_mag_1.Q0.n3 CLK_div_3_mag_1.Q0.t3 15.3826
R1777 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.t1 7.09905
R1778 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n3 6.86029
R1779 CLK_div_3_mag_1.Q0.n4 CLK_div_3_mag_1.Q0 5.01077
R1780 CLK_div_3_mag_1.Q0.n6 CLK_div_3_mag_1.Q0 3.41843
R1781 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n1 3.25053
R1782 CLK_div_3_mag_1.Q0.n1 CLK_div_3_mag_1.Q0.t0 2.2755
R1783 CLK_div_3_mag_1.Q0.n1 CLK_div_3_mag_1.Q0.n0 2.2755
R1784 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n6 2.2505
R1785 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n2 2.13459
R1786 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n5 1.74998
R1787 CLK_div_3_mag_1.Q0.n6 CLK_div_3_mag_1.Q0.n4 1.50381
R1788 CLK_div_3_mag_1.Q0.n4 CLK_div_3_mag_1.Q0 1.12067
R1789 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 37.1981
R1790 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_3_mag_1.JK_FF_mag_1.K.t3 31.4332
R1791 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 30.4613
R1792 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_3_mag_1.JK_FF_mag_1.K.t7 24.7562
R1793 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_3_mag_1.JK_FF_mag_1.K.t2 17.6611
R1794 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 15.3826
R1795 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K 12.0716
R1796 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n5 7.62076
R1797 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_3_mag_1.JK_FF_mag_1.K 6.09789
R1798 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 2.99416
R1799 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_3_mag_1.JK_FF_mag_1.K.t1 2.2755
R1800 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_3_mag_1.JK_FF_mag_1.K.n1 2.2755
R1801 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 2.2505
R1802 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K 2.24788
R1803 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 1.94903
R1804 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n4 1.81638
R1805 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n3 1.43706
R1806 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n7 0.4325
R1807 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 37.1981
R1808 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 31.4332
R1809 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 30.4613
R1810 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 24.7562
R1811 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 17.6611
R1812 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K.t2 15.3826
R1813 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 12.0716
R1814 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n5 7.62076
R1815 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R1816 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 2.99416
R1817 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t1 2.2755
R1818 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 2.2755
R1819 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2505
R1820 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.24788
R1821 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.94903
R1822 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.81638
R1823 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n3 1.43706
R1824 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n7 0.4325
R1825 CLK_div_3_mag_1.Q1.n5 CLK_div_3_mag_1.Q1.t7 36.935
R1826 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1.t5 31.4332
R1827 CLK_div_3_mag_1.Q1.n6 CLK_div_3_mag_1.Q1.t9 31.4332
R1828 CLK_div_3_mag_1.Q1.n3 CLK_div_3_mag_1.Q1.t10 30.4613
R1829 CLK_div_3_mag_1.Q1.n3 CLK_div_3_mag_1.Q1.t4 24.7562
R1830 CLK_div_3_mag_1.Q1.n5 CLK_div_3_mag_1.Q1.t3 18.1962
R1831 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1.t6 15.3826
R1832 CLK_div_3_mag_1.Q1.n6 CLK_div_3_mag_1.Q1.t8 15.3826
R1833 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1 8.5575
R1834 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.t1 7.09905
R1835 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n6 6.86029
R1836 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1 5.69501
R1837 CLK_div_3_mag_1.Q1.n7 CLK_div_3_mag_1.Q1 5.01077
R1838 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n1 3.25053
R1839 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n8 2.43532
R1840 CLK_div_3_mag_1.Q1.n1 CLK_div_3_mag_1.Q1.t2 2.2755
R1841 CLK_div_3_mag_1.Q1.n1 CLK_div_3_mag_1.Q1.n0 2.2755
R1842 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n5 2.13459
R1843 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n3 1.81638
R1844 CLK_div_3_mag_1.Q1.n8 CLK_div_3_mag_1.Q1.n7 1.45395
R1845 CLK_div_3_mag_1.Q1.n8 CLK_div_3_mag_1.Q1.n4 1.23718
R1846 CLK_div_3_mag_1.Q1.n7 CLK_div_3_mag_1.Q1 1.12067
R1847 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1 0.976433
R1848 CLK_div_3_mag_0.CLK.n8 CLK_div_3_mag_0.CLK.t3 36.935
R1849 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK.t6 36.935
R1850 CLK_div_3_mag_0.CLK.n12 CLK_div_3_mag_0.CLK.t12 36.935
R1851 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.t11 36.935
R1852 CLK_div_3_mag_0.CLK.n10 CLK_div_3_mag_0.CLK.t5 30.5752
R1853 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.t10 25.4744
R1854 CLK_div_3_mag_0.CLK.n6 CLK_div_3_mag_0.CLK.t8 25.4742
R1855 CLK_div_3_mag_0.CLK.n10 CLK_div_3_mag_0.CLK.t4 21.7814
R1856 CLK_div_3_mag_0.CLK.n8 CLK_div_3_mag_0.CLK.t14 18.1962
R1857 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK.t2 18.1962
R1858 CLK_div_3_mag_0.CLK.n12 CLK_div_3_mag_0.CLK.t9 18.1962
R1859 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.t7 18.1962
R1860 CLK_div_3_mag_0.CLK.n6 CLK_div_3_mag_0.CLK.t13 14.142
R1861 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.t15 14.1417
R1862 CLK_div_3_mag_0.CLK.n5 CLK_div_3_mag_0.CLK.t1 9.33985
R1863 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n11 7.41483
R1864 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK.n14 5.37091
R1865 CLK_div_3_mag_0.CLK.n5 CLK_div_3_mag_0.CLK.t0 5.17836
R1866 CLK_div_3_mag_0.CLK.n2 CLK_div_3_mag_0.CLK.n12 2.13265
R1867 CLK_div_3_mag_0.CLK.n2 CLK_div_3_mag_0.CLK 0.077103
R1868 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.n3 1.42996
R1869 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n2 1.11863
R1870 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.n3 1.19586
R1871 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n8 2.13265
R1872 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK.n10 1.80883
R1873 CLK_div_3_mag_0.CLK.n1 CLK_div_3_mag_0.CLK 2.63776
R1874 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK 2.51943
R1875 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK 2.13281
R1876 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK 2.13261
R1877 CLK_div_3_mag_0.CLK.n4 CLK_div_3_mag_0.CLK.n6 1.43004
R1878 CLK_div_3_mag_0.CLK.n3 CLK_div_3_mag_0.CLK 0.196041
R1879 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n4 0.196041
R1880 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n5 0.115328
R1881 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK 0.108371
R1882 CLK_div_3_mag_0.CLK.n4 CLK_div_3_mag_0.CLK.n15 1.19586
R1883 CLK_div_3_mag_0.CLK.n1 CLK_div_3_mag_0.CLK 1.11863
R1884 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.n0 1.01264
R1885 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK.n1 0.894314
R1886 CLK.n1 CLK.t5 36.935
R1887 CLK.n7 CLK.t11 36.935
R1888 CLK.n13 CLK.t7 36.935
R1889 CLK.n17 CLK.t8 36.935
R1890 CLK.n23 CLK.t3 30.5752
R1891 CLK.n30 CLK.t1 25.4744
R1892 CLK.n37 CLK.t12 25.4742
R1893 CLK.n23 CLK.t0 21.7814
R1894 CLK.n1 CLK.t13 18.1962
R1895 CLK.n7 CLK.t10 18.1962
R1896 CLK.n13 CLK.t2 18.1962
R1897 CLK.n17 CLK.t4 18.1962
R1898 CLK.n37 CLK.t6 14.142
R1899 CLK.n30 CLK.t9 14.1417
R1900 CLK.n25 CLK.n24 7.41483
R1901 CLK.n35 CLK.n34 5.37091
R1902 CLK.n12 CLK.n4 2.25107
R1903 CLK.n27 CLK.n16 2.25107
R1904 CLK.n33 CLK.n32 2.24352
R1905 CLK.n39 CLK.n36 2.24352
R1906 CLK.n20 CLK.n17 2.12464
R1907 CLK.n8 CLK.n7 2.12444
R1908 CLK.n2 CLK.n1 2.12188
R1909 CLK.n14 CLK.n13 2.12188
R1910 CLK.n24 CLK.n23 1.80883
R1911 CLK.n11 CLK.n10 1.71671
R1912 CLK.n25 CLK.n22 1.59838
R1913 CLK.n9 CLK.n8 1.50503
R1914 CLK.n21 CLK.n20 1.50503
R1915 CLK.n38 CLK.n37 1.42126
R1916 CLK.n31 CLK.n30 1.42118
R1917 CLK.n35 CLK.n12 0.882596
R1918 CLK.n34 CLK.n27 0.882596
R1919 CLK.n29 CLK 0.1605
R1920 CLK.n26 CLK.n25 0.118826
R1921 CLK.n24 CLK 0.108371
R1922 CLK.n34 CLK.n33 0.0733415
R1923 CLK.n36 CLK.n35 0.0733415
R1924 CLK CLK.n40 0.05925
R1925 CLK.n3 CLK 0.0457995
R1926 CLK.n5 CLK 0.0457995
R1927 CLK.n15 CLK 0.0457995
R1928 CLK.n18 CLK 0.0457995
R1929 CLK.n10 CLK.n9 0.0386356
R1930 CLK.n22 CLK.n21 0.0386356
R1931 CLK.n4 CLK.n3 0.0377414
R1932 CLK.n6 CLK.n5 0.0377414
R1933 CLK.n16 CLK.n15 0.0377414
R1934 CLK.n19 CLK.n18 0.0377414
R1935 CLK.n32 CLK.n29 0.03175
R1936 CLK.n40 CLK.n39 0.03175
R1937 CLK.n33 CLK.n28 0.0198632
R1938 CLK.n36 CLK.n0 0.0198632
R1939 CLK.n12 CLK.n11 0.0122182
R1940 CLK.n27 CLK.n26 0.0122182
R1941 CLK.n4 CLK.n2 0.00360345
R1942 CLK.n16 CLK.n14 0.00360345
R1943 CLK.n8 CLK.n6 0.00203726
R1944 CLK.n20 CLK.n19 0.00203726
R1945 CLK.n32 CLK.n31 0.00175
R1946 CLK.n39 CLK.n38 0.00175
R1947 RST.n26 RST.t12 37.2596
R1948 RST.n40 RST.t0 37.2594
R1949 RST.n34 RST.t11 36.935
R1950 RST.n21 RST.t6 36.935
R1951 RST.n12 RST.t3 36.935
R1952 RST.n10 RST.t5 36.935
R1953 RST.n16 RST.t15 36.935
R1954 RST.n5 RST.t10 36.859
R1955 RST.n34 RST.t7 18.1962
R1956 RST.n21 RST.t2 18.1962
R1957 RST.n12 RST.t1 18.1962
R1958 RST.n10 RST.t4 18.1962
R1959 RST.n16 RST.t14 18.1962
R1960 RST.n26 RST.t9 17.5947
R1961 RST.n40 RST.t13 17.594
R1962 RST.n3 RST.t8 17.236
R1963 RST.n39 RST.n18 6.53894
R1964 RST.n38 RST.n31 6.06869
R1965 RST.n14 RST.n13 5.39891
R1966 RST.n31 RST.n24 4.82595
R1967 RST.n38 RST.n37 4.82279
R1968 RST.n31 RST.n30 4.5933
R1969 RST.n50 RST.n49 4.52909
R1970 RST.n37 RST.n36 4.5005
R1971 RST.n24 RST.n23 4.5005
R1972 RST.n4 RST.n3 3.60685
R1973 RST.n15 RST.n14 3.52872
R1974 RST.n6 RST.n5 2.88526
R1975 RST.n46 RST.n45 2.8454
R1976 RST.n47 RST.n46 2.41332
R1977 RST.n50 RST.n48 2.25693
R1978 RST.n35 RST.n33 2.25022
R1979 RST.n22 RST.n20 2.25022
R1980 RST.n47 RST.n0 2.24413
R1981 RST.n45 RST.n43 2.24196
R1982 RST.n30 RST.n29 2.24196
R1983 RST.n13 RST.n12 2.13713
R1984 RST.n11 RST.n10 2.13713
R1985 RST.n17 RST.n16 2.1349
R1986 RST.n35 RST.n34 2.12393
R1987 RST.n22 RST.n21 2.12393
R1988 RST.n14 RST.n11 1.87041
R1989 RST RST.n17 1.81585
R1990 RST.n18 RST.n15 1.75158
R1991 RST.n18 RST 1.72336
R1992 RST.n8 RST.n7 1.51223
R1993 RST.n41 RST.n40 1.42237
R1994 RST.n27 RST.n26 1.42168
R1995 RST.n46 RST.n39 1.19738
R1996 RST.n15 RST.n9 1.12371
R1997 RST.n39 RST.n38 0.118716
R1998 RST.n17 RST 0.0687763
R1999 RST.n11 RST 0.06755
R2000 RST.n13 RST 0.0675495
R2001 RST.n32 RST 0.0584663
R2002 RST.n19 RST 0.0584663
R2003 RST.n42 RST 0.0394837
R2004 RST.n28 RST 0.0394837
R2005 RST.n1 RST 0.0394837
R2006 RST.n43 RST.n42 0.0377414
R2007 RST.n29 RST.n28 0.0377414
R2008 RST.n7 RST.n2 0.0367013
R2009 RST.n37 RST 0.0293
R2010 RST.n24 RST 0.0293
R2011 RST.n45 RST.n44 0.0238218
R2012 RST.n30 RST.n25 0.0238218
R2013 RST.n36 RST.n32 0.0196058
R2014 RST.n23 RST.n19 0.0196058
R2015 RST.n50 RST.n47 0.0152321
R2016 RST.n49 RST.n48 0.0073371
R2017 RST.n7 RST.n6 0.0051456
R2018 RST RST.n50 0.00437097
R2019 RST.n9 RST.n8 0.003875
R2020 RST.n43 RST.n41 0.00360345
R2021 RST.n29 RST.n27 0.00360345
R2022 RST.n36 RST.n35 0.00255119
R2023 RST.n23 RST.n22 0.00255119
R2024 RST.n2 RST.n1 0.00205172
R2025 RST.n6 RST.n4 0.00199457
R2026 RST.n33 RST 0.0017
R2027 RST.n20 RST 0.0017
R2028 CLK_div_3_mag_0.Q1.n5 CLK_div_3_mag_0.Q1.t9 36.935
R2029 CLK_div_3_mag_0.Q1.n2 CLK_div_3_mag_0.Q1.t8 31.4332
R2030 CLK_div_3_mag_0.Q1.n6 CLK_div_3_mag_0.Q1.t5 31.4332
R2031 CLK_div_3_mag_0.Q1.n3 CLK_div_3_mag_0.Q1.t4 30.4613
R2032 CLK_div_3_mag_0.Q1.n3 CLK_div_3_mag_0.Q1.t7 24.7562
R2033 CLK_div_3_mag_0.Q1.n5 CLK_div_3_mag_0.Q1.t6 18.1962
R2034 CLK_div_3_mag_0.Q1.n2 CLK_div_3_mag_0.Q1.t10 15.3826
R2035 CLK_div_3_mag_0.Q1.n6 CLK_div_3_mag_0.Q1.t3 15.3826
R2036 CLK_div_3_mag_0.Q1.n4 CLK_div_3_mag_0.Q1 8.5575
R2037 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.t1 7.09905
R2038 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n6 6.86029
R2039 CLK_div_3_mag_0.Q1.n2 CLK_div_3_mag_0.Q1 5.69501
R2040 CLK_div_3_mag_0.Q1.n7 CLK_div_3_mag_0.Q1 5.01077
R2041 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n1 3.25053
R2042 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n8 2.43532
R2043 CLK_div_3_mag_0.Q1.n1 CLK_div_3_mag_0.Q1.t0 2.2755
R2044 CLK_div_3_mag_0.Q1.n1 CLK_div_3_mag_0.Q1.n0 2.2755
R2045 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n5 2.13459
R2046 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q1.n3 1.81638
R2047 CLK_div_3_mag_0.Q1.n8 CLK_div_3_mag_0.Q1.n7 1.45395
R2048 CLK_div_3_mag_0.Q1.n8 CLK_div_3_mag_0.Q1.n4 1.23718
R2049 CLK_div_3_mag_0.Q1.n7 CLK_div_3_mag_0.Q1 1.12067
R2050 CLK_div_3_mag_0.Q1.n4 CLK_div_3_mag_0.Q1 0.976433
R2051 CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_10_mag_0.JK_FF_mag_2.K.t6 37.1986
R2052 CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_10_mag_0.JK_FF_mag_2.K.t8 31.528
R2053 CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_10_mag_0.JK_FF_mag_2.K.t3 30.6315
R2054 CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_10_mag_0.JK_FF_mag_2.K.t4 24.5953
R2055 CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_10_mag_0.JK_FF_mag_2.K.t5 17.6614
R2056 CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_10_mag_0.JK_FF_mag_2.K 17.0516
R2057 CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_10_mag_0.JK_FF_mag_2.K.t7 15.3826
R2058 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K.n1 7.62751
R2059 CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_10_mag_0.JK_FF_mag_2.K.n4 3.28711
R2060 CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_10_mag_0.JK_FF_mag_2.K.n7 2.99416
R2061 CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_10_mag_0.JK_FF_mag_2.K 2.81128
R2062 CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_10_mag_0.JK_FF_mag_2.K 2.67866
R2063 CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_10_mag_0.JK_FF_mag_2.K.t1 2.2755
R2064 CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_10_mag_0.JK_FF_mag_2.K.n6 2.2755
R2065 CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_10_mag_0.JK_FF_mag_2.K.n5 2.2505
R2066 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K.n3 1.80496
R2067 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K.n2 1.43709
R2068 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.K.n0 0.281955
R2069 Vdiv90.n4 Vdiv90.n3 9.28675
R2070 Vdiv90.n2 Vdiv90.n1 6.01414
R2071 Vdiv90.n2 Vdiv90.t2 6.01414
R2072 Vdiv90.n5 Vdiv90.n0 3.88449
R2073 Vdiv90.n4 Vdiv90.n2 3.74699
R2074 Vdiv90.n5 Vdiv90.n4 0.0331087
R2075 Vdiv90 Vdiv90.n5 0.00269512
C0 CLK_div_3_mag_1.or_2_mag_0.IN2 a_11779_8699# 7.48e-20
C1 CLK a_12061_10895# 0.00164f
C2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_14508_9798# 0.00378f
C3 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 0.69f
C4 CLK_div_10_mag_0.Q0 a_6026_4761# 0.0157f
C5 CLK_div_10_mag_0.Q3 a_13231_5814# 2.79e-20
C6 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C7 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK 0.235f
C8 RST a_4404_10895# 0.00123f
C9 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4738_4717# 0.0203f
C10 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4744_5858# 0.0202f
C11 a_13071_5814# a_13231_5814# 0.0504f
C12 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Q2 0.179f
C13 RST a_7191_4717# 0.00186f
C14 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00152f
C15 CLK_div_10_mag_0.JK_FF_mag_3.QB a_11342_5858# 2.96e-19
C16 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_14354_10895# 8.64e-19
C17 RST a_10363_9798# 3.96e-19
C18 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C19 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_10048_4717# 0.0202f
C20 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C21 CLK_div_10_mag_0.Q0 a_11342_5858# 6.06e-21
C22 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C23 VDD CLK_div_10_mag_0.JK_FF_mag_2.QB 0.913f
C24 RST CLK_div_10_mag_0.Q3 0.0395f
C25 VDD CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.514f
C26 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.and2_mag_0.OUT 0.144f
C27 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_8869_10895# 1.17e-20
C28 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_13790_10895# 0.0036f
C29 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C30 CLK_div_10_mag_0.Q0 a_5462_4761# 0.00859f
C31 a_7031_4717# a_7191_4717# 0.0504f
C32 RST a_3840_10895# 0.00114f
C33 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4174_4717# 1.5e-20
C34 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN Vdiv90 1.82e-19
C35 RST a_7031_4717# 0.00186f
C36 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C37 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.741f
C38 CLK_div_10_mag_0.JK_FF_mag_3.QB a_10778_5858# 3.25e-19
C39 CLK CLK_div_10_mag_0.Q2 8.71e-19
C40 CLK_div_3_mag_1.Q0 a_12221_10895# 0.00335f
C41 RST CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.96e-19
C42 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C43 CLK_div_3_mag_0.JK_FF_mag_1.QB a_5846_9798# 1.86e-20
C44 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C45 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_13225_4717# 1.46e-19
C46 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C47 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C48 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C49 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_8709_10895# 1.5e-20
C50 CLK CLK_div_10_mag_0.nor_3_mag_0.IN3 9.91e-21
C51 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0854f
C52 CLK_div_10_mag_0.Q0 a_4898_4717# 0.0101f
C53 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4014_4717# 1.17e-20
C54 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_11342_5858# 4.52e-20
C55 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_15124_7257# 5.39e-20
C56 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C57 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.312f
C58 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.251f
C59 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C60 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.999f
C61 RST a_6026_4761# 9.66e-19
C62 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00586f
C63 CLK_div_10_mag_0.JK_FF_mag_3.QB a_10214_5814# 0.00392f
C64 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_8889_5858# 0.00118f
C65 CLK_div_3_mag_1.Q0 a_12061_10895# 0.00789f
C66 CLK_div_3_mag_0.JK_FF_mag_1.QB a_5686_9798# 1.41e-20
C67 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C68 VDD CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C69 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.29e-19
C70 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8863_9798# 0.0203f
C71 a_11779_8699# CLK_div_10_mag_0.and2_mag_0.OUT 1.87e-19
C72 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.Q0 0.338f
C73 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.QB 0.103f
C74 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_8145_10895# 0.0203f
C75 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.113f
C76 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C77 CLK_div_10_mag_0.CLK CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.129f
C78 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.4f
C79 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_10778_5858# 0.0202f
C80 VDD CLK_div_3_mag_1.JK_FF_mag_1.QB 0.878f
C81 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_14964_7257# 9.16e-20
C82 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_11491_9798# 0.0202f
C83 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C84 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C85 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_12061_10895# 1.46e-19
C86 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q0 4.36e-20
C87 RST a_5462_4761# 9.41e-19
C88 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C89 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00174f
C90 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C91 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C92 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_2.K 9.73e-19
C93 CLK_div_3_mag_1.Q0 a_11497_10895# 0.0102f
C94 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_8325_5858# 0.011f
C95 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C96 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0798f
C97 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C98 a_10927_9798# CLK_div_3_mag_1.or_2_mag_0.IN2 4.9e-20
C99 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 9.71e-20
C100 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0215f
C101 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C102 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.QB 2.59e-21
C103 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8703_9798# 0.0732f
C104 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_7985_10895# 0.0733f
C105 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.or_2_mag_0.IN2 4.52e-20
C106 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.07f
C107 CLK a_11779_8699# 0.0103f
C108 RST a_10778_5858# 1.23e-20
C109 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C110 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C111 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C112 CLK_div_10_mag_0.and2_mag_0.OUT a_14923_5858# 1.54e-19
C113 VDD a_5846_9798# 2.21e-19
C114 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C115 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C116 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_2.K 0.0626f
C117 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_10927_9798# 4.52e-20
C118 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C119 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C120 RST a_4898_4717# 0.00186f
C121 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_7761_5858# 1.43e-19
C122 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C123 CLK_div_3_mag_1.Q0 a_11337_10895# 0.0101f
C124 VDD CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.468f
C125 CLK_div_3_mag_1.Q0 a_8869_10895# 1.38e-20
C126 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.K 0.0275f
C127 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C128 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 4.42e-19
C129 CLK a_12215_9798# 0.0101f
C130 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C131 CLK_div_10_mag_0.Q0 a_8889_5858# 9.26e-19
C132 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.7e-20
C133 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8139_9798# 0.00378f
C134 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C135 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_7421_10895# 0.00378f
C136 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C137 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C138 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C139 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C140 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.QB 1.33e-20
C141 a_11928_6955# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.29e-22
C142 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_5122_9798# 0.0697f
C143 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.K 0.289f
C144 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Q0 0.026f
C145 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.305f
C146 CLK_div_3_mag_1.JK_FF_mag_1.QB a_15072_9798# 0.00392f
C147 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_7197_5814# 0.00119f
C148 CLK_div_3_mag_1.Q0 a_10773_10895# 0.00859f
C149 CLK_div_3_mag_1.JK_FF_mag_1.QB a_14964_7257# 5.07e-21
C150 CLK_div_3_mag_1.Q0 a_10806_8231# 0.0134f
C151 CLK_div_3_mag_1.Q0 a_8709_10895# 1.09e-20
C152 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 0.338f
C153 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.11e-19
C154 VDD a_4437_8231# 0.165f
C155 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.17e-19
C156 CLK_div_3_mag_0.JK_FF_mag_1.K a_5686_9798# 0.00392f
C157 CLK a_12055_9798# 0.00939f
C158 RST CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0758f
C159 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C160 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00213f
C161 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C162 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.IN2 0.0655f
C163 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C164 VDD a_5122_9798# 3.14e-19
C165 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C166 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C167 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C168 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_7915_4717# 8.64e-19
C169 VDD CLK_div_3_mag_1.JK_FF_mag_1.K 2.41f
C170 CLK_div_3_mag_0.JK_FF_mag_1.K a_4437_8231# 0.00168f
C171 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_4558_9798# 0.0059f
C172 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_5852_10895# 1.17e-20
C173 CLK_div_10_mag_0.Q1 a_10772_4717# 3.6e-22
C174 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.Q2 0.98f
C175 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_10773_10895# 0.0036f
C176 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0384f
C177 CLK_div_3_mag_1.JK_FF_mag_1.QB a_14508_9798# 3.33e-19
C178 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_10806_8231# 1.4e-19
C179 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00511f
C180 CLK_div_3_mag_1.Q0 a_10209_10895# 0.0157f
C181 CLK_div_3_mag_1.JK_FF_mag_1.K Vdiv90 2.52e-19
C182 CLK_div_10_mag_0.Q0 a_7761_5858# 6.43e-21
C183 CLK a_11491_9798# 6.43e-21
C184 CLK_div_3_mag_0.JK_FF_mag_1.K a_5122_9798# 1.75e-19
C185 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0569f
C186 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K 8.36e-19
C187 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C188 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00722f
C189 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0905f
C190 VDD a_4558_9798# 3.14e-19
C191 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 4.39e-19
C192 VDD CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.431f
C193 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C194 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C195 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0854f
C196 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_5692_10895# 1.5e-20
C197 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_10927_9798# 0.069f
C198 CLK_div_10_mag_0.Q1 a_10208_4717# 0.00166f
C199 CLK_div_3_mag_1.JK_FF_mag_1.K a_15232_9798# 8.64e-19
C200 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C201 CLK_div_3_mag_1.JK_FF_mag_1.K a_15124_7257# 3.16e-19
C202 CLK_div_10_mag_0.Q0 a_7197_5814# 0.00939f
C203 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C204 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.337f
C205 CLK_div_3_mag_0.JK_FF_mag_1.K a_4558_9798# 2.96e-19
C206 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C207 a_10806_8231# CLK_div_10_mag_0.Q1 5.89e-19
C208 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Q3 0.124f
C209 CLK_div_10_mag_0.JK_FF_mag_2.K a_14923_5858# 0.0114f
C210 VDD CLK_div_10_mag_0.and2_mag_1.OUT 0.578f
C211 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C212 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C213 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C214 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_7011_9798# 4.52e-20
C215 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C216 VDD a_3994_9798# 3.56e-19
C217 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.nor_3_mag_0.IN3 1.41e-20
C218 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_5128_10895# 0.0203f
C219 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C220 CLK_div_10_mag_0.Q1 a_10048_4717# 0.00119f
C221 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_10363_9798# 0.00372f
C222 CLK_div_3_mag_1.Q0 a_12055_9798# 2.79e-20
C223 CLK_div_3_mag_0.Q0 a_5852_10895# 0.00335f
C224 CLK_div_3_mag_1.JK_FF_mag_1.QB a_13380_9798# 0.0112f
C225 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.178f
C226 RST CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00289f
C227 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_5872_5858# 0.00372f
C228 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB 0.878f
C229 CLK_div_3_mag_1.JK_FF_mag_1.K a_14964_7257# 3.16e-19
C230 CLK_div_10_mag_0.Q0 a_7037_5814# 0.0101f
C231 CLK_div_3_mag_0.JK_FF_mag_1.K a_3994_9798# 0.012f
C232 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_8709_10895# 1.46e-19
C233 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C234 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00178f
C235 CLK_div_10_mag_0.JK_FF_mag_2.K a_14359_5858# 2.96e-19
C236 RST CLK 0.0337f
C237 CLK CLK_div_10_mag_0.Q3 4.37e-20
C238 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0835f
C239 RST a_7761_5858# 1.37e-19
C240 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.K 0.783f
C241 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C242 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_4738_4717# 9.1e-19
C243 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_12055_9798# 0.00119f
C244 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C245 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C246 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C247 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C248 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4968_10895# 0.0733f
C249 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.131f
C250 CLK_div_3_mag_0.Q0 a_5692_10895# 0.00789f
C251 CLK_div_10_mag_0.Q1 a_9043_4761# 0.0157f
C252 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.or_2_mag_0.IN2 4.52e-20
C253 RST a_8863_9798# 6.26e-19
C254 RST CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0732f
C255 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_5308_5858# 0.069f
C256 CLK_div_10_mag_0.Q0 a_5872_5858# 0.069f
C257 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C258 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.64e-20
C259 CLK_div_10_mag_0.JK_FF_mag_2.K a_13795_5858# 3.25e-19
C260 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.193f
C261 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_12060_4761# 0.00372f
C262 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.25e-20
C263 RST a_7197_5814# 7.09e-19
C264 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_3.QB 5.7e-19
C265 RST CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 9.24e-20
C266 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C267 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C268 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_11491_9798# 1.43e-19
C269 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_4174_4717# 0.0731f
C270 RST CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0202f
C271 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4404_10895# 0.00378f
C272 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.K 0.487f
C273 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_14923_5858# 0.00118f
C274 a_10054_5814# a_10214_5814# 0.0504f
C275 CLK_div_10_mag_0.Q1 a_8479_4761# 0.00859f
C276 CLK_div_3_mag_0.Q0 a_5128_10895# 0.0102f
C277 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C278 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C279 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00481f
C280 RST a_8703_9798# 5.13e-19
C281 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_11928_6955# 0.069f
C282 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.175f
C283 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0334f
C284 CLK_div_10_mag_0.Q0 a_5308_5858# 6.06e-21
C285 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C286 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C287 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0147f
C288 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 0.0435f
C289 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.317f
C290 CLK_div_10_mag_0.JK_FF_mag_2.K a_13231_5814# 0.00486f
C291 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.or_2_mag_0.IN2 5.32e-19
C292 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_11496_4761# 0.069f
C293 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C294 RST a_7037_5814# 0.00109f
C295 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C296 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C297 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.QB 0.311f
C298 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_10927_9798# 0.011f
C299 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_4014_4717# 0.0202f
C300 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_12896_6955# 5.1e-20
C301 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.38e-19
C302 CLK_div_3_mag_1.JK_FF_mag_1.QB a_14514_10895# 0.00695f
C303 VDD CLK_div_10_mag_0.CLK 1.61f
C304 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.Q0 1.16f
C305 CLK_div_3_mag_1.Q0 a_10363_9798# 0.069f
C306 CLK_div_10_mag_0.Q1 a_7915_4717# 0.0101f
C307 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_14359_5858# 0.011f
C308 CLK_div_3_mag_0.Q0 a_4968_10895# 0.0101f
C309 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_11906_5858# 0.00372f
C310 VDD Vdiv90 0.105f
C311 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C312 RST a_8139_9798# 1.8e-19
C313 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C314 RST CLK_div_10_mag_0.JK_FF_mag_2.K 3.05f
C315 RST CLK_div_3_mag_1.Q0 0.337f
C316 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_2.K 2f
C317 CLK_div_10_mag_0.Q0 a_4738_4717# 0.0102f
C318 VDD CLK_div_3_mag_0.JK_FF_mag_1.K 2.36f
C319 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C320 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C321 CLK_div_10_mag_0.JK_FF_mag_2.K a_13071_5814# 0.00111f
C322 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_7421_10895# 0.0036f
C323 CLK_div_10_mag_0.and2_mag_1.OUT a_12896_6955# 3.92e-20
C324 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00311f
C325 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_10_mag_0.CLK 4.46e-19
C326 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_6026_4761# 0.00372f
C327 RST a_5872_5858# 0.00168f
C328 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_13949_4717# 8.64e-19
C329 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_4558_9798# 0.069f
C330 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_10363_9798# 0.00118f
C331 CLK_div_10_mag_0.JK_FF_mag_2.K a_7031_4717# 2.81e-19
C332 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5462_4761# 0.0036f
C333 CLK_div_3_mag_1.JK_FF_mag_1.QB a_14354_10895# 0.00696f
C334 VDD a_15232_9798# 5.99e-19
C335 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C336 RST CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.023f
C337 CLK_div_10_mag_0.Q1 a_7755_4717# 0.0102f
C338 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_13795_5858# 1.43e-19
C339 CLK_div_3_mag_0.Q0 a_4404_10895# 0.00859f
C340 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C341 VDD a_15124_7257# 0.0407f
C342 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_11342_5858# 0.069f
C343 RST a_7575_9798# 0.0011f
C344 CLK_div_10_mag_0.Q0 a_4174_4717# 0.00789f
C345 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C346 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.or_2_mag_0.IN2 3.81e-19
C347 RST CLK_div_10_mag_0.JK_FF_mag_0.K 1.55e-19
C348 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C349 CLK_div_10_mag_0.Q0 a_4180_5814# 2.79e-20
C350 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.125f
C351 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C352 a_15124_7257# Vdiv90 0.198f
C353 CLK_div_10_mag_0.JK_FF_mag_2.K a_11906_5858# 7.4e-19
C354 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_11337_10895# 8.64e-19
C355 CLK CLK_div_3_mag_1.or_2_mag_0.IN2 6.62e-20
C356 RST CLK_div_3_mag_0.Q0 0.163f
C357 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C358 CLK_div_10_mag_0.JK_FF_mag_0.K a_13071_5814# 8.64e-19
C359 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00157f
C360 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_5462_4761# 0.069f
C361 RST a_5308_5858# 0.00105f
C362 RST CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00352f
C363 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.652f
C364 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11496_4761# 0.0036f
C365 VDD a_15077_4761# 3.14e-19
C366 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_3994_9798# 0.00372f
C367 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C368 CLK_div_3_mag_1.JK_FF_mag_1.QB a_13790_10895# 0.00964f
C369 VDD a_15072_9798# 2.65e-19
C370 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_13231_5814# 0.00119f
C371 CLK_div_3_mag_0.Q0 a_3840_10895# 0.0157f
C372 CLK_div_10_mag_0.Q1 a_7191_4717# 0.00789f
C373 VDD a_14964_7257# 0.234f
C374 RST a_7011_9798# 0.00151f
C375 CLK_div_10_mag_0.Q0 a_4014_4717# 0.00335f
C376 CLK CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00302f
C377 VDD CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C378 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.2e-19
C379 RST CLK_div_10_mag_0.Q1 0.134f
C380 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 8.58e-20
C381 a_14964_7257# Vdiv90 0.0132f
C382 CLK_div_10_mag_0.JK_FF_mag_2.K a_11342_5858# 7.4e-19
C383 RST a_4738_4717# 8.64e-19
C384 RST CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00237f
C385 RST a_4744_5858# 7.59e-20
C386 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0263f
C387 VDD CLK_div_10_mag_0.JK_FF_mag_1.QB 0.92f
C388 VDD a_14513_4761# 3.14e-19
C389 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.or_2_mag_0.IN2 0.0445f
C390 CLK_div_3_mag_1.JK_FF_mag_1.QB a_13226_10895# 0.0811f
C391 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5692_10895# 1.46e-19
C392 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C393 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C394 VDD a_14508_9798# 3.14e-19
C395 CLK_div_10_mag_0.Q1 a_7031_4717# 0.00335f
C396 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.QB 0.307f
C397 VDD a_11928_6955# 3.14e-19
C398 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.Q0 5.62e-19
C399 VDD a_5410_8699# 5.92e-19
C400 a_15072_9798# a_15232_9798# 0.0504f
C401 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.28f
C402 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.15f
C403 CLK_div_10_mag_0.JK_FF_mag_2.K a_10778_5858# 3.12e-19
C404 a_14964_7257# a_15124_7257# 0.186f
C405 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_7761_5858# 0.00378f
C406 CLK_div_10_mag_0.JK_FF_mag_2.QB a_9043_4761# 0.0811f
C407 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C408 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 6.88e-21
C409 VDD a_12896_6955# 3.14e-19
C410 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0209f
C411 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C412 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C413 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.Q3 5.07e-21
C414 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C415 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C416 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C417 VDD a_13944_9798# 3.14e-19
C418 VDD a_10960_6955# 6e-19
C419 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.or_2_mag_0.IN2 0.0655f
C420 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.999f
C421 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q2 2.25e-19
C422 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_7197_5814# 0.0732f
C423 CLK_div_10_mag_0.JK_FF_mag_2.QB a_8479_4761# 0.00964f
C424 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_8325_5858# 0.0059f
C425 CLK_div_10_mag_0.JK_FF_mag_2.K a_10214_5814# 9.32e-19
C426 CLK CLK_div_10_mag_0.and2_mag_0.OUT 0.0104f
C427 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.0881f
C428 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C429 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C430 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_10208_4717# 1.46e-19
C431 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C432 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C433 VDD a_13789_4717# 2.21e-19
C434 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C435 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.652f
C436 VDD a_13380_9798# 3.56e-19
C437 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.159f
C438 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.98e-19
C439 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C440 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.or_2_mag_0.IN2 5.32e-19
C441 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_14359_5858# 5.94e-20
C442 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_3.QB 2.59e-21
C443 CLK_div_3_mag_1.JK_FF_mag_1.K a_11497_10895# 0.00695f
C444 CLK CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 7.81e-19
C445 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 0.198f
C446 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C447 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_15238_10895# 0.0202f
C448 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0151f
C449 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C450 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_7761_5858# 0.0697f
C451 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.QB 0.348f
C452 CLK_div_10_mag_0.JK_FF_mag_2.QB a_7915_4717# 0.00696f
C453 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_7037_5814# 0.0203f
C454 CLK_div_10_mag_0.JK_FF_mag_2.K a_10054_5814# 0.00111f
C455 CLK_div_10_mag_0.Q1 a_10778_5858# 1.25e-20
C456 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00243f
C457 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C458 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C459 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.27e-19
C460 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_10806_8231# 3.25e-19
C461 VDD a_15238_10895# 0.0132f
C462 CLK_div_3_mag_0.or_2_mag_0.IN2 a_4437_8231# 8.64e-19
C463 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C464 VDD a_13225_4717# 0.00299f
C465 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C466 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_4404_10895# 0.0036f
C467 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C468 CLK_div_3_mag_1.JK_FF_mag_1.QB a_12215_9798# 1.86e-20
C469 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.31f
C470 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_8479_4761# 0.00378f
C471 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C472 a_4738_4717# a_4898_4717# 0.0504f
C473 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.86e-19
C474 CLK_div_3_mag_1.JK_FF_mag_1.K a_11337_10895# 0.00696f
C475 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C476 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_11491_9798# 0.0697f
C477 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C478 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_15078_10895# 0.0731f
C479 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_10_mag_0.nor_3_mag_0.IN3 2.77e-19
C480 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_10_mag_0.Q1 9.34e-19
C481 RST CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0633f
C482 CLK_div_10_mag_0.JK_FF_mag_2.K a_8889_5858# 7.4e-19
C483 CLK_div_10_mag_0.JK_FF_mag_2.QB a_7755_4717# 0.00695f
C484 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00233f
C485 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C486 CLK_div_10_mag_0.Q1 a_10214_5814# 0.00939f
C487 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.013f
C488 VDD a_15078_10895# 0.00888f
C489 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_11779_8699# 0.069f
C490 VDD a_13065_4717# 0.00727f
C491 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_1.OUT 0.124f
C492 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.103f
C493 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C494 CLK_div_3_mag_1.JK_FF_mag_1.QB a_12055_9798# 1.41e-20
C495 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C496 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C497 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C498 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_7915_4717# 0.0733f
C499 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C500 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.K 0.00656f
C501 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_8139_9798# 0.0202f
C502 a_4558_9798# CLK_div_3_mag_0.or_2_mag_0.IN2 4.9e-20
C503 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C504 CLK_div_3_mag_1.JK_FF_mag_1.K a_10773_10895# 0.00964f
C505 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_10927_9798# 0.0059f
C506 CLK_div_3_mag_1.JK_FF_mag_1.K a_10806_8231# 0.00168f
C507 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_14514_10895# 9.1e-19
C508 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C509 CLK_div_10_mag_0.JK_FF_mag_2.K a_8325_5858# 7.4e-19
C510 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_1.OUT 0.0165f
C511 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C512 CLK_div_10_mag_0.Q1 a_10054_5814# 0.0101f
C513 VDD a_14514_10895# 0.0012f
C514 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C515 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C516 RST CLK_div_10_mag_0.JK_FF_mag_2.QB 0.183f
C517 VDD a_12060_4761# 0.00152f
C518 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C519 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0432f
C520 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C521 a_8703_9798# a_8863_9798# 0.0504f
C522 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C523 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C524 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C525 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C526 VDD a_12221_10895# 0.00743f
C527 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C528 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C529 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_7755_4717# 0.0203f
C530 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C531 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_7575_9798# 4.52e-20
C532 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.K 0.0659f
C533 CLK_div_3_mag_1.JK_FF_mag_1.K a_10209_10895# 0.0811f
C534 CLK_div_3_mag_1.Q0 CLK 0.149f
C535 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_14354_10895# 2.88e-20
C536 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C537 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.155f
C538 CLK_div_10_mag_0.JK_FF_mag_2.K a_7761_5858# 3.12e-19
C539 CLK_div_10_mag_0.Q1 a_8889_5858# 0.069f
C540 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C541 VDD a_14354_10895# 9.82e-19
C542 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C543 VDD a_11496_4761# 0.00152f
C544 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C545 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_13949_4717# 2.88e-20
C546 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C547 RST CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0172f
C548 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C549 a_13789_4717# a_13949_4717# 0.0504f
C550 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 4.42e-19
C551 CLK_div_3_mag_1.Q0 a_8863_9798# 3.69e-19
C552 a_7037_5814# a_7197_5814# 0.0504f
C553 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.K 1.41e-20
C554 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C555 VDD a_12061_10895# 0.00305f
C556 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_7191_4717# 1.5e-20
C557 CLK CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.471f
C558 a_10960_6955# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.36e-22
C559 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C560 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Q1 0.0529f
C561 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.268f
C562 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5872_5858# 0.00118f
C563 CLK_div_10_mag_0.JK_FF_mag_2.K a_7197_5814# 9.32e-19
C564 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C565 CLK_div_10_mag_0.Q1 a_8325_5858# 6.06e-21
C566 VDD a_13790_10895# 0.00149f
C567 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.065f
C568 VDD a_10932_4717# 0.00101f
C569 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_13789_4717# 9.1e-19
C570 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C571 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C572 VDD a_11497_10895# 2.21e-19
C573 VDD CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.441f
C574 CLK_div_3_mag_1.JK_FF_mag_1.K a_12055_9798# 0.00392f
C575 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.175f
C576 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C577 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.159f
C578 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_7031_4717# 1.17e-20
C579 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00675f
C580 a_11906_5858# CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C581 RST CLK_div_3_mag_1.JK_FF_mag_1.QB 0.59f
C582 a_5872_5858# CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C583 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.or_2_mag_0.IN2 1.82e-19
C584 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C585 CLK_div_10_mag_0.JK_FF_mag_2.K a_7037_5814# 0.00876f
C586 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.193f
C587 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C588 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5308_5858# 0.011f
C589 CLK CLK_div_10_mag_0.Q1 1.93e-19
C590 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C591 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C592 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C593 CLK_div_3_mag_0.JK_FF_mag_1.QB a_8145_10895# 0.00695f
C594 VDD a_13226_10895# 0.00149f
C595 VDD CLK_div_10_mag_0.Q2 2.86f
C596 VDD a_10772_4717# 0.00123f
C597 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_13225_4717# 0.0731f
C598 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_7915_4717# 2.88e-20
C599 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C600 RST CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.055f
C601 CLK_div_3_mag_1.JK_FF_mag_1.K a_11491_9798# 1.75e-19
C602 VDD CLK_div_10_mag_0.nor_3_mag_0.IN3 0.396f
C603 VDD a_8869_10895# 0.0132f
C604 RST a_5846_9798# 0.00222f
C605 VDD CLK_div_3_mag_0.or_2_mag_0.IN2 0.493f
C606 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.647f
C607 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_13795_5858# 0.00378f
C608 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.0881f
C609 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_4744_5858# 1.43e-19
C610 CLK_div_10_mag_0.nor_3_mag_0.IN3 Vdiv90 0.0263f
C611 CLK_div_10_mag_0.Q1 a_7197_5814# 2.79e-20
C612 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.QB 1e-19
C613 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C614 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C615 CLK_div_3_mag_0.JK_FF_mag_1.QB a_7985_10895# 0.00696f
C616 VDD a_10208_4717# 0.00891f
C617 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.or_2_mag_0.IN2 0.00761f
C618 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C619 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.QB 0.215f
C620 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_13065_4717# 0.0202f
C621 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C622 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.Q0 0.0116f
C623 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_7755_4717# 9.1e-19
C624 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C625 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.298f
C626 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_14513_4761# 0.00378f
C627 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_2.K 0.0156f
C628 CLK_div_10_mag_0.JK_FF_mag_2.QB a_10214_5814# 1.41e-20
C629 VDD a_10773_10895# 3.14e-19
C630 CLK_div_3_mag_1.JK_FF_mag_1.K a_10927_9798# 2.96e-19
C631 VDD a_10806_8231# 0.165f
C632 RST a_5686_9798# 0.00159f
C633 VDD a_8709_10895# 0.00888f
C634 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_13231_5814# 0.0732f
C635 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_14359_5858# 0.0059f
C636 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_4174_4717# 1.46e-19
C637 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11906_5858# 0.00118f
C638 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_13380_9798# 4.52e-20
C639 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C640 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_14964_7257# 2.85e-20
C641 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_4180_5814# 0.00119f
C642 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_1.OUT 2.11e-20
C643 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C644 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_15124_7257# 2.44e-20
C645 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.or_2_mag_0.IN2 1.82e-19
C646 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_12215_9798# 0.0203f
C647 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C648 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C649 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_3994_9798# 4.52e-20
C650 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C651 CLK_div_3_mag_0.JK_FF_mag_1.QB a_7421_10895# 0.00964f
C652 a_15078_10895# a_15238_10895# 0.0504f
C653 VDD a_10048_4717# 0.0132f
C654 a_13065_4717# a_13225_4717# 0.0504f
C655 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C656 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_7191_4717# 0.0731f
C657 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_13949_4717# 0.0733f
C658 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C659 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00229f
C660 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C661 CLK_div_10_mag_0.JK_FF_mag_2.QB a_10054_5814# 1.86e-20
C662 RST a_5122_9798# 5.71e-19
C663 CLK_div_3_mag_1.JK_FF_mag_1.K a_10363_9798# 0.012f
C664 VDD a_10209_10895# 3.14e-19
C665 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.K 0.0871f
C666 CLK_div_10_mag_0.and2_mag_1.OUT a_13795_5858# 5.94e-20
C667 VDD a_8145_10895# 0.0012f
C668 RST CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0783f
C669 CLK_div_3_mag_1.Q0 CLK_div_10_mag_0.Q1 1.5e-20
C670 VDD a_11779_8699# 5.92e-19
C671 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C672 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_8703_9798# 0.00119f
C673 RST CLK_div_3_mag_1.JK_FF_mag_1.K 0.428f
C674 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_10_mag_0.Q3 2.77e-19
C675 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_13795_5858# 0.0697f
C676 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_13071_5814# 0.0203f
C677 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_11342_5858# 0.011f
C678 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C679 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C680 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.283f
C681 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_14964_7257# 9.02e-19
C682 VDD a_5852_10895# 0.00743f
C683 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C684 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C685 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_12055_9798# 0.0732f
C686 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C687 CLK_div_3_mag_0.JK_FF_mag_1.QB a_6857_10895# 0.0811f
C688 VDD a_9043_4761# 0.00152f
C689 VDD a_12215_9798# 2.21e-19
C690 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C691 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_7031_4717# 0.0202f
C692 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_13789_4717# 0.0203f
C693 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C694 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00125f
C695 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_12896_6955# 0.069f
C696 CLK_div_10_mag_0.JK_FF_mag_2.QB a_8889_5858# 0.0114f
C697 RST a_4558_9798# 5.16e-19
C698 VDD a_7985_10895# 9.82e-19
C699 CLK_div_10_mag_0.Q2 a_11928_6955# 0.0112f
C700 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_8139_9798# 1.43e-19
C701 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_4898_4717# 8.64e-19
C702 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.11e-20
C703 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_0.K 0.0685f
C704 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_10778_5858# 1.43e-19
C705 VDD a_14923_5858# 3.56e-19
C706 VDD a_5692_10895# 0.00305f
C707 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_11491_9798# 0.00378f
C708 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0836f
C709 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.398f
C710 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_10806_8231# 0.132f
C711 CLK_div_3_mag_0.or_2_mag_0.IN2 a_5410_8699# 7.48e-20
C712 VDD a_8479_4761# 0.00152f
C713 CLK_div_10_mag_0.Q2 a_12896_6955# 0.0096f
C714 RST CLK_div_10_mag_0.and2_mag_1.OUT 4.25e-20
C715 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C716 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.and2_mag_1.OUT 0.00132f
C717 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C718 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C719 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.152f
C720 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_13225_4717# 1.5e-20
C721 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_10932_4717# 8.64e-19
C722 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00393f
C723 CLK_div_10_mag_0.JK_FF_mag_2.QB a_8325_5858# 2.96e-19
C724 VDD a_7421_10895# 0.00149f
C725 RST a_3994_9798# 5.16e-19
C726 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C727 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_7575_9798# 0.011f
C728 CLK_div_10_mag_0.Q2 a_10960_6955# 0.00929f
C729 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C730 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_10214_5814# 0.00119f
C731 VDD a_14359_5858# 3.14e-19
C732 VDD a_5128_10895# 2.21e-19
C733 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C734 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0378f
C735 VDD CLK_div_10_mag_0.JK_FF_mag_3.QB 0.911f
C736 RST CLK_div_3_mag_0.JK_FF_mag_1.QB 0.771f
C737 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_4968_10895# 8.64e-19
C738 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C739 VDD CLK_div_10_mag_0.Q0 5.08f
C740 VDD a_7915_4717# 0.00101f
C741 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C742 CLK_div_10_mag_0.Q2 a_13789_4717# 3.6e-22
C743 VDD a_11491_9798# 3.14e-19
C744 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00137f
C745 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_13065_4717# 1.17e-20
C746 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.Q0 0.149f
C747 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C748 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00545f
C749 CLK_div_10_mag_0.JK_FF_mag_2.QB a_7761_5858# 3.25e-19
C750 CLK_div_3_mag_0.JK_FF_mag_1.K a_5128_10895# 0.00695f
C751 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.198f
C752 VDD a_6857_10895# 0.00149f
C753 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_7011_9798# 0.00118f
C754 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_7985_10895# 8.64e-19
C755 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.or_2_mag_0.IN2 3.81e-19
C756 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C757 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C758 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C759 VDD a_13795_5858# 3.14e-19
C760 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C761 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C762 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.08e-20
C763 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.4e-19
C764 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK 0.00254f
C765 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00543f
C766 a_14354_10895# a_14514_10895# 0.0504f
C767 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_8325_5858# 4.52e-20
C768 VDD a_7755_4717# 0.00123f
C769 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C770 VDD a_10927_9798# 3.14e-19
C771 CLK_div_10_mag_0.Q2 a_13225_4717# 1.86e-20
C772 CLK_div_10_mag_0.JK_FF_mag_2.QB a_7197_5814# 0.00392f
C773 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_13790_10895# 0.069f
C774 CLK_div_3_mag_0.JK_FF_mag_1.K a_4968_10895# 0.00696f
C775 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.999f
C776 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_13944_9798# 0.069f
C777 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C778 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 RST 0.169f
C779 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C780 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_10_mag_0.and2_mag_0.OUT 2.97e-20
C781 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.or_2_mag_0.IN2 0.00761f
C782 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C783 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C784 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_5846_9798# 0.0203f
C785 a_12061_10895# a_12221_10895# 0.0504f
C786 VDD a_4404_10895# 3.14e-19
C787 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C788 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0545f
C789 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_7761_5858# 0.0202f
C790 VDD a_7191_4717# 0.00863f
C791 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_12221_10895# 0.0202f
C792 CLK_div_10_mag_0.Q2 a_13065_4717# 2.55e-20
C793 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.23f
C794 VDD a_10363_9798# 3.56e-19
C795 VDD RST 3.32f
C796 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C797 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 6.22e-20
C798 VDD CLK_div_10_mag_0.Q3 1.18f
C799 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_13226_10895# 0.00372f
C800 CLK_div_3_mag_0.JK_FF_mag_1.K a_4404_10895# 0.00964f
C801 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_13380_9798# 0.00372f
C802 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C803 RST CLK_div_10_mag_0.CLK 5.44e-19
C804 VDD a_13071_5814# 2.21e-19
C805 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_5686_9798# 0.0732f
C806 CLK CLK_div_3_mag_1.JK_FF_mag_1.QB 0.362f
C807 VDD a_3840_10895# 3.14e-19
C808 CLK_div_10_mag_0.Q3 Vdiv90 0.247f
C809 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 0.103f
C810 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0838f
C811 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C812 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_0.OUT 0.00117f
C813 RST CLK_div_3_mag_0.JK_FF_mag_1.K 0.477f
C814 a_4014_4717# a_4174_4717# 0.0504f
C815 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_12061_10895# 0.0731f
C816 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C817 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.QB 1.96f
C818 VDD a_7031_4717# 0.0123f
C819 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.54e-21
C820 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C821 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.21f
C822 CLK_div_10_mag_0.Q2 a_12060_4761# 0.0157f
C823 a_11928_6955# CLK_div_10_mag_0.JK_FF_mag_3.QB 1.45e-20
C824 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C825 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C826 a_4020_5814# a_4180_5814# 0.0504f
C827 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C828 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C829 CLK_div_3_mag_0.JK_FF_mag_1.K a_3840_10895# 0.0811f
C830 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C831 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C832 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C833 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.Q0 0.00335f
C834 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C835 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.QB 0.0147f
C836 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_5122_9798# 0.00378f
C837 Vdiv90 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.1e-22
C838 VDD a_11906_5858# 3.56e-19
C839 CLK_div_10_mag_0.Q3 a_15124_7257# 0.019f
C840 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00586f
C841 RST CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 9.24e-20
C842 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C843 VDD a_6026_4761# 0.00152f
C844 CLK_div_10_mag_0.Q0 a_12896_6955# 0.01f
C845 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_11497_10895# 9.1e-19
C846 CLK CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.0983f
C847 CLK_div_10_mag_0.Q2 a_11496_4761# 0.00859f
C848 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.45e-22
C849 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.94e-19
C850 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.207f
C851 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C852 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0334f
C853 CLK_div_10_mag_0.Q3 a_15077_4761# 0.0157f
C854 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_10_mag_0.and2_mag_0.OUT 2.77e-19
C855 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C856 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C857 VDD a_11342_5858# 3.14e-19
C858 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C859 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C860 a_10363_9798# CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C861 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C862 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C863 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.QB 1.96f
C864 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0378f
C865 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_11337_10895# 2.88e-20
C866 VDD a_5462_4761# 0.00152f
C867 a_10772_4717# a_10932_4717# 0.0504f
C868 CLK_div_10_mag_0.Q2 a_10932_4717# 0.0101f
C869 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C870 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C871 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00157f
C872 RST CLK_div_10_mag_0.JK_FF_mag_1.QB 0.163f
C873 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C874 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_15077_4761# 0.00372f
C875 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.305f
C876 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.0758f
C877 CLK_div_10_mag_0.Q3 a_14513_4761# 0.00859f
C878 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00943f
C879 RST CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 3.84e-20
C880 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C881 CLK CLK_div_3_mag_1.JK_FF_mag_1.K 2.11f
C882 VDD a_10778_5858# 3.14e-19
C883 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 4.85e-20
C884 a_11337_10895# a_11497_10895# 0.0504f
C885 a_10960_6955# CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.38e-20
C886 RST a_5410_8699# 5e-19
C887 VDD a_4898_4717# 0.00101f
C888 CLK_div_10_mag_0.Q0 a_13225_4717# 0.00164f
C889 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0501f
C890 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_4744_5858# 0.00378f
C891 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_1.OUT 0.0693f
C892 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C893 CLK_div_10_mag_0.Q2 a_10772_4717# 0.0102f
C894 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C895 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.QB 7.08e-20
C896 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C897 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_7575_9798# 0.069f
C898 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.69e-19
C899 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C900 CLK_div_3_mag_1.JK_FF_mag_1.K a_8863_9798# 1.09e-20
C901 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_14513_4761# 0.069f
C902 VDD CLK_div_3_mag_1.or_2_mag_0.IN2 0.492f
C903 RST a_13949_4717# 0.00127f
C904 CLK_div_10_mag_0.Q3 a_13949_4717# 0.0101f
C905 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Q2 3.87e-19
C906 RST a_13944_9798# 3.62e-19
C907 CLK CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 3.42e-19
C908 VDD a_10214_5814# 2.66e-19
C909 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C910 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 8.58e-20
C911 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C912 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C913 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_10773_10895# 0.069f
C914 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 0.215f
C915 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.264f
C916 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C917 CLK_div_10_mag_0.JK_FF_mag_1.QB a_6026_4761# 0.0811f
C918 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_4180_5814# 0.0732f
C919 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_5308_5858# 0.0059f
C920 CLK_div_10_mag_0.Q0 a_13065_4717# 0.00117f
C921 CLK_div_10_mag_0.Q2 a_10208_4717# 0.00789f
C922 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.41e-20
C923 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C924 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_14508_9798# 0.0202f
C925 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_7011_9798# 0.00372f
C926 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C927 VDD CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.458f
C928 CLK_div_3_mag_1.JK_FF_mag_1.K a_8703_9798# 8.77e-21
C929 RST CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00365f
C930 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0759f
C931 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_9043_4761# 0.00372f
C932 RST a_13789_4717# 0.00169f
C933 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C934 CLK_div_10_mag_0.Q3 a_13789_4717# 0.0102f
C935 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_5122_9798# 0.0202f
C936 RST CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.177f
C937 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C938 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C939 RST a_13380_9798# 7.24e-19
C940 VDD a_10054_5814# 0.00746f
C941 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C942 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_10209_10895# 0.00372f
C943 a_8709_10895# a_8869_10895# 0.0504f
C944 CLK_div_10_mag_0.JK_FF_mag_3.QB a_12060_4761# 0.0811f
C945 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C946 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_4020_5814# 0.0203f
C947 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_4744_5858# 0.0697f
C948 CLK_div_10_mag_0.JK_FF_mag_1.QB a_5462_4761# 0.00964f
C949 CLK_div_10_mag_0.Q2 a_10048_4717# 0.00335f
C950 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.647f
C951 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_13944_9798# 4.52e-20
C952 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0286f
C953 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C954 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K 2.37f
C955 RST a_13225_4717# 0.00186f
C956 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C957 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_8479_4761# 0.069f
C958 CLK_div_10_mag_0.Q3 a_13225_4717# 0.00789f
C959 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_4558_9798# 4.52e-20
C960 a_11779_8699# CLK_div_10_mag_0.Q2 1.71e-20
C961 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C962 CLK_div_3_mag_0.Q0 a_5686_9798# 2.79e-20
C963 VDD a_8889_5858# 3.56e-19
C964 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_14359_5858# 4.52e-20
C965 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_5852_10895# 0.0202f
C966 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C967 CLK_div_10_mag_0.JK_FF_mag_3.QB a_11496_4761# 0.00964f
C968 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_10778_5858# 0.00378f
C969 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.or_2_mag_0.IN2 0.0445f
C970 CLK_div_10_mag_0.JK_FF_mag_1.QB a_4898_4717# 0.00696f
C971 a_10048_4717# a_10208_4717# 0.0504f
C972 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C973 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C974 CLK_div_3_mag_0.Q0 a_4437_8231# 0.0134f
C975 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 0.69f
C976 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C977 CLK CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C978 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_4437_8231# 3.25e-19
C979 VDD CLK_div_10_mag_0.and2_mag_0.OUT 1.01f
C980 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C981 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C982 RST a_13065_4717# 0.00186f
C983 CLK_div_10_mag_0.Q3 a_13065_4717# 0.00335f
C984 VDD a_8325_5858# 3.14e-19
C985 CLK_div_3_mag_0.JK_FF_mag_1.QB a_8703_9798# 0.00392f
C986 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_5462_4761# 0.00378f
C987 CLK_div_10_mag_0.and2_mag_0.OUT Vdiv90 0.119f
C988 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0573f
C989 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_5692_10895# 0.0731f
C990 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_13795_5858# 0.0202f
C991 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_10214_5814# 0.0732f
C992 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_11342_5858# 0.0059f
C993 CLK_div_10_mag_0.JK_FF_mag_3.QB a_10932_4717# 0.00696f
C994 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C995 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_15238_10895# 1.17e-20
C996 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.038f
C997 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C998 VDD CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.654f
C999 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C1000 CLK_div_10_mag_0.nor_3_mag_0.IN3 a_14923_5858# 2.1e-20
C1001 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_8889_5858# 0.00372f
C1002 RST a_14514_10895# 8.64e-19
C1003 RST a_12060_4761# 9.66e-19
C1004 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_0.K 0.125f
C1005 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C1006 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C1007 VDD CLK 2.39f
C1008 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_11496_4761# 0.00378f
C1009 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C1010 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C1011 VDD a_7761_5858# 3.14e-19
C1012 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_11928_6955# 5.1e-20
C1013 CLK_div_3_mag_0.JK_FF_mag_1.QB a_8139_9798# 3.33e-19
C1014 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4898_4717# 0.0733f
C1015 RST a_12221_10895# 0.0049f
C1016 CLK_div_10_mag_0.and2_mag_0.OUT a_15124_7257# 0.00894f
C1017 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C1018 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_5128_10895# 9.1e-19
C1019 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_10778_5858# 0.0697f
C1020 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.QB 1.96f
C1021 CLK_div_10_mag_0.JK_FF_mag_3.QB a_10772_4717# 0.00695f
C1022 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_10054_5814# 0.0203f
C1023 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1f
C1024 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.and2_mag_1.OUT 2.57e-20
C1025 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_15078_10895# 1.5e-20
C1026 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C1027 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.Q0 0.622f
C1028 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C1029 VDD a_8863_9798# 5.99e-19
C1030 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C1031 CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00264f
C1032 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C1033 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_8325_5858# 0.069f
C1034 RST a_14354_10895# 0.00151f
C1035 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C1036 CLK_div_10_mag_0.CLK CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.419f
C1037 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C1038 RST a_11496_4761# 9.41e-19
C1039 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.652f
C1040 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C1041 RST CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.255f
C1042 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C1043 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C1044 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 3.25e-20
C1045 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_10932_4717# 0.0733f
C1046 VDD a_7197_5814# 2.66e-19
C1047 CLK_div_3_mag_0.Q0 a_3994_9798# 0.069f
C1048 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_10960_6955# 0.069f
C1049 RST CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0172f
C1050 VDD CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C1051 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C1052 RST a_12061_10895# 0.00487f
C1053 CLK_div_3_mag_0.JK_FF_mag_1.K a_8863_9798# 8.64e-19
C1054 CLK_div_10_mag_0.and2_mag_0.OUT a_14964_7257# 0.0294f
C1055 CLK a_15232_9798# 0.0101f
C1056 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_4968_10895# 2.88e-20
C1057 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C1058 a_7985_10895# a_8145_10895# 0.0504f
C1059 CLK a_15124_7257# 5.07e-21
C1060 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C1061 VDD CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C1062 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.109f
C1063 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_14514_10895# 0.0203f
C1064 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.and2_mag_1.OUT 8.51e-22
C1065 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C1066 VDD a_8703_9798# 2.65e-19
C1067 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_7421_10895# 0.069f
C1068 RST a_13790_10895# 8.68e-19
C1069 RST a_10932_4717# 0.00186f
C1070 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00718f
C1071 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C1072 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C1073 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.36e-19
C1074 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1075 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0352f
C1076 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1077 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_10772_4717# 0.0203f
C1078 a_5692_10895# a_5852_10895# 0.0504f
C1079 VDD a_7037_5814# 3.78e-19
C1080 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C1081 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_10363_9798# 4.52e-20
C1082 CLK_div_3_mag_0.JK_FF_mag_1.QB a_7011_9798# 0.0112f
C1083 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C1084 CLK a_15072_9798# 0.00939f
C1085 CLK_div_10_mag_0.and2_mag_0.OUT a_11928_6955# 0.00138f
C1086 RST a_11497_10895# 0.00343f
C1087 RST CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0198f
C1088 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00157f
C1089 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_8479_4761# 0.0036f
C1090 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_14354_10895# 0.0733f
C1091 CLK CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 7.03e-21
C1092 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.23f
C1093 VDD CLK_div_10_mag_0.JK_FF_mag_2.K 1.65f
C1094 VDD CLK_div_3_mag_1.Q0 1.29f
C1095 VDD a_8139_9798# 3.14e-19
C1096 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_15072_9798# 0.00119f
C1097 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_6857_10895# 0.00372f
C1098 RST a_13226_10895# 0.00192f
C1099 CLK_div_10_mag_0.and2_mag_0.OUT a_12896_6955# 0.00138f
C1100 a_12055_9798# a_12215_9798# 0.0504f
C1101 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.112f
C1102 RST CLK_div_10_mag_0.Q2 0.105f
C1103 RST a_10772_4717# 0.00169f
C1104 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5686_9798# 0.00119f
C1105 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.Q2 9.83e-19
C1106 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_10208_4717# 1.5e-20
C1107 Vdiv90 CLK_div_10_mag_0.JK_FF_mag_2.K 4.19e-19
C1108 VDD a_5872_5858# 3.56e-19
C1109 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C1110 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.Q0 0.00335f
C1111 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.49e-19
C1112 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K 0.0463f
C1113 CLK a_14508_9798# 6.43e-21
C1114 CLK_div_10_mag_0.Q2 a_13071_5814# 6.36e-19
C1115 RST a_11337_10895# 0.00327f
C1116 RST a_8869_10895# 0.00446f
C1117 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C1118 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.Q3 0.00442f
C1119 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C1120 RST CLK_div_3_mag_0.or_2_mag_0.IN2 0.00103f
C1121 CLK a_11928_6955# 1.71e-20
C1122 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.21f
C1123 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C1124 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00337f
C1125 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_4437_8231# 1.4e-19
C1126 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_13790_10895# 0.00378f
C1127 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C1128 VDD a_7575_9798# 3.14e-19
C1129 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C1130 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_14508_9798# 1.43e-19
C1131 VDD CLK_div_10_mag_0.JK_FF_mag_0.K 0.497f
C1132 RST a_10208_4717# 0.00186f
C1133 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_5122_9798# 1.43e-19
C1134 VDD CLK_div_3_mag_0.Q0 1.27f
C1135 a_15124_7257# CLK_div_10_mag_0.JK_FF_mag_2.K 3.02e-19
C1136 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_10048_4717# 1.17e-20
C1137 VDD a_5308_5858# 3.14e-19
C1138 VDD CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.467f
C1139 CLK_div_10_mag_0.JK_FF_mag_1.QB a_7197_5814# 1.41e-20
C1140 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_14508_9798# 0.0697f
C1141 RST a_10773_10895# 0.00382f
C1142 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C1143 CLK_div_10_mag_0.Q2 a_11906_5858# 0.069f
C1144 CLK a_13944_9798# 6.06e-21
C1145 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C1146 RST a_8709_10895# 0.00446f
C1147 CLK_div_3_mag_0.Q0 CLK_div_10_mag_0.CLK 0.00887f
C1148 CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 7.14e-19
C1149 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C1150 CLK_div_10_mag_0.CLK CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1e-19
C1151 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C1152 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C1153 VDD a_7011_9798# 3.56e-19
C1154 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.37f
C1155 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_8139_9798# 0.0697f
C1156 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_13944_9798# 0.011f
C1157 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0686f
C1158 CLK_div_10_mag_0.JK_FF_mag_2.K a_15077_4761# 0.0811f
C1159 VDD CLK_div_10_mag_0.Q1 4.08f
C1160 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C1161 RST a_10048_4717# 0.00186f
C1162 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_12221_10895# 1.17e-20
C1163 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_4558_9798# 0.011f
C1164 a_14964_7257# CLK_div_10_mag_0.JK_FF_mag_2.K 9.21e-20
C1165 VDD a_4738_4717# 0.00123f
C1166 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 6.71e-19
C1167 VDD CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C1168 VDD a_4744_5858# 3.14e-19
C1169 CLK_div_10_mag_0.JK_FF_mag_1.QB a_7037_5814# 1.86e-20
C1170 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C1171 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_13944_9798# 0.0059f
C1172 CLK a_13380_9798# 9.45e-19
C1173 RST a_10209_10895# 0.00371f
C1174 RST a_8145_10895# 0.00311f
C1175 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C1176 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0615f
C1177 CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C1178 CLK_div_10_mag_0.CLK a_4744_5858# 6.43e-21
C1179 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_7191_4717# 1.46e-19
C1180 RST CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0495f
C1181 CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_10_mag_0.JK_FF_mag_2.K 6.05e-19
C1182 RST a_5852_10895# 0.00325f
C1183 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_7575_9798# 0.0059f
C1184 RST CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0677f
C1185 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_13380_9798# 0.00118f
C1186 CLK_div_10_mag_0.JK_FF_mag_2.K a_14513_4761# 0.00964f
C1187 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1f
C1188 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C1189 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C1190 RST a_9043_4761# 9.66e-19
C1191 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_12061_10895# 1.5e-20
C1192 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_3994_9798# 0.00118f
C1193 CLK a_15238_10895# 0.00117f
C1194 VDD a_4174_4717# 0.00892f
C1195 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C1196 RST a_12215_9798# 7.78e-19
C1197 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C1198 a_4968_10895# a_5128_10895# 0.0504f
C1199 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 0.0435f
C1200 VDD a_4180_5814# 2.66e-19
C1201 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C1202 CLK_div_10_mag_0.JK_FF_mag_1.QB a_5872_5858# 0.0114f
C1203 CLK_div_10_mag_0.Q0 a_13795_5858# 6.43e-21
C1204 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_8869_10895# 0.0202f
C1205 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.647f
C1206 CLK_div_10_mag_0.CLK a_4174_4717# 0.00164f
C1207 RST a_7985_10895# 0.00359f
C1208 CLK_div_10_mag_0.CLK a_4180_5814# 0.00939f
C1209 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C1210 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C1211 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C1212 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 7.08e-20
C1213 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C1214 CLK_div_10_mag_0.Q0 a_7755_4717# 3.6e-22
C1215 CLK_div_10_mag_0.Q3 a_14923_5858# 0.069f
C1216 a_7755_4717# a_7915_4717# 0.0504f
C1217 RST a_5692_10895# 0.00302f
C1218 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C1219 CLK_div_10_mag_0.JK_FF_mag_2.K a_13949_4717# 0.00696f
C1220 RST CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0106f
C1221 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_4437_8231# 0.132f
C1222 CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.25f
C1223 RST a_8479_4761# 9.41e-19
C1224 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_11497_10895# 0.0203f
C1225 VDD a_4014_4717# 0.0132f
C1226 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C1227 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_10_mag_0.Q2 3.27e-19
C1228 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C1229 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1230 CLK_div_10_mag_0.JK_FF_mag_3.QB a_13231_5814# 1.41e-20
C1231 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C1232 CLK a_15078_10895# 0.00164f
C1233 RST a_12055_9798# 6.43e-19
C1234 CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C1235 VDD a_4020_5814# 0.00752f
C1236 CLK_div_10_mag_0.JK_FF_mag_1.QB a_5308_5858# 2.96e-19
C1237 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_4404_10895# 0.069f
C1238 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_10932_4717# 2.88e-20
C1239 CLK_div_10_mag_0.Q0 a_13231_5814# 0.00939f
C1240 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_8709_10895# 0.0731f
C1241 CLK_div_10_mag_0.CLK a_4014_4717# 0.00117f
C1242 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.29e-19
C1243 CLK_div_10_mag_0.Q2 a_10214_5814# 2.79e-20
C1244 RST a_7421_10895# 0.00439f
C1245 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_10_mag_0.Q1 4.44e-20
C1246 CLK CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 5.57e-19
C1247 CLK_div_10_mag_0.CLK a_4020_5814# 0.0101f
C1248 a_14923_5858# CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C1249 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_15078_10895# 1.46e-19
C1250 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_15232_9798# 0.0203f
C1251 a_8889_5858# CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C1252 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_14923_5858# 0.00372f
C1253 CLK_div_10_mag_0.Q0 a_7191_4717# 0.00166f
C1254 RST CLK_div_10_mag_0.JK_FF_mag_3.QB 0.179f
C1255 a_5686_9798# a_5846_9798# 0.0504f
C1256 RST a_5128_10895# 0.00232f
C1257 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.11f
C1258 CLK_div_10_mag_0.JK_FF_mag_2.K a_13789_4717# 0.00695f
C1259 RST CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.027f
C1260 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_5410_8699# 0.069f
C1261 CLK_div_10_mag_0.JK_FF_mag_0.K a_12896_6955# 0.0027f
C1262 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.QB 3.28e-19
C1263 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C1264 CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0432f
C1265 RST CLK_div_10_mag_0.Q0 0.293f
C1266 RST a_7915_4717# 0.00186f
C1267 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C1268 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.322f
C1269 CLK_div_10_mag_0.Q3 CLK_div_10_mag_0.Q0 0.149f
C1270 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_11337_10895# 0.0733f
C1271 CLK_div_10_mag_0.JK_FF_mag_3.QB a_13071_5814# 1.86e-20
C1272 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.38e-19
C1273 CLK_div_10_mag_0.JK_FF_mag_1.QB a_4738_4717# 0.00695f
C1274 RST a_11491_9798# 3.71e-19
C1275 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1276 CLK_div_10_mag_0.Q1 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C1277 CLK_div_10_mag_0.JK_FF_mag_1.QB a_4744_5858# 3.33e-19
C1278 CLK_div_10_mag_0.Q2 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C1279 CLK_div_10_mag_0.Q0 a_13071_5814# 0.0101f
C1280 CLK_div_10_mag_0.Q1 a_11928_6955# 0.0084f
C1281 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_10772_4717# 9.1e-19
C1282 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_8145_10895# 9.1e-19
C1283 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_3840_10895# 0.00372f
C1284 RST a_6857_10895# 0.00379f
C1285 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_14513_4761# 0.0036f
C1286 CLK_div_3_mag_1.or_2_mag_0.IN2 a_10806_8231# 8.64e-19
C1287 CLK a_12221_10895# 0.00117f
C1288 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_15072_9798# 0.0732f
C1289 RST a_13795_5858# 2.78e-19
C1290 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_14359_5858# 0.069f
C1291 CLK_div_10_mag_0.Q0 a_7031_4717# 0.001f
C1292 RST a_4968_10895# 0.00221f
C1293 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_5308_5858# 4.52e-20
C1294 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C1295 CLK_div_10_mag_0.Q0 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C1296 RST a_7755_4717# 0.00169f
C1297 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_10773_10895# 0.00378f
C1298 CLK_div_10_mag_0.JK_FF_mag_3.QB a_11906_5858# 0.0114f
C1299 RST a_10927_9798# 3.96e-19
C1300 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C1301 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C1302 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_10208_4717# 0.0731f
C1303 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_7985_10895# 2.88e-20
C1304 CLK_div_10_mag_0.JK_FF_mag_1.QB a_4180_5814# 0.00392f
C1305 CLK_div_10_mag_0.Q0 a_11906_5858# 9.45e-19
C1306 CLK_div_10_mag_0.Q1 a_10960_6955# 0.0105f
C1307 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_4898_4717# 2.88e-20
C1308 a_3994_9798# CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C1309 CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C1310 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C1311 RST CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.266f
C1312 a_15077_4761# VSS 0.0675f
C1313 a_14513_4761# VSS 0.0676f
C1314 a_13949_4717# VSS 0.0343f
C1315 a_13789_4717# VSS 0.0881f
C1316 a_13225_4717# VSS 0.0343f
C1317 a_13065_4717# VSS 0.0881f
C1318 a_12060_4761# VSS 0.0675f
C1319 a_11496_4761# VSS 0.0676f
C1320 a_10932_4717# VSS 0.0343f
C1321 a_10772_4717# VSS 0.0881f
C1322 a_10208_4717# VSS 0.0343f
C1323 a_10048_4717# VSS 0.0881f
C1324 a_9043_4761# VSS 0.0675f
C1325 a_8479_4761# VSS 0.0676f
C1326 a_7915_4717# VSS 0.0343f
C1327 a_7755_4717# VSS 0.0881f
C1328 a_7191_4717# VSS 0.0343f
C1329 a_7031_4717# VSS 0.0881f
C1330 a_6026_4761# VSS 0.0675f
C1331 a_5462_4761# VSS 0.0676f
C1332 a_4898_4717# VSS 0.0343f
C1333 a_4738_4717# VSS 0.0881f
C1334 a_4174_4717# VSS 0.0343f
C1335 a_4014_4717# VSS 0.0881f
C1336 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C1337 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.521f
C1338 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.416f
C1339 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.541f
C1340 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.416f
C1341 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.541f
C1342 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.416f
C1343 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.541f
C1344 a_14923_5858# VSS 0.0676f
C1345 a_14359_5858# VSS 0.0676f
C1346 a_13795_5858# VSS 0.0676f
C1347 a_13231_5814# VSS 0.0343f
C1348 a_13071_5814# VSS 0.0881f
C1349 a_11906_5858# VSS 0.0676f
C1350 a_11342_5858# VSS 0.0676f
C1351 a_10778_5858# VSS 0.0676f
C1352 a_10214_5814# VSS 0.0343f
C1353 a_10054_5814# VSS 0.0881f
C1354 a_8889_5858# VSS 0.0676f
C1355 a_8325_5858# VSS 0.0676f
C1356 a_7761_5858# VSS 0.0676f
C1357 a_7197_5814# VSS 0.0343f
C1358 a_7037_5814# VSS 0.0881f
C1359 a_5872_5858# VSS 0.0676f
C1360 a_5308_5858# VSS 0.0676f
C1361 a_4744_5858# VSS 0.0676f
C1362 a_4180_5814# VSS 0.0343f
C1363 a_4020_5814# VSS 0.0881f
C1364 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C1365 CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.755f
C1366 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C1367 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.808f
C1368 CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1369 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.414f
C1370 CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.693f
C1371 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.726f
C1372 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.809f
C1373 CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C1374 CLK_div_10_mag_0.JK_FF_mag_3.QB VSS 0.877f
C1375 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C1376 CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.696f
C1377 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.725f
C1378 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.81f
C1379 CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.509f
C1380 CLK_div_10_mag_0.JK_FF_mag_2.QB VSS 0.879f
C1381 CLK_div_10_mag_0.JK_FF_mag_2.K VSS 3.14f
C1382 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1383 CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.91f
C1384 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C1385 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.811f
C1386 CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.511f
C1387 CLK_div_10_mag_0.JK_FF_mag_1.QB VSS 0.899f
C1388 a_12896_6955# VSS 0.0679f
C1389 Vdiv90 VSS 0.519f
C1390 a_15124_7257# VSS 0.0371f
C1391 a_14964_7257# VSS 0.038f
C1392 a_11928_6955# VSS 0.0679f
C1393 a_10960_6955# VSS 0.0676f
C1394 CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.669f
C1395 CLK_div_10_mag_0.and2_mag_1.OUT VSS 0.706f
C1396 CLK_div_10_mag_0.JK_FF_mag_0.K VSS 0.633f
C1397 CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.435f
C1398 CLK_div_10_mag_0.Q0 VSS 3.5f
C1399 CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C1400 CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C1401 CLK_div_10_mag_0.Q2 VSS 2.22f
C1402 CLK_div_10_mag_0.Q1 VSS 2.63f
C1403 CLK_div_10_mag_0.Q3 VSS 1.96f
C1404 CLK_div_10_mag_0.and2_mag_0.OUT VSS 0.758f
C1405 CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS 0.337f
C1406 a_10806_8231# VSS 0.0247f
C1407 a_11779_8699# VSS 0.0676f
C1408 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.434f
C1409 a_4437_8231# VSS 0.0259f
C1410 CLK_div_3_mag_1.or_2_mag_0.IN2 VSS 0.416f
C1411 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C1412 a_5410_8699# VSS 0.0676f
C1413 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.436f
C1414 CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.42f
C1415 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.606f
C1416 CLK_div_10_mag_0.CLK VSS 2.59f
C1417 a_15232_9798# VSS 0.0881f
C1418 a_15072_9798# VSS 0.0343f
C1419 a_14508_9798# VSS 0.0676f
C1420 a_13944_9798# VSS 0.0676f
C1421 a_13380_9798# VSS 0.0676f
C1422 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C1423 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1424 a_12215_9798# VSS 0.0881f
C1425 a_12055_9798# VSS 0.0343f
C1426 a_11491_9798# VSS 0.0676f
C1427 a_10927_9798# VSS 0.0676f
C1428 a_10363_9798# VSS 0.0676f
C1429 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1430 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1431 a_8863_9798# VSS 0.0881f
C1432 a_8703_9798# VSS 0.0343f
C1433 a_8139_9798# VSS 0.0676f
C1434 a_7575_9798# VSS 0.0676f
C1435 a_7011_9798# VSS 0.0676f
C1436 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C1437 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1438 a_5846_9798# VSS 0.0881f
C1439 a_5686_9798# VSS 0.0343f
C1440 a_5122_9798# VSS 0.0676f
C1441 a_4558_9798# VSS 0.0676f
C1442 a_3994_9798# VSS 0.0676f
C1443 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1444 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1445 a_15238_10895# VSS 0.0881f
C1446 a_15078_10895# VSS 0.0343f
C1447 a_14514_10895# VSS 0.0881f
C1448 a_14354_10895# VSS 0.0343f
C1449 a_13790_10895# VSS 0.0676f
C1450 a_13226_10895# VSS 0.0675f
C1451 CLK_div_3_mag_1.JK_FF_mag_1.QB VSS 0.859f
C1452 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C1453 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.697f
C1454 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C1455 a_12221_10895# VSS 0.0881f
C1456 a_12061_10895# VSS 0.0343f
C1457 a_11497_10895# VSS 0.0881f
C1458 a_11337_10895# VSS 0.0343f
C1459 a_10773_10895# VSS 0.0676f
C1460 a_10209_10895# VSS 0.0675f
C1461 CLK_div_3_mag_1.JK_FF_mag_1.K VSS 4.56f
C1462 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.81f
C1463 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C1464 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C1465 a_8869_10895# VSS 0.0881f
C1466 a_8709_10895# VSS 0.0343f
C1467 a_8145_10895# VSS 0.0881f
C1468 a_7985_10895# VSS 0.0343f
C1469 a_7421_10895# VSS 0.0676f
C1470 a_6857_10895# VSS 0.0675f
C1471 CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.859f
C1472 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C1473 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.7f
C1474 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C1475 a_5852_10895# VSS 0.0881f
C1476 a_5692_10895# VSS 0.0343f
C1477 a_5128_10895# VSS 0.0881f
C1478 a_4968_10895# VSS 0.0343f
C1479 a_4404_10895# VSS 0.0676f
C1480 a_3840_10895# VSS 0.0675f
C1481 CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.55f
C1482 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.81f
C1483 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C1484 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C1485 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C1486 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.725f
C1487 CLK VSS 2.78f
C1488 CLK_div_3_mag_1.Q0 VSS 2.64f
C1489 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.54f
C1490 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C1491 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C1492 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.725f
C1493 CLK_div_3_mag_0.Q0 VSS 2.77f
C1494 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.54f
C1495 RST VSS 7.89f
C1496 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C1497 VDD VSS 0.146p
C1498 CLK_div_10_mag_0.JK_FF_mag_2.K.n0 VSS 0.0877f
C1499 CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VSS 0.0189f
C1500 CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VSS 0.0237f
C1501 CLK_div_10_mag_0.JK_FF_mag_2.K.n1 VSS 0.0561f
C1502 CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VSS 0.0333f
C1503 CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VSS 0.0212f
C1504 CLK_div_10_mag_0.JK_FF_mag_2.K.n2 VSS 0.0588f
C1505 CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VSS 0.0306f
C1506 CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VSS 0.0235f
C1507 CLK_div_10_mag_0.JK_FF_mag_2.K.n3 VSS 0.0604f
C1508 CLK_div_10_mag_0.JK_FF_mag_2.K.n4 VSS 1.13f
C1509 CLK_div_10_mag_0.JK_FF_mag_2.K.n5 VSS 0.378f
C1510 CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VSS 0.0148f
C1511 CLK_div_10_mag_0.JK_FF_mag_2.K.n6 VSS 0.0148f
C1512 CLK_div_10_mag_0.JK_FF_mag_2.K.n7 VSS 0.0349f
C1513 CLK_div_3_mag_0.Q1.t1 VSS 0.021f
C1514 CLK_div_3_mag_0.Q1.t0 VSS 0.0173f
C1515 CLK_div_3_mag_0.Q1.n0 VSS 0.0173f
C1516 CLK_div_3_mag_0.Q1.n1 VSS 0.0415f
C1517 CLK_div_3_mag_0.Q1.t8 VSS 0.0276f
C1518 CLK_div_3_mag_0.Q1.t10 VSS 0.0221f
C1519 CLK_div_3_mag_0.Q1.n2 VSS 0.0625f
C1520 CLK_div_3_mag_0.Q1.t7 VSS 0.0277f
C1521 CLK_div_3_mag_0.Q1.t4 VSS 0.0355f
C1522 CLK_div_3_mag_0.Q1.n3 VSS 0.0706f
C1523 CLK_div_3_mag_0.Q1.n4 VSS 0.321f
C1524 CLK_div_3_mag_0.Q1.t9 VSS 0.0385f
C1525 CLK_div_3_mag_0.Q1.t6 VSS 0.0254f
C1526 CLK_div_3_mag_0.Q1.n5 VSS 0.0684f
C1527 CLK_div_3_mag_0.Q1.t5 VSS 0.0276f
C1528 CLK_div_3_mag_0.Q1.t3 VSS 0.0221f
C1529 CLK_div_3_mag_0.Q1.n6 VSS 0.0642f
C1530 CLK_div_3_mag_0.Q1.n7 VSS 0.505f
C1531 CLK_div_3_mag_0.Q1.n8 VSS 0.209f
C1532 RST.n0 VSS 0.105f
C1533 RST.n1 VSS 0.00173f
C1534 RST.n2 VSS 0.00162f
C1535 RST.t8 VSS 0.0133f
C1536 RST.n3 VSS 0.0122f
C1537 RST.n4 VSS 0.00469f
C1538 RST.t10 VSS 0.0211f
C1539 RST.n5 VSS 0.0259f
C1540 RST.n6 VSS 2.05e-19
C1541 RST.n7 VSS 0.00172f
C1542 RST.n8 VSS 0.0108f
C1543 RST.n9 VSS 0.00863f
C1544 RST.t4 VSS 0.014f
C1545 RST.t5 VSS 0.0212f
C1546 RST.n10 VSS 0.0375f
C1547 RST.n11 VSS 0.0202f
C1548 RST.t1 VSS 0.014f
C1549 RST.t3 VSS 0.0212f
C1550 RST.n12 VSS 0.0375f
C1551 RST.n13 VSS 0.204f
C1552 RST.n14 VSS 0.636f
C1553 RST.n15 VSS 0.397f
C1554 RST.t14 VSS 0.014f
C1555 RST.t15 VSS 0.0212f
C1556 RST.n16 VSS 0.0375f
C1557 RST.n17 VSS 0.0195f
C1558 RST.n18 VSS 0.754f
C1559 RST.n19 VSS 0.00219f
C1560 RST.n20 VSS 0.00657f
C1561 RST.t6 VSS 0.0212f
C1562 RST.t2 VSS 0.0139f
C1563 RST.n21 VSS 0.0374f
C1564 RST.n22 VSS 0.00488f
C1565 RST.n23 VSS 0.00175f
C1566 RST.n24 VSS 0.139f
C1567 RST.n25 VSS 0.0061f
C1568 RST.t12 VSS 0.0214f
C1569 RST.t9 VSS 0.0136f
C1570 RST.n26 VSS 0.0376f
C1571 RST.n27 VSS 0.00489f
C1572 RST.n28 VSS 0.00325f
C1573 RST.n29 VSS 0.00172f
C1574 RST.n30 VSS 0.0834f
C1575 RST.n31 VSS 0.978f
C1576 RST.n32 VSS 0.00219f
C1577 RST.n33 VSS 0.00657f
C1578 RST.t11 VSS 0.0212f
C1579 RST.t7 VSS 0.0139f
C1580 RST.n34 VSS 0.0374f
C1581 RST.n35 VSS 0.00488f
C1582 RST.n36 VSS 0.00175f
C1583 RST.n37 VSS 0.139f
C1584 RST.n38 VSS 0.859f
C1585 RST.n39 VSS 0.59f
C1586 RST.t13 VSS 0.0136f
C1587 RST.t0 VSS 0.0214f
C1588 RST.n40 VSS 0.0376f
C1589 RST.n41 VSS 0.00489f
C1590 RST.n42 VSS 0.00325f
C1591 RST.n43 VSS 0.00172f
C1592 RST.n44 VSS 0.0061f
C1593 RST.n45 VSS 0.0517f
C1594 RST.n46 VSS 0.278f
C1595 RST.n47 VSS 0.2f
C1596 RST.n48 VSS 0.00143f
C1597 RST.n49 VSS 0.038f
C1598 RST.n50 VSS 0.0141f
C1599 CLK.n0 VSS 0.0189f
C1600 CLK.t5 VSS 0.053f
C1601 CLK.t13 VSS 0.0349f
C1602 CLK.n1 VSS 0.0936f
C1603 CLK.n2 VSS 0.0122f
C1604 CLK.n3 VSS 0.00879f
C1605 CLK.n4 VSS 0.00434f
C1606 CLK.n5 VSS 0.00879f
C1607 CLK.n6 VSS 0.00439f
C1608 CLK.t11 VSS 0.053f
C1609 CLK.t10 VSS 0.0349f
C1610 CLK.n7 VSS 0.0936f
C1611 CLK.n8 VSS 0.0122f
C1612 CLK.n9 VSS 0.0173f
C1613 CLK.n10 VSS 0.176f
C1614 CLK.n11 VSS 0.173f
C1615 CLK.n12 VSS 0.101f
C1616 CLK.t7 VSS 0.053f
C1617 CLK.t2 VSS 0.0349f
C1618 CLK.n13 VSS 0.0936f
C1619 CLK.n14 VSS 0.0122f
C1620 CLK.n15 VSS 0.00879f
C1621 CLK.n16 VSS 0.00434f
C1622 CLK.t8 VSS 0.053f
C1623 CLK.t4 VSS 0.0349f
C1624 CLK.n17 VSS 0.0936f
C1625 CLK.n18 VSS 0.00879f
C1626 CLK.n19 VSS 0.00439f
C1627 CLK.n20 VSS 0.0122f
C1628 CLK.n21 VSS 0.0173f
C1629 CLK.n22 VSS 0.164f
C1630 CLK.t0 VSS 0.0275f
C1631 CLK.t3 VSS 0.0491f
C1632 CLK.n23 VSS 0.0935f
C1633 CLK.n24 VSS 0.3f
C1634 CLK.n25 VSS 0.36f
C1635 CLK.n26 VSS 0.0135f
C1636 CLK.n27 VSS 0.101f
C1637 CLK.n28 VSS 0.0189f
C1638 CLK.n29 VSS 0.0315f
C1639 CLK.t1 VSS 0.0437f
C1640 CLK.t9 VSS 0.0113f
C1641 CLK.n30 VSS 0.0724f
C1642 CLK.n31 VSS 0.0154f
C1643 CLK.n32 VSS 0.00535f
C1644 CLK.n33 VSS 0.0114f
C1645 CLK.n34 VSS 0.669f
C1646 CLK.n35 VSS 0.669f
C1647 CLK.n36 VSS 0.0114f
C1648 CLK.t6 VSS 0.0113f
C1649 CLK.t12 VSS 0.0437f
C1650 CLK.n37 VSS 0.0724f
C1651 CLK.n38 VSS 0.0154f
C1652 CLK.n39 VSS 0.00535f
C1653 CLK.n40 VSS 0.0148f
C1654 CLK_div_3_mag_0.CLK.n0 VSS 0.52f
C1655 CLK_div_3_mag_0.CLK.n1 VSS 0.328f
C1656 CLK_div_3_mag_0.CLK.n2 VSS 0.0208f
C1657 CLK_div_3_mag_0.CLK.n3 VSS 0.0494f
C1658 CLK_div_3_mag_0.CLK.n4 VSS 0.0494f
C1659 CLK_div_3_mag_0.CLK.t1 VSS 0.0172f
C1660 CLK_div_3_mag_0.CLK.t0 VSS 0.0571f
C1661 CLK_div_3_mag_0.CLK.n5 VSS 0.198f
C1662 CLK_div_3_mag_0.CLK.t13 VSS 0.0109f
C1663 CLK_div_3_mag_0.CLK.t8 VSS 0.042f
C1664 CLK_div_3_mag_0.CLK.n6 VSS 0.0697f
C1665 CLK_div_3_mag_0.CLK.t6 VSS 0.0509f
C1666 CLK_div_3_mag_0.CLK.t2 VSS 0.0335f
C1667 CLK_div_3_mag_0.CLK.n7 VSS 0.09f
C1668 CLK_div_3_mag_0.CLK.t3 VSS 0.0509f
C1669 CLK_div_3_mag_0.CLK.t14 VSS 0.0335f
C1670 CLK_div_3_mag_0.CLK.n8 VSS 0.09f
C1671 CLK_div_3_mag_0.CLK.t11 VSS 0.0509f
C1672 CLK_div_3_mag_0.CLK.t7 VSS 0.0335f
C1673 CLK_div_3_mag_0.CLK.n9 VSS 0.09f
C1674 CLK_div_3_mag_0.CLK.t4 VSS 0.0264f
C1675 CLK_div_3_mag_0.CLK.t5 VSS 0.0472f
C1676 CLK_div_3_mag_0.CLK.n10 VSS 0.0899f
C1677 CLK_div_3_mag_0.CLK.n11 VSS 0.288f
C1678 CLK_div_3_mag_0.CLK.t12 VSS 0.0509f
C1679 CLK_div_3_mag_0.CLK.t9 VSS 0.0335f
C1680 CLK_div_3_mag_0.CLK.n12 VSS 0.09f
C1681 CLK_div_3_mag_0.CLK.t10 VSS 0.042f
C1682 CLK_div_3_mag_0.CLK.t15 VSS 0.0109f
C1683 CLK_div_3_mag_0.CLK.n13 VSS 0.0697f
C1684 CLK_div_3_mag_0.CLK.n14 VSS 0.67f
C1685 CLK_div_3_mag_0.CLK.n15 VSS 0.671f
C1686 CLK_div_3_mag_1.Q1.t1 VSS 0.021f
C1687 CLK_div_3_mag_1.Q1.t2 VSS 0.0173f
C1688 CLK_div_3_mag_1.Q1.n0 VSS 0.0173f
C1689 CLK_div_3_mag_1.Q1.n1 VSS 0.0415f
C1690 CLK_div_3_mag_1.Q1.t5 VSS 0.0276f
C1691 CLK_div_3_mag_1.Q1.t6 VSS 0.0221f
C1692 CLK_div_3_mag_1.Q1.n2 VSS 0.0625f
C1693 CLK_div_3_mag_1.Q1.t4 VSS 0.0277f
C1694 CLK_div_3_mag_1.Q1.t10 VSS 0.0355f
C1695 CLK_div_3_mag_1.Q1.n3 VSS 0.0706f
C1696 CLK_div_3_mag_1.Q1.n4 VSS 0.321f
C1697 CLK_div_3_mag_1.Q1.t7 VSS 0.0385f
C1698 CLK_div_3_mag_1.Q1.t3 VSS 0.0254f
C1699 CLK_div_3_mag_1.Q1.n5 VSS 0.0684f
C1700 CLK_div_3_mag_1.Q1.t9 VSS 0.0276f
C1701 CLK_div_3_mag_1.Q1.t8 VSS 0.0221f
C1702 CLK_div_3_mag_1.Q1.n6 VSS 0.0642f
C1703 CLK_div_3_mag_1.Q1.n7 VSS 0.505f
C1704 CLK_div_3_mag_1.Q1.n8 VSS 0.209f
C1705 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.07f
C1706 CLK_div_3_mag_0.JK_FF_mag_1.K.t1 VSS 0.0344f
C1707 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.0344f
C1708 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.0734f
C1709 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0774f
C1710 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.0493f
C1711 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.137f
C1712 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0552f
C1713 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0708f
C1714 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.141f
C1715 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.055f
C1716 CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VSS 0.044f
C1717 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 0.131f
C1718 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 1.18f
C1719 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.215f
C1720 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 VSS 2.07f
C1721 CLK_div_3_mag_1.JK_FF_mag_1.K.t1 VSS 0.0344f
C1722 CLK_div_3_mag_1.JK_FF_mag_1.K.n1 VSS 0.0344f
C1723 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 VSS 0.0734f
C1724 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 VSS 0.0774f
C1725 CLK_div_3_mag_1.JK_FF_mag_1.K.t2 VSS 0.0493f
C1726 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 VSS 0.137f
C1727 CLK_div_3_mag_1.JK_FF_mag_1.K.t7 VSS 0.0552f
C1728 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 VSS 0.0708f
C1729 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 VSS 0.141f
C1730 CLK_div_3_mag_1.JK_FF_mag_1.K.t3 VSS 0.055f
C1731 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VSS 0.044f
C1732 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 VSS 0.131f
C1733 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 VSS 1.18f
C1734 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 VSS 0.215f
C1735 CLK_div_3_mag_1.Q0.t1 VSS 0.025f
C1736 CLK_div_3_mag_1.Q0.t0 VSS 0.0206f
C1737 CLK_div_3_mag_1.Q0.n0 VSS 0.0206f
C1738 CLK_div_3_mag_1.Q0.n1 VSS 0.0494f
C1739 CLK_div_3_mag_1.Q0.t8 VSS 0.0459f
C1740 CLK_div_3_mag_1.Q0.t7 VSS 0.0302f
C1741 CLK_div_3_mag_1.Q0.n2 VSS 0.0814f
C1742 CLK_div_3_mag_1.Q0.t4 VSS 0.0329f
C1743 CLK_div_3_mag_1.Q0.t3 VSS 0.0263f
C1744 CLK_div_3_mag_1.Q0.n3 VSS 0.0764f
C1745 CLK_div_3_mag_1.Q0.n4 VSS 0.606f
C1746 CLK_div_3_mag_1.Q0.t6 VSS 0.0641f
C1747 CLK_div_3_mag_1.Q0.t5 VSS 0.0199f
C1748 CLK_div_3_mag_1.Q0.n5 VSS 0.0675f
C1749 CLK_div_3_mag_1.Q0.n6 VSS 0.447f
C1750 VDD.n0 VSS 0.0795f
C1751 VDD.t346 VSS 0.0229f
C1752 VDD.t383 VSS 0.00597f
C1753 VDD.n1 VSS 0.109f
C1754 VDD.n2 VSS 0.0852f
C1755 VDD.n3 VSS 0.00589f
C1756 VDD.t367 VSS 0.071f
C1757 VDD.n4 VSS 0.0365f
C1758 VDD.t460 VSS 0.00588f
C1759 VDD.n5 VSS 0.00586f
C1760 VDD.n6 VSS 0.0141f
C1761 VDD.n7 VSS 0.0573f
C1762 VDD.t459 VSS 0.0463f
C1763 VDD.t292 VSS 0.0531f
C1764 VDD.n8 VSS 0.0426f
C1765 VDD.t440 VSS 0.0523f
C1766 VDD.n9 VSS 0.00586f
C1767 VDD.n10 VSS 0.173f
C1768 VDD.n11 VSS 0.0139f
C1769 VDD.t267 VSS 0.00589f
C1770 VDD.n12 VSS 0.163f
C1771 VDD.t97 VSS 0.0271f
C1772 VDD.n13 VSS 0.00588f
C1773 VDD.t315 VSS 0.00589f
C1774 VDD.n14 VSS 0.00588f
C1775 VDD.n15 VSS 0.0292f
C1776 VDD.t403 VSS 0.0619f
C1777 VDD.n16 VSS 0.00588f
C1778 VDD.t34 VSS 0.00586f
C1779 VDD.t434 VSS 0.00589f
C1780 VDD.n17 VSS 0.0278f
C1781 VDD.t33 VSS 0.052f
C1782 VDD.t30 VSS 0.0403f
C1783 VDD.t121 VSS 0.00242f
C1784 VDD.n18 VSS 0.00242f
C1785 VDD.n19 VSS 0.00529f
C1786 VDD.t195 VSS 0.00589f
C1787 VDD.n20 VSS 0.00588f
C1788 VDD.n21 VSS 0.0292f
C1789 VDD.t171 VSS 0.0778f
C1790 VDD.n22 VSS 0.00588f
C1791 VDD.t424 VSS 0.00589f
C1792 VDD.n23 VSS 0.00588f
C1793 VDD.n24 VSS 0.00588f
C1794 VDD.t105 VSS 0.0767f
C1795 VDD.n25 VSS 0.0365f
C1796 VDD.t193 VSS 0.00589f
C1797 VDD.n26 VSS 0.00588f
C1798 VDD.t192 VSS 0.071f
C1799 VDD.t168 VSS 0.0778f
C1800 VDD.n27 VSS 0.0365f
C1801 VDD.t182 VSS 0.00589f
C1802 VDD.t205 VSS 0.00242f
C1803 VDD.n28 VSS 0.00242f
C1804 VDD.n29 VSS 0.00529f
C1805 VDD.t181 VSS 0.071f
C1806 VDD.t204 VSS 0.0867f
C1807 VDD.t347 VSS 0.0403f
C1808 VDD.n30 VSS 0.0365f
C1809 VDD.t254 VSS 0.00589f
C1810 VDD.t103 VSS 0.00242f
C1811 VDD.n31 VSS 0.00242f
C1812 VDD.n32 VSS 0.00529f
C1813 VDD.t253 VSS 0.071f
C1814 VDD.t102 VSS 0.0867f
C1815 VDD.t41 VSS 0.0403f
C1816 VDD.t287 VSS 0.0708f
C1817 VDD.n33 VSS 0.0365f
C1818 VDD.t288 VSS 0.0055f
C1819 VDD.t286 VSS 0.00505f
C1820 VDD.t471 VSS 0.00383f
C1821 VDD.n34 VSS 0.00987f
C1822 VDD.n35 VSS 0.00175f
C1823 VDD.t262 VSS 0.00505f
C1824 VDD.t479 VSS 0.00383f
C1825 VDD.n36 VSS 0.00987f
C1826 VDD.n37 VSS 0.00232f
C1827 VDD.n38 VSS 0.0012f
C1828 VDD.n39 VSS 6.06e-19
C1829 VDD.n40 VSS 0.0054f
C1830 VDD.n41 VSS 5.82e-19
C1831 VDD.t259 VSS 0.00491f
C1832 VDD.n42 VSS 0.00484f
C1833 VDD.t482 VSS 0.00382f
C1834 VDD.n43 VSS 0.00164f
C1835 VDD.n44 VSS 0.00518f
C1836 VDD.n45 VSS 0.00178f
C1837 VDD.n46 VSS 0.00147f
C1838 VDD.t279 VSS 0.00502f
C1839 VDD.t473 VSS 0.00383f
C1840 VDD.n47 VSS 0.0099f
C1841 VDD.n48 VSS 0.00186f
C1842 VDD.n49 VSS 0.00157f
C1843 VDD.n50 VSS 6.06e-19
C1844 VDD.n51 VSS 0.0191f
C1845 VDD.n52 VSS 0.074f
C1846 VDD.n53 VSS 0.108f
C1847 VDD.t477 VSS 0.00391f
C1848 VDD.t268 VSS 0.00496f
C1849 VDD.n54 VSS 0.00988f
C1850 VDD.n55 VSS 0.0036f
C1851 VDD.n56 VSS 0.00147f
C1852 VDD.t478 VSS 0.00383f
C1853 VDD.t265 VSS 0.00502f
C1854 VDD.n57 VSS 0.0099f
C1855 VDD.n58 VSS 0.00193f
C1856 VDD.n59 VSS 0.00152f
C1857 VDD.n60 VSS 6.06e-19
C1858 VDD.n61 VSS 0.0191f
C1859 VDD.n62 VSS 0.0249f
C1860 VDD.n63 VSS 0.12f
C1861 VDD.n64 VSS 0.0504f
C1862 VDD.n65 VSS 5.72e-19
C1863 VDD.n66 VSS 0.00473f
C1864 VDD.n67 VSS 0.0137f
C1865 VDD.n68 VSS 0.0336f
C1866 VDD.n69 VSS 0.0335f
C1867 VDD.n70 VSS 0.0344f
C1868 VDD.n71 VSS 0.0183f
C1869 VDD.n72 VSS 0.0335f
C1870 VDD.n73 VSS 0.0343f
C1871 VDD.n74 VSS 0.0203f
C1872 VDD.n75 VSS 0.0292f
C1873 VDD.n76 VSS 0.0271f
C1874 VDD.n77 VSS 0.0203f
C1875 VDD.n78 VSS 0.0555f
C1876 VDD.n79 VSS 0.0631f
C1877 VDD.t430 VSS 0.0767f
C1878 VDD.t423 VSS 0.071f
C1879 VDD.n80 VSS 0.0365f
C1880 VDD.n81 VSS 0.0203f
C1881 VDD.n82 VSS 0.0271f
C1882 VDD.n83 VSS 0.0292f
C1883 VDD.t203 VSS 0.00589f
C1884 VDD.n84 VSS 0.0271f
C1885 VDD.n85 VSS 0.0203f
C1886 VDD.n86 VSS 0.0365f
C1887 VDD.t202 VSS 0.071f
C1888 VDD.t178 VSS 0.0778f
C1889 VDD.t120 VSS 0.0867f
C1890 VDD.t194 VSS 0.071f
C1891 VDD.n87 VSS 0.0365f
C1892 VDD.n88 VSS 0.0203f
C1893 VDD.n89 VSS 0.0257f
C1894 VDD.n90 VSS 0.0241f
C1895 VDD.n91 VSS 0.0183f
C1896 VDD.n92 VSS 0.0365f
C1897 VDD.t433 VSS 0.0403f
C1898 VDD.n93 VSS 0.0547f
C1899 VDD.n94 VSS 0.0185f
C1900 VDD.n95 VSS 0.00588f
C1901 VDD.t393 VSS 0.0767f
C1902 VDD.n96 VSS 0.0365f
C1903 VDD.t111 VSS 0.00589f
C1904 VDD.n97 VSS 0.00588f
C1905 VDD.t110 VSS 0.071f
C1906 VDD.t65 VSS 0.0778f
C1907 VDD.n98 VSS 0.0365f
C1908 VDD.t101 VSS 0.00589f
C1909 VDD.t317 VSS 0.00242f
C1910 VDD.n99 VSS 0.00242f
C1911 VDD.n100 VSS 0.00529f
C1912 VDD.t100 VSS 0.071f
C1913 VDD.t316 VSS 0.0867f
C1914 VDD.t352 VSS 0.0403f
C1915 VDD.n101 VSS 0.0365f
C1916 VDD.t188 VSS 0.00589f
C1917 VDD.t399 VSS 0.00242f
C1918 VDD.n102 VSS 0.00242f
C1919 VDD.n103 VSS 0.00529f
C1920 VDD.t187 VSS 0.071f
C1921 VDD.t398 VSS 0.0867f
C1922 VDD.t162 VSS 0.0403f
C1923 VDD.t269 VSS 0.0708f
C1924 VDD.n104 VSS 0.0365f
C1925 VDD.t270 VSS 0.00631f
C1926 VDD.n105 VSS 0.0453f
C1927 VDD.n106 VSS 0.0335f
C1928 VDD.n107 VSS 0.0344f
C1929 VDD.n108 VSS 0.0183f
C1930 VDD.n109 VSS 0.0335f
C1931 VDD.n110 VSS 0.0343f
C1932 VDD.n111 VSS 0.0203f
C1933 VDD.n112 VSS 0.0292f
C1934 VDD.n113 VSS 0.0271f
C1935 VDD.n114 VSS 0.0203f
C1936 VDD.n115 VSS 0.0522f
C1937 VDD.n116 VSS 0.0417f
C1938 VDD.n117 VSS 0.0299f
C1939 VDD.t296 VSS 0.00589f
C1940 VDD.n118 VSS 0.0271f
C1941 VDD.n119 VSS 0.0203f
C1942 VDD.n120 VSS 0.0315f
C1943 VDD.t295 VSS 0.0565f
C1944 VDD.t62 VSS 0.0619f
C1945 VDD.t314 VSS 0.0418f
C1946 VDD.n121 VSS 0.0315f
C1947 VDD.n122 VSS 0.0203f
C1948 VDD.n123 VSS 0.0271f
C1949 VDD.n124 VSS 0.0292f
C1950 VDD.t1 VSS 0.00589f
C1951 VDD.t407 VSS 0.00242f
C1952 VDD.n125 VSS 0.00242f
C1953 VDD.n126 VSS 0.00529f
C1954 VDD.n127 VSS 0.0241f
C1955 VDD.t151 VSS 0.00589f
C1956 VDD.n128 VSS 0.00588f
C1957 VDD.n129 VSS 0.0289f
C1958 VDD.t396 VSS 0.0403f
C1959 VDD.t397 VSS 0.00589f
C1960 VDD.n130 VSS 0.00588f
C1961 VDD.n131 VSS 0.0289f
C1962 VDD.t28 VSS 0.0403f
C1963 VDD.t29 VSS 0.00589f
C1964 VDD.n132 VSS 0.00588f
C1965 VDD.n133 VSS 0.0289f
C1966 VDD.t447 VSS 0.00586f
C1967 VDD.n134 VSS 0.0207f
C1968 VDD.t104 VSS 0.15f
C1969 VDD.t201 VSS 0.0477f
C1970 VDD.n135 VSS 0.0553f
C1971 VDD.t345 VSS 0.152f
C1972 VDD.n136 VSS 0.0713f
C1973 VDD.t185 VSS 0.0753f
C1974 VDD.t186 VSS 0.00586f
C1975 VDD.n137 VSS 0.0279f
C1976 VDD.t184 VSS 0.00597f
C1977 VDD.n138 VSS 0.032f
C1978 VDD.n139 VSS 0.0193f
C1979 VDD.n140 VSS 0.083f
C1980 VDD.t183 VSS 0.049f
C1981 VDD.t446 VSS 0.0832f
C1982 VDD.n141 VSS 0.0543f
C1983 VDD.t390 VSS 0.0464f
C1984 VDD.n142 VSS 0.0365f
C1985 VDD.n143 VSS 0.0206f
C1986 VDD.n144 VSS 0.0274f
C1987 VDD.t96 VSS 0.00586f
C1988 VDD.n145 VSS 0.0207f
C1989 VDD.t95 VSS 0.0522f
C1990 VDD.n146 VSS 0.0855f
C1991 VDD.t165 VSS 0.0464f
C1992 VDD.n147 VSS 0.0365f
C1993 VDD.n148 VSS 0.0206f
C1994 VDD.n149 VSS 0.0274f
C1995 VDD.t308 VSS 0.00586f
C1996 VDD.n150 VSS 0.0207f
C1997 VDD.t307 VSS 0.0522f
C1998 VDD.n151 VSS 0.0855f
C1999 VDD.t400 VSS 0.0464f
C2000 VDD.t150 VSS 0.0708f
C2001 VDD.n152 VSS 0.0365f
C2002 VDD.n153 VSS 0.0206f
C2003 VDD.n154 VSS 0.0741f
C2004 VDD.n155 VSS 0.0623f
C2005 VDD.n156 VSS 0.0193f
C2006 VDD.n157 VSS 0.0203f
C2007 VDD.n158 VSS 0.0315f
C2008 VDD.t0 VSS 0.0565f
C2009 VDD.t406 VSS 0.069f
C2010 VDD.t159 VSS 0.032f
C2011 VDD.n159 VSS 0.0315f
C2012 VDD.t266 VSS 0.032f
C2013 VDD.n160 VSS 0.0902f
C2014 VDD.t152 VSS 0.0649f
C2015 VDD.t153 VSS 0.00586f
C2016 VDD.t124 VSS 0.0619f
C2017 VDD.n161 VSS 0.0315f
C2018 VDD.t177 VSS 0.00589f
C2019 VDD.n162 VSS 0.00588f
C2020 VDD.t176 VSS 0.0565f
C2021 VDD.t127 VSS 0.0619f
C2022 VDD.n163 VSS 0.0315f
C2023 VDD.n164 VSS 0.123f
C2024 VDD.t79 VSS 0.00589f
C2025 VDD.n165 VSS 0.00588f
C2026 VDD.n166 VSS 0.0315f
C2027 VDD.n167 VSS 0.136f
C2028 VDD.n168 VSS 0.00597f
C2029 VDD.n169 VSS 0.107f
C2030 VDD.n170 VSS 0.0841f
C2031 VDD.n171 VSS 0.00588f
C2032 VDD.n172 VSS 0.00588f
C2033 VDD.t35 VSS 0.0767f
C2034 VDD.n173 VSS 0.0365f
C2035 VDD.t134 VSS 0.00589f
C2036 VDD.n174 VSS 0.00588f
C2037 VDD.t133 VSS 0.071f
C2038 VDD.t331 VSS 0.0778f
C2039 VDD.n175 VSS 0.0365f
C2040 VDD.t222 VSS 0.00589f
C2041 VDD.t69 VSS 0.00242f
C2042 VDD.n176 VSS 0.00242f
C2043 VDD.n177 VSS 0.00529f
C2044 VDD.t221 VSS 0.071f
C2045 VDD.t68 VSS 0.0867f
C2046 VDD.t90 VSS 0.0403f
C2047 VDD.n178 VSS 0.0365f
C2048 VDD.t298 VSS 0.00589f
C2049 VDD.t22 VSS 0.00242f
C2050 VDD.n179 VSS 0.00242f
C2051 VDD.n180 VSS 0.00529f
C2052 VDD.t297 VSS 0.071f
C2053 VDD.t21 VSS 0.0867f
C2054 VDD.t323 VSS 0.0403f
C2055 VDD.t260 VSS 0.0708f
C2056 VDD.n181 VSS 0.0365f
C2057 VDD.t261 VSS 0.00631f
C2058 VDD.n182 VSS 0.0453f
C2059 VDD.n183 VSS 0.0335f
C2060 VDD.n184 VSS 0.0344f
C2061 VDD.n185 VSS 0.0183f
C2062 VDD.n186 VSS 0.0335f
C2063 VDD.n187 VSS 0.0343f
C2064 VDD.n188 VSS 0.0203f
C2065 VDD.n189 VSS 0.0292f
C2066 VDD.n190 VSS 0.0271f
C2067 VDD.n191 VSS 0.0203f
C2068 VDD.n192 VSS 0.0522f
C2069 VDD.t24 VSS 0.00586f
C2070 VDD.t78 VSS 0.0418f
C2071 VDD.t196 VSS 0.0271f
C2072 VDD.n193 VSS 0.163f
C2073 VDD.t312 VSS 0.0565f
C2074 VDD.t122 VSS 0.069f
C2075 VDD.t38 VSS 0.032f
C2076 VDD.t123 VSS 0.00242f
C2077 VDD.n194 VSS 0.00242f
C2078 VDD.n195 VSS 0.00529f
C2079 VDD.n196 VSS 0.0241f
C2080 VDD.t119 VSS 0.00589f
C2081 VDD.n197 VSS 0.0192f
C2082 VDD.n198 VSS 0.0183f
C2083 VDD.n199 VSS 0.0315f
C2084 VDD.t118 VSS 0.032f
C2085 VDD.n200 VSS 0.0902f
C2086 VDD.t23 VSS 0.0649f
C2087 VDD.n201 VSS 0.0181f
C2088 VDD.n202 VSS 0.037f
C2089 VDD.n203 VSS 0.0427f
C2090 VDD.n204 VSS 0.0748f
C2091 VDD.n205 VSS 0.00589f
C2092 VDD.t137 VSS 0.071f
C2093 VDD.n206 VSS 0.0365f
C2094 VDD.t422 VSS 0.00588f
C2095 VDD.t71 VSS 0.00599f
C2096 VDD.n207 VSS 0.0984f
C2097 VDD.t421 VSS 0.0463f
C2098 VDD.t2 VSS 0.0531f
C2099 VDD.n208 VSS 0.0918f
C2100 VDD.n209 VSS 0.00739f
C2101 VDD.n210 VSS 0.0141f
C2102 VDD.n211 VSS 0.0196f
C2103 VDD.t109 VSS 0.00599f
C2104 VDD.n212 VSS 0.00588f
C2105 VDD.n213 VSS 0.0247f
C2106 VDD.t223 VSS 0.0271f
C2107 VDD.t84 VSS 0.00242f
C2108 VDD.n214 VSS 0.00242f
C2109 VDD.n215 VSS 0.00529f
C2110 VDD.n216 VSS 0.0241f
C2111 VDD.n217 VSS 0.0149f
C2112 VDD.t334 VSS 0.0619f
C2113 VDD.n218 VSS 0.00588f
C2114 VDD.t426 VSS 0.00589f
C2115 VDD.t80 VSS 0.0619f
C2116 VDD.t425 VSS 0.0565f
C2117 VDD.n219 VSS 0.0315f
C2118 VDD.n220 VSS 0.024f
C2119 VDD.n221 VSS 0.025f
C2120 VDD.n222 VSS 0.0292f
C2121 VDD.n223 VSS 0.0203f
C2122 VDD.n224 VSS 0.0315f
C2123 VDD.t70 VSS 0.0418f
C2124 VDD.n225 VSS 0.163f
C2125 VDD.n226 VSS 0.00586f
C2126 VDD.n227 VSS 0.0265f
C2127 VDD.t5 VSS 0.0501f
C2128 VDD.t55 VSS 0.0523f
C2129 VDD.n228 VSS 0.0605f
C2130 VDD.t54 VSS 0.0527f
C2131 VDD.n229 VSS 0.0355f
C2132 VDD.n230 VSS 0.0171f
C2133 VDD.n231 VSS 0.158f
C2134 VDD.t281 VSS 0.00599f
C2135 VDD.n232 VSS 0.128f
C2136 VDD.t330 VSS 0.00615f
C2137 VDD.t329 VSS 0.0649f
C2138 VDD.n233 VSS 0.0902f
C2139 VDD.t280 VSS 0.032f
C2140 VDD.n234 VSS 0.0315f
C2141 VDD.t326 VSS 0.032f
C2142 VDD.t83 VSS 0.069f
C2143 VDD.t108 VSS 0.0565f
C2144 VDD.n235 VSS 0.0315f
C2145 VDD.n236 VSS 0.0203f
C2146 VDD.n237 VSS 0.097f
C2147 VDD.n238 VSS 0.0918f
C2148 VDD.n239 VSS 0.0345f
C2149 VDD.n240 VSS 0.0295f
C2150 VDD.n241 VSS 0.0993f
C2151 VDD.n242 VSS 0.0349f
C2152 VDD.n243 VSS 0.0288f
C2153 VDD.n244 VSS 0.0322f
C2154 VDD.t146 VSS 0.00242f
C2155 VDD.n245 VSS 0.00242f
C2156 VDD.n246 VSS 0.00529f
C2157 VDD.n247 VSS 0.019f
C2158 VDD.n248 VSS 0.00589f
C2159 VDD.n249 VSS 0.0259f
C2160 VDD.t147 VSS 0.0521f
C2161 VDD.n250 VSS 0.00586f
C2162 VDD.t412 VSS 0.00588f
C2163 VDD.t239 VSS 0.0712f
C2164 VDD.n251 VSS 0.00589f
C2165 VDD.t356 VSS 0.00242f
C2166 VDD.n252 VSS 0.00242f
C2167 VDD.n253 VSS 0.00529f
C2168 VDD.n254 VSS 0.00589f
C2169 VDD.n255 VSS 0.0344f
C2170 VDD.t272 VSS 0.071f
C2171 VDD.n256 VSS 7.94e-19
C2172 VDD.t480 VSS 0.00383f
C2173 VDD.n257 VSS 0.00526f
C2174 VDD.t271 VSS 0.00495f
C2175 VDD.n258 VSS 0.00471f
C2176 VDD.t475 VSS 0.00383f
C2177 VDD.t275 VSS 0.00505f
C2178 VDD.n259 VSS 0.00987f
C2179 VDD.n260 VSS 0.0656f
C2180 VDD.n261 VSS 0.0644f
C2181 VDD.n262 VSS 0.00285f
C2182 VDD.n263 VSS 0.0055f
C2183 VDD.n264 VSS 0.0155f
C2184 VDD.t136 VSS 0.00242f
C2185 VDD.n265 VSS 0.00242f
C2186 VDD.n266 VSS 0.00529f
C2187 VDD.n267 VSS 0.0336f
C2188 VDD.n268 VSS 0.0336f
C2189 VDD.n269 VSS 0.0365f
C2190 VDD.t135 VSS 0.0401f
C2191 VDD.t299 VSS 0.0867f
C2192 VDD.t309 VSS 0.0712f
C2193 VDD.t236 VSS 0.0867f
C2194 VDD.t355 VSS 0.0401f
C2195 VDD.n270 VSS 0.0365f
C2196 VDD.n271 VSS 0.0182f
C2197 VDD.n272 VSS 0.0336f
C2198 VDD.n273 VSS 0.0343f
C2199 VDD.t229 VSS 0.00588f
C2200 VDD.n274 VSS 0.00589f
C2201 VDD.n275 VSS 0.0271f
C2202 VDD.n276 VSS 0.0292f
C2203 VDD.n277 VSS 0.0204f
C2204 VDD.n278 VSS 0.0365f
C2205 VDD.t228 VSS 0.0776f
C2206 VDD.t230 VSS 0.0712f
C2207 VDD.t411 VSS 0.0765f
C2208 VDD.n279 VSS 0.0365f
C2209 VDD.n280 VSS 0.0204f
C2210 VDD.n281 VSS 0.0521f
C2211 VDD.t303 VSS 0.00588f
C2212 VDD.t233 VSS 0.0712f
C2213 VDD.n282 VSS 0.00589f
C2214 VDD.t418 VSS 0.0404f
C2215 VDD.n283 VSS 0.00589f
C2216 VDD.n284 VSS 0.00614f
C2217 VDD.t142 VSS 0.0521f
C2218 VDD.n285 VSS 0.0547f
C2219 VDD.n286 VSS 0.0279f
C2220 VDD.t322 VSS 0.00242f
C2221 VDD.n287 VSS 0.00242f
C2222 VDD.n288 VSS 0.00541f
C2223 VDD.n289 VSS 0.141f
C2224 VDD.n290 VSS 0.00589f
C2225 VDD.n291 VSS 0.0257f
C2226 VDD.n292 VSS 0.104f
C2227 VDD.n293 VSS 0.0182f
C2228 VDD.n294 VSS 0.0365f
C2229 VDD.t321 VSS 0.0401f
C2230 VDD.t304 VSS 0.0867f
C2231 VDD.t427 VSS 0.0712f
C2232 VDD.t242 VSS 0.0776f
C2233 VDD.n295 VSS 0.0365f
C2234 VDD.n296 VSS 0.0177f
C2235 VDD.t243 VSS 0.00597f
C2236 VDD.n297 VSS 0.109f
C2237 VDD.n298 VSS 0.0181f
C2238 VDD.t227 VSS 0.00588f
C2239 VDD.n299 VSS 0.0229f
C2240 VDD.n300 VSS 0.0204f
C2241 VDD.n301 VSS 0.0365f
C2242 VDD.t226 VSS 0.0776f
C2243 VDD.t215 VSS 0.0712f
C2244 VDD.t302 VSS 0.0765f
C2245 VDD.n302 VSS 0.0365f
C2246 VDD.n303 VSS 0.0204f
C2247 VDD.n304 VSS 0.0299f
C2248 VDD.n305 VSS 0.0416f
C2249 VDD.n306 VSS 0.0185f
C2250 VDD.n307 VSS 0.0547f
C2251 VDD.t443 VSS 0.0404f
C2252 VDD.t340 VSS 0.0776f
C2253 VDD.n308 VSS 0.00589f
C2254 VDD.n309 VSS 0.0257f
C2255 VDD.t341 VSS 0.00588f
C2256 VDD.n310 VSS 0.00589f
C2257 VDD.t209 VSS 0.0712f
C2258 VDD.n311 VSS 0.0365f
C2259 VDD.t75 VSS 0.00588f
C2260 VDD.n312 VSS 0.00589f
C2261 VDD.t74 VSS 0.0776f
C2262 VDD.t212 VSS 0.0712f
C2263 VDD.t413 VSS 0.0765f
C2264 VDD.n313 VSS 0.0365f
C2265 VDD.t414 VSS 0.00588f
C2266 VDD.t50 VSS 0.00588f
C2267 VDD.t342 VSS 0.0712f
C2268 VDD.n314 VSS 0.00589f
C2269 VDD.t89 VSS 0.00242f
C2270 VDD.n315 VSS 0.00242f
C2271 VDD.n316 VSS 0.00529f
C2272 VDD.n317 VSS 0.00589f
C2273 VDD.n318 VSS 0.0344f
C2274 VDD.t276 VSS 0.071f
C2275 VDD.n319 VSS 0.00631f
C2276 VDD.t141 VSS 0.00242f
C2277 VDD.n320 VSS 0.00242f
C2278 VDD.n321 VSS 0.00529f
C2279 VDD.n322 VSS 0.0336f
C2280 VDD.n323 VSS 0.0454f
C2281 VDD.n324 VSS 0.0365f
C2282 VDD.t140 VSS 0.0401f
C2283 VDD.t51 VSS 0.0867f
C2284 VDD.t337 VSS 0.0712f
C2285 VDD.t206 VSS 0.0867f
C2286 VDD.t88 VSS 0.0401f
C2287 VDD.n325 VSS 0.0365f
C2288 VDD.n326 VSS 0.0182f
C2289 VDD.n327 VSS 0.0336f
C2290 VDD.n328 VSS 0.0343f
C2291 VDD.t73 VSS 0.00588f
C2292 VDD.n329 VSS 0.00589f
C2293 VDD.n330 VSS 0.0271f
C2294 VDD.n331 VSS 0.0292f
C2295 VDD.n332 VSS 0.0204f
C2296 VDD.n333 VSS 0.0365f
C2297 VDD.t72 VSS 0.0776f
C2298 VDD.t289 VSS 0.0712f
C2299 VDD.t49 VSS 0.0765f
C2300 VDD.n334 VSS 0.0365f
C2301 VDD.n335 VSS 0.0204f
C2302 VDD.n336 VSS 0.0554f
C2303 VDD.n337 VSS 0.063f
C2304 VDD.n338 VSS 0.0204f
C2305 VDD.n339 VSS 0.0271f
C2306 VDD.n340 VSS 0.0292f
C2307 VDD.n341 VSS 0.0204f
C2308 VDD.n342 VSS 0.0271f
C2309 VDD.n343 VSS 0.0292f
C2310 VDD.n344 VSS 0.0204f
C2311 VDD.n345 VSS 0.0365f
C2312 VDD.t408 VSS 0.0712f
C2313 VDD.t415 VSS 0.0867f
C2314 VDD.t145 VSS 0.0401f
C2315 VDD.n346 VSS 0.0365f
C2316 VDD.n347 VSS 0.0136f
C2317 VDD.n348 VSS 0.0459f
C2318 VDD.n349 VSS 0.0521f
C2319 VDD.n350 VSS 0.0964f
C2320 VDD.n351 VSS 0.166f
C2321 VDD.n352 VSS 0.143f
C2322 VDD.n353 VSS 0.126f
C2323 VDD.t313 VSS 0.00599f
C2324 VDD.n354 VSS 0.097f
C2325 VDD.n355 VSS 0.0203f
C2326 VDD.n356 VSS 0.0292f
C2327 VDD.n357 VSS 0.0264f
C2328 VDD.n358 VSS 0.0732f
C2329 VDD.n359 VSS 0.0203f
C2330 VDD.n360 VSS 0.0292f
C2331 VDD.n361 VSS 0.0271f
C2332 VDD.n362 VSS 0.0178f
C2333 VDD.n363 VSS 0.00598f
C2334 VDD.n364 VSS 0.102f
C2335 VDD.n365 VSS 0.00588f
C2336 VDD.t154 VSS 0.0767f
C2337 VDD.n366 VSS 0.0365f
C2338 VDD.t175 VSS 0.00589f
C2339 VDD.n367 VSS 0.00588f
C2340 VDD.t174 VSS 0.071f
C2341 VDD.t130 VSS 0.0778f
C2342 VDD.n368 VSS 0.0365f
C2343 VDD.t200 VSS 0.00589f
C2344 VDD.t77 VSS 0.00242f
C2345 VDD.n369 VSS 0.00242f
C2346 VDD.n370 VSS 0.00529f
C2347 VDD.t199 VSS 0.071f
C2348 VDD.t76 VSS 0.0867f
C2349 VDD.t357 VSS 0.0403f
C2350 VDD.n371 VSS 0.0365f
C2351 VDD.t94 VSS 0.00589f
C2352 VDD.t158 VSS 0.00242f
C2353 VDD.n372 VSS 0.00242f
C2354 VDD.n373 VSS 0.00529f
C2355 VDD.t93 VSS 0.071f
C2356 VDD.t157 VSS 0.0867f
C2357 VDD.t25 VSS 0.0403f
C2358 VDD.t263 VSS 0.0708f
C2359 VDD.n374 VSS 0.0365f
C2360 VDD.t264 VSS 0.00631f
C2361 VDD.n375 VSS 0.0453f
C2362 VDD.n376 VSS 0.0335f
C2363 VDD.n377 VSS 0.0344f
C2364 VDD.n378 VSS 0.0183f
C2365 VDD.n379 VSS 0.0335f
C2366 VDD.n380 VSS 0.0343f
C2367 VDD.n381 VSS 0.0203f
C2368 VDD.n382 VSS 0.0292f
C2369 VDD.n383 VSS 0.0271f
C2370 VDD.n384 VSS 0.0203f
C2371 VDD.n385 VSS 0.0522f
C2372 VDD.n386 VSS 0.0349f
C2373 VDD.n387 VSS 0.0185f
C2374 VDD.n388 VSS 0.0259f
C2375 VDD.n389 VSS 0.0733f
C2376 VDD.n390 VSS 0.172f
C2377 VDD.n391 VSS 0.0722f
C2378 VDD.n392 VSS 0.0192f
C2379 VDD.n393 VSS 0.0605f
C2380 VDD.t114 VSS 0.0527f
C2381 VDD.n394 VSS 0.0355f
C2382 VDD.t218 VSS 0.0501f
C2383 VDD.n395 VSS 0.0918f
C2384 VDD.n396 VSS 0.0397f
C2385 VDD.n397 VSS 0.0467f
C2386 VDD.n398 VSS 0.0288f
C2387 VDD.n399 VSS 0.0443f
C2388 VDD.n400 VSS 0.0847f
C2389 VDD.t462 VSS 0.00588f
C2390 VDD.t384 VSS 0.0712f
C2391 VDD.n401 VSS 0.00589f
C2392 VDD.t351 VSS 0.00242f
C2393 VDD.n402 VSS 0.00242f
C2394 VDD.n403 VSS 0.00529f
C2395 VDD.n404 VSS 0.00589f
C2396 VDD.n405 VSS 0.0344f
C2397 VDD.t283 VSS 0.071f
C2398 VDD.n406 VSS 5.83e-19
C2399 VDD.t469 VSS 0.00383f
C2400 VDD.t255 VSS 0.00505f
C2401 VDD.n407 VSS 0.00987f
C2402 VDD.n408 VSS 0.0656f
C2403 VDD.n409 VSS 0.0648f
C2404 VDD.t474 VSS 0.00383f
C2405 VDD.t282 VSS 0.00495f
C2406 VDD.n410 VSS 0.00471f
C2407 VDD.n411 VSS 0.00526f
C2408 VDD.n412 VSS 8.32e-19
C2409 VDD.n413 VSS 0.0044f
C2410 VDD.n414 VSS 0.0055f
C2411 VDD.n415 VSS 0.0138f
C2412 VDD.t373 VSS 0.00242f
C2413 VDD.n416 VSS 0.00242f
C2414 VDD.n417 VSS 0.00529f
C2415 VDD.n418 VSS 0.0336f
C2416 VDD.n419 VSS 0.0336f
C2417 VDD.n420 VSS 0.0365f
C2418 VDD.t372 VSS 0.0401f
C2419 VDD.t456 VSS 0.0867f
C2420 VDD.t318 VSS 0.0712f
C2421 VDD.t247 VSS 0.0867f
C2422 VDD.t350 VSS 0.0401f
C2423 VDD.n421 VSS 0.0365f
C2424 VDD.n422 VSS 0.0182f
C2425 VDD.n423 VSS 0.0336f
C2426 VDD.n424 VSS 0.0343f
C2427 VDD.t17 VSS 0.00588f
C2428 VDD.n425 VSS 0.00589f
C2429 VDD.n426 VSS 0.0271f
C2430 VDD.n427 VSS 0.0292f
C2431 VDD.n428 VSS 0.0204f
C2432 VDD.n429 VSS 0.0365f
C2433 VDD.t16 VSS 0.0776f
C2434 VDD.t387 VSS 0.0712f
C2435 VDD.t461 VSS 0.0765f
C2436 VDD.n430 VSS 0.0365f
C2437 VDD.n431 VSS 0.0204f
C2438 VDD.n432 VSS 0.0508f
C2439 VDD.t45 VSS 0.00588f
C2440 VDD.n433 VSS 0.00589f
C2441 VDD.n434 VSS 0.022f
C2442 VDD.t85 VSS 0.0712f
C2443 VDD.n435 VSS 0.00589f
C2444 VDD.n436 VSS 0.00589f
C2445 VDD.n437 VSS 0.0279f
C2446 VDD.t448 VSS 0.0521f
C2447 VDD.n438 VSS 0.00614f
C2448 VDD.n439 VSS 0.0547f
C2449 VDD.t377 VSS 0.0404f
C2450 VDD.t46 VSS 0.0867f
C2451 VDD.t451 VSS 0.0401f
C2452 VDD.n440 VSS 0.0365f
C2453 VDD.n441 VSS 0.0182f
C2454 VDD.t452 VSS 0.00242f
C2455 VDD.n442 VSS 0.00242f
C2456 VDD.n443 VSS 0.00541f
C2457 VDD.n444 VSS 0.105f
C2458 VDD.n445 VSS 0.0257f
C2459 VDD.n446 VSS 0.0163f
C2460 VDD.n447 VSS 0.0365f
C2461 VDD.t382 VSS 0.0776f
C2462 VDD.t244 VSS 0.0712f
C2463 VDD.n448 VSS 0.00589f
C2464 VDD.n449 VSS 0.0194f
C2465 VDD.t15 VSS 0.00588f
C2466 VDD.n450 VSS 0.0234f
C2467 VDD.n451 VSS 0.0204f
C2468 VDD.n452 VSS 0.0365f
C2469 VDD.t14 VSS 0.0776f
C2470 VDD.t189 VSS 0.0712f
C2471 VDD.t44 VSS 0.0765f
C2472 VDD.n453 VSS 0.0365f
C2473 VDD.n454 VSS 0.0204f
C2474 VDD.n455 VSS 0.0284f
C2475 VDD.n456 VSS 0.0414f
C2476 VDD.n457 VSS 0.00586f
C2477 VDD.n458 VSS 0.00589f
C2478 VDD.n459 VSS 0.0259f
C2479 VDD.t362 VSS 0.0521f
C2480 VDD.n460 VSS 0.0136f
C2481 VDD.t438 VSS 0.0776f
C2482 VDD.n461 VSS 0.00589f
C2483 VDD.t366 VSS 0.00242f
C2484 VDD.n462 VSS 0.00242f
C2485 VDD.n463 VSS 0.00529f
C2486 VDD.n464 VSS 0.0459f
C2487 VDD.n465 VSS 0.019f
C2488 VDD.n466 VSS 0.0257f
C2489 VDD.t439 VSS 0.00588f
C2490 VDD.n467 VSS 0.00589f
C2491 VDD.t11 VSS 0.0712f
C2492 VDD.n468 VSS 0.0365f
C2493 VDD.t61 VSS 0.00588f
C2494 VDD.n469 VSS 0.00589f
C2495 VDD.t60 VSS 0.0776f
C2496 VDD.t18 VSS 0.0712f
C2497 VDD.t380 VSS 0.0765f
C2498 VDD.n470 VSS 0.0365f
C2499 VDD.t381 VSS 0.00588f
C2500 VDD.t113 VSS 0.00588f
C2501 VDD.t435 VSS 0.0712f
C2502 VDD.n471 VSS 0.00589f
C2503 VDD.t361 VSS 0.00242f
C2504 VDD.n472 VSS 0.00242f
C2505 VDD.n473 VSS 0.00529f
C2506 VDD.n474 VSS 0.00589f
C2507 VDD.n475 VSS 0.0344f
C2508 VDD.t256 VSS 0.071f
C2509 VDD.n476 VSS 0.00631f
C2510 VDD.t371 VSS 0.00242f
C2511 VDD.n477 VSS 0.00242f
C2512 VDD.n478 VSS 0.00529f
C2513 VDD.n479 VSS 0.0336f
C2514 VDD.n480 VSS 0.0454f
C2515 VDD.n481 VSS 0.0365f
C2516 VDD.t370 VSS 0.0401f
C2517 VDD.t115 VSS 0.0867f
C2518 VDD.t466 VSS 0.0712f
C2519 VDD.t8 VSS 0.0867f
C2520 VDD.t360 VSS 0.0401f
C2521 VDD.n482 VSS 0.0365f
C2522 VDD.n483 VSS 0.0182f
C2523 VDD.n484 VSS 0.0336f
C2524 VDD.n485 VSS 0.0343f
C2525 VDD.t59 VSS 0.00588f
C2526 VDD.n486 VSS 0.00589f
C2527 VDD.n487 VSS 0.0271f
C2528 VDD.n488 VSS 0.0292f
C2529 VDD.n489 VSS 0.0204f
C2530 VDD.n490 VSS 0.0365f
C2531 VDD.t58 VSS 0.0776f
C2532 VDD.t453 VSS 0.0712f
C2533 VDD.t112 VSS 0.0765f
C2534 VDD.n491 VSS 0.0365f
C2535 VDD.n492 VSS 0.0204f
C2536 VDD.n493 VSS 0.0554f
C2537 VDD.n494 VSS 0.063f
C2538 VDD.n495 VSS 0.0204f
C2539 VDD.n496 VSS 0.0271f
C2540 VDD.n497 VSS 0.0292f
C2541 VDD.n498 VSS 0.0204f
C2542 VDD.n499 VSS 0.0271f
C2543 VDD.n500 VSS 0.0292f
C2544 VDD.n501 VSS 0.0204f
C2545 VDD.n502 VSS 0.0365f
C2546 VDD.t250 VSS 0.0712f
C2547 VDD.t374 VSS 0.0867f
C2548 VDD.t365 VSS 0.0401f
C2549 VDD.n503 VSS 0.0365f
C2550 VDD.t463 VSS 0.0404f
C2551 VDD.n504 VSS 0.0547f
C2552 VDD.n505 VSS 0.0187f
C2553 VDD.n506 VSS 0.0842f
C2554 VDD.n507 VSS 0.184f
C2555 VDD.n508 VSS 0.183f
C2556 VDD.n509 VSS 0.149f
C2557 VDD.n510 VSS 0.0398f
C2558 VDD.n511 VSS 0.0484f
C2559 CLK_div_3_mag_0.Q0.t2 VSS 0.025f
C2560 CLK_div_3_mag_0.Q0.t0 VSS 0.0206f
C2561 CLK_div_3_mag_0.Q0.n0 VSS 0.0206f
C2562 CLK_div_3_mag_0.Q0.n1 VSS 0.0494f
C2563 CLK_div_3_mag_0.Q0.t5 VSS 0.0459f
C2564 CLK_div_3_mag_0.Q0.t4 VSS 0.0302f
C2565 CLK_div_3_mag_0.Q0.n2 VSS 0.0814f
C2566 CLK_div_3_mag_0.Q0.t7 VSS 0.0329f
C2567 CLK_div_3_mag_0.Q0.t6 VSS 0.0263f
C2568 CLK_div_3_mag_0.Q0.n3 VSS 0.0764f
C2569 CLK_div_3_mag_0.Q0.n4 VSS 0.606f
C2570 CLK_div_3_mag_0.Q0.t3 VSS 0.0641f
C2571 CLK_div_3_mag_0.Q0.t8 VSS 0.0199f
C2572 CLK_div_3_mag_0.Q0.n5 VSS 0.0675f
C2573 CLK_div_3_mag_0.Q0.n6 VSS 0.447f
.ends

