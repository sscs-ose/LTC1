** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/TG_TB.sch
**.subckt TG_TB
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
V3 IN VSS pulse(0 3.3 0 100p 100p 50u 100u)
.save i(v3)
V4 SEL VSS 0
.save i(v4)
x1 VDD SEL VSS OUT IN pex_TG
R1 OUT VSS 1k m=1
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_TG.spice
.control
save all

tran 100n 200u
plot v(OUT)
*************plot v(SEL)
plot v(IN)
*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
