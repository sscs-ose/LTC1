magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -28450 -15708 -4739 2632
<< metal1 >>
rect -23503 628 -22848 632
rect -23503 626 -13707 628
rect -10772 626 -9968 628
rect -23503 499 -9968 626
rect -23503 483 -16897 499
rect -23503 480 -23020 483
rect -23503 462 -23196 480
rect -23503 410 -23368 462
rect -23316 428 -23196 462
rect -23144 431 -23020 480
rect -22968 470 -16897 483
rect -22968 465 -19769 470
rect -22968 431 -21714 465
rect -23144 428 -21714 431
rect -23316 413 -21714 428
rect -21662 418 -19769 465
rect -19717 447 -16897 470
rect -16845 496 -9968 499
rect -16845 447 -16734 496
rect -19717 444 -16734 447
rect -16682 495 -9968 496
rect -16682 482 -10600 495
rect -16682 444 -16544 482
rect -19717 430 -16544 444
rect -16492 456 -10600 482
rect -16492 430 -13879 456
rect -19717 418 -13879 430
rect -21662 413 -13879 418
rect -23316 410 -13879 413
rect -23503 404 -13879 410
rect -13827 443 -10600 456
rect -10548 473 -9968 495
rect -10548 462 -10232 473
rect -10548 443 -10400 462
rect -13827 410 -10400 443
rect -10348 421 -10232 462
rect -10180 421 -9968 473
rect -10348 410 -9968 421
rect -13827 404 -9968 410
rect -23503 367 -9968 404
rect -23503 288 -22848 367
rect -23503 287 -23032 288
rect -23503 286 -23200 287
rect -23503 234 -23369 286
rect -23317 235 -23200 286
rect -23148 236 -23032 287
rect -22980 236 -22848 288
rect -23148 235 -22848 236
rect -23317 234 -22848 235
rect -23503 174 -22848 234
rect -21788 294 -21527 367
rect -21788 242 -21717 294
rect -21665 242 -21527 294
rect -21788 191 -21527 242
rect -19858 275 -19597 367
rect -19858 223 -19780 275
rect -19728 223 -19597 275
rect -19858 185 -19597 223
rect -16998 299 -16347 367
rect -16082 365 -9968 367
rect -16998 295 -16733 299
rect -16998 243 -16916 295
rect -16864 247 -16733 295
rect -16681 289 -16347 299
rect -16681 247 -16557 289
rect -16864 243 -16557 247
rect -16998 237 -16557 243
rect -16505 237 -16347 289
rect -16998 176 -16347 237
rect -13968 273 -13707 365
rect -13968 221 -13884 273
rect -13832 221 -13707 273
rect -13968 185 -13707 221
rect -10772 299 -9968 365
rect -10772 286 -10406 299
rect -10772 234 -10593 286
rect -10541 247 -10406 286
rect -10354 295 -9968 299
rect -10354 247 -10223 295
rect -10541 243 -10223 247
rect -10171 243 -9968 295
rect -10541 234 -9968 243
rect -10772 163 -9968 234
rect -13781 -13238 -13048 -13201
rect -13781 -13252 -13340 -13238
rect -13781 -13304 -13534 -13252
rect -13482 -13290 -13340 -13252
rect -13288 -13290 -13048 -13238
rect -13482 -13304 -13048 -13290
rect -13781 -13320 -13048 -13304
rect -20281 -13389 -19756 -13350
rect -13781 -13354 -13129 -13320
rect -20281 -13393 -19865 -13389
rect -20281 -13445 -20228 -13393
rect -20176 -13415 -19865 -13393
rect -20176 -13445 -20069 -13415
rect -20281 -13467 -20069 -13445
rect -20017 -13441 -19865 -13415
rect -19813 -13441 -19756 -13389
rect -20017 -13467 -19756 -13441
rect -20281 -13567 -19756 -13467
rect -17519 -13415 -17380 -13383
rect -17519 -13467 -17468 -13415
rect -17416 -13467 -17380 -13415
rect -17519 -13567 -17380 -13467
rect -15199 -13402 -15060 -13371
rect -15199 -13454 -15173 -13402
rect -15121 -13454 -15060 -13402
rect -15199 -13567 -15060 -13454
rect -13781 -13406 -13711 -13354
rect -13659 -13372 -13129 -13354
rect -13077 -13372 -13048 -13320
rect -13659 -13406 -13048 -13372
rect -13781 -13437 -13048 -13406
rect -13781 -13442 -13333 -13437
rect -13781 -13494 -13527 -13442
rect -13475 -13489 -13333 -13442
rect -13281 -13489 -13048 -13437
rect -13475 -13494 -13048 -13489
rect -13781 -13567 -13048 -13494
rect -12281 -13417 -12142 -13376
rect -12281 -13469 -12232 -13417
rect -12180 -13469 -12142 -13417
rect -12281 -13567 -12142 -13469
rect -8329 -13398 -7592 -13279
rect -8329 -13450 -8246 -13398
rect -8194 -13415 -7592 -13398
rect -8194 -13419 -7914 -13415
rect -8194 -13450 -8071 -13419
rect -8329 -13471 -8071 -13450
rect -8019 -13467 -7914 -13419
rect -7862 -13467 -7592 -13415
rect -8019 -13471 -7592 -13467
rect -8329 -13567 -7592 -13471
rect -20281 -13568 -7592 -13567
rect -20281 -13620 -20231 -13568
rect -20179 -13593 -7592 -13568
rect -20179 -13601 -19836 -13593
rect -20179 -13620 -20039 -13601
rect -20281 -13653 -20039 -13620
rect -19987 -13645 -19836 -13601
rect -19784 -13645 -8273 -13593
rect -8221 -13597 -7592 -13593
rect -8221 -13601 -7908 -13597
rect -8221 -13645 -8073 -13601
rect -19987 -13653 -8073 -13645
rect -8021 -13649 -7908 -13601
rect -7856 -13649 -7592 -13597
rect -8021 -13653 -7592 -13649
rect -20281 -13706 -7592 -13653
rect -20281 -13708 -19756 -13706
rect -8329 -13707 -7592 -13706
<< via1 >>
rect -23368 410 -23316 462
rect -23196 428 -23144 480
rect -23020 431 -22968 483
rect -21714 413 -21662 465
rect -19769 418 -19717 470
rect -16897 447 -16845 499
rect -16734 444 -16682 496
rect -16544 430 -16492 482
rect -13879 404 -13827 456
rect -10600 443 -10548 495
rect -10400 410 -10348 462
rect -10232 421 -10180 473
rect -23369 234 -23317 286
rect -23200 235 -23148 287
rect -23032 236 -22980 288
rect -21717 242 -21665 294
rect -19780 223 -19728 275
rect -16916 243 -16864 295
rect -16733 247 -16681 299
rect -16557 237 -16505 289
rect -13884 221 -13832 273
rect -10593 234 -10541 286
rect -10406 247 -10354 299
rect -10223 243 -10171 295
rect -13534 -13304 -13482 -13252
rect -13340 -13290 -13288 -13238
rect -20228 -13445 -20176 -13393
rect -20069 -13467 -20017 -13415
rect -19865 -13441 -19813 -13389
rect -17468 -13467 -17416 -13415
rect -15173 -13454 -15121 -13402
rect -13711 -13406 -13659 -13354
rect -13129 -13372 -13077 -13320
rect -13527 -13494 -13475 -13442
rect -13333 -13489 -13281 -13437
rect -12232 -13469 -12180 -13417
rect -8246 -13450 -8194 -13398
rect -8071 -13471 -8019 -13419
rect -7914 -13467 -7862 -13415
rect -20231 -13620 -20179 -13568
rect -20039 -13653 -19987 -13601
rect -19836 -13645 -19784 -13593
rect -8273 -13645 -8221 -13593
rect -8073 -13653 -8021 -13601
rect -7908 -13649 -7856 -13597
<< metal2 >>
rect -23503 486 -22848 632
rect -16998 502 -16347 628
rect -23503 483 -23022 486
rect -23503 465 -23198 483
rect -23503 409 -23370 465
rect -23314 427 -23198 465
rect -23142 430 -23022 483
rect -22966 430 -22848 486
rect -23142 427 -22848 430
rect -23314 409 -22848 427
rect -23503 291 -22848 409
rect -21737 468 -21637 495
rect -21737 412 -21716 468
rect -21660 412 -21637 468
rect -21737 389 -21637 412
rect -19792 473 -19692 500
rect -19792 417 -19771 473
rect -19715 417 -19692 473
rect -19792 394 -19692 417
rect -16998 446 -16899 502
rect -16843 499 -16347 502
rect -16843 446 -16736 499
rect -16998 443 -16736 446
rect -16680 485 -16347 499
rect -10772 498 -9968 628
rect -16680 443 -16546 485
rect -16998 429 -16546 443
rect -16490 429 -16347 485
rect -23503 290 -23034 291
rect -23503 289 -23202 290
rect -23503 233 -23371 289
rect -23315 234 -23202 289
rect -23146 235 -23034 290
rect -22978 235 -22848 291
rect -23146 234 -22848 235
rect -23315 233 -22848 234
rect -23503 174 -22848 233
rect -21740 297 -21640 324
rect -21740 241 -21719 297
rect -21663 241 -21640 297
rect -21740 218 -21640 241
rect -19803 278 -19703 305
rect -19803 222 -19782 278
rect -19726 222 -19703 278
rect -19803 199 -19703 222
rect -16998 302 -16347 429
rect -13902 459 -13802 486
rect -13902 403 -13881 459
rect -13825 403 -13802 459
rect -13902 380 -13802 403
rect -10772 442 -10602 498
rect -10546 476 -9968 498
rect -10546 465 -10234 476
rect -10546 442 -10402 465
rect -10772 409 -10402 442
rect -10346 420 -10234 465
rect -10178 420 -9968 476
rect -10346 409 -9968 420
rect -16998 298 -16735 302
rect -16998 242 -16918 298
rect -16862 246 -16735 298
rect -16679 292 -16347 302
rect -16679 246 -16559 292
rect -16862 242 -16559 246
rect -16998 236 -16559 242
rect -16503 236 -16347 292
rect -16998 176 -16347 236
rect -13907 276 -13807 303
rect -13907 220 -13886 276
rect -13830 220 -13807 276
rect -13907 198 -13807 220
rect -10772 302 -9968 409
rect -10772 289 -10408 302
rect -10772 233 -10595 289
rect -10539 246 -10408 289
rect -10352 298 -9968 302
rect -10352 246 -10225 298
rect -10539 242 -10225 246
rect -10169 242 -9968 298
rect -10539 233 -9968 242
rect -10772 163 -9968 233
rect -13781 -13235 -13048 -13201
rect -13781 -13249 -13342 -13235
rect -13781 -13305 -13536 -13249
rect -13480 -13291 -13342 -13249
rect -13286 -13291 -13048 -13235
rect -13480 -13305 -13048 -13291
rect -13781 -13317 -13048 -13305
rect -20281 -13386 -19756 -13350
rect -13781 -13351 -13131 -13317
rect -20281 -13390 -19867 -13386
rect -20281 -13446 -20230 -13390
rect -20174 -13412 -19867 -13390
rect -20174 -13446 -20071 -13412
rect -20281 -13468 -20071 -13446
rect -20015 -13442 -19867 -13412
rect -19811 -13442 -19756 -13386
rect -20015 -13468 -19756 -13442
rect -20281 -13565 -19756 -13468
rect -17491 -13412 -17391 -13385
rect -17491 -13468 -17470 -13412
rect -17414 -13468 -17391 -13412
rect -17491 -13490 -17391 -13468
rect -15196 -13399 -15096 -13372
rect -15196 -13455 -15175 -13399
rect -15119 -13455 -15096 -13399
rect -15196 -13477 -15096 -13455
rect -13781 -13407 -13713 -13351
rect -13657 -13373 -13131 -13351
rect -13075 -13373 -13048 -13317
rect -13657 -13407 -13048 -13373
rect -13781 -13434 -13048 -13407
rect -13781 -13439 -13335 -13434
rect -20281 -13621 -20233 -13565
rect -20177 -13590 -19756 -13565
rect -20177 -13598 -19838 -13590
rect -20177 -13621 -20041 -13598
rect -20281 -13654 -20041 -13621
rect -19985 -13646 -19838 -13598
rect -19782 -13646 -19756 -13590
rect -13781 -13495 -13529 -13439
rect -13473 -13490 -13335 -13439
rect -13279 -13490 -13048 -13434
rect -13473 -13495 -13048 -13490
rect -12255 -13414 -12155 -13387
rect -12255 -13470 -12234 -13414
rect -12178 -13470 -12155 -13414
rect -12255 -13492 -12155 -13470
rect -8329 -13395 -7592 -13279
rect -8329 -13451 -8248 -13395
rect -8192 -13412 -7592 -13395
rect -8192 -13416 -7916 -13412
rect -8192 -13451 -8073 -13416
rect -8329 -13472 -8073 -13451
rect -8017 -13468 -7916 -13416
rect -7860 -13468 -7592 -13412
rect -8017 -13472 -7592 -13468
rect -13781 -13635 -13048 -13495
rect -8329 -13590 -7592 -13472
rect -19985 -13654 -19756 -13646
rect -20281 -13708 -19756 -13654
rect -8329 -13646 -8275 -13590
rect -8219 -13594 -7592 -13590
rect -8219 -13598 -7910 -13594
rect -8219 -13646 -8075 -13598
rect -8329 -13654 -8075 -13646
rect -8019 -13650 -7910 -13598
rect -7854 -13650 -7592 -13594
rect -8019 -13654 -7592 -13650
rect -8329 -13707 -7592 -13654
<< via2 >>
rect -23022 483 -22966 486
rect -23198 480 -23142 483
rect -23370 462 -23314 465
rect -23370 410 -23368 462
rect -23368 410 -23316 462
rect -23316 410 -23314 462
rect -23198 428 -23196 480
rect -23196 428 -23144 480
rect -23144 428 -23142 480
rect -23022 431 -23020 483
rect -23020 431 -22968 483
rect -22968 431 -22966 483
rect -23022 430 -22966 431
rect -23198 427 -23142 428
rect -23370 409 -23314 410
rect -21716 465 -21660 468
rect -21716 413 -21714 465
rect -21714 413 -21662 465
rect -21662 413 -21660 465
rect -21716 412 -21660 413
rect -19771 470 -19715 473
rect -19771 418 -19769 470
rect -19769 418 -19717 470
rect -19717 418 -19715 470
rect -19771 417 -19715 418
rect -16899 499 -16843 502
rect -16899 447 -16897 499
rect -16897 447 -16845 499
rect -16845 447 -16843 499
rect -16899 446 -16843 447
rect -16736 496 -16680 499
rect -16736 444 -16734 496
rect -16734 444 -16682 496
rect -16682 444 -16680 496
rect -16736 443 -16680 444
rect -16546 482 -16490 485
rect -16546 430 -16544 482
rect -16544 430 -16492 482
rect -16492 430 -16490 482
rect -16546 429 -16490 430
rect -23371 286 -23315 289
rect -23371 234 -23369 286
rect -23369 234 -23317 286
rect -23317 234 -23315 286
rect -23202 287 -23146 290
rect -23202 235 -23200 287
rect -23200 235 -23148 287
rect -23148 235 -23146 287
rect -23034 288 -22978 291
rect -23034 236 -23032 288
rect -23032 236 -22980 288
rect -22980 236 -22978 288
rect -23034 235 -22978 236
rect -23202 234 -23146 235
rect -23371 233 -23315 234
rect -21719 294 -21663 297
rect -21719 242 -21717 294
rect -21717 242 -21665 294
rect -21665 242 -21663 294
rect -21719 241 -21663 242
rect -19782 275 -19726 278
rect -19782 223 -19780 275
rect -19780 223 -19728 275
rect -19728 223 -19726 275
rect -19782 222 -19726 223
rect -13881 456 -13825 459
rect -13881 404 -13879 456
rect -13879 404 -13827 456
rect -13827 404 -13825 456
rect -13881 403 -13825 404
rect -10602 495 -10546 498
rect -10602 443 -10600 495
rect -10600 443 -10548 495
rect -10548 443 -10546 495
rect -10234 473 -10178 476
rect -10602 442 -10546 443
rect -10402 462 -10346 465
rect -10402 410 -10400 462
rect -10400 410 -10348 462
rect -10348 410 -10346 462
rect -10234 421 -10232 473
rect -10232 421 -10180 473
rect -10180 421 -10178 473
rect -10234 420 -10178 421
rect -10402 409 -10346 410
rect -16735 299 -16679 302
rect -16918 295 -16862 298
rect -16918 243 -16916 295
rect -16916 243 -16864 295
rect -16864 243 -16862 295
rect -16735 247 -16733 299
rect -16733 247 -16681 299
rect -16681 247 -16679 299
rect -16735 246 -16679 247
rect -16559 289 -16503 292
rect -16918 242 -16862 243
rect -16559 237 -16557 289
rect -16557 237 -16505 289
rect -16505 237 -16503 289
rect -16559 236 -16503 237
rect -13886 273 -13830 276
rect -13886 221 -13884 273
rect -13884 221 -13832 273
rect -13832 221 -13830 273
rect -13886 220 -13830 221
rect -10408 299 -10352 302
rect -10595 286 -10539 289
rect -10595 234 -10593 286
rect -10593 234 -10541 286
rect -10541 234 -10539 286
rect -10408 247 -10406 299
rect -10406 247 -10354 299
rect -10354 247 -10352 299
rect -10408 246 -10352 247
rect -10225 295 -10169 298
rect -10225 243 -10223 295
rect -10223 243 -10171 295
rect -10171 243 -10169 295
rect -10225 242 -10169 243
rect -10595 233 -10539 234
rect -13342 -13238 -13286 -13235
rect -13536 -13252 -13480 -13249
rect -13536 -13304 -13534 -13252
rect -13534 -13304 -13482 -13252
rect -13482 -13304 -13480 -13252
rect -13342 -13290 -13340 -13238
rect -13340 -13290 -13288 -13238
rect -13288 -13290 -13286 -13238
rect -13342 -13291 -13286 -13290
rect -13536 -13305 -13480 -13304
rect -13131 -13320 -13075 -13317
rect -19867 -13389 -19811 -13386
rect -20230 -13393 -20174 -13390
rect -20230 -13445 -20228 -13393
rect -20228 -13445 -20176 -13393
rect -20176 -13445 -20174 -13393
rect -20230 -13446 -20174 -13445
rect -20071 -13415 -20015 -13412
rect -20071 -13467 -20069 -13415
rect -20069 -13467 -20017 -13415
rect -20017 -13467 -20015 -13415
rect -19867 -13441 -19865 -13389
rect -19865 -13441 -19813 -13389
rect -19813 -13441 -19811 -13389
rect -19867 -13442 -19811 -13441
rect -20071 -13468 -20015 -13467
rect -17470 -13415 -17414 -13412
rect -17470 -13467 -17468 -13415
rect -17468 -13467 -17416 -13415
rect -17416 -13467 -17414 -13415
rect -17470 -13468 -17414 -13467
rect -15175 -13402 -15119 -13399
rect -15175 -13454 -15173 -13402
rect -15173 -13454 -15121 -13402
rect -15121 -13454 -15119 -13402
rect -15175 -13455 -15119 -13454
rect -13713 -13354 -13657 -13351
rect -13713 -13406 -13711 -13354
rect -13711 -13406 -13659 -13354
rect -13659 -13406 -13657 -13354
rect -13131 -13372 -13129 -13320
rect -13129 -13372 -13077 -13320
rect -13077 -13372 -13075 -13320
rect -13131 -13373 -13075 -13372
rect -13713 -13407 -13657 -13406
rect -13335 -13437 -13279 -13434
rect -20233 -13568 -20177 -13565
rect -20233 -13620 -20231 -13568
rect -20231 -13620 -20179 -13568
rect -20179 -13620 -20177 -13568
rect -19838 -13593 -19782 -13590
rect -20233 -13621 -20177 -13620
rect -20041 -13601 -19985 -13598
rect -20041 -13653 -20039 -13601
rect -20039 -13653 -19987 -13601
rect -19987 -13653 -19985 -13601
rect -19838 -13645 -19836 -13593
rect -19836 -13645 -19784 -13593
rect -19784 -13645 -19782 -13593
rect -19838 -13646 -19782 -13645
rect -13529 -13442 -13473 -13439
rect -13529 -13494 -13527 -13442
rect -13527 -13494 -13475 -13442
rect -13475 -13494 -13473 -13442
rect -13335 -13489 -13333 -13437
rect -13333 -13489 -13281 -13437
rect -13281 -13489 -13279 -13437
rect -13335 -13490 -13279 -13489
rect -13529 -13495 -13473 -13494
rect -12234 -13417 -12178 -13414
rect -12234 -13469 -12232 -13417
rect -12232 -13469 -12180 -13417
rect -12180 -13469 -12178 -13417
rect -12234 -13470 -12178 -13469
rect -8248 -13398 -8192 -13395
rect -8248 -13450 -8246 -13398
rect -8246 -13450 -8194 -13398
rect -8194 -13450 -8192 -13398
rect -7916 -13415 -7860 -13412
rect -8248 -13451 -8192 -13450
rect -8073 -13419 -8017 -13416
rect -8073 -13471 -8071 -13419
rect -8071 -13471 -8019 -13419
rect -8019 -13471 -8017 -13419
rect -7916 -13467 -7914 -13415
rect -7914 -13467 -7862 -13415
rect -7862 -13467 -7860 -13415
rect -7916 -13468 -7860 -13467
rect -8073 -13472 -8017 -13471
rect -20041 -13654 -19985 -13653
rect -8275 -13593 -8219 -13590
rect -8275 -13645 -8273 -13593
rect -8273 -13645 -8221 -13593
rect -8221 -13645 -8219 -13593
rect -7910 -13597 -7854 -13594
rect -8275 -13646 -8219 -13645
rect -8075 -13601 -8019 -13598
rect -8075 -13653 -8073 -13601
rect -8073 -13653 -8021 -13601
rect -8021 -13653 -8019 -13601
rect -7910 -13649 -7908 -13597
rect -7908 -13649 -7856 -13597
rect -7856 -13649 -7854 -13597
rect -7910 -13650 -7854 -13649
rect -8075 -13654 -8019 -13653
<< metal3 >>
rect -23503 487 -22848 632
rect -16998 503 -16347 628
rect -23503 484 -23022 487
rect -23503 466 -23198 484
rect -23503 409 -23370 466
rect -23314 427 -23198 466
rect -23142 430 -23022 484
rect -22966 430 -22848 487
rect -23142 427 -22848 430
rect -23314 409 -22848 427
rect -23503 292 -22848 409
rect -21737 469 -21637 495
rect -21737 412 -21716 469
rect -21660 412 -21637 469
rect -21737 389 -21637 412
rect -19792 474 -19692 500
rect -19792 417 -19771 474
rect -19715 417 -19692 474
rect -19792 394 -19692 417
rect -16998 446 -16899 503
rect -16843 500 -16347 503
rect -16843 446 -16736 500
rect -16998 443 -16736 446
rect -16680 486 -16347 500
rect -10772 499 -9968 628
rect -16680 443 -16546 486
rect -16998 429 -16546 443
rect -16490 429 -16347 486
rect -23503 291 -23034 292
rect -23503 290 -23202 291
rect -23503 233 -23371 290
rect -23315 234 -23202 290
rect -23146 235 -23034 291
rect -22978 235 -22848 292
rect -23146 234 -22848 235
rect -23315 233 -22848 234
rect -23503 174 -22848 233
rect -21740 298 -21640 324
rect -21740 241 -21719 298
rect -21663 241 -21640 298
rect -21740 218 -21640 241
rect -19803 279 -19703 305
rect -19803 222 -19782 279
rect -19726 222 -19703 279
rect -19803 199 -19703 222
rect -16998 303 -16347 429
rect -13902 460 -13802 486
rect -13902 403 -13881 460
rect -13825 403 -13802 460
rect -13902 380 -13802 403
rect -10772 442 -10602 499
rect -10546 477 -9968 499
rect -10546 466 -10234 477
rect -10546 442 -10402 466
rect -10772 409 -10402 442
rect -10346 420 -10234 466
rect -10178 420 -9968 477
rect -10346 409 -9968 420
rect -10772 303 -9968 409
rect -16998 299 -16735 303
rect -16998 242 -16918 299
rect -16862 246 -16735 299
rect -16679 293 -16347 303
rect -16679 246 -16559 293
rect -16862 242 -16559 246
rect -16998 236 -16559 242
rect -16503 236 -16347 293
rect -16998 176 -16347 236
rect -13907 277 -13807 303
rect -13907 220 -13886 277
rect -13830 220 -13807 277
rect -13907 198 -13807 220
rect -10772 290 -10408 303
rect -10772 233 -10595 290
rect -10539 246 -10408 290
rect -10352 299 -9968 303
rect -10352 246 -10225 299
rect -10539 242 -10225 246
rect -10169 242 -9968 299
rect -10539 233 -9968 242
rect -10772 163 -9968 233
rect -13781 -13234 -13048 -13201
rect -13781 -13248 -13342 -13234
rect -13781 -13305 -13536 -13248
rect -13480 -13291 -13342 -13248
rect -13286 -13291 -13048 -13234
rect -13480 -13305 -13048 -13291
rect -13781 -13316 -13048 -13305
rect -13781 -13350 -13131 -13316
rect -20251 -13389 -20151 -13363
rect -19888 -13385 -19788 -13359
rect -20251 -13446 -20230 -13389
rect -20174 -13446 -20151 -13389
rect -20251 -13468 -20151 -13446
rect -20092 -13411 -19992 -13385
rect -20092 -13468 -20071 -13411
rect -20015 -13468 -19992 -13411
rect -19888 -13442 -19867 -13385
rect -19811 -13442 -19788 -13385
rect -19888 -13464 -19788 -13442
rect -17491 -13411 -17391 -13385
rect -20092 -13490 -19992 -13468
rect -17491 -13468 -17470 -13411
rect -17414 -13468 -17391 -13411
rect -17491 -13490 -17391 -13468
rect -15196 -13398 -15096 -13372
rect -15196 -13455 -15175 -13398
rect -15119 -13455 -15096 -13398
rect -15196 -13477 -15096 -13455
rect -13781 -13407 -13713 -13350
rect -13657 -13373 -13131 -13350
rect -13075 -13373 -13048 -13316
rect -13657 -13407 -13048 -13373
rect -13781 -13433 -13048 -13407
rect -13781 -13438 -13335 -13433
rect -13781 -13495 -13529 -13438
rect -13473 -13490 -13335 -13438
rect -13279 -13490 -13048 -13433
rect -13473 -13495 -13048 -13490
rect -12255 -13413 -12155 -13387
rect -12255 -13470 -12234 -13413
rect -12178 -13470 -12155 -13413
rect -12255 -13492 -12155 -13470
rect -8329 -13394 -7592 -13279
rect -8329 -13451 -8248 -13394
rect -8192 -13411 -7592 -13394
rect -8192 -13415 -7916 -13411
rect -8192 -13451 -8073 -13415
rect -8329 -13472 -8073 -13451
rect -8017 -13468 -7916 -13415
rect -7860 -13468 -7592 -13411
rect -8017 -13472 -7592 -13468
rect -20254 -13564 -20154 -13538
rect -20254 -13621 -20233 -13564
rect -20177 -13621 -20154 -13564
rect -20254 -13643 -20154 -13621
rect -20062 -13597 -19962 -13571
rect -20062 -13654 -20041 -13597
rect -19985 -13654 -19962 -13597
rect -20062 -13676 -19962 -13654
rect -19859 -13589 -19759 -13563
rect -19859 -13646 -19838 -13589
rect -19782 -13646 -19759 -13589
rect -13781 -13635 -13048 -13495
rect -8329 -13589 -7592 -13472
rect -19859 -13668 -19759 -13646
rect -8329 -13646 -8275 -13589
rect -8219 -13593 -7592 -13589
rect -8219 -13597 -7910 -13593
rect -8219 -13646 -8075 -13597
rect -8329 -13654 -8075 -13646
rect -8019 -13650 -7910 -13597
rect -7854 -13650 -7592 -13593
rect -8019 -13654 -7592 -13650
rect -8329 -13707 -7592 -13654
<< via3 >>
rect -23022 486 -22966 487
rect -23198 483 -23142 484
rect -23370 465 -23314 466
rect -23370 410 -23314 465
rect -23198 428 -23142 483
rect -23022 431 -22966 486
rect -21716 468 -21660 469
rect -21716 413 -21660 468
rect -19771 473 -19715 474
rect -19771 418 -19715 473
rect -16899 502 -16843 503
rect -16899 447 -16843 502
rect -16736 499 -16680 500
rect -16736 444 -16680 499
rect -16546 485 -16490 486
rect -16546 430 -16490 485
rect -23034 291 -22978 292
rect -23202 290 -23146 291
rect -23371 289 -23315 290
rect -23371 234 -23315 289
rect -23202 235 -23146 290
rect -23034 236 -22978 291
rect -21719 297 -21663 298
rect -21719 242 -21663 297
rect -19782 278 -19726 279
rect -19782 223 -19726 278
rect -13881 459 -13825 460
rect -13881 404 -13825 459
rect -10602 498 -10546 499
rect -10602 443 -10546 498
rect -10234 476 -10178 477
rect -10402 465 -10346 466
rect -10402 410 -10346 465
rect -10234 421 -10178 476
rect -16735 302 -16679 303
rect -16918 298 -16862 299
rect -16918 243 -16862 298
rect -16735 247 -16679 302
rect -16559 292 -16503 293
rect -16559 237 -16503 292
rect -13886 276 -13830 277
rect -13886 221 -13830 276
rect -10408 302 -10352 303
rect -10595 289 -10539 290
rect -10595 234 -10539 289
rect -10408 247 -10352 302
rect -10225 298 -10169 299
rect -10225 243 -10169 298
rect -13342 -13235 -13286 -13234
rect -13536 -13249 -13480 -13248
rect -13536 -13304 -13480 -13249
rect -13342 -13290 -13286 -13235
rect -13131 -13317 -13075 -13316
rect -20230 -13390 -20174 -13389
rect -20230 -13445 -20174 -13390
rect -20071 -13412 -20015 -13411
rect -20071 -13467 -20015 -13412
rect -19867 -13386 -19811 -13385
rect -19867 -13441 -19811 -13386
rect -17470 -13412 -17414 -13411
rect -17470 -13467 -17414 -13412
rect -15175 -13399 -15119 -13398
rect -15175 -13454 -15119 -13399
rect -13713 -13351 -13657 -13350
rect -13713 -13406 -13657 -13351
rect -13131 -13372 -13075 -13317
rect -13335 -13434 -13279 -13433
rect -13529 -13439 -13473 -13438
rect -13529 -13494 -13473 -13439
rect -13335 -13489 -13279 -13434
rect -12234 -13414 -12178 -13413
rect -12234 -13469 -12178 -13414
rect -8248 -13395 -8192 -13394
rect -8248 -13450 -8192 -13395
rect -7916 -13412 -7860 -13411
rect -8073 -13416 -8017 -13415
rect -8073 -13471 -8017 -13416
rect -7916 -13467 -7860 -13412
rect -20233 -13565 -20177 -13564
rect -20233 -13620 -20177 -13565
rect -20041 -13598 -19985 -13597
rect -20041 -13653 -19985 -13598
rect -19838 -13590 -19782 -13589
rect -19838 -13645 -19782 -13590
rect -8275 -13590 -8219 -13589
rect -8275 -13645 -8219 -13590
rect -7910 -13594 -7854 -13593
rect -8075 -13598 -8019 -13597
rect -8075 -13653 -8019 -13598
rect -7910 -13649 -7854 -13594
<< metal4 >>
rect -23503 489 -22848 632
rect -16998 505 -16347 628
rect -16998 503 -16898 505
rect -23503 487 -23021 489
rect -23503 486 -23022 487
rect -23503 484 -23197 486
rect -23503 468 -23198 484
rect -23503 466 -23369 468
rect -23503 410 -23370 466
rect -23313 428 -23198 468
rect -23141 431 -23022 486
rect -22965 433 -22848 489
rect -22966 431 -22848 433
rect -23141 430 -22848 431
rect -23142 428 -22848 430
rect -23313 412 -22848 428
rect -23314 410 -22848 412
rect -23503 294 -22848 410
rect -21737 471 -21637 495
rect -21737 469 -21715 471
rect -21737 413 -21716 469
rect -21659 415 -21637 471
rect -21660 413 -21637 415
rect -21737 389 -21637 413
rect -19792 476 -19692 500
rect -19792 474 -19770 476
rect -19792 418 -19771 474
rect -19714 420 -19692 476
rect -19715 418 -19692 420
rect -19792 394 -19692 418
rect -16998 447 -16899 503
rect -16842 502 -16347 505
rect -16842 500 -16735 502
rect -16842 449 -16736 500
rect -16843 447 -16736 449
rect -16998 444 -16736 447
rect -16679 488 -16347 502
rect -16679 486 -16545 488
rect -16679 446 -16546 486
rect -16680 444 -16546 446
rect -16998 430 -16546 444
rect -16489 432 -16347 488
rect -10772 501 -9968 628
rect -10772 499 -10601 501
rect -16490 430 -16347 432
rect -23503 293 -23033 294
rect -23503 292 -23201 293
rect -23503 290 -23370 292
rect -23314 291 -23201 292
rect -23145 292 -23033 293
rect -23503 234 -23371 290
rect -23314 236 -23202 291
rect -23145 237 -23034 292
rect -22977 238 -22848 294
rect -23315 235 -23202 236
rect -23146 236 -23034 237
rect -22978 236 -22848 238
rect -23146 235 -22848 236
rect -23315 234 -22848 235
rect -23503 174 -22848 234
rect -21740 300 -21640 324
rect -16998 305 -16347 430
rect -13902 462 -13802 486
rect -13902 460 -13880 462
rect -13902 404 -13881 460
rect -13824 406 -13802 462
rect -13825 404 -13802 406
rect -13902 380 -13802 404
rect -10772 443 -10602 499
rect -10545 479 -9968 501
rect -10545 477 -10233 479
rect -10545 468 -10234 477
rect -10545 466 -10401 468
rect -10545 445 -10402 466
rect -10546 443 -10402 445
rect -10772 410 -10402 443
rect -10345 421 -10234 468
rect -10177 423 -9968 479
rect -10178 421 -9968 423
rect -10345 412 -9968 421
rect -10346 410 -9968 412
rect -21740 298 -21718 300
rect -21740 242 -21719 298
rect -21662 244 -21640 300
rect -21663 242 -21640 244
rect -21740 218 -21640 242
rect -19803 281 -19703 305
rect -19803 279 -19781 281
rect -19803 223 -19782 279
rect -19725 225 -19703 281
rect -19726 223 -19703 225
rect -19803 199 -19703 223
rect -16998 303 -16734 305
rect -16998 301 -16735 303
rect -16998 299 -16917 301
rect -16998 243 -16918 299
rect -16861 247 -16735 301
rect -16678 295 -16347 305
rect -10772 305 -9968 410
rect -10772 303 -10407 305
rect -16678 293 -16558 295
rect -16678 249 -16559 293
rect -16679 247 -16559 249
rect -16861 245 -16559 247
rect -16862 243 -16559 245
rect -16998 237 -16559 243
rect -16502 239 -16347 295
rect -16503 237 -16347 239
rect -16998 176 -16347 237
rect -13907 279 -13807 303
rect -13907 277 -13885 279
rect -13907 221 -13886 277
rect -13829 223 -13807 279
rect -13830 221 -13807 223
rect -13907 198 -13807 221
rect -10772 292 -10408 303
rect -10772 290 -10594 292
rect -10772 234 -10595 290
rect -10538 247 -10408 292
rect -10351 301 -9968 305
rect -10351 299 -10224 301
rect -10351 249 -10225 299
rect -10352 247 -10225 249
rect -10538 243 -10225 247
rect -10168 245 -9968 301
rect -10169 243 -9968 245
rect -10538 236 -9968 243
rect -10539 234 -9968 236
rect -10772 163 -9968 234
rect -6954 -86 -6742 -20
rect -13781 -13232 -13048 -13201
rect -13781 -13234 -13341 -13232
rect -13781 -13246 -13342 -13234
rect -13781 -13248 -13535 -13246
rect -13781 -13304 -13536 -13248
rect -13479 -13290 -13342 -13246
rect -13285 -13288 -13048 -13232
rect -13286 -13290 -13048 -13288
rect -13479 -13302 -13048 -13290
rect -13480 -13304 -13048 -13302
rect -13781 -13314 -13048 -13304
rect -13781 -13316 -13130 -13314
rect -13781 -13348 -13131 -13316
rect -13781 -13350 -13712 -13348
rect -20281 -13383 -19756 -13350
rect -20281 -13385 -19866 -13383
rect -20281 -13387 -19867 -13385
rect -20281 -13389 -20229 -13387
rect -20281 -13445 -20230 -13389
rect -20173 -13409 -19867 -13387
rect -20173 -13411 -20070 -13409
rect -20173 -13443 -20071 -13411
rect -20174 -13445 -20071 -13443
rect -20281 -13467 -20071 -13445
rect -20014 -13441 -19867 -13409
rect -19810 -13439 -19756 -13383
rect -19811 -13441 -19756 -13439
rect -20014 -13465 -19756 -13441
rect -20015 -13467 -19756 -13465
rect -20281 -13562 -19756 -13467
rect -17491 -13409 -17391 -13385
rect -17491 -13411 -17469 -13409
rect -17491 -13467 -17470 -13411
rect -17413 -13465 -17391 -13409
rect -17414 -13467 -17391 -13465
rect -17491 -13490 -17391 -13467
rect -15196 -13396 -15096 -13372
rect -15196 -13398 -15174 -13396
rect -15196 -13454 -15175 -13398
rect -15118 -13452 -15096 -13396
rect -15119 -13454 -15096 -13452
rect -15196 -13477 -15096 -13454
rect -13781 -13406 -13713 -13350
rect -13656 -13372 -13131 -13348
rect -13074 -13370 -13048 -13314
rect -13075 -13372 -13048 -13370
rect -13656 -13404 -13048 -13372
rect -13657 -13406 -13048 -13404
rect -13781 -13431 -13048 -13406
rect -13781 -13433 -13334 -13431
rect -13781 -13436 -13335 -13433
rect -13781 -13438 -13528 -13436
rect -20281 -13564 -20232 -13562
rect -20281 -13620 -20233 -13564
rect -20176 -13587 -19756 -13562
rect -20176 -13589 -19837 -13587
rect -20176 -13595 -19838 -13589
rect -20176 -13597 -20040 -13595
rect -20176 -13618 -20041 -13597
rect -20177 -13620 -20041 -13618
rect -20281 -13653 -20041 -13620
rect -19984 -13645 -19838 -13595
rect -19781 -13643 -19756 -13587
rect -13781 -13494 -13529 -13438
rect -13472 -13489 -13335 -13436
rect -13278 -13487 -13048 -13431
rect -13279 -13489 -13048 -13487
rect -13472 -13492 -13048 -13489
rect -12255 -13411 -12155 -13387
rect -12255 -13413 -12233 -13411
rect -12255 -13469 -12234 -13413
rect -12177 -13467 -12155 -13411
rect -12178 -13469 -12155 -13467
rect -12255 -13492 -12155 -13469
rect -8329 -13392 -7592 -13279
rect -8329 -13394 -8247 -13392
rect -8329 -13450 -8248 -13394
rect -8191 -13409 -7592 -13392
rect -8191 -13411 -7915 -13409
rect -8191 -13413 -7916 -13411
rect -8191 -13415 -8072 -13413
rect -8191 -13448 -8073 -13415
rect -8192 -13450 -8073 -13448
rect -8329 -13471 -8073 -13450
rect -8016 -13467 -7916 -13413
rect -7859 -13465 -7592 -13409
rect -7860 -13467 -7592 -13465
rect -8016 -13469 -7592 -13467
rect -8017 -13471 -7592 -13469
rect -13473 -13494 -13048 -13492
rect -13781 -13635 -13048 -13494
rect -8329 -13587 -7592 -13471
rect -8329 -13589 -8274 -13587
rect -19782 -13645 -19756 -13643
rect -19984 -13651 -19756 -13645
rect -19985 -13653 -19756 -13651
rect -20281 -13708 -19756 -13653
rect -8329 -13645 -8275 -13589
rect -8218 -13591 -7592 -13587
rect -8218 -13593 -7909 -13591
rect -8218 -13595 -7910 -13593
rect -8218 -13597 -8074 -13595
rect -8218 -13643 -8075 -13597
rect -8219 -13645 -8075 -13643
rect -8329 -13653 -8075 -13645
rect -8018 -13649 -7910 -13595
rect -7853 -13647 -7592 -13591
rect -7854 -13649 -7592 -13647
rect -8018 -13651 -7592 -13649
rect -8019 -13653 -7592 -13651
rect -8329 -13707 -7592 -13653
<< via4 >>
rect -16898 503 -16842 505
rect -23021 487 -22965 489
rect -23197 484 -23141 486
rect -23369 466 -23313 468
rect -23369 412 -23314 466
rect -23314 412 -23313 466
rect -23197 430 -23142 484
rect -23142 430 -23141 484
rect -23021 433 -22966 487
rect -22966 433 -22965 487
rect -21715 469 -21659 471
rect -21715 415 -21660 469
rect -21660 415 -21659 469
rect -19770 474 -19714 476
rect -19770 420 -19715 474
rect -19715 420 -19714 474
rect -16898 449 -16843 503
rect -16843 449 -16842 503
rect -16735 500 -16679 502
rect -16735 446 -16680 500
rect -16680 446 -16679 500
rect -16545 486 -16489 488
rect -16545 432 -16490 486
rect -16490 432 -16489 486
rect -10601 499 -10545 501
rect -23370 290 -23314 292
rect -23201 291 -23145 293
rect -23033 292 -22977 294
rect -23370 236 -23315 290
rect -23315 236 -23314 290
rect -23201 237 -23146 291
rect -23146 237 -23145 291
rect -23033 238 -22978 292
rect -22978 238 -22977 292
rect -13880 460 -13824 462
rect -13880 406 -13825 460
rect -13825 406 -13824 460
rect -10601 445 -10546 499
rect -10546 445 -10545 499
rect -10233 477 -10177 479
rect -10401 466 -10345 468
rect -10401 412 -10346 466
rect -10346 412 -10345 466
rect -10233 423 -10178 477
rect -10178 423 -10177 477
rect -21718 298 -21662 300
rect -21718 244 -21663 298
rect -21663 244 -21662 298
rect -19781 279 -19725 281
rect -19781 225 -19726 279
rect -19726 225 -19725 279
rect -16734 303 -16678 305
rect -16917 299 -16861 301
rect -16917 245 -16862 299
rect -16862 245 -16861 299
rect -16734 249 -16679 303
rect -16679 249 -16678 303
rect -10407 303 -10351 305
rect -16558 293 -16502 295
rect -16558 239 -16503 293
rect -16503 239 -16502 293
rect -13885 277 -13829 279
rect -13885 223 -13830 277
rect -13830 223 -13829 277
rect -10594 290 -10538 292
rect -10594 236 -10539 290
rect -10539 236 -10538 290
rect -10407 249 -10352 303
rect -10352 249 -10351 303
rect -10224 299 -10168 301
rect -10224 245 -10169 299
rect -10169 245 -10168 299
rect -13341 -13234 -13285 -13232
rect -13535 -13248 -13479 -13246
rect -13535 -13302 -13480 -13248
rect -13480 -13302 -13479 -13248
rect -13341 -13288 -13286 -13234
rect -13286 -13288 -13285 -13234
rect -13130 -13316 -13074 -13314
rect -13712 -13350 -13656 -13348
rect -19866 -13385 -19810 -13383
rect -20229 -13389 -20173 -13387
rect -20229 -13443 -20174 -13389
rect -20174 -13443 -20173 -13389
rect -20070 -13411 -20014 -13409
rect -20070 -13465 -20015 -13411
rect -20015 -13465 -20014 -13411
rect -19866 -13439 -19811 -13385
rect -19811 -13439 -19810 -13385
rect -17469 -13411 -17413 -13409
rect -17469 -13465 -17414 -13411
rect -17414 -13465 -17413 -13411
rect -15174 -13398 -15118 -13396
rect -15174 -13452 -15119 -13398
rect -15119 -13452 -15118 -13398
rect -13712 -13404 -13657 -13350
rect -13657 -13404 -13656 -13350
rect -13130 -13370 -13075 -13316
rect -13075 -13370 -13074 -13316
rect -13334 -13433 -13278 -13431
rect -13528 -13438 -13472 -13436
rect -20232 -13564 -20176 -13562
rect -20232 -13618 -20177 -13564
rect -20177 -13618 -20176 -13564
rect -19837 -13589 -19781 -13587
rect -20040 -13597 -19984 -13595
rect -20040 -13651 -19985 -13597
rect -19985 -13651 -19984 -13597
rect -19837 -13643 -19782 -13589
rect -19782 -13643 -19781 -13589
rect -13528 -13492 -13473 -13438
rect -13473 -13492 -13472 -13438
rect -13334 -13487 -13279 -13433
rect -13279 -13487 -13278 -13433
rect -12233 -13413 -12177 -13411
rect -12233 -13467 -12178 -13413
rect -12178 -13467 -12177 -13413
rect -8247 -13394 -8191 -13392
rect -8247 -13448 -8192 -13394
rect -8192 -13448 -8191 -13394
rect -7915 -13411 -7859 -13409
rect -8072 -13415 -8016 -13413
rect -8072 -13469 -8017 -13415
rect -8017 -13469 -8016 -13415
rect -7915 -13465 -7860 -13411
rect -7860 -13465 -7859 -13411
rect -8274 -13589 -8218 -13587
rect -8274 -13643 -8219 -13589
rect -8219 -13643 -8218 -13589
rect -7909 -13593 -7853 -13591
rect -8074 -13597 -8018 -13595
rect -8074 -13651 -8019 -13597
rect -8019 -13651 -8018 -13597
rect -7909 -13647 -7854 -13593
rect -7854 -13647 -7853 -13593
<< metal5 >>
rect -16760 530 -16650 531
rect -23501 505 -9968 530
rect -23501 489 -16898 505
rect -23501 486 -23021 489
rect -23501 468 -23197 486
rect -23501 412 -23369 468
rect -23313 430 -23197 468
rect -23141 433 -23021 486
rect -22965 476 -16898 489
rect -22965 471 -19770 476
rect -22965 433 -21715 471
rect -23141 430 -21715 433
rect -23313 415 -21715 430
rect -21659 420 -19770 471
rect -19714 449 -16898 476
rect -16842 502 -9968 505
rect -16842 449 -16735 502
rect -19714 446 -16735 449
rect -16679 501 -9968 502
rect -16679 488 -10601 501
rect -16679 446 -16545 488
rect -19714 432 -16545 446
rect -16489 462 -10601 488
rect -16489 432 -13880 462
rect -19714 420 -13880 432
rect -21659 415 -13880 420
rect -23313 412 -13880 415
rect -23501 406 -13880 412
rect -13824 445 -10601 462
rect -10545 479 -9968 501
rect -10545 468 -10233 479
rect -10545 445 -10401 468
rect -13824 412 -10401 445
rect -10345 423 -10233 468
rect -10177 423 -9968 479
rect -10345 412 -9968 423
rect -13824 406 -9968 412
rect -23501 305 -9968 406
rect -23501 301 -16734 305
rect -23501 300 -16917 301
rect -23501 294 -21718 300
rect -23501 293 -23033 294
rect -23501 292 -23201 293
rect -23501 236 -23370 292
rect -23314 237 -23201 292
rect -23145 238 -23033 293
rect -22977 244 -21718 294
rect -21662 281 -16917 300
rect -21662 244 -19781 281
rect -22977 238 -19781 244
rect -23145 237 -19781 238
rect -23314 236 -19781 237
rect -23501 225 -19781 236
rect -19725 245 -16917 281
rect -16861 249 -16734 301
rect -16678 295 -10407 305
rect -16678 249 -16558 295
rect -16861 245 -16558 249
rect -19725 239 -16558 245
rect -16502 292 -10407 295
rect -16502 279 -10594 292
rect -16502 239 -13885 279
rect -19725 225 -13885 239
rect -23501 223 -13885 225
rect -13829 236 -10594 279
rect -10538 249 -10407 292
rect -10351 301 -9968 305
rect -10351 249 -10224 301
rect -10538 245 -10224 249
rect -10168 245 -9968 301
rect -10538 236 -9968 245
rect -13829 223 -9968 236
rect -23501 139 -9968 223
rect -23501 -351 -23157 139
rect -16822 -232 -16610 139
rect -10312 -325 -9968 139
rect -20280 -13278 -19942 -12580
rect -13607 -13201 -13269 -12580
rect -6955 -12839 -6739 -12505
rect -13781 -13232 -13048 -13201
rect -13781 -13246 -13341 -13232
rect -13781 -13278 -13535 -13246
rect -20280 -13302 -13535 -13278
rect -13479 -13288 -13341 -13246
rect -13285 -13278 -13048 -13232
rect -6955 -13278 -6741 -12839
rect -13285 -13288 -6741 -13278
rect -13479 -13302 -6741 -13288
rect -20280 -13314 -6741 -13302
rect -20280 -13348 -13130 -13314
rect -20280 -13350 -13712 -13348
rect -20281 -13383 -13712 -13350
rect -20281 -13387 -19866 -13383
rect -20281 -13443 -20229 -13387
rect -20173 -13409 -19866 -13387
rect -20173 -13443 -20070 -13409
rect -20281 -13465 -20070 -13443
rect -20014 -13439 -19866 -13409
rect -19810 -13396 -13712 -13383
rect -19810 -13409 -15174 -13396
rect -19810 -13439 -17469 -13409
rect -20014 -13465 -17469 -13439
rect -17413 -13452 -15174 -13409
rect -15118 -13404 -13712 -13396
rect -13656 -13370 -13130 -13348
rect -13074 -13370 -6741 -13314
rect -13656 -13392 -6741 -13370
rect -13656 -13404 -8247 -13392
rect -15118 -13411 -8247 -13404
rect -15118 -13431 -12233 -13411
rect -15118 -13436 -13334 -13431
rect -15118 -13452 -13528 -13436
rect -17413 -13465 -13528 -13452
rect -20281 -13492 -13528 -13465
rect -13472 -13487 -13334 -13436
rect -13278 -13467 -12233 -13431
rect -12177 -13448 -8247 -13411
rect -8191 -13409 -6741 -13392
rect -8191 -13413 -7915 -13409
rect -8191 -13448 -8072 -13413
rect -12177 -13467 -8072 -13448
rect -13278 -13469 -8072 -13467
rect -8016 -13465 -7915 -13413
rect -7859 -13465 -6741 -13409
rect -8016 -13469 -6741 -13465
rect -13278 -13487 -6741 -13469
rect -13472 -13492 -6741 -13487
rect -20281 -13562 -6741 -13492
rect -20281 -13618 -20232 -13562
rect -20176 -13587 -6741 -13562
rect -20176 -13595 -19837 -13587
rect -20176 -13618 -20040 -13595
rect -20281 -13651 -20040 -13618
rect -19984 -13643 -19837 -13595
rect -19781 -13616 -8274 -13587
rect -19781 -13643 -19756 -13616
rect -13781 -13635 -13048 -13616
rect -19984 -13651 -19756 -13643
rect -20281 -13708 -19756 -13651
rect -8329 -13643 -8274 -13616
rect -8218 -13591 -6741 -13587
rect -8218 -13595 -7909 -13591
rect -8218 -13643 -8074 -13595
rect -8329 -13651 -8074 -13643
rect -8018 -13647 -7909 -13595
rect -7853 -13616 -6741 -13591
rect -7853 -13647 -7592 -13616
rect -8018 -13651 -7592 -13647
rect -8329 -13707 -7592 -13651
use cap_mim_2p0fF_VGWXT2  cap_mim_2p0fF_VGWXT2_1
timestamp 1713185578
transform 1 0 -16596 0 1 -6380
box -9854 -6360 9854 6360
<< labels >>
flabel metal1 s -16715 433 -16715 433 0 FreeSans 2500 0 0 0 P
port 1 nsew
flabel metal1 s -13450 -13625 -13450 -13625 0 FreeSans 2500 0 0 0 M
port 2 nsew
<< end >>
