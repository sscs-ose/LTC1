magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1184 -1316 1184 1316
<< metal2 >>
rect -184 311 184 316
rect -184 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 184 311
rect -184 245 184 283
rect -184 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 184 245
rect -184 179 184 217
rect -184 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 184 179
rect -184 113 184 151
rect -184 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 184 113
rect -184 47 184 85
rect -184 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 184 47
rect -184 -19 184 19
rect -184 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 184 -19
rect -184 -85 184 -47
rect -184 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 184 -85
rect -184 -151 184 -113
rect -184 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 184 -151
rect -184 -217 184 -179
rect -184 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 184 -217
rect -184 -283 184 -245
rect -184 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 184 -283
rect -184 -316 184 -311
<< via2 >>
rect -179 283 -151 311
rect -113 283 -85 311
rect -47 283 -19 311
rect 19 283 47 311
rect 85 283 113 311
rect 151 283 179 311
rect -179 217 -151 245
rect -113 217 -85 245
rect -47 217 -19 245
rect 19 217 47 245
rect 85 217 113 245
rect 151 217 179 245
rect -179 151 -151 179
rect -113 151 -85 179
rect -47 151 -19 179
rect 19 151 47 179
rect 85 151 113 179
rect 151 151 179 179
rect -179 85 -151 113
rect -113 85 -85 113
rect -47 85 -19 113
rect 19 85 47 113
rect 85 85 113 113
rect 151 85 179 113
rect -179 19 -151 47
rect -113 19 -85 47
rect -47 19 -19 47
rect 19 19 47 47
rect 85 19 113 47
rect 151 19 179 47
rect -179 -47 -151 -19
rect -113 -47 -85 -19
rect -47 -47 -19 -19
rect 19 -47 47 -19
rect 85 -47 113 -19
rect 151 -47 179 -19
rect -179 -113 -151 -85
rect -113 -113 -85 -85
rect -47 -113 -19 -85
rect 19 -113 47 -85
rect 85 -113 113 -85
rect 151 -113 179 -85
rect -179 -179 -151 -151
rect -113 -179 -85 -151
rect -47 -179 -19 -151
rect 19 -179 47 -151
rect 85 -179 113 -151
rect 151 -179 179 -151
rect -179 -245 -151 -217
rect -113 -245 -85 -217
rect -47 -245 -19 -217
rect 19 -245 47 -217
rect 85 -245 113 -217
rect 151 -245 179 -217
rect -179 -311 -151 -283
rect -113 -311 -85 -283
rect -47 -311 -19 -283
rect 19 -311 47 -283
rect 85 -311 113 -283
rect 151 -311 179 -283
<< metal3 >>
rect -184 311 184 316
rect -184 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 184 311
rect -184 245 184 283
rect -184 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 184 245
rect -184 179 184 217
rect -184 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 184 179
rect -184 113 184 151
rect -184 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 184 113
rect -184 47 184 85
rect -184 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 184 47
rect -184 -19 184 19
rect -184 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 184 -19
rect -184 -85 184 -47
rect -184 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 184 -85
rect -184 -151 184 -113
rect -184 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 184 -151
rect -184 -217 184 -179
rect -184 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 184 -217
rect -184 -283 184 -245
rect -184 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 184 -283
rect -184 -316 184 -311
<< end >>
