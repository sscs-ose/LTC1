magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -2375 -1319 2375 1319
<< metal4 >>
rect -1372 311 1372 316
rect -1372 283 -1367 311
rect -1339 283 -1301 311
rect -1273 283 -1235 311
rect -1207 283 -1169 311
rect -1141 283 -1103 311
rect -1075 283 -1037 311
rect -1009 283 -971 311
rect -943 283 -905 311
rect -877 283 -839 311
rect -811 283 -773 311
rect -745 283 -707 311
rect -679 283 -641 311
rect -613 283 -575 311
rect -547 283 -509 311
rect -481 283 -443 311
rect -415 283 -377 311
rect -349 283 -311 311
rect -283 283 -245 311
rect -217 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 217 311
rect 245 283 283 311
rect 311 283 349 311
rect 377 283 415 311
rect 443 283 481 311
rect 509 283 547 311
rect 575 283 613 311
rect 641 283 679 311
rect 707 283 745 311
rect 773 283 811 311
rect 839 283 877 311
rect 905 283 943 311
rect 971 283 1009 311
rect 1037 283 1075 311
rect 1103 283 1141 311
rect 1169 283 1207 311
rect 1235 283 1273 311
rect 1301 283 1339 311
rect 1367 283 1372 311
rect -1372 245 1372 283
rect -1372 217 -1367 245
rect -1339 217 -1301 245
rect -1273 217 -1235 245
rect -1207 217 -1169 245
rect -1141 217 -1103 245
rect -1075 217 -1037 245
rect -1009 217 -971 245
rect -943 217 -905 245
rect -877 217 -839 245
rect -811 217 -773 245
rect -745 217 -707 245
rect -679 217 -641 245
rect -613 217 -575 245
rect -547 217 -509 245
rect -481 217 -443 245
rect -415 217 -377 245
rect -349 217 -311 245
rect -283 217 -245 245
rect -217 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 217 245
rect 245 217 283 245
rect 311 217 349 245
rect 377 217 415 245
rect 443 217 481 245
rect 509 217 547 245
rect 575 217 613 245
rect 641 217 679 245
rect 707 217 745 245
rect 773 217 811 245
rect 839 217 877 245
rect 905 217 943 245
rect 971 217 1009 245
rect 1037 217 1075 245
rect 1103 217 1141 245
rect 1169 217 1207 245
rect 1235 217 1273 245
rect 1301 217 1339 245
rect 1367 217 1372 245
rect -1372 179 1372 217
rect -1372 151 -1367 179
rect -1339 151 -1301 179
rect -1273 151 -1235 179
rect -1207 151 -1169 179
rect -1141 151 -1103 179
rect -1075 151 -1037 179
rect -1009 151 -971 179
rect -943 151 -905 179
rect -877 151 -839 179
rect -811 151 -773 179
rect -745 151 -707 179
rect -679 151 -641 179
rect -613 151 -575 179
rect -547 151 -509 179
rect -481 151 -443 179
rect -415 151 -377 179
rect -349 151 -311 179
rect -283 151 -245 179
rect -217 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 217 179
rect 245 151 283 179
rect 311 151 349 179
rect 377 151 415 179
rect 443 151 481 179
rect 509 151 547 179
rect 575 151 613 179
rect 641 151 679 179
rect 707 151 745 179
rect 773 151 811 179
rect 839 151 877 179
rect 905 151 943 179
rect 971 151 1009 179
rect 1037 151 1075 179
rect 1103 151 1141 179
rect 1169 151 1207 179
rect 1235 151 1273 179
rect 1301 151 1339 179
rect 1367 151 1372 179
rect -1372 113 1372 151
rect -1372 85 -1367 113
rect -1339 85 -1301 113
rect -1273 85 -1235 113
rect -1207 85 -1169 113
rect -1141 85 -1103 113
rect -1075 85 -1037 113
rect -1009 85 -971 113
rect -943 85 -905 113
rect -877 85 -839 113
rect -811 85 -773 113
rect -745 85 -707 113
rect -679 85 -641 113
rect -613 85 -575 113
rect -547 85 -509 113
rect -481 85 -443 113
rect -415 85 -377 113
rect -349 85 -311 113
rect -283 85 -245 113
rect -217 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 217 113
rect 245 85 283 113
rect 311 85 349 113
rect 377 85 415 113
rect 443 85 481 113
rect 509 85 547 113
rect 575 85 613 113
rect 641 85 679 113
rect 707 85 745 113
rect 773 85 811 113
rect 839 85 877 113
rect 905 85 943 113
rect 971 85 1009 113
rect 1037 85 1075 113
rect 1103 85 1141 113
rect 1169 85 1207 113
rect 1235 85 1273 113
rect 1301 85 1339 113
rect 1367 85 1372 113
rect -1372 47 1372 85
rect -1372 19 -1367 47
rect -1339 19 -1301 47
rect -1273 19 -1235 47
rect -1207 19 -1169 47
rect -1141 19 -1103 47
rect -1075 19 -1037 47
rect -1009 19 -971 47
rect -943 19 -905 47
rect -877 19 -839 47
rect -811 19 -773 47
rect -745 19 -707 47
rect -679 19 -641 47
rect -613 19 -575 47
rect -547 19 -509 47
rect -481 19 -443 47
rect -415 19 -377 47
rect -349 19 -311 47
rect -283 19 -245 47
rect -217 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 217 47
rect 245 19 283 47
rect 311 19 349 47
rect 377 19 415 47
rect 443 19 481 47
rect 509 19 547 47
rect 575 19 613 47
rect 641 19 679 47
rect 707 19 745 47
rect 773 19 811 47
rect 839 19 877 47
rect 905 19 943 47
rect 971 19 1009 47
rect 1037 19 1075 47
rect 1103 19 1141 47
rect 1169 19 1207 47
rect 1235 19 1273 47
rect 1301 19 1339 47
rect 1367 19 1372 47
rect -1372 -19 1372 19
rect -1372 -47 -1367 -19
rect -1339 -47 -1301 -19
rect -1273 -47 -1235 -19
rect -1207 -47 -1169 -19
rect -1141 -47 -1103 -19
rect -1075 -47 -1037 -19
rect -1009 -47 -971 -19
rect -943 -47 -905 -19
rect -877 -47 -839 -19
rect -811 -47 -773 -19
rect -745 -47 -707 -19
rect -679 -47 -641 -19
rect -613 -47 -575 -19
rect -547 -47 -509 -19
rect -481 -47 -443 -19
rect -415 -47 -377 -19
rect -349 -47 -311 -19
rect -283 -47 -245 -19
rect -217 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 217 -19
rect 245 -47 283 -19
rect 311 -47 349 -19
rect 377 -47 415 -19
rect 443 -47 481 -19
rect 509 -47 547 -19
rect 575 -47 613 -19
rect 641 -47 679 -19
rect 707 -47 745 -19
rect 773 -47 811 -19
rect 839 -47 877 -19
rect 905 -47 943 -19
rect 971 -47 1009 -19
rect 1037 -47 1075 -19
rect 1103 -47 1141 -19
rect 1169 -47 1207 -19
rect 1235 -47 1273 -19
rect 1301 -47 1339 -19
rect 1367 -47 1372 -19
rect -1372 -85 1372 -47
rect -1372 -113 -1367 -85
rect -1339 -113 -1301 -85
rect -1273 -113 -1235 -85
rect -1207 -113 -1169 -85
rect -1141 -113 -1103 -85
rect -1075 -113 -1037 -85
rect -1009 -113 -971 -85
rect -943 -113 -905 -85
rect -877 -113 -839 -85
rect -811 -113 -773 -85
rect -745 -113 -707 -85
rect -679 -113 -641 -85
rect -613 -113 -575 -85
rect -547 -113 -509 -85
rect -481 -113 -443 -85
rect -415 -113 -377 -85
rect -349 -113 -311 -85
rect -283 -113 -245 -85
rect -217 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 217 -85
rect 245 -113 283 -85
rect 311 -113 349 -85
rect 377 -113 415 -85
rect 443 -113 481 -85
rect 509 -113 547 -85
rect 575 -113 613 -85
rect 641 -113 679 -85
rect 707 -113 745 -85
rect 773 -113 811 -85
rect 839 -113 877 -85
rect 905 -113 943 -85
rect 971 -113 1009 -85
rect 1037 -113 1075 -85
rect 1103 -113 1141 -85
rect 1169 -113 1207 -85
rect 1235 -113 1273 -85
rect 1301 -113 1339 -85
rect 1367 -113 1372 -85
rect -1372 -151 1372 -113
rect -1372 -179 -1367 -151
rect -1339 -179 -1301 -151
rect -1273 -179 -1235 -151
rect -1207 -179 -1169 -151
rect -1141 -179 -1103 -151
rect -1075 -179 -1037 -151
rect -1009 -179 -971 -151
rect -943 -179 -905 -151
rect -877 -179 -839 -151
rect -811 -179 -773 -151
rect -745 -179 -707 -151
rect -679 -179 -641 -151
rect -613 -179 -575 -151
rect -547 -179 -509 -151
rect -481 -179 -443 -151
rect -415 -179 -377 -151
rect -349 -179 -311 -151
rect -283 -179 -245 -151
rect -217 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 217 -151
rect 245 -179 283 -151
rect 311 -179 349 -151
rect 377 -179 415 -151
rect 443 -179 481 -151
rect 509 -179 547 -151
rect 575 -179 613 -151
rect 641 -179 679 -151
rect 707 -179 745 -151
rect 773 -179 811 -151
rect 839 -179 877 -151
rect 905 -179 943 -151
rect 971 -179 1009 -151
rect 1037 -179 1075 -151
rect 1103 -179 1141 -151
rect 1169 -179 1207 -151
rect 1235 -179 1273 -151
rect 1301 -179 1339 -151
rect 1367 -179 1372 -151
rect -1372 -217 1372 -179
rect -1372 -245 -1367 -217
rect -1339 -245 -1301 -217
rect -1273 -245 -1235 -217
rect -1207 -245 -1169 -217
rect -1141 -245 -1103 -217
rect -1075 -245 -1037 -217
rect -1009 -245 -971 -217
rect -943 -245 -905 -217
rect -877 -245 -839 -217
rect -811 -245 -773 -217
rect -745 -245 -707 -217
rect -679 -245 -641 -217
rect -613 -245 -575 -217
rect -547 -245 -509 -217
rect -481 -245 -443 -217
rect -415 -245 -377 -217
rect -349 -245 -311 -217
rect -283 -245 -245 -217
rect -217 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 217 -217
rect 245 -245 283 -217
rect 311 -245 349 -217
rect 377 -245 415 -217
rect 443 -245 481 -217
rect 509 -245 547 -217
rect 575 -245 613 -217
rect 641 -245 679 -217
rect 707 -245 745 -217
rect 773 -245 811 -217
rect 839 -245 877 -217
rect 905 -245 943 -217
rect 971 -245 1009 -217
rect 1037 -245 1075 -217
rect 1103 -245 1141 -217
rect 1169 -245 1207 -217
rect 1235 -245 1273 -217
rect 1301 -245 1339 -217
rect 1367 -245 1372 -217
rect -1372 -283 1372 -245
rect -1372 -311 -1367 -283
rect -1339 -311 -1301 -283
rect -1273 -311 -1235 -283
rect -1207 -311 -1169 -283
rect -1141 -311 -1103 -283
rect -1075 -311 -1037 -283
rect -1009 -311 -971 -283
rect -943 -311 -905 -283
rect -877 -311 -839 -283
rect -811 -311 -773 -283
rect -745 -311 -707 -283
rect -679 -311 -641 -283
rect -613 -311 -575 -283
rect -547 -311 -509 -283
rect -481 -311 -443 -283
rect -415 -311 -377 -283
rect -349 -311 -311 -283
rect -283 -311 -245 -283
rect -217 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 217 -283
rect 245 -311 283 -283
rect 311 -311 349 -283
rect 377 -311 415 -283
rect 443 -311 481 -283
rect 509 -311 547 -283
rect 575 -311 613 -283
rect 641 -311 679 -283
rect 707 -311 745 -283
rect 773 -311 811 -283
rect 839 -311 877 -283
rect 905 -311 943 -283
rect 971 -311 1009 -283
rect 1037 -311 1075 -283
rect 1103 -311 1141 -283
rect 1169 -311 1207 -283
rect 1235 -311 1273 -283
rect 1301 -311 1339 -283
rect 1367 -311 1372 -283
rect -1372 -316 1372 -311
<< via4 >>
rect -1367 283 -1339 311
rect -1301 283 -1273 311
rect -1235 283 -1207 311
rect -1169 283 -1141 311
rect -1103 283 -1075 311
rect -1037 283 -1009 311
rect -971 283 -943 311
rect -905 283 -877 311
rect -839 283 -811 311
rect -773 283 -745 311
rect -707 283 -679 311
rect -641 283 -613 311
rect -575 283 -547 311
rect -509 283 -481 311
rect -443 283 -415 311
rect -377 283 -349 311
rect -311 283 -283 311
rect -245 283 -217 311
rect -179 283 -151 311
rect -113 283 -85 311
rect -47 283 -19 311
rect 19 283 47 311
rect 85 283 113 311
rect 151 283 179 311
rect 217 283 245 311
rect 283 283 311 311
rect 349 283 377 311
rect 415 283 443 311
rect 481 283 509 311
rect 547 283 575 311
rect 613 283 641 311
rect 679 283 707 311
rect 745 283 773 311
rect 811 283 839 311
rect 877 283 905 311
rect 943 283 971 311
rect 1009 283 1037 311
rect 1075 283 1103 311
rect 1141 283 1169 311
rect 1207 283 1235 311
rect 1273 283 1301 311
rect 1339 283 1367 311
rect -1367 217 -1339 245
rect -1301 217 -1273 245
rect -1235 217 -1207 245
rect -1169 217 -1141 245
rect -1103 217 -1075 245
rect -1037 217 -1009 245
rect -971 217 -943 245
rect -905 217 -877 245
rect -839 217 -811 245
rect -773 217 -745 245
rect -707 217 -679 245
rect -641 217 -613 245
rect -575 217 -547 245
rect -509 217 -481 245
rect -443 217 -415 245
rect -377 217 -349 245
rect -311 217 -283 245
rect -245 217 -217 245
rect -179 217 -151 245
rect -113 217 -85 245
rect -47 217 -19 245
rect 19 217 47 245
rect 85 217 113 245
rect 151 217 179 245
rect 217 217 245 245
rect 283 217 311 245
rect 349 217 377 245
rect 415 217 443 245
rect 481 217 509 245
rect 547 217 575 245
rect 613 217 641 245
rect 679 217 707 245
rect 745 217 773 245
rect 811 217 839 245
rect 877 217 905 245
rect 943 217 971 245
rect 1009 217 1037 245
rect 1075 217 1103 245
rect 1141 217 1169 245
rect 1207 217 1235 245
rect 1273 217 1301 245
rect 1339 217 1367 245
rect -1367 151 -1339 179
rect -1301 151 -1273 179
rect -1235 151 -1207 179
rect -1169 151 -1141 179
rect -1103 151 -1075 179
rect -1037 151 -1009 179
rect -971 151 -943 179
rect -905 151 -877 179
rect -839 151 -811 179
rect -773 151 -745 179
rect -707 151 -679 179
rect -641 151 -613 179
rect -575 151 -547 179
rect -509 151 -481 179
rect -443 151 -415 179
rect -377 151 -349 179
rect -311 151 -283 179
rect -245 151 -217 179
rect -179 151 -151 179
rect -113 151 -85 179
rect -47 151 -19 179
rect 19 151 47 179
rect 85 151 113 179
rect 151 151 179 179
rect 217 151 245 179
rect 283 151 311 179
rect 349 151 377 179
rect 415 151 443 179
rect 481 151 509 179
rect 547 151 575 179
rect 613 151 641 179
rect 679 151 707 179
rect 745 151 773 179
rect 811 151 839 179
rect 877 151 905 179
rect 943 151 971 179
rect 1009 151 1037 179
rect 1075 151 1103 179
rect 1141 151 1169 179
rect 1207 151 1235 179
rect 1273 151 1301 179
rect 1339 151 1367 179
rect -1367 85 -1339 113
rect -1301 85 -1273 113
rect -1235 85 -1207 113
rect -1169 85 -1141 113
rect -1103 85 -1075 113
rect -1037 85 -1009 113
rect -971 85 -943 113
rect -905 85 -877 113
rect -839 85 -811 113
rect -773 85 -745 113
rect -707 85 -679 113
rect -641 85 -613 113
rect -575 85 -547 113
rect -509 85 -481 113
rect -443 85 -415 113
rect -377 85 -349 113
rect -311 85 -283 113
rect -245 85 -217 113
rect -179 85 -151 113
rect -113 85 -85 113
rect -47 85 -19 113
rect 19 85 47 113
rect 85 85 113 113
rect 151 85 179 113
rect 217 85 245 113
rect 283 85 311 113
rect 349 85 377 113
rect 415 85 443 113
rect 481 85 509 113
rect 547 85 575 113
rect 613 85 641 113
rect 679 85 707 113
rect 745 85 773 113
rect 811 85 839 113
rect 877 85 905 113
rect 943 85 971 113
rect 1009 85 1037 113
rect 1075 85 1103 113
rect 1141 85 1169 113
rect 1207 85 1235 113
rect 1273 85 1301 113
rect 1339 85 1367 113
rect -1367 19 -1339 47
rect -1301 19 -1273 47
rect -1235 19 -1207 47
rect -1169 19 -1141 47
rect -1103 19 -1075 47
rect -1037 19 -1009 47
rect -971 19 -943 47
rect -905 19 -877 47
rect -839 19 -811 47
rect -773 19 -745 47
rect -707 19 -679 47
rect -641 19 -613 47
rect -575 19 -547 47
rect -509 19 -481 47
rect -443 19 -415 47
rect -377 19 -349 47
rect -311 19 -283 47
rect -245 19 -217 47
rect -179 19 -151 47
rect -113 19 -85 47
rect -47 19 -19 47
rect 19 19 47 47
rect 85 19 113 47
rect 151 19 179 47
rect 217 19 245 47
rect 283 19 311 47
rect 349 19 377 47
rect 415 19 443 47
rect 481 19 509 47
rect 547 19 575 47
rect 613 19 641 47
rect 679 19 707 47
rect 745 19 773 47
rect 811 19 839 47
rect 877 19 905 47
rect 943 19 971 47
rect 1009 19 1037 47
rect 1075 19 1103 47
rect 1141 19 1169 47
rect 1207 19 1235 47
rect 1273 19 1301 47
rect 1339 19 1367 47
rect -1367 -47 -1339 -19
rect -1301 -47 -1273 -19
rect -1235 -47 -1207 -19
rect -1169 -47 -1141 -19
rect -1103 -47 -1075 -19
rect -1037 -47 -1009 -19
rect -971 -47 -943 -19
rect -905 -47 -877 -19
rect -839 -47 -811 -19
rect -773 -47 -745 -19
rect -707 -47 -679 -19
rect -641 -47 -613 -19
rect -575 -47 -547 -19
rect -509 -47 -481 -19
rect -443 -47 -415 -19
rect -377 -47 -349 -19
rect -311 -47 -283 -19
rect -245 -47 -217 -19
rect -179 -47 -151 -19
rect -113 -47 -85 -19
rect -47 -47 -19 -19
rect 19 -47 47 -19
rect 85 -47 113 -19
rect 151 -47 179 -19
rect 217 -47 245 -19
rect 283 -47 311 -19
rect 349 -47 377 -19
rect 415 -47 443 -19
rect 481 -47 509 -19
rect 547 -47 575 -19
rect 613 -47 641 -19
rect 679 -47 707 -19
rect 745 -47 773 -19
rect 811 -47 839 -19
rect 877 -47 905 -19
rect 943 -47 971 -19
rect 1009 -47 1037 -19
rect 1075 -47 1103 -19
rect 1141 -47 1169 -19
rect 1207 -47 1235 -19
rect 1273 -47 1301 -19
rect 1339 -47 1367 -19
rect -1367 -113 -1339 -85
rect -1301 -113 -1273 -85
rect -1235 -113 -1207 -85
rect -1169 -113 -1141 -85
rect -1103 -113 -1075 -85
rect -1037 -113 -1009 -85
rect -971 -113 -943 -85
rect -905 -113 -877 -85
rect -839 -113 -811 -85
rect -773 -113 -745 -85
rect -707 -113 -679 -85
rect -641 -113 -613 -85
rect -575 -113 -547 -85
rect -509 -113 -481 -85
rect -443 -113 -415 -85
rect -377 -113 -349 -85
rect -311 -113 -283 -85
rect -245 -113 -217 -85
rect -179 -113 -151 -85
rect -113 -113 -85 -85
rect -47 -113 -19 -85
rect 19 -113 47 -85
rect 85 -113 113 -85
rect 151 -113 179 -85
rect 217 -113 245 -85
rect 283 -113 311 -85
rect 349 -113 377 -85
rect 415 -113 443 -85
rect 481 -113 509 -85
rect 547 -113 575 -85
rect 613 -113 641 -85
rect 679 -113 707 -85
rect 745 -113 773 -85
rect 811 -113 839 -85
rect 877 -113 905 -85
rect 943 -113 971 -85
rect 1009 -113 1037 -85
rect 1075 -113 1103 -85
rect 1141 -113 1169 -85
rect 1207 -113 1235 -85
rect 1273 -113 1301 -85
rect 1339 -113 1367 -85
rect -1367 -179 -1339 -151
rect -1301 -179 -1273 -151
rect -1235 -179 -1207 -151
rect -1169 -179 -1141 -151
rect -1103 -179 -1075 -151
rect -1037 -179 -1009 -151
rect -971 -179 -943 -151
rect -905 -179 -877 -151
rect -839 -179 -811 -151
rect -773 -179 -745 -151
rect -707 -179 -679 -151
rect -641 -179 -613 -151
rect -575 -179 -547 -151
rect -509 -179 -481 -151
rect -443 -179 -415 -151
rect -377 -179 -349 -151
rect -311 -179 -283 -151
rect -245 -179 -217 -151
rect -179 -179 -151 -151
rect -113 -179 -85 -151
rect -47 -179 -19 -151
rect 19 -179 47 -151
rect 85 -179 113 -151
rect 151 -179 179 -151
rect 217 -179 245 -151
rect 283 -179 311 -151
rect 349 -179 377 -151
rect 415 -179 443 -151
rect 481 -179 509 -151
rect 547 -179 575 -151
rect 613 -179 641 -151
rect 679 -179 707 -151
rect 745 -179 773 -151
rect 811 -179 839 -151
rect 877 -179 905 -151
rect 943 -179 971 -151
rect 1009 -179 1037 -151
rect 1075 -179 1103 -151
rect 1141 -179 1169 -151
rect 1207 -179 1235 -151
rect 1273 -179 1301 -151
rect 1339 -179 1367 -151
rect -1367 -245 -1339 -217
rect -1301 -245 -1273 -217
rect -1235 -245 -1207 -217
rect -1169 -245 -1141 -217
rect -1103 -245 -1075 -217
rect -1037 -245 -1009 -217
rect -971 -245 -943 -217
rect -905 -245 -877 -217
rect -839 -245 -811 -217
rect -773 -245 -745 -217
rect -707 -245 -679 -217
rect -641 -245 -613 -217
rect -575 -245 -547 -217
rect -509 -245 -481 -217
rect -443 -245 -415 -217
rect -377 -245 -349 -217
rect -311 -245 -283 -217
rect -245 -245 -217 -217
rect -179 -245 -151 -217
rect -113 -245 -85 -217
rect -47 -245 -19 -217
rect 19 -245 47 -217
rect 85 -245 113 -217
rect 151 -245 179 -217
rect 217 -245 245 -217
rect 283 -245 311 -217
rect 349 -245 377 -217
rect 415 -245 443 -217
rect 481 -245 509 -217
rect 547 -245 575 -217
rect 613 -245 641 -217
rect 679 -245 707 -217
rect 745 -245 773 -217
rect 811 -245 839 -217
rect 877 -245 905 -217
rect 943 -245 971 -217
rect 1009 -245 1037 -217
rect 1075 -245 1103 -217
rect 1141 -245 1169 -217
rect 1207 -245 1235 -217
rect 1273 -245 1301 -217
rect 1339 -245 1367 -217
rect -1367 -311 -1339 -283
rect -1301 -311 -1273 -283
rect -1235 -311 -1207 -283
rect -1169 -311 -1141 -283
rect -1103 -311 -1075 -283
rect -1037 -311 -1009 -283
rect -971 -311 -943 -283
rect -905 -311 -877 -283
rect -839 -311 -811 -283
rect -773 -311 -745 -283
rect -707 -311 -679 -283
rect -641 -311 -613 -283
rect -575 -311 -547 -283
rect -509 -311 -481 -283
rect -443 -311 -415 -283
rect -377 -311 -349 -283
rect -311 -311 -283 -283
rect -245 -311 -217 -283
rect -179 -311 -151 -283
rect -113 -311 -85 -283
rect -47 -311 -19 -283
rect 19 -311 47 -283
rect 85 -311 113 -283
rect 151 -311 179 -283
rect 217 -311 245 -283
rect 283 -311 311 -283
rect 349 -311 377 -283
rect 415 -311 443 -283
rect 481 -311 509 -283
rect 547 -311 575 -283
rect 613 -311 641 -283
rect 679 -311 707 -283
rect 745 -311 773 -283
rect 811 -311 839 -283
rect 877 -311 905 -283
rect 943 -311 971 -283
rect 1009 -311 1037 -283
rect 1075 -311 1103 -283
rect 1141 -311 1169 -283
rect 1207 -311 1235 -283
rect 1273 -311 1301 -283
rect 1339 -311 1367 -283
<< metal5 >>
rect -1375 311 1375 319
rect -1375 283 -1367 311
rect -1339 283 -1301 311
rect -1273 283 -1235 311
rect -1207 283 -1169 311
rect -1141 283 -1103 311
rect -1075 283 -1037 311
rect -1009 283 -971 311
rect -943 283 -905 311
rect -877 283 -839 311
rect -811 283 -773 311
rect -745 283 -707 311
rect -679 283 -641 311
rect -613 283 -575 311
rect -547 283 -509 311
rect -481 283 -443 311
rect -415 283 -377 311
rect -349 283 -311 311
rect -283 283 -245 311
rect -217 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 217 311
rect 245 283 283 311
rect 311 283 349 311
rect 377 283 415 311
rect 443 283 481 311
rect 509 283 547 311
rect 575 283 613 311
rect 641 283 679 311
rect 707 283 745 311
rect 773 283 811 311
rect 839 283 877 311
rect 905 283 943 311
rect 971 283 1009 311
rect 1037 283 1075 311
rect 1103 283 1141 311
rect 1169 283 1207 311
rect 1235 283 1273 311
rect 1301 283 1339 311
rect 1367 283 1375 311
rect -1375 245 1375 283
rect -1375 217 -1367 245
rect -1339 217 -1301 245
rect -1273 217 -1235 245
rect -1207 217 -1169 245
rect -1141 217 -1103 245
rect -1075 217 -1037 245
rect -1009 217 -971 245
rect -943 217 -905 245
rect -877 217 -839 245
rect -811 217 -773 245
rect -745 217 -707 245
rect -679 217 -641 245
rect -613 217 -575 245
rect -547 217 -509 245
rect -481 217 -443 245
rect -415 217 -377 245
rect -349 217 -311 245
rect -283 217 -245 245
rect -217 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 217 245
rect 245 217 283 245
rect 311 217 349 245
rect 377 217 415 245
rect 443 217 481 245
rect 509 217 547 245
rect 575 217 613 245
rect 641 217 679 245
rect 707 217 745 245
rect 773 217 811 245
rect 839 217 877 245
rect 905 217 943 245
rect 971 217 1009 245
rect 1037 217 1075 245
rect 1103 217 1141 245
rect 1169 217 1207 245
rect 1235 217 1273 245
rect 1301 217 1339 245
rect 1367 217 1375 245
rect -1375 179 1375 217
rect -1375 151 -1367 179
rect -1339 151 -1301 179
rect -1273 151 -1235 179
rect -1207 151 -1169 179
rect -1141 151 -1103 179
rect -1075 151 -1037 179
rect -1009 151 -971 179
rect -943 151 -905 179
rect -877 151 -839 179
rect -811 151 -773 179
rect -745 151 -707 179
rect -679 151 -641 179
rect -613 151 -575 179
rect -547 151 -509 179
rect -481 151 -443 179
rect -415 151 -377 179
rect -349 151 -311 179
rect -283 151 -245 179
rect -217 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 217 179
rect 245 151 283 179
rect 311 151 349 179
rect 377 151 415 179
rect 443 151 481 179
rect 509 151 547 179
rect 575 151 613 179
rect 641 151 679 179
rect 707 151 745 179
rect 773 151 811 179
rect 839 151 877 179
rect 905 151 943 179
rect 971 151 1009 179
rect 1037 151 1075 179
rect 1103 151 1141 179
rect 1169 151 1207 179
rect 1235 151 1273 179
rect 1301 151 1339 179
rect 1367 151 1375 179
rect -1375 113 1375 151
rect -1375 85 -1367 113
rect -1339 85 -1301 113
rect -1273 85 -1235 113
rect -1207 85 -1169 113
rect -1141 85 -1103 113
rect -1075 85 -1037 113
rect -1009 85 -971 113
rect -943 85 -905 113
rect -877 85 -839 113
rect -811 85 -773 113
rect -745 85 -707 113
rect -679 85 -641 113
rect -613 85 -575 113
rect -547 85 -509 113
rect -481 85 -443 113
rect -415 85 -377 113
rect -349 85 -311 113
rect -283 85 -245 113
rect -217 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 217 113
rect 245 85 283 113
rect 311 85 349 113
rect 377 85 415 113
rect 443 85 481 113
rect 509 85 547 113
rect 575 85 613 113
rect 641 85 679 113
rect 707 85 745 113
rect 773 85 811 113
rect 839 85 877 113
rect 905 85 943 113
rect 971 85 1009 113
rect 1037 85 1075 113
rect 1103 85 1141 113
rect 1169 85 1207 113
rect 1235 85 1273 113
rect 1301 85 1339 113
rect 1367 85 1375 113
rect -1375 47 1375 85
rect -1375 19 -1367 47
rect -1339 19 -1301 47
rect -1273 19 -1235 47
rect -1207 19 -1169 47
rect -1141 19 -1103 47
rect -1075 19 -1037 47
rect -1009 19 -971 47
rect -943 19 -905 47
rect -877 19 -839 47
rect -811 19 -773 47
rect -745 19 -707 47
rect -679 19 -641 47
rect -613 19 -575 47
rect -547 19 -509 47
rect -481 19 -443 47
rect -415 19 -377 47
rect -349 19 -311 47
rect -283 19 -245 47
rect -217 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 217 47
rect 245 19 283 47
rect 311 19 349 47
rect 377 19 415 47
rect 443 19 481 47
rect 509 19 547 47
rect 575 19 613 47
rect 641 19 679 47
rect 707 19 745 47
rect 773 19 811 47
rect 839 19 877 47
rect 905 19 943 47
rect 971 19 1009 47
rect 1037 19 1075 47
rect 1103 19 1141 47
rect 1169 19 1207 47
rect 1235 19 1273 47
rect 1301 19 1339 47
rect 1367 19 1375 47
rect -1375 -19 1375 19
rect -1375 -47 -1367 -19
rect -1339 -47 -1301 -19
rect -1273 -47 -1235 -19
rect -1207 -47 -1169 -19
rect -1141 -47 -1103 -19
rect -1075 -47 -1037 -19
rect -1009 -47 -971 -19
rect -943 -47 -905 -19
rect -877 -47 -839 -19
rect -811 -47 -773 -19
rect -745 -47 -707 -19
rect -679 -47 -641 -19
rect -613 -47 -575 -19
rect -547 -47 -509 -19
rect -481 -47 -443 -19
rect -415 -47 -377 -19
rect -349 -47 -311 -19
rect -283 -47 -245 -19
rect -217 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 217 -19
rect 245 -47 283 -19
rect 311 -47 349 -19
rect 377 -47 415 -19
rect 443 -47 481 -19
rect 509 -47 547 -19
rect 575 -47 613 -19
rect 641 -47 679 -19
rect 707 -47 745 -19
rect 773 -47 811 -19
rect 839 -47 877 -19
rect 905 -47 943 -19
rect 971 -47 1009 -19
rect 1037 -47 1075 -19
rect 1103 -47 1141 -19
rect 1169 -47 1207 -19
rect 1235 -47 1273 -19
rect 1301 -47 1339 -19
rect 1367 -47 1375 -19
rect -1375 -85 1375 -47
rect -1375 -113 -1367 -85
rect -1339 -113 -1301 -85
rect -1273 -113 -1235 -85
rect -1207 -113 -1169 -85
rect -1141 -113 -1103 -85
rect -1075 -113 -1037 -85
rect -1009 -113 -971 -85
rect -943 -113 -905 -85
rect -877 -113 -839 -85
rect -811 -113 -773 -85
rect -745 -113 -707 -85
rect -679 -113 -641 -85
rect -613 -113 -575 -85
rect -547 -113 -509 -85
rect -481 -113 -443 -85
rect -415 -113 -377 -85
rect -349 -113 -311 -85
rect -283 -113 -245 -85
rect -217 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 217 -85
rect 245 -113 283 -85
rect 311 -113 349 -85
rect 377 -113 415 -85
rect 443 -113 481 -85
rect 509 -113 547 -85
rect 575 -113 613 -85
rect 641 -113 679 -85
rect 707 -113 745 -85
rect 773 -113 811 -85
rect 839 -113 877 -85
rect 905 -113 943 -85
rect 971 -113 1009 -85
rect 1037 -113 1075 -85
rect 1103 -113 1141 -85
rect 1169 -113 1207 -85
rect 1235 -113 1273 -85
rect 1301 -113 1339 -85
rect 1367 -113 1375 -85
rect -1375 -151 1375 -113
rect -1375 -179 -1367 -151
rect -1339 -179 -1301 -151
rect -1273 -179 -1235 -151
rect -1207 -179 -1169 -151
rect -1141 -179 -1103 -151
rect -1075 -179 -1037 -151
rect -1009 -179 -971 -151
rect -943 -179 -905 -151
rect -877 -179 -839 -151
rect -811 -179 -773 -151
rect -745 -179 -707 -151
rect -679 -179 -641 -151
rect -613 -179 -575 -151
rect -547 -179 -509 -151
rect -481 -179 -443 -151
rect -415 -179 -377 -151
rect -349 -179 -311 -151
rect -283 -179 -245 -151
rect -217 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 217 -151
rect 245 -179 283 -151
rect 311 -179 349 -151
rect 377 -179 415 -151
rect 443 -179 481 -151
rect 509 -179 547 -151
rect 575 -179 613 -151
rect 641 -179 679 -151
rect 707 -179 745 -151
rect 773 -179 811 -151
rect 839 -179 877 -151
rect 905 -179 943 -151
rect 971 -179 1009 -151
rect 1037 -179 1075 -151
rect 1103 -179 1141 -151
rect 1169 -179 1207 -151
rect 1235 -179 1273 -151
rect 1301 -179 1339 -151
rect 1367 -179 1375 -151
rect -1375 -217 1375 -179
rect -1375 -245 -1367 -217
rect -1339 -245 -1301 -217
rect -1273 -245 -1235 -217
rect -1207 -245 -1169 -217
rect -1141 -245 -1103 -217
rect -1075 -245 -1037 -217
rect -1009 -245 -971 -217
rect -943 -245 -905 -217
rect -877 -245 -839 -217
rect -811 -245 -773 -217
rect -745 -245 -707 -217
rect -679 -245 -641 -217
rect -613 -245 -575 -217
rect -547 -245 -509 -217
rect -481 -245 -443 -217
rect -415 -245 -377 -217
rect -349 -245 -311 -217
rect -283 -245 -245 -217
rect -217 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 217 -217
rect 245 -245 283 -217
rect 311 -245 349 -217
rect 377 -245 415 -217
rect 443 -245 481 -217
rect 509 -245 547 -217
rect 575 -245 613 -217
rect 641 -245 679 -217
rect 707 -245 745 -217
rect 773 -245 811 -217
rect 839 -245 877 -217
rect 905 -245 943 -217
rect 971 -245 1009 -217
rect 1037 -245 1075 -217
rect 1103 -245 1141 -217
rect 1169 -245 1207 -217
rect 1235 -245 1273 -217
rect 1301 -245 1339 -217
rect 1367 -245 1375 -217
rect -1375 -283 1375 -245
rect -1375 -311 -1367 -283
rect -1339 -311 -1301 -283
rect -1273 -311 -1235 -283
rect -1207 -311 -1169 -283
rect -1141 -311 -1103 -283
rect -1075 -311 -1037 -283
rect -1009 -311 -971 -283
rect -943 -311 -905 -283
rect -877 -311 -839 -283
rect -811 -311 -773 -283
rect -745 -311 -707 -283
rect -679 -311 -641 -283
rect -613 -311 -575 -283
rect -547 -311 -509 -283
rect -481 -311 -443 -283
rect -415 -311 -377 -283
rect -349 -311 -311 -283
rect -283 -311 -245 -283
rect -217 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 217 -283
rect 245 -311 283 -283
rect 311 -311 349 -283
rect 377 -311 415 -283
rect 443 -311 481 -283
rect 509 -311 547 -283
rect 575 -311 613 -283
rect 641 -311 679 -283
rect 707 -311 745 -283
rect 773 -311 811 -283
rect 839 -311 877 -283
rect 905 -311 943 -283
rect 971 -311 1009 -283
rect 1037 -311 1075 -283
rect 1103 -311 1141 -283
rect 1169 -311 1207 -283
rect 1235 -311 1273 -283
rect 1301 -311 1339 -283
rect 1367 -311 1375 -283
rect -1375 -319 1375 -311
<< end >>
