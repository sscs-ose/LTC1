magic
tech gf180mcuC
magscale 1 10
timestamp 1691673501
<< nwell >>
rect -62 731 342 856
<< psubdiff >>
rect 10 -45 270 -32
rect 10 -91 23 -45
rect 69 -91 117 -45
rect 163 -91 211 -45
rect 257 -91 270 -45
rect 10 -104 270 -91
<< nsubdiff >>
rect -37 810 317 823
rect -37 764 -24 810
rect 22 764 70 810
rect 116 764 164 810
rect 210 764 258 810
rect 304 764 317 810
rect -37 751 317 764
<< psubdiffcont >>
rect 23 -91 69 -45
rect 117 -91 163 -45
rect 211 -91 257 -45
<< nsubdiffcont >>
rect -24 764 22 810
rect 70 764 116 810
rect 164 764 210 810
rect 258 764 304 810
<< polysilicon >>
rect -8 274 64 282
rect 112 274 168 446
rect -8 269 168 274
rect -8 223 5 269
rect 51 223 168 269
rect -8 218 168 223
rect -8 210 64 218
rect 112 173 168 218
<< polycontact >>
rect 5 223 51 269
<< metal1 >>
rect -62 810 342 843
rect -62 764 -24 810
rect 22 764 70 810
rect 116 764 164 810
rect 210 764 258 810
rect 304 764 342 810
rect -62 731 342 764
rect 37 609 83 731
rect 197 396 243 470
rect 197 350 340 396
rect -6 269 62 280
rect -60 223 5 269
rect 51 223 62 269
rect -6 212 62 223
rect 197 141 243 350
rect 37 -12 83 98
rect -10 -45 290 -12
rect -10 -91 23 -45
rect 69 -91 117 -45
rect 163 -91 211 -45
rect 257 -91 290 -45
rect -10 -124 290 -91
use nmos_3p3_GGGST2#3  nmos_3p3_GGGST2_0
timestamp 1691670445
transform 1 0 140 0 1 118
box -140 -118 140 118
use pmos_3p3_MNVUAR#3  pmos_3p3_MNVUAR_0
timestamp 1691670445
transform 1 0 140 0 1 540
box -202 -230 202 230
<< labels >>
flabel psubdiffcont 140 -68 140 -68 0 FreeSans 320 0 0 0 VSS
port 7 nsew
flabel metal1 140 790 140 790 0 FreeSans 320 0 0 0 VDD
port 9 nsew
flabel metal1 -40 246 -40 246 0 FreeSans 320 0 0 0 IN
port 4 nsew
flabel metal1 279 373 279 373 0 FreeSans 320 0 0 0 OUT
port 6 nsew
<< end >>
