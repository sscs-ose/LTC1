magic
tech gf180mcuC
magscale 1 10
timestamp 1695119997
<< polysilicon >>
rect 892 1016 2388 1072
rect 892 915 948 1016
rect 1052 915 1108 1016
rect 1212 915 1268 1016
rect 1372 915 1428 1016
rect 1532 915 1588 1016
rect 1692 915 1748 1016
rect 1852 915 1908 1016
rect 2012 915 2068 1016
rect 2172 915 2228 1016
rect 2332 915 2388 1016
rect 892 616 943 671
rect 659 598 943 616
rect 659 541 673 598
rect 726 549 943 598
rect 726 541 742 549
rect 659 516 742 541
rect 891 181 948 207
rect 831 166 948 181
rect 831 119 851 166
rect 897 158 948 166
rect 1052 158 1108 206
rect 1212 158 1268 206
rect 1372 158 1428 206
rect 1532 158 1588 206
rect 1692 158 1748 206
rect 1852 158 1908 206
rect 2012 158 2068 206
rect 2172 158 2228 206
rect 2332 158 2388 206
rect 897 119 2388 158
rect 831 103 2388 119
rect 832 102 2388 103
<< polycontact >>
rect 673 541 726 598
rect 851 119 897 166
<< metal1 >>
rect 314 926 719 1097
rect 804 920 2483 983
rect 620 616 695 617
rect 620 598 734 616
rect 285 565 360 575
rect 285 562 418 565
rect 285 504 299 562
rect 353 515 418 562
rect 620 541 673 598
rect 726 541 734 598
rect 620 517 734 541
rect 659 516 734 517
rect 353 504 360 515
rect 285 490 360 504
rect 804 250 872 920
rect 314 127 719 241
rect 831 169 913 181
rect 831 114 847 169
rect 900 114 913 169
rect 831 103 913 114
rect 966 151 1034 871
rect 1124 250 1192 920
rect 1285 151 1353 871
rect 1445 250 1513 920
rect 1605 151 1673 871
rect 1764 250 1832 920
rect 1924 151 1992 871
rect 2085 251 2153 920
rect 2246 545 2314 871
rect 2246 492 2251 545
rect 2307 492 2314 545
rect 2246 151 2314 492
rect 2405 680 2473 920
rect 2405 612 2689 680
rect 2405 251 2473 612
rect 2603 540 2690 551
rect 2603 488 2618 540
rect 2674 488 2690 540
rect 2603 474 2690 488
rect 966 101 2314 151
rect 967 83 2314 101
<< via1 >>
rect 299 504 353 562
rect 847 166 900 169
rect 847 119 851 166
rect 851 119 897 166
rect 897 119 900 166
rect 847 114 900 119
rect 2251 492 2307 545
rect 2618 488 2674 540
<< metal2 >>
rect 285 562 360 575
rect 285 504 299 562
rect 353 504 360 562
rect 285 490 360 504
rect 2239 547 2314 554
rect 2603 547 2690 551
rect 2239 545 2690 547
rect 2239 492 2251 545
rect 2307 540 2690 545
rect 2307 492 2618 540
rect 295 359 352 490
rect 2239 488 2618 492
rect 2674 488 2690 540
rect 2239 482 2690 488
rect 2239 478 2314 482
rect 2603 474 2690 482
rect 295 300 948 359
rect 885 181 944 300
rect 831 169 944 181
rect 831 114 847 169
rect 900 114 944 169
rect 831 112 944 114
rect 831 103 913 112
use inv_my_mag  inv_my_mag_0
timestamp 1695119997
transform 1 0 375 0 1 69
box -61 58 345 1028
use nmos_3p3_W9BEG7  nmos_3p3_W9BEG7_0
timestamp 1693575223
transform 1 0 1640 0 1 350
box -860 -168 860 168
use pmos_3p3_Q354KU  pmos_3p3_Q354KU_0
timestamp 1693575223
transform 1 0 1640 0 1 771
box -922 -230 922 230
<< labels >>
flabel via1 323 537 323 537 0 FreeSans 480 0 0 0 CLK
port 2 nsew
flabel metal1 505 1060 505 1060 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal1 498 179 498 179 0 FreeSans 480 0 0 0 VSS
port 4 nsew
flabel metal1 2663 654 2663 654 0 FreeSans 480 0 0 0 VIN
port 5 nsew
flabel via1 2640 510 2640 510 0 FreeSans 480 0 0 0 VOUT
port 6 nsew
<< end >>
