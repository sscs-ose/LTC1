* NGSPICE file created from CLK_div_10_mag_flat.ext - technology: gf180mcuC

.subckt CLK_div_10_mag_flat CLK VSS VDD Q0 Vdiv10 RST Q3 Q1 Q2
X0 JK_FF_mag_2.nand3_mag_2.OUT Q1.t3 VDD.t191 VDD.t190 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1 a_794_1309# CLK.t0 a_634_1309# VSS.t106 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2 Q1 JK_FF_mag_2.Qb a_5503_1353# VSS.t108 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand3_mag_1.IN1 VDD.t25 VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 a_4375_1353# JK_FF_mag_2.nand3_mag_0.OUT VSS.t49 VSS.t48 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X5 VDD Q0.t3 JK_FF_mag_0.nand3_mag_2.OUT VDD.t75 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X6 JK_FF_mag_2.nand2_mag_3.IN1 Q0.t4 VDD.t17 VDD.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.J.t3 VDD.t146 VDD.t145 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 VSS and2_mag_0.OUT Vdiv10.t0 VSS.t39 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X9 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 VDD.t128 VDD.t127 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X10 a_9510_2450# Q0.t5 VSS.t14 VSS.t13 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X11 a_2076_256# JK_FF_mag_1.nand3_mag_1.OUT VSS.t31 VSS.t30 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X12 nor_3_mag_0.IN3 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t82 VSS.t81 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X13 a_788_212# CLK.t1 a_628_212# VSS.t105 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X14 VDD JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_1.IN2 VDD.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X15 Q1 JK_FF_mag_2.nand2_mag_1.IN2 VDD.t60 VDD.t59 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X16 a_9845_1309# Q0.t6 a_9685_1309# VSS.t16 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X17 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand3_mag_1.OUT VDD.t65 VDD.t64 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 JK_FF_mag_2.nand3_mag_2.OUT Q1.t4 a_3805_212# VSS.t124 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X19 VDD RST.t0 JK_FF_mag_0.nand3_mag_1.OUT VDD.t82 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X20 JK_FF_mag_0.J and2_mag_2.GF_INV_MAG_0.IN VSS.t84 VSS.t83 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X21 VDD JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t52 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X22 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 VDD.t41 VDD.t40 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 a_9839_212# Q0.t7 a_9679_212# VSS.t17 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X24 a_9685_1309# JK_FF_mag_0.J VSS.t112 VSS.t111 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X25 and2_mag_0.GF_INV_MAG_0.IN Q2.t3 a_7574_2450# VSS.t15 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X26 VDD JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t35 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X27 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand3_mag_1.IN1 VDD.t224 VDD.t223 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X28 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 a_7546_212# VSS.t91 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X29 JK_FF_mag_1.nand3_mag_2.OUT Q0.t8 VDD.t173 VDD.t172 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X30 JK_FF_mag_1.Qb Q0.t9 a_2640_256# VSS.t115 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X31 VDD Q1.t5 JK_FF_mag_2.Qb VDD.t187 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X32 JK_FF_mag_2.nand3_mag_2.OUT VDD.t107 VDD.t109 VDD.t108 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X33 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.Qb a_6828_1309# VSS.t126 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X34 a_7574_2450# Q1.t6 VSS.t123 VSS.t122 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X35 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_11127_256# VSS.t132 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X36 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT VDD.t27 VDD.t26 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 VDD RST.t1 JK_FF_mag_1.nand3_mag_1.OUT VDD.t197 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X38 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.Qb VDD.t7 VDD.t6 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X39 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t69 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X40 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand2_mag_3.IN1 a_7956_1353# VSS.t88 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X41 and2_mag_0.OUT and2_mag_0.GF_INV_MAG_0.IN VDD.t226 VDD.t225 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X42 and2_mag_2.GF_INV_MAG_0.IN Q2.t4 VDD.t19 VDD.t18 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X43 a_10563_212# RST.t2 a_10403_212# VSS.t127 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X44 a_8520_1353# JK_FF_mag_3.nand2_mag_1.IN2 VSS.t98 VSS.t97 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X45 a_5657_256# JK_FF_mag_2.nand2_mag_4.IN2 VSS.t64 VSS.t63 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X46 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_2076_256# VSS.t58 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X47 VDD CLK.t2 JK_FF_mag_1.nand3_mag_0.OUT VDD.t169 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X48 JK_FF_mag_3.nand3_mag_2.OUT Q2.t5 VDD.t21 VDD.t20 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X49 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_2.OUT VDD.t43 VDD.t42 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X50 VDD Q2.t6 and2_mag_1.GF_INV_MAG_0.IN VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X51 JK_FF_mag_1.nand3_mag_2.OUT Q0.t10 a_788_212# VSS.t94 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X52 a_3645_212# VDD.t227 VSS.t76 VSS.t75 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X53 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.Qb a_3811_1309# VSS.t107 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X54 a_4939_1353# JK_FF_mag_2.nand3_mag_1.IN1 VSS.t20 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X55 JK_FF_mag_3.Qb JK_FF_mag_3.nand2_mag_4.IN2 VDD.t13 VDD.t12 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X56 VDD JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_4.IN2 VDD.t132 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X57 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN and2_mag_1.OUT VSS.t136 VSS.t135 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X58 a_1512_212# RST.t3 a_1352_212# VSS.t23 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X59 VDD Q0.t11 JK_FF_mag_0.nand3_mag_0.OUT VDD.t129 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X60 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t39 VDD.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X61 Vdiv10 Q3.t3 a_11738_2752# VDD.t124 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X62 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_3.IN1 a_4939_1353# VSS.t96 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X63 a_634_1309# VDD.t228 VSS.t78 VSS.t77 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X64 a_5503_1353# JK_FF_mag_2.nand2_mag_1.IN2 VSS.t53 VSS.t52 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X65 a_5093_256# JK_FF_mag_2.nand3_mag_1.OUT VSS.t56 VSS.t55 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X66 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand3_mag_1.OUT VDD.t49 VDD.t48 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X67 JK_FF_mag_0.nand2_mag_3.IN1 Q0.t12 VDD.t15 VDD.t14 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X68 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.J VDD.t166 VDD.t165 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X69 JK_FF_mag_3.nand3_mag_2.OUT Q2.t7 a_6822_212# VSS.t62 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X70 a_4369_212# JK_FF_mag_2.nand3_mag_2.OUT VSS.t36 VSS.t35 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X71 JK_FF_mag_2.nand2_mag_3.IN1 Q0.t13 VSS.t12 VSS.t11 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X72 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT a_10409_1353# VSS.t47 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X73 a_10973_1353# JK_FF_mag_0.nand3_mag_1.IN1 VSS.t34 VSS.t33 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X74 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.Qb VDD.t196 VDD.t195 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X75 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT a_1358_1353# VSS.t29 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X76 a_1922_1353# JK_FF_mag_1.nand3_mag_1.IN1 VSS.t139 VSS.t138 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X77 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 a_10563_212# VSS.t32 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X78 JK_FF_mag_2.Qb Q1.t7 a_5657_256# VSS.t121 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X79 and2_mag_1.OUT and2_mag_1.GF_INV_MAG_0.IN VDD.t215 VDD.t214 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X80 VDD JK_FF_mag_2.J.t4 Q3.t2 VDD.t147 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 a_1358_1353# JK_FF_mag_1.nand3_mag_0.OUT VSS.t22 VSS.t21 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X82 VDD RST.t4 JK_FF_mag_2.nand3_mag_1.OUT VDD.t28 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X83 VDD JK_FF_mag_1.Qb Q0.t1 VDD.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X84 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT VDD.t151 VDD.t150 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X85 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_1922_1353# VSS.t57 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X86 JK_FF_mag_3.nand2_mag_3.IN1 Q1.t8 VDD.t186 VDD.t185 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X87 VDD Q2.t8 JK_FF_mag_3.Qb VDD.t152 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X88 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t211 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X89 and2_mag_2.GF_INV_MAG_0.IN Q1.t9 a_8542_2450# VSS.t120 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X90 a_6828_1309# Q1.t10 a_6668_1309# VSS.t119 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X91 Q0 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t11 VDD.t10 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X92 JK_FF_mag_2.J JK_FF_mag_0.nand2_mag_4.IN2 VDD.t111 VDD.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X93 JK_FF_mag_0.nand3_mag_2.OUT Q3.t4 VDD.t79 VDD.t78 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X94 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.Qb VDD.t162 VDD.t161 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X95 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_2.OUT VDD.t91 VDD.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X96 a_6668_1309# VDD.t229 VSS.t74 VSS.t73 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X97 a_8674_256# JK_FF_mag_3.nand2_mag_4.IN2 VSS.t10 VSS.t9 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X98 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_3.IN1 a_5093_256# VSS.t95 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X99 a_4529_212# RST.t5 a_4369_212# VSS.t129 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X100 JK_FF_mag_1.nand2_mag_3.IN1 CLK.t3 VDD.t204 VDD.t203 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X101 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t51 VDD.t50 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X102 JK_FF_mag_1.Qb JK_FF_mag_1.nand2_mag_4.IN2 VDD.t164 VDD.t163 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X103 JK_FF_mag_1.nand3_mag_0.OUT VDD.t104 VDD.t106 VDD.t105 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X104 JK_FF_mag_0.J and2_mag_2.GF_INV_MAG_0.IN VDD.t115 VDD.t114 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X105 and2_mag_1.GF_INV_MAG_0.IN Q0.t14 VDD.t81 VDD.t80 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X106 a_8110_256# JK_FF_mag_3.nand3_mag_1.OUT VSS.t44 VSS.t43 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X107 a_3811_1309# Q0.t15 a_3651_1309# VSS.t60 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X108 JK_FF_mag_0.nand3_mag_2.OUT Q3.t5 a_9839_212# VSS.t59 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X109 a_7386_212# JK_FF_mag_3.nand3_mag_2.OUT VSS.t66 VSS.t65 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X110 JK_FF_mag_1.nand3_mag_2.OUT VDD.t101 VDD.t103 VDD.t102 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X111 VDD Q0.t16 JK_FF_mag_2.nand3_mag_2.OUT VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X112 a_11738_2752# and2_mag_0.OUT a_11578_2752# VDD.t44 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X113 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t222 VDD.t221 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X114 VDD Q2.t9 and2_mag_0.GF_INV_MAG_0.IN VDD.t155 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X115 VDD Q3.t6 JK_FF_mag_2.J.t2 VDD.t142 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X116 JK_FF_mag_0.nand2_mag_3.IN1 Q0.t17 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X117 VDD RST.t6 JK_FF_mag_3.nand3_mag_1.OUT VDD.t200 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X118 Q3 JK_FF_mag_2.J.t5 a_11537_1353# VSS.t37 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X119 a_11578_2752# nor_3_mag_0.IN3 VDD.t117 VDD.t116 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X120 a_10409_1353# JK_FF_mag_0.nand3_mag_0.OUT VSS.t102 VSS.t101 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X121 and2_mag_0.GF_INV_MAG_0.IN Q1.t11 VDD.t184 VDD.t183 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X122 Q0 JK_FF_mag_1.Qb a_2486_1353# VSS.t3 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X123 JK_FF_mag_3.nand3_mag_2.OUT VDD.t98 VDD.t100 VDD.t99 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X124 VDD Q1.t12 JK_FF_mag_3.nand3_mag_0.OUT VDD.t180 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X125 JK_FF_mag_3.Qb Q2.t10 a_8674_256# VSS.t24 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X126 a_628_212# VDD.t230 VSS.t72 VSS.t71 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X127 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_10973_1353# VSS.t131 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X128 VDD JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 VDD.t45 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X129 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand3_mag_1.IN1 VDD.t126 VDD.t125 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X130 a_2486_1353# JK_FF_mag_1.nand2_mag_1.IN2 VSS.t8 VSS.t7 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X131 a_11691_256# JK_FF_mag_0.nand2_mag_4.IN2 VSS.t80 VSS.t79 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X132 a_3805_212# Q0.t18 a_3645_212# VSS.t130 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X133 JK_FF_mag_3.nand3_mag_0.OUT VDD.t95 VDD.t97 VDD.t96 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X134 VDD JK_FF_mag_3.Qb Q2.t1 VDD.t192 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X135 Q3 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t141 VDD.t140 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X136 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 a_1512_212# VSS.t137 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X137 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT VDD.t32 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X138 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_0.OUT VDD.t168 VDD.t167 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X139 Vdiv10 Q3.t7 VSS.t93 VSS.t92 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X140 a_7546_212# RST.t7 a_7386_212# VSS.t128 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X141 JK_FF_mag_3.nand2_mag_3.IN1 Q1.t13 VSS.t118 VSS.t117 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X142 a_8542_2450# Q2.t11 VSS.t26 VSS.t25 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X143 a_11127_256# JK_FF_mag_0.nand3_mag_1.OUT VSS.t46 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X144 a_6662_212# VDD.t231 VSS.t70 VSS.t69 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X145 a_2640_256# JK_FF_mag_1.nand2_mag_4.IN2 VSS.t110 VSS.t109 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X146 nor_3_mag_0.IN3 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t113 VDD.t112 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X147 VDD JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_4.IN2 VDD.t121 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X148 VDD Q0.t19 JK_FF_mag_2.nand3_mag_0.OUT VDD.t205 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X149 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_2.OUT VDD.t9 VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X150 and2_mag_1.GF_INV_MAG_0.IN Q2.t12 a_9510_2450# VSS.t61 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X151 VDD JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 VDD.t61 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X152 a_10403_212# JK_FF_mag_0.nand3_mag_2.OUT VSS.t28 VSS.t27 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X153 VDD JK_FF_mag_2.Qb Q1.t1 VDD.t158 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X154 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_2.J.t6 a_9845_1309# VSS.t38 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X155 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_0.OUT VDD.t56 VDD.t55 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X156 VDD Q1.t14 JK_FF_mag_3.nand3_mag_2.OUT VDD.t177 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X157 and2_mag_0.OUT and2_mag_0.GF_INV_MAG_0.IN VSS.t141 VSS.t140 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X158 JK_FF_mag_1.nand2_mag_3.IN1 CLK.t4 VSS.t104 VSS.t103 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X159 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 VDD.t23 VDD.t22 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X160 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT VDD.t34 VDD.t33 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X161 a_3651_1309# JK_FF_mag_2.J.t7 VSS.t51 VSS.t50 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X162 JK_FF_mag_2.J Q3.t8 a_11691_256# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X163 a_1352_212# JK_FF_mag_1.nand3_mag_2.OUT VSS.t5 VSS.t4 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X164 JK_FF_mag_0.nand3_mag_2.OUT VDD.t92 VDD.t94 VDD.t93 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X165 Vdiv10 nor_3_mag_0.IN3 VSS.t86 VSS.t85 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X166 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_1.OUT a_7392_1353# VSS.t42 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X167 a_6822_212# Q1.t15 a_6662_212# VSS.t116 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X168 a_7956_1353# JK_FF_mag_3.nand3_mag_1.IN1 VSS.t90 VSS.t89 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X169 a_11537_1353# JK_FF_mag_0.nand2_mag_1.IN2 VSS.t100 VSS.t99 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X170 VDD Q1.t16 and2_mag_2.GF_INV_MAG_0.IN VDD.t174 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 a_4529_212# VSS.t18 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X172 Q2 JK_FF_mag_3.Qb a_8520_1353# VSS.t125 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X173 a_7392_1353# JK_FF_mag_3.nand3_mag_0.OUT VSS.t114 VSS.t113 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X174 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 VDD.t208 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X175 VDD Q0.t20 JK_FF_mag_1.Qb VDD.t72 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X176 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN and2_mag_1.OUT VDD.t217 VDD.t216 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X177 a_9679_212# VDD.t232 VSS.t68 VSS.t67 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X178 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand2_mag_3.IN1 a_8110_256# VSS.t87 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X179 VDD JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_1.IN2 VDD.t118 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X180 Q2 JK_FF_mag_3.nand2_mag_1.IN2 VDD.t139 VDD.t138 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X181 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.Qb a_794_1309# VSS.t2 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X182 VDD CLK.t5 JK_FF_mag_1.nand3_mag_2.OUT VDD.t218 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X183 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_1.OUT a_4375_1353# VSS.t54 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X184 JK_FF_mag_2.Qb JK_FF_mag_2.nand2_mag_4.IN2 VDD.t89 VDD.t88 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X185 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 VDD.t66 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X186 and2_mag_1.OUT and2_mag_1.GF_INV_MAG_0.IN VSS.t134 VSS.t133 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X187 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_2.J.t8 VDD.t58 VDD.t57 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 Q1.n8 Q1.t4 36.935
R1 Q1.n40 Q1.t10 36.935
R2 Q1.n0 Q1.t15 36.935
R3 Q1.n10 Q1.t7 31.528
R4 Q1.n23 Q1.t9 31.528
R5 Q1.n28 Q1.t11 30.9379
R6 Q1.n15 Q1.t8 25.5364
R7 Q1.n28 Q1.t6 21.6422
R8 Q1.n8 Q1.t3 18.1962
R9 Q1.n40 Q1.t12 18.1962
R10 Q1.n0 Q1.t14 18.1962
R11 Q1.n10 Q1.t5 15.3826
R12 Q1.n23 Q1.t16 15.3826
R13 Q1.n15 Q1.t13 14.0749
R14 Q1.n6 Q1.n3 7.09905
R15 Q1.n11 Q1.n10 6.86134
R16 Q1.n24 Q1.n23 5.62394
R17 Q1.n12 Q1.n9 5.01116
R18 Q1.n44 Q1.n43 4.5005
R19 Q1.n39 Q1.n38 4.5005
R20 Q1.n34 Q1.n33 3.81183
R21 Q1.n6 Q1.n5 3.25085
R22 Q1.n33 Q1.n26 3.06735
R23 Q1.n5 Q1.t1 2.2755
R24 Q1.n5 Q1.n4 2.2755
R25 Q1.n13 Q1.n7 2.2505
R26 Q1.n19 Q1.n18 2.24235
R27 Q1.n32 Q1.n31 2.24151
R28 Q1.n26 Q1.n25 2.2414
R29 Q1.n9 Q1.n8 2.13398
R30 Q1.n29 Q1.n28 2.12245
R31 Q1.n1 Q1.n0 2.12175
R32 Q1.n41 Q1.n40 2.12084
R33 Q1.n46 Q1.n44 1.71062
R34 Q1.n35 Q1.n34 1.54045
R35 Q1.n13 Q1.n12 1.5289
R36 Q1.n47 Q1.n46 1.49778
R37 Q1.n16 Q1.n15 1.42706
R38 Q1.n12 Q1.n11 1.12056
R39 Q1.n20 Q1.n19 0.962512
R40 Q1.n33 Q1.n32 0.961174
R41 Q1.n14 Q1 0.644908
R42 Q1.n17 Q1 0.1605
R43 Q1.n7 Q1.n6 0.0919062
R44 Q1.n11 Q1 0.0857632
R45 Q1.n9 Q1 0.0810725
R46 Q1.n30 Q1 0.0749415
R47 Q1.n7 Q1 0.073625
R48 Q1.n38 Q1 0.0473512
R49 Q1 Q1.n48 0.0473512
R50 Q1.n22 Q1 0.0460172
R51 Q1.n48 Q1.n47 0.0361897
R52 Q1.n44 Q1.n39 0.0328437
R53 Q1 Q1.n13 0.0322045
R54 Q1.n18 Q1.n17 0.03175
R55 Q1.n25 Q1.n22 0.028431
R56 Q1.n19 Q1.n14 0.0246174
R57 Q1.n26 Q1.n21 0.0234177
R58 Q1.n32 Q1.n27 0.0215128
R59 Q1.n31 Q1.n30 0.02075
R60 Q1.n20 Q1.n2 0.0168541
R61 Q1.n35 Q1.n20 0.0145871
R62 Q1.n46 Q1.n45 0.0131772
R63 Q1.n25 Q1.n24 0.0129138
R64 Q1.n31 Q1.n29 0.0095
R65 Q1.n43 Q1.n42 0.00515517
R66 Q1.n47 Q1.n1 0.00515517
R67 Q1.n39 Q1.n36 0.00471875
R68 Q1.n36 Q1.n35 0.00287694
R69 Q1.n38 Q1.n37 0.00205172
R70 Q1.n18 Q1.n16 0.00175
R71 Q1.n42 Q1.n41 0.00140935
R72 VDD.n207 VDD.n206 11185.2
R73 VDD.n154 VDD.n153 11185.2
R74 VDD.n131 VDD.t112 1105.93
R75 VDD.t69 VDD.t10 961.905
R76 VDD.t6 VDD.t26 961.905
R77 VDD.t135 VDD.t59 961.905
R78 VDD.t161 VDD.t55 961.905
R79 VDD.t118 VDD.t138 961.905
R80 VDD.t167 VDD.t195 961.905
R81 VDD.t66 VDD.t163 765.152
R82 VDD.t221 VDD.t33 765.152
R83 VDD.t172 VDD.t8 765.152
R84 VDD.t140 VDD.t211 765.152
R85 VDD.t52 VDD.t40 765.152
R86 VDD.t150 VDD.t57 765.152
R87 VDD.t208 VDD.t110 765.152
R88 VDD.t38 VDD.t50 765.152
R89 VDD.t78 VDD.t31 765.152
R90 VDD.t121 VDD.t12 765.152
R91 VDD.t127 VDD.t48 765.152
R92 VDD.t20 VDD.t90 765.152
R93 VDD.t132 VDD.t88 765.152
R94 VDD.t22 VDD.t64 765.152
R95 VDD.t190 VDD.t42 765.152
R96 VDD.n128 VDD.t116 747.159
R97 VDD.n206 VDD.t223 676.191
R98 VDD.t24 VDD.n182 676.191
R99 VDD.n153 VDD.t125 676.191
R100 VDD.t214 VDD.t216 645.307
R101 VDD.n207 VDD.t105 485.714
R102 VDD.n154 VDD.t96 485.714
R103 VDD VDD.n84 429.187
R104 VDD VDD.n137 427.092
R105 VDD.n143 VDD 427.092
R106 VDD.t203 VDD.n207 426.44
R107 VDD.t16 VDD.n196 426.44
R108 VDD.t185 VDD.n154 426.44
R109 VDD VDD.n132 425.019
R110 VDD.n84 VDD.t165 386.365
R111 VDD.n143 VDD.t18 386.365
R112 VDD.n137 VDD.t80 386.365
R113 VDD.t169 VDD.t6 380.952
R114 VDD.t205 VDD.t161 380.952
R115 VDD.t195 VDD.t180 380.952
R116 VDD.t155 VDD.n143 378.788
R117 VDD.n137 VDD.t174 378.788
R118 VDD.n132 VDD.t85 378.788
R119 VDD.t197 VDD.t221 303.031
R120 VDD.t218 VDD.t172 303.031
R121 VDD.t57 VDD.t129 303.031
R122 VDD.t82 VDD.t38 303.031
R123 VDD.t75 VDD.t78 303.031
R124 VDD.t200 VDD.t127 303.031
R125 VDD.t177 VDD.t20 303.031
R126 VDD.t28 VDD.t22 303.031
R127 VDD.t0 VDD.t190 303.031
R128 VDD.n206 VDD.t35 285.714
R129 VDD.n182 VDD.t61 285.714
R130 VDD.n153 VDD.t45 285.714
R131 VDD.n198 VDD.t3 242.857
R132 VDD.n200 VDD.t69 242.857
R133 VDD.t35 VDD.n202 242.857
R134 VDD.n205 VDD.t169 242.857
R135 VDD.n181 VDD.t158 242.857
R136 VDD.n183 VDD.t135 242.857
R137 VDD.n192 VDD.t61 242.857
R138 VDD.n193 VDD.t205 242.857
R139 VDD.n111 VDD.t192 242.857
R140 VDD.n112 VDD.t118 242.857
R141 VDD.t45 VDD.n152 242.857
R142 VDD.t180 VDD.n151 242.857
R143 VDD.n221 VDD.t72 193.183
R144 VDD.n223 VDD.t66 193.183
R145 VDD.n226 VDD.t197 193.183
R146 VDD.n229 VDD.t218 193.183
R147 VDD.n71 VDD.t147 193.183
R148 VDD.n77 VDD.t211 193.183
R149 VDD.n78 VDD.t52 193.183
R150 VDD.n83 VDD.t129 193.183
R151 VDD.n17 VDD.t142 193.183
R152 VDD.n19 VDD.t208 193.183
R153 VDD.n22 VDD.t82 193.183
R154 VDD.n25 VDD.t75 193.183
R155 VDD.n87 VDD.t152 193.183
R156 VDD.n89 VDD.t121 193.183
R157 VDD.n92 VDD.t200 193.183
R158 VDD.n95 VDD.t177 193.183
R159 VDD.n144 VDD.t155 193.183
R160 VDD.n142 VDD.t174 193.183
R161 VDD.n136 VDD.t85 193.183
R162 VDD.n157 VDD.t187 193.183
R163 VDD.n159 VDD.t132 193.183
R164 VDD.n162 VDD.t28 193.183
R165 VDD.n165 VDD.t0 193.183
R166 VDD.t44 VDD.t124 175.631
R167 VDD.t116 VDD.n127 153.678
R168 VDD.t10 VDD.n198 138.095
R169 VDD.t223 VDD.n200 138.095
R170 VDD.t26 VDD.n202 138.095
R171 VDD.t105 VDD.n205 138.095
R172 VDD.t59 VDD.n181 138.095
R173 VDD.n183 VDD.t24 138.095
R174 VDD.t55 VDD.n192 138.095
R175 VDD.n193 VDD.t145 138.095
R176 VDD.t138 VDD.n111 138.095
R177 VDD.n112 VDD.t125 138.095
R178 VDD.n152 VDD.t167 138.095
R179 VDD.n151 VDD.t96 138.095
R180 VDD.t163 VDD.n221 109.849
R181 VDD.t33 VDD.n223 109.849
R182 VDD.t8 VDD.n226 109.849
R183 VDD.n229 VDD.t102 109.849
R184 VDD.n71 VDD.t140 109.849
R185 VDD.t40 VDD.n77 109.849
R186 VDD.n78 VDD.t150 109.849
R187 VDD.t165 VDD.n83 109.849
R188 VDD.t110 VDD.n17 109.849
R189 VDD.t50 VDD.n19 109.849
R190 VDD.t31 VDD.n22 109.849
R191 VDD.n25 VDD.t93 109.849
R192 VDD.t12 VDD.n87 109.849
R193 VDD.t48 VDD.n89 109.849
R194 VDD.t90 VDD.n92 109.849
R195 VDD.n95 VDD.t99 109.849
R196 VDD.n144 VDD.t183 109.849
R197 VDD.t18 VDD.n142 109.849
R198 VDD.t80 VDD.n136 109.849
R199 VDD.t88 VDD.n157 109.849
R200 VDD.t64 VDD.n159 109.849
R201 VDD.t42 VDD.n162 109.849
R202 VDD.n165 VDD.t108 109.849
R203 VDD.n84 VDD.t14 59.702
R204 VDD.n143 VDD.t225 59.4064
R205 VDD.n137 VDD.t114 59.4064
R206 VDD.n132 VDD.t214 59.1138
R207 VDD.n128 VDD.t112 55.0852
R208 VDD.t216 VDD.n131 55.0852
R209 VDD.n26 VDD.t92 30.9379
R210 VDD.n28 VDD.t107 30.9379
R211 VDD.n49 VDD.t95 30.721
R212 VDD.n39 VDD.t104 30.7203
R213 VDD.n46 VDD.t98 30.3459
R214 VDD.n34 VDD.t101 30.0062
R215 VDD.n46 VDD.t231 24.8618
R216 VDD.n26 VDD.t232 24.5101
R217 VDD.n28 VDD.t227 24.5101
R218 VDD.n49 VDD.t229 24.4816
R219 VDD.n39 VDD.t228 24.4814
R220 VDD.n36 VDD.t230 24.4392
R221 VDD.n127 VDD.t44 21.9544
R222 VDD VDD.t203 10.5649
R223 VDD VDD.t16 10.5649
R224 VDD VDD.t185 10.5649
R225 VDD.n36 VDD.n35 8.0005
R226 VDD.n56 VDD.n55 6.39748
R227 VDD.n127 VDD 6.30126
R228 VDD.n209 VDD.n205 6.3005
R229 VDD.n212 VDD.n202 6.3005
R230 VDD.n215 VDD.n200 6.3005
R231 VDD.n218 VDD.n198 6.3005
R232 VDD.n230 VDD.n229 6.3005
R233 VDD.n233 VDD.n226 6.3005
R234 VDD.n236 VDD.n223 6.3005
R235 VDD.n239 VDD.n221 6.3005
R236 VDD.n59 VDD.n25 6.3005
R237 VDD.n62 VDD.n22 6.3005
R238 VDD.n65 VDD.n19 6.3005
R239 VDD.n68 VDD.n17 6.3005
R240 VDD.n83 VDD.n82 6.3005
R241 VDD.n79 VDD.n78 6.3005
R242 VDD.n77 VDD.n76 6.3005
R243 VDD.n72 VDD.n71 6.3005
R244 VDD.n96 VDD.n95 6.3005
R245 VDD.n99 VDD.n92 6.3005
R246 VDD.n102 VDD.n89 6.3005
R247 VDD.n105 VDD.n87 6.3005
R248 VDD VDD.n128 6.3005
R249 VDD.n131 VDD.n130 6.3005
R250 VDD.n136 VDD.n135 6.3005
R251 VDD.n142 VDD.n141 6.3005
R252 VDD.n145 VDD.n144 6.3005
R253 VDD.n151 VDD.n150 6.3005
R254 VDD.n152 VDD.n116 6.3005
R255 VDD.n113 VDD.n112 6.3005
R256 VDD.n111 VDD.n110 6.3005
R257 VDD.n166 VDD.n165 6.3005
R258 VDD.n169 VDD.n162 6.3005
R259 VDD.n172 VDD.n159 6.3005
R260 VDD.n175 VDD.n157 6.3005
R261 VDD.n194 VDD.n193 6.3005
R262 VDD.n192 VDD.n191 6.3005
R263 VDD.n184 VDD.n183 6.3005
R264 VDD.n181 VDD.n180 6.3005
R265 VDD.n45 VDD.n44 5.30657
R266 VDD.n230 VDD.t103 5.213
R267 VDD.n96 VDD.t100 5.213
R268 VDD.n166 VDD.t109 5.213
R269 VDD VDD.t204 5.16454
R270 VDD.n125 VDD.t217 5.14212
R271 VDD.n208 VDD.t106 5.13287
R272 VDD.n211 VDD.t27 5.13287
R273 VDD.n213 VDD.n201 5.13287
R274 VDD.n214 VDD.t224 5.13287
R275 VDD.n216 VDD.n199 5.13287
R276 VDD.n217 VDD.t11 5.13287
R277 VDD.n219 VDD.n197 5.13287
R278 VDD.n232 VDD.t9 5.13287
R279 VDD.n235 VDD.t34 5.13287
R280 VDD.n237 VDD.n222 5.13287
R281 VDD.n238 VDD.t164 5.13287
R282 VDD.n240 VDD.n220 5.13287
R283 VDD.n9 VDD.t166 5.13287
R284 VDD.n80 VDD.t151 5.13287
R285 VDD.n13 VDD.n12 5.13287
R286 VDD.n75 VDD.t41 5.13287
R287 VDD.n74 VDD.n14 5.13287
R288 VDD.n73 VDD.t141 5.13287
R289 VDD.n70 VDD.n15 5.13287
R290 VDD.n61 VDD.t32 5.13287
R291 VDD.n64 VDD.t51 5.13287
R292 VDD.n66 VDD.n18 5.13287
R293 VDD.n67 VDD.t111 5.13287
R294 VDD.n69 VDD.n16 5.13287
R295 VDD.n98 VDD.t91 5.13287
R296 VDD.n101 VDD.t49 5.13287
R297 VDD.n103 VDD.n88 5.13287
R298 VDD.n104 VDD.t13 5.13287
R299 VDD.n106 VDD.n86 5.13287
R300 VDD.n123 VDD.t81 5.13287
R301 VDD.n134 VDD.n124 5.13287
R302 VDD.n140 VDD.t19 5.13287
R303 VDD.n139 VDD.n122 5.13287
R304 VDD.n146 VDD.t184 5.13287
R305 VDD.n120 VDD.n119 5.13287
R306 VDD.n4 VDD.t97 5.13287
R307 VDD.n147 VDD.t168 5.13287
R308 VDD.n115 VDD.n5 5.13287
R309 VDD.n114 VDD.t126 5.13287
R310 VDD.n7 VDD.n6 5.13287
R311 VDD.n109 VDD.t139 5.13287
R312 VDD.n108 VDD.n8 5.13287
R313 VDD.n168 VDD.t43 5.13287
R314 VDD.n171 VDD.t65 5.13287
R315 VDD.n173 VDD.n158 5.13287
R316 VDD.n174 VDD.t89 5.13287
R317 VDD.n176 VDD.n156 5.13287
R318 VDD.n195 VDD.t146 5.13287
R319 VDD.n190 VDD.t56 5.13287
R320 VDD.n186 VDD.n0 5.13287
R321 VDD.n185 VDD.t25 5.13287
R322 VDD.n2 VDD.n1 5.13287
R323 VDD.n179 VDD.t60 5.13287
R324 VDD.n178 VDD.n3 5.13287
R325 VDD.n129 VDD.t113 5.09693
R326 VDD.n85 VDD.t15 5.09407
R327 VDD.n133 VDD.t215 5.09407
R328 VDD.n138 VDD.t115 5.09407
R329 VDD.n121 VDD.t226 5.09407
R330 VDD.n155 VDD.t186 5.09407
R331 VDD.n242 VDD.t17 5.09407
R332 VDD.n58 VDD.t94 4.8755
R333 VDD.n55 VDD.n45 4.84121
R334 VDD.n37 VDD.n36 4.5005
R335 VDD.n40 VDD.n38 4.5005
R336 VDD.n41 VDD.n38 4.5005
R337 VDD.n29 VDD.n27 4.5005
R338 VDD.n30 VDD.n27 4.5005
R339 VDD.n50 VDD.n48 4.5005
R340 VDD.n51 VDD.n48 4.5005
R341 VDD.n126 VDD.t117 3.94862
R342 VDD.n34 VDD.n33 3.61662
R343 VDD.n56 VDD.n26 2.88182
R344 VDD.n210 VDD.n204 2.85787
R345 VDD.n231 VDD.n228 2.85787
R346 VDD.n234 VDD.n225 2.85787
R347 VDD.n81 VDD.n11 2.85787
R348 VDD.n60 VDD.n24 2.85787
R349 VDD.n63 VDD.n21 2.85787
R350 VDD.n97 VDD.n94 2.85787
R351 VDD.n100 VDD.n91 2.85787
R352 VDD.n149 VDD.n118 2.85787
R353 VDD.n167 VDD.n164 2.85787
R354 VDD.n170 VDD.n161 2.85787
R355 VDD.n189 VDD.n188 2.85787
R356 VDD.n204 VDD.t7 2.2755
R357 VDD.n204 VDD.n203 2.2755
R358 VDD.n228 VDD.t173 2.2755
R359 VDD.n228 VDD.n227 2.2755
R360 VDD.n225 VDD.t222 2.2755
R361 VDD.n225 VDD.n224 2.2755
R362 VDD.n11 VDD.t58 2.2755
R363 VDD.n11 VDD.n10 2.2755
R364 VDD.n24 VDD.t79 2.2755
R365 VDD.n24 VDD.n23 2.2755
R366 VDD.n21 VDD.t39 2.2755
R367 VDD.n21 VDD.n20 2.2755
R368 VDD.n94 VDD.t21 2.2755
R369 VDD.n94 VDD.n93 2.2755
R370 VDD.n91 VDD.t128 2.2755
R371 VDD.n91 VDD.n90 2.2755
R372 VDD.n118 VDD.t196 2.2755
R373 VDD.n118 VDD.n117 2.2755
R374 VDD.n164 VDD.t191 2.2755
R375 VDD.n164 VDD.n163 2.2755
R376 VDD.n161 VDD.t23 2.2755
R377 VDD.n161 VDD.n160 2.2755
R378 VDD.n188 VDD.t162 2.2755
R379 VDD.n188 VDD.n187 2.2755
R380 VDD.n43 VDD.n42 2.2439
R381 VDD.n53 VDD.n52 2.2439
R382 VDD.n32 VDD.n31 2.24362
R383 VDD.n29 VDD.n28 2.12257
R384 VDD.n47 VDD.n46 1.81789
R385 VDD.n208 VDD 1.77285
R386 VDD VDD.n9 1.77285
R387 VDD VDD.n123 1.77285
R388 VDD.n140 VDD 1.77285
R389 VDD VDD.n4 1.77285
R390 VDD VDD.n195 1.77285
R391 VDD.n44 VDD.n43 1.62565
R392 VDD.n54 VDD.n53 1.62565
R393 VDD.n50 VDD.n49 1.39782
R394 VDD.n40 VDD.n39 1.39728
R395 VDD.n70 VDD.n69 1.16167
R396 VDD.n44 VDD.n37 1.12171
R397 VDD.n54 VDD.n47 1.12171
R398 VDD.n241 VDD.n240 1.07428
R399 VDD.n107 VDD.n106 1.07428
R400 VDD.n177 VDD.n176 1.07428
R401 VDD.n36 VDD.n34 0.840632
R402 VDD.n148 VDD.n146 0.715235
R403 VDD.n55 VDD.n54 0.5228
R404 VDD VDD.n126 0.498723
R405 VDD.n45 VDD.n32 0.497812
R406 VDD.n59 VDD.n58 0.337997
R407 VDD VDD.n125 0.334577
R408 VDD.n58 VDD.n57 0.333658
R409 VDD.n130 VDD.n129 0.317357
R410 VDD.n235 VDD.n234 0.233919
R411 VDD.n232 VDD.n231 0.233919
R412 VDD.n64 VDD.n63 0.233919
R413 VDD.n61 VDD.n60 0.233919
R414 VDD.n101 VDD.n100 0.233919
R415 VDD.n98 VDD.n97 0.233919
R416 VDD.n171 VDD.n170 0.233919
R417 VDD.n168 VDD.n167 0.233919
R418 VDD.n134 VDD.n133 0.170231
R419 VDD.n139 VDD.n138 0.170231
R420 VDD.n121 VDD.n120 0.170231
R421 VDD VDD.n126 0.16613
R422 VDD.n129 VDD 0.147133
R423 VDD.n241 VDD.n219 0.143501
R424 VDD.n108 VDD.n107 0.143501
R425 VDD.n178 VDD.n177 0.143501
R426 VDD.n217 VDD.n216 0.141016
R427 VDD.n214 VDD.n213 0.141016
R428 VDD.n238 VDD.n237 0.141016
R429 VDD.n67 VDD.n66 0.141016
R430 VDD.n74 VDD.n73 0.141016
R431 VDD.n75 VDD.n13 0.141016
R432 VDD.n104 VDD.n103 0.141016
R433 VDD.n109 VDD.n7 0.141016
R434 VDD.n115 VDD.n114 0.141016
R435 VDD.n174 VDD.n173 0.141016
R436 VDD.n179 VDD.n2 0.141016
R437 VDD.n186 VDD.n185 0.141016
R438 VDD.n107 VDD.n85 0.138896
R439 VDD.n177 VDD.n155 0.138896
R440 VDD.n242 VDD 0.127858
R441 VDD.n211 VDD 0.122435
R442 VDD VDD.n80 0.122435
R443 VDD.n190 VDD 0.122435
R444 VDD VDD.n210 0.111984
R445 VDD.n81 VDD 0.111984
R446 VDD.n149 VDD 0.111984
R447 VDD VDD.n189 0.111984
R448 VDD.n47 VDD 0.110941
R449 VDD.n219 VDD.n218 0.107339
R450 VDD.n216 VDD.n215 0.107339
R451 VDD.n213 VDD.n212 0.107339
R452 VDD.n240 VDD.n239 0.107339
R453 VDD.n237 VDD.n236 0.107339
R454 VDD.n69 VDD.n68 0.107339
R455 VDD.n66 VDD.n65 0.107339
R456 VDD.n72 VDD.n70 0.107339
R457 VDD.n76 VDD.n74 0.107339
R458 VDD.n79 VDD.n13 0.107339
R459 VDD.n106 VDD.n105 0.107339
R460 VDD.n103 VDD.n102 0.107339
R461 VDD.n135 VDD.n134 0.107339
R462 VDD.n141 VDD.n139 0.107339
R463 VDD.n145 VDD.n120 0.107339
R464 VDD.n110 VDD.n108 0.107339
R465 VDD.n113 VDD.n7 0.107339
R466 VDD.n116 VDD.n115 0.107339
R467 VDD.n176 VDD.n175 0.107339
R468 VDD.n173 VDD.n172 0.107339
R469 VDD.n180 VDD.n178 0.107339
R470 VDD.n184 VDD.n2 0.107339
R471 VDD.n191 VDD.n186 0.107339
R472 VDD.n210 VDD 0.106177
R473 VDD.n234 VDD 0.106177
R474 VDD.n231 VDD 0.106177
R475 VDD.n63 VDD 0.106177
R476 VDD.n60 VDD 0.106177
R477 VDD VDD.n81 0.106177
R478 VDD.n100 VDD 0.106177
R479 VDD.n97 VDD 0.106177
R480 VDD VDD.n149 0.106177
R481 VDD.n170 VDD 0.106177
R482 VDD.n167 VDD 0.106177
R483 VDD.n189 VDD 0.106177
R484 VDD.n35 VDD 0.0839415
R485 VDD VDD.n148 0.082371
R486 VDD.n41 VDD 0.0816915
R487 VDD.n209 VDD.n208 0.080629
R488 VDD.n233 VDD.n232 0.080629
R489 VDD.n62 VDD.n61 0.080629
R490 VDD.n82 VDD.n9 0.080629
R491 VDD.n99 VDD.n98 0.080629
R492 VDD.n150 VDD.n4 0.080629
R493 VDD.n169 VDD.n168 0.080629
R494 VDD.n195 VDD.n194 0.080629
R495 VDD.n51 VDD 0.0805665
R496 VDD VDD.n217 0.0794677
R497 VDD VDD.n214 0.0794677
R498 VDD VDD.n211 0.0794677
R499 VDD VDD.n238 0.0794677
R500 VDD VDD.n235 0.0794677
R501 VDD VDD.n67 0.0794677
R502 VDD VDD.n64 0.0794677
R503 VDD.n73 VDD 0.0794677
R504 VDD VDD.n75 0.0794677
R505 VDD.n80 VDD 0.0794677
R506 VDD VDD.n104 0.0794677
R507 VDD VDD.n101 0.0794677
R508 VDD VDD.n109 0.0794677
R509 VDD.n114 VDD 0.0794677
R510 VDD.n147 VDD 0.0794677
R511 VDD VDD.n174 0.0794677
R512 VDD VDD.n171 0.0794677
R513 VDD VDD.n179 0.0794677
R514 VDD.n185 VDD 0.0794677
R515 VDD VDD.n190 0.0794677
R516 VDD VDD.n125 0.0794623
R517 VDD VDD.n123 0.0759839
R518 VDD VDD.n140 0.0759839
R519 VDD.n146 VDD 0.0759839
R520 VDD.n30 VDD 0.0738165
R521 VDD.n57 VDD.n56 0.0725
R522 VDD.n85 VDD 0.0709717
R523 VDD.n133 VDD 0.0709717
R524 VDD.n138 VDD 0.0709717
R525 VDD VDD.n121 0.0709717
R526 VDD.n155 VDD 0.0709717
R527 VDD VDD.n242 0.0709717
R528 VDD.n57 VDD 0.0493298
R529 VDD.n148 VDD.n147 0.0405645
R530 VDD.n42 VDD.n41 0.0275
R531 VDD.n35 VDD.n33 0.0275
R532 VDD.n52 VDD.n51 0.026375
R533 VDD.n43 VDD.n38 0.025705
R534 VDD.n53 VDD.n48 0.025705
R535 VDD.n31 VDD.n30 0.02075
R536 VDD.n32 VDD.n27 0.0169383
R537 VDD VDD.n241 0.0115377
R538 VDD.n31 VDD.n29 0.0095
R539 VDD.n135 VDD 0.00514516
R540 VDD.n141 VDD 0.00514516
R541 VDD VDD.n145 0.00514516
R542 VDD.n52 VDD.n50 0.003875
R543 VDD.n42 VDD.n40 0.00275
R544 VDD.n130 VDD 0.00219811
R545 VDD.n218 VDD 0.00166129
R546 VDD.n215 VDD 0.00166129
R547 VDD.n212 VDD 0.00166129
R548 VDD VDD.n209 0.00166129
R549 VDD.n239 VDD 0.00166129
R550 VDD.n236 VDD 0.00166129
R551 VDD VDD.n233 0.00166129
R552 VDD VDD.n230 0.00166129
R553 VDD.n68 VDD 0.00166129
R554 VDD.n65 VDD 0.00166129
R555 VDD VDD.n62 0.00166129
R556 VDD VDD.n59 0.00166129
R557 VDD VDD.n72 0.00166129
R558 VDD.n76 VDD 0.00166129
R559 VDD VDD.n79 0.00166129
R560 VDD.n82 VDD 0.00166129
R561 VDD.n105 VDD 0.00166129
R562 VDD.n102 VDD 0.00166129
R563 VDD VDD.n99 0.00166129
R564 VDD VDD.n96 0.00166129
R565 VDD.n110 VDD 0.00166129
R566 VDD VDD.n113 0.00166129
R567 VDD VDD.n116 0.00166129
R568 VDD.n150 VDD 0.00166129
R569 VDD.n175 VDD 0.00166129
R570 VDD.n172 VDD 0.00166129
R571 VDD VDD.n169 0.00166129
R572 VDD VDD.n166 0.00166129
R573 VDD.n180 VDD 0.00166129
R574 VDD VDD.n184 0.00166129
R575 VDD.n191 VDD 0.00166129
R576 VDD.n194 VDD 0.00166129
R577 VDD.n37 VDD.n33 0.001625
R578 CLK.n9 CLK.t0 36.935
R579 CLK.n3 CLK.t1 36.935
R580 CLK.n14 CLK.t3 25.5361
R581 CLK.n9 CLK.t2 18.1962
R582 CLK.n3 CLK.t5 18.1962
R583 CLK.n14 CLK.t4 14.0734
R584 CLK.n5 CLK.n2 4.5005
R585 CLK.n5 CLK.n4 4.5005
R586 CLK.n8 CLK.n7 4.5005
R587 CLK.n10 CLK.n7 4.5005
R588 CLK.n16 CLK.n15 4.5005
R589 CLK.n17 CLK.n16 4.5005
R590 CLK.n12 CLK.n11 2.25107
R591 CLK.n13 CLK.n0 2.24235
R592 CLK.n4 CLK.n3 2.12175
R593 CLK.n10 CLK.n9 2.12075
R594 CLK.n7 CLK.n6 1.74297
R595 CLK.n6 CLK.n1 1.49778
R596 CLK.n15 CLK.n14 1.42775
R597 CLK.n13 CLK.n12 0.97145
R598 CLK CLK.n17 0.158
R599 CLK.n8 CLK 0.0473512
R600 CLK.n2 CLK 0.0473512
R601 CLK.n11 CLK.n8 0.0361897
R602 CLK.n2 CLK.n1 0.0361897
R603 CLK.n17 CLK.n0 0.03175
R604 CLK.n16 CLK.n13 0.0246174
R605 CLK.n6 CLK.n5 0.0131772
R606 CLK.n12 CLK.n7 0.0122182
R607 CLK.n11 CLK.n10 0.00515517
R608 CLK.n4 CLK.n1 0.00515517
R609 CLK.n15 CLK.n0 0.00175
R610 VSS.n79 VSS.n74 18801.2
R611 VSS.n114 VSS.t71 6810.9
R612 VSS.n40 VSS.t92 6265.15
R613 VSS.n55 VSS.n12 3893.61
R614 VSS.n78 VSS.n75 3893.61
R615 VSS.n100 VSS.n97 3893.61
R616 VSS.n14 VSS.t81 3606.54
R617 VSS.n13 VSS.t85 3112.87
R618 VSS.t133 VSS.t135 3055.32
R619 VSS.n12 VSS.t67 2628.58
R620 VSS.n75 VSS.t69 2628.58
R621 VSS.n97 VSS.t75 2628.58
R622 VSS.n12 VSS.t24 2622.37
R623 VSS.n75 VSS.t121 2622.37
R624 VSS.n97 VSS.t115 2622.37
R625 VSS.t132 VSS.t79 2510.52
R626 VSS.t59 VSS.t27 2510.52
R627 VSS.t87 VSS.t9 2510.52
R628 VSS.t62 VSS.t65 2510.52
R629 VSS.t95 VSS.t63 2510.52
R630 VSS.t124 VSS.t35 2510.52
R631 VSS.t58 VSS.t109 2510.52
R632 VSS.t94 VSS.t4 2510.52
R633 VSS.t140 VSS.t25 2307.56
R634 VSS.t99 VSS.t131 2307.56
R635 VSS.t47 VSS.t33 2307.56
R636 VSS.t0 VSS.t111 2307.56
R637 VSS.t88 VSS.t97 2307.56
R638 VSS.t89 VSS.t42 2307.56
R639 VSS.t126 VSS.t113 2307.56
R640 VSS.t96 VSS.t52 2307.56
R641 VSS.t19 VSS.t54 2307.56
R642 VSS.t107 VSS.t48 2307.56
R643 VSS.t57 VSS.t7 2307.56
R644 VSS.t138 VSS.t29 2307.56
R645 VSS.t2 VSS.t21 2307.56
R646 VSS.t37 VSS.n40 2084.8
R647 VSS.t125 VSS.n56 1713.53
R648 VSS.t108 VSS.n79 1713.53
R649 VSS.t3 VSS.n101 1713.53
R650 VSS.n56 VSS.n55 1565.03
R651 VSS.n79 VSS.n78 1565.03
R652 VSS.n101 VSS.n100 1565.03
R653 VSS.t92 VSS.t39 1151.9
R654 VSS.t127 VSS.t32 994.264
R655 VSS.t17 VSS.t59 994.264
R656 VSS.t128 VSS.t91 994.264
R657 VSS.t116 VSS.t62 994.264
R658 VSS.t129 VSS.t18 994.264
R659 VSS.t130 VSS.t124 994.264
R660 VSS.t23 VSS.t137 994.264
R661 VSS.t105 VSS.t94 994.264
R662 VSS.t16 VSS.t38 913.885
R663 VSS.t119 VSS.t126 913.885
R664 VSS.t60 VSS.t107 913.885
R665 VSS.t106 VSS.t2 913.885
R666 VSS.n27 VSS.t83 838.187
R667 VSS.t39 VSS.n39 671.942
R668 VSS.n3 VSS.t6 596.558
R669 VSS.n4 VSS.t132 596.558
R670 VSS.n5 VSS.t127 596.558
R671 VSS.n6 VSS.t17 596.558
R672 VSS.t24 VSS.n8 596.558
R673 VSS.n9 VSS.t87 596.558
R674 VSS.n10 VSS.t128 596.558
R675 VSS.n11 VSS.t116 596.558
R676 VSS.t121 VSS.n70 596.558
R677 VSS.n71 VSS.t95 596.558
R678 VSS.n72 VSS.t129 596.558
R679 VSS.n73 VSS.t130 596.558
R680 VSS.t115 VSS.n93 596.558
R681 VSS.n94 VSS.t58 596.558
R682 VSS.n95 VSS.t23 596.558
R683 VSS.n96 VSS.t105 596.558
R684 VSS.n16 VSS.t61 548.331
R685 VSS.n17 VSS.t120 548.331
R686 VSS.n19 VSS.t15 548.331
R687 VSS.n41 VSS.t37 548.331
R688 VSS.n46 VSS.t131 548.331
R689 VSS.n47 VSS.t47 548.331
R690 VSS.n52 VSS.t16 548.331
R691 VSS.n59 VSS.t125 548.331
R692 VSS.n60 VSS.t88 548.331
R693 VSS.n65 VSS.t42 548.331
R694 VSS.n66 VSS.t119 548.331
R695 VSS.n82 VSS.t108 548.331
R696 VSS.n83 VSS.t96 548.331
R697 VSS.n88 VSS.t54 548.331
R698 VSS.n89 VSS.t60 548.331
R699 VSS.n104 VSS.t3 548.331
R700 VSS.n105 VSS.t57 548.331
R701 VSS.n110 VSS.t29 548.331
R702 VSS.n111 VSS.t106 548.331
R703 VSS.n39 VSS.t85 479.959
R704 VSS.t79 VSS.n3 397.707
R705 VSS.n4 VSS.t45 397.707
R706 VSS.t27 VSS.n5 397.707
R707 VSS.t67 VSS.n6 397.707
R708 VSS.t9 VSS.n8 397.707
R709 VSS.n9 VSS.t43 397.707
R710 VSS.t65 VSS.n10 397.707
R711 VSS.t69 VSS.n11 397.707
R712 VSS.t63 VSS.n70 397.707
R713 VSS.n71 VSS.t55 397.707
R714 VSS.t35 VSS.n72 397.707
R715 VSS.t75 VSS.n73 397.707
R716 VSS.t109 VSS.n93 397.707
R717 VSS.n94 VSS.t30 397.707
R718 VSS.t4 VSS.n95 397.707
R719 VSS.t71 VSS.n96 397.707
R720 VSS.t13 VSS.n16 365.555
R721 VSS.t25 VSS.n17 365.555
R722 VSS.n19 VSS.t122 365.555
R723 VSS.n41 VSS.t99 365.555
R724 VSS.t33 VSS.n46 365.555
R725 VSS.n47 VSS.t101 365.555
R726 VSS.t111 VSS.n52 365.555
R727 VSS.t97 VSS.n59 365.555
R728 VSS.n60 VSS.t89 365.555
R729 VSS.t113 VSS.n65 365.555
R730 VSS.n66 VSS.t73 365.555
R731 VSS.t52 VSS.n82 365.555
R732 VSS.n83 VSS.t19 365.555
R733 VSS.t48 VSS.n88 365.555
R734 VSS.n89 VSS.t50 365.555
R735 VSS.t7 VSS.n104 365.555
R736 VSS.n105 VSS.t138 365.555
R737 VSS.t21 VSS.n110 365.555
R738 VSS.n111 VSS.t77 365.555
R739 VSS.n26 VSS.t13 165.642
R740 VSS.t81 VSS.n13 150.845
R741 VSS.t135 VSS.n14 150.845
R742 VSS.n55 VSS.n54 119.948
R743 VSS.n78 VSS.n77 119.948
R744 VSS.n100 VSS.n99 119.948
R745 VSS.n15 VSS.t133 34.2711
R746 VSS.n18 VSS.t140 34.2711
R747 VSS.n54 VSS.t0 34.2711
R748 VSS.n77 VSS.t117 34.2711
R749 VSS.n99 VSS.t11 34.2711
R750 VSS.n27 VSS.n26 27.0388
R751 VSS.n114 VSS.t103 22.8476
R752 VSS.n115 VSS.n114 16.6241
R753 VSS.n37 VSS.t86 9.37686
R754 VSS.n115 VSS.t104 9.3736
R755 VSS.n98 VSS.t12 9.3736
R756 VSS.n76 VSS.t118 9.3736
R757 VSS.n53 VSS.t1 9.3736
R758 VSS.n31 VSS.t134 9.30652
R759 VSS.n25 VSS.t84 9.30652
R760 VSS.n21 VSS.t141 9.30652
R761 VSS.n35 VSS.t82 9.30518
R762 VSS.n33 VSS.t136 9.25414
R763 VSS VSS.t123 7.30633
R764 VSS.n150 VSS.t80 7.19156
R765 VSS.n148 VSS.t46 7.19156
R766 VSS.n141 VSS.t10 7.19156
R767 VSS.n139 VSS.t44 7.19156
R768 VSS.n132 VSS.t64 7.19156
R769 VSS.n130 VSS.t56 7.19156
R770 VSS.n123 VSS.t110 7.19156
R771 VSS.n121 VSS.t31 7.19156
R772 VSS.n80 VSS.t53 7.19156
R773 VSS.n85 VSS.t20 7.19156
R774 VSS.n86 VSS.t49 7.19156
R775 VSS.n57 VSS.t98 7.19156
R776 VSS.n62 VSS.t90 7.19156
R777 VSS.n63 VSS.t114 7.19156
R778 VSS.n43 VSS.t100 7.19156
R779 VSS.n44 VSS.t34 7.19156
R780 VSS.n49 VSS.t102 7.19156
R781 VSS.n102 VSS.t8 7.19156
R782 VSS.n107 VSS.t139 7.19156
R783 VSS.n108 VSS.t22 7.19156
R784 VSS.n29 VSS.t14 6.88656
R785 VSS.n23 VSS.t26 6.88656
R786 VSS.n1 VSS.n0 6.01414
R787 VSS.n1 VSS.t93 6.01414
R788 VSS.n146 VSS.t28 5.91399
R789 VSS.n144 VSS.t68 5.91399
R790 VSS.n137 VSS.t66 5.91399
R791 VSS.n135 VSS.t70 5.91399
R792 VSS.n128 VSS.t36 5.91399
R793 VSS.n126 VSS.t76 5.91399
R794 VSS.n119 VSS.t5 5.91399
R795 VSS.n117 VSS.t72 5.91399
R796 VSS.n91 VSS.t51 5.91399
R797 VSS.n68 VSS.t74 5.91399
R798 VSS.n50 VSS.t112 5.91399
R799 VSS.n113 VSS.t78 5.91399
R800 VSS.n39 VSS.n38 5.2005
R801 VSS.n36 VSS.n13 5.2005
R802 VSS.n34 VSS.n14 5.2005
R803 VSS.n32 VSS.n15 5.2005
R804 VSS.n30 VSS.n16 5.2005
R805 VSS.n28 VSS.n27 5.2005
R806 VSS.n22 VSS.n18 5.2005
R807 VSS.n20 VSS.n19 5.2005
R808 VSS.n24 VSS.n17 5.2005
R809 VSS.n42 VSS.n41 5.2005
R810 VSS.n46 VSS.n45 5.2005
R811 VSS.n48 VSS.n47 5.2005
R812 VSS.n52 VSS.n51 5.2005
R813 VSS.n54 VSS.n53 5.2005
R814 VSS.n59 VSS.n58 5.2005
R815 VSS.n61 VSS.n60 5.2005
R816 VSS.n65 VSS.n64 5.2005
R817 VSS.n67 VSS.n66 5.2005
R818 VSS.n77 VSS.n76 5.2005
R819 VSS.n82 VSS.n81 5.2005
R820 VSS.n84 VSS.n83 5.2005
R821 VSS.n88 VSS.n87 5.2005
R822 VSS.n90 VSS.n89 5.2005
R823 VSS.n99 VSS.n98 5.2005
R824 VSS.n104 VSS.n103 5.2005
R825 VSS.n106 VSS.n105 5.2005
R826 VSS.n110 VSS.n109 5.2005
R827 VSS.n112 VSS.n111 5.2005
R828 VSS.n118 VSS.n96 5.2005
R829 VSS.n120 VSS.n95 5.2005
R830 VSS.n122 VSS.n94 5.2005
R831 VSS.n124 VSS.n93 5.2005
R832 VSS.n127 VSS.n73 5.2005
R833 VSS.n129 VSS.n72 5.2005
R834 VSS.n131 VSS.n71 5.2005
R835 VSS.n133 VSS.n70 5.2005
R836 VSS.n136 VSS.n11 5.2005
R837 VSS.n138 VSS.n10 5.2005
R838 VSS.n140 VSS.n9 5.2005
R839 VSS.n142 VSS.n8 5.2005
R840 VSS.n145 VSS.n6 5.2005
R841 VSS.n147 VSS.n5 5.2005
R842 VSS.n149 VSS.n4 5.2005
R843 VSS.n151 VSS.n3 5.2005
R844 VSS.n2 VSS.n1 3.36323
R845 VSS VSS.n2 2.40845
R846 VSS.n117 VSS.n116 1.03335
R847 VSS.n125 VSS.n92 0.845914
R848 VSS.n134 VSS.n69 0.845914
R849 VSS.n143 VSS.n7 0.845914
R850 VSS.n143 VSS 0.519858
R851 VSS.n134 VSS 0.519858
R852 VSS.n148 VSS.n147 0.480225
R853 VSS.n146 VSS.n145 0.480225
R854 VSS.n139 VSS.n138 0.480225
R855 VSS.n137 VSS.n136 0.480225
R856 VSS.n130 VSS.n129 0.480225
R857 VSS.n128 VSS.n127 0.480225
R858 VSS.n121 VSS.n120 0.480225
R859 VSS.n119 VSS.n118 0.480225
R860 VSS.n31 VSS.n30 0.396455
R861 VSS.n21 VSS.n20 0.396455
R862 VSS.n25 VSS.n24 0.396455
R863 VSS.n37 VSS 0.379596
R864 VSS.n80 VSS 0.343161
R865 VSS VSS.n85 0.343161
R866 VSS.n57 VSS 0.343161
R867 VSS VSS.n62 0.343161
R868 VSS VSS.n43 0.343161
R869 VSS.n44 VSS 0.343161
R870 VSS.n102 VSS 0.343161
R871 VSS VSS.n107 0.343161
R872 VSS.n150 VSS 0.343161
R873 VSS.n141 VSS 0.343161
R874 VSS.n132 VSS 0.343161
R875 VSS.n123 VSS 0.343161
R876 VSS.n35 VSS 0.310668
R877 VSS.n90 VSS 0.289491
R878 VSS.n67 VSS 0.289491
R879 VSS.n51 VSS 0.289491
R880 VSS.n112 VSS 0.289491
R881 VSS.n23 VSS 0.27984
R882 VSS.n29 VSS 0.27984
R883 VSS.n33 VSS 0.250123
R884 VSS.n34 VSS.n33 0.247195
R885 VSS VSS.n29 0.243604
R886 VSS VSS.n23 0.243604
R887 VSS.n125 VSS 0.21683
R888 VSS.n86 VSS 0.191234
R889 VSS.n63 VSS 0.191234
R890 VSS VSS.n49 0.191234
R891 VSS.n108 VSS 0.191234
R892 VSS.n144 VSS.n143 0.187931
R893 VSS.n135 VSS.n134 0.187931
R894 VSS.n126 VSS.n125 0.187931
R895 VSS.n36 VSS.n35 0.152211
R896 VSS.n38 VSS.n2 0.138903
R897 VSS.n116 VSS 0.137685
R898 VSS VSS.n92 0.137685
R899 VSS VSS.n69 0.137685
R900 VSS VSS.n7 0.137685
R901 VSS.n81 VSS.n80 0.118573
R902 VSS.n85 VSS.n84 0.118573
R903 VSS.n87 VSS.n86 0.118573
R904 VSS.n58 VSS.n57 0.118573
R905 VSS.n62 VSS.n61 0.118573
R906 VSS.n64 VSS.n63 0.118573
R907 VSS.n43 VSS.n42 0.118573
R908 VSS.n45 VSS.n44 0.118573
R909 VSS.n49 VSS.n48 0.118573
R910 VSS.n103 VSS.n102 0.118573
R911 VSS.n107 VSS.n106 0.118573
R912 VSS.n109 VSS.n108 0.118573
R913 VSS.n151 VSS.n150 0.118573
R914 VSS.n149 VSS.n148 0.118573
R915 VSS.n142 VSS.n141 0.118573
R916 VSS.n140 VSS.n139 0.118573
R917 VSS.n133 VSS.n132 0.118573
R918 VSS.n131 VSS.n130 0.118573
R919 VSS.n124 VSS.n123 0.118573
R920 VSS.n122 VSS.n121 0.118573
R921 VSS.n91 VSS 0.115271
R922 VSS.n68 VSS 0.115271
R923 VSS VSS.n50 0.115271
R924 VSS.n113 VSS 0.115271
R925 VSS VSS.n146 0.115271
R926 VSS VSS.n144 0.115271
R927 VSS VSS.n137 0.115271
R928 VSS VSS.n135 0.115271
R929 VSS VSS.n128 0.115271
R930 VSS VSS.n126 0.115271
R931 VSS VSS.n119 0.115271
R932 VSS VSS.n117 0.115271
R933 VSS VSS.n37 0.113945
R934 VSS.n92 VSS.n91 0.10206
R935 VSS.n69 VSS.n68 0.10206
R936 VSS.n50 VSS.n7 0.10206
R937 VSS.n116 VSS.n113 0.10206
R938 VSS.n32 VSS.n31 0.0675755
R939 VSS.n22 VSS.n21 0.0675755
R940 VSS.n28 VSS.n25 0.0675755
R941 VSS.n81 VSS 0.00545413
R942 VSS.n84 VSS 0.00545413
R943 VSS.n87 VSS 0.00545413
R944 VSS.n58 VSS 0.00545413
R945 VSS.n61 VSS 0.00545413
R946 VSS.n64 VSS 0.00545413
R947 VSS.n42 VSS 0.00545413
R948 VSS.n45 VSS 0.00545413
R949 VSS.n48 VSS 0.00545413
R950 VSS.n103 VSS 0.00545413
R951 VSS.n106 VSS 0.00545413
R952 VSS.n109 VSS 0.00545413
R953 VSS VSS.n151 0.00545413
R954 VSS VSS.n149 0.00545413
R955 VSS VSS.n142 0.00545413
R956 VSS VSS.n140 0.00545413
R957 VSS VSS.n133 0.00545413
R958 VSS VSS.n131 0.00545413
R959 VSS VSS.n124 0.00545413
R960 VSS VSS.n122 0.00545413
R961 VSS VSS.n90 0.00380275
R962 VSS VSS.n67 0.00380275
R963 VSS.n51 VSS 0.00380275
R964 VSS.n30 VSS 0.00380275
R965 VSS.n20 VSS 0.00380275
R966 VSS.n24 VSS 0.00380275
R967 VSS VSS.n112 0.00380275
R968 VSS.n147 VSS 0.00380275
R969 VSS.n145 VSS 0.00380275
R970 VSS.n138 VSS 0.00380275
R971 VSS.n136 VSS 0.00380275
R972 VSS.n129 VSS 0.00380275
R973 VSS.n127 VSS 0.00380275
R974 VSS.n120 VSS 0.00380275
R975 VSS.n118 VSS 0.00380275
R976 VSS.n38 VSS 0.00352521
R977 VSS VSS.n115 0.00219811
R978 VSS.n98 VSS 0.00219811
R979 VSS.n76 VSS 0.00219811
R980 VSS.n53 VSS 0.00219811
R981 VSS VSS.n36 0.00219811
R982 VSS VSS.n34 0.00219811
R983 VSS VSS.n32 0.00219811
R984 VSS VSS.n22 0.00219811
R985 VSS VSS.n28 0.00219811
R986 Q0.n33 Q0.t10 36.935
R987 Q0.n16 Q0.t6 36.935
R988 Q0.n9 Q0.t7 36.935
R989 Q0.n47 Q0.t15 36.935
R990 Q0.n0 Q0.t18 36.935
R991 Q0.n35 Q0.t9 31.528
R992 Q0.n22 Q0.t14 30.7203
R993 Q0.n40 Q0.t4 25.5364
R994 Q0.n3 Q0.t12 25.5364
R995 Q0.n22 Q0.t5 21.6135
R996 Q0.n33 Q0.t8 18.1962
R997 Q0.n16 Q0.t11 18.1962
R998 Q0.n9 Q0.t3 18.1962
R999 Q0.n47 Q0.t19 18.1962
R1000 Q0.n0 Q0.t16 18.1962
R1001 Q0.n35 Q0.t20 15.3826
R1002 Q0.n40 Q0.t13 14.0749
R1003 Q0.n3 Q0.t17 14.0749
R1004 Q0.n45 Q0.n27 9.89892
R1005 Q0.n31 Q0.n28 7.09905
R1006 Q0.n36 Q0.n35 6.86134
R1007 Q0.n27 Q0.n26 6.01475
R1008 Q0.n37 Q0.n34 5.01116
R1009 Q0.n31 Q0.n30 3.25085
R1010 Q0.n30 Q0.t1 2.2755
R1011 Q0.n30 Q0.n29 2.2755
R1012 Q0.n19 Q0.n18 2.25107
R1013 Q0.n50 Q0.n49 2.25107
R1014 Q0.n38 Q0.n32 2.2505
R1015 Q0.n26 Q0.n25 2.24299
R1016 Q0.n7 Q0.n6 2.24235
R1017 Q0.n44 Q0.n43 2.24235
R1018 Q0.n34 Q0.n33 2.13398
R1019 Q0.n10 Q0.n9 2.12175
R1020 Q0.n1 Q0.n0 2.12175
R1021 Q0.n17 Q0.n16 2.12075
R1022 Q0.n48 Q0.n47 2.12075
R1023 Q0.n14 Q0.n13 1.74297
R1024 Q0.n53 Q0.n51 1.74297
R1025 Q0.n38 Q0.n37 1.5289
R1026 Q0.n13 Q0.n11 1.49778
R1027 Q0.n54 Q0.n53 1.49778
R1028 Q0.n41 Q0.n40 1.42706
R1029 Q0.n4 Q0.n3 1.42706
R1030 Q0.n23 Q0.n22 1.3985
R1031 Q0.n50 Q0.n45 1.1676
R1032 Q0.n37 Q0.n36 1.12056
R1033 Q0.n20 Q0.n19 0.928385
R1034 Q0.n39 Q0 0.628836
R1035 Q0.n27 Q0.n20 0.286289
R1036 Q0.n42 Q0 0.1605
R1037 Q0.n5 Q0 0.1605
R1038 Q0.n32 Q0.n31 0.0919062
R1039 Q0.n36 Q0 0.0857632
R1040 Q0.n34 Q0 0.0810725
R1041 Q0.n24 Q0 0.0805665
R1042 Q0.n32 Q0 0.073625
R1043 Q0.n15 Q0 0.0473512
R1044 Q0.n8 Q0 0.0473512
R1045 Q0.n46 Q0 0.0473512
R1046 Q0 Q0.n55 0.0473512
R1047 Q0.n20 Q0.n7 0.0435648
R1048 Q0.n18 Q0.n15 0.0361897
R1049 Q0.n11 Q0.n8 0.0361897
R1050 Q0.n49 Q0.n46 0.0361897
R1051 Q0.n55 Q0.n54 0.0361897
R1052 Q0.n43 Q0.n42 0.03175
R1053 Q0.n6 Q0.n5 0.03175
R1054 Q0 Q0.n38 0.0289903
R1055 Q0.n45 Q0.n44 0.0277753
R1056 Q0.n25 Q0.n24 0.0275
R1057 Q0.n26 Q0.n21 0.0266571
R1058 Q0.n7 Q0.n2 0.0246174
R1059 Q0.n44 Q0.n39 0.0246174
R1060 Q0.n13 Q0.n12 0.0131772
R1061 Q0.n53 Q0.n52 0.0131772
R1062 Q0.n19 Q0.n14 0.0122182
R1063 Q0.n51 Q0.n50 0.0122182
R1064 Q0.n18 Q0.n17 0.00515517
R1065 Q0.n11 Q0.n10 0.00515517
R1066 Q0.n49 Q0.n48 0.00515517
R1067 Q0.n54 Q0.n1 0.00515517
R1068 Q0.n25 Q0.n23 0.00275
R1069 Q0.n43 Q0.n41 0.00175
R1070 Q0.n6 Q0.n4 0.00175
R1071 JK_FF_mag_2.J.n2 JK_FF_mag_2.J.t6 37.1986
R1072 JK_FF_mag_2.J.n1 JK_FF_mag_2.J.t5 31.528
R1073 JK_FF_mag_2.J.n3 JK_FF_mag_2.J.t3 30.6315
R1074 JK_FF_mag_2.J.n3 JK_FF_mag_2.J.t7 24.5953
R1075 JK_FF_mag_2.J.n2 JK_FF_mag_2.J.t8 17.6614
R1076 JK_FF_mag_2.J.n4 JK_FF_mag_2.J 17.0516
R1077 JK_FF_mag_2.J.n1 JK_FF_mag_2.J.t4 15.3826
R1078 JK_FF_mag_2.J JK_FF_mag_2.J.n1 7.62751
R1079 JK_FF_mag_2.J.n5 JK_FF_mag_2.J.n4 3.28711
R1080 JK_FF_mag_2.J.n0 JK_FF_mag_2.J.n7 2.99416
R1081 JK_FF_mag_2.J.n4 JK_FF_mag_2.J 2.81128
R1082 JK_FF_mag_2.J.n5 JK_FF_mag_2.J 2.67866
R1083 JK_FF_mag_2.J.n7 JK_FF_mag_2.J.t2 2.2755
R1084 JK_FF_mag_2.J.n7 JK_FF_mag_2.J.n6 2.2755
R1085 JK_FF_mag_2.J.n0 JK_FF_mag_2.J.n5 2.2505
R1086 JK_FF_mag_2.J JK_FF_mag_2.J.n3 1.80496
R1087 JK_FF_mag_2.J JK_FF_mag_2.J.n2 1.43709
R1088 JK_FF_mag_2.J JK_FF_mag_2.J.n0 0.290136
R1089 Vdiv10.n4 Vdiv10.n3 9.28675
R1090 Vdiv10.n2 Vdiv10.n1 6.01414
R1091 Vdiv10.n2 Vdiv10.t0 6.01414
R1092 Vdiv10.n5 Vdiv10.n0 3.87666
R1093 Vdiv10.n4 Vdiv10.n2 3.74699
R1094 Vdiv10.n5 Vdiv10.n4 0.0409348
R1095 Vdiv10 Vdiv10.n5 0.0031087
R1096 RST.n10 RST.t7 36.935
R1097 RST.n12 RST.t2 36.935
R1098 RST.n0 RST.t3 36.935
R1099 RST.n5 RST.t5 36.859
R1100 RST.n10 RST.t6 18.1962
R1101 RST.n12 RST.t0 18.1962
R1102 RST.n0 RST.t1 18.1962
R1103 RST.n4 RST.t4 17.236
R1104 RST.n14 RST.n13 5.39891
R1105 RST.n9 RST.n8 4.5005
R1106 RST.n3 RST.n2 4.5005
R1107 RST.n9 RST.n1 4.5005
R1108 RST.n4 RST.n1 3.60685
R1109 RST.n15 RST.n14 3.52872
R1110 RST RST.n15 3.47443
R1111 RST.n6 RST.n5 2.88526
R1112 RST.n13 RST.n12 2.13713
R1113 RST.n11 RST.n10 2.13713
R1114 RST.n16 RST.n0 2.13533
R1115 RST.n14 RST.n11 1.87041
R1116 RST.n16 RST 1.81616
R1117 RST.n7 RST.n2 1.51223
R1118 RST.n15 RST.n9 1.12371
R1119 RST.n5 RST.n4 0.865351
R1120 RST RST.n16 0.0693483
R1121 RST.n11 RST 0.06755
R1122 RST.n13 RST 0.0675495
R1123 RST.n3 RST 0.0394837
R1124 RST.n8 RST.n7 0.0367013
R1125 RST.n7 RST.n6 0.0051456
R1126 RST.n9 RST.n2 0.003875
R1127 RST.n8 RST.n3 0.00205172
R1128 RST.n6 RST.n1 0.00199457
R1129 Q2.n8 Q2.t7 36.935
R1130 Q2.n2 Q2.t3 31.528
R1131 Q2.n5 Q2.t12 31.528
R1132 Q2.n10 Q2.t10 31.528
R1133 Q2.n0 Q2.t4 30.6315
R1134 Q2.n0 Q2.t11 21.7275
R1135 Q2.n8 Q2.t5 18.1962
R1136 Q2.n2 Q2.t9 15.3826
R1137 Q2.n5 Q2.t6 15.3826
R1138 Q2.n10 Q2.t8 15.3826
R1139 Q2.n17 Q2.n14 7.09905
R1140 Q2.n6 Q2.n5 6.86647
R1141 Q2.n3 Q2.n2 6.86646
R1142 Q2.n11 Q2.n10 6.86134
R1143 Q2.n7 Q2.n6 5.61236
R1144 Q2.n12 Q2.n9 5.01116
R1145 Q2.n17 Q2.n16 3.25085
R1146 Q2.n4 Q2.n3 3.00879
R1147 Q2.n7 Q2.n4 2.84996
R1148 Q2.n16 Q2.t1 2.2755
R1149 Q2.n16 Q2.n15 2.2755
R1150 Q2.n18 Q2.n13 2.25648
R1151 Q2.n9 Q2.n8 2.13398
R1152 Q2.n1 Q2.n0 1.80477
R1153 Q2.n4 Q2.n1 1.67937
R1154 Q2.n13 Q2.n12 1.52473
R1155 Q2.n13 Q2.n7 1.44626
R1156 Q2.n12 Q2.n11 1.12056
R1157 Q2.n1 Q2 0.105737
R1158 Q2.n18 Q2.n17 0.0919062
R1159 Q2.n3 Q2 0.0878146
R1160 Q2.n6 Q2 0.0878108
R1161 Q2.n11 Q2 0.0857632
R1162 Q2.n9 Q2 0.0810725
R1163 Q2 Q2.n18 0.073625
R1164 Q3.n1 Q3.t3 39.7867
R1165 Q3.n6 Q3.t5 36.935
R1166 Q3.n8 Q3.t8 31.528
R1167 Q3.n1 Q3.t7 30.2921
R1168 Q3.n6 Q3.t4 18.1962
R1169 Q3.n8 Q3.t6 15.3826
R1170 Q3.n15 Q3.n12 7.09905
R1171 Q3.n9 Q3.n8 6.86134
R1172 Q3.n10 Q3.n7 5.01116
R1173 Q3.n3 Q3.n0 4.5005
R1174 Q3.n2 Q3.n0 4.5005
R1175 Q3.n15 Q3.n14 3.25085
R1176 Q3.n14 Q3.t2 2.2755
R1177 Q3.n14 Q3.n13 2.2755
R1178 Q3.n16 Q3.n11 2.2505
R1179 Q3.n5 Q3.n4 2.2422
R1180 Q3.n7 Q3.n6 2.13398
R1181 Q3.n11 Q3.n5 1.73784
R1182 Q3.n11 Q3.n10 1.52239
R1183 Q3.n2 Q3.n1 1.38211
R1184 Q3.n10 Q3.n9 1.12056
R1185 Q3.n16 Q3.n15 0.0919062
R1186 Q3.n9 Q3 0.0857632
R1187 Q3.n7 Q3 0.0810725
R1188 Q3 Q3.n16 0.073625
R1189 Q3.n5 Q3.n0 0.025038
R1190 Q3.n4 Q3.n3 0.0239247
R1191 Q3.n3 Q3 0.0214589
R1192 Q3.n4 Q3.n2 0.00913014
C0 a_7956_1353# Q0 6.06e-21
C1 JK_FF_mag_3.nand3_mag_0.OUT Q2 0.00125f
C2 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C3 JK_FF_mag_0.nand2_mag_3.IN1 and2_mag_1.GF_INV_MAG_0.IN 0.00213f
C4 JK_FF_mag_3.nand3_mag_1.IN1 a_7574_2450# 2.36e-22
C5 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_2.J 0.0334f
C6 a_9510_2450# and2_mag_1.GF_INV_MAG_0.IN 0.069f
C7 a_634_1309# CLK 0.0101f
C8 a_3645_212# VDD 0.0123f
C9 JK_FF_mag_2.nand3_mag_0.OUT VDD 0.647f
C10 a_788_212# JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C11 a_7392_1353# RST 1.23e-20
C12 JK_FF_mag_3.Qb Q1 0.311f
C13 a_1352_212# a_1512_212# 0.0504f
C14 JK_FF_mag_2.J JK_FF_mag_0.J 0.0156f
C15 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_2.J 0.346f
C16 a_6662_212# Q2 0.00335f
C17 VDD a_4375_1353# 3.14e-19
C18 JK_FF_mag_0.nand3_mag_1.OUT a_9679_212# 1.17e-20
C19 a_10403_212# a_10563_212# 0.0504f
C20 JK_FF_mag_0.nand3_mag_0.OUT a_9845_1309# 0.0732f
C21 Q3 and2_mag_0.OUT 0.124f
C22 and2_mag_1.OUT Q2 0.0165f
C23 CLK VDD 1.09f
C24 a_11738_2752# nor_3_mag_0.IN3 2.44e-20
C25 JK_FF_mag_1.nand2_mag_3.IN1 RST 0.0675f
C26 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.Qb 0.28f
C27 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.Qb 0.0378f
C28 and2_mag_1.OUT Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C29 JK_FF_mag_1.nand2_mag_3.IN1 Q0 0.0228f
C30 JK_FF_mag_2.J and2_mag_1.GF_INV_MAG_0.IN 9.73e-19
C31 VDD a_3811_1309# 2.66e-19
C32 JK_FF_mag_2.Qb JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C33 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C34 JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.395f
C35 JK_FF_mag_3.nand2_mag_3.IN1 a_7956_1353# 0.011f
C36 JK_FF_mag_0.J a_9685_1309# 8.64e-19
C37 JK_FF_mag_0.nand3_mag_0.OUT a_9685_1309# 0.0203f
C38 and2_mag_0.GF_INV_MAG_0.IN Q1 0.0995f
C39 a_5503_1353# Q0 9.26e-19
C40 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_0.OUT 0.122f
C41 a_794_1309# JK_FF_mag_1.Qb 0.00392f
C42 JK_FF_mag_2.Qb a_4375_1353# 3.25e-19
C43 a_4939_1353# JK_FF_mag_2.nand3_mag_1.OUT 4.52e-20
C44 JK_FF_mag_3.nand3_mag_2.OUT Q1 0.235f
C45 a_794_1309# Q0 2.79e-20
C46 JK_FF_mag_3.nand3_mag_1.OUT RST 0.266f
C47 JK_FF_mag_3.Qb a_7546_212# 0.00696f
C48 JK_FF_mag_2.J Q1 0.0871f
C49 JK_FF_mag_2.nand3_mag_1.IN1 a_4375_1353# 0.0697f
C50 VDD a_3651_1309# 3.78e-19
C51 JK_FF_mag_3.nand3_mag_1.OUT Q0 0.00395f
C52 JK_FF_mag_3.nand2_mag_3.IN1 a_7392_1353# 1.43e-19
C53 JK_FF_mag_3.nand3_mag_0.OUT VDD 0.741f
C54 JK_FF_mag_0.nand2_mag_3.IN1 Q3 0.0263f
C55 JK_FF_mag_3.nand3_mag_1.IN1 and2_mag_0.GF_INV_MAG_0.IN 1.36e-19
C56 CLK a_1358_1353# 6.43e-21
C57 a_10403_212# Q2 3.6e-22
C58 JK_FF_mag_0.J RST 1.55e-19
C59 JK_FF_mag_3.Qb a_8520_1353# 0.0114f
C60 JK_FF_mag_0.nand3_mag_0.OUT RST 0.00229f
C61 JK_FF_mag_2.Qb a_3811_1309# 0.00392f
C62 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand3_mag_1.IN1 0.00157f
C63 JK_FF_mag_0.nand2_mag_4.IN2 Q3 0.0635f
C64 JK_FF_mag_0.J Q0 0.487f
C65 JK_FF_mag_0.nand3_mag_0.OUT Q0 0.27f
C66 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_2.J 0.0432f
C67 a_1512_212# JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C68 JK_FF_mag_3.nand2_mag_4.IN2 a_8520_1353# 4.52e-20
C69 JK_FF_mag_3.nand2_mag_3.IN1 a_6828_1309# 0.00119f
C70 a_6662_212# VDD 0.0132f
C71 a_4939_1353# VDD 3.14e-19
C72 a_628_212# JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C73 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand3_mag_1.OUT 0.159f
C74 a_11127_256# VDD 3.14e-19
C75 and2_mag_1.GF_INV_MAG_0.IN nor_3_mag_0.IN3 4.85e-20
C76 and2_mag_1.OUT VDD 0.576f
C77 JK_FF_mag_0.J and2_mag_2.GF_INV_MAG_0.IN 0.125f
C78 and2_mag_1.GF_INV_MAG_0.IN Q0 0.0979f
C79 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_2.Qb 2.81e-20
C80 JK_FF_mag_3.nand3_mag_2.OUT a_7546_212# 2.88e-20
C81 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN Q2 0.00311f
C82 a_1352_212# RST 8.64e-19
C83 JK_FF_mag_2.J Q3 2f
C84 a_1352_212# JK_FF_mag_1.Qb 0.00695f
C85 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_1.OUT 0.159f
C86 Q1 RST 0.133f
C87 a_1352_212# Q0 0.0102f
C88 a_3805_212# Q1 0.00789f
C89 Q3 a_9845_1309# 2.79e-20
C90 JK_FF_mag_2.J JK_FF_mag_1.nand3_mag_1.OUT 4.24e-20
C91 JK_FF_mag_2.J a_8520_1353# 7.4e-19
C92 Q0 Q1 1.16f
C93 a_9839_212# Q3 0.00789f
C94 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.00157f
C95 and2_mag_1.GF_INV_MAG_0.IN and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C96 a_5657_256# Q1 0.0157f
C97 a_4939_1353# JK_FF_mag_2.Qb 2.96e-19
C98 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_0.J 1.41e-20
C99 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.J 0.00488f
C100 JK_FF_mag_1.nand3_mag_0.OUT CLK 0.267f
C101 JK_FF_mag_2.nand2_mag_3.IN1 VDD 1.03f
C102 a_4939_1353# JK_FF_mag_2.nand3_mag_1.IN1 0.0059f
C103 JK_FF_mag_3.nand3_mag_1.IN1 RST 0.177f
C104 CLK JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C105 a_6822_212# JK_FF_mag_3.nand3_mag_1.OUT 1.5e-20
C106 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C107 JK_FF_mag_3.nand3_mag_1.IN1 Q0 0.0126f
C108 and2_mag_2.GF_INV_MAG_0.IN Q1 0.303f
C109 a_10403_212# VDD 2.21e-19
C110 JK_FF_mag_2.nand3_mag_2.OUT Q1 0.338f
C111 a_4369_212# RST 0.00169f
C112 a_788_212# JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C113 Q0 a_4369_212# 3.6e-22
C114 JK_FF_mag_0.nand3_mag_1.OUT and2_mag_1.OUT 0.00243f
C115 JK_FF_mag_0.nand3_mag_1.OUT a_11127_256# 0.00378f
C116 a_7546_212# RST 0.00186f
C117 Q3 RST 0.0395f
C118 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.Qb 0.28f
C119 JK_FF_mag_3.nand2_mag_3.IN1 Q1 0.447f
C120 Q3 nor_3_mag_0.IN3 0.00442f
C121 Q2 VDD 2.85f
C122 Q0 Q3 0.149f
C123 JK_FF_mag_1.nand3_mag_1.OUT RST 0.261f
C124 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand3_mag_1.IN1 0.231f
C125 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.Qb 0.25f
C126 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD 0.51f
C127 JK_FF_mag_2.nand3_mag_2.OUT a_4369_212# 9.1e-19
C128 Q0 a_8520_1353# 9.45e-19
C129 JK_FF_mag_1.nand3_mag_1.OUT Q0 0.0343f
C130 JK_FF_mag_0.nand3_mag_1.OUT a_10563_212# 0.0733f
C131 JK_FF_mag_2.nand2_mag_1.IN2 RST 9.24e-20
C132 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_1.IN1 0.231f
C133 JK_FF_mag_2.nand2_mag_1.IN2 Q0 0.0205f
C134 a_6822_212# Q1 0.00166f
C135 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C136 a_7956_1353# JK_FF_mag_3.nand3_mag_1.OUT 4.52e-20
C137 JK_FF_mag_0.nand3_mag_1.OUT a_10403_212# 0.0203f
C138 JK_FF_mag_2.nand3_mag_1.OUT VDD 0.999f
C139 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.J 0.00586f
C140 a_6668_1309# a_6828_1309# 0.0504f
C141 a_634_1309# VDD 0.00752f
C142 a_2486_1353# RST 6.14e-19
C143 JK_FF_mag_1.Qb a_2486_1353# 0.0114f
C144 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.J 8.2e-19
C145 a_5093_256# RST 9.41e-19
C146 Q0 a_2486_1353# 0.069f
C147 a_7392_1353# JK_FF_mag_3.nand3_mag_1.OUT 0.0202f
C148 a_9679_212# a_9839_212# 0.0504f
C149 JK_FF_mag_0.nand3_mag_1.OUT Q2 2.45e-22
C150 JK_FF_mag_3.nand2_mag_3.IN1 a_8520_1353# 0.00118f
C151 a_10409_1353# and2_mag_1.OUT 5.94e-20
C152 a_1922_1353# RST 6.14e-19
C153 JK_FF_mag_1.Qb a_1922_1353# 2.96e-19
C154 JK_FF_mag_0.nand3_mag_1.IN1 and2_mag_1.OUT 4.42e-19
C155 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.Qb 0.25f
C156 JK_FF_mag_0.nand3_mag_1.OUT Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.25e-20
C157 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_2.J 0.11f
C158 a_794_1309# JK_FF_mag_1.nand2_mag_3.IN1 0.00119f
C159 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_1.IN2 2.11e-19
C160 Q0 a_1922_1353# 6.06e-21
C161 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C162 a_9839_212# JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C163 Q2 a_7386_212# 0.0102f
C164 a_10563_212# JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C165 a_3645_212# JK_FF_mag_2.J 2.81e-19
C166 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.J 0.1f
C167 JK_FF_mag_2.nand2_mag_4.IN2 RST 0.0172f
C168 JK_FF_mag_1.nand2_mag_1.IN2 RST 0.00434f
C169 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.Qb 0.0592f
C170 a_11691_256# Q3 0.0157f
C171 and2_mag_1.OUT and2_mag_0.OUT 0.0693f
C172 JK_FF_mag_2.nand2_mag_4.IN2 Q0 6.82e-19
C173 a_9679_212# RST 0.00186f
C174 JK_FF_mag_2.Qb VDD 0.912f
C175 a_628_212# a_788_212# 0.0504f
C176 JK_FF_mag_2.J a_4375_1353# 3.12e-19
C177 JK_FF_mag_1.nand2_mag_1.IN2 Q0 0.108f
C178 JK_FF_mag_2.nand2_mag_4.IN2 a_5657_256# 0.00372f
C179 JK_FF_mag_3.Qb JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C180 JK_FF_mag_3.nand2_mag_1.IN2 Q2 0.113f
C181 a_9679_212# Q0 0.00117f
C182 a_7392_1353# Q1 1.25e-20
C183 a_7956_1353# JK_FF_mag_3.nand3_mag_1.IN1 0.0059f
C184 JK_FF_mag_2.nand3_mag_1.IN1 VDD 0.652f
C185 VDD a_1358_1353# 3.14e-19
C186 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT 0.768f
C187 JK_FF_mag_1.nand2_mag_4.IN2 a_2640_256# 0.00372f
C188 a_10973_1353# Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 5.94e-20
C189 a_6668_1309# Q1 0.0101f
C190 JK_FF_mag_0.nand3_mag_2.OUT RST 0.0759f
C191 a_2076_256# RST 9.41e-19
C192 JK_FF_mag_2.J a_3811_1309# 9.32e-19
C193 a_2076_256# JK_FF_mag_1.Qb 0.00964f
C194 JK_FF_mag_0.nand3_mag_2.OUT Q0 0.235f
C195 JK_FF_mag_0.nand3_mag_1.OUT VDD 0.994f
C196 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_2.J 1.54e-19
C197 a_628_212# Q0 0.00335f
C198 a_2076_256# Q0 0.00859f
C199 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.J 0.106f
C200 a_6828_1309# Q1 0.00939f
C201 a_7392_1353# JK_FF_mag_3.nand3_mag_1.IN1 0.0697f
C202 JK_FF_mag_0.nand2_mag_1.IN2 Q3 0.11f
C203 a_11578_2752# Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 9.16e-20
C204 Vdiv10 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.82e-19
C205 a_5503_1353# Q1 0.069f
C206 JK_FF_mag_0.nand2_mag_3.IN1 and2_mag_1.OUT 0.00718f
C207 JK_FF_mag_0.nand3_mag_1.IN1 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.29e-19
C208 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.Qb 0.0378f
C209 a_11127_256# JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C210 a_9510_2450# and2_mag_1.OUT 3.92e-20
C211 JK_FF_mag_2.J a_3651_1309# 0.00876f
C212 a_788_212# CLK 0.00164f
C213 a_3645_212# RST 0.00186f
C214 a_634_1309# JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C215 JK_FF_mag_2.nand3_mag_0.OUT RST 3.84e-20
C216 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_1.Qb 2.81e-20
C217 a_3645_212# a_3805_212# 0.0504f
C218 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C219 a_8542_2450# Q2 0.0112f
C220 and2_mag_1.GF_INV_MAG_0.IN JK_FF_mag_0.J 0.0275f
C221 VDD a_7386_212# 0.00123f
C222 JK_FF_mag_0.nand3_mag_0.OUT and2_mag_1.GF_INV_MAG_0.IN 1.98e-19
C223 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_2.J 0.00602f
C224 a_3645_212# Q0 0.001f
C225 Q2 a_8110_256# 0.00859f
C226 JK_FF_mag_2.nand3_mag_0.OUT Q0 0.298f
C227 JK_FF_mag_0.nand2_mag_4.IN2 a_11127_256# 0.069f
C228 JK_FF_mag_3.nand3_mag_1.OUT Q1 0.00335f
C229 a_4375_1353# RST 1.23e-20
C230 a_11537_1353# VDD 3.56e-19
C231 Q0 a_4375_1353# 6.43e-21
C232 CLK JK_FF_mag_1.Qb 0.307f
C233 CLK RST 5.44e-19
C234 JK_FF_mag_3.nand3_mag_2.OUT a_6662_212# 0.0202f
C235 Q2 and2_mag_0.OUT 0.179f
C236 JK_FF_mag_0.J Q1 0.0685f
C237 JK_FF_mag_1.nand3_mag_1.IN1 a_1922_1353# 0.0059f
C238 a_7574_2450# Q2 0.00929f
C239 JK_FF_mag_1.nand3_mag_0.OUT VDD 0.741f
C240 a_11738_2752# Q3 0.019f
C241 JK_FF_mag_2.nand3_mag_1.OUT a_4529_212# 0.0733f
C242 CLK Q0 0.149f
C243 a_4939_1353# JK_FF_mag_2.J 7.4e-19
C244 JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.397f
C245 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C246 JK_FF_mag_2.nand3_mag_2.OUT a_3645_212# 0.0202f
C247 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN and2_mag_0.OUT 0.0654f
C248 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C249 VDD JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C250 a_10973_1353# VDD 3.14e-19
C251 JK_FF_mag_1.Qb a_3811_1309# 1.41e-20
C252 a_11127_256# JK_FF_mag_2.J 0.00964f
C253 JK_FF_mag_1.nand2_mag_4.IN2 RST 0.019f
C254 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.Qb 0.198f
C255 Q0 a_3811_1309# 0.00939f
C256 JK_FF_mag_1.nand2_mag_4.IN2 Q0 0.0635f
C257 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_1.OUT 0.16f
C258 a_8674_256# Q2 0.0157f
C259 and2_mag_1.GF_INV_MAG_0.IN Q1 1.17e-19
C260 a_11578_2752# VDD 0.234f
C261 Vdiv10 VDD 0.0712f
C262 JK_FF_mag_1.Qb a_3651_1309# 1.86e-20
C263 a_10409_1353# VDD 3.14e-19
C264 JK_FF_mag_3.nand3_mag_1.OUT a_7546_212# 0.0733f
C265 a_10563_212# JK_FF_mag_2.J 0.00696f
C266 JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.652f
C267 JK_FF_mag_3.Qb Q2 1.96f
C268 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C269 JK_FF_mag_3.nand3_mag_0.OUT RST 3.84e-20
C270 Q0 a_3651_1309# 0.0101f
C271 VDD a_4529_212# 0.00101f
C272 a_5503_1353# JK_FF_mag_2.nand2_mag_1.IN2 0.00372f
C273 JK_FF_mag_3.nand3_mag_0.OUT Q0 0.0285f
C274 JK_FF_mag_0.nand2_mag_3.IN1 Q2 0.0569f
C275 JK_FF_mag_1.nand3_mag_0.OUT a_1358_1353# 0.00378f
C276 a_9510_2450# Q2 0.0096f
C277 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.J 0.0905f
C278 JK_FF_mag_3.nand2_mag_4.IN2 Q2 0.0635f
C279 a_8542_2450# VDD 3.14e-19
C280 JK_FF_mag_0.nand2_mag_3.IN1 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00943f
C281 JK_FF_mag_0.nand3_mag_0.OUT Q3 8.98e-19
C282 VDD a_8110_256# 0.00152f
C283 a_10403_212# JK_FF_mag_2.J 0.00695f
C284 a_6662_212# RST 0.00186f
C285 JK_FF_mag_1.nand2_mag_3.IN1 a_2486_1353# 0.00118f
C286 JK_FF_mag_3.nand3_mag_1.IN1 Q1 0.00152f
C287 and2_mag_1.OUT RST 4.25e-20
C288 JK_FF_mag_0.nand3_mag_1.OUT a_10973_1353# 4.52e-20
C289 and2_mag_0.OUT VDD 0.911f
C290 a_7574_2450# VDD 6e-19
C291 and2_mag_0.GF_INV_MAG_0.IN Q2 0.322f
C292 JK_FF_mag_2.Qb a_4529_212# 0.00696f
C293 and2_mag_1.OUT Q0 2.11e-20
C294 Q1 a_4369_212# 0.0102f
C295 JK_FF_mag_3.nand3_mag_2.OUT Q2 0.338f
C296 JK_FF_mag_1.nand2_mag_3.IN1 a_1922_1353# 0.011f
C297 JK_FF_mag_2.nand3_mag_1.IN1 a_4529_212# 8.64e-19
C298 JK_FF_mag_2.J Q2 0.0626f
C299 a_10563_212# RST 0.00127f
C300 JK_FF_mag_0.nand3_mag_1.OUT a_10409_1353# 0.0202f
C301 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_0.OUT 0.0854f
C302 a_8674_256# VDD 0.00152f
C303 a_9839_212# Q2 1.86e-20
C304 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C305 a_1352_212# JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C306 JK_FF_mag_2.nand2_mag_3.IN1 RST 0.0568f
C307 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_1.Qb 7.08e-20
C308 a_3805_212# JK_FF_mag_2.nand2_mag_3.IN1 1.46e-19
C309 JK_FF_mag_1.nand3_mag_1.IN1 CLK 9.71e-20
C310 JK_FF_mag_3.Qb VDD 0.911f
C311 JK_FF_mag_2.nand2_mag_3.IN1 Q0 1.3f
C312 Q2 a_9685_1309# 6.36e-19
C313 JK_FF_mag_3.nand3_mag_1.IN1 a_7546_212# 8.64e-19
C314 a_10403_212# RST 0.00169f
C315 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C316 JK_FF_mag_2.nand2_mag_1.IN2 Q1 0.108f
C317 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_3.IN1 0.36f
C318 JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.14f
C319 a_1512_212# VDD 0.00101f
C320 a_9510_2450# VDD 3.14e-19
C321 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.J 0.0334f
C322 JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.395f
C323 a_5503_1353# JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C324 JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C325 JK_FF_mag_0.nand3_mag_1.OUT and2_mag_0.OUT 3.38e-19
C326 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C327 Q2 RST 0.105f
C328 a_2640_256# VDD 0.00152f
C329 a_6662_212# a_6822_212# 0.0504f
C330 JK_FF_mag_3.Qb JK_FF_mag_2.Qb 2.59e-21
C331 a_2076_256# JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C332 and2_mag_0.GF_INV_MAG_0.IN VDD 0.455f
C333 Q2 nor_3_mag_0.IN3 3.87e-19
C334 Q0 Q2 0.622f
C335 Q1 a_5093_256# 0.00859f
C336 a_10973_1353# JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C337 JK_FF_mag_3.nand3_mag_2.OUT VDD 0.768f
C338 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN nor_3_mag_0.IN3 0.11f
C339 JK_FF_mag_2.J VDD 1.65f
C340 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.00233f
C341 a_11537_1353# and2_mag_0.OUT 1.54e-19
C342 Vdiv10 a_11578_2752# 0.0132f
C343 a_9839_212# VDD 0.00299f
C344 and2_mag_2.GF_INV_MAG_0.IN Q2 0.103f
C345 a_10409_1353# JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C346 JK_FF_mag_2.nand3_mag_1.OUT RST 0.266f
C347 a_3805_212# JK_FF_mag_2.nand3_mag_1.OUT 1.5e-20
C348 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C349 JK_FF_mag_2.nand3_mag_1.OUT Q0 0.00481f
C350 VDD a_9685_1309# 2.21e-19
C351 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C352 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C353 JK_FF_mag_1.nand2_mag_3.IN1 CLK 0.407f
C354 a_788_212# VDD 0.00892f
C355 JK_FF_mag_2.Qb JK_FF_mag_2.J 0.0838f
C356 JK_FF_mag_3.Qb a_7386_212# 0.00695f
C357 JK_FF_mag_3.nand2_mag_3.IN1 Q2 0.0209f
C358 JK_FF_mag_2.nand2_mag_4.IN2 Q1 0.0635f
C359 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.J 0.0432f
C360 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 0.321f
C361 a_11578_2752# and2_mag_0.OUT 0.0294f
C362 Vdiv10 and2_mag_0.OUT 0.119f
C363 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C364 a_794_1309# CLK 0.00939f
C365 a_7392_1353# JK_FF_mag_3.nand3_mag_0.OUT 0.00378f
C366 a_11537_1353# JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C367 VDD RST 1.15f
C368 JK_FF_mag_0.nand3_mag_1.IN1 and2_mag_0.OUT 6.69e-19
C369 JK_FF_mag_1.Qb VDD 0.916f
C370 a_3805_212# VDD 0.00863f
C371 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_2.J 0.251f
C372 nor_3_mag_0.IN3 VDD 0.395f
C373 JK_FF_mag_0.nand2_mag_4.IN2 a_11537_1353# 4.52e-20
C374 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.Qb 0.0591f
C375 Q0 VDD 4.98f
C376 a_6668_1309# JK_FF_mag_3.nand3_mag_0.OUT 0.0203f
C377 a_5657_256# VDD 0.00152f
C378 a_6822_212# Q2 0.00789f
C379 a_8542_2450# and2_mag_0.OUT 0.00138f
C380 JK_FF_mag_0.nand3_mag_1.OUT a_9839_212# 1.5e-20
C381 JK_FF_mag_1.nand3_mag_1.OUT a_1922_1353# 4.52e-20
C382 a_1512_212# JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C383 a_6828_1309# JK_FF_mag_3.nand3_mag_0.OUT 0.0732f
C384 a_10973_1353# JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C385 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C386 JK_FF_mag_3.nand3_mag_2.OUT a_7386_212# 9.1e-19
C387 and2_mag_2.GF_INV_MAG_0.IN VDD 0.43f
C388 JK_FF_mag_2.nand3_mag_2.OUT VDD 0.748f
C389 JK_FF_mag_2.Qb RST 0.179f
C390 JK_FF_mag_2.Qb JK_FF_mag_1.Qb 2.59e-21
C391 a_11537_1353# JK_FF_mag_2.J 0.0114f
C392 JK_FF_mag_2.nand3_mag_0.OUT Q1 7.24e-19
C393 a_3645_212# Q1 0.00335f
C394 a_10409_1353# JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C395 JK_FF_mag_2.Qb Q0 0.348f
C396 a_9679_212# Q3 0.00335f
C397 JK_FF_mag_2.nand3_mag_1.IN1 RST 0.177f
C398 JK_FF_mag_3.nand2_mag_1.IN2 and2_mag_0.GF_INV_MAG_0.IN 6.88e-21
C399 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C400 JK_FF_mag_1.Qb a_1358_1353# 3.33e-19
C401 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C402 a_5657_256# JK_FF_mag_2.Qb 0.0811f
C403 JK_FF_mag_0.nand2_mag_4.IN2 Vdiv10 3.1e-22
C404 JK_FF_mag_2.nand3_mag_1.IN1 Q0 0.0129f
C405 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C406 JK_FF_mag_3.Qb a_8542_2450# 1.45e-20
C407 JK_FF_mag_3.Qb a_8110_256# 0.00964f
C408 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_2.J 0.00488f
C409 JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.07f
C410 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C411 a_10973_1353# JK_FF_mag_2.J 2.96e-19
C412 JK_FF_mag_0.nand3_mag_1.OUT RST 0.255f
C413 a_6662_212# JK_FF_mag_3.nand3_mag_1.OUT 1.17e-20
C414 JK_FF_mag_0.nand3_mag_2.OUT Q3 0.338f
C415 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.Qb 0.103f
C416 JK_FF_mag_3.nand2_mag_4.IN2 a_8542_2450# 1.29e-22
C417 JK_FF_mag_0.nand3_mag_1.OUT Q0 9.9e-19
C418 JK_FF_mag_3.nand2_mag_4.IN2 a_8110_256# 0.069f
C419 JK_FF_mag_3.Qb and2_mag_0.OUT 1.33e-20
C420 Q1 a_3811_1309# 2.79e-20
C421 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_1.IN1 0.00157f
C422 a_628_212# JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C423 a_2076_256# JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C424 JK_FF_mag_2.J a_11578_2752# 9.21e-20
C425 JK_FF_mag_2.J Vdiv10 4.19e-19
C426 JK_FF_mag_0.nand2_mag_3.IN1 and2_mag_0.OUT 0.065f
C427 a_10409_1353# JK_FF_mag_2.J 3.25e-19
C428 a_9510_2450# and2_mag_0.OUT 0.00138f
C429 JK_FF_mag_0.nand2_mag_1.IN2 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.42e-19
C430 a_6822_212# VDD 0.00891f
C431 a_7386_212# RST 0.00169f
C432 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_2.J 0.038f
C433 a_788_212# JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C434 JK_FF_mag_1.nand2_mag_1.IN2 a_2486_1353# 0.00372f
C435 and2_mag_1.OUT JK_FF_mag_0.J 2.57e-20
C436 a_8542_2450# and2_mag_0.GF_INV_MAG_0.IN 5.1e-20
C437 JK_FF_mag_0.nand3_mag_0.OUT and2_mag_1.OUT 1.29e-19
C438 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.Qb 3.49e-19
C439 JK_FF_mag_2.nand2_mag_4.IN2 a_5093_256# 0.069f
C440 a_8674_256# JK_FF_mag_3.Qb 0.0811f
C441 a_5503_1353# JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C442 a_11537_1353# nor_3_mag_0.IN3 2.1e-20
C443 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.nand3_mag_1.IN1 1.54e-21
C444 JK_FF_mag_3.nand3_mag_0.OUT Q1 0.273f
C445 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.Qb 0.343f
C446 a_8674_256# JK_FF_mag_3.nand2_mag_4.IN2 0.00372f
C447 JK_FF_mag_3.nand2_mag_1.IN2 RST 9.24e-20
C448 and2_mag_0.GF_INV_MAG_0.IN and2_mag_0.OUT 0.125f
C449 a_11691_256# VDD 3.14e-19
C450 JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.652f
C451 a_7574_2450# and2_mag_0.GF_INV_MAG_0.IN 0.069f
C452 and2_mag_1.OUT and2_mag_1.GF_INV_MAG_0.IN 0.124f
C453 JK_FF_mag_1.nand2_mag_1.IN2 a_1922_1353# 0.069f
C454 JK_FF_mag_1.nand3_mag_0.OUT Q0 7.24e-19
C455 JK_FF_mag_1.nand3_mag_2.OUT RST 0.0495f
C456 JK_FF_mag_1.Qb JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C457 JK_FF_mag_3.nand2_mag_1.IN2 Q0 0.0215f
C458 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_3.Qb 7.08e-20
C459 Q0 JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C460 JK_FF_mag_2.J and2_mag_0.OUT 0.00656f
C461 a_11738_2752# Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 5.39e-20
C462 a_6828_1309# Q2 2.79e-20
C463 a_6662_212# Q1 0.00119f
C464 JK_FF_mag_1.nand3_mag_1.OUT CLK 6.64e-19
C465 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.Qb 0.198f
C466 a_4939_1353# Q1 6.06e-21
C467 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_0.OUT 0.122f
C468 and2_mag_1.OUT Q1 8.51e-22
C469 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C470 a_10409_1353# RST 2.78e-19
C471 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C472 Vdiv10 nor_3_mag_0.IN3 0.0263f
C473 a_11578_2752# nor_3_mag_0.IN3 9.02e-19
C474 JK_FF_mag_0.nand3_mag_1.IN1 RST 0.152f
C475 a_10409_1353# Q0 6.43e-21
C476 a_4529_212# RST 0.00186f
C477 JK_FF_mag_3.nand3_mag_1.OUT Q2 0.0352f
C478 JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C479 JK_FF_mag_0.nand3_mag_1.IN1 Q0 5.11e-19
C480 a_7956_1353# VDD 3.14e-19
C481 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.Qb 0.103f
C482 JK_FF_mag_1.nand3_mag_1.IN1 a_1358_1353# 0.0697f
C483 JK_FF_mag_3.Qb JK_FF_mag_2.J 0.0835f
C484 a_8110_256# RST 9.41e-19
C485 JK_FF_mag_0.J Q2 0.289f
C486 JK_FF_mag_3.Qb a_9845_1309# 1.41e-20
C487 JK_FF_mag_0.nand3_mag_0.OUT Q2 8.27e-19
C488 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_2.J 0.283f
C489 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C490 JK_FF_mag_2.nand2_mag_3.IN1 Q1 0.018f
C491 JK_FF_mag_0.nand2_mag_3.IN1 a_9845_1309# 0.00119f
C492 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_2.J 0.00586f
C493 a_7392_1353# VDD 3.14e-19
C494 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_2.J 0.199f
C495 a_9679_212# JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C496 a_9839_212# JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C497 JK_FF_mag_2.nand3_mag_2.OUT a_4529_212# 2.88e-20
C498 JK_FF_mag_1.nand2_mag_4.IN2 a_2486_1353# 4.52e-20
C499 a_6668_1309# VDD 0.00746f
C500 nor_3_mag_0.IN3 and2_mag_0.OUT 0.144f
C501 Q0 and2_mag_0.OUT 0.026f
C502 and2_mag_1.OUT Q3 0.00132f
C503 a_11738_2752# VDD 0.0407f
C504 and2_mag_1.GF_INV_MAG_0.IN Q2 0.305f
C505 a_11127_256# Q3 0.00859f
C506 a_634_1309# a_794_1309# 0.0504f
C507 a_8542_2450# and2_mag_2.GF_INV_MAG_0.IN 0.069f
C508 JK_FF_mag_3.Qb a_9685_1309# 1.86e-20
C509 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN and2_mag_1.GF_INV_MAG_0.IN 3.38e-19
C510 JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.18f
C511 a_6828_1309# VDD 2.66e-19
C512 a_4939_1353# JK_FF_mag_2.nand2_mag_1.IN2 0.069f
C513 a_8674_256# RST 9.66e-19
C514 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_2.J 0.0151f
C515 a_5503_1353# VDD 3.56e-19
C516 and2_mag_2.GF_INV_MAG_0.IN and2_mag_0.OUT 0.0758f
C517 Q2 Q1 0.98f
C518 a_10563_212# Q3 0.0101f
C519 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C520 JK_FF_mag_2.J a_9845_1309# 0.00486f
C521 a_794_1309# VDD 2.66e-19
C522 JK_FF_mag_3.Qb RST 0.179f
C523 JK_FF_mag_3.nand2_mag_3.IN1 a_8110_256# 0.0036f
C524 a_6668_1309# JK_FF_mag_2.Qb 1.86e-20
C525 JK_FF_mag_3.nand3_mag_1.OUT VDD 0.999f
C526 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C527 JK_FF_mag_1.nand2_mag_1.IN2 CLK 1.48e-20
C528 JK_FF_mag_3.Qb Q0 0.0615f
C529 JK_FF_mag_0.nand2_mag_3.IN1 RST 0.00237f
C530 a_1512_212# RST 0.00186f
C531 a_1512_212# JK_FF_mag_1.Qb 0.00696f
C532 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C533 a_6828_1309# JK_FF_mag_2.Qb 1.41e-20
C534 JK_FF_mag_0.nand2_mag_3.IN1 nor_3_mag_0.IN3 4.39e-19
C535 JK_FF_mag_3.nand3_mag_1.IN1 Q2 0.00545f
C536 a_10403_212# Q3 0.0102f
C537 JK_FF_mag_3.nand2_mag_4.IN2 RST 0.0172f
C538 JK_FF_mag_0.nand2_mag_3.IN1 Q0 0.529f
C539 a_1512_212# Q0 0.0101f
C540 a_9510_2450# Q0 0.01f
C541 JK_FF_mag_0.nand2_mag_4.IN2 RST 2.96e-19
C542 JK_FF_mag_3.nand2_mag_3.IN1 and2_mag_0.OUT 6.22e-20
C543 JK_FF_mag_2.J a_9685_1309# 0.00111f
C544 JK_FF_mag_3.nand2_mag_4.IN2 Q0 6.82e-19
C545 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C546 JK_FF_mag_0.J VDD 0.496f
C547 JK_FF_mag_0.nand3_mag_0.OUT VDD 0.648f
C548 JK_FF_mag_1.nand2_mag_3.IN1 a_1358_1353# 1.43e-19
C549 a_11537_1353# JK_FF_mag_0.nand2_mag_1.IN2 0.00372f
C550 a_5503_1353# JK_FF_mag_2.Qb 0.0114f
C551 JK_FF_mag_2.nand3_mag_1.OUT Q1 0.0343f
C552 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C553 a_9685_1309# a_9845_1309# 0.0504f
C554 JK_FF_mag_3.Qb and2_mag_2.GF_INV_MAG_0.IN 1e-19
C555 a_2640_256# RST 9.66e-19
C556 a_628_212# CLK 0.00117f
C557 a_2640_256# JK_FF_mag_1.Qb 0.0811f
C558 a_9510_2450# and2_mag_2.GF_INV_MAG_0.IN 5.1e-20
C559 Q2 a_7546_212# 0.0101f
C560 a_2640_256# Q0 0.0157f
C561 and2_mag_1.GF_INV_MAG_0.IN VDD 0.44f
C562 Q2 Q3 9.83e-19
C563 and2_mag_0.GF_INV_MAG_0.IN Q0 4.36e-20
C564 JK_FF_mag_3.nand3_mag_2.OUT RST 0.0758f
C565 JK_FF_mag_3.nand2_mag_1.IN2 a_7956_1353# 0.069f
C566 JK_FF_mag_2.nand3_mag_0.OUT a_4375_1353# 0.00378f
C567 a_10973_1353# JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C568 JK_FF_mag_2.J RST 3.04f
C569 JK_FF_mag_2.J JK_FF_mag_1.Qb 9.14e-19
C570 JK_FF_mag_1.nand2_mag_4.IN2 a_2076_256# 0.069f
C571 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN Q3 0.00357f
C572 JK_FF_mag_2.J Q0 0.783f
C573 Q2 a_8520_1353# 0.069f
C574 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.Qb 0.28f
C575 a_1352_212# VDD 0.00123f
C576 a_9839_212# RST 0.00186f
C577 JK_FF_mag_2.nand3_mag_1.OUT a_4369_212# 0.0203f
C578 Q0 a_9845_1309# 0.00939f
C579 JK_FF_mag_2.nand2_mag_3.IN1 a_5093_256# 0.0036f
C580 Q1 VDD 4.07f
C581 a_9839_212# Q0 0.00164f
C582 and2_mag_0.GF_INV_MAG_0.IN and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C583 JK_FF_mag_2.nand3_mag_0.OUT a_3811_1309# 0.0732f
C584 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C585 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C586 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.J 0.0286f
C587 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.J 0.00174f
C588 Q0 a_9685_1309# 0.0101f
C589 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C590 JK_FF_mag_3.nand3_mag_1.IN1 VDD 0.652f
C591 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_0.OUT 0.0894f
C592 a_788_212# Q0 0.00789f
C593 JK_FF_mag_3.nand3_mag_1.OUT a_7386_212# 0.0203f
C594 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C595 JK_FF_mag_2.nand3_mag_0.OUT a_3651_1309# 0.0203f
C596 JK_FF_mag_3.nand2_mag_3.IN1 and2_mag_0.GF_INV_MAG_0.IN 0.00137f
C597 JK_FF_mag_2.Qb Q1 1.96f
C598 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand3_mag_1.OUT 0.00975f
C599 VDD a_4369_212# 0.00123f
C600 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C601 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.J 0.0501f
C602 a_794_1309# JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C603 a_11738_2752# Vdiv10 0.198f
C604 a_11738_2752# a_11578_2752# 0.186f
C605 JK_FF_mag_1.Qb RST 0.144f
C606 a_3805_212# RST 0.00186f
C607 JK_FF_mag_2.nand3_mag_1.IN1 Q1 0.00335f
C608 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C609 JK_FF_mag_0.nand2_mag_1.IN2 and2_mag_0.OUT 0.00178f
C610 Q0 RST 0.154f
C611 JK_FF_mag_1.Qb Q0 1.96f
C612 VDD a_7546_212# 0.00101f
C613 a_3805_212# Q0 0.00166f
C614 Q3 VDD 1.18f
C615 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand3_mag_1.OUT 0.00975f
C616 a_5657_256# RST 9.66e-19
C617 a_1512_212# JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C618 a_3651_1309# a_3811_1309# 0.0504f
C619 JK_FF_mag_0.nand3_mag_2.OUT a_10563_212# 2.88e-20
C620 JK_FF_mag_1.nand3_mag_1.OUT VDD 0.999f
C621 JK_FF_mag_0.nand2_mag_4.IN2 a_11691_256# 0.00372f
C622 VDD a_8520_1353# 3.56e-19
C623 JK_FF_mag_3.nand3_mag_2.OUT a_6822_212# 0.0731f
C624 JK_FF_mag_2.Qb a_4369_212# 0.00695f
C625 JK_FF_mag_2.nand3_mag_1.OUT a_5093_256# 0.00378f
C626 JK_FF_mag_2.nand3_mag_2.OUT RST 0.0763f
C627 JK_FF_mag_2.nand2_mag_1.IN2 VDD 0.397f
C628 JK_FF_mag_2.nand3_mag_2.OUT a_3805_212# 0.0731f
C629 and2_mag_2.GF_INV_MAG_0.IN Q0 0.0116f
C630 JK_FF_mag_2.nand3_mag_2.OUT Q0 0.233f
C631 JK_FF_mag_0.nand3_mag_2.OUT a_10403_212# 9.1e-19
C632 a_11738_2752# and2_mag_0.OUT 0.00894f
C633 Q1 a_7386_212# 3.6e-22
C634 a_7956_1353# JK_FF_mag_3.Qb 2.96e-19
C635 a_9679_212# Q2 2.55e-20
C636 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C637 a_11691_256# JK_FF_mag_2.J 0.0811f
C638 JK_FF_mag_0.nand3_mag_0.OUT a_10409_1353# 0.00378f
C639 JK_FF_mag_3.nand2_mag_3.IN1 RST 0.055f
C640 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.J 0.00264f
C641 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C642 JK_FF_mag_3.nand3_mag_1.OUT a_8110_256# 0.00378f
C643 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C644 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand3_mag_0.OUT 0.0854f
C645 VDD a_2486_1353# 3.56e-19
C646 JK_FF_mag_3.nand2_mag_3.IN1 Q0 0.857f
C647 JK_FF_mag_1.nand3_mag_1.OUT a_1358_1353# 0.0202f
C648 a_7392_1353# JK_FF_mag_3.Qb 3.25e-19
C649 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.Qb 0.0591f
C650 a_1352_212# JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C651 VDD a_5093_256# 0.00152f
C652 JK_FF_mag_3.nand2_mag_1.IN2 Q1 5.37e-19
C653 JK_FF_mag_2.nand2_mag_3.IN1 a_4375_1353# 1.43e-19
C654 JK_FF_mag_0.nand3_mag_2.OUT Q2 9.98e-19
C655 JK_FF_mag_0.nand3_mag_1.OUT Q3 0.0345f
C656 a_11578_2752# and2_mag_1.GF_INV_MAG_0.IN 2.85e-20
C657 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand3_mag_1.IN1 0.109f
C658 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand3_mag_1.OUT 0.122f
C659 JK_FF_mag_3.nand3_mag_1.OUT a_7574_2450# 3.38e-20
C660 VDD a_1922_1353# 3.14e-19
C661 a_6822_212# RST 0.00186f
C662 a_6828_1309# JK_FF_mag_3.Qb 0.00392f
C663 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_2.J 0.0592f
C664 JK_FF_mag_2.nand2_mag_3.IN1 a_3811_1309# 0.00119f
C665 a_7386_212# a_7546_212# 0.0504f
C666 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand3_mag_1.IN1 0.109f
C667 JK_FF_mag_0.J and2_mag_0.OUT 0.0659f
C668 a_7956_1353# JK_FF_mag_2.J 7.4e-19
C669 JK_FF_mag_0.nand3_mag_0.OUT and2_mag_0.OUT 8.94e-19
C670 JK_FF_mag_2.Qb a_5093_256# 0.00964f
C671 a_11537_1353# Q3 0.069f
C672 Q1 a_4529_212# 0.0101f
C673 JK_FF_mag_1.nand3_mag_1.IN1 RST 0.189f
C674 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.Qb 0.0384f
C675 JK_FF_mag_2.nand2_mag_4.IN2 VDD 0.395f
C676 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.Qb 0.25f
C677 a_7392_1353# JK_FF_mag_2.J 3.12e-19
C678 and2_mag_1.GF_INV_MAG_0.IN and2_mag_0.OUT 0.0496f
C679 a_8542_2450# Q1 0.0084f
C680 JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.397f
C681 JK_FF_mag_1.nand3_mag_1.IN1 Q0 0.00356f
C682 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_2.nand2_mag_3.IN1 4.27e-20
C683 a_9679_212# VDD 0.00727f
C684 a_6668_1309# JK_FF_mag_2.J 0.00111f
C685 JK_FF_mag_2.J a_11738_2752# 3.02e-19
C686 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C687 JK_FF_mag_3.Qb JK_FF_mag_0.J 5.7e-19
C688 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand3_mag_1.OUT 0.122f
C689 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_3.Qb 2.81e-20
C690 a_3645_212# JK_FF_mag_2.nand3_mag_1.OUT 1.17e-20
C691 JK_FF_mag_3.nand2_mag_1.IN2 a_8520_1353# 0.00372f
C692 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_0.OUT 0.0622f
C693 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C694 Q1 and2_mag_0.OUT 0.0529f
C695 JK_FF_mag_2.J JK_FF_mag_1.nand2_mag_3.IN1 1.48e-19
C696 a_6828_1309# JK_FF_mag_2.J 9.32e-19
C697 a_7574_2450# Q1 0.0105f
C698 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.J 0.0836f
C699 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C700 a_9510_2450# JK_FF_mag_0.J 0.0027f
C701 a_4369_212# a_4529_212# 0.0504f
C702 JK_FF_mag_3.nand2_mag_3.IN1 a_6822_212# 1.46e-19
C703 JK_FF_mag_2.nand3_mag_1.OUT a_4375_1353# 0.0202f
C704 JK_FF_mag_0.nand3_mag_2.OUT VDD 0.792f
C705 a_4939_1353# JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C706 a_628_212# VDD 0.0132f
C707 a_2076_256# VDD 0.00152f
C708 Vdiv10 Q3 0.242f
C709 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.Qb 0.198f
C710 a_5503_1353# JK_FF_mag_2.J 7.4e-19
C711 JK_FF_mag_0.nand2_mag_1.IN2 nor_3_mag_0.IN3 7.14e-19
C712 JK_FF_mag_3.nand3_mag_1.OUT and2_mag_0.GF_INV_MAG_0.IN 5.7e-20
C713 JK_FF_mag_0.nand3_mag_1.IN1 Q3 0.00393f
C714 JK_FF_mag_0.nand2_mag_1.IN2 Q0 5.08e-20
C715 a_11691_256# VSS 0.0675f
C716 a_11127_256# VSS 0.0676f
C717 a_10563_212# VSS 0.0343f
C718 a_10403_212# VSS 0.0881f
C719 a_9839_212# VSS 0.0343f
C720 a_9679_212# VSS 0.0881f
C721 a_8674_256# VSS 0.0675f
C722 a_8110_256# VSS 0.0676f
C723 a_7546_212# VSS 0.0343f
C724 a_7386_212# VSS 0.0881f
C725 a_6822_212# VSS 0.0343f
C726 a_6662_212# VSS 0.0881f
C727 a_5657_256# VSS 0.0675f
C728 a_5093_256# VSS 0.0676f
C729 a_4529_212# VSS 0.0343f
C730 a_4369_212# VSS 0.0881f
C731 a_3805_212# VSS 0.0343f
C732 a_3645_212# VSS 0.0881f
C733 a_2640_256# VSS 0.0675f
C734 a_2076_256# VSS 0.0676f
C735 a_1512_212# VSS 0.0343f
C736 a_1352_212# VSS 0.0881f
C737 a_788_212# VSS 0.0343f
C738 a_628_212# VSS 0.0881f
C739 JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C740 JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C741 JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.415f
C742 JK_FF_mag_3.nand3_mag_2.OUT VSS 0.539f
C743 JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C744 JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C745 JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.415f
C746 RST VSS 2.72f
C747 JK_FF_mag_1.nand3_mag_2.OUT VSS 0.539f
C748 a_11537_1353# VSS 0.0676f
C749 a_10973_1353# VSS 0.0676f
C750 a_10409_1353# VSS 0.0676f
C751 a_9845_1309# VSS 0.0343f
C752 a_9685_1309# VSS 0.0881f
C753 a_8520_1353# VSS 0.0676f
C754 a_7956_1353# VSS 0.0676f
C755 a_7392_1353# VSS 0.0676f
C756 a_6828_1309# VSS 0.0343f
C757 a_6668_1309# VSS 0.0881f
C758 a_5503_1353# VSS 0.0676f
C759 a_4939_1353# VSS 0.0676f
C760 a_4375_1353# VSS 0.0676f
C761 a_3811_1309# VSS 0.0343f
C762 a_3651_1309# VSS 0.0881f
C763 a_2486_1353# VSS 0.0676f
C764 a_1922_1353# VSS 0.0676f
C765 a_1358_1353# VSS 0.0676f
C766 a_794_1309# VSS 0.0343f
C767 a_634_1309# VSS 0.0881f
C768 JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C769 JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C770 JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C771 JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C772 JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C773 JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.413f
C774 JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.692f
C775 JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.724f
C776 JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C777 JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C778 JK_FF_mag_3.Qb VSS 0.877f
C779 JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C780 JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.695f
C781 JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.724f
C782 JK_FF_mag_2.nand3_mag_1.OUT VSS 0.809f
C783 JK_FF_mag_2.nand3_mag_0.OUT VSS 0.509f
C784 JK_FF_mag_2.Qb VSS 0.879f
C785 JK_FF_mag_2.J VSS 3.11f
C786 JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C787 JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.954f
C788 JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.724f
C789 JK_FF_mag_1.nand3_mag_1.OUT VSS 0.809f
C790 JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C791 JK_FF_mag_1.Qb VSS 0.901f
C792 CLK VSS 0.855f
C793 a_9510_2450# VSS 0.0679f
C794 Vdiv10 VSS 0.464f
C795 a_11738_2752# VSS 0.0371f
C796 a_11578_2752# VSS 0.038f
C797 a_8542_2450# VSS 0.0679f
C798 a_7574_2450# VSS 0.0676f
C799 Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.669f
C800 and2_mag_1.OUT VSS 0.706f
C801 JK_FF_mag_0.J VSS 0.634f
C802 and2_mag_1.GF_INV_MAG_0.IN VSS 0.435f
C803 Q0 VSS 3.75f
C804 and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C805 and2_mag_0.GF_INV_MAG_0.IN VSS 0.436f
C806 Q2 VSS 2.3f
C807 Q1 VSS 2.8f
C808 Q3 VSS 1.93f
C809 and2_mag_0.OUT VSS 0.91f
C810 nor_3_mag_0.IN3 VSS 0.337f
C811 VDD VSS 68.9f
C812 Q2.t11 VSS 0.0181f
C813 Q2.t4 VSS 0.0326f
C814 Q2.n0 VSS 0.062f
C815 Q2.n1 VSS 0.052f
C816 Q2.t9 VSS 0.0202f
C817 Q2.t3 VSS 0.0253f
C818 Q2.n2 VSS 0.0584f
C819 Q2.n3 VSS 0.135f
C820 Q2.n4 VSS 0.311f
C821 Q2.t6 VSS 0.0202f
C822 Q2.t12 VSS 0.0253f
C823 Q2.n5 VSS 0.0584f
C824 Q2.n6 VSS 0.261f
C825 Q2.n7 VSS 0.294f
C826 Q2.t5 VSS 0.0231f
C827 Q2.t7 VSS 0.0351f
C828 Q2.n8 VSS 0.0623f
C829 Q2.n9 VSS 0.244f
C830 Q2.t8 VSS 0.0202f
C831 Q2.t10 VSS 0.0253f
C832 Q2.n10 VSS 0.0584f
C833 Q2.n11 VSS 0.0363f
C834 Q2.n12 VSS 0.465f
C835 Q2.n13 VSS 0.144f
C836 Q2.n14 VSS 0.0191f
C837 Q2.t1 VSS 0.0158f
C838 Q2.n15 VSS 0.0158f
C839 Q2.n16 VSS 0.0433f
C840 Q2.n17 VSS 0.14f
C841 Q2.n18 VSS 0.0142f
C842 RST.t1 VSS 0.0207f
C843 RST.t3 VSS 0.0314f
C844 RST.n0 VSS 0.0555f
C845 RST.n1 VSS 0.00695f
C846 RST.n2 VSS 0.016f
C847 RST.n3 VSS 0.00256f
C848 RST.t4 VSS 0.0197f
C849 RST.n4 VSS 0.0181f
C850 RST.t5 VSS 0.0313f
C851 RST.n5 VSS 0.0384f
C852 RST.n6 VSS 3.04e-19
C853 RST.n7 VSS 0.00255f
C854 RST.n8 VSS 0.00241f
C855 RST.n9 VSS 0.0128f
C856 RST.t6 VSS 0.0207f
C857 RST.t7 VSS 0.0314f
C858 RST.n10 VSS 0.0555f
C859 RST.n11 VSS 0.0299f
C860 RST.t0 VSS 0.0207f
C861 RST.t2 VSS 0.0314f
C862 RST.n12 VSS 0.0555f
C863 RST.n13 VSS 0.303f
C864 RST.n14 VSS 0.943f
C865 RST.n15 VSS 0.781f
C866 RST.n16 VSS 0.0289f
C867 JK_FF_mag_2.J.n0 VSS 0.0867f
C868 JK_FF_mag_2.J.t4 VSS 0.0183f
C869 JK_FF_mag_2.J.t5 VSS 0.0229f
C870 JK_FF_mag_2.J.n1 VSS 0.0543f
C871 JK_FF_mag_2.J.t6 VSS 0.0322f
C872 JK_FF_mag_2.J.t8 VSS 0.0205f
C873 JK_FF_mag_2.J.n2 VSS 0.0569f
C874 JK_FF_mag_2.J.t3 VSS 0.0296f
C875 JK_FF_mag_2.J.t7 VSS 0.0228f
C876 JK_FF_mag_2.J.n3 VSS 0.0585f
C877 JK_FF_mag_2.J.n4 VSS 1.1f
C878 JK_FF_mag_2.J.n5 VSS 0.366f
C879 JK_FF_mag_2.J.t2 VSS 0.0143f
C880 JK_FF_mag_2.J.n6 VSS 0.0143f
C881 JK_FF_mag_2.J.n7 VSS 0.0338f
C882 Q0.t16 VSS 0.0237f
C883 Q0.t18 VSS 0.0359f
C884 Q0.n0 VSS 0.0634f
C885 Q0.n1 VSS 0.00818f
C886 Q0.n2 VSS 0.0103f
C887 Q0.t12 VSS 0.0297f
C888 Q0.t17 VSS 0.00758f
C889 Q0.n3 VSS 0.0491f
C890 Q0.n4 VSS 0.0104f
C891 Q0.n5 VSS 0.0213f
C892 Q0.n6 VSS 0.00363f
C893 Q0.n7 VSS 0.00321f
C894 Q0.n8 VSS 0.00596f
C895 Q0.t3 VSS 0.0237f
C896 Q0.t7 VSS 0.0359f
C897 Q0.n9 VSS 0.0634f
C898 Q0.n10 VSS 0.00818f
C899 Q0.n11 VSS 0.00298f
C900 Q0.n12 VSS 0.0116f
C901 Q0.n13 VSS 0.117f
C902 Q0.n14 VSS 0.119f
C903 Q0.n15 VSS 0.00596f
C904 Q0.t11 VSS 0.0237f
C905 Q0.t6 VSS 0.0359f
C906 Q0.n16 VSS 0.0634f
C907 Q0.n17 VSS 0.00818f
C908 Q0.n18 VSS 0.00294f
C909 Q0.n19 VSS 0.0719f
C910 Q0.n20 VSS 0.0942f
C911 Q0.n21 VSS 0.00938f
C912 Q0.t14 VSS 0.0334f
C913 Q0.t5 VSS 0.0184f
C914 Q0.n22 VSS 0.0634f
C915 Q0.n23 VSS 0.0127f
C916 Q0.n24 VSS 0.0102f
C917 Q0.n25 VSS 0.00403f
C918 Q0.n26 VSS 0.136f
C919 Q0.n27 VSS 0.825f
C920 Q0.n28 VSS 0.0195f
C921 Q0.t1 VSS 0.0161f
C922 Q0.n29 VSS 0.0161f
C923 Q0.n30 VSS 0.0443f
C924 Q0.n31 VSS 0.143f
C925 Q0.n32 VSS 0.0145f
C926 Q0.t8 VSS 0.0237f
C927 Q0.t10 VSS 0.0359f
C928 Q0.n33 VSS 0.0638f
C929 Q0.n34 VSS 0.25f
C930 Q0.t20 VSS 0.0206f
C931 Q0.t9 VSS 0.0258f
C932 Q0.n35 VSS 0.0598f
C933 Q0.n36 VSS 0.0371f
C934 Q0.n37 VSS 0.476f
C935 Q0.n38 VSS 0.121f
C936 Q0.n39 VSS 0.0507f
C937 Q0.t4 VSS 0.0297f
C938 Q0.t13 VSS 0.00758f
C939 Q0.n40 VSS 0.0491f
C940 Q0.n41 VSS 0.0104f
C941 Q0.n42 VSS 0.0213f
C942 Q0.n43 VSS 0.00363f
C943 Q0.n44 VSS 0.00183f
C944 Q0.n45 VSS 0.754f
C945 Q0.n46 VSS 0.00596f
C946 Q0.t19 VSS 0.0237f
C947 Q0.t15 VSS 0.0359f
C948 Q0.n47 VSS 0.0634f
C949 Q0.n48 VSS 0.00818f
C950 Q0.n49 VSS 0.00294f
C951 Q0.n50 VSS 0.0843f
C952 Q0.n51 VSS 0.119f
C953 Q0.n52 VSS 0.0116f
C954 Q0.n53 VSS 0.117f
C955 Q0.n54 VSS 0.00298f
C956 Q0.n55 VSS 0.00596f
C957 VDD.t146 VSS 0.00515f
C958 VDD.t61 VSS 0.0237f
C959 VDD.n0 VSS 0.00514f
C960 VDD.t25 VSS 0.00515f
C961 VDD.n1 VSS 0.00514f
C962 VDD.n2 VSS 0.0255f
C963 VDD.t158 VSS 0.0541f
C964 VDD.n3 VSS 0.00514f
C965 VDD.t186 VSS 0.00513f
C966 VDD.t97 VSS 0.00515f
C967 VDD.n4 VSS 0.0243f
C968 VDD.t96 VSS 0.028f
C969 VDD.t125 VSS 0.0365f
C970 VDD.n5 VSS 0.00514f
C971 VDD.t126 VSS 0.00515f
C972 VDD.n6 VSS 0.00514f
C973 VDD.n7 VSS 0.0255f
C974 VDD.t192 VSS 0.0541f
C975 VDD.n8 VSS 0.00514f
C976 VDD.t15 VSS 0.00513f
C977 VDD.t166 VSS 0.00515f
C978 VDD.n9 VSS 0.0243f
C979 VDD.t14 VSS 0.0454f
C980 VDD.t129 VSS 0.0352f
C981 VDD.t58 VSS 0.00212f
C982 VDD.n10 VSS 0.00212f
C983 VDD.n11 VSS 0.00462f
C984 VDD.t151 VSS 0.00515f
C985 VDD.n12 VSS 0.00514f
C986 VDD.n13 VSS 0.0255f
C987 VDD.t211 VSS 0.068f
C988 VDD.n14 VSS 0.00514f
C989 VDD.t141 VSS 0.00515f
C990 VDD.n15 VSS 0.00514f
C991 VDD.n16 VSS 0.00514f
C992 VDD.t142 VSS 0.067f
C993 VDD.n17 VSS 0.0319f
C994 VDD.t111 VSS 0.00515f
C995 VDD.n18 VSS 0.00514f
C996 VDD.t110 VSS 0.0621f
C997 VDD.t208 VSS 0.068f
C998 VDD.n19 VSS 0.0319f
C999 VDD.t51 VSS 0.00515f
C1000 VDD.t39 VSS 0.00212f
C1001 VDD.n20 VSS 0.00212f
C1002 VDD.n21 VSS 0.00462f
C1003 VDD.t50 VSS 0.0621f
C1004 VDD.t38 VSS 0.0758f
C1005 VDD.t82 VSS 0.0352f
C1006 VDD.n22 VSS 0.0319f
C1007 VDD.t32 VSS 0.00515f
C1008 VDD.t79 VSS 0.00212f
C1009 VDD.n23 VSS 0.00212f
C1010 VDD.n24 VSS 0.00462f
C1011 VDD.t31 VSS 0.0621f
C1012 VDD.t78 VSS 0.0758f
C1013 VDD.t75 VSS 0.0352f
C1014 VDD.t93 VSS 0.0619f
C1015 VDD.n25 VSS 0.0319f
C1016 VDD.t94 VSS 0.00481f
C1017 VDD.t92 VSS 0.00442f
C1018 VDD.t232 VSS 0.00335f
C1019 VDD.n26 VSS 0.00862f
C1020 VDD.n27 VSS 0.00153f
C1021 VDD.t107 VSS 0.00442f
C1022 VDD.t227 VSS 0.00335f
C1023 VDD.n28 VSS 0.00863f
C1024 VDD.n29 VSS 0.00203f
C1025 VDD.n30 VSS 0.00105f
C1026 VDD.n31 VSS 5.29e-19
C1027 VDD.n32 VSS 0.00472f
C1028 VDD.n33 VSS 5.09e-19
C1029 VDD.t101 VSS 0.00429f
C1030 VDD.n34 VSS 0.00423f
C1031 VDD.t230 VSS 0.00334f
C1032 VDD.n35 VSS 0.00143f
C1033 VDD.n36 VSS 0.00453f
C1034 VDD.n37 VSS 0.00156f
C1035 VDD.n38 VSS 0.00128f
C1036 VDD.t104 VSS 0.00439f
C1037 VDD.t228 VSS 0.00335f
C1038 VDD.n39 VSS 0.00865f
C1039 VDD.n40 VSS 0.00162f
C1040 VDD.n41 VSS 0.00137f
C1041 VDD.n42 VSS 5.29e-19
C1042 VDD.n43 VSS 0.0167f
C1043 VDD.n44 VSS 0.0647f
C1044 VDD.n45 VSS 0.0945f
C1045 VDD.t231 VSS 0.00341f
C1046 VDD.t98 VSS 0.00434f
C1047 VDD.n46 VSS 0.00864f
C1048 VDD.n47 VSS 0.00315f
C1049 VDD.n48 VSS 0.00128f
C1050 VDD.t229 VSS 0.00335f
C1051 VDD.t95 VSS 0.00439f
C1052 VDD.n49 VSS 0.00865f
C1053 VDD.n50 VSS 0.00168f
C1054 VDD.n51 VSS 0.00133f
C1055 VDD.n52 VSS 5.29e-19
C1056 VDD.n53 VSS 0.0167f
C1057 VDD.n54 VSS 0.0218f
C1058 VDD.n55 VSS 0.105f
C1059 VDD.n56 VSS 0.0441f
C1060 VDD.n57 VSS 0.00417f
C1061 VDD.n58 VSS 0.012f
C1062 VDD.n59 VSS 0.0294f
C1063 VDD.n60 VSS 0.0293f
C1064 VDD.n61 VSS 0.0301f
C1065 VDD.n62 VSS 0.016f
C1066 VDD.n63 VSS 0.0293f
C1067 VDD.n64 VSS 0.03f
C1068 VDD.n65 VSS 0.0178f
C1069 VDD.n66 VSS 0.0255f
C1070 VDD.n67 VSS 0.0237f
C1071 VDD.n68 VSS 0.0178f
C1072 VDD.n69 VSS 0.0485f
C1073 VDD.n70 VSS 0.0552f
C1074 VDD.t147 VSS 0.067f
C1075 VDD.t140 VSS 0.0621f
C1076 VDD.n71 VSS 0.0319f
C1077 VDD.n72 VSS 0.0178f
C1078 VDD.n73 VSS 0.0237f
C1079 VDD.n74 VSS 0.0255f
C1080 VDD.t41 VSS 0.00515f
C1081 VDD.n75 VSS 0.0237f
C1082 VDD.n76 VSS 0.0178f
C1083 VDD.n77 VSS 0.0319f
C1084 VDD.t40 VSS 0.0621f
C1085 VDD.t52 VSS 0.068f
C1086 VDD.t57 VSS 0.0758f
C1087 VDD.t150 VSS 0.0621f
C1088 VDD.n78 VSS 0.0319f
C1089 VDD.n79 VSS 0.0178f
C1090 VDD.n80 VSS 0.0224f
C1091 VDD.n81 VSS 0.021f
C1092 VDD.n82 VSS 0.016f
C1093 VDD.n83 VSS 0.0319f
C1094 VDD.t165 VSS 0.0352f
C1095 VDD.n84 VSS 0.0478f
C1096 VDD.n85 VSS 0.0161f
C1097 VDD.n86 VSS 0.00514f
C1098 VDD.t152 VSS 0.067f
C1099 VDD.n87 VSS 0.0319f
C1100 VDD.t13 VSS 0.00515f
C1101 VDD.n88 VSS 0.00514f
C1102 VDD.t12 VSS 0.0621f
C1103 VDD.t121 VSS 0.068f
C1104 VDD.n89 VSS 0.0319f
C1105 VDD.t49 VSS 0.00515f
C1106 VDD.t128 VSS 0.00212f
C1107 VDD.n90 VSS 0.00212f
C1108 VDD.n91 VSS 0.00462f
C1109 VDD.t48 VSS 0.0621f
C1110 VDD.t127 VSS 0.0758f
C1111 VDD.t200 VSS 0.0352f
C1112 VDD.n92 VSS 0.0319f
C1113 VDD.t91 VSS 0.00515f
C1114 VDD.t21 VSS 0.00212f
C1115 VDD.n93 VSS 0.00212f
C1116 VDD.n94 VSS 0.00462f
C1117 VDD.t90 VSS 0.0621f
C1118 VDD.t20 VSS 0.0758f
C1119 VDD.t177 VSS 0.0352f
C1120 VDD.t99 VSS 0.0619f
C1121 VDD.n95 VSS 0.0319f
C1122 VDD.t100 VSS 0.00552f
C1123 VDD.n96 VSS 0.0396f
C1124 VDD.n97 VSS 0.0293f
C1125 VDD.n98 VSS 0.0301f
C1126 VDD.n99 VSS 0.016f
C1127 VDD.n100 VSS 0.0293f
C1128 VDD.n101 VSS 0.03f
C1129 VDD.n102 VSS 0.0178f
C1130 VDD.n103 VSS 0.0255f
C1131 VDD.n104 VSS 0.0237f
C1132 VDD.n105 VSS 0.0178f
C1133 VDD.n106 VSS 0.0456f
C1134 VDD.n107 VSS 0.0364f
C1135 VDD.n108 VSS 0.0261f
C1136 VDD.t139 VSS 0.00515f
C1137 VDD.n109 VSS 0.0237f
C1138 VDD.n110 VSS 0.0178f
C1139 VDD.n111 VSS 0.0275f
C1140 VDD.t138 VSS 0.0494f
C1141 VDD.t118 VSS 0.0541f
C1142 VDD.n112 VSS 0.0275f
C1143 VDD.n113 VSS 0.0178f
C1144 VDD.n114 VSS 0.0237f
C1145 VDD.n115 VSS 0.0255f
C1146 VDD.n116 VSS 0.0178f
C1147 VDD.t196 VSS 0.00212f
C1148 VDD.n117 VSS 0.00212f
C1149 VDD.n118 VSS 0.00462f
C1150 VDD.t184 VSS 0.00515f
C1151 VDD.n119 VSS 0.00514f
C1152 VDD.n120 VSS 0.0253f
C1153 VDD.t226 VSS 0.00513f
C1154 VDD.n121 VSS 0.0181f
C1155 VDD.t225 VSS 0.0456f
C1156 VDD.t174 VSS 0.0406f
C1157 VDD.n122 VSS 0.00514f
C1158 VDD.t115 VSS 0.00513f
C1159 VDD.t81 VSS 0.00515f
C1160 VDD.n123 VSS 0.024f
C1161 VDD.t114 VSS 0.0456f
C1162 VDD.t85 VSS 0.0406f
C1163 VDD.n124 VSS 0.00514f
C1164 VDD.t215 VSS 0.00513f
C1165 VDD.t217 VSS 0.00522f
C1166 VDD.n125 VSS 0.028f
C1167 VDD.t112 VSS 0.0658f
C1168 VDD.t113 VSS 0.00513f
C1169 VDD.t117 VSS 0.02f
C1170 VDD.n126 VSS 0.0401f
C1171 VDD.t124 VSS 0.131f
C1172 VDD.t44 VSS 0.0417f
C1173 VDD.n127 VSS 0.0484f
C1174 VDD.t116 VSS 0.133f
C1175 VDD.n128 VSS 0.0623f
C1176 VDD.n129 VSS 0.0243f
C1177 VDD.n130 VSS 0.0169f
C1178 VDD.n131 VSS 0.0725f
C1179 VDD.t216 VSS 0.0429f
C1180 VDD.t214 VSS 0.0727f
C1181 VDD.n132 VSS 0.0475f
C1182 VDD.n133 VSS 0.0181f
C1183 VDD.n134 VSS 0.0253f
C1184 VDD.n135 VSS 0.018f
C1185 VDD.n136 VSS 0.0319f
C1186 VDD.t80 VSS 0.0352f
C1187 VDD.n137 VSS 0.0748f
C1188 VDD.n138 VSS 0.0181f
C1189 VDD.n139 VSS 0.0253f
C1190 VDD.t19 VSS 0.00515f
C1191 VDD.n140 VSS 0.024f
C1192 VDD.n141 VSS 0.018f
C1193 VDD.n142 VSS 0.0319f
C1194 VDD.t18 VSS 0.0352f
C1195 VDD.n143 VSS 0.0748f
C1196 VDD.t155 VSS 0.0406f
C1197 VDD.t183 VSS 0.0619f
C1198 VDD.n144 VSS 0.0319f
C1199 VDD.n145 VSS 0.018f
C1200 VDD.n146 VSS 0.0648f
C1201 VDD.t168 VSS 0.00515f
C1202 VDD.n147 VSS 0.0169f
C1203 VDD.n148 VSS 0.0545f
C1204 VDD.n149 VSS 0.021f
C1205 VDD.n150 VSS 0.016f
C1206 VDD.n151 VSS 0.0275f
C1207 VDD.t180 VSS 0.028f
C1208 VDD.t195 VSS 0.0603f
C1209 VDD.t167 VSS 0.0494f
C1210 VDD.n152 VSS 0.0275f
C1211 VDD.t45 VSS 0.0237f
C1212 VDD.n153 VSS 0.143f
C1213 VDD.n154 VSS 0.0789f
C1214 VDD.t185 VSS 0.0567f
C1215 VDD.n155 VSS 0.0161f
C1216 VDD.n156 VSS 0.00514f
C1217 VDD.t187 VSS 0.067f
C1218 VDD.n157 VSS 0.0319f
C1219 VDD.t89 VSS 0.00515f
C1220 VDD.n158 VSS 0.00514f
C1221 VDD.t88 VSS 0.0621f
C1222 VDD.t132 VSS 0.068f
C1223 VDD.n159 VSS 0.0319f
C1224 VDD.t65 VSS 0.00515f
C1225 VDD.t23 VSS 0.00212f
C1226 VDD.n160 VSS 0.00212f
C1227 VDD.n161 VSS 0.00462f
C1228 VDD.t64 VSS 0.0621f
C1229 VDD.t22 VSS 0.0758f
C1230 VDD.t28 VSS 0.0352f
C1231 VDD.n162 VSS 0.0319f
C1232 VDD.t43 VSS 0.00515f
C1233 VDD.t191 VSS 0.00212f
C1234 VDD.n163 VSS 0.00212f
C1235 VDD.n164 VSS 0.00462f
C1236 VDD.t42 VSS 0.0621f
C1237 VDD.t190 VSS 0.0758f
C1238 VDD.t0 VSS 0.0352f
C1239 VDD.t108 VSS 0.0619f
C1240 VDD.n165 VSS 0.0319f
C1241 VDD.t109 VSS 0.00552f
C1242 VDD.n166 VSS 0.0396f
C1243 VDD.n167 VSS 0.0293f
C1244 VDD.n168 VSS 0.0301f
C1245 VDD.n169 VSS 0.016f
C1246 VDD.n170 VSS 0.0293f
C1247 VDD.n171 VSS 0.03f
C1248 VDD.n172 VSS 0.0178f
C1249 VDD.n173 VSS 0.0255f
C1250 VDD.n174 VSS 0.0237f
C1251 VDD.n175 VSS 0.0178f
C1252 VDD.n176 VSS 0.0456f
C1253 VDD.n177 VSS 0.0364f
C1254 VDD.n178 VSS 0.0261f
C1255 VDD.t60 VSS 0.00515f
C1256 VDD.n179 VSS 0.0237f
C1257 VDD.n180 VSS 0.0178f
C1258 VDD.n181 VSS 0.0275f
C1259 VDD.t59 VSS 0.0494f
C1260 VDD.t135 VSS 0.0541f
C1261 VDD.n182 VSS 0.143f
C1262 VDD.t24 VSS 0.0365f
C1263 VDD.n183 VSS 0.0275f
C1264 VDD.n184 VSS 0.0178f
C1265 VDD.n185 VSS 0.0237f
C1266 VDD.n186 VSS 0.0255f
C1267 VDD.t56 VSS 0.00515f
C1268 VDD.t162 VSS 0.00212f
C1269 VDD.n187 VSS 0.00212f
C1270 VDD.n188 VSS 0.00462f
C1271 VDD.n189 VSS 0.021f
C1272 VDD.n190 VSS 0.0224f
C1273 VDD.n191 VSS 0.0178f
C1274 VDD.n192 VSS 0.0275f
C1275 VDD.t55 VSS 0.0494f
C1276 VDD.t161 VSS 0.0603f
C1277 VDD.t205 VSS 0.028f
C1278 VDD.t145 VSS 0.028f
C1279 VDD.n193 VSS 0.0275f
C1280 VDD.n194 VSS 0.016f
C1281 VDD.n195 VSS 0.0243f
C1282 VDD.n196 VSS 0.0789f
C1283 VDD.t16 VSS 0.0567f
C1284 VDD.t17 VSS 0.00513f
C1285 VDD.n197 VSS 0.00514f
C1286 VDD.t3 VSS 0.0541f
C1287 VDD.n198 VSS 0.0275f
C1288 VDD.t11 VSS 0.00515f
C1289 VDD.n199 VSS 0.00514f
C1290 VDD.t10 VSS 0.0494f
C1291 VDD.t69 VSS 0.0541f
C1292 VDD.n200 VSS 0.0275f
C1293 VDD.t224 VSS 0.00515f
C1294 VDD.n201 VSS 0.00514f
C1295 VDD.n202 VSS 0.0275f
C1296 VDD.t27 VSS 0.00515f
C1297 VDD.t7 VSS 0.00212f
C1298 VDD.n203 VSS 0.00212f
C1299 VDD.n204 VSS 0.00462f
C1300 VDD.t26 VSS 0.0494f
C1301 VDD.t6 VSS 0.0603f
C1302 VDD.t169 VSS 0.028f
C1303 VDD.n205 VSS 0.0275f
C1304 VDD.t106 VSS 0.00515f
C1305 VDD.t223 VSS 0.0365f
C1306 VDD.t35 VSS 0.0237f
C1307 VDD.n206 VSS 0.143f
C1308 VDD.t105 VSS 0.028f
C1309 VDD.n207 VSS 0.0789f
C1310 VDD.t203 VSS 0.0567f
C1311 VDD.t204 VSS 0.00537f
C1312 VDD.n208 VSS 0.0243f
C1313 VDD.n209 VSS 0.016f
C1314 VDD.n210 VSS 0.021f
C1315 VDD.n211 VSS 0.0224f
C1316 VDD.n212 VSS 0.0178f
C1317 VDD.n213 VSS 0.0255f
C1318 VDD.n214 VSS 0.0237f
C1319 VDD.n215 VSS 0.0178f
C1320 VDD.n216 VSS 0.0255f
C1321 VDD.n217 VSS 0.0237f
C1322 VDD.n218 VSS 0.0178f
C1323 VDD.n219 VSS 0.0261f
C1324 VDD.n220 VSS 0.00514f
C1325 VDD.t72 VSS 0.067f
C1326 VDD.n221 VSS 0.0319f
C1327 VDD.t164 VSS 0.00515f
C1328 VDD.n222 VSS 0.00514f
C1329 VDD.t163 VSS 0.0621f
C1330 VDD.t66 VSS 0.068f
C1331 VDD.n223 VSS 0.0319f
C1332 VDD.t34 VSS 0.00515f
C1333 VDD.t222 VSS 0.00212f
C1334 VDD.n224 VSS 0.00212f
C1335 VDD.n225 VSS 0.00462f
C1336 VDD.t33 VSS 0.0621f
C1337 VDD.t221 VSS 0.0758f
C1338 VDD.t197 VSS 0.0352f
C1339 VDD.n226 VSS 0.0319f
C1340 VDD.t9 VSS 0.00515f
C1341 VDD.t173 VSS 0.00212f
C1342 VDD.n227 VSS 0.00212f
C1343 VDD.n228 VSS 0.00462f
C1344 VDD.t8 VSS 0.0621f
C1345 VDD.t172 VSS 0.0758f
C1346 VDD.t218 VSS 0.0352f
C1347 VDD.t102 VSS 0.0619f
C1348 VDD.n229 VSS 0.0319f
C1349 VDD.t103 VSS 0.00552f
C1350 VDD.n230 VSS 0.0396f
C1351 VDD.n231 VSS 0.0293f
C1352 VDD.n232 VSS 0.0301f
C1353 VDD.n233 VSS 0.016f
C1354 VDD.n234 VSS 0.0293f
C1355 VDD.n235 VSS 0.03f
C1356 VDD.n236 VSS 0.0178f
C1357 VDD.n237 VSS 0.0255f
C1358 VDD.n238 VSS 0.0237f
C1359 VDD.n239 VSS 0.0178f
C1360 VDD.n240 VSS 0.0456f
C1361 VDD.n241 VSS 0.0324f
C1362 VDD.n242 VSS 0.0158f
C1363 Q1.t14 VSS 0.028f
C1364 Q1.t15 VSS 0.0425f
C1365 Q1.n0 VSS 0.075f
C1366 Q1.n1 VSS 0.00967f
C1367 Q1.n2 VSS 0.00683f
C1368 Q1.n3 VSS 0.0231f
C1369 Q1.t1 VSS 0.0191f
C1370 Q1.n4 VSS 0.0191f
C1371 Q1.n5 VSS 0.0523f
C1372 Q1.n6 VSS 0.169f
C1373 Q1.n7 VSS 0.0172f
C1374 Q1.t3 VSS 0.028f
C1375 Q1.t4 VSS 0.0425f
C1376 Q1.n8 VSS 0.0754f
C1377 Q1.n9 VSS 0.296f
C1378 Q1.t5 VSS 0.0244f
C1379 Q1.t7 VSS 0.0305f
C1380 Q1.n10 VSS 0.0706f
C1381 Q1.n11 VSS 0.0439f
C1382 Q1.n12 VSS 0.563f
C1383 Q1.n13 VSS 0.143f
C1384 Q1.n14 VSS 0.0612f
C1385 Q1.t8 VSS 0.0351f
C1386 Q1.t13 VSS 0.00896f
C1387 Q1.n15 VSS 0.0581f
C1388 Q1.n16 VSS 0.0123f
C1389 Q1.n17 VSS 0.0252f
C1390 Q1.n18 VSS 0.00429f
C1391 Q1.n19 VSS 0.0873f
C1392 Q1.n20 VSS 0.0832f
C1393 Q1.n21 VSS 0.0124f
C1394 Q1.n22 VSS 0.00623f
C1395 Q1.t16 VSS 0.0244f
C1396 Q1.t9 VSS 0.0305f
C1397 Q1.n23 VSS 0.0687f
C1398 Q1.n24 VSS 0.0303f
C1399 Q1.n25 VSS 0.00345f
C1400 Q1.n26 VSS 0.25f
C1401 Q1.n27 VSS 0.0134f
C1402 Q1.t11 VSS 0.0398f
C1403 Q1.t6 VSS 0.0217f
C1404 Q1.n28 VSS 0.0748f
C1405 Q1.n29 VSS 0.0179f
C1406 Q1.n30 VSS 0.0097f
C1407 Q1.n31 VSS 0.00476f
C1408 Q1.n32 VSS 0.0852f
C1409 Q1.n33 VSS 0.501f
C1410 Q1.n34 VSS 0.132f
C1411 Q1.n35 VSS 2.25e-19
C1412 Q1.n36 VSS -7.03e-19
C1413 Q1.n37 VSS 0.00306f
C1414 Q1.n38 VSS 0.00412f
C1415 Q1.n39 VSS 0.00381f
C1416 Q1.t12 VSS 0.028f
C1417 Q1.t10 VSS 0.0425f
C1418 Q1.n40 VSS 0.075f
C1419 Q1.n41 VSS 0.00914f
C1420 Q1.n42 VSS 5.31e-19
C1421 Q1.n43 VSS 0.00332f
C1422 Q1.n44 VSS 0.14f
C1423 Q1.n45 VSS 0.0137f
C1424 Q1.n46 VSS 0.136f
C1425 Q1.n47 VSS 0.00352f
C1426 Q1.n48 VSS 0.00705f
.ends

