** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/LSB_V1 _PEX_TB.sch
**.subckt LSB_V1 _PEX_TB
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
V6 B4 VSS pulse(0 3.3 0 10p 10p 400n 800n)
.save i(v6)
V7 B5 VSS pulse(0 3.3 0 10p 10p 800n 1.6u)
.save i(v7)
V8 B6 VSS pulse(0 3.3 0 10p 10p 1.6u 3.2u)
.save i(v8)
V10 B3 VSS pulse(0 3.3 0 10p 10p 200n 400n)
.save i(v10)
V11 B2 VSS pulse(0 3.3 0 10p 10p 100n 200n)
.save i(v11)
V12 B1 VSS pulse(0 3.3 0 10p 10p 50n 100n)
.save i(v12)
I0 VDD ITAIL 2.5u
R1 VDD OUT+ 10k m=1
R2 VDD OUT- 10k m=1
V3 net1 VSS 0
.save i(v3)
V4 net2 VSS 0
.save i(v4)
V5 net3 VSS 0
.save i(v5)
V9 net4 VSS 3.3
.save i(v9)
V13 net5 VSS 0
.save i(v13)
V14 net6 VSS 0
.save i(v14)
x1 VDD VSS B1 B2 B3 B4 B5 B6 ITAIL OUT+ OUT- net8 net9 net10 net11 net12 net13 pex_LSBs_magic
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_LSBs_magic.spice
.option savecurrents
.control
save all
op

tran 10n 3.2u
plot v(OUT+) v(OUT-)
write LSB_TB.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
