magic
tech gf180mcuC
magscale 1 10
timestamp 1691396512
<< pwell >>
rect -460 -804 460 804
<< nmos >>
rect -348 336 -292 736
rect -188 336 -132 736
rect -28 336 28 736
rect 132 336 188 736
rect 292 336 348 736
rect -348 -200 -292 200
rect -188 -200 -132 200
rect -28 -200 28 200
rect 132 -200 188 200
rect 292 -200 348 200
rect -348 -736 -292 -336
rect -188 -736 -132 -336
rect -28 -736 28 -336
rect 132 -736 188 -336
rect 292 -736 348 -336
<< ndiff >>
rect -436 723 -348 736
rect -436 349 -423 723
rect -377 349 -348 723
rect -436 336 -348 349
rect -292 723 -188 736
rect -292 349 -263 723
rect -217 349 -188 723
rect -292 336 -188 349
rect -132 723 -28 736
rect -132 349 -103 723
rect -57 349 -28 723
rect -132 336 -28 349
rect 28 723 132 736
rect 28 349 57 723
rect 103 349 132 723
rect 28 336 132 349
rect 188 723 292 736
rect 188 349 217 723
rect 263 349 292 723
rect 188 336 292 349
rect 348 723 436 736
rect 348 349 377 723
rect 423 349 436 723
rect 348 336 436 349
rect -436 187 -348 200
rect -436 -187 -423 187
rect -377 -187 -348 187
rect -436 -200 -348 -187
rect -292 187 -188 200
rect -292 -187 -263 187
rect -217 -187 -188 187
rect -292 -200 -188 -187
rect -132 187 -28 200
rect -132 -187 -103 187
rect -57 -187 -28 187
rect -132 -200 -28 -187
rect 28 187 132 200
rect 28 -187 57 187
rect 103 -187 132 187
rect 28 -200 132 -187
rect 188 187 292 200
rect 188 -187 217 187
rect 263 -187 292 187
rect 188 -200 292 -187
rect 348 187 436 200
rect 348 -187 377 187
rect 423 -187 436 187
rect 348 -200 436 -187
rect -436 -349 -348 -336
rect -436 -723 -423 -349
rect -377 -723 -348 -349
rect -436 -736 -348 -723
rect -292 -349 -188 -336
rect -292 -723 -263 -349
rect -217 -723 -188 -349
rect -292 -736 -188 -723
rect -132 -349 -28 -336
rect -132 -723 -103 -349
rect -57 -723 -28 -349
rect -132 -736 -28 -723
rect 28 -349 132 -336
rect 28 -723 57 -349
rect 103 -723 132 -349
rect 28 -736 132 -723
rect 188 -349 292 -336
rect 188 -723 217 -349
rect 263 -723 292 -349
rect 188 -736 292 -723
rect 348 -349 436 -336
rect 348 -723 377 -349
rect 423 -723 436 -349
rect 348 -736 436 -723
<< ndiffc >>
rect -423 349 -377 723
rect -263 349 -217 723
rect -103 349 -57 723
rect 57 349 103 723
rect 217 349 263 723
rect 377 349 423 723
rect -423 -187 -377 187
rect -263 -187 -217 187
rect -103 -187 -57 187
rect 57 -187 103 187
rect 217 -187 263 187
rect 377 -187 423 187
rect -423 -723 -377 -349
rect -263 -723 -217 -349
rect -103 -723 -57 -349
rect 57 -723 103 -349
rect 217 -723 263 -349
rect 377 -723 423 -349
<< polysilicon >>
rect -348 736 -292 780
rect -188 736 -132 780
rect -28 736 28 780
rect 132 736 188 780
rect 292 736 348 780
rect -348 292 -292 336
rect -188 292 -132 336
rect -28 292 28 336
rect 132 292 188 336
rect 292 292 348 336
rect -348 200 -292 244
rect -188 200 -132 244
rect -28 200 28 244
rect 132 200 188 244
rect 292 200 348 244
rect -348 -244 -292 -200
rect -188 -244 -132 -200
rect -28 -244 28 -200
rect 132 -244 188 -200
rect 292 -244 348 -200
rect -348 -336 -292 -292
rect -188 -336 -132 -292
rect -28 -336 28 -292
rect 132 -336 188 -292
rect 292 -336 348 -292
rect -348 -780 -292 -736
rect -188 -780 -132 -736
rect -28 -780 28 -736
rect 132 -780 188 -736
rect 292 -780 348 -736
<< metal1 >>
rect -423 723 -377 734
rect -423 338 -377 349
rect -263 723 -217 734
rect -263 338 -217 349
rect -103 723 -57 734
rect -103 338 -57 349
rect 57 723 103 734
rect 57 338 103 349
rect 217 723 263 734
rect 217 338 263 349
rect 377 723 423 734
rect 377 338 423 349
rect -423 187 -377 198
rect -423 -198 -377 -187
rect -263 187 -217 198
rect -263 -198 -217 -187
rect -103 187 -57 198
rect -103 -198 -57 -187
rect 57 187 103 198
rect 57 -198 103 -187
rect 217 187 263 198
rect 217 -198 263 -187
rect 377 187 423 198
rect 377 -198 423 -187
rect -423 -349 -377 -338
rect -423 -734 -377 -723
rect -263 -349 -217 -338
rect -263 -734 -217 -723
rect -103 -349 -57 -338
rect -103 -734 -57 -723
rect 57 -349 103 -338
rect 57 -734 103 -723
rect 217 -349 263 -338
rect 217 -734 263 -723
rect 377 -349 423 -338
rect 377 -734 423 -723
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 2 l 0.280 m 3 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
