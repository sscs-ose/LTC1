magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -3230 -1349 3230 1349
<< metal3 >>
rect -2230 344 2230 349
rect -2230 316 -2225 344
rect -2197 316 -2159 344
rect -2131 316 -2093 344
rect -2065 316 -2027 344
rect -1999 316 -1961 344
rect -1933 316 -1895 344
rect -1867 316 -1829 344
rect -1801 316 -1763 344
rect -1735 316 -1697 344
rect -1669 316 -1631 344
rect -1603 316 -1565 344
rect -1537 316 -1499 344
rect -1471 316 -1433 344
rect -1405 316 -1367 344
rect -1339 316 -1301 344
rect -1273 316 -1235 344
rect -1207 316 -1169 344
rect -1141 316 -1103 344
rect -1075 316 -1037 344
rect -1009 316 -971 344
rect -943 316 -905 344
rect -877 316 -839 344
rect -811 316 -773 344
rect -745 316 -707 344
rect -679 316 -641 344
rect -613 316 -575 344
rect -547 316 -509 344
rect -481 316 -443 344
rect -415 316 -377 344
rect -349 316 -311 344
rect -283 316 -245 344
rect -217 316 -179 344
rect -151 316 -113 344
rect -85 316 -47 344
rect -19 316 19 344
rect 47 316 85 344
rect 113 316 151 344
rect 179 316 217 344
rect 245 316 283 344
rect 311 316 349 344
rect 377 316 415 344
rect 443 316 481 344
rect 509 316 547 344
rect 575 316 613 344
rect 641 316 679 344
rect 707 316 745 344
rect 773 316 811 344
rect 839 316 877 344
rect 905 316 943 344
rect 971 316 1009 344
rect 1037 316 1075 344
rect 1103 316 1141 344
rect 1169 316 1207 344
rect 1235 316 1273 344
rect 1301 316 1339 344
rect 1367 316 1405 344
rect 1433 316 1471 344
rect 1499 316 1537 344
rect 1565 316 1603 344
rect 1631 316 1669 344
rect 1697 316 1735 344
rect 1763 316 1801 344
rect 1829 316 1867 344
rect 1895 316 1933 344
rect 1961 316 1999 344
rect 2027 316 2065 344
rect 2093 316 2131 344
rect 2159 316 2197 344
rect 2225 316 2230 344
rect -2230 278 2230 316
rect -2230 250 -2225 278
rect -2197 250 -2159 278
rect -2131 250 -2093 278
rect -2065 250 -2027 278
rect -1999 250 -1961 278
rect -1933 250 -1895 278
rect -1867 250 -1829 278
rect -1801 250 -1763 278
rect -1735 250 -1697 278
rect -1669 250 -1631 278
rect -1603 250 -1565 278
rect -1537 250 -1499 278
rect -1471 250 -1433 278
rect -1405 250 -1367 278
rect -1339 250 -1301 278
rect -1273 250 -1235 278
rect -1207 250 -1169 278
rect -1141 250 -1103 278
rect -1075 250 -1037 278
rect -1009 250 -971 278
rect -943 250 -905 278
rect -877 250 -839 278
rect -811 250 -773 278
rect -745 250 -707 278
rect -679 250 -641 278
rect -613 250 -575 278
rect -547 250 -509 278
rect -481 250 -443 278
rect -415 250 -377 278
rect -349 250 -311 278
rect -283 250 -245 278
rect -217 250 -179 278
rect -151 250 -113 278
rect -85 250 -47 278
rect -19 250 19 278
rect 47 250 85 278
rect 113 250 151 278
rect 179 250 217 278
rect 245 250 283 278
rect 311 250 349 278
rect 377 250 415 278
rect 443 250 481 278
rect 509 250 547 278
rect 575 250 613 278
rect 641 250 679 278
rect 707 250 745 278
rect 773 250 811 278
rect 839 250 877 278
rect 905 250 943 278
rect 971 250 1009 278
rect 1037 250 1075 278
rect 1103 250 1141 278
rect 1169 250 1207 278
rect 1235 250 1273 278
rect 1301 250 1339 278
rect 1367 250 1405 278
rect 1433 250 1471 278
rect 1499 250 1537 278
rect 1565 250 1603 278
rect 1631 250 1669 278
rect 1697 250 1735 278
rect 1763 250 1801 278
rect 1829 250 1867 278
rect 1895 250 1933 278
rect 1961 250 1999 278
rect 2027 250 2065 278
rect 2093 250 2131 278
rect 2159 250 2197 278
rect 2225 250 2230 278
rect -2230 212 2230 250
rect -2230 184 -2225 212
rect -2197 184 -2159 212
rect -2131 184 -2093 212
rect -2065 184 -2027 212
rect -1999 184 -1961 212
rect -1933 184 -1895 212
rect -1867 184 -1829 212
rect -1801 184 -1763 212
rect -1735 184 -1697 212
rect -1669 184 -1631 212
rect -1603 184 -1565 212
rect -1537 184 -1499 212
rect -1471 184 -1433 212
rect -1405 184 -1367 212
rect -1339 184 -1301 212
rect -1273 184 -1235 212
rect -1207 184 -1169 212
rect -1141 184 -1103 212
rect -1075 184 -1037 212
rect -1009 184 -971 212
rect -943 184 -905 212
rect -877 184 -839 212
rect -811 184 -773 212
rect -745 184 -707 212
rect -679 184 -641 212
rect -613 184 -575 212
rect -547 184 -509 212
rect -481 184 -443 212
rect -415 184 -377 212
rect -349 184 -311 212
rect -283 184 -245 212
rect -217 184 -179 212
rect -151 184 -113 212
rect -85 184 -47 212
rect -19 184 19 212
rect 47 184 85 212
rect 113 184 151 212
rect 179 184 217 212
rect 245 184 283 212
rect 311 184 349 212
rect 377 184 415 212
rect 443 184 481 212
rect 509 184 547 212
rect 575 184 613 212
rect 641 184 679 212
rect 707 184 745 212
rect 773 184 811 212
rect 839 184 877 212
rect 905 184 943 212
rect 971 184 1009 212
rect 1037 184 1075 212
rect 1103 184 1141 212
rect 1169 184 1207 212
rect 1235 184 1273 212
rect 1301 184 1339 212
rect 1367 184 1405 212
rect 1433 184 1471 212
rect 1499 184 1537 212
rect 1565 184 1603 212
rect 1631 184 1669 212
rect 1697 184 1735 212
rect 1763 184 1801 212
rect 1829 184 1867 212
rect 1895 184 1933 212
rect 1961 184 1999 212
rect 2027 184 2065 212
rect 2093 184 2131 212
rect 2159 184 2197 212
rect 2225 184 2230 212
rect -2230 146 2230 184
rect -2230 118 -2225 146
rect -2197 118 -2159 146
rect -2131 118 -2093 146
rect -2065 118 -2027 146
rect -1999 118 -1961 146
rect -1933 118 -1895 146
rect -1867 118 -1829 146
rect -1801 118 -1763 146
rect -1735 118 -1697 146
rect -1669 118 -1631 146
rect -1603 118 -1565 146
rect -1537 118 -1499 146
rect -1471 118 -1433 146
rect -1405 118 -1367 146
rect -1339 118 -1301 146
rect -1273 118 -1235 146
rect -1207 118 -1169 146
rect -1141 118 -1103 146
rect -1075 118 -1037 146
rect -1009 118 -971 146
rect -943 118 -905 146
rect -877 118 -839 146
rect -811 118 -773 146
rect -745 118 -707 146
rect -679 118 -641 146
rect -613 118 -575 146
rect -547 118 -509 146
rect -481 118 -443 146
rect -415 118 -377 146
rect -349 118 -311 146
rect -283 118 -245 146
rect -217 118 -179 146
rect -151 118 -113 146
rect -85 118 -47 146
rect -19 118 19 146
rect 47 118 85 146
rect 113 118 151 146
rect 179 118 217 146
rect 245 118 283 146
rect 311 118 349 146
rect 377 118 415 146
rect 443 118 481 146
rect 509 118 547 146
rect 575 118 613 146
rect 641 118 679 146
rect 707 118 745 146
rect 773 118 811 146
rect 839 118 877 146
rect 905 118 943 146
rect 971 118 1009 146
rect 1037 118 1075 146
rect 1103 118 1141 146
rect 1169 118 1207 146
rect 1235 118 1273 146
rect 1301 118 1339 146
rect 1367 118 1405 146
rect 1433 118 1471 146
rect 1499 118 1537 146
rect 1565 118 1603 146
rect 1631 118 1669 146
rect 1697 118 1735 146
rect 1763 118 1801 146
rect 1829 118 1867 146
rect 1895 118 1933 146
rect 1961 118 1999 146
rect 2027 118 2065 146
rect 2093 118 2131 146
rect 2159 118 2197 146
rect 2225 118 2230 146
rect -2230 80 2230 118
rect -2230 52 -2225 80
rect -2197 52 -2159 80
rect -2131 52 -2093 80
rect -2065 52 -2027 80
rect -1999 52 -1961 80
rect -1933 52 -1895 80
rect -1867 52 -1829 80
rect -1801 52 -1763 80
rect -1735 52 -1697 80
rect -1669 52 -1631 80
rect -1603 52 -1565 80
rect -1537 52 -1499 80
rect -1471 52 -1433 80
rect -1405 52 -1367 80
rect -1339 52 -1301 80
rect -1273 52 -1235 80
rect -1207 52 -1169 80
rect -1141 52 -1103 80
rect -1075 52 -1037 80
rect -1009 52 -971 80
rect -943 52 -905 80
rect -877 52 -839 80
rect -811 52 -773 80
rect -745 52 -707 80
rect -679 52 -641 80
rect -613 52 -575 80
rect -547 52 -509 80
rect -481 52 -443 80
rect -415 52 -377 80
rect -349 52 -311 80
rect -283 52 -245 80
rect -217 52 -179 80
rect -151 52 -113 80
rect -85 52 -47 80
rect -19 52 19 80
rect 47 52 85 80
rect 113 52 151 80
rect 179 52 217 80
rect 245 52 283 80
rect 311 52 349 80
rect 377 52 415 80
rect 443 52 481 80
rect 509 52 547 80
rect 575 52 613 80
rect 641 52 679 80
rect 707 52 745 80
rect 773 52 811 80
rect 839 52 877 80
rect 905 52 943 80
rect 971 52 1009 80
rect 1037 52 1075 80
rect 1103 52 1141 80
rect 1169 52 1207 80
rect 1235 52 1273 80
rect 1301 52 1339 80
rect 1367 52 1405 80
rect 1433 52 1471 80
rect 1499 52 1537 80
rect 1565 52 1603 80
rect 1631 52 1669 80
rect 1697 52 1735 80
rect 1763 52 1801 80
rect 1829 52 1867 80
rect 1895 52 1933 80
rect 1961 52 1999 80
rect 2027 52 2065 80
rect 2093 52 2131 80
rect 2159 52 2197 80
rect 2225 52 2230 80
rect -2230 14 2230 52
rect -2230 -14 -2225 14
rect -2197 -14 -2159 14
rect -2131 -14 -2093 14
rect -2065 -14 -2027 14
rect -1999 -14 -1961 14
rect -1933 -14 -1895 14
rect -1867 -14 -1829 14
rect -1801 -14 -1763 14
rect -1735 -14 -1697 14
rect -1669 -14 -1631 14
rect -1603 -14 -1565 14
rect -1537 -14 -1499 14
rect -1471 -14 -1433 14
rect -1405 -14 -1367 14
rect -1339 -14 -1301 14
rect -1273 -14 -1235 14
rect -1207 -14 -1169 14
rect -1141 -14 -1103 14
rect -1075 -14 -1037 14
rect -1009 -14 -971 14
rect -943 -14 -905 14
rect -877 -14 -839 14
rect -811 -14 -773 14
rect -745 -14 -707 14
rect -679 -14 -641 14
rect -613 -14 -575 14
rect -547 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 19 14
rect 47 -14 85 14
rect 113 -14 151 14
rect 179 -14 217 14
rect 245 -14 283 14
rect 311 -14 349 14
rect 377 -14 415 14
rect 443 -14 481 14
rect 509 -14 547 14
rect 575 -14 613 14
rect 641 -14 679 14
rect 707 -14 745 14
rect 773 -14 811 14
rect 839 -14 877 14
rect 905 -14 943 14
rect 971 -14 1009 14
rect 1037 -14 1075 14
rect 1103 -14 1141 14
rect 1169 -14 1207 14
rect 1235 -14 1273 14
rect 1301 -14 1339 14
rect 1367 -14 1405 14
rect 1433 -14 1471 14
rect 1499 -14 1537 14
rect 1565 -14 1603 14
rect 1631 -14 1669 14
rect 1697 -14 1735 14
rect 1763 -14 1801 14
rect 1829 -14 1867 14
rect 1895 -14 1933 14
rect 1961 -14 1999 14
rect 2027 -14 2065 14
rect 2093 -14 2131 14
rect 2159 -14 2197 14
rect 2225 -14 2230 14
rect -2230 -52 2230 -14
rect -2230 -80 -2225 -52
rect -2197 -80 -2159 -52
rect -2131 -80 -2093 -52
rect -2065 -80 -2027 -52
rect -1999 -80 -1961 -52
rect -1933 -80 -1895 -52
rect -1867 -80 -1829 -52
rect -1801 -80 -1763 -52
rect -1735 -80 -1697 -52
rect -1669 -80 -1631 -52
rect -1603 -80 -1565 -52
rect -1537 -80 -1499 -52
rect -1471 -80 -1433 -52
rect -1405 -80 -1367 -52
rect -1339 -80 -1301 -52
rect -1273 -80 -1235 -52
rect -1207 -80 -1169 -52
rect -1141 -80 -1103 -52
rect -1075 -80 -1037 -52
rect -1009 -80 -971 -52
rect -943 -80 -905 -52
rect -877 -80 -839 -52
rect -811 -80 -773 -52
rect -745 -80 -707 -52
rect -679 -80 -641 -52
rect -613 -80 -575 -52
rect -547 -80 -509 -52
rect -481 -80 -443 -52
rect -415 -80 -377 -52
rect -349 -80 -311 -52
rect -283 -80 -245 -52
rect -217 -80 -179 -52
rect -151 -80 -113 -52
rect -85 -80 -47 -52
rect -19 -80 19 -52
rect 47 -80 85 -52
rect 113 -80 151 -52
rect 179 -80 217 -52
rect 245 -80 283 -52
rect 311 -80 349 -52
rect 377 -80 415 -52
rect 443 -80 481 -52
rect 509 -80 547 -52
rect 575 -80 613 -52
rect 641 -80 679 -52
rect 707 -80 745 -52
rect 773 -80 811 -52
rect 839 -80 877 -52
rect 905 -80 943 -52
rect 971 -80 1009 -52
rect 1037 -80 1075 -52
rect 1103 -80 1141 -52
rect 1169 -80 1207 -52
rect 1235 -80 1273 -52
rect 1301 -80 1339 -52
rect 1367 -80 1405 -52
rect 1433 -80 1471 -52
rect 1499 -80 1537 -52
rect 1565 -80 1603 -52
rect 1631 -80 1669 -52
rect 1697 -80 1735 -52
rect 1763 -80 1801 -52
rect 1829 -80 1867 -52
rect 1895 -80 1933 -52
rect 1961 -80 1999 -52
rect 2027 -80 2065 -52
rect 2093 -80 2131 -52
rect 2159 -80 2197 -52
rect 2225 -80 2230 -52
rect -2230 -118 2230 -80
rect -2230 -146 -2225 -118
rect -2197 -146 -2159 -118
rect -2131 -146 -2093 -118
rect -2065 -146 -2027 -118
rect -1999 -146 -1961 -118
rect -1933 -146 -1895 -118
rect -1867 -146 -1829 -118
rect -1801 -146 -1763 -118
rect -1735 -146 -1697 -118
rect -1669 -146 -1631 -118
rect -1603 -146 -1565 -118
rect -1537 -146 -1499 -118
rect -1471 -146 -1433 -118
rect -1405 -146 -1367 -118
rect -1339 -146 -1301 -118
rect -1273 -146 -1235 -118
rect -1207 -146 -1169 -118
rect -1141 -146 -1103 -118
rect -1075 -146 -1037 -118
rect -1009 -146 -971 -118
rect -943 -146 -905 -118
rect -877 -146 -839 -118
rect -811 -146 -773 -118
rect -745 -146 -707 -118
rect -679 -146 -641 -118
rect -613 -146 -575 -118
rect -547 -146 -509 -118
rect -481 -146 -443 -118
rect -415 -146 -377 -118
rect -349 -146 -311 -118
rect -283 -146 -245 -118
rect -217 -146 -179 -118
rect -151 -146 -113 -118
rect -85 -146 -47 -118
rect -19 -146 19 -118
rect 47 -146 85 -118
rect 113 -146 151 -118
rect 179 -146 217 -118
rect 245 -146 283 -118
rect 311 -146 349 -118
rect 377 -146 415 -118
rect 443 -146 481 -118
rect 509 -146 547 -118
rect 575 -146 613 -118
rect 641 -146 679 -118
rect 707 -146 745 -118
rect 773 -146 811 -118
rect 839 -146 877 -118
rect 905 -146 943 -118
rect 971 -146 1009 -118
rect 1037 -146 1075 -118
rect 1103 -146 1141 -118
rect 1169 -146 1207 -118
rect 1235 -146 1273 -118
rect 1301 -146 1339 -118
rect 1367 -146 1405 -118
rect 1433 -146 1471 -118
rect 1499 -146 1537 -118
rect 1565 -146 1603 -118
rect 1631 -146 1669 -118
rect 1697 -146 1735 -118
rect 1763 -146 1801 -118
rect 1829 -146 1867 -118
rect 1895 -146 1933 -118
rect 1961 -146 1999 -118
rect 2027 -146 2065 -118
rect 2093 -146 2131 -118
rect 2159 -146 2197 -118
rect 2225 -146 2230 -118
rect -2230 -184 2230 -146
rect -2230 -212 -2225 -184
rect -2197 -212 -2159 -184
rect -2131 -212 -2093 -184
rect -2065 -212 -2027 -184
rect -1999 -212 -1961 -184
rect -1933 -212 -1895 -184
rect -1867 -212 -1829 -184
rect -1801 -212 -1763 -184
rect -1735 -212 -1697 -184
rect -1669 -212 -1631 -184
rect -1603 -212 -1565 -184
rect -1537 -212 -1499 -184
rect -1471 -212 -1433 -184
rect -1405 -212 -1367 -184
rect -1339 -212 -1301 -184
rect -1273 -212 -1235 -184
rect -1207 -212 -1169 -184
rect -1141 -212 -1103 -184
rect -1075 -212 -1037 -184
rect -1009 -212 -971 -184
rect -943 -212 -905 -184
rect -877 -212 -839 -184
rect -811 -212 -773 -184
rect -745 -212 -707 -184
rect -679 -212 -641 -184
rect -613 -212 -575 -184
rect -547 -212 -509 -184
rect -481 -212 -443 -184
rect -415 -212 -377 -184
rect -349 -212 -311 -184
rect -283 -212 -245 -184
rect -217 -212 -179 -184
rect -151 -212 -113 -184
rect -85 -212 -47 -184
rect -19 -212 19 -184
rect 47 -212 85 -184
rect 113 -212 151 -184
rect 179 -212 217 -184
rect 245 -212 283 -184
rect 311 -212 349 -184
rect 377 -212 415 -184
rect 443 -212 481 -184
rect 509 -212 547 -184
rect 575 -212 613 -184
rect 641 -212 679 -184
rect 707 -212 745 -184
rect 773 -212 811 -184
rect 839 -212 877 -184
rect 905 -212 943 -184
rect 971 -212 1009 -184
rect 1037 -212 1075 -184
rect 1103 -212 1141 -184
rect 1169 -212 1207 -184
rect 1235 -212 1273 -184
rect 1301 -212 1339 -184
rect 1367 -212 1405 -184
rect 1433 -212 1471 -184
rect 1499 -212 1537 -184
rect 1565 -212 1603 -184
rect 1631 -212 1669 -184
rect 1697 -212 1735 -184
rect 1763 -212 1801 -184
rect 1829 -212 1867 -184
rect 1895 -212 1933 -184
rect 1961 -212 1999 -184
rect 2027 -212 2065 -184
rect 2093 -212 2131 -184
rect 2159 -212 2197 -184
rect 2225 -212 2230 -184
rect -2230 -250 2230 -212
rect -2230 -278 -2225 -250
rect -2197 -278 -2159 -250
rect -2131 -278 -2093 -250
rect -2065 -278 -2027 -250
rect -1999 -278 -1961 -250
rect -1933 -278 -1895 -250
rect -1867 -278 -1829 -250
rect -1801 -278 -1763 -250
rect -1735 -278 -1697 -250
rect -1669 -278 -1631 -250
rect -1603 -278 -1565 -250
rect -1537 -278 -1499 -250
rect -1471 -278 -1433 -250
rect -1405 -278 -1367 -250
rect -1339 -278 -1301 -250
rect -1273 -278 -1235 -250
rect -1207 -278 -1169 -250
rect -1141 -278 -1103 -250
rect -1075 -278 -1037 -250
rect -1009 -278 -971 -250
rect -943 -278 -905 -250
rect -877 -278 -839 -250
rect -811 -278 -773 -250
rect -745 -278 -707 -250
rect -679 -278 -641 -250
rect -613 -278 -575 -250
rect -547 -278 -509 -250
rect -481 -278 -443 -250
rect -415 -278 -377 -250
rect -349 -278 -311 -250
rect -283 -278 -245 -250
rect -217 -278 -179 -250
rect -151 -278 -113 -250
rect -85 -278 -47 -250
rect -19 -278 19 -250
rect 47 -278 85 -250
rect 113 -278 151 -250
rect 179 -278 217 -250
rect 245 -278 283 -250
rect 311 -278 349 -250
rect 377 -278 415 -250
rect 443 -278 481 -250
rect 509 -278 547 -250
rect 575 -278 613 -250
rect 641 -278 679 -250
rect 707 -278 745 -250
rect 773 -278 811 -250
rect 839 -278 877 -250
rect 905 -278 943 -250
rect 971 -278 1009 -250
rect 1037 -278 1075 -250
rect 1103 -278 1141 -250
rect 1169 -278 1207 -250
rect 1235 -278 1273 -250
rect 1301 -278 1339 -250
rect 1367 -278 1405 -250
rect 1433 -278 1471 -250
rect 1499 -278 1537 -250
rect 1565 -278 1603 -250
rect 1631 -278 1669 -250
rect 1697 -278 1735 -250
rect 1763 -278 1801 -250
rect 1829 -278 1867 -250
rect 1895 -278 1933 -250
rect 1961 -278 1999 -250
rect 2027 -278 2065 -250
rect 2093 -278 2131 -250
rect 2159 -278 2197 -250
rect 2225 -278 2230 -250
rect -2230 -316 2230 -278
rect -2230 -344 -2225 -316
rect -2197 -344 -2159 -316
rect -2131 -344 -2093 -316
rect -2065 -344 -2027 -316
rect -1999 -344 -1961 -316
rect -1933 -344 -1895 -316
rect -1867 -344 -1829 -316
rect -1801 -344 -1763 -316
rect -1735 -344 -1697 -316
rect -1669 -344 -1631 -316
rect -1603 -344 -1565 -316
rect -1537 -344 -1499 -316
rect -1471 -344 -1433 -316
rect -1405 -344 -1367 -316
rect -1339 -344 -1301 -316
rect -1273 -344 -1235 -316
rect -1207 -344 -1169 -316
rect -1141 -344 -1103 -316
rect -1075 -344 -1037 -316
rect -1009 -344 -971 -316
rect -943 -344 -905 -316
rect -877 -344 -839 -316
rect -811 -344 -773 -316
rect -745 -344 -707 -316
rect -679 -344 -641 -316
rect -613 -344 -575 -316
rect -547 -344 -509 -316
rect -481 -344 -443 -316
rect -415 -344 -377 -316
rect -349 -344 -311 -316
rect -283 -344 -245 -316
rect -217 -344 -179 -316
rect -151 -344 -113 -316
rect -85 -344 -47 -316
rect -19 -344 19 -316
rect 47 -344 85 -316
rect 113 -344 151 -316
rect 179 -344 217 -316
rect 245 -344 283 -316
rect 311 -344 349 -316
rect 377 -344 415 -316
rect 443 -344 481 -316
rect 509 -344 547 -316
rect 575 -344 613 -316
rect 641 -344 679 -316
rect 707 -344 745 -316
rect 773 -344 811 -316
rect 839 -344 877 -316
rect 905 -344 943 -316
rect 971 -344 1009 -316
rect 1037 -344 1075 -316
rect 1103 -344 1141 -316
rect 1169 -344 1207 -316
rect 1235 -344 1273 -316
rect 1301 -344 1339 -316
rect 1367 -344 1405 -316
rect 1433 -344 1471 -316
rect 1499 -344 1537 -316
rect 1565 -344 1603 -316
rect 1631 -344 1669 -316
rect 1697 -344 1735 -316
rect 1763 -344 1801 -316
rect 1829 -344 1867 -316
rect 1895 -344 1933 -316
rect 1961 -344 1999 -316
rect 2027 -344 2065 -316
rect 2093 -344 2131 -316
rect 2159 -344 2197 -316
rect 2225 -344 2230 -316
rect -2230 -349 2230 -344
<< via3 >>
rect -2225 316 -2197 344
rect -2159 316 -2131 344
rect -2093 316 -2065 344
rect -2027 316 -1999 344
rect -1961 316 -1933 344
rect -1895 316 -1867 344
rect -1829 316 -1801 344
rect -1763 316 -1735 344
rect -1697 316 -1669 344
rect -1631 316 -1603 344
rect -1565 316 -1537 344
rect -1499 316 -1471 344
rect -1433 316 -1405 344
rect -1367 316 -1339 344
rect -1301 316 -1273 344
rect -1235 316 -1207 344
rect -1169 316 -1141 344
rect -1103 316 -1075 344
rect -1037 316 -1009 344
rect -971 316 -943 344
rect -905 316 -877 344
rect -839 316 -811 344
rect -773 316 -745 344
rect -707 316 -679 344
rect -641 316 -613 344
rect -575 316 -547 344
rect -509 316 -481 344
rect -443 316 -415 344
rect -377 316 -349 344
rect -311 316 -283 344
rect -245 316 -217 344
rect -179 316 -151 344
rect -113 316 -85 344
rect -47 316 -19 344
rect 19 316 47 344
rect 85 316 113 344
rect 151 316 179 344
rect 217 316 245 344
rect 283 316 311 344
rect 349 316 377 344
rect 415 316 443 344
rect 481 316 509 344
rect 547 316 575 344
rect 613 316 641 344
rect 679 316 707 344
rect 745 316 773 344
rect 811 316 839 344
rect 877 316 905 344
rect 943 316 971 344
rect 1009 316 1037 344
rect 1075 316 1103 344
rect 1141 316 1169 344
rect 1207 316 1235 344
rect 1273 316 1301 344
rect 1339 316 1367 344
rect 1405 316 1433 344
rect 1471 316 1499 344
rect 1537 316 1565 344
rect 1603 316 1631 344
rect 1669 316 1697 344
rect 1735 316 1763 344
rect 1801 316 1829 344
rect 1867 316 1895 344
rect 1933 316 1961 344
rect 1999 316 2027 344
rect 2065 316 2093 344
rect 2131 316 2159 344
rect 2197 316 2225 344
rect -2225 250 -2197 278
rect -2159 250 -2131 278
rect -2093 250 -2065 278
rect -2027 250 -1999 278
rect -1961 250 -1933 278
rect -1895 250 -1867 278
rect -1829 250 -1801 278
rect -1763 250 -1735 278
rect -1697 250 -1669 278
rect -1631 250 -1603 278
rect -1565 250 -1537 278
rect -1499 250 -1471 278
rect -1433 250 -1405 278
rect -1367 250 -1339 278
rect -1301 250 -1273 278
rect -1235 250 -1207 278
rect -1169 250 -1141 278
rect -1103 250 -1075 278
rect -1037 250 -1009 278
rect -971 250 -943 278
rect -905 250 -877 278
rect -839 250 -811 278
rect -773 250 -745 278
rect -707 250 -679 278
rect -641 250 -613 278
rect -575 250 -547 278
rect -509 250 -481 278
rect -443 250 -415 278
rect -377 250 -349 278
rect -311 250 -283 278
rect -245 250 -217 278
rect -179 250 -151 278
rect -113 250 -85 278
rect -47 250 -19 278
rect 19 250 47 278
rect 85 250 113 278
rect 151 250 179 278
rect 217 250 245 278
rect 283 250 311 278
rect 349 250 377 278
rect 415 250 443 278
rect 481 250 509 278
rect 547 250 575 278
rect 613 250 641 278
rect 679 250 707 278
rect 745 250 773 278
rect 811 250 839 278
rect 877 250 905 278
rect 943 250 971 278
rect 1009 250 1037 278
rect 1075 250 1103 278
rect 1141 250 1169 278
rect 1207 250 1235 278
rect 1273 250 1301 278
rect 1339 250 1367 278
rect 1405 250 1433 278
rect 1471 250 1499 278
rect 1537 250 1565 278
rect 1603 250 1631 278
rect 1669 250 1697 278
rect 1735 250 1763 278
rect 1801 250 1829 278
rect 1867 250 1895 278
rect 1933 250 1961 278
rect 1999 250 2027 278
rect 2065 250 2093 278
rect 2131 250 2159 278
rect 2197 250 2225 278
rect -2225 184 -2197 212
rect -2159 184 -2131 212
rect -2093 184 -2065 212
rect -2027 184 -1999 212
rect -1961 184 -1933 212
rect -1895 184 -1867 212
rect -1829 184 -1801 212
rect -1763 184 -1735 212
rect -1697 184 -1669 212
rect -1631 184 -1603 212
rect -1565 184 -1537 212
rect -1499 184 -1471 212
rect -1433 184 -1405 212
rect -1367 184 -1339 212
rect -1301 184 -1273 212
rect -1235 184 -1207 212
rect -1169 184 -1141 212
rect -1103 184 -1075 212
rect -1037 184 -1009 212
rect -971 184 -943 212
rect -905 184 -877 212
rect -839 184 -811 212
rect -773 184 -745 212
rect -707 184 -679 212
rect -641 184 -613 212
rect -575 184 -547 212
rect -509 184 -481 212
rect -443 184 -415 212
rect -377 184 -349 212
rect -311 184 -283 212
rect -245 184 -217 212
rect -179 184 -151 212
rect -113 184 -85 212
rect -47 184 -19 212
rect 19 184 47 212
rect 85 184 113 212
rect 151 184 179 212
rect 217 184 245 212
rect 283 184 311 212
rect 349 184 377 212
rect 415 184 443 212
rect 481 184 509 212
rect 547 184 575 212
rect 613 184 641 212
rect 679 184 707 212
rect 745 184 773 212
rect 811 184 839 212
rect 877 184 905 212
rect 943 184 971 212
rect 1009 184 1037 212
rect 1075 184 1103 212
rect 1141 184 1169 212
rect 1207 184 1235 212
rect 1273 184 1301 212
rect 1339 184 1367 212
rect 1405 184 1433 212
rect 1471 184 1499 212
rect 1537 184 1565 212
rect 1603 184 1631 212
rect 1669 184 1697 212
rect 1735 184 1763 212
rect 1801 184 1829 212
rect 1867 184 1895 212
rect 1933 184 1961 212
rect 1999 184 2027 212
rect 2065 184 2093 212
rect 2131 184 2159 212
rect 2197 184 2225 212
rect -2225 118 -2197 146
rect -2159 118 -2131 146
rect -2093 118 -2065 146
rect -2027 118 -1999 146
rect -1961 118 -1933 146
rect -1895 118 -1867 146
rect -1829 118 -1801 146
rect -1763 118 -1735 146
rect -1697 118 -1669 146
rect -1631 118 -1603 146
rect -1565 118 -1537 146
rect -1499 118 -1471 146
rect -1433 118 -1405 146
rect -1367 118 -1339 146
rect -1301 118 -1273 146
rect -1235 118 -1207 146
rect -1169 118 -1141 146
rect -1103 118 -1075 146
rect -1037 118 -1009 146
rect -971 118 -943 146
rect -905 118 -877 146
rect -839 118 -811 146
rect -773 118 -745 146
rect -707 118 -679 146
rect -641 118 -613 146
rect -575 118 -547 146
rect -509 118 -481 146
rect -443 118 -415 146
rect -377 118 -349 146
rect -311 118 -283 146
rect -245 118 -217 146
rect -179 118 -151 146
rect -113 118 -85 146
rect -47 118 -19 146
rect 19 118 47 146
rect 85 118 113 146
rect 151 118 179 146
rect 217 118 245 146
rect 283 118 311 146
rect 349 118 377 146
rect 415 118 443 146
rect 481 118 509 146
rect 547 118 575 146
rect 613 118 641 146
rect 679 118 707 146
rect 745 118 773 146
rect 811 118 839 146
rect 877 118 905 146
rect 943 118 971 146
rect 1009 118 1037 146
rect 1075 118 1103 146
rect 1141 118 1169 146
rect 1207 118 1235 146
rect 1273 118 1301 146
rect 1339 118 1367 146
rect 1405 118 1433 146
rect 1471 118 1499 146
rect 1537 118 1565 146
rect 1603 118 1631 146
rect 1669 118 1697 146
rect 1735 118 1763 146
rect 1801 118 1829 146
rect 1867 118 1895 146
rect 1933 118 1961 146
rect 1999 118 2027 146
rect 2065 118 2093 146
rect 2131 118 2159 146
rect 2197 118 2225 146
rect -2225 52 -2197 80
rect -2159 52 -2131 80
rect -2093 52 -2065 80
rect -2027 52 -1999 80
rect -1961 52 -1933 80
rect -1895 52 -1867 80
rect -1829 52 -1801 80
rect -1763 52 -1735 80
rect -1697 52 -1669 80
rect -1631 52 -1603 80
rect -1565 52 -1537 80
rect -1499 52 -1471 80
rect -1433 52 -1405 80
rect -1367 52 -1339 80
rect -1301 52 -1273 80
rect -1235 52 -1207 80
rect -1169 52 -1141 80
rect -1103 52 -1075 80
rect -1037 52 -1009 80
rect -971 52 -943 80
rect -905 52 -877 80
rect -839 52 -811 80
rect -773 52 -745 80
rect -707 52 -679 80
rect -641 52 -613 80
rect -575 52 -547 80
rect -509 52 -481 80
rect -443 52 -415 80
rect -377 52 -349 80
rect -311 52 -283 80
rect -245 52 -217 80
rect -179 52 -151 80
rect -113 52 -85 80
rect -47 52 -19 80
rect 19 52 47 80
rect 85 52 113 80
rect 151 52 179 80
rect 217 52 245 80
rect 283 52 311 80
rect 349 52 377 80
rect 415 52 443 80
rect 481 52 509 80
rect 547 52 575 80
rect 613 52 641 80
rect 679 52 707 80
rect 745 52 773 80
rect 811 52 839 80
rect 877 52 905 80
rect 943 52 971 80
rect 1009 52 1037 80
rect 1075 52 1103 80
rect 1141 52 1169 80
rect 1207 52 1235 80
rect 1273 52 1301 80
rect 1339 52 1367 80
rect 1405 52 1433 80
rect 1471 52 1499 80
rect 1537 52 1565 80
rect 1603 52 1631 80
rect 1669 52 1697 80
rect 1735 52 1763 80
rect 1801 52 1829 80
rect 1867 52 1895 80
rect 1933 52 1961 80
rect 1999 52 2027 80
rect 2065 52 2093 80
rect 2131 52 2159 80
rect 2197 52 2225 80
rect -2225 -14 -2197 14
rect -2159 -14 -2131 14
rect -2093 -14 -2065 14
rect -2027 -14 -1999 14
rect -1961 -14 -1933 14
rect -1895 -14 -1867 14
rect -1829 -14 -1801 14
rect -1763 -14 -1735 14
rect -1697 -14 -1669 14
rect -1631 -14 -1603 14
rect -1565 -14 -1537 14
rect -1499 -14 -1471 14
rect -1433 -14 -1405 14
rect -1367 -14 -1339 14
rect -1301 -14 -1273 14
rect -1235 -14 -1207 14
rect -1169 -14 -1141 14
rect -1103 -14 -1075 14
rect -1037 -14 -1009 14
rect -971 -14 -943 14
rect -905 -14 -877 14
rect -839 -14 -811 14
rect -773 -14 -745 14
rect -707 -14 -679 14
rect -641 -14 -613 14
rect -575 -14 -547 14
rect -509 -14 -481 14
rect -443 -14 -415 14
rect -377 -14 -349 14
rect -311 -14 -283 14
rect -245 -14 -217 14
rect -179 -14 -151 14
rect -113 -14 -85 14
rect -47 -14 -19 14
rect 19 -14 47 14
rect 85 -14 113 14
rect 151 -14 179 14
rect 217 -14 245 14
rect 283 -14 311 14
rect 349 -14 377 14
rect 415 -14 443 14
rect 481 -14 509 14
rect 547 -14 575 14
rect 613 -14 641 14
rect 679 -14 707 14
rect 745 -14 773 14
rect 811 -14 839 14
rect 877 -14 905 14
rect 943 -14 971 14
rect 1009 -14 1037 14
rect 1075 -14 1103 14
rect 1141 -14 1169 14
rect 1207 -14 1235 14
rect 1273 -14 1301 14
rect 1339 -14 1367 14
rect 1405 -14 1433 14
rect 1471 -14 1499 14
rect 1537 -14 1565 14
rect 1603 -14 1631 14
rect 1669 -14 1697 14
rect 1735 -14 1763 14
rect 1801 -14 1829 14
rect 1867 -14 1895 14
rect 1933 -14 1961 14
rect 1999 -14 2027 14
rect 2065 -14 2093 14
rect 2131 -14 2159 14
rect 2197 -14 2225 14
rect -2225 -80 -2197 -52
rect -2159 -80 -2131 -52
rect -2093 -80 -2065 -52
rect -2027 -80 -1999 -52
rect -1961 -80 -1933 -52
rect -1895 -80 -1867 -52
rect -1829 -80 -1801 -52
rect -1763 -80 -1735 -52
rect -1697 -80 -1669 -52
rect -1631 -80 -1603 -52
rect -1565 -80 -1537 -52
rect -1499 -80 -1471 -52
rect -1433 -80 -1405 -52
rect -1367 -80 -1339 -52
rect -1301 -80 -1273 -52
rect -1235 -80 -1207 -52
rect -1169 -80 -1141 -52
rect -1103 -80 -1075 -52
rect -1037 -80 -1009 -52
rect -971 -80 -943 -52
rect -905 -80 -877 -52
rect -839 -80 -811 -52
rect -773 -80 -745 -52
rect -707 -80 -679 -52
rect -641 -80 -613 -52
rect -575 -80 -547 -52
rect -509 -80 -481 -52
rect -443 -80 -415 -52
rect -377 -80 -349 -52
rect -311 -80 -283 -52
rect -245 -80 -217 -52
rect -179 -80 -151 -52
rect -113 -80 -85 -52
rect -47 -80 -19 -52
rect 19 -80 47 -52
rect 85 -80 113 -52
rect 151 -80 179 -52
rect 217 -80 245 -52
rect 283 -80 311 -52
rect 349 -80 377 -52
rect 415 -80 443 -52
rect 481 -80 509 -52
rect 547 -80 575 -52
rect 613 -80 641 -52
rect 679 -80 707 -52
rect 745 -80 773 -52
rect 811 -80 839 -52
rect 877 -80 905 -52
rect 943 -80 971 -52
rect 1009 -80 1037 -52
rect 1075 -80 1103 -52
rect 1141 -80 1169 -52
rect 1207 -80 1235 -52
rect 1273 -80 1301 -52
rect 1339 -80 1367 -52
rect 1405 -80 1433 -52
rect 1471 -80 1499 -52
rect 1537 -80 1565 -52
rect 1603 -80 1631 -52
rect 1669 -80 1697 -52
rect 1735 -80 1763 -52
rect 1801 -80 1829 -52
rect 1867 -80 1895 -52
rect 1933 -80 1961 -52
rect 1999 -80 2027 -52
rect 2065 -80 2093 -52
rect 2131 -80 2159 -52
rect 2197 -80 2225 -52
rect -2225 -146 -2197 -118
rect -2159 -146 -2131 -118
rect -2093 -146 -2065 -118
rect -2027 -146 -1999 -118
rect -1961 -146 -1933 -118
rect -1895 -146 -1867 -118
rect -1829 -146 -1801 -118
rect -1763 -146 -1735 -118
rect -1697 -146 -1669 -118
rect -1631 -146 -1603 -118
rect -1565 -146 -1537 -118
rect -1499 -146 -1471 -118
rect -1433 -146 -1405 -118
rect -1367 -146 -1339 -118
rect -1301 -146 -1273 -118
rect -1235 -146 -1207 -118
rect -1169 -146 -1141 -118
rect -1103 -146 -1075 -118
rect -1037 -146 -1009 -118
rect -971 -146 -943 -118
rect -905 -146 -877 -118
rect -839 -146 -811 -118
rect -773 -146 -745 -118
rect -707 -146 -679 -118
rect -641 -146 -613 -118
rect -575 -146 -547 -118
rect -509 -146 -481 -118
rect -443 -146 -415 -118
rect -377 -146 -349 -118
rect -311 -146 -283 -118
rect -245 -146 -217 -118
rect -179 -146 -151 -118
rect -113 -146 -85 -118
rect -47 -146 -19 -118
rect 19 -146 47 -118
rect 85 -146 113 -118
rect 151 -146 179 -118
rect 217 -146 245 -118
rect 283 -146 311 -118
rect 349 -146 377 -118
rect 415 -146 443 -118
rect 481 -146 509 -118
rect 547 -146 575 -118
rect 613 -146 641 -118
rect 679 -146 707 -118
rect 745 -146 773 -118
rect 811 -146 839 -118
rect 877 -146 905 -118
rect 943 -146 971 -118
rect 1009 -146 1037 -118
rect 1075 -146 1103 -118
rect 1141 -146 1169 -118
rect 1207 -146 1235 -118
rect 1273 -146 1301 -118
rect 1339 -146 1367 -118
rect 1405 -146 1433 -118
rect 1471 -146 1499 -118
rect 1537 -146 1565 -118
rect 1603 -146 1631 -118
rect 1669 -146 1697 -118
rect 1735 -146 1763 -118
rect 1801 -146 1829 -118
rect 1867 -146 1895 -118
rect 1933 -146 1961 -118
rect 1999 -146 2027 -118
rect 2065 -146 2093 -118
rect 2131 -146 2159 -118
rect 2197 -146 2225 -118
rect -2225 -212 -2197 -184
rect -2159 -212 -2131 -184
rect -2093 -212 -2065 -184
rect -2027 -212 -1999 -184
rect -1961 -212 -1933 -184
rect -1895 -212 -1867 -184
rect -1829 -212 -1801 -184
rect -1763 -212 -1735 -184
rect -1697 -212 -1669 -184
rect -1631 -212 -1603 -184
rect -1565 -212 -1537 -184
rect -1499 -212 -1471 -184
rect -1433 -212 -1405 -184
rect -1367 -212 -1339 -184
rect -1301 -212 -1273 -184
rect -1235 -212 -1207 -184
rect -1169 -212 -1141 -184
rect -1103 -212 -1075 -184
rect -1037 -212 -1009 -184
rect -971 -212 -943 -184
rect -905 -212 -877 -184
rect -839 -212 -811 -184
rect -773 -212 -745 -184
rect -707 -212 -679 -184
rect -641 -212 -613 -184
rect -575 -212 -547 -184
rect -509 -212 -481 -184
rect -443 -212 -415 -184
rect -377 -212 -349 -184
rect -311 -212 -283 -184
rect -245 -212 -217 -184
rect -179 -212 -151 -184
rect -113 -212 -85 -184
rect -47 -212 -19 -184
rect 19 -212 47 -184
rect 85 -212 113 -184
rect 151 -212 179 -184
rect 217 -212 245 -184
rect 283 -212 311 -184
rect 349 -212 377 -184
rect 415 -212 443 -184
rect 481 -212 509 -184
rect 547 -212 575 -184
rect 613 -212 641 -184
rect 679 -212 707 -184
rect 745 -212 773 -184
rect 811 -212 839 -184
rect 877 -212 905 -184
rect 943 -212 971 -184
rect 1009 -212 1037 -184
rect 1075 -212 1103 -184
rect 1141 -212 1169 -184
rect 1207 -212 1235 -184
rect 1273 -212 1301 -184
rect 1339 -212 1367 -184
rect 1405 -212 1433 -184
rect 1471 -212 1499 -184
rect 1537 -212 1565 -184
rect 1603 -212 1631 -184
rect 1669 -212 1697 -184
rect 1735 -212 1763 -184
rect 1801 -212 1829 -184
rect 1867 -212 1895 -184
rect 1933 -212 1961 -184
rect 1999 -212 2027 -184
rect 2065 -212 2093 -184
rect 2131 -212 2159 -184
rect 2197 -212 2225 -184
rect -2225 -278 -2197 -250
rect -2159 -278 -2131 -250
rect -2093 -278 -2065 -250
rect -2027 -278 -1999 -250
rect -1961 -278 -1933 -250
rect -1895 -278 -1867 -250
rect -1829 -278 -1801 -250
rect -1763 -278 -1735 -250
rect -1697 -278 -1669 -250
rect -1631 -278 -1603 -250
rect -1565 -278 -1537 -250
rect -1499 -278 -1471 -250
rect -1433 -278 -1405 -250
rect -1367 -278 -1339 -250
rect -1301 -278 -1273 -250
rect -1235 -278 -1207 -250
rect -1169 -278 -1141 -250
rect -1103 -278 -1075 -250
rect -1037 -278 -1009 -250
rect -971 -278 -943 -250
rect -905 -278 -877 -250
rect -839 -278 -811 -250
rect -773 -278 -745 -250
rect -707 -278 -679 -250
rect -641 -278 -613 -250
rect -575 -278 -547 -250
rect -509 -278 -481 -250
rect -443 -278 -415 -250
rect -377 -278 -349 -250
rect -311 -278 -283 -250
rect -245 -278 -217 -250
rect -179 -278 -151 -250
rect -113 -278 -85 -250
rect -47 -278 -19 -250
rect 19 -278 47 -250
rect 85 -278 113 -250
rect 151 -278 179 -250
rect 217 -278 245 -250
rect 283 -278 311 -250
rect 349 -278 377 -250
rect 415 -278 443 -250
rect 481 -278 509 -250
rect 547 -278 575 -250
rect 613 -278 641 -250
rect 679 -278 707 -250
rect 745 -278 773 -250
rect 811 -278 839 -250
rect 877 -278 905 -250
rect 943 -278 971 -250
rect 1009 -278 1037 -250
rect 1075 -278 1103 -250
rect 1141 -278 1169 -250
rect 1207 -278 1235 -250
rect 1273 -278 1301 -250
rect 1339 -278 1367 -250
rect 1405 -278 1433 -250
rect 1471 -278 1499 -250
rect 1537 -278 1565 -250
rect 1603 -278 1631 -250
rect 1669 -278 1697 -250
rect 1735 -278 1763 -250
rect 1801 -278 1829 -250
rect 1867 -278 1895 -250
rect 1933 -278 1961 -250
rect 1999 -278 2027 -250
rect 2065 -278 2093 -250
rect 2131 -278 2159 -250
rect 2197 -278 2225 -250
rect -2225 -344 -2197 -316
rect -2159 -344 -2131 -316
rect -2093 -344 -2065 -316
rect -2027 -344 -1999 -316
rect -1961 -344 -1933 -316
rect -1895 -344 -1867 -316
rect -1829 -344 -1801 -316
rect -1763 -344 -1735 -316
rect -1697 -344 -1669 -316
rect -1631 -344 -1603 -316
rect -1565 -344 -1537 -316
rect -1499 -344 -1471 -316
rect -1433 -344 -1405 -316
rect -1367 -344 -1339 -316
rect -1301 -344 -1273 -316
rect -1235 -344 -1207 -316
rect -1169 -344 -1141 -316
rect -1103 -344 -1075 -316
rect -1037 -344 -1009 -316
rect -971 -344 -943 -316
rect -905 -344 -877 -316
rect -839 -344 -811 -316
rect -773 -344 -745 -316
rect -707 -344 -679 -316
rect -641 -344 -613 -316
rect -575 -344 -547 -316
rect -509 -344 -481 -316
rect -443 -344 -415 -316
rect -377 -344 -349 -316
rect -311 -344 -283 -316
rect -245 -344 -217 -316
rect -179 -344 -151 -316
rect -113 -344 -85 -316
rect -47 -344 -19 -316
rect 19 -344 47 -316
rect 85 -344 113 -316
rect 151 -344 179 -316
rect 217 -344 245 -316
rect 283 -344 311 -316
rect 349 -344 377 -316
rect 415 -344 443 -316
rect 481 -344 509 -316
rect 547 -344 575 -316
rect 613 -344 641 -316
rect 679 -344 707 -316
rect 745 -344 773 -316
rect 811 -344 839 -316
rect 877 -344 905 -316
rect 943 -344 971 -316
rect 1009 -344 1037 -316
rect 1075 -344 1103 -316
rect 1141 -344 1169 -316
rect 1207 -344 1235 -316
rect 1273 -344 1301 -316
rect 1339 -344 1367 -316
rect 1405 -344 1433 -316
rect 1471 -344 1499 -316
rect 1537 -344 1565 -316
rect 1603 -344 1631 -316
rect 1669 -344 1697 -316
rect 1735 -344 1763 -316
rect 1801 -344 1829 -316
rect 1867 -344 1895 -316
rect 1933 -344 1961 -316
rect 1999 -344 2027 -316
rect 2065 -344 2093 -316
rect 2131 -344 2159 -316
rect 2197 -344 2225 -316
<< metal4 >>
rect -2230 344 2230 349
rect -2230 316 -2225 344
rect -2197 316 -2159 344
rect -2131 316 -2093 344
rect -2065 316 -2027 344
rect -1999 316 -1961 344
rect -1933 316 -1895 344
rect -1867 316 -1829 344
rect -1801 316 -1763 344
rect -1735 316 -1697 344
rect -1669 316 -1631 344
rect -1603 316 -1565 344
rect -1537 316 -1499 344
rect -1471 316 -1433 344
rect -1405 316 -1367 344
rect -1339 316 -1301 344
rect -1273 316 -1235 344
rect -1207 316 -1169 344
rect -1141 316 -1103 344
rect -1075 316 -1037 344
rect -1009 316 -971 344
rect -943 316 -905 344
rect -877 316 -839 344
rect -811 316 -773 344
rect -745 316 -707 344
rect -679 316 -641 344
rect -613 316 -575 344
rect -547 316 -509 344
rect -481 316 -443 344
rect -415 316 -377 344
rect -349 316 -311 344
rect -283 316 -245 344
rect -217 316 -179 344
rect -151 316 -113 344
rect -85 316 -47 344
rect -19 316 19 344
rect 47 316 85 344
rect 113 316 151 344
rect 179 316 217 344
rect 245 316 283 344
rect 311 316 349 344
rect 377 316 415 344
rect 443 316 481 344
rect 509 316 547 344
rect 575 316 613 344
rect 641 316 679 344
rect 707 316 745 344
rect 773 316 811 344
rect 839 316 877 344
rect 905 316 943 344
rect 971 316 1009 344
rect 1037 316 1075 344
rect 1103 316 1141 344
rect 1169 316 1207 344
rect 1235 316 1273 344
rect 1301 316 1339 344
rect 1367 316 1405 344
rect 1433 316 1471 344
rect 1499 316 1537 344
rect 1565 316 1603 344
rect 1631 316 1669 344
rect 1697 316 1735 344
rect 1763 316 1801 344
rect 1829 316 1867 344
rect 1895 316 1933 344
rect 1961 316 1999 344
rect 2027 316 2065 344
rect 2093 316 2131 344
rect 2159 316 2197 344
rect 2225 316 2230 344
rect -2230 278 2230 316
rect -2230 250 -2225 278
rect -2197 250 -2159 278
rect -2131 250 -2093 278
rect -2065 250 -2027 278
rect -1999 250 -1961 278
rect -1933 250 -1895 278
rect -1867 250 -1829 278
rect -1801 250 -1763 278
rect -1735 250 -1697 278
rect -1669 250 -1631 278
rect -1603 250 -1565 278
rect -1537 250 -1499 278
rect -1471 250 -1433 278
rect -1405 250 -1367 278
rect -1339 250 -1301 278
rect -1273 250 -1235 278
rect -1207 250 -1169 278
rect -1141 250 -1103 278
rect -1075 250 -1037 278
rect -1009 250 -971 278
rect -943 250 -905 278
rect -877 250 -839 278
rect -811 250 -773 278
rect -745 250 -707 278
rect -679 250 -641 278
rect -613 250 -575 278
rect -547 250 -509 278
rect -481 250 -443 278
rect -415 250 -377 278
rect -349 250 -311 278
rect -283 250 -245 278
rect -217 250 -179 278
rect -151 250 -113 278
rect -85 250 -47 278
rect -19 250 19 278
rect 47 250 85 278
rect 113 250 151 278
rect 179 250 217 278
rect 245 250 283 278
rect 311 250 349 278
rect 377 250 415 278
rect 443 250 481 278
rect 509 250 547 278
rect 575 250 613 278
rect 641 250 679 278
rect 707 250 745 278
rect 773 250 811 278
rect 839 250 877 278
rect 905 250 943 278
rect 971 250 1009 278
rect 1037 250 1075 278
rect 1103 250 1141 278
rect 1169 250 1207 278
rect 1235 250 1273 278
rect 1301 250 1339 278
rect 1367 250 1405 278
rect 1433 250 1471 278
rect 1499 250 1537 278
rect 1565 250 1603 278
rect 1631 250 1669 278
rect 1697 250 1735 278
rect 1763 250 1801 278
rect 1829 250 1867 278
rect 1895 250 1933 278
rect 1961 250 1999 278
rect 2027 250 2065 278
rect 2093 250 2131 278
rect 2159 250 2197 278
rect 2225 250 2230 278
rect -2230 212 2230 250
rect -2230 184 -2225 212
rect -2197 184 -2159 212
rect -2131 184 -2093 212
rect -2065 184 -2027 212
rect -1999 184 -1961 212
rect -1933 184 -1895 212
rect -1867 184 -1829 212
rect -1801 184 -1763 212
rect -1735 184 -1697 212
rect -1669 184 -1631 212
rect -1603 184 -1565 212
rect -1537 184 -1499 212
rect -1471 184 -1433 212
rect -1405 184 -1367 212
rect -1339 184 -1301 212
rect -1273 184 -1235 212
rect -1207 184 -1169 212
rect -1141 184 -1103 212
rect -1075 184 -1037 212
rect -1009 184 -971 212
rect -943 184 -905 212
rect -877 184 -839 212
rect -811 184 -773 212
rect -745 184 -707 212
rect -679 184 -641 212
rect -613 184 -575 212
rect -547 184 -509 212
rect -481 184 -443 212
rect -415 184 -377 212
rect -349 184 -311 212
rect -283 184 -245 212
rect -217 184 -179 212
rect -151 184 -113 212
rect -85 184 -47 212
rect -19 184 19 212
rect 47 184 85 212
rect 113 184 151 212
rect 179 184 217 212
rect 245 184 283 212
rect 311 184 349 212
rect 377 184 415 212
rect 443 184 481 212
rect 509 184 547 212
rect 575 184 613 212
rect 641 184 679 212
rect 707 184 745 212
rect 773 184 811 212
rect 839 184 877 212
rect 905 184 943 212
rect 971 184 1009 212
rect 1037 184 1075 212
rect 1103 184 1141 212
rect 1169 184 1207 212
rect 1235 184 1273 212
rect 1301 184 1339 212
rect 1367 184 1405 212
rect 1433 184 1471 212
rect 1499 184 1537 212
rect 1565 184 1603 212
rect 1631 184 1669 212
rect 1697 184 1735 212
rect 1763 184 1801 212
rect 1829 184 1867 212
rect 1895 184 1933 212
rect 1961 184 1999 212
rect 2027 184 2065 212
rect 2093 184 2131 212
rect 2159 184 2197 212
rect 2225 184 2230 212
rect -2230 146 2230 184
rect -2230 118 -2225 146
rect -2197 118 -2159 146
rect -2131 118 -2093 146
rect -2065 118 -2027 146
rect -1999 118 -1961 146
rect -1933 118 -1895 146
rect -1867 118 -1829 146
rect -1801 118 -1763 146
rect -1735 118 -1697 146
rect -1669 118 -1631 146
rect -1603 118 -1565 146
rect -1537 118 -1499 146
rect -1471 118 -1433 146
rect -1405 118 -1367 146
rect -1339 118 -1301 146
rect -1273 118 -1235 146
rect -1207 118 -1169 146
rect -1141 118 -1103 146
rect -1075 118 -1037 146
rect -1009 118 -971 146
rect -943 118 -905 146
rect -877 118 -839 146
rect -811 118 -773 146
rect -745 118 -707 146
rect -679 118 -641 146
rect -613 118 -575 146
rect -547 118 -509 146
rect -481 118 -443 146
rect -415 118 -377 146
rect -349 118 -311 146
rect -283 118 -245 146
rect -217 118 -179 146
rect -151 118 -113 146
rect -85 118 -47 146
rect -19 118 19 146
rect 47 118 85 146
rect 113 118 151 146
rect 179 118 217 146
rect 245 118 283 146
rect 311 118 349 146
rect 377 118 415 146
rect 443 118 481 146
rect 509 118 547 146
rect 575 118 613 146
rect 641 118 679 146
rect 707 118 745 146
rect 773 118 811 146
rect 839 118 877 146
rect 905 118 943 146
rect 971 118 1009 146
rect 1037 118 1075 146
rect 1103 118 1141 146
rect 1169 118 1207 146
rect 1235 118 1273 146
rect 1301 118 1339 146
rect 1367 118 1405 146
rect 1433 118 1471 146
rect 1499 118 1537 146
rect 1565 118 1603 146
rect 1631 118 1669 146
rect 1697 118 1735 146
rect 1763 118 1801 146
rect 1829 118 1867 146
rect 1895 118 1933 146
rect 1961 118 1999 146
rect 2027 118 2065 146
rect 2093 118 2131 146
rect 2159 118 2197 146
rect 2225 118 2230 146
rect -2230 80 2230 118
rect -2230 52 -2225 80
rect -2197 52 -2159 80
rect -2131 52 -2093 80
rect -2065 52 -2027 80
rect -1999 52 -1961 80
rect -1933 52 -1895 80
rect -1867 52 -1829 80
rect -1801 52 -1763 80
rect -1735 52 -1697 80
rect -1669 52 -1631 80
rect -1603 52 -1565 80
rect -1537 52 -1499 80
rect -1471 52 -1433 80
rect -1405 52 -1367 80
rect -1339 52 -1301 80
rect -1273 52 -1235 80
rect -1207 52 -1169 80
rect -1141 52 -1103 80
rect -1075 52 -1037 80
rect -1009 52 -971 80
rect -943 52 -905 80
rect -877 52 -839 80
rect -811 52 -773 80
rect -745 52 -707 80
rect -679 52 -641 80
rect -613 52 -575 80
rect -547 52 -509 80
rect -481 52 -443 80
rect -415 52 -377 80
rect -349 52 -311 80
rect -283 52 -245 80
rect -217 52 -179 80
rect -151 52 -113 80
rect -85 52 -47 80
rect -19 52 19 80
rect 47 52 85 80
rect 113 52 151 80
rect 179 52 217 80
rect 245 52 283 80
rect 311 52 349 80
rect 377 52 415 80
rect 443 52 481 80
rect 509 52 547 80
rect 575 52 613 80
rect 641 52 679 80
rect 707 52 745 80
rect 773 52 811 80
rect 839 52 877 80
rect 905 52 943 80
rect 971 52 1009 80
rect 1037 52 1075 80
rect 1103 52 1141 80
rect 1169 52 1207 80
rect 1235 52 1273 80
rect 1301 52 1339 80
rect 1367 52 1405 80
rect 1433 52 1471 80
rect 1499 52 1537 80
rect 1565 52 1603 80
rect 1631 52 1669 80
rect 1697 52 1735 80
rect 1763 52 1801 80
rect 1829 52 1867 80
rect 1895 52 1933 80
rect 1961 52 1999 80
rect 2027 52 2065 80
rect 2093 52 2131 80
rect 2159 52 2197 80
rect 2225 52 2230 80
rect -2230 14 2230 52
rect -2230 -14 -2225 14
rect -2197 -14 -2159 14
rect -2131 -14 -2093 14
rect -2065 -14 -2027 14
rect -1999 -14 -1961 14
rect -1933 -14 -1895 14
rect -1867 -14 -1829 14
rect -1801 -14 -1763 14
rect -1735 -14 -1697 14
rect -1669 -14 -1631 14
rect -1603 -14 -1565 14
rect -1537 -14 -1499 14
rect -1471 -14 -1433 14
rect -1405 -14 -1367 14
rect -1339 -14 -1301 14
rect -1273 -14 -1235 14
rect -1207 -14 -1169 14
rect -1141 -14 -1103 14
rect -1075 -14 -1037 14
rect -1009 -14 -971 14
rect -943 -14 -905 14
rect -877 -14 -839 14
rect -811 -14 -773 14
rect -745 -14 -707 14
rect -679 -14 -641 14
rect -613 -14 -575 14
rect -547 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 19 14
rect 47 -14 85 14
rect 113 -14 151 14
rect 179 -14 217 14
rect 245 -14 283 14
rect 311 -14 349 14
rect 377 -14 415 14
rect 443 -14 481 14
rect 509 -14 547 14
rect 575 -14 613 14
rect 641 -14 679 14
rect 707 -14 745 14
rect 773 -14 811 14
rect 839 -14 877 14
rect 905 -14 943 14
rect 971 -14 1009 14
rect 1037 -14 1075 14
rect 1103 -14 1141 14
rect 1169 -14 1207 14
rect 1235 -14 1273 14
rect 1301 -14 1339 14
rect 1367 -14 1405 14
rect 1433 -14 1471 14
rect 1499 -14 1537 14
rect 1565 -14 1603 14
rect 1631 -14 1669 14
rect 1697 -14 1735 14
rect 1763 -14 1801 14
rect 1829 -14 1867 14
rect 1895 -14 1933 14
rect 1961 -14 1999 14
rect 2027 -14 2065 14
rect 2093 -14 2131 14
rect 2159 -14 2197 14
rect 2225 -14 2230 14
rect -2230 -52 2230 -14
rect -2230 -80 -2225 -52
rect -2197 -80 -2159 -52
rect -2131 -80 -2093 -52
rect -2065 -80 -2027 -52
rect -1999 -80 -1961 -52
rect -1933 -80 -1895 -52
rect -1867 -80 -1829 -52
rect -1801 -80 -1763 -52
rect -1735 -80 -1697 -52
rect -1669 -80 -1631 -52
rect -1603 -80 -1565 -52
rect -1537 -80 -1499 -52
rect -1471 -80 -1433 -52
rect -1405 -80 -1367 -52
rect -1339 -80 -1301 -52
rect -1273 -80 -1235 -52
rect -1207 -80 -1169 -52
rect -1141 -80 -1103 -52
rect -1075 -80 -1037 -52
rect -1009 -80 -971 -52
rect -943 -80 -905 -52
rect -877 -80 -839 -52
rect -811 -80 -773 -52
rect -745 -80 -707 -52
rect -679 -80 -641 -52
rect -613 -80 -575 -52
rect -547 -80 -509 -52
rect -481 -80 -443 -52
rect -415 -80 -377 -52
rect -349 -80 -311 -52
rect -283 -80 -245 -52
rect -217 -80 -179 -52
rect -151 -80 -113 -52
rect -85 -80 -47 -52
rect -19 -80 19 -52
rect 47 -80 85 -52
rect 113 -80 151 -52
rect 179 -80 217 -52
rect 245 -80 283 -52
rect 311 -80 349 -52
rect 377 -80 415 -52
rect 443 -80 481 -52
rect 509 -80 547 -52
rect 575 -80 613 -52
rect 641 -80 679 -52
rect 707 -80 745 -52
rect 773 -80 811 -52
rect 839 -80 877 -52
rect 905 -80 943 -52
rect 971 -80 1009 -52
rect 1037 -80 1075 -52
rect 1103 -80 1141 -52
rect 1169 -80 1207 -52
rect 1235 -80 1273 -52
rect 1301 -80 1339 -52
rect 1367 -80 1405 -52
rect 1433 -80 1471 -52
rect 1499 -80 1537 -52
rect 1565 -80 1603 -52
rect 1631 -80 1669 -52
rect 1697 -80 1735 -52
rect 1763 -80 1801 -52
rect 1829 -80 1867 -52
rect 1895 -80 1933 -52
rect 1961 -80 1999 -52
rect 2027 -80 2065 -52
rect 2093 -80 2131 -52
rect 2159 -80 2197 -52
rect 2225 -80 2230 -52
rect -2230 -118 2230 -80
rect -2230 -146 -2225 -118
rect -2197 -146 -2159 -118
rect -2131 -146 -2093 -118
rect -2065 -146 -2027 -118
rect -1999 -146 -1961 -118
rect -1933 -146 -1895 -118
rect -1867 -146 -1829 -118
rect -1801 -146 -1763 -118
rect -1735 -146 -1697 -118
rect -1669 -146 -1631 -118
rect -1603 -146 -1565 -118
rect -1537 -146 -1499 -118
rect -1471 -146 -1433 -118
rect -1405 -146 -1367 -118
rect -1339 -146 -1301 -118
rect -1273 -146 -1235 -118
rect -1207 -146 -1169 -118
rect -1141 -146 -1103 -118
rect -1075 -146 -1037 -118
rect -1009 -146 -971 -118
rect -943 -146 -905 -118
rect -877 -146 -839 -118
rect -811 -146 -773 -118
rect -745 -146 -707 -118
rect -679 -146 -641 -118
rect -613 -146 -575 -118
rect -547 -146 -509 -118
rect -481 -146 -443 -118
rect -415 -146 -377 -118
rect -349 -146 -311 -118
rect -283 -146 -245 -118
rect -217 -146 -179 -118
rect -151 -146 -113 -118
rect -85 -146 -47 -118
rect -19 -146 19 -118
rect 47 -146 85 -118
rect 113 -146 151 -118
rect 179 -146 217 -118
rect 245 -146 283 -118
rect 311 -146 349 -118
rect 377 -146 415 -118
rect 443 -146 481 -118
rect 509 -146 547 -118
rect 575 -146 613 -118
rect 641 -146 679 -118
rect 707 -146 745 -118
rect 773 -146 811 -118
rect 839 -146 877 -118
rect 905 -146 943 -118
rect 971 -146 1009 -118
rect 1037 -146 1075 -118
rect 1103 -146 1141 -118
rect 1169 -146 1207 -118
rect 1235 -146 1273 -118
rect 1301 -146 1339 -118
rect 1367 -146 1405 -118
rect 1433 -146 1471 -118
rect 1499 -146 1537 -118
rect 1565 -146 1603 -118
rect 1631 -146 1669 -118
rect 1697 -146 1735 -118
rect 1763 -146 1801 -118
rect 1829 -146 1867 -118
rect 1895 -146 1933 -118
rect 1961 -146 1999 -118
rect 2027 -146 2065 -118
rect 2093 -146 2131 -118
rect 2159 -146 2197 -118
rect 2225 -146 2230 -118
rect -2230 -184 2230 -146
rect -2230 -212 -2225 -184
rect -2197 -212 -2159 -184
rect -2131 -212 -2093 -184
rect -2065 -212 -2027 -184
rect -1999 -212 -1961 -184
rect -1933 -212 -1895 -184
rect -1867 -212 -1829 -184
rect -1801 -212 -1763 -184
rect -1735 -212 -1697 -184
rect -1669 -212 -1631 -184
rect -1603 -212 -1565 -184
rect -1537 -212 -1499 -184
rect -1471 -212 -1433 -184
rect -1405 -212 -1367 -184
rect -1339 -212 -1301 -184
rect -1273 -212 -1235 -184
rect -1207 -212 -1169 -184
rect -1141 -212 -1103 -184
rect -1075 -212 -1037 -184
rect -1009 -212 -971 -184
rect -943 -212 -905 -184
rect -877 -212 -839 -184
rect -811 -212 -773 -184
rect -745 -212 -707 -184
rect -679 -212 -641 -184
rect -613 -212 -575 -184
rect -547 -212 -509 -184
rect -481 -212 -443 -184
rect -415 -212 -377 -184
rect -349 -212 -311 -184
rect -283 -212 -245 -184
rect -217 -212 -179 -184
rect -151 -212 -113 -184
rect -85 -212 -47 -184
rect -19 -212 19 -184
rect 47 -212 85 -184
rect 113 -212 151 -184
rect 179 -212 217 -184
rect 245 -212 283 -184
rect 311 -212 349 -184
rect 377 -212 415 -184
rect 443 -212 481 -184
rect 509 -212 547 -184
rect 575 -212 613 -184
rect 641 -212 679 -184
rect 707 -212 745 -184
rect 773 -212 811 -184
rect 839 -212 877 -184
rect 905 -212 943 -184
rect 971 -212 1009 -184
rect 1037 -212 1075 -184
rect 1103 -212 1141 -184
rect 1169 -212 1207 -184
rect 1235 -212 1273 -184
rect 1301 -212 1339 -184
rect 1367 -212 1405 -184
rect 1433 -212 1471 -184
rect 1499 -212 1537 -184
rect 1565 -212 1603 -184
rect 1631 -212 1669 -184
rect 1697 -212 1735 -184
rect 1763 -212 1801 -184
rect 1829 -212 1867 -184
rect 1895 -212 1933 -184
rect 1961 -212 1999 -184
rect 2027 -212 2065 -184
rect 2093 -212 2131 -184
rect 2159 -212 2197 -184
rect 2225 -212 2230 -184
rect -2230 -250 2230 -212
rect -2230 -278 -2225 -250
rect -2197 -278 -2159 -250
rect -2131 -278 -2093 -250
rect -2065 -278 -2027 -250
rect -1999 -278 -1961 -250
rect -1933 -278 -1895 -250
rect -1867 -278 -1829 -250
rect -1801 -278 -1763 -250
rect -1735 -278 -1697 -250
rect -1669 -278 -1631 -250
rect -1603 -278 -1565 -250
rect -1537 -278 -1499 -250
rect -1471 -278 -1433 -250
rect -1405 -278 -1367 -250
rect -1339 -278 -1301 -250
rect -1273 -278 -1235 -250
rect -1207 -278 -1169 -250
rect -1141 -278 -1103 -250
rect -1075 -278 -1037 -250
rect -1009 -278 -971 -250
rect -943 -278 -905 -250
rect -877 -278 -839 -250
rect -811 -278 -773 -250
rect -745 -278 -707 -250
rect -679 -278 -641 -250
rect -613 -278 -575 -250
rect -547 -278 -509 -250
rect -481 -278 -443 -250
rect -415 -278 -377 -250
rect -349 -278 -311 -250
rect -283 -278 -245 -250
rect -217 -278 -179 -250
rect -151 -278 -113 -250
rect -85 -278 -47 -250
rect -19 -278 19 -250
rect 47 -278 85 -250
rect 113 -278 151 -250
rect 179 -278 217 -250
rect 245 -278 283 -250
rect 311 -278 349 -250
rect 377 -278 415 -250
rect 443 -278 481 -250
rect 509 -278 547 -250
rect 575 -278 613 -250
rect 641 -278 679 -250
rect 707 -278 745 -250
rect 773 -278 811 -250
rect 839 -278 877 -250
rect 905 -278 943 -250
rect 971 -278 1009 -250
rect 1037 -278 1075 -250
rect 1103 -278 1141 -250
rect 1169 -278 1207 -250
rect 1235 -278 1273 -250
rect 1301 -278 1339 -250
rect 1367 -278 1405 -250
rect 1433 -278 1471 -250
rect 1499 -278 1537 -250
rect 1565 -278 1603 -250
rect 1631 -278 1669 -250
rect 1697 -278 1735 -250
rect 1763 -278 1801 -250
rect 1829 -278 1867 -250
rect 1895 -278 1933 -250
rect 1961 -278 1999 -250
rect 2027 -278 2065 -250
rect 2093 -278 2131 -250
rect 2159 -278 2197 -250
rect 2225 -278 2230 -250
rect -2230 -316 2230 -278
rect -2230 -344 -2225 -316
rect -2197 -344 -2159 -316
rect -2131 -344 -2093 -316
rect -2065 -344 -2027 -316
rect -1999 -344 -1961 -316
rect -1933 -344 -1895 -316
rect -1867 -344 -1829 -316
rect -1801 -344 -1763 -316
rect -1735 -344 -1697 -316
rect -1669 -344 -1631 -316
rect -1603 -344 -1565 -316
rect -1537 -344 -1499 -316
rect -1471 -344 -1433 -316
rect -1405 -344 -1367 -316
rect -1339 -344 -1301 -316
rect -1273 -344 -1235 -316
rect -1207 -344 -1169 -316
rect -1141 -344 -1103 -316
rect -1075 -344 -1037 -316
rect -1009 -344 -971 -316
rect -943 -344 -905 -316
rect -877 -344 -839 -316
rect -811 -344 -773 -316
rect -745 -344 -707 -316
rect -679 -344 -641 -316
rect -613 -344 -575 -316
rect -547 -344 -509 -316
rect -481 -344 -443 -316
rect -415 -344 -377 -316
rect -349 -344 -311 -316
rect -283 -344 -245 -316
rect -217 -344 -179 -316
rect -151 -344 -113 -316
rect -85 -344 -47 -316
rect -19 -344 19 -316
rect 47 -344 85 -316
rect 113 -344 151 -316
rect 179 -344 217 -316
rect 245 -344 283 -316
rect 311 -344 349 -316
rect 377 -344 415 -316
rect 443 -344 481 -316
rect 509 -344 547 -316
rect 575 -344 613 -316
rect 641 -344 679 -316
rect 707 -344 745 -316
rect 773 -344 811 -316
rect 839 -344 877 -316
rect 905 -344 943 -316
rect 971 -344 1009 -316
rect 1037 -344 1075 -316
rect 1103 -344 1141 -316
rect 1169 -344 1207 -316
rect 1235 -344 1273 -316
rect 1301 -344 1339 -316
rect 1367 -344 1405 -316
rect 1433 -344 1471 -316
rect 1499 -344 1537 -316
rect 1565 -344 1603 -316
rect 1631 -344 1669 -316
rect 1697 -344 1735 -316
rect 1763 -344 1801 -316
rect 1829 -344 1867 -316
rect 1895 -344 1933 -316
rect 1961 -344 1999 -316
rect 2027 -344 2065 -316
rect 2093 -344 2131 -316
rect 2159 -344 2197 -316
rect 2225 -344 2230 -316
rect -2230 -349 2230 -344
<< end >>
