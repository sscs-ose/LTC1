magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2245 -22745 2245 22745
<< psubdiff >>
rect -245 20723 245 20745
rect -245 -20723 -223 20723
rect 223 -20723 245 20723
rect -245 -20745 245 -20723
<< psubdiffcont >>
rect -223 -20723 223 20723
<< metal1 >>
rect -234 20723 234 20734
rect -234 -20723 -223 20723
rect 223 -20723 234 20723
rect -234 -20734 234 -20723
<< end >>
