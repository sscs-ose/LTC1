magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1547 -1019 1085 1019
<< metal3 >>
rect -547 14 85 19
rect -547 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 85 14
rect -547 -19 85 -14
<< via3 >>
rect -542 -14 -514 14
rect -476 -14 -448 14
rect -410 -14 -382 14
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
rect 52 -14 80 14
<< metal4 >>
rect -547 14 85 19
rect -547 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 85 14
rect -547 -19 85 -14
<< end >>
