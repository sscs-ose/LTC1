magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2000 -2000 17064 59600
<< isosubstrate >>
rect 2267 55971 14818 57307
rect 4664 55935 7604 55971
rect 9908 55935 12848 55971
rect 10564 42616 14743 43682
rect 11970 40982 14743 42616
<< nwell >>
rect 354 55007 1644 56793
rect 873 54844 1644 55007
rect 873 53312 2754 54844
<< psubdiff >>
rect 2331 56054 2421 57134
rect 14645 56144 14735 57134
<< nsubdiff >>
rect 437 56688 1561 56710
rect 437 56642 459 56688
rect 975 56642 1305 56688
rect 1539 56642 1561 56688
rect 437 56620 1561 56642
rect 437 56556 527 56620
rect 1471 56534 1561 56620
rect 1471 56300 1493 56534
rect 1539 56300 1561 56534
rect 1471 56064 1561 56300
rect 1471 55548 1493 56064
rect 1539 55548 1561 56064
rect 1471 55312 1561 55548
rect 1471 55266 1493 55312
rect 1539 55266 1561 55312
rect 1471 55180 1561 55266
<< nsubdiffcont >>
rect 459 56642 975 56688
rect 1305 56642 1539 56688
rect 1493 56300 1539 56534
rect 1493 55548 1539 56064
rect 1493 55266 1539 55312
<< metal1 >>
rect 0 11002 122 57527
rect 704 57263 14134 57339
rect 448 56688 999 56699
rect 448 56642 459 56688
rect 975 56642 999 56688
rect 448 56631 999 56642
rect 448 56545 516 56631
rect 861 56225 937 56383
rect 1061 56315 1217 57263
rect 2342 56807 14724 57213
rect 1273 56688 1550 56699
rect 1273 56642 1305 56688
rect 1539 56642 1550 56688
rect 1273 56631 1550 56642
rect 1482 56534 1550 56631
rect 1482 56300 1493 56534
rect 1539 56300 1550 56534
rect 1482 56285 1550 56300
rect 2342 56471 2410 56807
rect 14350 56531 14560 56747
rect 14656 56471 14724 56807
rect 861 56149 1827 56225
rect 1482 56064 1550 56089
rect 1482 55548 1493 56064
rect 1539 55548 1550 56064
rect 1751 55723 1827 56149
rect 2342 56065 14724 56471
rect 6096 55741 6172 55773
rect 11340 55741 11416 55773
rect 1751 55647 2385 55723
rect 1482 55520 1550 55548
rect 448 55403 937 55471
rect 1143 55403 2667 55471
rect 1482 55312 1550 55345
rect 1482 55266 1493 55312
rect 1539 55266 1550 55312
rect 448 55169 516 55255
rect 1482 55169 1550 55266
rect 184 54724 921 55169
rect 184 53815 921 54260
rect 704 52943 3794 53019
rect 14408 48804 14564 49320
rect 3185 46133 3365 46520
rect 11589 46426 11742 47954
rect 14408 47836 14564 48352
rect 12241 46467 13567 46957
rect 10470 43143 10761 43639
rect 11846 43134 14677 43588
rect 11846 42659 12064 43134
rect 12064 41075 14677 41529
rect 11017 40804 11890 40910
rect 1913 40670 14134 40746
rect 1596 40504 5746 40580
rect 11416 40534 13842 40610
rect 10644 40398 13988 40474
rect 184 40250 954 40318
rect 6306 39057 6382 39459
rect 6306 38877 6504 39057
rect 8439 36834 13242 36910
rect 8293 36698 13102 36774
rect 2066 36562 2469 36638
rect 4461 36562 9150 36638
rect 1822 36426 3271 36502
rect 3659 36426 9010 36502
rect 2482 36290 12686 36366
rect 1310 36154 13754 36230
rect 3386 36018 13515 36094
rect 13919 35890 14119 38520
rect 1367 29741 6612 29841
rect 8696 29741 13699 29841
rect 1547 29561 6856 29661
rect 8452 29561 13519 29661
rect 2340 29319 3888 29481
rect 2340 24880 2502 29319
rect 3726 24880 3888 29319
rect 4112 24880 4274 29481
rect 4960 29319 5648 29481
rect 5486 24880 5648 29319
rect 5877 29319 7420 29481
rect 5877 24880 6039 29319
rect 7258 24880 7420 29319
rect 7646 29319 9190 29481
rect 7646 24880 7808 29319
rect 9028 24880 9190 29319
rect 9415 29319 10106 29481
rect 9415 24880 9577 29319
rect 10794 24880 10956 29481
rect 11181 29319 12729 29481
rect 11181 24880 11343 29319
rect 12567 24880 12729 29319
rect 14942 11002 15064 57557
rect 0 1217 268 11002
rect 14734 1217 15064 11002
rect 0 846 15064 1217
rect 0 708 122 846
rect 14942 708 15064 846
<< metal2 >>
rect 704 55400 780 57339
rect 1225 55400 1301 57600
rect 32 51200 122 52600
rect 184 38400 584 55169
rect 32 36800 122 38200
rect 704 36800 1104 53019
rect 1454 40579 1530 57339
rect 1184 40503 1530 40579
rect 1596 40504 1672 57339
rect 1886 53031 1962 57163
rect 2098 53666 2174 57600
rect 2670 56531 13350 56747
rect 3500 55849 13350 55925
rect 2309 54460 2385 55741
rect 2605 55399 4238 55475
rect 4162 54692 4238 55399
rect 8030 54829 8106 55849
rect 8499 54829 8575 55849
rect 8714 54973 8790 55849
rect 8937 54829 9013 55849
rect 9406 54829 9482 55849
rect 13274 55581 13350 55849
rect 4162 54616 13350 54692
rect 2098 53590 2347 53666
rect 3470 52943 3546 54152
rect 4162 53451 4238 54616
rect 8030 53870 8106 54616
rect 3769 53379 4238 53451
rect 3769 53361 4163 53379
rect 3769 52989 3863 53361
rect 4938 52615 5014 53418
rect 6766 52615 6842 53418
rect 7254 52615 7330 53418
rect 8718 52839 8794 54616
rect 9149 52777 9549 54200
rect 13274 53870 13350 54616
rect 9149 51265 9425 52777
rect 4594 46620 4994 50281
rect 5513 49080 5913 50281
rect 6416 49080 6816 50281
rect 3158 46020 4378 46520
rect 7427 46020 7627 49561
rect 7714 49080 8114 50281
rect 8416 49080 8816 50281
rect 9149 48662 9549 51265
rect 9713 46200 9931 48031
rect 10566 46330 10642 48046
rect 11589 47774 11742 49911
rect 10566 46254 10964 46330
rect 9713 44800 10470 46200
rect 10888 46170 10964 46254
rect 10888 44770 11093 46170
rect 1184 39027 1260 40503
rect 1913 39057 1989 40746
rect 4941 39057 5017 40746
rect 5670 39027 5746 40580
rect 7157 39057 7233 40746
rect 2393 37771 2783 37951
rect 165 28632 383 36600
rect 1310 32888 1386 36230
rect 1822 34267 1898 36502
rect 2066 34267 2142 36638
rect 2393 36562 2469 37771
rect 3195 36426 3271 37951
rect 2482 34267 2558 36366
rect 3427 36230 3503 38524
rect 3659 36426 3735 37951
rect 4147 37771 4537 37951
rect 4461 36562 4537 37771
rect 3092 36154 3503 36230
rect 3092 34499 3168 36154
rect 3386 34267 3462 36094
rect 4594 34267 4670 36094
rect 5498 34267 5574 36366
rect 5914 34267 5990 36638
rect 6158 34267 6234 36502
rect 6670 32888 6746 36230
rect 3020 30770 4243 30870
rect 4472 30770 6002 30870
rect 1444 30201 1544 30690
rect 1007 30101 1544 30201
rect 165 27223 586 28632
rect 1007 28401 1107 30101
rect 1688 30021 1788 30690
rect 1187 29921 1788 30021
rect 1187 28401 1287 29921
rect 1367 28401 1467 29829
rect 1547 28401 1655 29649
rect 3496 29366 3596 30690
rect 4143 29301 4243 30770
rect 4948 29301 5048 30690
rect 5902 29301 6002 30770
rect 6512 29753 6612 30690
rect 6756 29573 6856 30690
rect 7332 28015 7732 41648
rect 11017 40975 11093 44770
rect 11426 41647 11658 41827
rect 11200 40995 11290 41175
rect 11426 41080 11502 41647
rect 11626 41173 12060 41353
rect 11426 41004 11596 41080
rect 10644 38878 10720 40474
rect 10888 39057 10964 40746
rect 11200 39596 11276 40995
rect 8293 36698 8369 38700
rect 11520 38517 11596 41004
rect 8439 36834 8515 37951
rect 8318 32888 8394 36230
rect 8671 35882 8747 38486
rect 8895 37771 9566 37951
rect 8830 34267 8906 36502
rect 9074 34267 9150 36638
rect 9490 34267 9566 37771
rect 11690 37712 11890 40910
rect 11984 40398 12060 41173
rect 11690 37512 12090 37712
rect 10394 34267 10470 36094
rect 11602 34267 11678 36094
rect 11890 34499 12090 37512
rect 12406 36800 12624 44065
rect 13096 41773 13608 42996
rect 13766 40534 13842 57339
rect 13912 40398 13988 57339
rect 14058 40670 14134 57339
rect 14204 51352 14280 57600
rect 14204 45825 14280 49606
rect 13303 38507 13754 38687
rect 12506 34267 12582 36366
rect 12922 34267 12998 36774
rect 13166 34267 13242 36910
rect 13439 36018 13515 38035
rect 13678 32888 13754 38507
rect 9062 30770 10592 30870
rect 10821 30770 12044 30870
rect 8452 29573 8552 30690
rect 8696 29753 8796 30690
rect 9062 29301 9162 30770
rect 10016 29301 10116 30690
rect 10821 29301 10921 30770
rect 11468 29366 11568 30690
rect 13520 30021 13620 30690
rect 13764 30201 13864 30690
rect 13764 30101 14059 30201
rect 13520 29921 13879 30021
rect 13411 28401 13519 29649
rect 13599 28401 13699 29829
rect 13779 28401 13879 29921
rect 13959 28401 14059 30101
rect 165 14114 383 27223
rect 14380 17400 14780 56747
rect 14942 51200 15032 52600
rect 14942 36800 15032 38200
rect 14380 14400 14834 17400
rect 165 12894 870 14114
rect 165 1600 383 12894
rect 14634 12293 14834 14400
rect 14169 11223 14834 12293
use comp018green_esd_cdm  comp018green_esd_cdm_0
timestamp 1713338890
transform 1 0 4583 0 -1 49459
box -205 -83 5981 8547
use comp018green_inpath_cms_smt  comp018green_inpath_cms_smt_0
timestamp 1713338890
transform 1 0 848 0 -1 55852
box -144 -83 13504 14940
use comp018green_out_paddrv_16T  comp018green_out_paddrv_16T_0
timestamp 1713338890
transform 1 0 794 0 1 1465
box -360 -1465 13796 27678
use comp018green_out_predrv  comp018green_out_predrv_0
timestamp 1713338890
transform -1 0 7577 0 -1 35969
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_1
timestamp 1713338890
transform 1 0 479 0 -1 35969
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_2
timestamp 1713338890
transform 1 0 7487 0 -1 35969
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_3
timestamp 1713338890
transform -1 0 14585 0 -1 35969
box -83 -83 3677 6020
use comp018green_out_sigbuf_a  comp018green_out_sigbuf_a_0
timestamp 1713338890
transform -1 0 11282 0 1 37501
box -83 -83 2701 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_0
timestamp 1713338890
transform 1 0 798 0 1 37501
box -83 -803 2795 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_1
timestamp 1713338890
transform -1 0 6132 0 1 37501
box -83 -803 2795 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_2
timestamp 1713338890
transform 1 0 6042 0 1 37501
box -83 -803 2795 2911
use comp018green_sigbuf_1  comp018green_sigbuf_1_0
timestamp 1713338890
transform 1 0 11192 0 1 37501
box -83 -83 2889 2911
use M1_NWELL_CDNS_40661953145322  M1_NWELL_CDNS_40661953145322_0
timestamp 1713338890
transform 1 0 999 0 1 55135
box -645 -128 645 128
use M1_NWELL_CDNS_40661953145377  M1_NWELL_CDNS_40661953145377_0
timestamp 1713338890
transform 1 0 482 0 1 55900
box -128 -739 128 739
use M1_PSUB_CDNS_69033583165549  M1_PSUB_CDNS_69033583165549_0
timestamp 1713338890
transform 0 -1 8533 1 0 56099
box -45 -6202 45 6202
use M1_PSUB_CDNS_69033583165549  M1_PSUB_CDNS_69033583165549_1
timestamp 1713338890
transform 0 -1 8533 1 0 57179
box -45 -6202 45 6202
use M1_PSUB_CDNS_69033583165550  M1_PSUB_CDNS_69033583165550_0
timestamp 1713338890
transform 1 0 7502 0 1 1121
box -7237 -107 7237 107
use M1_PSUB_CDNS_69033583165552  M1_PSUB_CDNS_69033583165552_0
timestamp 1713338890
transform 1 0 11300 0 1 43149
box -558 -501 558 501
use M1_PSUB_CDNS_69033583165559  M1_PSUB_CDNS_69033583165559_0
timestamp 1713338890
transform 1 0 12098 0 1 42332
box -45 -1267 45 1267
use M1_PSUB_CDNS_69033583165559  M1_PSUB_CDNS_69033583165559_1
timestamp 1713338890
transform 1 0 14615 0 1 42332
box -45 -1267 45 1267
use M1_PSUB_CDNS_69033583165568  M1_PSUB_CDNS_69033583165568_0
timestamp 1713338890
transform 1 0 14690 0 1 56639
box -45 -421 45 421
use M1_PSUB_CDNS_69033583165568  M1_PSUB_CDNS_69033583165568_1
timestamp 1713338890
transform 1 0 2376 0 1 56639
box -45 -421 45 421
use M1_PSUB_CDNS_69033583165569  M1_PSUB_CDNS_69033583165569_0
timestamp 1713338890
transform 1 0 13333 0 1 41110
box -1173 -45 1173 45
use M1_PSUB_CDNS_69033583165569  M1_PSUB_CDNS_69033583165569_1
timestamp 1713338890
transform 1 0 13333 0 1 43554
box -1173 -45 1173 45
use M1_PSUB_CDNS_69033583165608  M1_PSUB_CDNS_69033583165608_0
timestamp 1713338890
transform -1 0 234 0 1 6174
box -45 -4839 45 4839
use M1_PSUB_CDNS_69033583165608  M1_PSUB_CDNS_69033583165608_1
timestamp 1713338890
transform 1 0 14768 0 1 6174
box -45 -4839 45 4839
use M2_M1_CDNS_69033583165515  M2_M1_CDNS_69033583165515_0
timestamp 1713338890
transform 1 0 13278 0 1 40288
box -506 -38 506 38
use M2_M1_CDNS_69033583165518  M2_M1_CDNS_69033583165518_0
timestamp 1713338890
transform 1 0 13952 0 1 57301
box -142 -38 142 38
use M2_M1_CDNS_69033583165521  M2_M1_CDNS_69033583165521_0
timestamp 1713338890
transform 1 0 14980 0 1 51893
box -38 -610 38 610
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_0
timestamp 1713338890
transform 1 0 1457 0 1 29791
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_1
timestamp 1713338890
transform 1 0 1637 0 1 29611
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_2
timestamp 1713338890
transform 1 0 3586 0 1 29404
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_3
timestamp 1713338890
transform 1 0 1400 0 1 36192
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_4
timestamp 1713338890
transform 1 0 1912 0 1 36464
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_5
timestamp 1713338890
transform 1 0 2572 0 1 36328
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_6
timestamp 1713338890
transform 1 0 1686 0 1 40542
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_7
timestamp 1713338890
transform 1 0 2003 0 1 40708
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_8
timestamp 1713338890
transform -1 0 3749 0 1 36464
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_9
timestamp 1713338890
transform 1 0 3181 0 1 36464
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_10
timestamp 1713338890
transform 1 0 3476 0 1 36056
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_11
timestamp 1713338890
transform -1 0 4580 0 1 36056
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_12
timestamp 1713338890
transform -1 0 4551 0 1 36600
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_13
timestamp 1713338890
transform -1 0 5484 0 1 36328
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_14
timestamp 1713338890
transform 1 0 5656 0 1 40542
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_15
timestamp 1713338890
transform -1 0 4927 0 1 40708
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_16
timestamp 1713338890
transform -1 0 5900 0 1 36600
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_17
timestamp 1713338890
transform -1 0 6144 0 1 36464
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_18
timestamp 1713338890
transform 1 0 6766 0 1 29611
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_19
timestamp 1713338890
transform 1 0 6522 0 1 29791
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_20
timestamp 1713338890
transform 1 0 8786 0 1 29791
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_21
timestamp 1713338890
transform 1 0 8542 0 1 29611
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_22
timestamp 1713338890
transform -1 0 11480 0 1 29404
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_23
timestamp 1713338890
transform 0 -1 8477 1 0 36924
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_24
timestamp 1713338890
transform -1 0 9060 0 1 36600
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_25
timestamp 1713338890
transform 1 0 8920 0 1 36464
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_26
timestamp 1713338890
transform 1 0 8383 0 1 36736
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_27
timestamp 1713338890
transform 1 0 8657 0 1 35920
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_28
timestamp 1713338890
transform 1 0 8408 0 1 36192
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_29
timestamp 1713338890
transform -1 0 6656 0 1 36192
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_30
timestamp 1713338890
transform 1 0 9580 0 1 36328
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_31
timestamp 1713338890
transform 1 0 10484 0 1 36056
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_32
timestamp 1713338890
transform -1 0 11588 0 1 36056
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_33
timestamp 1713338890
transform -1 0 7143 0 1 40708
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_34
timestamp 1713338890
transform 0 -1 11558 1 0 38607
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_35
timestamp 1713338890
transform 1 0 10734 0 1 40436
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_36
timestamp 1713338890
transform 1 0 10978 0 1 40708
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_37
timestamp 1713338890
transform 1 0 12074 0 1 40436
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_38
timestamp 1713338890
transform 1 0 11506 0 1 40572
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_39
timestamp 1713338890
transform 1 0 11792 0 1 40857
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_40
timestamp 1713338890
transform -1 0 13429 0 1 29611
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_41
timestamp 1713338890
transform -1 0 13609 0 1 29791
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_42
timestamp 1713338890
transform 1 0 13425 0 1 36056
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_43
timestamp 1713338890
transform -1 0 12596 0 1 36328
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_44
timestamp 1713338890
transform -1 0 13664 0 1 36192
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_45
timestamp 1713338890
transform 1 0 13152 0 1 36872
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_46
timestamp 1713338890
transform 1 0 13012 0 1 36736
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_47
timestamp 1713338890
transform 0 -1 14096 1 0 40760
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_48
timestamp 1713338890
transform 1 0 13898 0 1 40436
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_49
timestamp 1713338890
transform 1 0 13752 0 1 40572
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_50
timestamp 1713338890
transform 1 0 12512 0 1 44027
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_51
timestamp 1713338890
transform 1 0 3456 0 1 52981
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_52
timestamp 1713338890
transform 1 0 3773 0 1 52981
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_53
timestamp 1713338890
transform 1 0 7344 0 1 52653
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_54
timestamp 1713338890
transform 1 0 2683 0 1 55437
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_55
timestamp 1713338890
transform 1 0 1564 0 1 57301
box -90 -38 90 38
use M2_M1_CDNS_69033583165525  M2_M1_CDNS_69033583165525_0
timestamp 1713338890
transform 1 0 4980 0 1 52653
box -246 -38 246 38
use M2_M1_CDNS_69033583165525  M2_M1_CDNS_69033583165525_1
timestamp 1713338890
transform 1 0 6684 0 1 52653
box -246 -38 246 38
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_0
timestamp 1713338890
transform 1 0 2760 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_1
timestamp 1713338890
transform 1 0 3760 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_2
timestamp 1713338890
transform 1 0 4260 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_3
timestamp 1713338890
transform 1 0 5260 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_4
timestamp 1713338890
transform 1 0 5760 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_5
timestamp 1713338890
transform 1 0 6760 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_6
timestamp 1713338890
transform 1 0 7260 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_7
timestamp 1713338890
transform 1 0 8260 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_8
timestamp 1713338890
transform 1 0 8760 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_9
timestamp 1713338890
transform 1 0 10260 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_10
timestamp 1713338890
transform 1 0 9760 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_11
timestamp 1713338890
transform 1 0 11260 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_12
timestamp 1713338890
transform 1 0 11760 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_13
timestamp 1713338890
transform 1 0 12760 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_14
timestamp 1713338890
transform 1 0 13260 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_15
timestamp 1713338890
transform 1 0 14470 0 1 56637
box -90 -90 90 90
use M2_M1_CDNS_69033583165539  M2_M1_CDNS_69033583165539_0
timestamp 1713338890
transform 1 0 84 0 1 37493
box -38 -662 38 662
use M2_M1_CDNS_69033583165539  M2_M1_CDNS_69033583165539_1
timestamp 1713338890
transform 1 0 3646 0 1 42293
box -38 -662 38 662
use M2_M1_CDNS_69033583165539  M2_M1_CDNS_69033583165539_2
timestamp 1713338890
transform 1 0 14980 0 1 37493
box -38 -662 38 662
use M2_M1_CDNS_69033583165539  M2_M1_CDNS_69033583165539_3
timestamp 1713338890
transform 1 0 3646 0 1 43893
box -38 -662 38 662
use M2_M1_CDNS_69033583165539  M2_M1_CDNS_69033583165539_4
timestamp 1713338890
transform 1 0 84 0 1 51893
box -38 -662 38 662
use M2_M1_CDNS_69033583165540  M2_M1_CDNS_69033583165540_0
timestamp 1713338890
transform 1 0 524 0 1 31953
box -38 -1910 38 1910
use M2_M1_CDNS_69033583165540  M2_M1_CDNS_69033583165540_1
timestamp 1713338890
transform 1 0 14540 0 1 31953
box -38 -1910 38 1910
use M2_M1_CDNS_69033583165541  M2_M1_CDNS_69033583165541_0
timestamp 1713338890
transform 1 0 10941 0 1 37542
box -610 -38 610 38
use M2_M1_CDNS_69033583165548  M2_M1_CDNS_69033583165548_0
timestamp 1713338890
transform 1 0 8066 0 1 56268
box -5556 -162 5556 162
use M2_M1_CDNS_69033583165548  M2_M1_CDNS_69033583165548_1
timestamp 1713338890
transform 1 0 8066 0 1 57010
box -5556 -162 5556 162
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_0
timestamp 1713338890
transform 1 0 3302 0 1 31884
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_1
timestamp 1713338890
transform 1 0 3790 0 1 31834
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_2
timestamp 1713338890
transform 1 0 4266 0 1 31834
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_3
timestamp 1713338890
transform 1 0 4754 0 1 31884
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_4
timestamp 1713338890
transform 1 0 5242 0 1 31884
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_5
timestamp 1713338890
transform 1 0 5658 0 1 31884
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_6
timestamp 1713338890
transform 1 0 9406 0 1 31884
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_7
timestamp 1713338890
transform 1 0 9822 0 1 31884
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_8
timestamp 1713338890
transform 1 0 10310 0 1 31884
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_9
timestamp 1713338890
transform 1 0 10798 0 1 31834
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_10
timestamp 1713338890
transform 1 0 11274 0 1 31834
box -38 -818 38 818
use M2_M1_CDNS_69033583165555  M2_M1_CDNS_69033583165555_11
timestamp 1713338890
transform 1 0 11762 0 1 31884
box -38 -818 38 818
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_0
timestamp 1713338890
transform 1 0 843 0 1 38018
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_1
timestamp 1713338890
transform 1 0 3465 0 1 38018
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_2
timestamp 1713338890
transform 1 0 6087 0 1 39264
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_3
timestamp 1713338890
transform 1 0 6087 0 1 38018
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_4
timestamp 1713338890
transform 1 0 8709 0 1 38018
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_5
timestamp 1713338890
transform 1 0 10365 0 1 39294
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_6
timestamp 1713338890
transform 1 0 11238 0 1 39294
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_7
timestamp 1713338890
transform 1 0 10820 0 1 48866
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_8
timestamp 1713338890
transform 1 0 3508 0 1 53877
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_9
timestamp 1713338890
transform 1 0 8756 0 1 53877
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_10
timestamp 1713338890
transform 1 0 8752 0 1 55335
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_11
timestamp 1713338890
transform 1 0 8537 0 1 55335
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_12
timestamp 1713338890
transform 1 0 8975 0 1 55335
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_13
timestamp 1713338890
transform 1 0 8068 0 1 55335
box -38 -506 38 506
use M2_M1_CDNS_69033583165558  M2_M1_CDNS_69033583165558_14
timestamp 1713338890
transform 1 0 9444 0 1 55335
box -38 -506 38 506
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_0
timestamp 1713338890
transform 1 0 1809 0 1 39502
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_1
timestamp 1713338890
transform 1 0 5121 0 1 39472
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_2
timestamp 1713338890
transform 1 0 7053 0 1 39472
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_3
timestamp 1713338890
transform 1 0 11039 0 1 47432
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_4
timestamp 1713338890
transform 1 0 4976 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_5
timestamp 1713338890
transform 1 0 5464 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_6
timestamp 1713338890
transform 1 0 5952 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_7
timestamp 1713338890
transform 1 0 6316 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_8
timestamp 1713338890
transform 1 0 6804 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_9
timestamp 1713338890
transform 1 0 7292 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_10
timestamp 1713338890
transform 1 0 10220 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_11
timestamp 1713338890
transform 1 0 10708 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_12
timestamp 1713338890
transform 1 0 11196 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_13
timestamp 1713338890
transform 1 0 11560 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_14
timestamp 1713338890
transform 1 0 12048 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165563  M2_M1_CDNS_69033583165563_15
timestamp 1713338890
transform 1 0 12536 0 1 53716
box -38 -298 38 298
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_0
timestamp 1713338890
transform 1 0 6134 0 1 53825
box -38 -454 38 454
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_1
timestamp 1713338890
transform 1 0 11378 0 1 53825
box -38 -454 38 454
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_2
timestamp 1713338890
transform 1 0 4788 0 1 55287
box -38 -454 38 454
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_3
timestamp 1713338890
transform 1 0 6134 0 1 55287
box -38 -454 38 454
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_4
timestamp 1713338890
transform 1 0 7480 0 1 55287
box -38 -454 38 454
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_5
timestamp 1713338890
transform 1 0 10032 0 1 55287
box -38 -454 38 454
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_6
timestamp 1713338890
transform 1 0 11378 0 1 55287
box -38 -454 38 454
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_7
timestamp 1713338890
transform 1 0 12724 0 1 55287
box -38 -454 38 454
use M2_M1_CDNS_69033583165565  M2_M1_CDNS_69033583165565_8
timestamp 1713338890
transform 1 0 13312 0 1 55287
box -38 -454 38 454
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_0
timestamp 1713338890
transform 1 0 4200 0 1 53773
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_1
timestamp 1713338890
transform 1 0 4788 0 1 53773
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_2
timestamp 1713338890
transform 1 0 7480 0 1 53773
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_3
timestamp 1713338890
transform 1 0 8068 0 1 53773
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_4
timestamp 1713338890
transform 1 0 10032 0 1 53773
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_5
timestamp 1713338890
transform 1 0 12724 0 1 53773
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_6
timestamp 1713338890
transform 1 0 13312 0 1 53773
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_7
timestamp 1713338890
transform 1 0 4976 0 1 55368
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_8
timestamp 1713338890
transform 1 0 5464 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_9
timestamp 1713338890
transform 1 0 5952 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_10
timestamp 1713338890
transform 1 0 6316 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_11
timestamp 1713338890
transform 1 0 6804 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_12
timestamp 1713338890
transform 1 0 7292 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_13
timestamp 1713338890
transform 1 0 10220 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_14
timestamp 1713338890
transform 1 0 11560 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_15
timestamp 1713338890
transform 1 0 10708 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_16
timestamp 1713338890
transform 1 0 11196 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_17
timestamp 1713338890
transform 1 0 12536 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165567  M2_M1_CDNS_69033583165567_18
timestamp 1713338890
transform 1 0 12048 0 1 55377
box -38 -402 38 402
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_0
timestamp 1713338890
transform 1 0 2104 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_1
timestamp 1713338890
transform 1 0 1860 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_2
timestamp 1713338890
transform 1 0 2520 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_3
timestamp 1713338890
transform 1 0 4193 0 1 29391
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_4
timestamp 1713338890
transform -1 0 4998 0 1 29391
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_5
timestamp 1713338890
transform -1 0 5952 0 1 29391
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_6
timestamp 1713338890
transform -1 0 5536 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_7
timestamp 1713338890
transform 1 0 5952 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_8
timestamp 1713338890
transform 1 0 6196 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_9
timestamp 1713338890
transform 1 0 2745 0 1 37861
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_10
timestamp 1713338890
transform 1 0 3233 0 1 37861
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_11
timestamp 1713338890
transform -1 0 3697 0 1 37861
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_12
timestamp 1713338890
transform -1 0 4185 0 1 37861
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_13
timestamp 1713338890
transform 1 0 9114 0 1 29391
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_14
timestamp 1713338890
transform 1 0 10068 0 1 29391
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_15
timestamp 1713338890
transform -1 0 10873 0 1 29391
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_16
timestamp 1713338890
transform 1 0 9112 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_17
timestamp 1713338890
transform -1 0 8868 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_18
timestamp 1713338890
transform 1 0 9528 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_19
timestamp 1713338890
transform 1 0 8933 0 1 37861
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_20
timestamp 1713338890
transform -1 0 8331 0 1 38610
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_21
timestamp 1713338890
transform -1 0 8477 0 1 37861
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_22
timestamp 1713338890
transform 1 0 10682 0 1 38968
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_23
timestamp 1713338890
transform 1 0 10926 0 1 38968
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_24
timestamp 1713338890
transform 1 0 11055 0 1 40894
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_25
timestamp 1713338890
transform 1 0 11324 0 1 41085
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_26
timestamp 1713338890
transform 1 0 11609 0 1 41263
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_27
timestamp 1713338890
transform 1 0 11609 0 1 41737
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_28
timestamp 1713338890
transform -1 0 12544 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_29
timestamp 1713338890
transform -1 0 12960 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_30
timestamp 1713338890
transform -1 0 13204 0 1 34357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_31
timestamp 1713338890
transform 1 0 13477 0 1 37945
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_32
timestamp 1713338890
transform 1 0 13341 0 1 38597
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_33
timestamp 1713338890
transform 1 0 13134 0 1 41863
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_34
timestamp 1713338890
transform 1 0 13134 0 1 42790
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_35
timestamp 1713338890
transform 1 0 13570 0 1 42790
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_36
timestamp 1713338890
transform 1 0 13570 0 1 41863
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_37
timestamp 1713338890
transform 1 0 14242 0 1 45915
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_38
timestamp 1713338890
transform 1 0 11656 0 1 47864
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_39
timestamp 1713338890
transform 1 0 2347 0 1 55633
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_40
timestamp 1713338890
transform 1 0 742 0 1 57249
box -38 -90 38 90
use M2_M1_CDNS_69033583165571  M2_M1_CDNS_69033583165571_0
timestamp 1713338890
transform 1 0 14472 0 1 48094
box -92 -254 92 254
use M2_M1_CDNS_69033583165571  M2_M1_CDNS_69033583165571_1
timestamp 1713338890
transform 1 0 14472 0 1 49062
box -92 -254 92 254
use M2_M1_CDNS_69033583165572  M2_M1_CDNS_69033583165572_0
timestamp 1713338890
transform 1 0 12460 0 1 46940
box -200 -38 200 38
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_0
timestamp 1713338890
transform 1 0 5713 0 1 49268
box -194 -142 194 142
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_1
timestamp 1713338890
transform 1 0 6616 0 1 49268
box -194 -142 194 142
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_2
timestamp 1713338890
transform 1 0 7914 0 1 49268
box -194 -142 194 142
use M2_M1_CDNS_69033583165574  M2_M1_CDNS_69033583165574_3
timestamp 1713338890
transform 1 0 8616 0 1 49268
box -194 -142 194 142
use M2_M1_CDNS_69033583165575  M2_M1_CDNS_69033583165575_0
timestamp 1713338890
transform 1 0 2270 0 1 36600
box -194 -38 194 38
use M2_M1_CDNS_69033583165575  M2_M1_CDNS_69033583165575_1
timestamp 1713338890
transform 1 0 384 0 1 40280
box -194 -38 194 38
use M2_M1_CDNS_69033583165575  M2_M1_CDNS_69033583165575_2
timestamp 1713338890
transform 1 0 8616 0 1 50243
box -194 -38 194 38
use M2_M1_CDNS_69033583165575  M2_M1_CDNS_69033583165575_3
timestamp 1713338890
transform 1 0 7914 0 1 50243
box -194 -38 194 38
use M2_M1_CDNS_69033583165575  M2_M1_CDNS_69033583165575_4
timestamp 1713338890
transform 1 0 904 0 1 52981
box -194 -38 194 38
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_0
timestamp 1713338890
transform 1 0 1006 0 1 31572
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_1
timestamp 1713338890
transform 1 0 2398 0 1 31572
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_2
timestamp 1713338890
transform 1 0 2814 0 1 31572
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_3
timestamp 1713338890
transform 1 0 7050 0 1 31572
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_4
timestamp 1713338890
transform 1 0 8014 0 1 31572
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_5
timestamp 1713338890
transform 1 0 12250 0 1 31572
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_6
timestamp 1713338890
transform 1 0 12666 0 1 31572
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_7
timestamp 1713338890
transform 1 0 14058 0 1 31572
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165581  M2_M1_CDNS_69033583165581_0
timestamp 1713338890
transform 1 0 4028 0 1 34620
box -38 -1338 38 1338
use M2_M1_CDNS_69033583165581  M2_M1_CDNS_69033583165581_1
timestamp 1713338890
transform 1 0 11036 0 1 34620
box -38 -1338 38 1338
use M2_M1_CDNS_69033583165584  M2_M1_CDNS_69033583165584_0
timestamp 1713338890
transform 1 0 762 0 1 35244
box -38 -714 38 714
use M2_M1_CDNS_69033583165584  M2_M1_CDNS_69033583165584_1
timestamp 1713338890
transform 1 0 3130 0 1 35244
box -38 -714 38 714
use M2_M1_CDNS_69033583165584  M2_M1_CDNS_69033583165584_2
timestamp 1713338890
transform 1 0 4926 0 1 35244
box -38 -714 38 714
use M2_M1_CDNS_69033583165584  M2_M1_CDNS_69033583165584_3
timestamp 1713338890
transform 1 0 10138 0 1 35244
box -38 -714 38 714
use M2_M1_CDNS_69033583165584  M2_M1_CDNS_69033583165584_4
timestamp 1713338890
transform 1 0 11934 0 1 35244
box -38 -714 38 714
use M2_M1_CDNS_69033583165586  M2_M1_CDNS_69033583165586_0
timestamp 1713338890
transform 1 0 524 0 1 35036
box -38 -922 38 922
use M2_M1_CDNS_69033583165586  M2_M1_CDNS_69033583165586_1
timestamp 1713338890
transform 1 0 4028 0 1 31915
box -38 -922 38 922
use M2_M1_CDNS_69033583165586  M2_M1_CDNS_69033583165586_2
timestamp 1713338890
transform 1 0 11036 0 1 31915
box -38 -922 38 922
use M2_M1_CDNS_69033583165587  M2_M1_CDNS_69033583165587_0
timestamp 1713338890
transform 1 0 2758 0 1 41044
box -922 -38 922 38
use M2_M1_CDNS_69033583165587  M2_M1_CDNS_69033583165587_1
timestamp 1713338890
transform 1 0 8810 0 1 40288
box -922 -38 922 38
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_0
timestamp 1713338890
transform 1 0 1494 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_1
timestamp 1713338890
transform 1 0 1738 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_2
timestamp 1713338890
transform 1 0 3058 0 1 30676
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_3
timestamp 1713338890
transform 1 0 3546 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_4
timestamp 1713338890
transform 1 0 4510 0 1 30676
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_5
timestamp 1713338890
transform 1 0 4998 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_6
timestamp 1713338890
transform 1 0 6806 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_7
timestamp 1713338890
transform 1 0 6562 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_8
timestamp 1713338890
transform 1 0 8746 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_9
timestamp 1713338890
transform 1 0 8502 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_10
timestamp 1713338890
transform -1 0 10066 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_11
timestamp 1713338890
transform -1 0 10554 0 1 30676
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_12
timestamp 1713338890
transform -1 0 11518 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_13
timestamp 1713338890
transform -1 0 12006 0 1 30676
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_14
timestamp 1713338890
transform -1 0 13814 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_15
timestamp 1713338890
transform -1 0 13570 0 1 30496
box -38 -194 38 194
use M2_M1_CDNS_69033583165592  M2_M1_CDNS_69033583165592_0
timestamp 1713338890
transform 1 0 2662 0 1 30081
box -662 -38 662 38
use M2_M1_CDNS_69033583165592  M2_M1_CDNS_69033583165592_1
timestamp 1713338890
transform 1 0 12599 0 1 30081
box -662 -38 662 38
use M2_M1_CDNS_69033583165593  M2_M1_CDNS_69033583165593_0
timestamp 1713338890
transform 1 0 3459 0 1 40288
box -1026 -38 1026 38
use M2_M1_CDNS_69033583165595  M2_M1_CDNS_69033583165595_0
timestamp 1713338890
transform 1 0 4334 0 1 50243
box -2482 -38 2482 38
use M2_M1_CDNS_69033583165596  M2_M1_CDNS_69033583165596_0
timestamp 1713338890
transform 1 0 4794 0 1 48654
box -162 -782 162 782
use M2_M1_CDNS_69033583165597  M2_M1_CDNS_69033583165597_0
timestamp 1713338890
transform 1 0 3646 0 1 47242
box -38 -558 38 558
use M2_M1_CDNS_69033583165598  M2_M1_CDNS_69033583165598_0
timestamp 1713338890
transform 1 0 3275 0 1 46270
box -90 -246 90 246
use M2_M1_CDNS_69033583165601  M2_M1_CDNS_69033583165601_0
timestamp 1713338890
transform 1 0 384 0 1 54036
box -162 -162 162 162
use M2_M1_CDNS_69033583165601  M2_M1_CDNS_69033583165601_1
timestamp 1713338890
transform 1 0 384 0 1 54945
box -162 -162 162 162
use M2_M1_CDNS_69033583165702  M2_M1_CDNS_69033583165702_0
timestamp 1713338890
transform 1 0 3798 0 1 55811
box -298 -38 298 38
use M3_M2_CDNS_69033583165547  M3_M2_CDNS_69033583165547_0
timestamp 1713338890
transform 1 0 8066 0 1 56268
box -5576 -180 5576 180
use M3_M2_CDNS_69033583165547  M3_M2_CDNS_69033583165547_1
timestamp 1713338890
transform 1 0 8066 0 1 57010
box -5576 -180 5576 180
use M3_M2_CDNS_69033583165553  M3_M2_CDNS_69033583165553_0
timestamp 1713338890
transform 1 0 13331 0 1 42380
box -150 -598 150 598
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_0
timestamp 1713338890
transform 1 0 3302 0 1 31884
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_1
timestamp 1713338890
transform 1 0 3790 0 1 31833
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_2
timestamp 1713338890
transform 1 0 4266 0 1 31833
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_3
timestamp 1713338890
transform 1 0 4754 0 1 31884
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_4
timestamp 1713338890
transform 1 0 5242 0 1 31884
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_5
timestamp 1713338890
transform 1 0 5658 0 1 31884
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_6
timestamp 1713338890
transform 1 0 9822 0 1 31884
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_7
timestamp 1713338890
transform 1 0 10310 0 1 31884
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_8
timestamp 1713338890
transform 1 0 9406 0 1 31884
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_9
timestamp 1713338890
transform 1 0 10798 0 1 31833
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_10
timestamp 1713338890
transform 1 0 11274 0 1 31833
box -38 -819 38 819
use M3_M2_CDNS_69033583165554  M3_M2_CDNS_69033583165554_11
timestamp 1713338890
transform 1 0 11762 0 1 31884
box -38 -819 38 819
use M3_M2_CDNS_69033583165556  M3_M2_CDNS_69033583165556_0
timestamp 1713338890
transform 1 0 10960 0 1 37542
box -535 -38 535 38
use M3_M2_CDNS_69033583165556  M3_M2_CDNS_69033583165556_1
timestamp 1713338890
transform 1 0 13283 0 1 40288
box -535 -38 535 38
use M3_M2_CDNS_69033583165557  M3_M2_CDNS_69033583165557_0
timestamp 1713338890
transform 1 0 6087 0 1 39229
box -38 -535 38 535
use M3_M2_CDNS_69033583165557  M3_M2_CDNS_69033583165557_1
timestamp 1713338890
transform 1 0 10365 0 1 39235
box -38 -535 38 535
use M3_M2_CDNS_69033583165557  M3_M2_CDNS_69033583165557_2
timestamp 1713338890
transform 1 0 11238 0 1 39235
box -38 -535 38 535
use M3_M2_CDNS_69033583165557  M3_M2_CDNS_69033583165557_3
timestamp 1713338890
transform 1 0 3646 0 1 47235
box -38 -535 38 535
use M3_M2_CDNS_69033583165557  M3_M2_CDNS_69033583165557_4
timestamp 1713338890
transform 1 0 10820 0 1 48835
box -38 -535 38 535
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_0
timestamp 1713338890
transform 1 0 904 0 1 37493
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_1
timestamp 1713338890
transform 1 0 384 0 1 39093
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_2
timestamp 1713338890
transform 1 0 14580 0 1 29500
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_3
timestamp 1713338890
transform 1 0 14580 0 1 40693
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_4
timestamp 1713338890
transform 1 0 14580 0 1 47093
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_5
timestamp 1713338890
transform 1 0 384 0 1 50293
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_6
timestamp 1713338890
transform 1 0 904 0 1 51893
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_7
timestamp 1713338890
transform 1 0 9349 0 1 53493
box -180 -677 180 677
use M3_M2_CDNS_69033583165560  M3_M2_CDNS_69033583165560_8
timestamp 1713338890
transform 1 0 14580 0 1 55100
box -180 -677 180 677
use M3_M2_CDNS_69033583165561  M3_M2_CDNS_69033583165561_0
timestamp 1713338890
transform 1 0 84 0 1 37500
box -38 -677 38 677
use M3_M2_CDNS_69033583165561  M3_M2_CDNS_69033583165561_1
timestamp 1713338890
transform 1 0 3646 0 1 42293
box -38 -677 38 677
use M3_M2_CDNS_69033583165561  M3_M2_CDNS_69033583165561_2
timestamp 1713338890
transform 1 0 6087 0 1 37493
box -38 -677 38 677
use M3_M2_CDNS_69033583165561  M3_M2_CDNS_69033583165561_3
timestamp 1713338890
transform 1 0 14980 0 1 37493
box -38 -677 38 677
use M3_M2_CDNS_69033583165561  M3_M2_CDNS_69033583165561_4
timestamp 1713338890
transform 1 0 3646 0 1 43893
box -38 -677 38 677
use M3_M2_CDNS_69033583165561  M3_M2_CDNS_69033583165561_5
timestamp 1713338890
transform 1 0 84 0 1 51900
box -38 -677 38 677
use M3_M2_CDNS_69033583165561  M3_M2_CDNS_69033583165561_6
timestamp 1713338890
transform 1 0 1924 0 1 53493
box -38 -677 38 677
use M3_M2_CDNS_69033583165562  M3_M2_CDNS_69033583165562_0
timestamp 1713338890
transform 1 0 11668 0 1 49762
box -94 -150 94 150
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_0
timestamp 1713338890
transform 1 0 4788 0 1 53706
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_1
timestamp 1713338890
transform 1 0 6134 0 1 53706
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_2
timestamp 1713338890
transform 1 0 7480 0 1 53706
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_3
timestamp 1713338890
transform 1 0 10032 0 1 53706
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_4
timestamp 1713338890
transform 1 0 11378 0 1 53706
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_5
timestamp 1713338890
transform 1 0 12724 0 1 53706
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_6
timestamp 1713338890
transform 1 0 4788 0 1 55287
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_7
timestamp 1713338890
transform 1 0 6134 0 1 55287
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_8
timestamp 1713338890
transform 1 0 7480 0 1 55287
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_9
timestamp 1713338890
transform 1 0 10032 0 1 55287
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_10
timestamp 1713338890
transform 1 0 11378 0 1 55287
box -38 -464 38 464
use M3_M2_CDNS_69033583165564  M3_M2_CDNS_69033583165564_11
timestamp 1713338890
transform 1 0 12724 0 1 55287
box -38 -464 38 464
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_0
timestamp 1713338890
transform 1 0 4976 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_1
timestamp 1713338890
transform 1 0 5464 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_2
timestamp 1713338890
transform 1 0 5952 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_3
timestamp 1713338890
transform 1 0 6316 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_4
timestamp 1713338890
transform 1 0 6804 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_5
timestamp 1713338890
transform 1 0 7292 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_6
timestamp 1713338890
transform 1 0 10220 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_7
timestamp 1713338890
transform 1 0 10708 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_8
timestamp 1713338890
transform 1 0 11196 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_9
timestamp 1713338890
transform 1 0 11560 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_10
timestamp 1713338890
transform 1 0 12048 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_11
timestamp 1713338890
transform 1 0 12536 0 1 53716
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_12
timestamp 1713338890
transform 1 0 4976 0 1 55368
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_13
timestamp 1713338890
transform 1 0 5464 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_14
timestamp 1713338890
transform 1 0 5952 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_15
timestamp 1713338890
transform 1 0 6316 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_16
timestamp 1713338890
transform 1 0 6804 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_17
timestamp 1713338890
transform 1 0 7292 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_18
timestamp 1713338890
transform 1 0 10220 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_19
timestamp 1713338890
transform 1 0 11560 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_20
timestamp 1713338890
transform 1 0 10708 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_21
timestamp 1713338890
transform 1 0 11196 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_22
timestamp 1713338890
transform 1 0 12048 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165566  M3_M2_CDNS_69033583165566_23
timestamp 1713338890
transform 1 0 12536 0 1 55377
box -38 -393 38 393
use M3_M2_CDNS_69033583165573  M3_M2_CDNS_69033583165573_0
timestamp 1713338890
transform 1 0 1809 0 1 39448
box -38 -322 38 322
use M3_M2_CDNS_69033583165573  M3_M2_CDNS_69033583165573_1
timestamp 1713338890
transform 1 0 5121 0 1 39448
box -38 -322 38 322
use M3_M2_CDNS_69033583165573  M3_M2_CDNS_69033583165573_2
timestamp 1713338890
transform 1 0 7053 0 1 39448
box -38 -322 38 322
use M3_M2_CDNS_69033583165573  M3_M2_CDNS_69033583165573_3
timestamp 1713338890
transform 1 0 11039 0 1 47432
box -38 -322 38 322
use M3_M2_CDNS_69033583165576  M3_M2_CDNS_69033583165576_0
timestamp 1713338890
transform 1 0 11055 0 1 45474
box -38 -662 38 662
use M3_M2_CDNS_69033583165576  M3_M2_CDNS_69033583165576_1
timestamp 1713338890
transform 1 0 10926 0 1 45474
box -38 -662 38 662
use M3_M2_CDNS_69033583165577  M3_M2_CDNS_69033583165577_0
timestamp 1713338890
transform 1 0 10514 0 1 48008
box -90 -38 90 38
use M3_M2_CDNS_69033583165578  M3_M2_CDNS_69033583165578_0
timestamp 1713338890
transform 1 0 1006 0 1 31599
box -38 -1103 38 1103
use M3_M2_CDNS_69033583165578  M3_M2_CDNS_69033583165578_1
timestamp 1713338890
transform 1 0 2398 0 1 31599
box -38 -1103 38 1103
use M3_M2_CDNS_69033583165578  M3_M2_CDNS_69033583165578_2
timestamp 1713338890
transform 1 0 2814 0 1 31599
box -38 -1103 38 1103
use M3_M2_CDNS_69033583165578  M3_M2_CDNS_69033583165578_3
timestamp 1713338890
transform 1 0 7050 0 1 31599
box -38 -1103 38 1103
use M3_M2_CDNS_69033583165578  M3_M2_CDNS_69033583165578_4
timestamp 1713338890
transform 1 0 8014 0 1 31599
box -38 -1103 38 1103
use M3_M2_CDNS_69033583165578  M3_M2_CDNS_69033583165578_5
timestamp 1713338890
transform 1 0 12250 0 1 31599
box -38 -1103 38 1103
use M3_M2_CDNS_69033583165578  M3_M2_CDNS_69033583165578_6
timestamp 1713338890
transform 1 0 12666 0 1 31599
box -38 -1103 38 1103
use M3_M2_CDNS_69033583165578  M3_M2_CDNS_69033583165578_7
timestamp 1713338890
transform 1 0 14058 0 1 31599
box -38 -1103 38 1103
use M3_M2_CDNS_69033583165580  M3_M2_CDNS_69033583165580_0
timestamp 1713338890
transform 1 0 4028 0 1 34851
box -38 -1245 38 1245
use M3_M2_CDNS_69033583165580  M3_M2_CDNS_69033583165580_1
timestamp 1713338890
transform 1 0 11036 0 1 34851
box -38 -1245 38 1245
use M3_M2_CDNS_69033583165582  M3_M2_CDNS_69033583165582_0
timestamp 1713338890
transform 1 0 762 0 1 35244
box -38 -748 38 748
use M3_M2_CDNS_69033583165582  M3_M2_CDNS_69033583165582_1
timestamp 1713338890
transform 1 0 3130 0 1 35244
box -38 -748 38 748
use M3_M2_CDNS_69033583165582  M3_M2_CDNS_69033583165582_2
timestamp 1713338890
transform 1 0 4926 0 1 35244
box -38 -748 38 748
use M3_M2_CDNS_69033583165582  M3_M2_CDNS_69033583165582_3
timestamp 1713338890
transform 1 0 8709 0 1 35244
box -38 -748 38 748
use M3_M2_CDNS_69033583165582  M3_M2_CDNS_69033583165582_4
timestamp 1713338890
transform 1 0 10138 0 1 35244
box -38 -748 38 748
use M3_M2_CDNS_69033583165582  M3_M2_CDNS_69033583165582_5
timestamp 1713338890
transform 1 0 11934 0 1 35244
box -38 -748 38 748
use M3_M2_CDNS_69033583165583  M3_M2_CDNS_69033583165583_0
timestamp 1713338890
transform 1 0 524 0 1 35036
box -38 -961 38 961
use M3_M2_CDNS_69033583165583  M3_M2_CDNS_69033583165583_1
timestamp 1713338890
transform 1 0 4028 0 1 31954
box -38 -961 38 961
use M3_M2_CDNS_69033583165583  M3_M2_CDNS_69033583165583_2
timestamp 1713338890
transform 1 0 11036 0 1 31954
box -38 -961 38 961
use M3_M2_CDNS_69033583165585  M3_M2_CDNS_69033583165585_0
timestamp 1713338890
transform 1 0 8877 0 1 40288
box -890 -38 890 38
use M3_M2_CDNS_69033583165589  M3_M2_CDNS_69033583165589_0
timestamp 1713338890
transform 1 0 14580 0 1 19100
box -180 -1458 180 1458
use M3_M2_CDNS_69033583165589  M3_M2_CDNS_69033583165589_1
timestamp 1713338890
transform 1 0 14580 0 1 15900
box -180 -1458 180 1458
use M3_M2_CDNS_69033583165589  M3_M2_CDNS_69033583165589_2
timestamp 1713338890
transform 1 0 14580 0 1 22300
box -180 -1458 180 1458
use M3_M2_CDNS_69033583165589  M3_M2_CDNS_69033583165589_3
timestamp 1713338890
transform 1 0 14580 0 1 25500
box -180 -1458 180 1458
use M3_M2_CDNS_69033583165589  M3_M2_CDNS_69033583165589_4
timestamp 1713338890
transform 1 0 14580 0 1 31900
box -180 -1458 180 1458
use M3_M2_CDNS_69033583165590  M3_M2_CDNS_69033583165590_0
timestamp 1713338890
transform 1 0 274 0 1 27900
box -109 -677 109 677
use M3_M2_CDNS_69033583165590  M3_M2_CDNS_69033583165590_1
timestamp 1713338890
transform 1 0 12515 0 1 37493
box -109 -677 109 677
use M3_M2_CDNS_69033583165591  M3_M2_CDNS_69033583165591_0
timestamp 1713338890
transform 1 0 2662 0 1 30081
box -677 -38 677 38
use M3_M2_CDNS_69033583165591  M3_M2_CDNS_69033583165591_1
timestamp 1713338890
transform 1 0 12599 0 1 30081
box -677 -38 677 38
use M3_M2_CDNS_69033583165594  M3_M2_CDNS_69033583165594_0
timestamp 1713338890
transform 1 0 3460 0 1 40288
box -1103 -38 1103 38
use M3_M2_CDNS_69033583165600  M3_M2_CDNS_69033583165600_0
timestamp 1713338890
transform 1 0 14980 0 1 51893
box -38 -606 38 606
use M3_M2_CDNS_69033583165600  M3_M2_CDNS_69033583165600_1
timestamp 1713338890
transform 1 0 1924 0 1 56639
box -38 -606 38 606
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_0
timestamp 1713338890
transform 1 0 274 0 1 3100
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_1
timestamp 1713338890
transform 1 0 274 0 1 6300
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_2
timestamp 1713338890
transform 1 0 274 0 1 9500
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_3
timestamp 1713338890
transform 1 0 274 0 1 35100
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165606  M3_M2_CDNS_69033583165606_0
timestamp 1713338890
transform 1 0 524 0 1 31900
box -38 -1458 38 1458
use M3_M2_CDNS_69033583165607  M3_M2_CDNS_69033583165607_0
timestamp 1713338890
transform 1 0 2797 0 1 41044
box -961 -38 961 38
use nmoscap_6p0_CDNS_4066195314522  nmoscap_6p0_CDNS_4066195314522_0
timestamp 1713338890
transform 0 1 12482 1 0 42516
box -218 -350 818 692
use nmoscap_6p0_CDNS_4066195314522  nmoscap_6p0_CDNS_4066195314522_1
timestamp 1713338890
transform 0 1 12482 1 0 41548
box -218 -350 818 692
use nmoscap_6p0_CDNS_4066195314522  nmoscap_6p0_CDNS_4066195314522_2
timestamp 1713338890
transform 0 1 13622 1 0 42516
box -218 -350 818 692
use nmoscap_6p0_CDNS_4066195314522  nmoscap_6p0_CDNS_4066195314522_3
timestamp 1713338890
transform 0 1 13622 1 0 41548
box -218 -350 818 692
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_0
timestamp 1713338890
transform 0 1 7260 1 0 56489
box -218 -350 518 1092
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_1
timestamp 1713338890
transform 0 1 2760 1 0 56489
box -218 -350 518 1092
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_2
timestamp 1713338890
transform 0 1 5760 1 0 56489
box -218 -350 518 1092
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_3
timestamp 1713338890
transform 0 1 4260 1 0 56489
box -218 -350 518 1092
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_4
timestamp 1713338890
transform 0 1 10260 1 0 56489
box -218 -350 518 1092
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_5
timestamp 1713338890
transform 0 1 11760 1 0 56489
box -218 -350 518 1092
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_6
timestamp 1713338890
transform 0 1 13260 1 0 56489
box -218 -350 518 1092
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_7
timestamp 1713338890
transform 0 1 8760 1 0 56489
box -218 -350 518 1092
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_0
timestamp 1713338890
transform 1 0 11458 0 1 41627
box -216 -216 416 416
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_1
timestamp 1713338890
transform 1 0 11458 0 1 41163
box -216 -216 416 416
use ppolyf_u_CDNS_4066195314551  ppolyf_u_CDNS_4066195314551_0
timestamp 1713338890
transform 0 -1 1219 1 0 55401
box 0 0 984 160
use ppolyf_u_CDNS_4066195314551  ppolyf_u_CDNS_4066195314551_1
timestamp 1713338890
transform 0 -1 939 1 0 55401
box 0 0 984 160
<< labels >>
rlabel metal2 s 2136 57487 2136 57487 4 PD
port 1 nsew
rlabel metal2 s 7532 28487 7532 28487 4 PAD
port 2 nsew
rlabel metal2 s 1263 57483 1263 57483 4 PU
port 3 nsew
rlabel metal2 s 14242 57528 14242 57528 4 Y
port 4 nsew
rlabel metal2 s 1047 29559 1047 29559 4 ndrive_x_<0>
port 5 nsew
rlabel metal2 s 1231 29559 1231 29559 4 ndrive_y_<0>
port 6 nsew
rlabel metal2 s 1408 29559 1408 29559 4 ndrive_x_<1>
port 7 nsew
rlabel metal2 s 1594 29559 1594 29559 4 ndrive_Y_<1>
port 8 nsew
rlabel metal2 s 13463 29559 13463 29559 4 ndrive_x_<2>
port 9 nsew
rlabel metal2 s 13647 29559 13647 29559 4 ndrive_y_<2>
port 10 nsew
rlabel metal2 s 13824 29559 13824 29559 4 ndrive_x_<3>
port 11 nsew
rlabel metal2 s 14010 29559 14010 29559 4 ndrive_Y_<3>
port 12 nsew
rlabel metal2 s 3547 29559 3547 29559 4 pdrive_x_<0>
port 13 nsew
rlabel metal2 s 4188 29559 4188 29559 4 pdrive_y_<0>
port 14 nsew
rlabel metal2 s 4995 29559 4995 29559 4 pdrive_y_<1>
port 15 nsew
rlabel metal2 s 5954 29559 5954 29559 4 pdrive_x_<1>
port 16 nsew
rlabel metal2 s 9110 29559 9110 29559 4 pdrive_x_<2>
port 17 nsew
rlabel metal2 s 10062 29559 10062 29559 4 pdrive_y_<2>
port 18 nsew
rlabel metal2 s 10870 29559 10870 29559 4 pdrive_y_<3>
port 19 nsew
rlabel metal2 s 11512 29559 11512 29559 4 pdrive_x_<3>
port 20 nsew
<< end >>
