magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1073 -2666 1073 2666
<< metal1 >>
rect -73 1660 73 1666
rect -73 1634 -67 1660
rect -41 1634 -13 1660
rect 13 1634 41 1660
rect 67 1634 73 1660
rect -73 1606 73 1634
rect -73 1580 -67 1606
rect -41 1580 -13 1606
rect 13 1580 41 1606
rect 67 1580 73 1606
rect -73 1552 73 1580
rect -73 1526 -67 1552
rect -41 1526 -13 1552
rect 13 1526 41 1552
rect 67 1526 73 1552
rect -73 1498 73 1526
rect -73 1472 -67 1498
rect -41 1472 -13 1498
rect 13 1472 41 1498
rect 67 1472 73 1498
rect -73 1444 73 1472
rect -73 1418 -67 1444
rect -41 1418 -13 1444
rect 13 1418 41 1444
rect 67 1418 73 1444
rect -73 1390 73 1418
rect -73 1364 -67 1390
rect -41 1364 -13 1390
rect 13 1364 41 1390
rect 67 1364 73 1390
rect -73 1336 73 1364
rect -73 1310 -67 1336
rect -41 1310 -13 1336
rect 13 1310 41 1336
rect 67 1310 73 1336
rect -73 1282 73 1310
rect -73 1256 -67 1282
rect -41 1256 -13 1282
rect 13 1256 41 1282
rect 67 1256 73 1282
rect -73 1228 73 1256
rect -73 1202 -67 1228
rect -41 1202 -13 1228
rect 13 1202 41 1228
rect 67 1202 73 1228
rect -73 1174 73 1202
rect -73 1148 -67 1174
rect -41 1148 -13 1174
rect 13 1148 41 1174
rect 67 1148 73 1174
rect -73 1120 73 1148
rect -73 1094 -67 1120
rect -41 1094 -13 1120
rect 13 1094 41 1120
rect 67 1094 73 1120
rect -73 1066 73 1094
rect -73 1040 -67 1066
rect -41 1040 -13 1066
rect 13 1040 41 1066
rect 67 1040 73 1066
rect -73 1012 73 1040
rect -73 986 -67 1012
rect -41 986 -13 1012
rect 13 986 41 1012
rect 67 986 73 1012
rect -73 958 73 986
rect -73 932 -67 958
rect -41 932 -13 958
rect 13 932 41 958
rect 67 932 73 958
rect -73 904 73 932
rect -73 878 -67 904
rect -41 878 -13 904
rect 13 878 41 904
rect 67 878 73 904
rect -73 850 73 878
rect -73 824 -67 850
rect -41 824 -13 850
rect 13 824 41 850
rect 67 824 73 850
rect -73 796 73 824
rect -73 770 -67 796
rect -41 770 -13 796
rect 13 770 41 796
rect 67 770 73 796
rect -73 742 73 770
rect -73 716 -67 742
rect -41 716 -13 742
rect 13 716 41 742
rect 67 716 73 742
rect -73 688 73 716
rect -73 662 -67 688
rect -41 662 -13 688
rect 13 662 41 688
rect 67 662 73 688
rect -73 634 73 662
rect -73 608 -67 634
rect -41 608 -13 634
rect 13 608 41 634
rect 67 608 73 634
rect -73 580 73 608
rect -73 554 -67 580
rect -41 554 -13 580
rect 13 554 41 580
rect 67 554 73 580
rect -73 526 73 554
rect -73 500 -67 526
rect -41 500 -13 526
rect 13 500 41 526
rect 67 500 73 526
rect -73 472 73 500
rect -73 446 -67 472
rect -41 446 -13 472
rect 13 446 41 472
rect 67 446 73 472
rect -73 418 73 446
rect -73 392 -67 418
rect -41 392 -13 418
rect 13 392 41 418
rect 67 392 73 418
rect -73 364 73 392
rect -73 338 -67 364
rect -41 338 -13 364
rect 13 338 41 364
rect 67 338 73 364
rect -73 310 73 338
rect -73 284 -67 310
rect -41 284 -13 310
rect 13 284 41 310
rect 67 284 73 310
rect -73 256 73 284
rect -73 230 -67 256
rect -41 230 -13 256
rect 13 230 41 256
rect 67 230 73 256
rect -73 202 73 230
rect -73 176 -67 202
rect -41 176 -13 202
rect 13 176 41 202
rect 67 176 73 202
rect -73 148 73 176
rect -73 122 -67 148
rect -41 122 -13 148
rect 13 122 41 148
rect 67 122 73 148
rect -73 94 73 122
rect -73 68 -67 94
rect -41 68 -13 94
rect 13 68 41 94
rect 67 68 73 94
rect -73 40 73 68
rect -73 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 73 40
rect -73 -14 73 14
rect -73 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 73 -14
rect -73 -68 73 -40
rect -73 -94 -67 -68
rect -41 -94 -13 -68
rect 13 -94 41 -68
rect 67 -94 73 -68
rect -73 -122 73 -94
rect -73 -148 -67 -122
rect -41 -148 -13 -122
rect 13 -148 41 -122
rect 67 -148 73 -122
rect -73 -176 73 -148
rect -73 -202 -67 -176
rect -41 -202 -13 -176
rect 13 -202 41 -176
rect 67 -202 73 -176
rect -73 -230 73 -202
rect -73 -256 -67 -230
rect -41 -256 -13 -230
rect 13 -256 41 -230
rect 67 -256 73 -230
rect -73 -284 73 -256
rect -73 -310 -67 -284
rect -41 -310 -13 -284
rect 13 -310 41 -284
rect 67 -310 73 -284
rect -73 -338 73 -310
rect -73 -364 -67 -338
rect -41 -364 -13 -338
rect 13 -364 41 -338
rect 67 -364 73 -338
rect -73 -392 73 -364
rect -73 -418 -67 -392
rect -41 -418 -13 -392
rect 13 -418 41 -392
rect 67 -418 73 -392
rect -73 -446 73 -418
rect -73 -472 -67 -446
rect -41 -472 -13 -446
rect 13 -472 41 -446
rect 67 -472 73 -446
rect -73 -500 73 -472
rect -73 -526 -67 -500
rect -41 -526 -13 -500
rect 13 -526 41 -500
rect 67 -526 73 -500
rect -73 -554 73 -526
rect -73 -580 -67 -554
rect -41 -580 -13 -554
rect 13 -580 41 -554
rect 67 -580 73 -554
rect -73 -608 73 -580
rect -73 -634 -67 -608
rect -41 -634 -13 -608
rect 13 -634 41 -608
rect 67 -634 73 -608
rect -73 -662 73 -634
rect -73 -688 -67 -662
rect -41 -688 -13 -662
rect 13 -688 41 -662
rect 67 -688 73 -662
rect -73 -716 73 -688
rect -73 -742 -67 -716
rect -41 -742 -13 -716
rect 13 -742 41 -716
rect 67 -742 73 -716
rect -73 -770 73 -742
rect -73 -796 -67 -770
rect -41 -796 -13 -770
rect 13 -796 41 -770
rect 67 -796 73 -770
rect -73 -824 73 -796
rect -73 -850 -67 -824
rect -41 -850 -13 -824
rect 13 -850 41 -824
rect 67 -850 73 -824
rect -73 -878 73 -850
rect -73 -904 -67 -878
rect -41 -904 -13 -878
rect 13 -904 41 -878
rect 67 -904 73 -878
rect -73 -932 73 -904
rect -73 -958 -67 -932
rect -41 -958 -13 -932
rect 13 -958 41 -932
rect 67 -958 73 -932
rect -73 -986 73 -958
rect -73 -1012 -67 -986
rect -41 -1012 -13 -986
rect 13 -1012 41 -986
rect 67 -1012 73 -986
rect -73 -1040 73 -1012
rect -73 -1066 -67 -1040
rect -41 -1066 -13 -1040
rect 13 -1066 41 -1040
rect 67 -1066 73 -1040
rect -73 -1094 73 -1066
rect -73 -1120 -67 -1094
rect -41 -1120 -13 -1094
rect 13 -1120 41 -1094
rect 67 -1120 73 -1094
rect -73 -1148 73 -1120
rect -73 -1174 -67 -1148
rect -41 -1174 -13 -1148
rect 13 -1174 41 -1148
rect 67 -1174 73 -1148
rect -73 -1202 73 -1174
rect -73 -1228 -67 -1202
rect -41 -1228 -13 -1202
rect 13 -1228 41 -1202
rect 67 -1228 73 -1202
rect -73 -1256 73 -1228
rect -73 -1282 -67 -1256
rect -41 -1282 -13 -1256
rect 13 -1282 41 -1256
rect 67 -1282 73 -1256
rect -73 -1310 73 -1282
rect -73 -1336 -67 -1310
rect -41 -1336 -13 -1310
rect 13 -1336 41 -1310
rect 67 -1336 73 -1310
rect -73 -1364 73 -1336
rect -73 -1390 -67 -1364
rect -41 -1390 -13 -1364
rect 13 -1390 41 -1364
rect 67 -1390 73 -1364
rect -73 -1418 73 -1390
rect -73 -1444 -67 -1418
rect -41 -1444 -13 -1418
rect 13 -1444 41 -1418
rect 67 -1444 73 -1418
rect -73 -1472 73 -1444
rect -73 -1498 -67 -1472
rect -41 -1498 -13 -1472
rect 13 -1498 41 -1472
rect 67 -1498 73 -1472
rect -73 -1526 73 -1498
rect -73 -1552 -67 -1526
rect -41 -1552 -13 -1526
rect 13 -1552 41 -1526
rect 67 -1552 73 -1526
rect -73 -1580 73 -1552
rect -73 -1606 -67 -1580
rect -41 -1606 -13 -1580
rect 13 -1606 41 -1580
rect 67 -1606 73 -1580
rect -73 -1634 73 -1606
rect -73 -1660 -67 -1634
rect -41 -1660 -13 -1634
rect 13 -1660 41 -1634
rect 67 -1660 73 -1634
rect -73 -1666 73 -1660
<< via1 >>
rect -67 1634 -41 1660
rect -13 1634 13 1660
rect 41 1634 67 1660
rect -67 1580 -41 1606
rect -13 1580 13 1606
rect 41 1580 67 1606
rect -67 1526 -41 1552
rect -13 1526 13 1552
rect 41 1526 67 1552
rect -67 1472 -41 1498
rect -13 1472 13 1498
rect 41 1472 67 1498
rect -67 1418 -41 1444
rect -13 1418 13 1444
rect 41 1418 67 1444
rect -67 1364 -41 1390
rect -13 1364 13 1390
rect 41 1364 67 1390
rect -67 1310 -41 1336
rect -13 1310 13 1336
rect 41 1310 67 1336
rect -67 1256 -41 1282
rect -13 1256 13 1282
rect 41 1256 67 1282
rect -67 1202 -41 1228
rect -13 1202 13 1228
rect 41 1202 67 1228
rect -67 1148 -41 1174
rect -13 1148 13 1174
rect 41 1148 67 1174
rect -67 1094 -41 1120
rect -13 1094 13 1120
rect 41 1094 67 1120
rect -67 1040 -41 1066
rect -13 1040 13 1066
rect 41 1040 67 1066
rect -67 986 -41 1012
rect -13 986 13 1012
rect 41 986 67 1012
rect -67 932 -41 958
rect -13 932 13 958
rect 41 932 67 958
rect -67 878 -41 904
rect -13 878 13 904
rect 41 878 67 904
rect -67 824 -41 850
rect -13 824 13 850
rect 41 824 67 850
rect -67 770 -41 796
rect -13 770 13 796
rect 41 770 67 796
rect -67 716 -41 742
rect -13 716 13 742
rect 41 716 67 742
rect -67 662 -41 688
rect -13 662 13 688
rect 41 662 67 688
rect -67 608 -41 634
rect -13 608 13 634
rect 41 608 67 634
rect -67 554 -41 580
rect -13 554 13 580
rect 41 554 67 580
rect -67 500 -41 526
rect -13 500 13 526
rect 41 500 67 526
rect -67 446 -41 472
rect -13 446 13 472
rect 41 446 67 472
rect -67 392 -41 418
rect -13 392 13 418
rect 41 392 67 418
rect -67 338 -41 364
rect -13 338 13 364
rect 41 338 67 364
rect -67 284 -41 310
rect -13 284 13 310
rect 41 284 67 310
rect -67 230 -41 256
rect -13 230 13 256
rect 41 230 67 256
rect -67 176 -41 202
rect -13 176 13 202
rect 41 176 67 202
rect -67 122 -41 148
rect -13 122 13 148
rect 41 122 67 148
rect -67 68 -41 94
rect -13 68 13 94
rect 41 68 67 94
rect -67 14 -41 40
rect -13 14 13 40
rect 41 14 67 40
rect -67 -40 -41 -14
rect -13 -40 13 -14
rect 41 -40 67 -14
rect -67 -94 -41 -68
rect -13 -94 13 -68
rect 41 -94 67 -68
rect -67 -148 -41 -122
rect -13 -148 13 -122
rect 41 -148 67 -122
rect -67 -202 -41 -176
rect -13 -202 13 -176
rect 41 -202 67 -176
rect -67 -256 -41 -230
rect -13 -256 13 -230
rect 41 -256 67 -230
rect -67 -310 -41 -284
rect -13 -310 13 -284
rect 41 -310 67 -284
rect -67 -364 -41 -338
rect -13 -364 13 -338
rect 41 -364 67 -338
rect -67 -418 -41 -392
rect -13 -418 13 -392
rect 41 -418 67 -392
rect -67 -472 -41 -446
rect -13 -472 13 -446
rect 41 -472 67 -446
rect -67 -526 -41 -500
rect -13 -526 13 -500
rect 41 -526 67 -500
rect -67 -580 -41 -554
rect -13 -580 13 -554
rect 41 -580 67 -554
rect -67 -634 -41 -608
rect -13 -634 13 -608
rect 41 -634 67 -608
rect -67 -688 -41 -662
rect -13 -688 13 -662
rect 41 -688 67 -662
rect -67 -742 -41 -716
rect -13 -742 13 -716
rect 41 -742 67 -716
rect -67 -796 -41 -770
rect -13 -796 13 -770
rect 41 -796 67 -770
rect -67 -850 -41 -824
rect -13 -850 13 -824
rect 41 -850 67 -824
rect -67 -904 -41 -878
rect -13 -904 13 -878
rect 41 -904 67 -878
rect -67 -958 -41 -932
rect -13 -958 13 -932
rect 41 -958 67 -932
rect -67 -1012 -41 -986
rect -13 -1012 13 -986
rect 41 -1012 67 -986
rect -67 -1066 -41 -1040
rect -13 -1066 13 -1040
rect 41 -1066 67 -1040
rect -67 -1120 -41 -1094
rect -13 -1120 13 -1094
rect 41 -1120 67 -1094
rect -67 -1174 -41 -1148
rect -13 -1174 13 -1148
rect 41 -1174 67 -1148
rect -67 -1228 -41 -1202
rect -13 -1228 13 -1202
rect 41 -1228 67 -1202
rect -67 -1282 -41 -1256
rect -13 -1282 13 -1256
rect 41 -1282 67 -1256
rect -67 -1336 -41 -1310
rect -13 -1336 13 -1310
rect 41 -1336 67 -1310
rect -67 -1390 -41 -1364
rect -13 -1390 13 -1364
rect 41 -1390 67 -1364
rect -67 -1444 -41 -1418
rect -13 -1444 13 -1418
rect 41 -1444 67 -1418
rect -67 -1498 -41 -1472
rect -13 -1498 13 -1472
rect 41 -1498 67 -1472
rect -67 -1552 -41 -1526
rect -13 -1552 13 -1526
rect 41 -1552 67 -1526
rect -67 -1606 -41 -1580
rect -13 -1606 13 -1580
rect 41 -1606 67 -1580
rect -67 -1660 -41 -1634
rect -13 -1660 13 -1634
rect 41 -1660 67 -1634
<< metal2 >>
rect -73 1660 73 1666
rect -73 1634 -67 1660
rect -41 1634 -13 1660
rect 13 1634 41 1660
rect 67 1634 73 1660
rect -73 1606 73 1634
rect -73 1580 -67 1606
rect -41 1580 -13 1606
rect 13 1580 41 1606
rect 67 1580 73 1606
rect -73 1552 73 1580
rect -73 1526 -67 1552
rect -41 1526 -13 1552
rect 13 1526 41 1552
rect 67 1526 73 1552
rect -73 1498 73 1526
rect -73 1472 -67 1498
rect -41 1472 -13 1498
rect 13 1472 41 1498
rect 67 1472 73 1498
rect -73 1444 73 1472
rect -73 1418 -67 1444
rect -41 1418 -13 1444
rect 13 1418 41 1444
rect 67 1418 73 1444
rect -73 1390 73 1418
rect -73 1364 -67 1390
rect -41 1364 -13 1390
rect 13 1364 41 1390
rect 67 1364 73 1390
rect -73 1336 73 1364
rect -73 1310 -67 1336
rect -41 1310 -13 1336
rect 13 1310 41 1336
rect 67 1310 73 1336
rect -73 1282 73 1310
rect -73 1256 -67 1282
rect -41 1256 -13 1282
rect 13 1256 41 1282
rect 67 1256 73 1282
rect -73 1228 73 1256
rect -73 1202 -67 1228
rect -41 1202 -13 1228
rect 13 1202 41 1228
rect 67 1202 73 1228
rect -73 1174 73 1202
rect -73 1148 -67 1174
rect -41 1148 -13 1174
rect 13 1148 41 1174
rect 67 1148 73 1174
rect -73 1120 73 1148
rect -73 1094 -67 1120
rect -41 1094 -13 1120
rect 13 1094 41 1120
rect 67 1094 73 1120
rect -73 1066 73 1094
rect -73 1040 -67 1066
rect -41 1040 -13 1066
rect 13 1040 41 1066
rect 67 1040 73 1066
rect -73 1012 73 1040
rect -73 986 -67 1012
rect -41 986 -13 1012
rect 13 986 41 1012
rect 67 986 73 1012
rect -73 958 73 986
rect -73 932 -67 958
rect -41 932 -13 958
rect 13 932 41 958
rect 67 932 73 958
rect -73 904 73 932
rect -73 878 -67 904
rect -41 878 -13 904
rect 13 878 41 904
rect 67 878 73 904
rect -73 850 73 878
rect -73 824 -67 850
rect -41 824 -13 850
rect 13 824 41 850
rect 67 824 73 850
rect -73 796 73 824
rect -73 770 -67 796
rect -41 770 -13 796
rect 13 770 41 796
rect 67 770 73 796
rect -73 742 73 770
rect -73 716 -67 742
rect -41 716 -13 742
rect 13 716 41 742
rect 67 716 73 742
rect -73 688 73 716
rect -73 662 -67 688
rect -41 662 -13 688
rect 13 662 41 688
rect 67 662 73 688
rect -73 634 73 662
rect -73 608 -67 634
rect -41 608 -13 634
rect 13 608 41 634
rect 67 608 73 634
rect -73 580 73 608
rect -73 554 -67 580
rect -41 554 -13 580
rect 13 554 41 580
rect 67 554 73 580
rect -73 526 73 554
rect -73 500 -67 526
rect -41 500 -13 526
rect 13 500 41 526
rect 67 500 73 526
rect -73 472 73 500
rect -73 446 -67 472
rect -41 446 -13 472
rect 13 446 41 472
rect 67 446 73 472
rect -73 418 73 446
rect -73 392 -67 418
rect -41 392 -13 418
rect 13 392 41 418
rect 67 392 73 418
rect -73 364 73 392
rect -73 338 -67 364
rect -41 338 -13 364
rect 13 338 41 364
rect 67 338 73 364
rect -73 310 73 338
rect -73 284 -67 310
rect -41 284 -13 310
rect 13 284 41 310
rect 67 284 73 310
rect -73 256 73 284
rect -73 230 -67 256
rect -41 230 -13 256
rect 13 230 41 256
rect 67 230 73 256
rect -73 202 73 230
rect -73 176 -67 202
rect -41 176 -13 202
rect 13 176 41 202
rect 67 176 73 202
rect -73 148 73 176
rect -73 122 -67 148
rect -41 122 -13 148
rect 13 122 41 148
rect 67 122 73 148
rect -73 94 73 122
rect -73 68 -67 94
rect -41 68 -13 94
rect 13 68 41 94
rect 67 68 73 94
rect -73 40 73 68
rect -73 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 73 40
rect -73 -14 73 14
rect -73 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 73 -14
rect -73 -68 73 -40
rect -73 -94 -67 -68
rect -41 -94 -13 -68
rect 13 -94 41 -68
rect 67 -94 73 -68
rect -73 -122 73 -94
rect -73 -148 -67 -122
rect -41 -148 -13 -122
rect 13 -148 41 -122
rect 67 -148 73 -122
rect -73 -176 73 -148
rect -73 -202 -67 -176
rect -41 -202 -13 -176
rect 13 -202 41 -176
rect 67 -202 73 -176
rect -73 -230 73 -202
rect -73 -256 -67 -230
rect -41 -256 -13 -230
rect 13 -256 41 -230
rect 67 -256 73 -230
rect -73 -284 73 -256
rect -73 -310 -67 -284
rect -41 -310 -13 -284
rect 13 -310 41 -284
rect 67 -310 73 -284
rect -73 -338 73 -310
rect -73 -364 -67 -338
rect -41 -364 -13 -338
rect 13 -364 41 -338
rect 67 -364 73 -338
rect -73 -392 73 -364
rect -73 -418 -67 -392
rect -41 -418 -13 -392
rect 13 -418 41 -392
rect 67 -418 73 -392
rect -73 -446 73 -418
rect -73 -472 -67 -446
rect -41 -472 -13 -446
rect 13 -472 41 -446
rect 67 -472 73 -446
rect -73 -500 73 -472
rect -73 -526 -67 -500
rect -41 -526 -13 -500
rect 13 -526 41 -500
rect 67 -526 73 -500
rect -73 -554 73 -526
rect -73 -580 -67 -554
rect -41 -580 -13 -554
rect 13 -580 41 -554
rect 67 -580 73 -554
rect -73 -608 73 -580
rect -73 -634 -67 -608
rect -41 -634 -13 -608
rect 13 -634 41 -608
rect 67 -634 73 -608
rect -73 -662 73 -634
rect -73 -688 -67 -662
rect -41 -688 -13 -662
rect 13 -688 41 -662
rect 67 -688 73 -662
rect -73 -716 73 -688
rect -73 -742 -67 -716
rect -41 -742 -13 -716
rect 13 -742 41 -716
rect 67 -742 73 -716
rect -73 -770 73 -742
rect -73 -796 -67 -770
rect -41 -796 -13 -770
rect 13 -796 41 -770
rect 67 -796 73 -770
rect -73 -824 73 -796
rect -73 -850 -67 -824
rect -41 -850 -13 -824
rect 13 -850 41 -824
rect 67 -850 73 -824
rect -73 -878 73 -850
rect -73 -904 -67 -878
rect -41 -904 -13 -878
rect 13 -904 41 -878
rect 67 -904 73 -878
rect -73 -932 73 -904
rect -73 -958 -67 -932
rect -41 -958 -13 -932
rect 13 -958 41 -932
rect 67 -958 73 -932
rect -73 -986 73 -958
rect -73 -1012 -67 -986
rect -41 -1012 -13 -986
rect 13 -1012 41 -986
rect 67 -1012 73 -986
rect -73 -1040 73 -1012
rect -73 -1066 -67 -1040
rect -41 -1066 -13 -1040
rect 13 -1066 41 -1040
rect 67 -1066 73 -1040
rect -73 -1094 73 -1066
rect -73 -1120 -67 -1094
rect -41 -1120 -13 -1094
rect 13 -1120 41 -1094
rect 67 -1120 73 -1094
rect -73 -1148 73 -1120
rect -73 -1174 -67 -1148
rect -41 -1174 -13 -1148
rect 13 -1174 41 -1148
rect 67 -1174 73 -1148
rect -73 -1202 73 -1174
rect -73 -1228 -67 -1202
rect -41 -1228 -13 -1202
rect 13 -1228 41 -1202
rect 67 -1228 73 -1202
rect -73 -1256 73 -1228
rect -73 -1282 -67 -1256
rect -41 -1282 -13 -1256
rect 13 -1282 41 -1256
rect 67 -1282 73 -1256
rect -73 -1310 73 -1282
rect -73 -1336 -67 -1310
rect -41 -1336 -13 -1310
rect 13 -1336 41 -1310
rect 67 -1336 73 -1310
rect -73 -1364 73 -1336
rect -73 -1390 -67 -1364
rect -41 -1390 -13 -1364
rect 13 -1390 41 -1364
rect 67 -1390 73 -1364
rect -73 -1418 73 -1390
rect -73 -1444 -67 -1418
rect -41 -1444 -13 -1418
rect 13 -1444 41 -1418
rect 67 -1444 73 -1418
rect -73 -1472 73 -1444
rect -73 -1498 -67 -1472
rect -41 -1498 -13 -1472
rect 13 -1498 41 -1472
rect 67 -1498 73 -1472
rect -73 -1526 73 -1498
rect -73 -1552 -67 -1526
rect -41 -1552 -13 -1526
rect 13 -1552 41 -1526
rect 67 -1552 73 -1526
rect -73 -1580 73 -1552
rect -73 -1606 -67 -1580
rect -41 -1606 -13 -1580
rect 13 -1606 41 -1580
rect 67 -1606 73 -1580
rect -73 -1634 73 -1606
rect -73 -1660 -67 -1634
rect -41 -1660 -13 -1634
rect 13 -1660 41 -1634
rect 67 -1660 73 -1634
rect -73 -1666 73 -1660
<< end >>
