magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2407 -2051 15369 49415
<< nwell >>
rect 2170 27627 10792 29165
<< psubdiff >>
rect 2253 25802 2343 25866
rect 10619 25802 10709 25866
rect 2253 25780 10709 25802
rect 2253 25734 2275 25780
rect 6739 25734 6975 25780
rect 7209 25734 7445 25780
rect 7679 25734 8009 25780
rect 10687 25734 10709 25780
rect 2253 25712 10709 25734
<< psubdiffcont >>
rect 2275 25734 6739 25780
rect 6975 25734 7209 25780
rect 7445 25734 7679 25780
rect 8009 25734 10687 25780
<< polysilicon >>
rect 2665 27601 2805 27745
rect 2909 27601 3049 27745
rect 3153 27601 3293 27745
rect 3397 27601 3537 27745
rect 2665 27517 3537 27601
rect 3641 27601 3781 27745
rect 3885 27601 4025 27745
rect 4129 27601 4269 27745
rect 3641 27517 4269 27601
rect 4545 27601 4685 27745
rect 4789 27601 4929 27745
rect 5033 27601 5173 27745
rect 4545 27517 5173 27601
rect 5277 27601 5417 27745
rect 5521 27601 5661 27745
rect 5765 27601 5905 27745
rect 5277 27517 5905 27601
rect 6009 27601 6149 27745
rect 6253 27601 6393 27745
rect 6497 27601 6637 27745
rect 6009 27517 6637 27601
rect 6741 27601 6881 27745
rect 6985 27601 7125 27745
rect 7229 27601 7369 27745
rect 6741 27517 7369 27601
rect 7473 27601 7613 27745
rect 7717 27601 7857 27745
rect 7961 27601 8101 27745
rect 7473 27517 8101 27601
rect 8205 27601 8345 27745
rect 8449 27601 8589 27745
rect 8693 27601 8833 27745
rect 8205 27517 8833 27601
rect 8937 27601 9077 27745
rect 9181 27601 9321 27745
rect 9425 27601 9565 27745
rect 8937 27517 9565 27601
rect 9669 27601 9809 27745
rect 9913 27601 10053 27745
rect 10157 27601 10297 27745
rect 9669 27517 10297 27601
rect 5191 27194 5819 27278
rect 4129 27050 4269 27150
rect 5191 27050 5331 27194
rect 5435 27050 5575 27194
rect 5679 27050 5819 27194
rect 5923 27194 6551 27278
rect 5923 27050 6063 27194
rect 6167 27050 6307 27194
rect 6411 27050 6551 27194
rect 6655 27194 7283 27278
rect 6655 27050 6795 27194
rect 6899 27050 7039 27194
rect 7143 27050 7283 27194
rect 7387 27194 8015 27278
rect 7387 27050 7527 27194
rect 7631 27050 7771 27194
rect 7875 27050 8015 27194
<< metal1 >>
rect -1 27593 67 30038
rect 2264 28917 2332 29003
rect 2575 27789 2651 29071
rect 2819 27729 2895 28789
rect 3063 27789 3139 29071
rect 3307 27729 3383 28789
rect 3551 27789 3627 29071
rect 3795 27729 3871 28789
rect 4039 27789 4115 29071
rect 4283 27729 4359 28789
rect 4455 27789 4531 29071
rect 2819 27653 3627 27729
rect 3795 27653 4359 27729
rect 4699 27729 4775 28789
rect 4943 27789 5019 29071
rect 5187 27729 5263 28789
rect 5431 27789 5507 29071
rect 5675 27729 5751 28789
rect 5919 27789 5995 29071
rect 6163 27729 6239 28789
rect 6407 27789 6483 29071
rect 6651 27729 6727 28789
rect 6895 27789 6971 29071
rect 7139 27729 7215 28789
rect 7383 27789 7459 29071
rect 7627 27729 7703 28789
rect 7871 27789 7947 29071
rect 8115 27729 8191 28789
rect 8359 27789 8435 29071
rect 8603 27729 8679 28789
rect 8847 27789 8923 29071
rect 9091 27729 9167 28789
rect 9335 27789 9411 29071
rect 9579 27729 9655 28789
rect 9823 27789 9899 29071
rect 10067 27729 10143 28789
rect 10311 27789 10387 29071
rect 10630 28917 10698 29003
rect 4699 27653 10433 27729
rect 3551 27597 3627 27653
rect -1 27393 3464 27593
rect 3388 27146 3464 27393
rect 3551 27521 4224 27597
rect 4283 27593 4359 27653
rect 3551 27274 3627 27521
rect 4283 27517 10275 27593
rect 3551 27198 6516 27274
rect 3388 27070 4223 27146
rect 2264 25791 2332 25877
rect 4039 25791 4115 27006
rect 4283 26006 4359 27198
rect 6652 27142 6728 27517
rect 10357 27142 10433 27653
rect 5345 27066 6728 27142
rect 6809 27066 10433 27142
rect 5101 25791 5177 27006
rect 5345 26006 5421 27066
rect 5589 25791 5665 27006
rect 5833 26006 5909 27066
rect 6077 25791 6153 27006
rect 6321 26006 6397 27066
rect 6565 25791 6641 27006
rect 2264 25780 6759 25791
rect 2264 25734 2275 25780
rect 6739 25734 6759 25780
rect 2264 25723 6759 25734
rect 6809 25617 6885 27066
rect 7053 25791 7129 27006
rect 7297 25979 7373 27066
rect 7541 25791 7617 27006
rect 7785 25979 7861 27066
rect 8029 25791 8105 27006
rect 10630 25791 10698 25877
rect 6935 25780 7247 25791
rect 6935 25734 6975 25780
rect 7209 25734 7247 25780
rect 6935 25723 7247 25734
rect 7423 25780 7735 25791
rect 7423 25734 7445 25780
rect 7679 25734 7735 25780
rect 7423 25723 7735 25734
rect 7911 25780 10698 25791
rect 7911 25734 8009 25780
rect 10687 25734 10698 25780
rect 7911 25723 10698 25734
rect 1213 25417 11749 25617
use comp018green_esd_rc_v5p0  comp018green_esd_rc_v5p0_0
timestamp 1713338890
transform 1 0 -356 0 -1 46507
box -51 491 13725 17038
use M1_NWELL_CDNS_40661953145107  M1_NWELL_CDNS_40661953145107_0
timestamp 1713338890
transform 1 0 6481 0 1 29037
box -4311 -128 4311 128
use M1_NWELL_CDNS_40661953145111  M1_NWELL_CDNS_40661953145111_0
timestamp 1713338890
transform 1 0 2298 0 1 28319
box -128 -692 128 692
use M1_NWELL_CDNS_40661953145111  M1_NWELL_CDNS_40661953145111_1
timestamp 1713338890
transform 1 0 10664 0 1 28319
box -128 -692 128 692
use M1_POLY2_CDNS_69033583165343  M1_POLY2_CDNS_69033583165343_0
timestamp 1713338890
transform 1 0 7421 0 1 27559
box -2862 -42 2862 42
use M1_POLY2_CDNS_69033583165344  M1_POLY2_CDNS_69033583165344_0
timestamp 1713338890
transform 1 0 5871 0 1 27236
box -653 -42 653 42
use M1_POLY2_CDNS_69033583165344  M1_POLY2_CDNS_69033583165344_1
timestamp 1713338890
transform 1 0 7335 0 1 27236
box -653 -42 653 42
use M1_POLY2_CDNS_69033583165345  M1_POLY2_CDNS_69033583165345_0
timestamp 1713338890
transform 1 0 3955 0 1 27559
box -277 -42 277 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_0
timestamp 1713338890
transform 1 0 4142 0 1 27108
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165347  M1_POLY2_CDNS_69033583165347_0
timestamp 1713338890
transform 1 0 3101 0 1 27559
box -371 -42 371 42
use M1_PSUB_CDNS_69033583165349  M1_PSUB_CDNS_69033583165349_0
timestamp 1713338890
transform 1 0 2298 0 -1 26522
box -45 -656 45 656
use M1_PSUB_CDNS_69033583165349  M1_PSUB_CDNS_69033583165349_1
timestamp 1713338890
transform 1 0 10664 0 -1 26522
box -45 -656 45 656
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_0
timestamp 1713338890
transform 1 0 1313 0 1 25517
box -92 -92 92 92
use M2_M1_CDNS_69033583165348  M2_M1_CDNS_69033583165348_1
timestamp 1713338890
transform 1 0 11649 0 1 25517
box -92 -92 92 92
use nmos_6p0_CDNS_406619531458  nmos_6p0_CDNS_406619531458_0
timestamp 1713338890
transform 1 0 5191 0 1 26006
box -88 -44 1448 1044
use nmos_6p0_CDNS_406619531458  nmos_6p0_CDNS_406619531458_1
timestamp 1713338890
transform 1 0 6655 0 1 26006
box -88 -44 1448 1044
use nmos_6p0_CDNS_406619531459  nmos_6p0_CDNS_406619531459_0
timestamp 1713338890
transform 1 0 4129 0 1 26006
box -88 -44 228 1044
use nmos_clamp_20_50_4  nmos_clamp_20_50_4_0
timestamp 1713338890
transform 1 0 0 0 1 0
box -51 -51 13013 25617
use pmos_6p0_CDNS_406619531452  pmos_6p0_CDNS_406619531452_0
timestamp 1713338890
transform 1 0 2665 0 1 27789
box -208 -120 1080 1120
use pmos_6p0_CDNS_406619531455  pmos_6p0_CDNS_406619531455_0
timestamp 1713338890
transform 1 0 4545 0 1 27789
box -208 -120 5960 1120
use pmos_6p0_CDNS_406619531456  pmos_6p0_CDNS_406619531456_0
timestamp 1713338890
transform 1 0 3641 0 1 27789
box -208 -120 836 1120
use top_route_1  top_route_1_0
timestamp 1713338890
transform 1 0 43 0 1 25617
box 0 0 12876 21798
<< end >>
