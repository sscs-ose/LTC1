magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -564 -3269 8904 3605
<< nwell >>
rect 1846 1263 2990 1605
rect 1846 1262 3249 1263
rect 1846 1261 6517 1262
rect 1846 -1140 6904 1261
rect 1846 -1142 3249 -1140
rect 6505 -1141 6904 -1140
rect 1846 -1269 2990 -1142
<< pmos >>
rect 6413 166 6581 266
rect 6413 -243 6581 -146
rect 6415 -656 6583 -556
rect 2256 -994 2356 -826
rect 2620 -998 2720 -830
<< pdiff >>
rect 6325 239 6413 266
rect 6325 193 6338 239
rect 6384 193 6413 239
rect 6325 166 6413 193
rect 6581 239 6669 266
rect 6581 193 6610 239
rect 6656 193 6669 239
rect 6581 166 6669 193
rect 6336 -173 6413 -146
rect 6336 -219 6338 -173
rect 6384 -219 6413 -173
rect 6336 -243 6413 -219
rect 6581 -173 6661 -146
rect 6581 -219 6610 -173
rect 6656 -219 6661 -173
rect 6581 -243 6661 -219
rect 6327 -583 6415 -556
rect 6327 -629 6340 -583
rect 6386 -629 6415 -583
rect 6327 -656 6415 -629
rect 6583 -583 6671 -556
rect 6583 -629 6612 -583
rect 6658 -629 6671 -583
rect 6583 -656 6671 -629
rect 2256 -751 2356 -738
rect 2256 -797 2283 -751
rect 2329 -797 2356 -751
rect 2256 -826 2356 -797
rect 2620 -755 2720 -742
rect 2620 -801 2647 -755
rect 2693 -801 2720 -755
rect 2620 -830 2720 -801
rect 2256 -1023 2356 -994
rect 2256 -1069 2283 -1023
rect 2329 -1069 2356 -1023
rect 2256 -1082 2356 -1069
rect 2620 -1027 2720 -998
rect 2620 -1073 2647 -1027
rect 2693 -1073 2720 -1027
rect 2620 -1086 2720 -1073
<< pdiffc >>
rect 6338 193 6384 239
rect 6610 193 6656 239
rect 6338 -219 6384 -173
rect 6610 -219 6656 -173
rect 6340 -629 6386 -583
rect 6612 -629 6658 -583
rect 2283 -797 2329 -751
rect 2647 -801 2693 -755
rect 2283 -1069 2329 -1023
rect 2647 -1073 2693 -1027
<< nsubdiff >>
rect 1877 1547 2941 1568
rect 1877 1501 1902 1547
rect 1948 1501 2022 1547
rect 2068 1501 2142 1547
rect 2188 1501 2262 1547
rect 2308 1501 2382 1547
rect 2428 1501 2502 1547
rect 2548 1501 2622 1547
rect 2668 1501 2742 1547
rect 2788 1501 2941 1547
rect 1877 1480 2941 1501
rect 1877 1006 1965 1480
rect 2846 1465 2941 1480
rect 2846 1419 2869 1465
rect 2915 1419 2941 1465
rect 2846 1326 2941 1419
rect 2846 1280 2869 1326
rect 2915 1280 2941 1326
rect 2846 1167 2941 1280
rect 2846 1142 6859 1167
rect 2846 1096 2869 1142
rect 2915 1096 3038 1142
rect 3084 1096 3207 1142
rect 3253 1096 3407 1142
rect 3453 1096 3526 1142
rect 3572 1096 3645 1142
rect 3691 1096 3764 1142
rect 3810 1096 3883 1142
rect 3929 1096 4002 1142
rect 4048 1096 4121 1142
rect 4167 1096 4240 1142
rect 4286 1096 4359 1142
rect 4405 1096 4478 1142
rect 4524 1096 4597 1142
rect 4643 1096 4716 1142
rect 4762 1096 4835 1142
rect 4881 1096 4954 1142
rect 5000 1096 5073 1142
rect 5119 1096 5192 1142
rect 5238 1096 5311 1142
rect 5357 1096 5430 1142
rect 5476 1096 5549 1142
rect 5595 1096 5668 1142
rect 5714 1096 5787 1142
rect 5833 1096 5906 1142
rect 5952 1096 6025 1142
rect 6071 1096 6144 1142
rect 6190 1096 6263 1142
rect 6309 1141 6859 1142
rect 6309 1096 6403 1141
rect 2846 1095 6403 1096
rect 6449 1095 6561 1141
rect 6607 1095 6859 1141
rect 2846 1072 6859 1095
rect 1877 960 1897 1006
rect 1943 960 1965 1006
rect 1877 883 1965 960
rect 1877 837 1897 883
rect 1943 837 1965 883
rect 2937 996 3031 1072
rect 2937 950 2961 996
rect 3007 950 3031 996
rect 2937 887 3031 950
rect 1877 769 1965 837
rect 1877 723 1897 769
rect 1943 723 1965 769
rect 1877 646 1965 723
rect 2937 841 2961 887
rect 3007 841 3031 887
rect 2937 778 3031 841
rect 6752 1034 6859 1072
rect 6752 988 6774 1034
rect 6820 988 6859 1034
rect 6752 915 6859 988
rect 6752 869 6774 915
rect 6820 869 6859 915
rect 2937 732 2961 778
rect 3007 732 3031 778
rect 1877 600 1897 646
rect 1943 600 1965 646
rect 2937 647 3031 732
rect 6752 796 6859 869
rect 6752 750 6774 796
rect 6820 750 6859 796
rect 6752 677 6859 750
rect 1877 529 1965 600
rect 1877 483 1897 529
rect 1943 483 1965 529
rect 1877 406 1965 483
rect 1877 360 1897 406
rect 1943 360 1965 406
rect 1877 289 1965 360
rect 1877 243 1897 289
rect 1943 243 1965 289
rect 1877 166 1965 243
rect 1877 120 1897 166
rect 1943 120 1965 166
rect 2937 601 2961 647
rect 3007 601 3031 647
rect 2937 517 3031 601
rect 6752 631 6774 677
rect 6820 631 6859 677
rect 6752 558 6859 631
rect 2937 471 2961 517
rect 3007 471 3031 517
rect 2937 386 3031 471
rect 6752 512 6774 558
rect 6820 512 6859 558
rect 6752 439 6859 512
rect 6752 393 6774 439
rect 6820 393 6859 439
rect 2937 340 2961 386
rect 3007 340 3031 386
rect 2937 255 3031 340
rect 6752 320 6859 393
rect 6752 274 6774 320
rect 6820 274 6859 320
rect 2937 209 2961 255
rect 3007 209 3031 255
rect 1877 49 1965 120
rect 2937 125 3031 209
rect 6752 201 6859 274
rect 2937 79 2961 125
rect 3007 79 3031 125
rect 1877 3 1897 49
rect 1943 3 1965 49
rect 1877 -74 1965 3
rect 1877 -120 1897 -74
rect 1943 -120 1965 -74
rect 2937 16 3031 79
rect 6752 155 6774 201
rect 6820 155 6859 201
rect 6752 82 6859 155
rect 2937 -30 2961 16
rect 3007 -30 3031 16
rect 6752 36 6774 82
rect 6820 36 6859 82
rect 2937 -93 3031 -30
rect 1877 -191 1965 -120
rect 1877 -237 1897 -191
rect 1943 -237 1965 -191
rect 1877 -314 1965 -237
rect 1877 -360 1897 -314
rect 1943 -360 1965 -314
rect 2937 -139 2961 -93
rect 3007 -139 3031 -93
rect 2937 -245 3031 -139
rect 6752 -37 6859 36
rect 6752 -83 6774 -37
rect 6820 -83 6859 -37
rect 6752 -156 6859 -83
rect 6752 -202 6774 -156
rect 6820 -202 6859 -156
rect 2937 -291 2961 -245
rect 3007 -291 3031 -245
rect 1877 -431 1965 -360
rect 1877 -477 1897 -431
rect 1943 -477 1965 -431
rect 1877 -554 1965 -477
rect 2937 -398 3031 -291
rect 6752 -275 6859 -202
rect 6752 -321 6774 -275
rect 6820 -321 6859 -275
rect 2937 -444 2961 -398
rect 3007 -444 3031 -398
rect 6752 -394 6859 -321
rect 1877 -600 1897 -554
rect 1943 -600 1965 -554
rect 1877 -681 1965 -600
rect 1877 -727 1897 -681
rect 1943 -727 1965 -681
rect 1877 -1157 1965 -727
rect 2937 -572 3031 -444
rect 6752 -440 6774 -394
rect 6820 -440 6859 -394
rect 6752 -513 6859 -440
rect 2937 -618 2961 -572
rect 3007 -618 3031 -572
rect 2937 -702 3031 -618
rect 6752 -559 6774 -513
rect 6820 -559 6859 -513
rect 6752 -632 6859 -559
rect 2937 -748 2961 -702
rect 3007 -748 3031 -702
rect 2937 -811 3031 -748
rect 6752 -678 6774 -632
rect 6820 -678 6859 -632
rect 6752 -751 6859 -678
rect 2937 -857 2961 -811
rect 3007 -857 3031 -811
rect 2937 -882 3031 -857
rect 2823 -901 3031 -882
rect 6752 -797 6774 -751
rect 6820 -797 6859 -751
rect 6752 -901 6859 -797
rect 2823 -924 6859 -901
rect 2823 -927 3416 -924
rect 2823 -973 3112 -927
rect 3158 -973 3282 -927
rect 3328 -970 3416 -927
rect 3462 -970 3535 -924
rect 3581 -970 3654 -924
rect 3700 -970 3773 -924
rect 3819 -970 3892 -924
rect 3938 -970 4011 -924
rect 4057 -970 4130 -924
rect 4176 -970 4249 -924
rect 4295 -970 4368 -924
rect 4414 -970 4487 -924
rect 4533 -970 4606 -924
rect 4652 -970 4725 -924
rect 4771 -970 4844 -924
rect 4890 -970 4963 -924
rect 5009 -970 5082 -924
rect 5128 -970 5201 -924
rect 5247 -970 5320 -924
rect 5366 -970 5439 -924
rect 5485 -970 5558 -924
rect 5604 -970 5677 -924
rect 5723 -970 5796 -924
rect 5842 -970 5915 -924
rect 5961 -970 6034 -924
rect 6080 -970 6153 -924
rect 6199 -970 6272 -924
rect 6318 -970 6423 -924
rect 6469 -970 6567 -924
rect 6613 -970 6791 -924
rect 6837 -970 6859 -924
rect 3328 -973 6859 -970
rect 2823 -993 6859 -973
rect 2823 -1157 2895 -993
rect 1877 -1178 2895 -1157
rect 1877 -1224 1902 -1178
rect 1948 -1224 2022 -1178
rect 2068 -1224 2142 -1178
rect 2188 -1224 2262 -1178
rect 2308 -1224 2382 -1178
rect 2428 -1224 2502 -1178
rect 2548 -1224 2622 -1178
rect 2668 -1224 2742 -1178
rect 2788 -1224 2895 -1178
rect 1877 -1245 2895 -1224
<< nsubdiffcont >>
rect 1902 1501 1948 1547
rect 2022 1501 2068 1547
rect 2142 1501 2188 1547
rect 2262 1501 2308 1547
rect 2382 1501 2428 1547
rect 2502 1501 2548 1547
rect 2622 1501 2668 1547
rect 2742 1501 2788 1547
rect 2869 1419 2915 1465
rect 2869 1280 2915 1326
rect 2869 1096 2915 1142
rect 3038 1096 3084 1142
rect 3207 1096 3253 1142
rect 3407 1096 3453 1142
rect 3526 1096 3572 1142
rect 3645 1096 3691 1142
rect 3764 1096 3810 1142
rect 3883 1096 3929 1142
rect 4002 1096 4048 1142
rect 4121 1096 4167 1142
rect 4240 1096 4286 1142
rect 4359 1096 4405 1142
rect 4478 1096 4524 1142
rect 4597 1096 4643 1142
rect 4716 1096 4762 1142
rect 4835 1096 4881 1142
rect 4954 1096 5000 1142
rect 5073 1096 5119 1142
rect 5192 1096 5238 1142
rect 5311 1096 5357 1142
rect 5430 1096 5476 1142
rect 5549 1096 5595 1142
rect 5668 1096 5714 1142
rect 5787 1096 5833 1142
rect 5906 1096 5952 1142
rect 6025 1096 6071 1142
rect 6144 1096 6190 1142
rect 6263 1096 6309 1142
rect 6403 1095 6449 1141
rect 6561 1095 6607 1141
rect 1897 960 1943 1006
rect 1897 837 1943 883
rect 2961 950 3007 996
rect 1897 723 1943 769
rect 2961 841 3007 887
rect 6774 988 6820 1034
rect 6774 869 6820 915
rect 2961 732 3007 778
rect 1897 600 1943 646
rect 6774 750 6820 796
rect 1897 483 1943 529
rect 1897 360 1943 406
rect 1897 243 1943 289
rect 1897 120 1943 166
rect 2961 601 3007 647
rect 6774 631 6820 677
rect 2961 471 3007 517
rect 6774 512 6820 558
rect 6774 393 6820 439
rect 2961 340 3007 386
rect 6774 274 6820 320
rect 2961 209 3007 255
rect 2961 79 3007 125
rect 1897 3 1943 49
rect 1897 -120 1943 -74
rect 6774 155 6820 201
rect 2961 -30 3007 16
rect 6774 36 6820 82
rect 1897 -237 1943 -191
rect 1897 -360 1943 -314
rect 2961 -139 3007 -93
rect 6774 -83 6820 -37
rect 6774 -202 6820 -156
rect 2961 -291 3007 -245
rect 1897 -477 1943 -431
rect 6774 -321 6820 -275
rect 2961 -444 3007 -398
rect 1897 -600 1943 -554
rect 1897 -727 1943 -681
rect 6774 -440 6820 -394
rect 2961 -618 3007 -572
rect 6774 -559 6820 -513
rect 2961 -748 3007 -702
rect 6774 -678 6820 -632
rect 2961 -857 3007 -811
rect 6774 -797 6820 -751
rect 3112 -973 3158 -927
rect 3282 -973 3328 -927
rect 3416 -970 3462 -924
rect 3535 -970 3581 -924
rect 3654 -970 3700 -924
rect 3773 -970 3819 -924
rect 3892 -970 3938 -924
rect 4011 -970 4057 -924
rect 4130 -970 4176 -924
rect 4249 -970 4295 -924
rect 4368 -970 4414 -924
rect 4487 -970 4533 -924
rect 4606 -970 4652 -924
rect 4725 -970 4771 -924
rect 4844 -970 4890 -924
rect 4963 -970 5009 -924
rect 5082 -970 5128 -924
rect 5201 -970 5247 -924
rect 5320 -970 5366 -924
rect 5439 -970 5485 -924
rect 5558 -970 5604 -924
rect 5677 -970 5723 -924
rect 5796 -970 5842 -924
rect 5915 -970 5961 -924
rect 6034 -970 6080 -924
rect 6153 -970 6199 -924
rect 6272 -970 6318 -924
rect 6423 -970 6469 -924
rect 6567 -970 6613 -924
rect 6791 -970 6837 -924
rect 1902 -1224 1948 -1178
rect 2022 -1224 2068 -1178
rect 2142 -1224 2188 -1178
rect 2262 -1224 2308 -1178
rect 2382 -1224 2428 -1178
rect 2502 -1224 2548 -1178
rect 2622 -1224 2668 -1178
rect 2742 -1224 2788 -1178
<< polysilicon >>
rect 2141 1242 2234 1306
rect 2141 1196 2169 1242
rect 2215 1196 2234 1242
rect 2141 1137 2234 1196
rect 2502 1305 2595 1306
rect 2502 1242 2620 1305
rect 2502 1196 2530 1242
rect 2576 1196 2620 1242
rect 2502 1137 2620 1196
rect 2720 1137 2764 1305
rect 2403 820 2461 876
rect 2448 774 2461 820
rect 2763 813 2813 876
rect 2719 794 2737 799
rect 2740 794 2745 799
rect 2403 708 2461 774
rect 2798 767 2813 813
rect 2763 708 2813 767
rect 3194 771 3362 799
rect 3194 736 3253 771
rect 3197 725 3253 736
rect 3299 725 3362 771
rect 3197 673 3362 725
rect 3713 754 3881 769
rect 3713 718 3769 754
rect 3815 718 3881 754
rect 4529 753 4697 771
rect 4529 718 4584 753
rect 3769 707 3815 708
rect 4573 707 4584 718
rect 4630 718 4697 753
rect 5317 753 5485 777
rect 4630 707 4641 718
rect 3785 674 3793 705
rect 4573 675 4641 707
rect 5317 707 5392 753
rect 5438 707 5485 753
rect 5317 703 5485 707
rect 5589 753 5757 777
rect 5589 707 5654 753
rect 5700 707 5757 753
rect 5589 703 5757 707
rect 6413 774 6581 802
rect 6413 728 6472 774
rect 6518 728 6581 774
rect 6413 690 6581 728
rect 2159 543 2217 604
rect 2524 546 2575 604
rect 2159 497 2180 543
rect 2226 535 2261 540
rect 2524 500 2540 546
rect 2586 526 2619 530
rect 3197 530 3362 573
rect 2159 164 2217 497
rect 2524 436 2575 500
rect 2524 164 2598 436
rect 3985 527 4153 537
rect 3985 481 4039 527
rect 4085 481 4153 527
rect 3985 463 4153 481
rect 4257 527 4425 537
rect 4257 481 4316 527
rect 4362 481 4425 527
rect 4257 463 4425 481
rect 5045 527 5213 530
rect 5045 481 5119 527
rect 5165 481 5213 527
rect 5045 465 5213 481
rect 5861 527 6030 530
rect 5861 481 5939 527
rect 5985 481 6030 527
rect 5861 468 6030 481
rect 3191 356 3359 384
rect 3191 321 3250 356
rect 3193 310 3250 321
rect 3296 310 3359 356
rect 3193 258 3359 310
rect 3713 344 3881 361
rect 3713 308 3786 344
rect 3832 308 3881 344
rect 4529 349 4697 364
rect 4529 308 4587 349
rect 4633 308 4697 349
rect 5317 349 5485 371
rect 4587 302 4633 303
rect 5317 303 5372 349
rect 5418 303 5485 349
rect 3786 297 3832 298
rect 5317 297 5485 303
rect 5589 353 5757 371
rect 5589 307 5652 353
rect 5698 307 5757 353
rect 5589 297 5757 307
rect 6413 364 6581 392
rect 6413 318 6472 364
rect 6518 318 6581 364
rect 6413 266 6581 318
rect 3194 116 3359 158
rect 3985 131 4153 141
rect 2403 9 2477 60
rect 2445 -37 2477 9
rect 2403 -108 2477 -37
rect 2719 -2 2813 60
rect 2719 -48 2752 -2
rect 2798 -48 2813 -2
rect 2719 -108 2813 -48
rect 3985 85 4044 131
rect 4090 85 4153 131
rect 3985 67 4153 85
rect 4257 131 4425 141
rect 4257 85 4321 131
rect 4367 85 4425 131
rect 4257 67 4425 85
rect 5045 84 5098 121
rect 5144 84 5213 121
rect 5045 57 5213 84
rect 5861 85 5931 121
rect 6413 122 6581 166
rect 5977 85 6029 121
rect 5861 65 6029 85
rect 3194 -51 3362 -23
rect 3194 -86 3253 -51
rect 3195 -97 3253 -86
rect 3299 -97 3362 -51
rect 3195 -149 3362 -97
rect 3985 -66 4153 -47
rect 3985 -112 4047 -66
rect 4093 -112 4153 -66
rect 3985 -121 4153 -112
rect 4257 -66 4425 -47
rect 6413 -48 6581 -20
rect 4257 -112 4335 -66
rect 4381 -112 4425 -66
rect 5045 -66 5213 -52
rect 5045 -102 5126 -66
rect 4257 -121 4425 -112
rect 5172 -102 5213 -66
rect 5861 -66 6029 -52
rect 5861 -102 5939 -66
rect 5126 -113 5172 -112
rect 5985 -102 6029 -66
rect 6413 -94 6472 -48
rect 6518 -94 6581 -48
rect 5939 -113 5985 -112
rect 6413 -146 6581 -94
rect 2159 -398 2216 -340
rect 2159 -444 2180 -398
rect 2226 -401 2259 -399
rect 2520 -404 2593 -340
rect 2159 -508 2216 -444
rect 2520 -450 2537 -404
rect 2583 -450 2593 -404
rect 2520 -508 2593 -450
rect 3195 -293 3362 -249
rect 3713 -281 3881 -253
rect 3713 -327 3772 -281
rect 3818 -327 3881 -281
rect 3713 -345 3881 -327
rect 4529 -279 4697 -251
rect 4529 -325 4588 -279
rect 4634 -325 4697 -279
rect 4529 -343 4697 -325
rect 5317 -290 5485 -287
rect 5317 -336 5379 -290
rect 5425 -336 5485 -290
rect 5317 -361 5485 -336
rect 5589 -290 5757 -287
rect 5589 -336 5656 -290
rect 5702 -336 5757 -290
rect 5589 -361 5757 -336
rect 3195 -463 3363 -435
rect 3195 -498 3254 -463
rect 3197 -509 3254 -498
rect 3300 -509 3363 -463
rect 3197 -561 3363 -509
rect 3985 -470 4153 -452
rect 3985 -516 4050 -470
rect 4096 -516 4153 -470
rect 3985 -526 4153 -516
rect 4257 -466 4425 -452
rect 4257 -512 4330 -466
rect 4376 -512 4425 -466
rect 5045 -470 5213 -456
rect 5045 -512 5115 -470
rect 4257 -526 4425 -512
rect 5161 -512 5213 -470
rect 5861 -471 6029 -456
rect 5861 -512 5928 -471
rect 5115 -517 5161 -516
rect 5974 -512 6029 -471
rect 6415 -458 6583 -430
rect 6415 -504 6474 -458
rect 6520 -504 6583 -458
rect 5928 -518 5974 -517
rect 6415 -556 6583 -504
rect 2138 -826 2231 -825
rect 2138 -889 2256 -826
rect 2138 -935 2166 -889
rect 2212 -935 2256 -889
rect 2138 -994 2256 -935
rect 2356 -994 2400 -826
rect 2502 -830 2595 -829
rect 3197 -703 3363 -661
rect 5317 -695 5485 -680
rect 3713 -741 3782 -699
rect 3828 -741 3881 -699
rect 3713 -757 3881 -741
rect 4529 -741 4599 -697
rect 4645 -741 4697 -697
rect 4529 -755 4697 -741
rect 5317 -741 5372 -695
rect 5418 -741 5485 -695
rect 5317 -754 5485 -741
rect 5589 -695 5757 -680
rect 5589 -741 5667 -695
rect 5713 -741 5757 -695
rect 6415 -700 6583 -656
rect 5589 -754 5757 -741
rect 2502 -893 2620 -830
rect 2502 -939 2530 -893
rect 2576 -939 2620 -893
rect 2502 -998 2620 -939
rect 2720 -998 2764 -830
<< polycontact >>
rect 2169 1196 2215 1242
rect 2530 1196 2576 1242
rect 2402 774 2448 820
rect 2752 767 2798 813
rect 3253 725 3299 771
rect 3769 708 3815 754
rect 4584 707 4630 753
rect 5392 707 5438 753
rect 5654 707 5700 753
rect 6472 728 6518 774
rect 2180 497 2226 543
rect 2540 500 2586 546
rect 4039 481 4085 527
rect 4316 481 4362 527
rect 5119 481 5165 527
rect 5939 481 5985 527
rect 3250 310 3296 356
rect 3786 298 3832 344
rect 4587 303 4633 349
rect 5372 303 5418 349
rect 5652 307 5698 353
rect 6472 318 6518 364
rect 2399 -37 2445 9
rect 2752 -48 2798 -2
rect 4044 85 4090 131
rect 4321 85 4367 131
rect 5098 84 5144 130
rect 5931 85 5977 131
rect 3253 -97 3299 -51
rect 4047 -112 4093 -66
rect 4335 -112 4381 -66
rect 5126 -112 5172 -66
rect 5939 -112 5985 -66
rect 6472 -94 6518 -48
rect 2180 -444 2226 -398
rect 2537 -450 2583 -404
rect 3772 -327 3818 -281
rect 4588 -325 4634 -279
rect 5379 -336 5425 -290
rect 5656 -336 5702 -290
rect 3254 -509 3300 -463
rect 4050 -516 4096 -470
rect 4330 -512 4376 -466
rect 5115 -516 5161 -470
rect 5928 -517 5974 -471
rect 6474 -504 6520 -458
rect 2166 -935 2212 -889
rect 3782 -741 3828 -695
rect 4599 -741 4645 -695
rect 5372 -741 5418 -695
rect 5667 -741 5713 -695
rect 2530 -939 2576 -893
<< metal1 >>
rect 1880 1547 2937 1566
rect 1880 1501 1902 1547
rect 1948 1501 2022 1547
rect 2068 1501 2142 1547
rect 2188 1501 2262 1547
rect 2308 1501 2382 1547
rect 2428 1501 2502 1547
rect 2548 1501 2622 1547
rect 2668 1501 2742 1547
rect 2788 1501 2937 1547
rect 1880 1485 2937 1501
rect 1880 1027 1962 1485
rect 2180 1382 2236 1485
rect 2527 1382 2589 1485
rect 2848 1465 2937 1485
rect 2848 1419 2869 1465
rect 2915 1419 2937 1465
rect 2140 1336 2356 1382
rect 2501 1380 2717 1382
rect 2140 1333 2357 1336
rect 2501 1333 2718 1380
rect 2140 1242 2235 1333
rect 2140 1196 2169 1242
rect 2215 1196 2235 1242
rect 2140 1108 2235 1196
rect 2501 1242 2596 1333
rect 2501 1196 2530 1242
rect 2576 1196 2596 1242
rect 2501 1108 2596 1196
rect 2848 1326 2937 1419
rect 2848 1280 2869 1326
rect 2915 1280 2937 1326
rect 2848 1163 2937 1280
rect 2848 1142 6839 1163
rect 2140 1061 2357 1108
rect 2501 1061 2718 1108
rect 2848 1096 2869 1142
rect 2915 1096 3038 1142
rect 3084 1096 3207 1142
rect 3253 1096 3407 1142
rect 3453 1096 3526 1142
rect 3572 1096 3645 1142
rect 3691 1096 3764 1142
rect 3810 1096 3883 1142
rect 3929 1096 4002 1142
rect 4048 1096 4121 1142
rect 4167 1096 4240 1142
rect 4286 1096 4359 1142
rect 4405 1096 4478 1142
rect 4524 1096 4597 1142
rect 4643 1096 4716 1142
rect 4762 1096 4835 1142
rect 4881 1096 4954 1142
rect 5000 1096 5073 1142
rect 5119 1096 5192 1142
rect 5238 1096 5311 1142
rect 5357 1096 5430 1142
rect 5476 1096 5549 1142
rect 5595 1096 5668 1142
rect 5714 1096 5787 1142
rect 5833 1096 5906 1142
rect 5952 1096 6025 1142
rect 6071 1096 6144 1142
rect 6190 1096 6263 1142
rect 6309 1141 6839 1142
rect 6309 1096 6403 1141
rect 2848 1095 6403 1096
rect 6449 1095 6561 1141
rect 6607 1095 6839 1141
rect 2848 1074 6839 1095
rect 1879 1006 1962 1027
rect 1879 960 1897 1006
rect 1943 960 1962 1006
rect 2943 996 3027 1074
rect 1879 883 1962 960
rect 2054 951 2134 952
rect 2265 951 2344 964
rect 2616 951 2719 966
rect 1879 837 1897 883
rect 1943 837 1962 883
rect 1879 769 1962 837
rect 1879 723 1897 769
rect 1943 723 1962 769
rect 1879 646 1962 723
rect 1879 600 1897 646
rect 1943 600 1962 646
rect 1879 529 1962 600
rect 1879 483 1897 529
rect 1943 483 1962 529
rect 1879 406 1962 483
rect 1879 360 1897 406
rect 1943 360 1962 406
rect 1879 289 1962 360
rect 1879 243 1897 289
rect 1943 243 1962 289
rect 1879 166 1962 243
rect 1879 120 1897 166
rect 1943 120 1962 166
rect 1879 49 1962 120
rect 1879 3 1897 49
rect 1943 3 1962 49
rect 1879 -74 1962 3
rect 1879 -120 1897 -74
rect 1943 -120 1962 -74
rect 1879 -191 1962 -120
rect 1879 -237 1897 -191
rect 1943 -237 1962 -191
rect 1879 -314 1962 -237
rect 1879 -360 1897 -314
rect 1943 -360 1962 -314
rect 1879 -431 1962 -360
rect 1879 -477 1897 -431
rect 1943 -477 1962 -431
rect 1879 -554 1962 -477
rect 1879 -600 1897 -554
rect 1943 -600 1962 -554
rect 1523 -657 1630 -623
rect 1436 -671 1630 -657
rect 1436 -723 1553 -671
rect 1605 -723 1630 -671
rect 1436 -737 1630 -723
rect 1523 -762 1630 -737
rect 1879 -681 1962 -600
rect 1879 -727 1897 -681
rect 1943 -727 1962 -681
rect 2008 899 2070 951
rect 2122 905 2357 951
rect 2122 899 2134 905
rect 2008 887 2134 899
rect 2008 272 2054 887
rect 2265 886 2344 905
rect 2616 899 2644 951
rect 2696 899 2719 951
rect 2616 887 2719 899
rect 2943 950 2961 996
rect 3007 950 3027 996
rect 2943 887 3027 950
rect 2943 841 2961 887
rect 3007 841 3027 887
rect 2374 823 2807 831
rect 2374 771 2398 823
rect 2450 816 2807 823
rect 2450 771 2742 816
rect 2794 813 2807 816
rect 2374 765 2742 771
rect 2798 767 2807 813
rect 2374 763 2460 765
rect 2730 764 2742 765
rect 2794 764 2807 767
rect 2730 752 2807 764
rect 2943 804 3027 841
rect 3910 890 3957 1074
rect 4454 890 4500 1074
rect 5242 890 5289 1074
rect 5786 890 5832 1074
rect 3910 844 5832 890
rect 2943 803 3156 804
rect 2943 778 3444 803
rect 2943 732 2961 778
rect 3007 771 3444 778
rect 3007 749 3253 771
rect 3007 732 3027 749
rect 2943 679 3027 732
rect 2261 647 3027 679
rect 2261 633 2961 647
rect 2943 601 2961 633
rect 3007 601 3027 647
rect 2164 546 2246 558
rect 2164 494 2178 546
rect 2230 494 2246 546
rect 2164 482 2246 494
rect 2529 548 2609 560
rect 2529 496 2536 548
rect 2588 496 2609 548
rect 2529 484 2609 496
rect 2943 517 3027 601
rect 3118 736 3253 749
rect 3118 574 3171 736
rect 3236 725 3253 736
rect 3299 736 3444 771
rect 3299 725 3316 736
rect 3236 709 3316 725
rect 3389 710 3444 736
rect 3758 755 3826 766
rect 3389 575 3443 710
rect 3758 703 3766 755
rect 3818 703 3826 755
rect 3758 677 3826 703
rect 3613 652 3691 669
rect 3613 649 3626 652
rect 3390 574 3443 575
rect 3537 600 3626 649
rect 3678 600 3691 652
rect 3537 586 3691 600
rect 3910 647 3957 844
rect 4167 651 4245 668
rect 2943 471 2961 517
rect 3007 471 3027 517
rect 2261 400 2357 407
rect 2261 361 2284 400
rect 2272 348 2284 361
rect 2336 348 2357 400
rect 2621 361 2717 407
rect 2943 388 3027 471
rect 2943 386 3439 388
rect 2272 336 2357 348
rect 2638 272 2684 361
rect 2008 226 2684 272
rect 2943 340 2961 386
rect 3007 356 3439 386
rect 3007 340 3250 356
rect 2943 333 3250 340
rect 2943 255 3027 333
rect 3113 321 3250 333
rect 3113 259 3167 321
rect 3233 310 3250 321
rect 3296 321 3439 356
rect 3296 310 3313 321
rect 3233 294 3313 310
rect 2008 -137 2054 226
rect 2943 209 2961 255
rect 3007 209 3027 255
rect 2943 135 3027 209
rect 3114 160 3167 259
rect 3386 160 3439 321
rect 2261 125 3027 135
rect 2261 89 2961 125
rect 2943 79 2961 89
rect 3007 79 3027 125
rect 2378 12 2456 24
rect 2378 -40 2396 12
rect 2448 6 2456 12
rect 2943 16 3027 79
rect 2734 6 2811 10
rect 2448 -2 2811 6
rect 2448 -40 2747 -2
rect 2378 -52 2456 -40
rect 2734 -54 2747 -40
rect 2799 -54 2811 -2
rect 2734 -66 2811 -54
rect 2943 -30 2961 16
rect 3007 -17 3027 16
rect 3007 -19 3161 -17
rect 3007 -30 3439 -19
rect 2943 -51 3439 -30
rect 2943 -72 3253 -51
rect 2943 -93 3027 -72
rect 2008 -183 2357 -137
rect 2008 -647 2054 -183
rect 2633 -189 2645 -137
rect 2697 -189 2709 -137
rect 2633 -201 2709 -189
rect 2943 -139 2961 -93
rect 3007 -139 3027 -93
rect 2943 -245 3027 -139
rect 2943 -265 2961 -245
rect 2261 -291 2961 -265
rect 3007 -291 3027 -245
rect 3116 -86 3253 -72
rect 3116 -248 3169 -86
rect 3236 -97 3253 -86
rect 3299 -86 3439 -51
rect 3299 -97 3316 -86
rect 3236 -113 3316 -97
rect 3389 -111 3439 -86
rect 3389 -248 3442 -111
rect 2261 -311 3027 -291
rect 2173 -387 2255 -383
rect 2169 -395 2255 -387
rect 2169 -398 2191 -395
rect 2169 -444 2180 -398
rect 2169 -447 2191 -444
rect 2243 -447 2255 -395
rect 2169 -455 2255 -447
rect 2173 -459 2255 -455
rect 2505 -401 2593 -389
rect 2505 -453 2535 -401
rect 2587 -453 2593 -401
rect 2505 -466 2593 -453
rect 2943 -398 3027 -311
rect 2943 -444 2961 -398
rect 3007 -431 3027 -398
rect 3007 -444 3440 -431
rect 2943 -463 3440 -444
rect 2943 -486 3254 -463
rect 2270 -589 2282 -537
rect 2334 -589 2346 -537
rect 2621 -583 2717 -537
rect 2943 -572 3027 -486
rect 2270 -601 2346 -589
rect 2648 -647 2694 -583
rect 2008 -693 2694 -647
rect 2943 -618 2961 -572
rect 3007 -618 3027 -572
rect 1879 -1157 1962 -727
rect 2943 -702 3027 -618
rect 3119 -498 3254 -486
rect 3119 -659 3172 -498
rect 3237 -509 3254 -498
rect 3300 -498 3440 -463
rect 3300 -509 3317 -498
rect 3237 -525 3317 -509
rect 3390 -522 3440 -498
rect 3390 -659 3443 -522
rect 3537 -568 3583 586
rect 3910 409 3956 647
rect 4167 599 4180 651
rect 4232 599 4245 651
rect 4167 585 4245 599
rect 4028 530 4096 555
rect 4028 478 4036 530
rect 4088 478 4096 530
rect 4028 469 4096 478
rect 4305 530 4373 555
rect 4305 478 4313 530
rect 4365 478 4373 530
rect 4305 469 4373 478
rect 4454 465 4500 844
rect 4573 753 4641 764
rect 4573 701 4581 753
rect 4633 701 4641 753
rect 4573 675 4641 701
rect 5242 672 5289 844
rect 5381 753 5449 764
rect 5381 701 5389 753
rect 5441 701 5449 753
rect 5381 675 5449 701
rect 5643 753 5711 764
rect 5643 701 5651 753
rect 5703 701 5711 753
rect 5643 675 5711 701
rect 4712 652 4790 669
rect 4712 600 4725 652
rect 4777 600 4790 652
rect 4712 586 4790 600
rect 4957 651 5035 668
rect 4957 599 4970 651
rect 5022 599 5035 651
rect 4957 585 5035 599
rect 5108 530 5176 555
rect 5108 478 5116 530
rect 5168 478 5176 530
rect 5108 469 5176 478
rect 5242 475 5288 672
rect 5496 644 5574 661
rect 5496 592 5509 644
rect 5561 592 5574 644
rect 5496 578 5574 592
rect 5786 475 5832 844
rect 6756 1034 6839 1074
rect 6756 988 6774 1034
rect 6820 988 6839 1034
rect 6756 915 6839 988
rect 6756 869 6774 915
rect 6820 869 6839 915
rect 6337 800 6658 807
rect 6756 800 6839 869
rect 6337 796 6839 800
rect 6337 774 6774 796
rect 6337 739 6472 774
rect 6043 651 6121 668
rect 6043 599 6056 651
rect 6108 648 6121 651
rect 6108 599 6240 648
rect 6043 598 6240 599
rect 6043 585 6121 598
rect 4454 419 4983 465
rect 4454 409 4500 419
rect 3910 363 4500 409
rect 3775 345 3843 356
rect 3775 293 3783 345
rect 3835 293 3843 345
rect 3775 267 3843 293
rect 3638 258 3684 262
rect 3629 241 3707 258
rect 3629 189 3642 241
rect 3694 189 3707 241
rect 3629 175 3707 189
rect 3638 -157 3684 175
rect 3630 -174 3708 -157
rect 3630 -226 3643 -174
rect 3695 -226 3708 -174
rect 3630 -240 3708 -226
rect 3638 -244 3684 -240
rect 3761 -278 3829 -253
rect 3761 -330 3769 -278
rect 3821 -330 3829 -278
rect 3761 -339 3829 -330
rect 3910 -361 3956 363
rect 4165 239 4243 256
rect 4165 187 4178 239
rect 4230 187 4243 239
rect 4165 173 4243 187
rect 4033 134 4101 159
rect 4033 82 4041 134
rect 4093 82 4101 134
rect 4033 73 4101 82
rect 4310 134 4378 159
rect 4310 82 4318 134
rect 4370 82 4378 134
rect 4310 73 4378 82
rect 4036 -65 4104 -54
rect 4036 -117 4044 -65
rect 4096 -117 4104 -65
rect 4036 -143 4104 -117
rect 4324 -65 4392 -54
rect 4324 -117 4332 -65
rect 4384 -117 4392 -65
rect 4324 -143 4392 -117
rect 4164 -193 4242 -176
rect 4164 -245 4177 -193
rect 4229 -245 4242 -193
rect 4164 -259 4242 -245
rect 4454 -361 4500 363
rect 4937 402 4983 419
rect 5242 429 5832 475
rect 5928 530 5996 555
rect 5928 478 5936 530
rect 5988 478 5996 530
rect 5928 469 5996 478
rect 5242 402 5288 429
rect 4576 350 4644 361
rect 4937 356 5288 402
rect 4576 298 4584 350
rect 4636 298 4644 350
rect 4576 272 4644 298
rect 4708 239 4786 256
rect 4708 187 4721 239
rect 4773 187 4786 239
rect 4708 173 4786 187
rect 4942 237 5020 254
rect 4942 185 4955 237
rect 5007 185 5020 237
rect 4942 184 5020 185
rect 4942 171 4970 184
rect 5016 171 5020 184
rect 5087 133 5155 158
rect 5087 81 5095 133
rect 5147 81 5155 133
rect 5087 72 5155 81
rect 5115 -65 5183 -54
rect 4708 -133 4786 -116
rect 5115 -117 5123 -65
rect 5175 -117 5183 -65
rect 4708 -185 4721 -133
rect 4773 -185 4786 -133
rect 4708 -199 4786 -185
rect 4951 -142 5029 -125
rect 4951 -194 4964 -142
rect 5016 -194 5029 -142
rect 5115 -143 5183 -117
rect 4951 -208 5029 -194
rect 4577 -276 4645 -251
rect 4577 -328 4585 -276
rect 4637 -328 4645 -276
rect 4577 -337 4645 -328
rect 3910 -407 4500 -361
rect 5242 -363 5288 356
rect 5361 350 5429 361
rect 5361 298 5369 350
rect 5421 298 5429 350
rect 5361 272 5429 298
rect 5641 354 5709 365
rect 5641 302 5649 354
rect 5701 302 5709 354
rect 5641 276 5709 302
rect 5496 222 5574 239
rect 5496 170 5509 222
rect 5561 170 5574 222
rect 5496 156 5574 170
rect 5495 -176 5573 -159
rect 5495 -228 5508 -176
rect 5560 -228 5573 -176
rect 5495 -242 5573 -228
rect 5368 -287 5436 -262
rect 5368 -339 5376 -287
rect 5428 -339 5436 -287
rect 5368 -348 5436 -339
rect 5645 -287 5713 -262
rect 5645 -339 5653 -287
rect 5705 -339 5713 -287
rect 5645 -348 5713 -339
rect 3638 -568 3684 -558
rect 3537 -585 3699 -568
rect 3537 -631 3634 -585
rect 3621 -637 3634 -631
rect 3686 -637 3699 -585
rect 3621 -651 3699 -637
rect 3638 -654 3684 -651
rect 2943 -748 2961 -702
rect 3007 -748 3027 -702
rect 2137 -751 2353 -749
rect 2137 -797 2283 -751
rect 2329 -797 2354 -751
rect 2137 -798 2354 -797
rect 2501 -755 2717 -753
rect 2137 -889 2232 -798
rect 2137 -935 2166 -889
rect 2212 -935 2232 -889
rect 2137 -1023 2232 -935
rect 2501 -801 2647 -755
rect 2693 -801 2718 -755
rect 2501 -802 2718 -801
rect 2501 -893 2596 -802
rect 2943 -811 3027 -748
rect 3771 -692 3839 -667
rect 3771 -744 3779 -692
rect 3831 -744 3839 -692
rect 3771 -753 3839 -744
rect 2943 -857 2961 -811
rect 3007 -857 3027 -811
rect 2943 -882 3027 -857
rect 2501 -939 2530 -893
rect 2576 -939 2596 -893
rect 2137 -1069 2283 -1023
rect 2329 -1069 2354 -1023
rect 2137 -1070 2354 -1069
rect 2501 -1027 2596 -939
rect 2823 -901 3027 -882
rect 2823 -903 3078 -901
rect 3910 -903 3956 -407
rect 4454 -424 4500 -407
rect 4934 -409 5288 -363
rect 4934 -424 4980 -409
rect 4039 -469 4107 -458
rect 4039 -521 4047 -469
rect 4099 -521 4107 -469
rect 4039 -547 4107 -521
rect 4319 -465 4387 -454
rect 4319 -517 4327 -465
rect 4379 -517 4387 -465
rect 4319 -543 4387 -517
rect 4454 -470 4980 -424
rect 5242 -421 5288 -409
rect 5786 -421 5832 429
rect 6058 256 6104 262
rect 6042 239 6120 256
rect 6042 187 6055 239
rect 6107 187 6120 239
rect 6042 186 6120 187
rect 6042 173 6058 186
rect 6104 173 6120 186
rect 5920 134 5988 159
rect 5920 82 5928 134
rect 5980 82 5988 134
rect 5920 73 5988 82
rect 5928 -65 5996 -54
rect 5928 -117 5936 -65
rect 5988 -117 5996 -65
rect 5928 -143 5996 -117
rect 6035 -194 6058 -178
rect 6104 -194 6113 -178
rect 6035 -195 6113 -194
rect 6035 -247 6048 -195
rect 6100 -247 6113 -195
rect 6035 -261 6113 -247
rect 5104 -469 5172 -458
rect 4163 -598 4241 -581
rect 4163 -650 4176 -598
rect 4228 -650 4241 -598
rect 4163 -664 4241 -650
rect 4454 -903 4500 -470
rect 5104 -521 5112 -469
rect 5164 -521 5172 -469
rect 5104 -547 5172 -521
rect 5242 -467 5832 -421
rect 4720 -587 4798 -570
rect 4720 -639 4733 -587
rect 4785 -639 4798 -587
rect 4720 -653 4798 -639
rect 4956 -590 5034 -573
rect 4956 -642 4969 -590
rect 5021 -642 5034 -590
rect 4956 -656 5034 -642
rect 4588 -692 4656 -667
rect 4588 -744 4596 -692
rect 4648 -744 4656 -692
rect 4588 -753 4656 -744
rect 5242 -903 5288 -467
rect 5485 -591 5563 -574
rect 5485 -643 5498 -591
rect 5550 -643 5563 -591
rect 5485 -657 5563 -643
rect 5361 -692 5429 -667
rect 5361 -744 5369 -692
rect 5421 -744 5429 -692
rect 5361 -753 5429 -744
rect 5656 -692 5724 -667
rect 5656 -744 5664 -692
rect 5716 -744 5724 -692
rect 5656 -753 5724 -744
rect 5786 -903 5832 -467
rect 5917 -470 5985 -459
rect 5917 -522 5925 -470
rect 5977 -522 5985 -470
rect 5917 -548 5985 -522
rect 6058 -583 6104 -558
rect 6190 -583 6240 598
rect 6337 579 6385 739
rect 6455 728 6472 739
rect 6518 750 6774 774
rect 6820 750 6839 796
rect 6518 739 6658 750
rect 6518 728 6535 739
rect 6455 712 6535 728
rect 6608 578 6658 739
rect 6756 677 6839 750
rect 6756 631 6774 677
rect 6820 631 6839 677
rect 6756 558 6839 631
rect 6756 512 6774 558
rect 6820 512 6839 558
rect 6756 439 6839 512
rect 6337 390 6658 397
rect 6756 393 6774 439
rect 6820 393 6839 439
rect 6756 390 6839 393
rect 6337 364 6839 390
rect 6337 329 6472 364
rect 6337 239 6385 329
rect 6455 318 6472 329
rect 6518 340 6839 364
rect 6518 329 6658 340
rect 6518 318 6535 329
rect 6455 302 6535 318
rect 6337 193 6338 239
rect 6384 193 6385 239
rect 6337 169 6385 193
rect 6608 239 6658 329
rect 6608 193 6610 239
rect 6656 193 6658 239
rect 6338 168 6384 169
rect 6608 168 6658 193
rect 6756 320 6839 340
rect 6756 274 6774 320
rect 6820 274 6839 320
rect 6756 201 6839 274
rect 6756 155 6774 201
rect 6820 155 6839 201
rect 6756 82 6839 155
rect 6756 36 6774 82
rect 6820 36 6839 82
rect 6337 -29 6658 -15
rect 6756 -29 6839 36
rect 6337 -37 6839 -29
rect 6337 -48 6774 -37
rect 6337 -83 6472 -48
rect 6337 -173 6385 -83
rect 6455 -94 6472 -83
rect 6518 -79 6774 -48
rect 6518 -83 6658 -79
rect 6518 -94 6535 -83
rect 6455 -110 6535 -94
rect 6337 -219 6338 -173
rect 6384 -219 6385 -173
rect 6337 -243 6385 -219
rect 6608 -173 6658 -83
rect 6608 -219 6610 -173
rect 6656 -219 6658 -173
rect 6608 -243 6658 -219
rect 6756 -83 6774 -79
rect 6820 -83 6839 -37
rect 6756 -156 6839 -83
rect 6756 -202 6774 -156
rect 6820 -202 6839 -156
rect 6756 -275 6839 -202
rect 6756 -321 6774 -275
rect 6820 -321 6839 -275
rect 6756 -394 6839 -321
rect 6058 -611 6240 -583
rect 6035 -628 6240 -611
rect 6035 -680 6048 -628
rect 6100 -633 6240 -628
rect 6339 -433 6660 -425
rect 6756 -433 6774 -394
rect 6339 -440 6774 -433
rect 6820 -440 6839 -394
rect 6339 -458 6839 -440
rect 6339 -493 6474 -458
rect 6339 -583 6387 -493
rect 6457 -504 6474 -493
rect 6520 -483 6839 -458
rect 6520 -493 6660 -483
rect 6520 -504 6537 -493
rect 6457 -520 6537 -504
rect 6339 -629 6340 -583
rect 6386 -629 6387 -583
rect 6100 -680 6113 -633
rect 6339 -653 6387 -629
rect 6610 -583 6660 -493
rect 6610 -629 6612 -583
rect 6658 -629 6660 -583
rect 6340 -654 6386 -653
rect 6610 -654 6660 -629
rect 6756 -513 6839 -483
rect 6756 -559 6774 -513
rect 6820 -559 6839 -513
rect 6756 -632 6839 -559
rect 6035 -694 6113 -680
rect 6756 -678 6774 -632
rect 6820 -678 6839 -632
rect 6756 -751 6839 -678
rect 6756 -797 6774 -751
rect 6820 -797 6839 -751
rect 6756 -903 6839 -797
rect 2823 -924 6856 -903
rect 2823 -927 3416 -924
rect 2823 -973 3112 -927
rect 3158 -973 3282 -927
rect 3328 -970 3416 -927
rect 3462 -970 3535 -924
rect 3581 -970 3654 -924
rect 3700 -970 3773 -924
rect 3819 -970 3892 -924
rect 3938 -970 4011 -924
rect 4057 -970 4130 -924
rect 4176 -970 4249 -924
rect 4295 -970 4368 -924
rect 4414 -970 4487 -924
rect 4533 -970 4606 -924
rect 4652 -970 4725 -924
rect 4771 -970 4844 -924
rect 4890 -970 4963 -924
rect 5009 -970 5082 -924
rect 5128 -970 5201 -924
rect 5247 -970 5320 -924
rect 5366 -970 5439 -924
rect 5485 -970 5558 -924
rect 5604 -970 5677 -924
rect 5723 -970 5796 -924
rect 5842 -970 5915 -924
rect 5961 -970 6034 -924
rect 6080 -970 6153 -924
rect 6199 -970 6272 -924
rect 6318 -970 6423 -924
rect 6469 -970 6567 -924
rect 6613 -970 6791 -924
rect 6837 -970 6856 -924
rect 3328 -973 6856 -970
rect 2823 -992 6856 -973
rect 2137 -1157 2195 -1070
rect 2501 -1073 2647 -1027
rect 2693 -1073 2718 -1027
rect 2501 -1074 2718 -1073
rect 2501 -1157 2570 -1074
rect 2656 -1157 2703 -1074
rect 2823 -1157 2895 -992
rect 1877 -1178 2895 -1157
rect 1877 -1224 1902 -1178
rect 1948 -1224 2022 -1178
rect 2068 -1224 2142 -1178
rect 2188 -1224 2262 -1178
rect 2308 -1224 2382 -1178
rect 2428 -1224 2502 -1178
rect 2548 -1224 2622 -1178
rect 2668 -1224 2742 -1178
rect 2788 -1224 2895 -1178
rect 1877 -1245 2895 -1224
<< via1 >>
rect 1553 -723 1605 -671
rect 2070 899 2122 951
rect 2644 899 2696 951
rect 2398 820 2450 823
rect 2398 774 2402 820
rect 2402 774 2448 820
rect 2448 774 2450 820
rect 2398 771 2450 774
rect 2742 813 2794 816
rect 2742 767 2752 813
rect 2752 767 2794 813
rect 2742 764 2794 767
rect 2178 543 2230 546
rect 2178 497 2180 543
rect 2180 497 2226 543
rect 2226 497 2230 543
rect 2178 494 2230 497
rect 2536 546 2588 548
rect 2536 500 2540 546
rect 2540 500 2586 546
rect 2586 500 2588 546
rect 2536 496 2588 500
rect 3766 754 3818 755
rect 3766 708 3769 754
rect 3769 708 3815 754
rect 3815 708 3818 754
rect 3766 703 3818 708
rect 3626 600 3678 652
rect 2284 348 2336 400
rect 2396 9 2448 12
rect 2396 -37 2399 9
rect 2399 -37 2445 9
rect 2445 -37 2448 9
rect 2396 -40 2448 -37
rect 2747 -48 2752 -2
rect 2752 -48 2798 -2
rect 2798 -48 2799 -2
rect 2747 -54 2799 -48
rect 2645 -189 2697 -137
rect 2191 -398 2243 -395
rect 2191 -444 2226 -398
rect 2226 -444 2243 -398
rect 2191 -447 2243 -444
rect 2535 -404 2587 -401
rect 2535 -450 2537 -404
rect 2537 -450 2583 -404
rect 2583 -450 2587 -404
rect 2535 -453 2587 -450
rect 2282 -589 2334 -537
rect 4180 599 4232 651
rect 4036 527 4088 530
rect 4036 481 4039 527
rect 4039 481 4085 527
rect 4085 481 4088 527
rect 4036 478 4088 481
rect 4313 527 4365 530
rect 4313 481 4316 527
rect 4316 481 4362 527
rect 4362 481 4365 527
rect 4313 478 4365 481
rect 4581 707 4584 753
rect 4584 707 4630 753
rect 4630 707 4633 753
rect 4581 701 4633 707
rect 5389 707 5392 753
rect 5392 707 5438 753
rect 5438 707 5441 753
rect 5389 701 5441 707
rect 5651 707 5654 753
rect 5654 707 5700 753
rect 5700 707 5703 753
rect 5651 701 5703 707
rect 4725 600 4777 652
rect 4970 599 5022 651
rect 5116 527 5168 530
rect 5116 481 5119 527
rect 5119 481 5165 527
rect 5165 481 5168 527
rect 5116 478 5168 481
rect 5509 592 5561 644
rect 6056 599 6108 651
rect 3783 344 3835 345
rect 3783 298 3786 344
rect 3786 298 3832 344
rect 3832 298 3835 344
rect 3783 293 3835 298
rect 3642 189 3694 241
rect 3643 -226 3695 -174
rect 3769 -281 3821 -278
rect 3769 -327 3772 -281
rect 3772 -327 3818 -281
rect 3818 -327 3821 -281
rect 3769 -330 3821 -327
rect 4178 187 4230 239
rect 4041 131 4093 134
rect 4041 85 4044 131
rect 4044 85 4090 131
rect 4090 85 4093 131
rect 4041 82 4093 85
rect 4318 131 4370 134
rect 4318 85 4321 131
rect 4321 85 4367 131
rect 4367 85 4370 131
rect 4318 82 4370 85
rect 4044 -66 4096 -65
rect 4044 -112 4047 -66
rect 4047 -112 4093 -66
rect 4093 -112 4096 -66
rect 4044 -117 4096 -112
rect 4332 -66 4384 -65
rect 4332 -112 4335 -66
rect 4335 -112 4381 -66
rect 4381 -112 4384 -66
rect 4332 -117 4384 -112
rect 4177 -245 4229 -193
rect 5936 527 5988 530
rect 5936 481 5939 527
rect 5939 481 5985 527
rect 5985 481 5988 527
rect 5936 478 5988 481
rect 4584 349 4636 350
rect 4584 303 4587 349
rect 4587 303 4633 349
rect 4633 303 4636 349
rect 4584 298 4636 303
rect 4721 187 4773 239
rect 4955 185 5007 237
rect 5095 130 5147 133
rect 5095 84 5098 130
rect 5098 84 5144 130
rect 5144 84 5147 130
rect 5095 81 5147 84
rect 5123 -66 5175 -65
rect 5123 -112 5126 -66
rect 5126 -112 5172 -66
rect 5172 -112 5175 -66
rect 5123 -117 5175 -112
rect 4721 -185 4773 -133
rect 4964 -194 5016 -142
rect 4585 -279 4637 -276
rect 4585 -325 4588 -279
rect 4588 -325 4634 -279
rect 4634 -325 4637 -279
rect 4585 -328 4637 -325
rect 5369 349 5421 350
rect 5369 303 5372 349
rect 5372 303 5418 349
rect 5418 303 5421 349
rect 5369 298 5421 303
rect 5649 353 5701 354
rect 5649 307 5652 353
rect 5652 307 5698 353
rect 5698 307 5701 353
rect 5649 302 5701 307
rect 5509 170 5561 222
rect 5508 -228 5560 -176
rect 5376 -290 5428 -287
rect 5376 -336 5379 -290
rect 5379 -336 5425 -290
rect 5425 -336 5428 -290
rect 5376 -339 5428 -336
rect 5653 -290 5705 -287
rect 5653 -336 5656 -290
rect 5656 -336 5702 -290
rect 5702 -336 5705 -290
rect 5653 -339 5705 -336
rect 3634 -637 3686 -585
rect 3779 -695 3831 -692
rect 3779 -741 3782 -695
rect 3782 -741 3828 -695
rect 3828 -741 3831 -695
rect 3779 -744 3831 -741
rect 4047 -470 4099 -469
rect 4047 -516 4050 -470
rect 4050 -516 4096 -470
rect 4096 -516 4099 -470
rect 4047 -521 4099 -516
rect 4327 -466 4379 -465
rect 4327 -512 4330 -466
rect 4330 -512 4376 -466
rect 4376 -512 4379 -466
rect 4327 -517 4379 -512
rect 6055 187 6107 239
rect 5928 131 5980 134
rect 5928 85 5931 131
rect 5931 85 5977 131
rect 5977 85 5980 131
rect 5928 82 5980 85
rect 5936 -66 5988 -65
rect 5936 -112 5939 -66
rect 5939 -112 5985 -66
rect 5985 -112 5988 -66
rect 5936 -117 5988 -112
rect 6048 -247 6100 -195
rect 4176 -650 4228 -598
rect 5112 -470 5164 -469
rect 5112 -516 5115 -470
rect 5115 -516 5161 -470
rect 5161 -516 5164 -470
rect 5112 -521 5164 -516
rect 4733 -639 4785 -587
rect 4969 -642 5021 -590
rect 4596 -695 4648 -692
rect 4596 -741 4599 -695
rect 4599 -741 4645 -695
rect 4645 -741 4648 -695
rect 4596 -744 4648 -741
rect 5498 -643 5550 -591
rect 5369 -695 5421 -692
rect 5369 -741 5372 -695
rect 5372 -741 5418 -695
rect 5418 -741 5421 -695
rect 5369 -744 5421 -741
rect 5664 -695 5716 -692
rect 5664 -741 5667 -695
rect 5667 -741 5713 -695
rect 5713 -741 5716 -695
rect 5664 -744 5716 -741
rect 5925 -471 5977 -470
rect 5925 -517 5928 -471
rect 5928 -517 5974 -471
rect 5974 -517 5977 -471
rect 5925 -522 5977 -517
rect 6048 -680 6100 -628
<< metal2 >>
rect 2054 953 2137 966
rect 2054 897 2068 953
rect 2124 897 2137 953
rect 2054 885 2137 897
rect 2444 831 2524 1329
rect 2374 823 2524 831
rect 2374 771 2398 823
rect 2450 771 2524 823
rect 2374 763 2524 771
rect 2444 560 2524 763
rect 2622 963 2684 965
rect 2622 951 2698 963
rect 2622 899 2644 951
rect 2696 899 2698 951
rect 2622 876 2698 899
rect 2622 688 2684 876
rect 2740 816 2912 828
rect 3689 820 6250 893
rect 2740 764 2742 816
rect 2794 764 2912 816
rect 2740 752 2912 764
rect 2622 626 2776 688
rect 2093 546 2238 558
rect 2093 494 2178 546
rect 2230 494 2238 546
rect 2093 482 2238 494
rect 2444 548 2599 560
rect 2444 496 2536 548
rect 2588 496 2599 548
rect 2444 484 2599 496
rect 2093 -383 2173 482
rect 2233 400 2339 412
rect 2233 390 2284 400
rect 2231 348 2284 390
rect 2336 348 2339 400
rect 2231 336 2339 348
rect 2231 -212 2287 336
rect 2444 80 2524 484
rect 2714 156 2776 626
rect 2602 94 2776 156
rect 2444 24 2525 80
rect 2378 12 2525 24
rect 2378 -40 2396 12
rect 2448 -40 2525 12
rect 2378 -52 2525 -40
rect 2231 -268 2382 -212
rect 2093 -395 2255 -383
rect 2093 -447 2191 -395
rect 2243 -447 2255 -395
rect 2093 -459 2255 -447
rect 1523 -657 1630 -623
rect 2093 -657 2173 -459
rect 2326 -522 2382 -268
rect 2444 -389 2525 -52
rect 2602 -125 2664 94
rect 2832 10 2912 752
rect 3758 755 3826 820
rect 3758 703 3766 755
rect 3818 703 3826 755
rect 3758 694 3826 703
rect 4573 753 4641 820
rect 4573 701 4581 753
rect 4633 701 4641 753
rect 4573 692 4641 701
rect 5381 753 5449 820
rect 5381 701 5389 753
rect 5441 701 5449 753
rect 5381 692 5449 701
rect 5643 753 5711 820
rect 5643 701 5651 753
rect 5703 701 5711 753
rect 5643 692 5711 701
rect 3613 654 3691 669
rect 3613 652 3624 654
rect 3612 598 3624 652
rect 3680 598 3691 654
rect 3612 586 3691 598
rect 4167 653 4245 668
rect 4712 660 4790 669
rect 4167 597 4178 653
rect 4234 597 4245 653
rect 3612 445 3685 586
rect 4167 585 4245 597
rect 4711 654 4790 660
rect 4711 598 4723 654
rect 4779 598 4790 654
rect 4711 586 4790 598
rect 4957 653 5035 668
rect 4957 597 4968 653
rect 5024 597 5035 653
rect 4028 530 4096 540
rect 4028 478 4036 530
rect 4088 478 4096 530
rect 4028 445 4096 478
rect 4305 530 4373 540
rect 4305 478 4313 530
rect 4365 478 4373 530
rect 4305 445 4373 478
rect 4711 445 4784 586
rect 4957 585 5035 597
rect 5496 646 5574 661
rect 5496 590 5507 646
rect 5563 590 5574 646
rect 5496 578 5574 590
rect 6043 653 6121 668
rect 6043 597 6054 653
rect 6110 597 6121 653
rect 6043 585 6121 597
rect 5108 530 5176 540
rect 5108 478 5116 530
rect 5168 478 5176 530
rect 5108 445 5176 478
rect 5928 530 5996 540
rect 5928 478 5936 530
rect 5988 478 5996 530
rect 5928 445 5996 478
rect 2734 -2 2912 10
rect 2734 -54 2747 -2
rect 2799 -54 2912 -2
rect 2734 -66 2912 -54
rect 2602 -134 2752 -125
rect 2602 -190 2641 -134
rect 2697 -190 2752 -134
rect 2602 -201 2752 -190
rect 2444 -401 2593 -389
rect 2444 -453 2535 -401
rect 2587 -453 2593 -401
rect 2444 -465 2593 -453
rect 2444 -466 2525 -465
rect 2680 -522 2752 -201
rect 2326 -525 2752 -522
rect 2280 -537 2752 -525
rect 2280 -589 2282 -537
rect 2334 -589 2752 -537
rect 2280 -601 2752 -589
rect 2832 -657 2912 -66
rect 3500 372 6041 445
rect 3500 -356 3573 372
rect 3775 345 3843 372
rect 3775 293 3783 345
rect 3835 293 3843 345
rect 3775 284 3843 293
rect 4576 350 4644 372
rect 4576 298 4584 350
rect 4636 298 4644 350
rect 4576 289 4644 298
rect 5361 350 5429 372
rect 5361 298 5369 350
rect 5421 298 5429 350
rect 5361 289 5429 298
rect 5641 354 5709 372
rect 5641 302 5649 354
rect 5701 302 5709 354
rect 5641 293 5709 302
rect 3629 243 3707 258
rect 3629 187 3640 243
rect 3696 187 3707 243
rect 3629 175 3707 187
rect 4165 241 4243 256
rect 4165 185 4176 241
rect 4232 185 4243 241
rect 4165 173 4243 185
rect 4708 241 4786 256
rect 4708 185 4719 241
rect 4775 185 4786 241
rect 4708 173 4786 185
rect 4942 239 5020 254
rect 6042 241 6120 256
rect 4942 183 4953 239
rect 5009 183 5020 239
rect 4942 171 5020 183
rect 5496 224 5574 239
rect 5496 168 5507 224
rect 5563 168 5574 224
rect 6042 185 6053 241
rect 6109 185 6120 241
rect 6042 173 6120 185
rect 5496 156 5574 168
rect 4033 134 4101 144
rect 4033 82 4041 134
rect 4093 82 4101 134
rect 4033 49 4101 82
rect 4310 134 4378 144
rect 4310 82 4318 134
rect 4370 82 4378 134
rect 4310 49 4378 82
rect 5087 133 5155 143
rect 5087 81 5095 133
rect 5147 81 5155 133
rect 5087 49 5155 81
rect 5920 134 5988 144
rect 5920 82 5928 134
rect 5980 82 5988 134
rect 5920 49 5988 82
rect 6177 49 6250 820
rect 3634 -24 6250 49
rect 3634 -157 3707 -24
rect 4036 -65 4104 -24
rect 4036 -117 4044 -65
rect 4096 -117 4104 -65
rect 4036 -126 4104 -117
rect 4324 -65 4392 -24
rect 4324 -117 4332 -65
rect 4384 -117 4392 -65
rect 5115 -65 5183 -24
rect 4324 -126 4392 -117
rect 4708 -131 4786 -116
rect 5115 -117 5123 -65
rect 5175 -117 5183 -65
rect 3630 -172 3708 -157
rect 3630 -228 3641 -172
rect 3697 -228 3708 -172
rect 3630 -240 3708 -228
rect 4164 -191 4242 -176
rect 3634 -242 3707 -240
rect 4164 -247 4175 -191
rect 4231 -247 4242 -191
rect 4708 -187 4719 -131
rect 4775 -187 4786 -131
rect 4708 -199 4786 -187
rect 4951 -140 5029 -125
rect 5115 -126 5183 -117
rect 5928 -65 5996 -24
rect 5928 -117 5936 -65
rect 5988 -117 5996 -65
rect 5928 -126 5996 -117
rect 4951 -196 4962 -140
rect 5018 -196 5029 -140
rect 4951 -208 5029 -196
rect 5495 -174 5573 -159
rect 5495 -230 5506 -174
rect 5562 -230 5573 -174
rect 5495 -242 5573 -230
rect 6035 -193 6113 -178
rect 4164 -259 4242 -247
rect 6035 -249 6046 -193
rect 6102 -249 6113 -193
rect 6035 -261 6113 -249
rect 3761 -278 3829 -268
rect 3761 -330 3769 -278
rect 3821 -330 3829 -278
rect 3761 -356 3829 -330
rect 4577 -276 4645 -266
rect 4577 -328 4585 -276
rect 4637 -328 4645 -276
rect 4577 -356 4645 -328
rect 5368 -287 5436 -277
rect 5368 -339 5376 -287
rect 5428 -339 5436 -287
rect 5368 -356 5436 -339
rect 5645 -287 5713 -277
rect 5645 -339 5653 -287
rect 5705 -339 5713 -287
rect 5645 -356 5713 -339
rect 3500 -429 6046 -356
rect 3625 -568 3698 -429
rect 4039 -469 4107 -429
rect 4039 -521 4047 -469
rect 4099 -521 4107 -469
rect 4039 -530 4107 -521
rect 4319 -465 4387 -429
rect 4319 -517 4327 -465
rect 4379 -517 4387 -465
rect 4319 -526 4387 -517
rect 5104 -469 5172 -429
rect 5104 -521 5112 -469
rect 5164 -521 5172 -469
rect 5104 -530 5172 -521
rect 5917 -470 5985 -429
rect 5917 -522 5925 -470
rect 5977 -522 5985 -470
rect 5917 -531 5985 -522
rect 3621 -583 3699 -568
rect 3621 -639 3632 -583
rect 3688 -639 3699 -583
rect 3621 -651 3699 -639
rect 4163 -596 4241 -581
rect 1523 -671 2912 -657
rect 4163 -652 4174 -596
rect 4230 -652 4241 -596
rect 4163 -664 4241 -652
rect 4720 -585 4798 -570
rect 4720 -641 4731 -585
rect 4787 -641 4798 -585
rect 4720 -653 4798 -641
rect 4956 -588 5034 -573
rect 4956 -644 4967 -588
rect 5023 -644 5034 -588
rect 4956 -656 5034 -644
rect 5485 -589 5563 -574
rect 5485 -645 5496 -589
rect 5552 -645 5563 -589
rect 5485 -657 5563 -645
rect 6035 -626 6113 -611
rect 1523 -723 1553 -671
rect 1605 -723 2912 -671
rect 6035 -682 6046 -626
rect 6102 -682 6113 -626
rect 1523 -737 2912 -723
rect 3771 -692 3839 -682
rect 1523 -762 1630 -737
rect 2093 -895 2173 -737
rect 3771 -744 3779 -692
rect 3831 -744 3839 -692
rect 3771 -777 3839 -744
rect 4588 -692 4656 -682
rect 4588 -744 4596 -692
rect 4648 -744 4656 -692
rect 4588 -777 4656 -744
rect 5361 -692 5429 -682
rect 5361 -744 5369 -692
rect 5421 -744 5429 -692
rect 5361 -777 5429 -744
rect 5656 -692 5724 -682
rect 5656 -744 5664 -692
rect 5716 -744 5724 -692
rect 6035 -694 6113 -682
rect 5656 -777 5724 -744
rect 6177 -777 6250 -24
rect 3689 -850 6250 -777
<< via2 >>
rect 2068 951 2124 953
rect 2068 899 2070 951
rect 2070 899 2122 951
rect 2122 899 2124 951
rect 2068 897 2124 899
rect 3624 652 3680 654
rect 3624 600 3626 652
rect 3626 600 3678 652
rect 3678 600 3680 652
rect 3624 598 3680 600
rect 4178 651 4234 653
rect 4178 599 4180 651
rect 4180 599 4232 651
rect 4232 599 4234 651
rect 4178 597 4234 599
rect 4723 652 4779 654
rect 4723 600 4725 652
rect 4725 600 4777 652
rect 4777 600 4779 652
rect 4723 598 4779 600
rect 4968 651 5024 653
rect 4968 599 4970 651
rect 4970 599 5022 651
rect 5022 599 5024 651
rect 4968 597 5024 599
rect 5507 644 5563 646
rect 5507 592 5509 644
rect 5509 592 5561 644
rect 5561 592 5563 644
rect 5507 590 5563 592
rect 6054 651 6110 653
rect 6054 599 6056 651
rect 6056 599 6108 651
rect 6108 599 6110 651
rect 6054 597 6110 599
rect 2641 -137 2697 -134
rect 2641 -189 2645 -137
rect 2645 -189 2697 -137
rect 2641 -190 2697 -189
rect 3640 241 3696 243
rect 3640 189 3642 241
rect 3642 189 3694 241
rect 3694 189 3696 241
rect 3640 187 3696 189
rect 4176 239 4232 241
rect 4176 187 4178 239
rect 4178 187 4230 239
rect 4230 187 4232 239
rect 4176 185 4232 187
rect 4719 239 4775 241
rect 4719 187 4721 239
rect 4721 187 4773 239
rect 4773 187 4775 239
rect 4719 185 4775 187
rect 4953 237 5009 239
rect 4953 185 4955 237
rect 4955 185 5007 237
rect 5007 185 5009 237
rect 4953 183 5009 185
rect 5507 222 5563 224
rect 5507 170 5509 222
rect 5509 170 5561 222
rect 5561 170 5563 222
rect 5507 168 5563 170
rect 6053 239 6109 241
rect 6053 187 6055 239
rect 6055 187 6107 239
rect 6107 187 6109 239
rect 6053 185 6109 187
rect 3641 -174 3697 -172
rect 3641 -226 3643 -174
rect 3643 -226 3695 -174
rect 3695 -226 3697 -174
rect 3641 -228 3697 -226
rect 4175 -193 4231 -191
rect 4175 -245 4177 -193
rect 4177 -245 4229 -193
rect 4229 -245 4231 -193
rect 4175 -247 4231 -245
rect 4719 -133 4775 -131
rect 4719 -185 4721 -133
rect 4721 -185 4773 -133
rect 4773 -185 4775 -133
rect 4719 -187 4775 -185
rect 4962 -142 5018 -140
rect 4962 -194 4964 -142
rect 4964 -194 5016 -142
rect 5016 -194 5018 -142
rect 4962 -196 5018 -194
rect 5506 -176 5562 -174
rect 5506 -228 5508 -176
rect 5508 -228 5560 -176
rect 5560 -228 5562 -176
rect 5506 -230 5562 -228
rect 6046 -195 6102 -193
rect 6046 -247 6048 -195
rect 6048 -247 6100 -195
rect 6100 -247 6102 -195
rect 6046 -249 6102 -247
rect 3632 -585 3688 -583
rect 3632 -637 3634 -585
rect 3634 -637 3686 -585
rect 3686 -637 3688 -585
rect 3632 -639 3688 -637
rect 4174 -598 4230 -596
rect 4174 -650 4176 -598
rect 4176 -650 4228 -598
rect 4228 -650 4230 -598
rect 4174 -652 4230 -650
rect 4731 -587 4787 -585
rect 4731 -639 4733 -587
rect 4733 -639 4785 -587
rect 4785 -639 4787 -587
rect 4731 -641 4787 -639
rect 4967 -590 5023 -588
rect 4967 -642 4969 -590
rect 4969 -642 5021 -590
rect 5021 -642 5023 -590
rect 4967 -644 5023 -642
rect 5496 -591 5552 -589
rect 5496 -643 5498 -591
rect 5498 -643 5550 -591
rect 5550 -643 5552 -591
rect 5496 -645 5552 -643
rect 6046 -628 6102 -626
rect 6046 -680 6048 -628
rect 6048 -680 6100 -628
rect 6100 -680 6102 -628
rect 6046 -682 6102 -680
<< metal3 >>
rect 2037 953 2137 966
rect 2037 897 2068 953
rect 2124 897 2137 953
rect 2037 885 2137 897
rect 3620 899 6257 956
rect 2037 -361 2128 885
rect 3620 747 3677 899
rect 3088 674 3691 747
rect 3088 -117 3161 674
rect 3613 654 3691 674
rect 4729 669 4786 899
rect 3613 598 3624 654
rect 3680 598 3691 654
rect 3613 586 3691 598
rect 4167 653 4245 668
rect 4167 597 4178 653
rect 4234 597 4245 653
rect 4167 568 4245 597
rect 4712 654 4790 669
rect 4712 598 4723 654
rect 4779 598 4790 654
rect 4712 586 4790 598
rect 4957 653 5035 668
rect 5505 661 5562 899
rect 4957 597 4968 653
rect 5024 597 5035 653
rect 4957 585 5035 597
rect 5496 646 5574 661
rect 5496 590 5507 646
rect 5563 590 5574 646
rect 4172 477 4232 568
rect 4964 477 5024 585
rect 5496 578 5574 590
rect 6043 653 6121 668
rect 6043 597 6054 653
rect 6110 597 6121 653
rect 6043 585 6121 597
rect 6051 477 6111 585
rect 3639 417 6111 477
rect 3639 258 3699 417
rect 3629 243 3707 258
rect 4706 256 4766 417
rect 3629 187 3640 243
rect 3696 187 3707 243
rect 3629 175 3707 187
rect 4165 241 4243 256
rect 4165 185 4176 241
rect 4232 185 4243 241
rect 4165 173 4243 185
rect 4706 241 4786 256
rect 4706 185 4719 241
rect 4775 185 4786 241
rect 4706 173 4786 185
rect 4942 239 5020 254
rect 5509 239 5569 417
rect 6042 241 6120 256
rect 4942 183 4953 239
rect 5009 183 5020 239
rect 2621 -125 3161 -117
rect 2619 -127 3161 -125
rect 2614 -134 3161 -127
rect 2614 -190 2641 -134
rect 2697 -190 3161 -134
rect 4181 35 4241 173
rect 4942 171 5020 183
rect 5496 224 5574 239
rect 4953 35 5013 171
rect 5496 168 5507 224
rect 5563 168 5574 224
rect 6042 185 6053 241
rect 6109 185 6120 241
rect 6042 173 6120 185
rect 5496 156 5574 168
rect 6049 53 6109 173
rect 6200 53 6257 899
rect 6049 35 6257 53
rect 4181 -4 6257 35
rect 4181 -25 6109 -4
rect 4181 -138 4241 -25
rect 4708 -131 4786 -116
rect 4953 -125 5013 -25
rect 3630 -172 3708 -157
rect 2614 -206 2729 -190
rect 3630 -228 3641 -172
rect 3697 -228 3708 -172
rect 3630 -257 3708 -228
rect 4164 -191 4242 -138
rect 4164 -247 4175 -191
rect 4231 -247 4242 -191
rect 4708 -187 4719 -131
rect 4775 -187 4786 -131
rect 4708 -199 4786 -187
rect 4951 -140 5029 -125
rect 4951 -196 4962 -140
rect 5018 -196 5029 -140
rect 3635 -361 3692 -257
rect 4164 -259 4242 -247
rect 2037 -379 3692 -361
rect 4713 -379 4770 -199
rect 4951 -208 5029 -196
rect 5495 -174 5573 -159
rect 5495 -230 5506 -174
rect 5562 -230 5573 -174
rect 6049 -178 6109 -25
rect 5495 -242 5573 -230
rect 6035 -193 6113 -178
rect 5507 -379 5564 -242
rect 6035 -249 6046 -193
rect 6102 -249 6113 -193
rect 6035 -261 6113 -249
rect 2037 -436 6107 -379
rect 2037 -452 4230 -436
rect 3621 -583 3699 -568
rect 4173 -581 4230 -452
rect 3621 -639 3632 -583
rect 3688 -639 3699 -583
rect 3621 -697 3699 -639
rect 4163 -596 4241 -581
rect 4163 -652 4174 -596
rect 4230 -652 4241 -596
rect 4163 -664 4241 -652
rect 4720 -585 4798 -570
rect 4965 -573 5022 -436
rect 4720 -641 4731 -585
rect 4787 -641 4798 -585
rect 4720 -653 4798 -641
rect 4956 -588 5034 -573
rect 4956 -644 4967 -588
rect 5023 -644 5034 -588
rect 3641 -843 3699 -697
rect 4733 -843 4791 -653
rect 4956 -656 5034 -644
rect 5485 -589 5563 -574
rect 5485 -645 5496 -589
rect 5552 -645 5563 -589
rect 6050 -611 6107 -436
rect 5485 -657 5563 -645
rect 6035 -626 6113 -611
rect 5498 -843 5556 -657
rect 6035 -682 6046 -626
rect 6102 -682 6113 -626
rect 6035 -694 6113 -682
rect 3641 -901 5556 -843
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_0
timestamp 1713185578
transform 0 1 2309 -1 0 -424
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_1
timestamp 1713185578
transform 1 0 3797 0 1 -606
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_2
timestamp 1713185578
transform 1 0 5945 0 1 -606
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_3
timestamp 1713185578
transform 0 1 2669 -1 0 -424
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_4
timestamp 1713185578
transform 1 0 5945 0 1 -196
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_5
timestamp 1713185578
transform 1 0 5129 0 1 -196
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_6
timestamp 1713185578
transform 0 1 2669 -1 0 792
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_7
timestamp 1713185578
transform 0 1 2669 -1 0 -24
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_8
timestamp 1713185578
transform 0 1 2309 -1 0 -24
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_9
timestamp 1713185578
transform 0 1 2309 -1 0 792
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_10
timestamp 1713185578
transform 1 0 5129 0 1 -606
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_11
timestamp 1713185578
transform 1 0 4613 0 1 -606
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_12
timestamp 1713185578
transform 1 0 4613 0 1 -196
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_13
timestamp 1713185578
transform 1 0 3797 0 1 -196
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_14
timestamp 1713185578
transform 1 0 5129 0 1 214
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_15
timestamp 1713185578
transform 1 0 5945 0 1 214
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_16
timestamp 1713185578
transform 1 0 5129 0 1 624
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_17
timestamp 1713185578
transform 1 0 5945 0 1 624
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_18
timestamp 1713185578
transform 1 0 3797 0 1 214
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_19
timestamp 1713185578
transform 1 0 3797 0 1 624
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_20
timestamp 1713185578
transform 1 0 4613 0 1 214
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_21
timestamp 1713185578
transform 1 0 4613 0 1 624
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_23
timestamp 1713185578
transform 0 -1 2670 1 0 -914
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_24
timestamp 1713185578
transform 0 -1 2306 1 0 -910
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_25
timestamp 1713185578
transform 0 -1 2309 1 0 1221
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_26
timestamp 1713185578
transform 0 -1 2668 1 0 1221
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_27
timestamp 1713185578
transform 1 0 3281 0 1 -609
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_28
timestamp 1713185578
transform 1 0 3281 0 1 624
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_29
timestamp 1713185578
transform 1 0 3277 0 1 210
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_30
timestamp 1713185578
transform 1 0 3279 0 1 -198
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_31
timestamp 1713185578
transform 1 0 6499 0 1 -606
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_32
timestamp 1713185578
transform 1 0 6497 0 1 626
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_33
timestamp 1713185578
transform 1 0 6497 0 1 216
box -258 -180 258 180
use pmos_3p3_HMKTA7  pmos_3p3_HMKTA7_34
timestamp 1713185578
transform 1 0 6497 0 1 -196
box -258 -180 258 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_0
timestamp 1713185578
transform 1 0 4205 0 1 -606
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_1
timestamp 1713185578
transform 1 0 5537 0 1 -196
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_2
timestamp 1713185578
transform 0 1 2669 -1 0 384
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_3
timestamp 1713185578
transform 0 1 2309 -1 0 384
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_4
timestamp 1713185578
transform 1 0 5537 0 1 -606
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_5
timestamp 1713185578
transform 1 0 4205 0 1 -196
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_6
timestamp 1713185578
transform 1 0 5537 0 1 214
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_7
timestamp 1713185578
transform 1 0 5537 0 1 624
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_8
timestamp 1713185578
transform 1 0 4205 0 1 214
box -394 -180 394 180
use pmos_3p3_HVHTA7  pmos_3p3_HVHTA7_9
timestamp 1713185578
transform 1 0 4205 0 1 624
box -394 -180 394 180
<< labels >>
flabel metal1 s 2710 935 2710 935 0 FreeSans 625 90 0 0 M2
port 1 nsew
flabel metal1 s 2182 927 2182 927 0 FreeSans 625 90 0 0 M4
port 2 nsew
flabel metal1 s 1483 -706 1483 -706 0 FreeSans 1250 0 0 0 VCTRL
port 3 nsew
<< end >>
