magic
tech gf180mcuC
magscale 1 10
timestamp 1693309239
<< pwell >>
rect -3324 -188 3324 188
<< nmos >>
rect -3212 -120 -3112 120
rect -3008 -120 -2908 120
rect -2804 -120 -2704 120
rect -2600 -120 -2500 120
rect -2396 -120 -2296 120
rect -2192 -120 -2092 120
rect -1988 -120 -1888 120
rect -1784 -120 -1684 120
rect -1580 -120 -1480 120
rect -1376 -120 -1276 120
rect -1172 -120 -1072 120
rect -968 -120 -868 120
rect -764 -120 -664 120
rect -560 -120 -460 120
rect -356 -120 -256 120
rect -152 -120 -52 120
rect 52 -120 152 120
rect 256 -120 356 120
rect 460 -120 560 120
rect 664 -120 764 120
rect 868 -120 968 120
rect 1072 -120 1172 120
rect 1276 -120 1376 120
rect 1480 -120 1580 120
rect 1684 -120 1784 120
rect 1888 -120 1988 120
rect 2092 -120 2192 120
rect 2296 -120 2396 120
rect 2500 -120 2600 120
rect 2704 -120 2804 120
rect 2908 -120 3008 120
rect 3112 -120 3212 120
<< ndiff >>
rect -3300 107 -3212 120
rect -3300 -107 -3287 107
rect -3241 -107 -3212 107
rect -3300 -120 -3212 -107
rect -3112 107 -3008 120
rect -3112 -107 -3083 107
rect -3037 -107 -3008 107
rect -3112 -120 -3008 -107
rect -2908 107 -2804 120
rect -2908 -107 -2879 107
rect -2833 -107 -2804 107
rect -2908 -120 -2804 -107
rect -2704 107 -2600 120
rect -2704 -107 -2675 107
rect -2629 -107 -2600 107
rect -2704 -120 -2600 -107
rect -2500 107 -2396 120
rect -2500 -107 -2471 107
rect -2425 -107 -2396 107
rect -2500 -120 -2396 -107
rect -2296 107 -2192 120
rect -2296 -107 -2267 107
rect -2221 -107 -2192 107
rect -2296 -120 -2192 -107
rect -2092 107 -1988 120
rect -2092 -107 -2063 107
rect -2017 -107 -1988 107
rect -2092 -120 -1988 -107
rect -1888 107 -1784 120
rect -1888 -107 -1859 107
rect -1813 -107 -1784 107
rect -1888 -120 -1784 -107
rect -1684 107 -1580 120
rect -1684 -107 -1655 107
rect -1609 -107 -1580 107
rect -1684 -120 -1580 -107
rect -1480 107 -1376 120
rect -1480 -107 -1451 107
rect -1405 -107 -1376 107
rect -1480 -120 -1376 -107
rect -1276 107 -1172 120
rect -1276 -107 -1247 107
rect -1201 -107 -1172 107
rect -1276 -120 -1172 -107
rect -1072 107 -968 120
rect -1072 -107 -1043 107
rect -997 -107 -968 107
rect -1072 -120 -968 -107
rect -868 107 -764 120
rect -868 -107 -839 107
rect -793 -107 -764 107
rect -868 -120 -764 -107
rect -664 107 -560 120
rect -664 -107 -635 107
rect -589 -107 -560 107
rect -664 -120 -560 -107
rect -460 107 -356 120
rect -460 -107 -431 107
rect -385 -107 -356 107
rect -460 -120 -356 -107
rect -256 107 -152 120
rect -256 -107 -227 107
rect -181 -107 -152 107
rect -256 -120 -152 -107
rect -52 107 52 120
rect -52 -107 -23 107
rect 23 -107 52 107
rect -52 -120 52 -107
rect 152 107 256 120
rect 152 -107 181 107
rect 227 -107 256 107
rect 152 -120 256 -107
rect 356 107 460 120
rect 356 -107 385 107
rect 431 -107 460 107
rect 356 -120 460 -107
rect 560 107 664 120
rect 560 -107 589 107
rect 635 -107 664 107
rect 560 -120 664 -107
rect 764 107 868 120
rect 764 -107 793 107
rect 839 -107 868 107
rect 764 -120 868 -107
rect 968 107 1072 120
rect 968 -107 997 107
rect 1043 -107 1072 107
rect 968 -120 1072 -107
rect 1172 107 1276 120
rect 1172 -107 1201 107
rect 1247 -107 1276 107
rect 1172 -120 1276 -107
rect 1376 107 1480 120
rect 1376 -107 1405 107
rect 1451 -107 1480 107
rect 1376 -120 1480 -107
rect 1580 107 1684 120
rect 1580 -107 1609 107
rect 1655 -107 1684 107
rect 1580 -120 1684 -107
rect 1784 107 1888 120
rect 1784 -107 1813 107
rect 1859 -107 1888 107
rect 1784 -120 1888 -107
rect 1988 107 2092 120
rect 1988 -107 2017 107
rect 2063 -107 2092 107
rect 1988 -120 2092 -107
rect 2192 107 2296 120
rect 2192 -107 2221 107
rect 2267 -107 2296 107
rect 2192 -120 2296 -107
rect 2396 107 2500 120
rect 2396 -107 2425 107
rect 2471 -107 2500 107
rect 2396 -120 2500 -107
rect 2600 107 2704 120
rect 2600 -107 2629 107
rect 2675 -107 2704 107
rect 2600 -120 2704 -107
rect 2804 107 2908 120
rect 2804 -107 2833 107
rect 2879 -107 2908 107
rect 2804 -120 2908 -107
rect 3008 107 3112 120
rect 3008 -107 3037 107
rect 3083 -107 3112 107
rect 3008 -120 3112 -107
rect 3212 107 3300 120
rect 3212 -107 3241 107
rect 3287 -107 3300 107
rect 3212 -120 3300 -107
<< ndiffc >>
rect -3287 -107 -3241 107
rect -3083 -107 -3037 107
rect -2879 -107 -2833 107
rect -2675 -107 -2629 107
rect -2471 -107 -2425 107
rect -2267 -107 -2221 107
rect -2063 -107 -2017 107
rect -1859 -107 -1813 107
rect -1655 -107 -1609 107
rect -1451 -107 -1405 107
rect -1247 -107 -1201 107
rect -1043 -107 -997 107
rect -839 -107 -793 107
rect -635 -107 -589 107
rect -431 -107 -385 107
rect -227 -107 -181 107
rect -23 -107 23 107
rect 181 -107 227 107
rect 385 -107 431 107
rect 589 -107 635 107
rect 793 -107 839 107
rect 997 -107 1043 107
rect 1201 -107 1247 107
rect 1405 -107 1451 107
rect 1609 -107 1655 107
rect 1813 -107 1859 107
rect 2017 -107 2063 107
rect 2221 -107 2267 107
rect 2425 -107 2471 107
rect 2629 -107 2675 107
rect 2833 -107 2879 107
rect 3037 -107 3083 107
rect 3241 -107 3287 107
<< polysilicon >>
rect -3212 120 -3112 164
rect -3008 120 -2908 164
rect -2804 120 -2704 164
rect -2600 120 -2500 164
rect -2396 120 -2296 164
rect -2192 120 -2092 164
rect -1988 120 -1888 164
rect -1784 120 -1684 164
rect -1580 120 -1480 164
rect -1376 120 -1276 164
rect -1172 120 -1072 164
rect -968 120 -868 164
rect -764 120 -664 164
rect -560 120 -460 164
rect -356 120 -256 164
rect -152 120 -52 164
rect 52 120 152 164
rect 256 120 356 164
rect 460 120 560 164
rect 664 120 764 164
rect 868 120 968 164
rect 1072 120 1172 164
rect 1276 120 1376 164
rect 1480 120 1580 164
rect 1684 120 1784 164
rect 1888 120 1988 164
rect 2092 120 2192 164
rect 2296 120 2396 164
rect 2500 120 2600 164
rect 2704 120 2804 164
rect 2908 120 3008 164
rect 3112 120 3212 164
rect -3212 -164 -3112 -120
rect -3008 -164 -2908 -120
rect -2804 -164 -2704 -120
rect -2600 -164 -2500 -120
rect -2396 -164 -2296 -120
rect -2192 -164 -2092 -120
rect -1988 -164 -1888 -120
rect -1784 -164 -1684 -120
rect -1580 -164 -1480 -120
rect -1376 -164 -1276 -120
rect -1172 -164 -1072 -120
rect -968 -164 -868 -120
rect -764 -164 -664 -120
rect -560 -164 -460 -120
rect -356 -164 -256 -120
rect -152 -164 -52 -120
rect 52 -164 152 -120
rect 256 -164 356 -120
rect 460 -164 560 -120
rect 664 -164 764 -120
rect 868 -164 968 -120
rect 1072 -164 1172 -120
rect 1276 -164 1376 -120
rect 1480 -164 1580 -120
rect 1684 -164 1784 -120
rect 1888 -164 1988 -120
rect 2092 -164 2192 -120
rect 2296 -164 2396 -120
rect 2500 -164 2600 -120
rect 2704 -164 2804 -120
rect 2908 -164 3008 -120
rect 3112 -164 3212 -120
<< metal1 >>
rect -3287 107 -3241 118
rect -3287 -118 -3241 -107
rect -3083 107 -3037 118
rect -3083 -118 -3037 -107
rect -2879 107 -2833 118
rect -2879 -118 -2833 -107
rect -2675 107 -2629 118
rect -2675 -118 -2629 -107
rect -2471 107 -2425 118
rect -2471 -118 -2425 -107
rect -2267 107 -2221 118
rect -2267 -118 -2221 -107
rect -2063 107 -2017 118
rect -2063 -118 -2017 -107
rect -1859 107 -1813 118
rect -1859 -118 -1813 -107
rect -1655 107 -1609 118
rect -1655 -118 -1609 -107
rect -1451 107 -1405 118
rect -1451 -118 -1405 -107
rect -1247 107 -1201 118
rect -1247 -118 -1201 -107
rect -1043 107 -997 118
rect -1043 -118 -997 -107
rect -839 107 -793 118
rect -839 -118 -793 -107
rect -635 107 -589 118
rect -635 -118 -589 -107
rect -431 107 -385 118
rect -431 -118 -385 -107
rect -227 107 -181 118
rect -227 -118 -181 -107
rect -23 107 23 118
rect -23 -118 23 -107
rect 181 107 227 118
rect 181 -118 227 -107
rect 385 107 431 118
rect 385 -118 431 -107
rect 589 107 635 118
rect 589 -118 635 -107
rect 793 107 839 118
rect 793 -118 839 -107
rect 997 107 1043 118
rect 997 -118 1043 -107
rect 1201 107 1247 118
rect 1201 -118 1247 -107
rect 1405 107 1451 118
rect 1405 -118 1451 -107
rect 1609 107 1655 118
rect 1609 -118 1655 -107
rect 1813 107 1859 118
rect 1813 -118 1859 -107
rect 2017 107 2063 118
rect 2017 -118 2063 -107
rect 2221 107 2267 118
rect 2221 -118 2267 -107
rect 2425 107 2471 118
rect 2425 -118 2471 -107
rect 2629 107 2675 118
rect 2629 -118 2675 -107
rect 2833 107 2879 118
rect 2833 -118 2879 -107
rect 3037 107 3083 118
rect 3037 -118 3083 -107
rect 3241 107 3287 118
rect 3241 -118 3287 -107
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1.2 l 0.5 m 1 nf 32 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
