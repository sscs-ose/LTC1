* NGSPICE file created from Delay_Cell_flat.ext - technology: gf180mcuC

.subckt Delay_Cell_PEX VDD VSS VCONT IN INB OUT OUTB EN 
X0 a_667_n765# EN.t0 VSS.t4 VSS.t3 nfet_03v3 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.56u
X1 VDD OUTB.t4 OUT.t0 VDD.t1 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X2 VDD a_86_130# a_86_130# VDD.t6 pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.56u
X3 OUTB OUT.t4 VDD.t11 VDD.t10 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X4 a_502_130# a_86_130# VDD.t5 VDD.t4 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X5 a_502_130# OUTB.t0 OUTB.t1 VDD.t0 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.56u
X6 a_86_130# VCONT.t0 VSS.t6 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X7 OUTB INB.t0 a_667_n765# VSS.t7 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X8 a_667_n765# IN.t0 OUT.t3 VSS.t11 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X9 OUT OUT.t1 a_502_130# VDD.t9 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X10 VSS VCONT.t1 a_86_130# VSS.t8 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X11 VSS EN.t1 a_667_n765# VSS.t0 nfet_03v3 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.56u
R0 EN EN.t1 13.1944
R1 EN EN.t0 13.1748
R2 VSS.n90 VSS.n89 231.117
R3 VSS.n38 VSS.t11 207.873
R4 VSS.n35 VSS.t7 163.899
R5 VSS.n6 VSS.n5 154.945
R6 VSS.n142 VSS.t5 123.924
R7 VSS.n139 VSS.t8 79.9513
R8 VSS.n44 VSS.t0 55.9661
R9 VSS.n27 VSS.n26 39.9759
R10 VSS.n112 VSS.n111 31.9808
R11 VSS.n47 VSS.t3 11.9931
R12 VSS.n1 VSS.n0 6.267
R13 VSS.n1 VSS.t4 5.44487
R14 VSS.n109 VSS.n108 4.26137
R15 VSS.n29 VSS.n25 4.26137
R16 VSS.n4 VSS.t6 3.07947
R17 VSS.n3 VSS.n2 3.06207
R18 VSS.n4 VSS.n3 2.83323
R19 VSS.n120 VSS.n119 2.60211
R20 VSS.n150 VSS.n149 2.60211
R21 VSS.n61 VSS.n60 2.6005
R22 VSS.n60 VSS.n59 2.6005
R23 VSS.n34 VSS.n33 2.6005
R24 VSS.n33 VSS.n32 2.6005
R25 VSS.n37 VSS.n36 2.6005
R26 VSS.n36 VSS.n35 2.6005
R27 VSS.n40 VSS.n39 2.6005
R28 VSS.n39 VSS.n38 2.6005
R29 VSS.n43 VSS.n42 2.6005
R30 VSS.n42 VSS.n41 2.6005
R31 VSS.n46 VSS.n45 2.6005
R32 VSS.n45 VSS.n44 2.6005
R33 VSS.n49 VSS.n48 2.6005
R34 VSS.n48 VSS.n47 2.6005
R35 VSS.n52 VSS.n51 2.6005
R36 VSS.n51 VSS.n50 2.6005
R37 VSS.n55 VSS.n54 2.6005
R38 VSS.n54 VSS.n53 2.6005
R39 VSS.n58 VSS.n57 2.6005
R40 VSS.n57 VSS.n56 2.6005
R41 VSS.n64 VSS.n63 2.6005
R42 VSS.n63 VSS.n62 2.6005
R43 VSS.n67 VSS.n66 2.6005
R44 VSS.n66 VSS.n65 2.6005
R45 VSS.n70 VSS.n69 2.6005
R46 VSS.n69 VSS.n68 2.6005
R47 VSS.n73 VSS.n72 2.6005
R48 VSS.n72 VSS.n71 2.6005
R49 VSS.n76 VSS.n75 2.6005
R50 VSS.n75 VSS.n74 2.6005
R51 VSS.n79 VSS.n78 2.6005
R52 VSS.n78 VSS.n77 2.6005
R53 VSS.n82 VSS.n81 2.6005
R54 VSS.n81 VSS.n80 2.6005
R55 VSS.n85 VSS.n84 2.6005
R56 VSS.n84 VSS.n83 2.6005
R57 VSS.n88 VSS.n87 2.6005
R58 VSS.n87 VSS.n86 2.6005
R59 VSS.n22 VSS.n21 2.6005
R60 VSS.n21 VSS.n20 2.6005
R61 VSS.n19 VSS.n18 2.6005
R62 VSS.n18 VSS.n17 2.6005
R63 VSS.n16 VSS.n15 2.6005
R64 VSS.n15 VSS.n14 2.6005
R65 VSS.n13 VSS.n12 2.6005
R66 VSS.n12 VSS.n11 2.6005
R67 VSS.n10 VSS.n9 2.6005
R68 VSS.n9 VSS.n8 2.6005
R69 VSS.n24 VSS.n23 2.6005
R70 VSS.n117 VSS.n116 2.6005
R71 VSS.n30 VSS.n29 2.6005
R72 VSS.n7 VSS.n6 2.6005
R73 VSS.n123 VSS.n122 2.6005
R74 VSS.n122 VSS.n121 2.6005
R75 VSS.n126 VSS.n125 2.6005
R76 VSS.n125 VSS.n124 2.6005
R77 VSS.n129 VSS.n128 2.6005
R78 VSS.n128 VSS.n127 2.6005
R79 VSS.n132 VSS.n131 2.6005
R80 VSS.n131 VSS.n130 2.6005
R81 VSS.n135 VSS.n134 2.6005
R82 VSS.n134 VSS.n133 2.6005
R83 VSS.n138 VSS.n137 2.6005
R84 VSS.n137 VSS.n136 2.6005
R85 VSS.n141 VSS.n140 2.6005
R86 VSS.n140 VSS.n139 2.6005
R87 VSS.n144 VSS.n143 2.6005
R88 VSS.n143 VSS.n142 2.6005
R89 VSS.n147 VSS.n146 2.6005
R90 VSS.n146 VSS.n145 2.6005
R91 VSS.n115 VSS.n114 2.6005
R92 VSS.n152 VSS.n151 2.6005
R93 VSS.n110 VSS.n109 2.6005
R94 VSS.n97 VSS.n96 2.6005
R95 VSS.n96 VSS.n95 2.6005
R96 VSS.n100 VSS.n99 2.6005
R97 VSS.n99 VSS.n98 2.6005
R98 VSS.n103 VSS.n102 2.6005
R99 VSS.n102 VSS.n101 2.6005
R100 VSS.n106 VSS.n105 2.6005
R101 VSS.n105 VSS.n104 2.6005
R102 VSS.n94 VSS.n93 2.6005
R103 VSS.n93 VSS.n92 2.6005
R104 VSS.n91 VSS.n90 2.6005
R105 VSS.n114 VSS.n113 1.95163
R106 VSS.n29 VSS.n28 1.951
R107 VSS.n3 VSS.n1 0.45756
R108 VSS.n28 VSS.n27 0.32628
R109 VSS.n113 VSS.n112 0.32628
R110 VSS.n94 VSS.n91 0.200589
R111 VSS.n10 VSS.n7 0.198982
R112 VSS.n126 VSS.n123 0.181382
R113 VSS.n129 VSS.n126 0.181382
R114 VSS.n132 VSS.n129 0.181382
R115 VSS.n135 VSS.n132 0.181382
R116 VSS.n138 VSS.n135 0.181382
R117 VSS.n141 VSS.n138 0.181382
R118 VSS.n144 VSS.n141 0.181382
R119 VSS.n147 VSS.n144 0.181382
R120 VSS.n37 VSS.n34 0.179626
R121 VSS.n40 VSS.n37 0.179626
R122 VSS.n43 VSS.n40 0.179626
R123 VSS.n46 VSS.n43 0.179626
R124 VSS.n49 VSS.n46 0.179626
R125 VSS.n52 VSS.n49 0.179626
R126 VSS.n55 VSS.n52 0.179626
R127 VSS.n58 VSS.n55 0.179626
R128 VSS.n61 VSS.n58 0.179626
R129 VSS.n67 VSS.n64 0.179626
R130 VSS.n70 VSS.n67 0.179626
R131 VSS.n73 VSS.n70 0.179626
R132 VSS.n76 VSS.n73 0.179626
R133 VSS.n79 VSS.n76 0.179626
R134 VSS.n82 VSS.n79 0.179626
R135 VSS.n85 VSS.n82 0.179626
R136 VSS.n88 VSS.n85 0.179626
R137 VSS VSS.n4 0.170912
R138 VSS.n13 VSS.n10 0.165232
R139 VSS.n16 VSS.n13 0.165232
R140 VSS.n19 VSS.n16 0.165232
R141 VSS.n22 VSS.n19 0.165232
R142 VSS.n30 VSS.n24 0.165232
R143 VSS.n97 VSS.n94 0.165232
R144 VSS.n100 VSS.n97 0.165232
R145 VSS.n103 VSS.n100 0.165232
R146 VSS.n106 VSS.n103 0.165232
R147 VSS.n115 VSS.n110 0.165232
R148 VSS.n120 VSS.n117 0.163625
R149 VSS.n152 VSS.n150 0.163625
R150 VSS.n123 VSS.n120 0.154029
R151 VSS VSS.n153 0.1445
R152 VSS.n150 VSS.n147 0.130206
R153 VSS.n91 VSS.n88 0.128073
R154 VSS.n31 VSS.n22 0.120232
R155 VSS.n107 VSS.n106 0.120232
R156 VSS.n153 VSS.n115 0.0953214
R157 VSS.n149 VSS.n148 0.076587
R158 VSS.n119 VSS.n118 0.076587
R159 VSS.n153 VSS.n152 0.0704107
R160 VSS.n34 VSS.n31 0.0511796
R161 VSS.n107 VSS.n61 0.0511796
R162 VSS.n31 VSS.n30 0.0455
R163 VSS.n110 VSS.n107 0.0455
R164 OUTB.n3 OUTB.t4 21.1283
R165 OUTB.n4 OUTB.t0 20.6862
R166 OUTB.n5 OUTB.n0 10.6918
R167 OUTB.n3 OUTB.n2 2.85009
R168 OUTB.n2 OUTB.t1 0.9105
R169 OUTB.n2 OUTB.n1 0.9105
R170 OUTB OUTB.n5 0.0611522
R171 OUTB.n5 OUTB.n4 0.0458582
R172 OUTB.n4 OUTB.n3 0.0448662
R173 OUT.n0 OUT.t4 21.2967
R174 OUT.n0 OUT.t1 20.6887
R175 OUT OUT.t3 11.0126
R176 OUT.n3 OUT.n2 2.6005
R177 OUT.n2 OUT.t0 0.9105
R178 OUT.n2 OUT.n1 0.9105
R179 OUT OUT.n3 0.26932
R180 OUT.n3 OUT.n0 0.196036
R181 VDD.n22 VDD.t0 57.1978
R182 VDD.n37 VDD.t4 52.4314
R183 VDD.n75 VDD.t9 47.6649
R184 VDD.n25 VDD.t10 20.9729
R185 VDD.n40 VDD.t6 20.0196
R186 VDD.n72 VDD.t1 10.4867
R187 VDD.n4 VDD.n3 3.43154
R188 VDD.n48 VDD.n47 3.15124
R189 VDD.n39 VDD.n38 3.1505
R190 VDD.n38 VDD.n37 3.1505
R191 VDD.n21 VDD.n20 3.1505
R192 VDD.n20 VDD.n19 3.1505
R193 VDD.n24 VDD.n23 3.1505
R194 VDD.n23 VDD.n22 3.1505
R195 VDD.n27 VDD.n26 3.1505
R196 VDD.n26 VDD.n25 3.1505
R197 VDD.n30 VDD.n29 3.1505
R198 VDD.n29 VDD.n28 3.1505
R199 VDD.n33 VDD.n32 3.1505
R200 VDD.n32 VDD.n31 3.1505
R201 VDD.n36 VDD.n35 3.1505
R202 VDD.n35 VDD.n34 3.1505
R203 VDD.n42 VDD.n41 3.1505
R204 VDD.n41 VDD.n40 3.1505
R205 VDD.n45 VDD.n44 3.1505
R206 VDD.n44 VDD.n43 3.1505
R207 VDD.n14 VDD.n7 3.1505
R208 VDD.n58 VDD.n57 3.1505
R209 VDD.n55 VDD.n54 3.1505
R210 VDD.n11 VDD.n10 3.1505
R211 VDD.n13 VDD.n12 3.1505
R212 VDD.n62 VDD.n61 3.1505
R213 VDD.n61 VDD.n60 3.1505
R214 VDD.n18 VDD.n17 3.1505
R215 VDD.n17 VDD.n16 3.1505
R216 VDD.n83 VDD.n82 3.1505
R217 VDD.n82 VDD.n81 3.1505
R218 VDD.n89 VDD.n88 3.1505
R219 VDD.n88 VDD.n87 3.1505
R220 VDD.n65 VDD.n64 3.1505
R221 VDD.n64 VDD.n63 3.1505
R222 VDD.n68 VDD.n67 3.1505
R223 VDD.n67 VDD.n66 3.1505
R224 VDD.n71 VDD.n70 3.1505
R225 VDD.n70 VDD.n69 3.1505
R226 VDD.n74 VDD.n73 3.1505
R227 VDD.n73 VDD.n72 3.1505
R228 VDD.n77 VDD.n76 3.1505
R229 VDD.n76 VDD.n75 3.1505
R230 VDD.n80 VDD.n79 3.1505
R231 VDD.n79 VDD.n78 3.1505
R232 VDD.n86 VDD.n85 3.1505
R233 VDD.n85 VDD.n84 3.1505
R234 VDD.n53 VDD.n52 3.1505
R235 VDD.n100 VDD.n99 3.1505
R236 VDD.n96 VDD.n95 3.1505
R237 VDD.n94 VDD.n93 3.1505
R238 VDD.n50 VDD.n49 3.1505
R239 VDD.n92 VDD.n91 3.1505
R240 VDD.n91 VDD.n90 3.1505
R241 VDD.n47 VDD.n46 3.1505
R242 VDD VDD.n4 2.88121
R243 VDD.n4 VDD.n1 2.42843
R244 VDD.n57 VDD.n56 2.26657
R245 VDD.n99 VDD.n98 2.22072
R246 VDD.n52 VDD.n51 2.11587
R247 VDD.n10 VDD.n8 1.98264
R248 VDD.n7 VDD.n6 1.87092
R249 VDD.n10 VDD.n9 1.29756
R250 VDD.n1 VDD.t5 0.9105
R251 VDD.n1 VDD.n0 0.9105
R252 VDD.n3 VDD.t11 0.9105
R253 VDD.n3 VDD.n2 0.9105
R254 VDD.n6 VDD.n5 0.854386
R255 VDD.n61 VDD.n59 0.467167
R256 VDD.n98 VDD.n97 0.46673
R257 VDD.n42 VDD.n39 0.135872
R258 VDD.n86 VDD.n83 0.135872
R259 VDD.n36 VDD.n33 0.133641
R260 VDD.n80 VDD.n77 0.133641
R261 VDD.n24 VDD.n21 0.132897
R262 VDD.n27 VDD.n24 0.132897
R263 VDD.n30 VDD.n27 0.132897
R264 VDD.n68 VDD.n65 0.132897
R265 VDD.n71 VDD.n68 0.132897
R266 VDD.n74 VDD.n71 0.132897
R267 VDD.n33 VDD.n30 0.132153
R268 VDD.n77 VDD.n74 0.132153
R269 VDD VDD.n101 0.131
R270 VDD.n58 VDD.n55 0.128861
R271 VDD.n100 VDD.n96 0.128861
R272 VDD.n96 VDD.n94 0.128861
R273 VDD.n13 VDD.n11 0.128123
R274 VDD.n45 VDD.n42 0.126946
R275 VDD.n89 VDD.n86 0.126946
R276 VDD.n101 VDD.n53 0.113369
R277 VDD.n14 VDD.n13 0.110418
R278 VDD.n53 VDD.n50 0.110418
R279 VDD.n39 VDD.n36 0.109839
R280 VDD.n83 VDD.n80 0.109839
R281 VDD.n48 VDD.n45 0.100169
R282 VDD.n92 VDD.n89 0.0971881
R283 VDD.n94 VDD.n92 0.0853361
R284 VDD.n62 VDD.n58 0.0816475
R285 VDD.n18 VDD.n14 0.0794344
R286 VDD.n17 VDD.n15 0.0782778
R287 VDD.n50 VDD.n48 0.0750082
R288 VDD.n65 VDD.n62 0.068186
R289 VDD.n21 VDD.n18 0.0644669
R290 VDD.n101 VDD.n100 0.0152541
R291 VCONT VCONT.t1 14.3672
R292 VCONT VCONT.t0 14.3281
R293 INB INB.t0 14.2767
R294 IN IN.t0 14.2771
C0 OUT a_86_130# 0.12f
C1 a_667_n765# EN 0.0983f
C2 a_667_n765# OUTB 0.058f
C3 EN OUTB 0.00122f
C4 IN OUT 0.01f
C5 OUT VCONT 3.14e-20
C6 a_667_n765# a_502_130# 0.0117f
C7 a_667_n765# VDD 0.00461f
C8 EN a_502_130# 4.03e-19
C9 OUTB a_502_130# 0.307f
C10 VCONT a_86_130# 0.0632f
C11 a_667_n765# INB 0.0188f
C12 VDD EN 0.00648f
C13 VDD OUTB 1.11f
C14 IN VCONT 8.86e-19
C15 INB OUTB 0.0123f
C16 VDD a_502_130# 0.654f
C17 INB a_502_130# 7.89e-19
C18 VDD INB 0.00406f
C19 a_667_n765# OUT 0.164f
C20 EN OUT 0.00964f
C21 OUT OUTB 0.259f
C22 a_667_n765# a_86_130# 3.09e-20
C23 EN a_86_130# 9.47e-20
C24 OUT a_502_130# 0.47f
C25 OUTB a_86_130# 6.04e-19
C26 a_667_n765# IN 0.0232f
C27 a_667_n765# VCONT 8.19e-20
C28 VDD OUT 1.27f
C29 EN IN 0.017f
C30 EN VCONT 0.0155f
C31 IN OUTB 0.00173f
C32 INB OUT 0.00118f
C33 a_86_130# a_502_130# 0.0116f
C34 VDD a_86_130# 1.22f
C35 IN a_502_130# 8.21e-19
C36 VDD IN 0.00413f
C37 VDD VCONT 0.0094f
C38 IN INB 0.0543f
.ends

