magic
tech gf180mcuC
magscale 1 10
timestamp 1693477706
<< nwell >>
rect -296 -270 296 270
<< pmos >>
rect -122 -140 -52 140
rect 52 -140 122 140
<< pdiff >>
rect -210 127 -122 140
rect -210 -127 -197 127
rect -151 -127 -122 127
rect -210 -140 -122 -127
rect -52 127 52 140
rect -52 -127 -23 127
rect 23 -127 52 127
rect -52 -140 52 -127
rect 122 127 210 140
rect 122 -127 151 127
rect 197 -127 210 127
rect 122 -140 210 -127
<< pdiffc >>
rect -197 -127 -151 127
rect -23 -127 23 127
rect 151 -127 197 127
<< polysilicon >>
rect -122 140 -52 184
rect 52 140 122 184
rect -122 -184 -52 -140
rect 52 -184 122 -140
<< metal1 >>
rect -197 127 -151 138
rect -197 -138 -151 -127
rect -23 127 23 138
rect -23 -138 23 -127
rect 151 127 197 138
rect 151 -138 197 -127
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 1.4 l 0.35 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
