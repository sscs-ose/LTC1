magic
tech gf180mcuC
magscale 1 10
timestamp 1689999765
<< nwell >>
rect 20 676 828 754
rect 20 287 1232 676
rect 828 254 1232 287
rect 828 235 1032 254
<< pwell >>
rect 82 10 766 246
rect 886 11 1174 209
<< nmos >>
rect 194 78 250 178
rect 598 78 654 178
rect 1002 85 1058 135
<< pmos >>
rect 194 417 250 517
rect 598 417 654 517
rect 1002 384 1058 484
<< ndiff >>
rect 106 165 194 178
rect 106 91 119 165
rect 165 91 194 165
rect 106 78 194 91
rect 250 165 338 178
rect 250 91 279 165
rect 325 91 338 165
rect 250 78 338 91
rect 510 165 598 178
rect 510 91 523 165
rect 569 91 598 165
rect 510 78 598 91
rect 654 165 742 178
rect 654 91 683 165
rect 729 91 742 165
rect 654 78 742 91
rect 910 135 982 146
rect 1078 135 1150 146
rect 910 133 1002 135
rect 910 87 923 133
rect 969 87 1002 133
rect 910 85 1002 87
rect 1058 133 1150 135
rect 1058 87 1091 133
rect 1137 87 1150 133
rect 1058 85 1150 87
rect 910 74 982 85
rect 1078 74 1150 85
<< pdiff >>
rect 106 504 194 517
rect 106 430 119 504
rect 165 430 194 504
rect 106 417 194 430
rect 250 504 338 517
rect 250 430 279 504
rect 325 430 338 504
rect 250 417 338 430
rect 510 504 598 517
rect 510 430 523 504
rect 569 430 598 504
rect 510 417 598 430
rect 654 504 742 517
rect 654 430 683 504
rect 729 430 742 504
rect 654 417 742 430
rect 914 471 1002 484
rect 914 397 927 471
rect 973 397 1002 471
rect 914 384 1002 397
rect 1058 471 1146 484
rect 1058 397 1087 471
rect 1133 397 1146 471
rect 1058 384 1146 397
<< ndiffc >>
rect 119 91 165 165
rect 279 91 325 165
rect 523 91 569 165
rect 683 91 729 165
rect 923 87 969 133
rect 1091 87 1137 133
<< pdiffc >>
rect 119 430 165 504
rect 279 430 325 504
rect 523 430 569 504
rect 683 430 729 504
rect 927 397 973 471
rect 1087 397 1133 471
<< psubdiff >>
rect 46 -46 873 -40
rect 46 -54 1202 -46
rect 46 -100 69 -54
rect 776 -59 1202 -54
rect 776 -100 873 -59
rect 46 -108 873 -100
rect 1182 -108 1202 -59
rect 46 -113 1202 -108
rect 797 -116 1202 -113
rect 854 -123 1202 -116
<< nsubdiff >>
rect 49 714 790 729
rect 49 662 70 714
rect 769 662 790 714
rect 49 645 790 662
rect 868 632 1160 649
rect 868 581 888 632
rect 1138 581 1160 632
rect 868 564 1160 581
<< psubdiffcont >>
rect 69 -100 776 -54
rect 873 -108 1182 -59
<< nsubdiffcont >>
rect 70 662 769 714
rect 888 581 1138 632
<< polysilicon >>
rect 194 517 250 561
rect 598 517 654 561
rect -18 429 71 442
rect -18 370 -5 429
rect 58 391 71 429
rect 1002 484 1058 528
rect 194 391 250 417
rect 58 370 250 391
rect -18 355 250 370
rect 194 178 250 355
rect 383 281 472 294
rect 383 222 396 281
rect 459 244 472 281
rect 598 244 654 417
rect 1002 322 1058 384
rect 459 222 654 244
rect 943 308 1058 322
rect 943 249 957 308
rect 1020 249 1058 308
rect 943 235 1058 249
rect 383 207 654 222
rect 598 178 654 207
rect 1002 135 1058 235
rect 194 34 250 78
rect 598 34 654 78
rect 1002 41 1058 85
<< polycontact >>
rect -5 370 58 429
rect 396 222 459 281
rect 957 249 1020 308
<< metal1 >>
rect 20 714 1232 754
rect 20 662 70 714
rect 769 662 1232 714
rect 20 636 1232 662
rect 119 504 165 636
rect -18 429 71 442
rect -18 370 -5 429
rect 58 370 71 429
rect 119 419 165 430
rect 279 504 325 515
rect 523 504 569 515
rect 325 449 523 495
rect 279 419 325 430
rect -18 355 71 370
rect 523 363 569 430
rect 683 504 729 636
rect 828 632 1232 636
rect 828 581 888 632
rect 1138 581 1232 632
rect 828 563 1232 581
rect 683 419 729 430
rect 904 471 974 563
rect 904 397 927 471
rect 973 397 974 471
rect 904 382 974 397
rect 1086 471 1150 484
rect 1086 397 1087 471
rect 1133 397 1150 471
rect 523 317 729 363
rect 383 285 472 294
rect -18 281 472 285
rect -18 239 396 281
rect 383 222 396 239
rect 459 222 472 281
rect 383 207 472 222
rect 683 291 729 317
rect 828 308 1032 316
rect 828 291 957 308
rect 683 249 957 291
rect 1020 249 1032 308
rect 683 245 1032 249
rect 119 165 165 176
rect 119 -19 165 91
rect 279 165 325 176
rect 523 165 569 176
rect 325 107 523 153
rect 279 80 325 91
rect 523 80 569 91
rect 683 165 729 245
rect 828 235 1032 245
rect 1086 281 1150 397
rect 1086 234 1263 281
rect 683 80 729 91
rect 901 133 982 138
rect 1086 133 1150 234
rect 901 87 923 133
rect 969 87 982 133
rect 1080 87 1091 133
rect 1137 87 1150 133
rect 20 -24 828 -19
rect 901 -24 982 87
rect 1086 86 1150 87
rect 20 -54 1232 -24
rect 20 -100 69 -54
rect 776 -59 1232 -54
rect 776 -100 873 -59
rect 20 -108 873 -100
rect 1182 -108 1232 -59
rect 20 -137 1232 -108
<< labels >>
flabel nsubdiffcont 363 679 433 702 0 FreeSans 640 0 0 0 VDD
port 1 nsew
flabel psubdiffcont 404 -88 474 -65 0 FreeSans 640 0 0 0 VSS
port 2 nsew
flabel metal1 21 255 91 278 0 FreeSans 640 0 0 0 B
port 4 nsew
flabel polycontact 20 400 20 400 0 FreeSans 640 0 0 0 A
port 6 nsew
flabel metal1 1240 260 1240 260 0 FreeSans 640 0 0 0 OUT
port 7 nsew
flabel nsubdiffcont 1013 607 1013 607 0 FreeSans 640 0 0 0 Inverter_0.VDD
flabel psubdiffcont 1027 -85 1027 -85 0 FreeSans 640 0 0 0 Inverter_0.VSS
flabel metal1 851 276 851 276 0 FreeSans 640 0 0 0 Inverter_0.IN
flabel metal1 1218 249 1218 249 0 FreeSans 640 0 0 0 Inverter_0.OUT
<< end >>
