magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1161 1019 1161
<< metal2 >>
rect -19 156 19 161
rect -19 128 -14 156
rect 14 128 19 156
rect -19 85 19 128
rect -19 57 -14 85
rect 14 57 19 85
rect -19 14 19 57
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -57 19 -14
rect -19 -85 -14 -57
rect 14 -85 19 -57
rect -19 -128 19 -85
rect -19 -156 -14 -128
rect 14 -156 19 -128
rect -19 -161 19 -156
<< via2 >>
rect -14 128 14 156
rect -14 57 14 85
rect -14 -14 14 14
rect -14 -85 14 -57
rect -14 -156 14 -128
<< metal3 >>
rect -19 156 19 161
rect -19 128 -14 156
rect 14 128 19 156
rect -19 85 19 128
rect -19 57 -14 85
rect 14 57 19 85
rect -19 14 19 57
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -57 19 -14
rect -19 -85 -14 -57
rect 14 -85 19 -57
rect -19 -128 19 -85
rect -19 -156 -14 -128
rect 14 -156 19 -128
rect -19 -161 19 -156
<< end >>
