* NGSPICE file created from pll_1_mag_flat.ext - technology: gf180mcuC

.subckt pll_1_mag_flat IPD_ pd VCO_op_bar IPD+ pu LP_ext VCO_op Vref RST_DIV EN VDD_VCO
+ VDD VSS
X0 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.OUTB.t16 VCO_mag_0.Delay_Cell_mag_0.IN VDD_VCO.t117 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X1 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t448 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2 a_72321_5529# VDD.t688 VSS.t481 VSS.t480 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VCO_op.t8 VDD.t398 VDD.t397 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 LF_mag_0.res_48k_mag_0.B VSS.t433 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X5 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t347 VDD.t346 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 a_68145_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t145 VSS.t144 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X7 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_0.OUT a_65581_17830# VSS.t352 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X8 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t2 VDD.t271 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X9 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t669 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X10 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t494 VDD.t496 VDD.t495 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 a_74333_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t163 VSS.t162 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X12 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_69327_6404# VSS.t249 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X13 VCO_op_bar VCO_mag_0.GF_INV16_1.IN VDD_VCO.t155 VDD_VCO.t154 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.35u
X14 VSS VCO_mag_0.VCONT.t45 a_67077_14631.t11 VSS.t609 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X15 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD.t238 VDD.t230 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X16 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD.t241 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X17 VDD RST_DIV.t0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t598 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X18 a_69891_6404# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t553 VSS.t552 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X19 VSS EN.t0 a_59138_17829# VSS.t547 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X20 VDD_VCO a_67077_18370.t10 a_67077_18370.t11 VDD_VCO.t50 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X21 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 VDD.t594 VDD.t593 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X22 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.CLK VCO_mag_0.VCONT.t38 VSS.t515 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X23 PFD_layout_0.DFF__0.nand2_2.IN2 PFD_layout_0.DFF__0.nand2_1.IN1 a_61538_21913# VSS.t275 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X24 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_64776_7545# VSS.t450 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X25 VDD_VCO VCO_mag_0.GF_INV1_0.OUT VCO_mag_0.GF_INV16_2.IN VDD_VCO.t164 pfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X26 VCO_mag_0.Delay_Cell_mag_0.INB VCO_mag_0.Delay_Cell_mag_2.OUT.t16 VSS.t663 VSS.t662 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X27 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.INB a_65581_14091# VSS.t609 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X28 VSS PFD_layout_0.buffer_loading_mag_1.IN a_62430_23292# VSS.t208 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X29 VDD a_63591_22645# pd.t7 VDD.t206 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X30 a_60147_8532# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t248 VSS.t247 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X31 VCO_mag_0.VCONT a2x1mux_mag_0.SEL LF_mag_0.VCNTL.t19 VSS.t105 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X32 a_63436_4432# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_63276_4432# VSS.t143 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X33 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_73056_7541# VSS.t213 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X34 a_63648_7545# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t497 VSS.t496 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X35 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_67501_6446# VSS.t572 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X36 LF_mag_0.res_48k_mag_0.B VSS.t432 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X37 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t445 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X38 a_73620_7541# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t603 VSS.t602 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X39 VDD RST_DIV.t1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t601 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X40 a_63452_24694# PFD_layout_0.nand2_0.IN1 VDD.t62 VDD.t61 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X41 PFD_layout_0.DFF__0.nand2_1.IN1 PFD_layout_0.DFF__0.CLK VDD.t245 VDD.t244 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X42 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.INB a_58943_20071# VDD_VCO.t33 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X43 a_67618_24851# IPD+.t4 VSS.t151 VSS.t150 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X44 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_1.INB.t16 a_59138_17829# VSS.t542 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X45 VSS CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t330 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X46 LF_mag_0.res_48k_mag_0.B VSS.t431 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X47 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_2.OUT.t17 VDD_VCO.t189 VDD_VCO.t113 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X48 a_70615_6448# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t112 VSS.t111 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X49 a_60304_24408# PFD_layout_0.DFF__1.CLK VSS.t230 VSS.t229 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X50 a_58943_16333# a_60634_14631.t12 VDD_VCO.t64 VDD_VCO.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X51 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VCO_op.t9 VDD.t400 VDD.t399 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X52 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t213 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X53 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_70188_5529# VSS.t528 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X54 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_74184_7541# VSS.t130 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X55 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT LP_ext.t9 VDD.t357 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X56 PFD_layout_0.DFF__0.nand2_2.IN2 PFD_layout_0.DFF__0.inv_0.OUT VDD.t658 VDD.t657 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X57 LF_mag_0.res_48k_mag_0.B VSS.t430 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X58 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t221 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X59 pu a_63452_24694# VDD.t20 VDD.t19 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X60 VDD_VCO VCO_mag_0.Delay_Cell_mag_0.OUTB.t16 VCO_mag_0.Delay_Cell_mag_0.OUT VDD_VCO.t40 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X61 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t338 VDD.t337 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X62 a_70752_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t369 VSS.t368 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X63 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.t2 VDD.t652 VDD.t651 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X64 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 a_72487_4432# VSS.t445 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X65 a_64776_7545# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t88 VSS.t87 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X66 a_63591_22645# PFD_layout_0.buffer_loading_mag_1.IN VSS.t207 VSS.t206 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X67 LF_mag_0.res_48k_mag_0.B VSS.t429 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X68 a_73051_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t325 VSS.t233 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X69 a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT a2x1mux_mag_0.Transmission_gate_mag_0.CLK VSS.t514 VSS.t513 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X70 a_65386_16333# VCO_mag_0.Delay_Cell_mag_0.OUTB.t10 VCO_mag_0.Delay_Cell_mag_0.OUTB.t11 VDD_VCO.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X71 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t606 VSS.t605 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X72 PFD_layout_0.DFF__0.inv_0.OUT PFD_layout_0.DFF__0.nand2_3.OUT VSS.t154 VSS.t153 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X73 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_72152_3335# VSS.t443 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X74 a_63276_4432# VDD.t689 VSS.t479 VSS.t478 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X75 a_73056_7541# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t215 VSS.t214 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X76 VCO_mag_0.Delay_Cell_mag_0.IN VCO_mag_0.Delay_Cell_mag_2.OUTB.t17 VSS.t188 VSS.t187 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X77 VSS EN.t1 a_65581_14091# VSS.t583 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X78 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_65128_4432# VSS.t251 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X79 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.INB a_65581_14091# VSS.t583 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X80 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t39 VDD.t38 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X81 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_71316_5529# VSS.t653 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X82 a_64212_7545# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t668 VSS.t667 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X83 PFD_layout_0.DFF__0.nand2_1.IN1 PFD_layout_0.buffer_mag_0.OUT a_60305_23482# VSS.t266 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X84 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_2.OUT.t18 VDD_VCO.t190 VDD_VCO.t109 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X85 LF_mag_0.res_48k_mag_0.B VSS.t428 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X86 VDD a_63452_24694# pu.t6 VDD.t16 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X87 PFD_layout_0.DFF__1.nand2_2.IN1 VDD.t491 VDD.t493 VDD.t492 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X88 a_67806_9704# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_67646_9704# VSS.t332 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X89 a_74184_7541# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t346 VSS.t345 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X90 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_1.INB.t6 a_65386_20072# VDD_VCO.t131 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X91 LF_mag_0.res_48k_mag_0.B VSS.t427 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X92 a_70188_5529# RST_DIV.t2 a_70028_5529# VSS.t594 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X93 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t334 VDD.t333 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X94 LF_mag_0.res_48k_mag_0.B VSS.t426 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X95 LF_mag_0.res_48k_mag_0.B VSS.t425 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X96 a_72487_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_72327_4432# VSS.t445 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X97 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t391 VDD.t390 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X98 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 VDD.t235 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X99 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD.t300 VDD.t299 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X100 LF_mag_0.res_48k_mag_0.B VSS.t424 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X101 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__1.nand2_5.OUT a_59418_24365# VSS.t158 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X102 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t232 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X103 VDD VCO_op.t10 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t401 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X104 VCO_mag_0.VCONT CP_mag_0.inv_0.OUT a_67611_25266# VDD.t153 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.56u
X105 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.OUTB.t18 VCO_mag_0.Delay_Cell_mag_0.IN VDD_VCO.t114 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X106 LF_mag_0.res_48k_mag_0.B VSS.t423 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X107 LF_mag_0.VCNTL a2x1mux_mag_0.SEL VCO_mag_0.VCONT.t20 VSS.t104 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X108 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t592 VDD.t591 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X109 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t358 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_73051_4432# VSS.t233 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X111 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD.t296 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X112 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 a_69333_7501# VSS.t577 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X113 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_61552_8823# VSS.t246 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X114 VDD_VCO VCO_mag_0.Delay_Cell_mag_1.INB.t18 VCO_mag_0.Delay_Cell_mag_1.IN VDD_VCO.t125 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X115 a_73615_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t319 VSS.t233 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X116 a_63452_24694# PFD_layout_0.nand2_0.IN1 VSS.t75 VSS.t74 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X117 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT LF_mag_0.VCNTL.t9 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X118 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t267 VDD.t266 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X119 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__1.nand2_1.IN1 VDD.t420 VDD.t419 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X120 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t502 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X121 VCO_op_bar VCO_mag_0.GF_INV16_1.IN VDD_VCO.t153 VDD_VCO.t152 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X122 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VSS.t331 VSS.t330 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X123 a_58357_44128# a_58117_42026# VDD.t253 ppolyf_u r_width=0.8u r_length=10u
X124 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.IN.t16 VCO_mag_0.Delay_Cell_mag_2.INB VDD_VCO.t24 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X125 a_65386_20072# VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.IN VDD_VCO.t140 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X126 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.DFF__1.nand2_2.OUT VDD.t45 VDD.t44 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X127 VDD_VCO a_67077_14631.t12 a_65386_16333# VDD_VCO.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X128 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t218 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X129 pu a_63452_24694# VSS.t15 VSS.t14 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X130 a_58943_20071# VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.INB VDD_VCO.t32 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X131 VSS VCO_mag_0.GF_INV1_1.OUT VCO_mag_0.GF_INV16_1.IN VSS.t289 nfet_03v3 ad=0.308p pd=2.28u as=0.182p ps=1.22u w=0.7u l=0.35u
X132 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t510 VDD.t509 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X133 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__1.nand2_3.OUT a_61533_24598# VSS.t541 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X134 a_66937_6402# RST_DIV.t3 a_66777_6402# VSS.t595 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X135 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t572 VDD.t571 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X136 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD.t506 VDD.t505 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X137 pd a_63591_22645# VSS.t228 VSS.t227 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X138 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.IN.t3 VDD_VCO.t29 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X139 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t387 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X140 LF_mag_0.res_48k_mag_0.B VSS.t422 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X141 VCO_mag_0.GF_INV16_1.IN VCO_mag_0.GF_INV1_1.OUT VSS.t288 VSS.t287 nfet_03v3 ad=0.182p pd=1.22u as=0.308p ps=2.28u w=0.7u l=0.35u
X142 LF_mag_0.VCNTL a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT VCO_mag_0.VCONT.t9 VDD.t2 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X143 a_66053_6402# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.t3 VSS.t176 VSS.t175 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X144 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t217 VDD.t216 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X145 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VCO_op.t11 VDD.t405 VDD.t404 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X146 a_58943_20071# VCO_mag_0.Delay_Cell_mag_2.IN.t14 VCO_mag_0.Delay_Cell_mag_2.IN.t15 VDD_VCO.t25 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X147 a_70028_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t534 VSS.t533 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X148 VDD RST_DIV.t4 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t604 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X149 LF_mag_0.res_48k_mag_0.B a_58597_42026# VDD.t645 ppolyf_u r_width=0.8u r_length=10u
X150 VDD IPD_.t4 a_67611_25266# VDD.t98 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.56u
X151 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t425 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X152 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t616 VDD.t615 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X153 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t191 VDD.t190 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X154 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_0.OUTB.t17 a_65581_17830# VSS.t36 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X155 VSS a_63452_24694# pu.t2 VSS.t11 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X156 LF_mag_0.res_48k_mag_0.B VSS.t421 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X157 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT LF_mag_0.VCNTL.t7 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X158 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD.t422 VDD.t421 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X159 a_57397_44128# a_57157_42026# VDD.t650 ppolyf_u r_width=0.8u r_length=10u
X160 a_66777_6402# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t49 VSS.t48 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X161 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.OUTB.t18 VDD_VCO.t87 VDD_VCO.t86 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X162 VDD PFD_layout_0.nand2_0.IN1 PFD_layout_0.DFF__1.QB VDD.t58 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X163 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.IN.t17 a_59138_14091# VSS.t635 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X164 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD.t310 VDD.t309 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X165 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VDD.t668 VDD.t667 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X166 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VCO_op.t12 VDD.t407 VDD.t406 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X167 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.CLK LP_ext.t18 VSS.t512 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X168 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t415 VDD.t414 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X169 VCO_mag_0.GF_INV1_1.OUT VCO_mag_0.Delay_Cell_mag_1.IN VDD_VCO.t139 VDD_VCO.t138 pfet_03v3 ad=0.165p pd=1.64u as=0.165p ps=1.64u w=0.35u l=0.35u
X170 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t642 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_66937_6402# VSS.t317 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X172 a_60301_26043# PFD_layout_0.DFF__1.nand2_2.OUT VSS.t55 VSS.t54 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X173 VDD_VCO a_67077_18370.t13 a_65386_20072# VDD_VCO.t46 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X174 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t120 VDD.t119 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X175 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VSS.t47 VSS.t46 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X176 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_70598_4432# VSS.t237 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X177 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD.t114 VDD.t113 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X178 LF_mag_0.res_48k_mag_0.B VSS.t420 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X179 LF_mag_0.res_48k_mag_0.B VSS.t419 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X180 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD.t330 VDD.t329 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X181 a_66213_6402# VCO_op.t13 a_66053_6402# VSS.t357 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X182 LF_mag_0.VCNTL a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT VCO_mag_0.VCONT.t8 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X183 VSS PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.OUT VSS.t43 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X184 VDD PFD_layout_0.DFF__0.QB PFD_layout_0.buffer_loading_mag_1.IN VDD.t451 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X185 a_57877_44128# a_57637_42026# VDD.t566 ppolyf_u r_width=0.8u r_length=10u
X186 VDD VCO_op.t14 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t408 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X187 VDD_VCO VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.OUTB.t3 VDD_VCO.t95 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X188 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT VCO_mag_0.VCONT.t28 VDD.t356 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X189 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_2.OUTB.t10 a_58943_16333# VDD_VCO.t113 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X190 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD.t636 VDD.t635 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X191 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t326 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X192 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_66219_7499# VSS.t294 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X193 LF_mag_0.res_48k_mag_0.B VSS.t418 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X194 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_70034_4432# VSS.t367 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X195 a_69304_5529# VDD.t690 VSS.t477 VSS.t476 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X196 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t103 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X197 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t620 VDD.t619 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X198 a_61544_9654# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD.t372 VDD.t371 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X199 a_65386_16333# VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.OUT VDD_VCO.t40 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X200 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t499 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X201 a_63591_22645# PFD_layout_0.buffer_loading_mag_1.IN VDD.t186 VDD.t185 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X202 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t66 VDD.t65 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X203 a_65581_17830# VCO_mag_0.Delay_Cell_mag_0.OUTB.t19 VCO_mag_0.Delay_Cell_mag_1.INB.t14 VSS.t164 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X204 a_71248_9766# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT VDD.t550 VDD.t549 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X205 LF_mag_0.res_48k_mag_0.B VSS.t417 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X206 a_61538_21913# PFD_layout_0.DFF__0.inv_0.OUT VSS.t641 VSS.t275 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X207 VSS VCO_mag_0.VCONT.t46 a_67077_18370.t2 VSS.t350 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X208 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t491 VSS.t490 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X209 VDD VCO_op.t15 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t411 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X210 a_62430_23292# PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.QB VSS.t517 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X211 a2x1mux_mag_0.Transmission_gate_mag_0.CLK a2x1mux_mag_0.SEL VDD.t88 VDD.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X212 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.IN a_65581_14091# VSS.t59 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X213 VSS VCO_mag_0.GF_INV16_1.IN VCO_op_bar.t3 VSS.t304 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X214 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD.t595 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X215 VCO_mag_0.GF_INV1_1.OUT VCO_mag_0.Delay_Cell_mag_1.IN VSS.t261 VSS.t260 nfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.35u
X216 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT VDD.t395 VDD.t394 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X217 a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT a2x1mux_mag_0.SEL VDD.t86 VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X218 a_59138_17829# VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_2.INB VSS.t259 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X219 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t522 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X220 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.OUTB.t20 VCO_mag_0.Delay_Cell_mag_2.OUT.t3 VDD_VCO.t110 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X221 a_63802_6404# RST_DIV.t5 a_63642_6404# VSS.t596 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X222 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t622 VDD.t621 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X223 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_73210_6400# VSS.t601 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X224 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_2.OUTB.t8 a_58943_16333# VDD_VCO.t109 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X225 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t323 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X226 VDD PFD_layout_0.nand2_0.IN1 a_63452_24694# VDD.t55 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X227 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_66447_5529# VSS.t314 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X228 a_67011_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t334 VSS.t333 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X229 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.IN VSS.t344 VSS.t343 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X230 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD.t368 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X231 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT VCO_mag_0.VCONT.t27 VDD.t355 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X232 a_59138_17829# VCO_mag_0.Delay_Cell_mag_1.INB.t19 VCO_mag_0.Delay_Cell_mag_2.IN.t6 VSS.t544 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X233 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.OUT.t19 VCO_mag_0.Delay_Cell_mag_2.OUTB.t15 VDD_VCO.t106 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X234 VDD a_63591_22645# pd.t6 VDD.t203 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X235 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_68511_9745# VSS.t324 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X236 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_67171_5529# VSS.t91 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X237 VSS PFD_layout_0.buffer_mag_0.IN PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VSS.t340 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X238 VSS VCO_mag_0.VCONT.t47 a_60634_18369.t3 VSS.t573 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X239 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t312 VDD.t311 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X240 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t6 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X241 VDD_VCO VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.INB.t11 VDD_VCO.t135 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X242 a_67735_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X243 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_69470_4432# VSS.t620 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X244 a_57877_44128# a_58117_42026# VDD.t151 ppolyf_u r_width=0.8u r_length=10u
X245 a_70034_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t608 VSS.t607 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X246 VDD_VCO VCO_mag_0.GF_INV16_2.IN VCO_op.t7 VDD_VCO.t17 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.35u
X247 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t198 VDD.t197 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X248 a_59138_14091# VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.OUTB.t3 VSS.t35 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X249 a_67611_25266# IPD_.t5 VDD.t559 VDD.t558 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.56u
X250 VSS EN.t2 a_65581_17830# VSS.t352 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X251 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.IN a_65386_20072# VDD_VCO.t134 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X252 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t488 VDD.t490 VDD.t489 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X253 a_65581_14091# EN.t3 VSS.t588 VSS.t58 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X254 a_60305_23482# PFD_layout_0.DFF__0.CLK VSS.t253 VSS.t252 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X255 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT LP_ext.t6 VDD.t354 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X256 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 VSS.t272 VSS.t271 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X257 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t150 VDD.t149 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X258 pu a_63452_24694# VDD.t15 VDD.t14 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X259 PFD_layout_0.DFF__0.inv_0.OUT PFD_layout_0.DFF__0.nand2_3.OUT VDD.t139 VDD.t138 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X260 VDD_VCO a_60634_18369.t6 a_60634_18369.t7 VDD_VCO.t77 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X261 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN VDD.t626 VDD.t625 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X262 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD.t444 VDD.t443 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X263 LF_mag_0.res_48k_mag_0.B VSS.t416 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X264 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_68299_5529# VSS.t313 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X265 a_69327_6404# VCO_op.t16 a_69167_6404# VSS.t79 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X266 a_63591_22645# PFD_layout_0.buffer_loading_mag_1.IN VSS.t205 VSS.t204 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X267 a_65581_14091# VCO_mag_0.Delay_Cell_mag_0.IN VCO_mag_0.Delay_Cell_mag_0.OUT VSS.t58 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X268 LF_mag_0.res_48k_mag_0.B VSS.t415 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X269 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD.t442 VDD.t441 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X270 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t612 VDD.t611 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X271 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VCO_op.t17 VSS.t81 VSS.t80 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X272 VDD VCO_op.t18 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t67 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X273 a_67171_5529# RST_DIV.t6 a_67011_5529# VSS.t597 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X274 a_59418_24365# VDD.t691 VSS.t475 VSS.t474 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X275 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VSS.t312 VSS.t311 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X276 a_69470_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_69310_4432# VSS.t310 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X277 LF_mag_0.res_48k_mag_0.B VSS.t414 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X278 VDD PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.buffer_mag_0.IN VDD.t182 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X279 VCO_mag_0.GF_INV16_2.IN VCO_mag_0.GF_INV1_0.OUT VSS.t522 VSS.t521 nfet_03v3 ad=0.182p pd=1.22u as=0.308p ps=2.28u w=0.7u l=0.35u
X280 a_59138_14091# EN.t4 VSS.t590 VSS.t589 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X281 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD.t291 VDD.t290 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X282 a_67501_6446# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t349 VSS.t348 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X283 LF_mag_0.res_48k_mag_0.B VSS.t413 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X284 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_71179_6448# VSS.t245 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X285 VSS VCO_mag_0.VCONT.t49 a_60634_18369.t2 VSS.t542 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X286 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VDD.t568 VDD.t567 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X287 a_56917_44128# a_57157_42026# VDD.t396 ppolyf_u r_width=0.8u r_length=10u
X288 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.CLK LP_ext.t17 VSS.t511 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X289 VSS PFD_layout_0.nand2_0.IN1 a_63452_24694# VSS.t71 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X290 a_59138_14091# VCO_mag_0.Delay_Cell_mag_2.IN.t18 VCO_mag_0.Delay_Cell_mag_2.OUT.t15 VSS.t589 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X291 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 VDD.t627 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X292 LF_mag_0.res_48k_mag_0.B VSS.t412 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X293 LF_mag_0.res_48k_mag_0.B VSS.t411 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X294 CP_mag_0.inv_0.OUT pu.t8 VDD.t649 VDD.t648 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X295 a_69167_6404# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT VSS.t356 VSS.t355 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X296 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_68065_6446# VSS.t286 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X297 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t542 VDD.t541 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X298 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.OUT a_65386_16333# VDD_VCO.t86 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X299 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.IN.t19 VDD_VCO.t182 VDD_VCO.t33 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X300 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.IN a_65386_20072# VDD_VCO.t133 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X301 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT VDD.t393 VDD.t392 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X302 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t424 VDD.t423 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X303 a_61533_24598# PFD_layout_0.DFF__1.nand2_1.IN1 VSS.t362 VSS.t361 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X304 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_64718_5529# VSS.t279 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X305 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_73774_6444# VSS.t485 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X306 VCO_mag_0.Delay_Cell_mag_0.IN VCO_mag_0.Delay_Cell_mag_2.OUTB.t22 VDD_VCO.t108 VDD_VCO.t107 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X307 LF_mag_0.res_48k_mag_0.B VSS.t410 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X308 LF_mag_0.res_48k_mag_0.B VSS.t409 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X309 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.INB a_58943_20071# VDD_VCO.t28 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X310 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VSS.t503 VSS.t502 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X311 LF_mag_0.res_48k_mag_0.B VSS.t408 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X312 VSS a_63591_22645# pd.t2 VSS.t224 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X313 VDD PFD_layout_0.DFF__1.QB PFD_layout_0.nand2_0.IN1 VDD.t194 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X314 a_72152_3335# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VSS.t444 VSS.t443 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X315 LF_mag_0.res_48k_mag_0.B VSS.t407 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X316 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_63430_5529# VSS.t442 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X317 a_57397_44128# a_57637_42026# VDD.t584 ppolyf_u r_width=0.8u r_length=10u
X318 PFD_layout_0.DFF__1.nand2_2.OUT PFD_layout_0.DFF__1.nand2_2.IN2 VDD.t470 VDD.t469 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X319 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT LF_mag_0.VCNTL.t5 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X320 VDD_VCO VCO_mag_0.GF_INV16_1.IN VCO_op_bar.t5 VDD_VCO.t149 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.35u
X321 LF_mag_0.res_48k_mag_0.B VSS.t406 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X322 a_63994_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t161 VSS.t160 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X323 PFD_layout_0.DFF__0.CLK PFD_layout_0.VDIV VSS.t139 VSS.t138 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X324 a_71179_6448# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t555 VSS.t554 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X325 PFD_layout_0.DFF__0.nand2_2.OUT PFD_layout_0.DFF__0.nand2_2.IN2 VDD.t92 VDD.t91 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X326 a_65128_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t600 VSS.t599 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X327 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD.t664 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X328 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_66783_7543# VSS.t347 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X329 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.OUT VDD_VCO.t159 VDD_VCO.t94 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X330 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t546 VDD.t545 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X331 a_71316_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t321 VSS.t320 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X332 pu a_63452_24694# VSS.t10 VSS.t9 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X333 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VDD.t37 VDD.t36 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X334 VSS CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 PFD_layout_0.VDIV VSS.t638 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X335 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_64154_5529# VSS.t256 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X336 a_65386_16333# VCO_mag_0.Delay_Cell_mag_0.OUTB.t8 VCO_mag_0.Delay_Cell_mag_0.OUTB.t9 VDD_VCO.t95 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X337 VSS PFD_layout_0.buffer_loading_mag_1.IN a_65208_24138# VSS.t201 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X338 PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.QB a_62434_21795# VSS.t446 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X339 a_67646_9704# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS.t323 VSS.t322 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X340 a_68065_6446# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t235 VSS.t234 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X341 PFD_layout_0.DFF__1.inv_0.OUT PFD_layout_0.DFF__1.nand2_3.OUT VDD.t557 VDD.t556 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X342 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t661 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X343 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_66453_4432# VSS.t281 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X344 VDD RST_DIV.t7 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t607 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X345 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t109 VDD.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X346 VDD PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.OUT VDD.t33 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X347 VSS VCO_mag_0.GF_INV16_2.IN VCO_op.t3 VSS.t29 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X348 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t296 VSS.t295 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X349 LF_mag_0.res_48k_mag_0.B VSS.t405 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X350 a_72327_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS.t551 VSS.t445 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X351 a_73774_6444# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t212 VSS.t211 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X352 PFD_layout_0.DFF__1.QB PFD_layout_0.DFF__1.nand2_5.OUT VDD.t146 VDD.t145 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X353 VCO_mag_0.Delay_Cell_mag_0.INB VCO_mag_0.Delay_Cell_mag_2.OUT.t20 VDD_VCO.t194 VDD_VCO.t193 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X354 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD.t367 VDD.t366 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X355 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_1.IN VDD_VCO.t132 VDD_VCO.t131 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X356 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 a_74179_4432# VSS.t233 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X357 VCO_op VCO_mag_0.GF_INV16_2.IN VSS.t28 VSS.t27 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X358 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD.t365 VDD.t364 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X359 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t552 VDD.t551 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X360 LF_mag_0.res_48k_mag_0.B VSS.t404 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X361 VCO_op VCO_mag_0.GF_INV16_2.IN VSS.t26 VSS.t25 nfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X362 VSS PFD_layout_0.nand2_0.IN1 a_62429_24598# VSS.t68 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X363 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD.t231 VDD.t230 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X364 a_69333_7501# VCO_op.t19 a_69173_7501# VSS.t82 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X365 a_61552_8823# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VSS.t329 VSS.t246 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X366 LF_mag_0.res_48k_mag_0.B VSS.t403 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X367 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 VDD.t130 VDD.t129 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X368 a_66783_7543# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t359 VSS.t358 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X369 LF_mag_0.VCNTL.t20 a_56677_42026# VDD.t656 ppolyf_u r_width=0.8u r_length=10u
X370 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_70461_7545# VSS.t624 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X371 PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.nand2_2.IN2 VDD.t90 VDD.t89 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X372 a_58943_16333# VCO_mag_0.Delay_Cell_mag_2.OUT.t12 VCO_mag_0.Delay_Cell_mag_2.OUT.t13 VDD_VCO.t110 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X373 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VSS.t441 VSS.t440 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X374 a_71025_7545# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t136 VSS.t135 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X375 VSS VCO_mag_0.GF_INV1_0.OUT VCO_mag_0.GF_INV16_2.IN VSS.t518 nfet_03v3 ad=0.308p pd=2.28u as=0.182p ps=1.22u w=0.7u l=0.35u
X376 VDD_VCO a_60634_14631.t6 a_60634_14631.t7 VDD_VCO.t70 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X377 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t540 VDD.t539 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X378 a_59584_26036# PFD_layout_0.DFF__1.nand2_2.IN2 VSS.t463 VSS.t462 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X379 VCO_mag_0.VCONT a2x1mux_mag_0.SEL LF_mag_0.VCNTL.t17 VSS.t103 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X380 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT LP_ext.t5 VDD.t353 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X381 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VSS.t285 VSS.t284 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X382 VDD_VCO VCO_mag_0.Delay_Cell_mag_1.INB.t20 VCO_mag_0.Delay_Cell_mag_1.IN VDD_VCO.t140 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X383 VDD VCO_op.t20 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t70 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X384 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J VDD.t583 VDD.t582 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X385 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.OUT VDD_VCO.t158 VDD_VCO.t93 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X386 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t163 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X387 a_74179_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t532 VSS.t233 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X388 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.IN.t20 VCO_mag_0.Delay_Cell_mag_2.INB VDD_VCO.t32 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X389 a_58943_16333# VCO_mag_0.Delay_Cell_mag_2.OUTB.t6 VCO_mag_0.Delay_Cell_mag_2.OUTB.t7 VDD_VCO.t106 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X390 VDD PFD_layout_0.buffer_loading_mag_1.IN a_63591_22645# VDD.t179 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X391 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VDD.t632 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X392 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD.t361 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X393 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t155 VDD.t154 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X394 VSS EN.t5 a_59138_14091# VSS.t34 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X395 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD.t295 VDD.t294 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X396 VDD PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.nand2_2.IN1 VDD.t531 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X397 VDD_VCO a_67077_14631.t14 a_65386_16333# VDD_VCO.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X398 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_70216_3335# VSS.t308 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X399 LF_mag_0.res_48k_mag_0.B VSS.t402 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X400 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_73205_5529# VSS.t318 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X401 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VDD.t521 VDD.t520 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X402 a_69173_7501# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT VSS.t354 VSS.t353 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X403 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.IN VDD.t384 VDD.t383 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X404 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t548 VDD.t547 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X405 VDD PFD_layout_0.DFF__1.nand2_1.IN1 PFD_layout_0.DFF__1.nand2_2.IN2 VDD.t416 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X406 LF_mag_0.VCNTL a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT VCO_mag_0.VCONT.t7 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X407 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS.t449 VSS.t448 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X408 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT a_61106_7416# VDD.t26 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X409 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t43 VDD.t42 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X410 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_1.INB.t4 a_65386_20072# VDD_VCO.t129 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X411 VDD RST_DIV.t8 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t672 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X412 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_69897_7545# VSS.t110 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X413 VSS CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t578 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X414 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t159 VDD.t158 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X415 PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.DFF__0.nand2_5.OUT a_59419_23525# VSS.t516 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X416 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_2.INB a_59138_14091# VSS.t34 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X417 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_60307_8532# VSS.t283 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X418 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS.t483 VSS.t482 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X419 LF_mag_0.res_48k_mag_0.B VSS.t401 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X420 a_70461_7545# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t78 VSS.t77 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X421 LF_mag_0.res_48k_mag_0.B VSS.t400 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X422 VDD PFD_layout_0.buffer_mag_0.IN PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VDD.t380 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X423 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.IN.t2 VDD_VCO.t25 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X424 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT VCO_mag_0.VCONT.t26 VDD.t352 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X425 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t588 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X426 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VCO_op.t21 VSS.t84 VSS.t83 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X427 VDD PFD_layout_0.DFF__0.nand2_3.OUT PFD_layout_0.DFF__0.nand2_5.OUT VDD.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X428 a_58943_20071# a_60634_18369.t14 VDD_VCO.t183 VDD_VCO.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X429 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t157 VDD.t156 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X430 a_63452_24694# PFD_layout_0.nand2_0.IN1 VDD.t54 VDD.t53 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X431 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 a_71025_7545# VSS.t598 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X432 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_1.IN a_59138_17829# VSS.t258 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X433 VDD VCO_op.t22 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X434 VDD_VCO a_60634_14631.t15 a_58943_16333# VDD_VCO.t61 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X435 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.OUTB.t23 VDD_VCO.t105 VDD_VCO.t104 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X436 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t538 VDD.t537 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X437 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VDD.t345 VDD.t344 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X438 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_60140_9217# VSS.t501 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X439 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t508 VDD.t507 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X440 VDD VCO_op.t23 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t76 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X441 VCO_op_bar VCO_mag_0.GF_INV16_1.IN VSS.t303 VSS.t302 nfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X442 a_70598_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t527 VSS.t526 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X443 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VDD.t32 VDD.t31 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X444 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_72486_6400# VSS.t328 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X445 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t517 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X446 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.CLK VCO_mag_0.VCONT.t37 VSS.t510 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X447 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.IN.t21 a_59138_14091# VSS.t191 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X448 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_74380_2641# VDD.t270 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X449 a_73050_6400# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t538 VSS.t537 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X450 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.OUT.t21 VCO_mag_0.Delay_Cell_mag_0.INB VDD_VCO.t195 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X451 VDD PFD_layout_0.nand2_0.IN1 a_63452_24694# VDD.t50 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X452 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t128 VSS.t127 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X453 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_71162_4432# VSS.t619 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X454 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t485 VDD.t487 VDD.t486 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X455 a_66219_7499# VCO_op.t24 a_66059_7499# VSS.t85 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X456 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT VCO_mag_0.VCONT.t25 VDD.t351 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X457 a_65581_17830# EN.t6 VSS.t593 VSS.t164 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X458 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.t4 VDD.t170 VDD.t169 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X459 VDD IPD_.t2 IPD_.t3 VDD.t95 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.56u
X460 a_65386_20072# VCO_mag_0.Delay_Cell_mag_1.INB.t2 VCO_mag_0.Delay_Cell_mag_1.INB.t3 VDD_VCO.t126 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X461 a_69897_7545# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t218 VSS.t217 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X462 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t187 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X463 LF_mag_0.res_48k_mag_0.B VSS.t399 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X464 VSS PFD_layout_0.buffer_loading_mag_1.IN a_63591_22645# VSS.t198 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X465 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD.t306 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X466 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t614 VDD.t613 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X467 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t534 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X468 LF_mag_0.res_48k_mag_0.B VSS.t398 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X469 PFD_layout_0.DFF__1.CLK Vref.t0 VDD.t302 VDD.t301 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X470 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 VSS.t142 VSS.t141 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X471 a_62918_6404# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J VSS.t568 VSS.t559 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X472 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT VDD.t118 VDD.t117 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X473 VDD_VCO a_60634_14631.t16 a_58943_16333# VDD_VCO.t67 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X474 a_72486_6400# VCO_op.t25 a_72326_6400# VSS.t86 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X475 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VCO_op.t26 VDD.t576 VDD.t575 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X476 a_74380_2641# CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 a_74220_2641# VDD.t655 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X477 PFD_layout_0.buffer_mag_0.IN PFD_layout_0.nand2_0.IN1 VDD.t49 VDD.t48 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X478 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.OUTB.t20 VDD_VCO.t89 VDD_VCO.t88 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X479 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J VDD.t581 VDD.t580 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X480 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_72492_7497# VSS.t129 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X481 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD.t110 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X482 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_63078_6404# VSS.t500 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X483 a_65581_17830# VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_1.IN VSS.t119 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X484 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD.t229 VDD.t228 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X485 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VDD.t47 VDD.t46 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X486 a_71162_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t489 VSS.t488 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X487 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t639 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X488 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.OUTB.t6 a_65386_16333# VDD_VCO.t94 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X489 a_63452_24694# PFD_layout_0.nand2_0.IN1 VSS.t67 VSS.t66 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X490 a_73210_6400# RST_DIV.t9 a_73050_6400# VSS.t654 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X491 a_63642_6404# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t53 VSS.t52 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X492 a_59585_21854# PFD_layout_0.DFF__0.nand2_2.IN2 VSS.t109 VSS.t108 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X493 a_63016_9651# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t460 VDD.t459 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X494 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD.t458 VDD.t457 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X495 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t482 VDD.t484 VDD.t483 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X496 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD.t322 VDD.t321 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X497 a_66059_7499# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.t5 VSS.t190 VSS.t189 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X498 a_66447_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_66287_5529# VSS.t439 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X499 LF_mag_0.res_48k_mag_0.B VSS.t397 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X500 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t374 VDD.t373 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X501 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t193 VDD.t192 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X502 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.IN VDD.t379 VDD.t378 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X503 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t613 VSS.t612 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X504 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VSS.t42 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X505 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.OUTB.t24 VCO_mag_0.Delay_Cell_mag_2.OUT.t1 VDD_VCO.t101 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X506 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t84 VDD.t83 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X507 a_68511_9745# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t244 VSS.t243 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X508 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN VDD.t544 VDD.t543 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X509 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t25 VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X510 pd a_63591_22645# VSS.t222 VSS.t221 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X511 a_72492_7497# VCO_op.t27 a_72332_7497# VSS.t558 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X512 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t386 VDD.t385 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X513 PFD_layout_0.nand2_0.IN1 PFD_layout_0.DFF__1.nand2_2.IN2 VDD.t468 VDD.t467 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X514 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.CLK LP_ext.t15 VSS.t509 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X515 LF_mag_0.res_48k_mag_0.B VSS.t396 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X516 VSS PFD_layout_0.nand2_0.IN1 a_63452_24694# VSS.t63 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X517 VDD PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.nand2_3.OUT VDD.t263 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X518 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS.t366 VSS.t365 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X519 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t160 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X520 LF_mag_0.res_48k_mag_0.B VSS.t395 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X521 VSS IPD+.t2 IPD+.t3 VSS.t457 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X522 a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT a2x1mux_mag_0.Transmission_gate_mag_0.CLK VDD.t528 VDD.t527 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X523 LF_mag_0.res_48k_mag_0.B VSS.t394 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X524 a_63078_6404# VCO_op.t28 a_62918_6404# VSS.t559 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X525 a_59138_17829# VCO_mag_0.Delay_Cell_mag_1.INB.t22 VCO_mag_0.Delay_Cell_mag_2.IN.t5 VSS.t121 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X526 VCO_mag_0.Delay_Cell_mag_0.INB VCO_mag_0.Delay_Cell_mag_2.OUT.t22 VSS.t665 VSS.t664 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X527 pd a_63591_22645# VDD.t202 VDD.t201 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X528 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.OUT.t23 VCO_mag_0.Delay_Cell_mag_2.OUTB.t12 VDD_VCO.t100 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X529 LF_mag_0.VCNTL a2x1mux_mag_0.SEL VCO_mag_0.VCONT.t19 VSS.t102 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X530 VDD VCO_op.t29 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t577 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X531 a_66287_5529# VDD.t692 VSS.t473 VSS.t472 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X532 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t647 VDD.t646 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X533 VCO_mag_0.GF_INV1_0.OUT VCO_mag_0.Delay_Cell_mag_1.INB.t23 VSS.t546 VSS.t545 nfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.35u
X534 a_58943_16333# a_60634_14631.t17 VDD_VCO.t71 VDD_VCO.t70 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X535 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN VDD.t574 VDD.t573 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X536 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD.t318 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X537 a_65208_24138# PFD_layout_0.nand2_0.IN1 PFD_layout_0.buffer_mag_0.IN VSS.t62 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X538 a_62434_21795# PFD_layout_0.DFF__0.nand2_2.IN2 VSS.t107 VSS.t106 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X539 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.INB.t24 VDD_VCO.t171 VDD_VCO.t134 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X540 VCO_op_bar VCO_mag_0.GF_INV16_1.IN VSS.t301 VSS.t300 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X541 a_68299_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t493 VSS.t492 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X542 VDD_VCO VCO_mag_0.Delay_Cell_mag_0.OUTB.t22 VCO_mag_0.Delay_Cell_mag_0.OUT VDD_VCO.t90 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X543 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 a_63016_9651# VDD.t610 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X544 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS.t487 VSS.t486 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X545 a_56917_44128# a_56677_42026# VDD.t168 ppolyf_u r_width=0.8u r_length=10u
X546 VSS a_63591_22645# pd.t0 VSS.t219 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X547 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.OUTB.t4 a_65386_16333# VDD_VCO.t93 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X548 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VDD.t167 VDD.t166 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X549 VDD RST_DIV.t10 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t675 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X550 VSS CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t19 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X551 LF_mag_0.VCNTL.t21 VSS.t137 cap_mim_2f0_m4m5_noshield c_width=42.5u c_length=42.5u
X552 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X553 a_65581_17830# a_65581_17830# a_65581_17830# VSS.t123 nfet_03v3 ad=0.26p pd=1.52u as=4p ps=24u w=1u l=0.56u
X554 LF_mag_0.res_48k_mag_0.B VSS.t393 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X555 VDD_VCO VCO_mag_0.Delay_Cell_mag_2.OUT.t24 VCO_mag_0.Delay_Cell_mag_0.INB VDD_VCO.t175 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X556 a_69310_4432# VDD.t693 VSS.t471 VSS.t470 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X557 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t438 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X558 a_65581_14091# VCO_mag_0.Delay_Cell_mag_0.INB VCO_mag_0.Delay_Cell_mag_0.OUTB.t13 VSS.t618 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X559 a_62429_24598# PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__1.QB VSS.t157 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X560 VDD PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__1.nand2_1.IN1 VDD.t260 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X561 a_59138_17829# VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_2.INB VSS.t193 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X562 VCO_mag_0.Delay_Cell_mag_0.IN VCO_mag_0.Delay_Cell_mag_2.OUTB.t25 VSS.t186 VSS.t185 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X563 LF_mag_0.res_48k_mag_0.B VSS.t392 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X564 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.IN VSS.t339 VSS.t338 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X565 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_2.IN.t12 a_58943_20071# VDD_VCO.t22 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X566 a_62924_7501# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J VSS.t567 VSS.t566 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X567 LF_mag_0.VCNTL a2x1mux_mag_0.SEL VCO_mag_0.VCONT.t18 VSS.t101 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X568 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t21 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X569 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.OUT.t10 a_58943_16333# VDD_VCO.t104 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X570 a_65581_17830# a_65581_17830# a_65581_17830# VSS.t159 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.56u
X571 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_63084_7501# VSS.t447 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X572 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t284 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X573 LF_mag_0.res_48k_mag_0.B VSS.t391 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X574 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t82 VDD.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X575 a_64718_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t453 VSS.t452 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X576 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_60147_7030# VSS.t499 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X577 a_67017_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t626 VSS.t625 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X578 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD.t437 VDD.t436 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X579 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.INB.t25 VDD_VCO.t172 VDD_VCO.t133 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X580 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VDD.t631 VDD.t630 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X581 a_63430_5529# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_63270_5529# VSS.t140 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X582 a_59138_14091# a_59138_14091# a_59138_14091# VSS.t531 nfet_03v3 ad=0.44p pd=2.88u as=4p ps=24u w=1u l=0.56u
X583 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_71408_9766# VDD.t516 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X584 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t148 VDD.t147 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X585 PFD_layout_0.DFF__0.nand2_2.IN1 VDD.t479 VDD.t481 VDD.t480 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X586 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.inv_0.OUT VDD.t10 VDD.t9 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X587 VSS PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.OUT VSS.t38 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X588 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD.t638 VDD.t637 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X589 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD.t287 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X590 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_65282_5529# VSS.t438 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X591 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.IN.t23 VDD_VCO.t122 VDD_VCO.t28 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X592 LF_mag_0.res_48k_mag_0.B VSS.t390 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X593 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_64366_6448# VSS.t174 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X594 PFD_layout_0.nand2_0.IN1 PFD_layout_0.DFF__1.QB a_62433_26095# VSS.t216 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X595 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_67581_4432# VSS.t3 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X596 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t340 VDD.t339 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X597 a_59419_23525# VDD.t694 VSS.t469 VSS.t468 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X598 a_65386_20072# a_67077_18370.t15 VDD_VCO.t55 VDD_VCO.t43 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X599 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t249 VDD.t248 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X600 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_74338_6444# VSS.t327 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X601 a_64930_6448# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t168 VSS.t167 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X602 VCO_mag_0.VCONT a2x1mux_mag_0.SEL LF_mag_0.VCNTL.t14 VSS.t100 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X603 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_2.IN.t10 a_58943_20071# VDD_VCO.t20 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X604 VSS VCO_mag_0.VCONT.t52 a_67077_14631.t9 VSS.t570 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X605 a_64154_5529# RST_DIV.t11 a_63994_5529# VSS.t655 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X606 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT LP_ext.t2 VDD.t350 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X607 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_73769_5529# VSS.t543 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X608 LF_mag_0.res_48k_mag_0.B VSS.t389 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X609 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD.t317 VDD.t316 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X610 a_66453_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_66293_4432# VSS.t437 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X611 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.nand2_1.IN1 VDD.t278 VDD.t277 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X612 VSS VCO_mag_0.Delay_Cell_mag_2.OUT.t26 VCO_mag_0.Delay_Cell_mag_0.INB VSS.t627 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X613 a_65581_14091# a_65581_14091# a_65581_14091# VSS.t570 nfet_03v3 ad=0.26p pd=1.52u as=4p ps=24u w=1u l=0.56u
X614 a_63084_7501# VCO_op.t30 a_62924_7501# VSS.t560 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X615 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_72481_5529# VSS.t270 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X616 a_73045_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t615 VSS.t614 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X617 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN VSS.t557 VSS.t556 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X618 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD.t240 VDD.t239 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X619 a_63270_5529# VDD.t695 VSS.t467 VSS.t466 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X620 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_67347_7543# VSS.t571 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X621 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t107 VDD.t106 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X622 IPD+ IPD+.t0 VSS.t149 VSS.t148 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X623 a_67911_7543# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t170 VSS.t169 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X624 VSS CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN VSS.t454 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X625 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t313 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X626 VSS VCO_mag_0.VCONT.t53 a_60634_14631.t2 VSS.t530 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X627 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t576 VSS.t575 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X628 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_67017_4432# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X629 a_65282_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t637 VSS.t636 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X630 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.nand2_1.IN1 a_61537_25977# VSS.t360 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X631 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.OUT a_65386_16333# VDD_VCO.t88 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X632 a_64366_6448# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t525 VSS.t524 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X633 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_0.OUTB.t24 a_65581_17830# VSS.t165 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X634 a_67581_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t90 VSS.t89 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X635 a_59138_14091# a_59138_14091# a_59138_14091# VSS.t530 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.56u
X636 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t281 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X637 a_73769_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t232 VSS.t231 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X638 LF_mag_0.res_48k_mag_0.B VSS.t388 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X639 a_66293_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VSS.t156 VSS.t155 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X640 a_65581_14091# a_65581_14091# a_65581_14091# VSS.t569 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.56u
X641 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_64930_6448# VSS.t498 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X642 a_72481_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_72321_5529# VSS.t436 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X643 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_68145_4432# VSS.t280 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X644 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT VDD.t116 VDD.t115 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X645 a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT a2x1mux_mag_0.SEL VSS.t99 VSS.t98 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X646 a_65386_20072# a_67077_18370.t16 VDD_VCO.t56 VDD_VCO.t50 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X647 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_74333_5529# VSS.t269 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X648 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t268 VSS.t267 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X649 VSS VCO_mag_0.Delay_Cell_mag_2.OUTB.t26 VCO_mag_0.Delay_Cell_mag_0.IN VSS.t182 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X650 VSS PFD_layout_0.buffer_mag_0.IN PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VSS.t335 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X651 a_58943_16333# VCO_mag_0.Delay_Cell_mag_2.OUT.t8 VCO_mag_0.Delay_Cell_mag_2.OUT.t9 VDD_VCO.t101 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X652 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD.t435 VDD.t434 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X653 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t472 VDD.t471 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X654 VDD PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.QB VDD.t176 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X655 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN VDD.t358 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X656 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VDD.t660 VDD.t659 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X657 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t336 VDD.t335 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X658 a2x1mux_mag_0.Transmission_gate_mag_0.CLK a2x1mux_mag_0.SEL VSS.t97 VSS.t96 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X659 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.CLK VCO_mag_0.VCONT.t36 VSS.t508 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X660 a_70216_3335# CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VSS.t309 VSS.t308 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X661 a_73205_5529# RST_DIV.t12 a_73045_5529# VSS.t656 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X662 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN VSS.t617 VSS.t616 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X663 VCO_mag_0.VCONT pd.t8 a_67618_24851# VSS.t238 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X664 a_65581_17830# VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_1.IN VSS.t351 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X665 a_61106_7416# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT VDD.t1 VDD.t0 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X666 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_1.INB.t26 a_59138_17829# VSS.t547 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X667 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t463 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X668 a_60307_8532# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_60147_8532# VSS.t326 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X669 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_67911_7543# VSS.t293 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X670 VDD_VCO VCO_mag_0.GF_INV1_1.OUT VCO_mag_0.GF_INV16_1.IN VDD_VCO.t143 pfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X671 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t247 VDD.t246 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X672 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_63648_7545# VSS.t523 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X673 a_58943_16333# VCO_mag_0.Delay_Cell_mag_2.OUTB.t4 VCO_mag_0.Delay_Cell_mag_2.OUTB.t5 VDD_VCO.t100 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X674 LF_mag_0.res_48k_mag_0.B VSS.t387 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X675 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_63436_4432# VSS.t250 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X676 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_1.IN VDD_VCO.t130 VDD_VCO.t129 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X677 VDD_VCO a_67077_14631.t4 a_67077_14631.t5 VDD_VCO.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X678 PFD_layout_0.DFF__0.nand2_3.OUT PFD_layout_0.buffer_mag_0.OUT a_60302_21847# VSS.t265 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X679 VSS VCO_mag_0.GF_INV16_2.IN VCO_op.t0 VSS.t22 nfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X680 VSS VCO_mag_0.VCONT.t54 a_60634_14631.t1 VSS.t33 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X681 a_64000_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t114 VSS.t113 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X682 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_73620_7541# VSS.t484 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X683 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t332 VDD.t331 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X684 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT LF_mag_0.VCNTL.t3 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X685 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN VDD.t41 VDD.t40 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X686 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_71184_3335# VSS.t308 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X687 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t172 VSS.t171 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X688 VCO_mag_0.GF_INV16_1.IN VCO_mag_0.GF_INV1_1.OUT VDD_VCO.t142 VDD_VCO.t141 pfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X689 LF_mag_0.res_48k_mag_0.B VSS.t386 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X690 LF_mag_0.res_48k_mag_0.B VSS.t385 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X691 a_65386_16333# VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.OUT VDD_VCO.t90 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X692 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_2.INB a_59138_14091# VSS.t33 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X693 a_60140_9217# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t242 VSS.t241 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X694 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_70615_6448# VSS.t623 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X695 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.nand2_3.OUT a_61534_23292# VSS.t152 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X696 VDD_VCO a_60634_18369.t4 a_60634_18369.t5 VDD_VCO.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X697 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_64564_4432# VSS.t278 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X698 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT VSS.t536 VSS.t535 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X699 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t563 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X700 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_70752_5529# VSS.t236 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X701 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.IN a_65581_14091# VSS.t57 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X702 VDD_VCO VCO_mag_0.GF_INV16_1.IN VCO_op_bar.t4 VDD_VCO.t146 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X703 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_1.IN a_59138_17829# VSS.t257 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X704 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.CLK VCO_mag_0.VCONT.t35 VSS.t507 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X705 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.OUTB.t27 VDD_VCO.t99 VDD_VCO.t98 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X706 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VCO_op.t31 VSS.t562 VSS.t561 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X707 PFD_layout_0.DFF__0.nand2_3.OUT PFD_layout_0.DFF__0.nand2_2.OUT VDD.t280 VDD.t279 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X708 VSS VCO_mag_0.Delay_Cell_mag_2.OUT.t27 VCO_mag_0.Delay_Cell_mag_0.INB VSS.t630 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X709 LF_mag_0.res_48k_mag_0.B VSS.t384 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X710 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t341 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X711 a_71184_3335# CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VSS.t652 VSS.t308 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X712 VCO_mag_0.VCONT a2x1mux_mag_0.SEL LF_mag_0.VCNTL.t13 VSS.t95 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X713 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_64212_7545# VSS.t173 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X714 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VDD.t454 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X715 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_64000_4432# VSS.t451 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X716 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VCO_op.t32 a_67806_9704# VSS.t563 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X717 a_64564_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t255 VSS.t254 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X718 VDD_VCO a_67077_14631.t2 a_67077_14631.t3 VDD_VCO.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X719 a_65581_14091# VCO_mag_0.Delay_Cell_mag_0.INB VCO_mag_0.Delay_Cell_mag_0.OUTB.t12 VSS.t117 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X720 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t515 VDD.t514 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X721 LF_mag_0.res_48k_mag_0.B VSS.t383 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X722 CP_mag_0.inv_0.OUT pu.t9 VSS.t634 VSS.t633 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X723 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t585 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X724 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.CLK LP_ext.t12 VSS.t506 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X725 VDD_VCO VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.INB.t8 VDD_VCO.t126 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X726 VDD PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__1.nand2_2.OUT VDD.t250 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X727 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT LP_ext.t1 VDD.t349 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X728 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN VSS.t51 VSS.t50 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X729 a_72326_6400# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT VSS.t134 VSS.t133 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X730 a_74220_2641# CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD.t498 VDD.t497 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X731 VDD PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.DFF__0.nand2_2.OUT VDD.t303 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X732 a_65386_20072# VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.IN VDD_VCO.t125 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X733 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD.t293 VDD.t292 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X734 pd a_63591_22645# VDD.t200 VDD.t199 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X735 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN VSS.t529 VSS.t486 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X736 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t64 VDD.t63 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X737 LF_mag_0.VCNTL a2x1mux_mag_0.SEL VCO_mag_0.VCONT.t17 VSS.t94 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X738 a_58943_20071# VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.INB VDD_VCO.t24 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X739 VCO_mag_0.GF_INV1_0.OUT VCO_mag_0.Delay_Cell_mag_1.INB.t27 VDD_VCO.t85 VDD_VCO.t84 pfet_03v3 ad=0.165p pd=1.64u as=0.165p ps=1.64u w=0.35u l=0.35u
X740 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t102 VDD.t101 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X741 PFD_layout_0.DFF__1.nand2_1.IN1 PFD_layout_0.DFF__1.CLK VDD.t210 VDD.t209 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X742 VSS VCO_mag_0.GF_INV16_1.IN VCO_op_bar.t0 VSS.t297 nfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X743 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VCO_op.t33 VSS.t565 VSS.t564 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X744 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_73615_4432# VSS.t233 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X745 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t431 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X746 VSS VCO_mag_0.Delay_Cell_mag_2.OUTB.t28 VCO_mag_0.Delay_Cell_mag_0.IN VSS.t179 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X747 VDD PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.OUT VDD.t28 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X748 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t80 VDD.t79 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X749 VDD PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.nand2_1.IN1 VDD.t257 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X750 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VSS.t435 VSS.t434 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X751 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t61 VSS.t60 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X752 LF_mag_0.res_48k_mag_0.B VSS.t382 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X753 PFD_layout_0.DFF__1.nand2_1.IN1 PFD_layout_0.buffer_mag_0.OUT a_60304_24408# VSS.t264 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X754 VCO_mag_0.VCONT a2x1mux_mag_0.SEL LF_mag_0.VCNTL.t11 VSS.t93 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X755 VCO_mag_0.Delay_Cell_mag_0.INB VCO_mag_0.Delay_Cell_mag_2.OUT.t28 VDD_VCO.t179 VDD_VCO.t178 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X756 VDD PFD_layout_0.DFF__0.nand2_1.IN1 PFD_layout_0.DFF__0.nand2_2.IN2 VDD.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X757 LF_mag_0.res_48k_mag_0.B VSS.t381 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X758 a_58943_20071# VCO_mag_0.Delay_Cell_mag_2.IN.t8 VCO_mag_0.Delay_Cell_mag_2.IN.t9 VDD_VCO.t29 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X759 LF_mag_0.res_48k_mag_0.B VSS.t380 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X760 VDD a_63452_24694# pu.t4 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X761 LF_mag_0.res_48k_mag_0.B VSS.t379 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X762 a_72332_7497# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT VSS.t132 VSS.t131 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X763 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t687 VDD.t686 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X764 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t685 VDD.t684 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X765 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t476 VDD.t478 VDD.t477 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X766 a_62433_26095# PFD_layout_0.DFF__1.nand2_2.IN2 VSS.t461 VSS.t460 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X767 a_67618_24851# pd.t9 VCO_mag_0.VCONT.t10 VSS.t37 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X768 PFD_layout_0.DFF__1.inv_0.OUT PFD_layout_0.DFF__1.nand2_3.OUT VSS.t540 VSS.t539 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X769 PFD_layout_0.DFF__0.CLK PFD_layout_0.VDIV VDD.t122 VDD.t121 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X770 PFD_layout_0.DFF__1.nand2_2.OUT PFD_layout_0.DFF__1.nand2_2.IN1 a_59584_26036# VSS.t262 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X771 LF_mag_0.VCNTL a2x1mux_mag_0.SEL VCO_mag_0.VCONT.t16 VSS.t92 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X772 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t512 VDD.t511 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X773 VDD PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__1.nand2_2.IN1 VDD.t142 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X774 VDD_VCO a_60634_18369.t15 a_58943_20071# VDD_VCO.t82 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X775 VSS VCO_mag_0.VCONT.t58 a_67077_18370.t0 VSS.t123 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X776 VDD_VCO a_67077_18370.t17 a_65386_20072# VDD_VCO.t48 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X777 VDD RST_DIV.t13 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t678 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X778 VDD_VCO a_60634_14631.t4 a_60634_14631.t5 VDD_VCO.t63 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X779 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_69464_5529# VSS.t651 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X780 LF_mag_0.res_48k_mag_0.B VSS.t378 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X781 a_59138_17829# EN.t7 VSS.t194 VSS.t193 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X782 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t178 VSS.t177 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X783 VDD_VCO VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.OUTB.t0 VDD_VCO.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X784 VCO_mag_0.Delay_Cell_mag_0.IN VCO_mag_0.Delay_Cell_mag_2.OUTB.t29 VDD_VCO.t97 VDD_VCO.t96 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X785 VDD PFD_layout_0.buffer_mag_0.IN PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VDD.t375 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X786 VDD PFD_layout_0.buffer_loading_mag_1.IN a_63591_22645# VDD.t173 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X787 a_61537_25977# PFD_layout_0.DFF__1.inv_0.OUT VSS.t5 VSS.t4 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X788 LF_mag_0.VCNTL a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT VCO_mag_0.VCONT.t6 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X789 a_65386_16333# a_67077_14631.t15 VDD_VCO.t7 VDD_VCO.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X790 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_66213_6402# VSS.t282 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X791 VDD PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.DFF__1.nand2_5.OUT VDD.t553 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X792 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_70051_6404# VSS.t76 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X793 VDD PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__1.nand2_3.OUT VDD.t254 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X794 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD.t227 VDD.t226 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X795 VDD_VCO VCO_mag_0.GF_INV16_2.IN VCO_op.t6 VDD_VCO.t14 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X796 a_65581_17830# VCO_mag_0.Delay_Cell_mag_0.OUTB.t25 VCO_mag_0.Delay_Cell_mag_1.INB.t12 VSS.t166 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X797 VSS a_63452_24694# pu.t0 VSS.t6 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X798 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t570 VDD.t569 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X799 VCO_mag_0.GF_INV16_2.IN VCO_mag_0.GF_INV1_0.OUT VDD_VCO.t163 VDD_VCO.t162 pfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X800 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t462 VDD.t461 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X801 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_2.INB VDD_VCO.t23 VDD_VCO.t22 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X802 a_60147_7030# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t240 VSS.t239 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X803 a_69464_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_69304_5529# VSS.t307 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X804 VCO_op VCO_mag_0.GF_INV16_2.IN VDD_VCO.t13 VDD_VCO.t12 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X805 LF_mag_0.res_48k_mag_0.B VSS.t377 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X806 VSS IPD+.t6 a_67618_24851# VSS.t548 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X807 VCO_op VCO_mag_0.GF_INV16_2.IN VDD_VCO.t11 VDD_VCO.t10 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.35u
X808 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT a_61544_9654# VDD.t513 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X809 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT VSS.t1 VSS.t0 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X810 VDD_VCO a_60634_18369.t16 a_58943_20071# VDD_VCO.t80 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X811 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t126 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X812 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.CLK LP_ext.t11 VSS.t505 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X813 PFD_layout_0.DFF__0.QB PFD_layout_0.DFF__0.nand2_5.OUT VDD.t530 VDD.t529 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X814 a_59138_17829# a_59138_17829# a_59138_17829# VSS.t574 nfet_03v3 ad=0.44p pd=2.88u as=4p ps=24u w=1u l=0.56u
X815 a_71408_9766# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_71248_9766# VDD.t466 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X816 LF_mag_0.res_48k_mag_0.B VSS.t376 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X817 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t132 VDD.t131 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X818 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD.t428 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X819 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.OUT.t6 a_58943_16333# VDD_VCO.t98 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X820 LF_mag_0.res_48k_mag_0.B VSS.t375 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X821 VDD RST_DIV.t14 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t681 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X822 a_74338_6444# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t465 VSS.t464 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X823 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_0.OUT a_65581_17830# VSS.t350 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X824 LF_mag_0.res_48k_mag_0.B VSS.t374 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X825 LF_mag_0.res_48k_mag_0.B VSS.t373 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X826 VDD CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t560 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X827 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t618 VDD.t617 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X828 a_60302_21847# PFD_layout_0.DFF__0.nand2_2.OUT VSS.t277 VSS.t276 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X829 a_59138_14091# VCO_mag_0.Delay_Cell_mag_2.IN.t25 VCO_mag_0.Delay_Cell_mag_2.OUT.t5 VSS.t192 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X830 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_63802_6404# VSS.t666 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X831 LF_mag_0.VCNTL a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT VCO_mag_0.VCONT.t5 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X832 VDD_VCO a_67077_18370.t4 a_67077_18370.t5 VDD_VCO.t43 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X833 LF_mag_0.res_48k_mag_0.B VSS.t372 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X834 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 VDD.t269 VDD.t268 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X835 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_2.INB VDD_VCO.t21 VDD_VCO.t20 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X836 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t624 VDD.t623 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X837 a_65386_16333# a_67077_14631.t17 VDD_VCO.t9 VDD_VCO.t8 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X838 LF_mag_0.res_48k_mag_0.B VSS.t371 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X839 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.CLK VCO_mag_0.VCONT.t34 VSS.t504 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X840 a_58357_44128# a_58597_42026# VDD.t27 ppolyf_u r_width=0.8u r_length=10u
X841 LF_mag_0.res_48k_mag_0.B VSS.t370 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X842 VDD CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t123 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X843 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t473 VDD.t475 VDD.t474 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X844 a_61534_23292# PFD_layout_0.DFF__0.nand2_1.IN1 VSS.t274 VSS.t273 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X845 LP_ext a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT VCO_mag_0.VCONT.t24 VDD.t348 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X846 a_65386_20072# VCO_mag_0.Delay_Cell_mag_1.INB.t0 VCO_mag_0.Delay_Cell_mag_1.INB.t1 VDD_VCO.t135 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X847 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t622 VSS.t621 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X848 a_67347_7543# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t316 VSS.t315 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X849 a_67611_25266# CP_mag_0.inv_0.OUT VCO_mag_0.VCONT.t21 VDD.t152 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.56u
X850 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.buffer_mag_0.OUT a_60301_26043# VSS.t263 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X851 a_59138_14091# VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.OUTB.t0 VSS.t32 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X852 a_70051_6404# RST_DIV.t15 a_69891_6404# VSS.t657 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X853 IPD_ IPD_.t0 VDD.t94 VDD.t93 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.56u
X854 VSS PFD_layout_0.buffer_loading_mag_1.IN a_63591_22645# VSS.t195 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X855 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t654 VDD.t653 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X856 a_63591_22645# PFD_layout_0.buffer_loading_mag_1.IN VDD.t172 VDD.t171 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X857 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_67735_5529# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X858 PFD_layout_0.DFF__1.CLK Vref.t1 VSS.t364 VSS.t363 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X859 a_59138_17829# a_59138_17829# a_59138_17829# VSS.t573 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.56u
X860 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t212 VDD.t211 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X861 PFD_layout_0.DFF__0.nand2_2.OUT PFD_layout_0.DFF__0.nand2_2.IN1 a_59585_21854# VSS.t292 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X862 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT LF_mag_0.VCNTL.t0 VDD.t2 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X863 a_65581_14091# VCO_mag_0.Delay_Cell_mag_0.IN VCO_mag_0.Delay_Cell_mag_0.OUT VSS.t56 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X864 a_58943_20071# a_60634_18369.t17 VDD_VCO.t188 VDD_VCO.t77 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X865 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD.t225 VDD.t224 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X866 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VDD.t141 VDD.t140 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 VCO_mag_0.Delay_Cell_mag_2.OUTB.n20 VCO_mag_0.Delay_Cell_mag_2.OUTB.t24 22.2916
R1 VCO_mag_0.Delay_Cell_mag_2.OUTB.n14 VCO_mag_0.Delay_Cell_mag_2.OUTB.t8 22.1612
R2 VCO_mag_0.Delay_Cell_mag_2.OUTB.n23 VCO_mag_0.Delay_Cell_mag_2.OUTB.t28 19.1891
R3 VCO_mag_0.Delay_Cell_mag_2.OUTB.n24 VCO_mag_0.Delay_Cell_mag_2.OUTB.t17 19.1891
R4 VCO_mag_0.Delay_Cell_mag_2.OUTB.n25 VCO_mag_0.Delay_Cell_mag_2.OUTB.t26 19.1891
R5 VCO_mag_0.Delay_Cell_mag_2.OUTB.n26 VCO_mag_0.Delay_Cell_mag_2.OUTB.t25 18.6676
R6 VCO_mag_0.Delay_Cell_mag_2.OUTB.t24 VCO_mag_0.Delay_Cell_mag_2.OUTB.n19 17.311
R7 VCO_mag_0.Delay_Cell_mag_2.OUTB.n24 VCO_mag_0.Delay_Cell_mag_2.OUTB.n23 16.9365
R8 VCO_mag_0.Delay_Cell_mag_2.OUTB.n25 VCO_mag_0.Delay_Cell_mag_2.OUTB.n24 16.9365
R9 VCO_mag_0.Delay_Cell_mag_2.OUTB.n26 VCO_mag_0.Delay_Cell_mag_2.OUTB.n25 16.6457
R10 VCO_mag_0.Delay_Cell_mag_2.OUTB.n16 VCO_mag_0.Delay_Cell_mag_2.OUTB.t4 15.1219
R11 VCO_mag_0.Delay_Cell_mag_2.OUTB.n15 VCO_mag_0.Delay_Cell_mag_2.OUTB.n14 14.0791
R12 VCO_mag_0.Delay_Cell_mag_2.OUTB.n21 VCO_mag_0.Delay_Cell_mag_2.OUTB.n20 14.0791
R13 VCO_mag_0.Delay_Cell_mag_2.OUTB.n22 VCO_mag_0.Delay_Cell_mag_2.OUTB.n21 14.0791
R14 VCO_mag_0.Delay_Cell_mag_2.OUTB.n23 VCO_mag_0.Delay_Cell_mag_2.OUTB.t18 11.6805
R15 VCO_mag_0.Delay_Cell_mag_2.OUTB.n24 VCO_mag_0.Delay_Cell_mag_2.OUTB.t22 11.6805
R16 VCO_mag_0.Delay_Cell_mag_2.OUTB.n25 VCO_mag_0.Delay_Cell_mag_2.OUTB.t16 11.6805
R17 VCO_mag_0.Delay_Cell_mag_2.OUTB.n26 VCO_mag_0.Delay_Cell_mag_2.OUTB.t29 11.4719
R18 VCO_mag_0.Delay_Cell_mag_2.OUTB.n20 VCO_mag_0.Delay_Cell_mag_2.OUTB.t27 8.213
R19 VCO_mag_0.Delay_Cell_mag_2.OUTB.n21 VCO_mag_0.Delay_Cell_mag_2.OUTB.t20 8.213
R20 VCO_mag_0.Delay_Cell_mag_2.OUTB.n22 VCO_mag_0.Delay_Cell_mag_2.OUTB.t23 8.213
R21 VCO_mag_0.Delay_Cell_mag_2.OUTB.n15 VCO_mag_0.Delay_Cell_mag_2.OUTB.t10 8.08264
R22 VCO_mag_0.Delay_Cell_mag_2.OUTB.n14 VCO_mag_0.Delay_Cell_mag_2.OUTB.t6 8.08264
R23 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_2.OUTB.n26 7.24687
R24 VCO_mag_0.Delay_Cell_mag_2.OUTB.n16 VCO_mag_0.Delay_Cell_mag_2.OUTB.n15 7.03979
R25 VCO_mag_0.Delay_Cell_mag_2.OUTB.n10 VCO_mag_0.Delay_Cell_mag_2.OUTB.n9 4.70398
R26 VCO_mag_0.Delay_Cell_mag_2.OUTB.n11 VCO_mag_0.Delay_Cell_mag_2.OUTB.n10 4.4843
R27 VCO_mag_0.Delay_Cell_mag_2.OUTB.n17 VCO_mag_0.Delay_Cell_mag_2.OUTB.n16 4.0005
R28 VCO_mag_0.Delay_Cell_mag_2.OUTB.n19 VCO_mag_0.Delay_Cell_mag_2.OUTB.n1 3.3342
R29 VCO_mag_0.Delay_Cell_mag_2.OUTB.n10 VCO_mag_0.Delay_Cell_mag_2.OUTB.n7 3.1505
R30 VCO_mag_0.Delay_Cell_mag_2.OUTB.n17 VCO_mag_0.Delay_Cell_mag_2.OUTB.n13 2.94411
R31 VCO_mag_0.Delay_Cell_mag_2.OUTB.n19 VCO_mag_0.Delay_Cell_mag_2.OUTB.n3 2.9292
R32 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_2.OUTB.n22 2.70347
R33 VCO_mag_0.Delay_Cell_mag_2.OUTB.n11 VCO_mag_0.Delay_Cell_mag_2.OUTB.n5 2.6005
R34 VCO_mag_0.Delay_Cell_mag_2.OUTB.n5 VCO_mag_0.Delay_Cell_mag_2.OUTB.t12 1.8205
R35 VCO_mag_0.Delay_Cell_mag_2.OUTB.n5 VCO_mag_0.Delay_Cell_mag_2.OUTB.n4 1.8205
R36 VCO_mag_0.Delay_Cell_mag_2.OUTB.n3 VCO_mag_0.Delay_Cell_mag_2.OUTB.t15 1.8205
R37 VCO_mag_0.Delay_Cell_mag_2.OUTB.n3 VCO_mag_0.Delay_Cell_mag_2.OUTB.n2 1.8205
R38 VCO_mag_0.Delay_Cell_mag_2.OUTB.n1 VCO_mag_0.Delay_Cell_mag_2.OUTB.t7 1.8205
R39 VCO_mag_0.Delay_Cell_mag_2.OUTB.n1 VCO_mag_0.Delay_Cell_mag_2.OUTB.n0 1.8205
R40 VCO_mag_0.Delay_Cell_mag_2.OUTB.n13 VCO_mag_0.Delay_Cell_mag_2.OUTB.t5 1.8205
R41 VCO_mag_0.Delay_Cell_mag_2.OUTB.n13 VCO_mag_0.Delay_Cell_mag_2.OUTB.n12 1.8205
R42 VCO_mag_0.Delay_Cell_mag_2.OUTB.n7 VCO_mag_0.Delay_Cell_mag_2.OUTB.t0 1.6385
R43 VCO_mag_0.Delay_Cell_mag_2.OUTB.n7 VCO_mag_0.Delay_Cell_mag_2.OUTB.n6 1.6385
R44 VCO_mag_0.Delay_Cell_mag_2.OUTB.n9 VCO_mag_0.Delay_Cell_mag_2.OUTB.t3 1.6385
R45 VCO_mag_0.Delay_Cell_mag_2.OUTB.n9 VCO_mag_0.Delay_Cell_mag_2.OUTB.n8 1.6385
R46 VCO_mag_0.Delay_Cell_mag_2.OUTB.n19 VCO_mag_0.Delay_Cell_mag_2.OUTB.n18 0.845717
R47 VCO_mag_0.Delay_Cell_mag_2.OUTB.n18 VCO_mag_0.Delay_Cell_mag_2.OUTB.n17 0.335065
R48 VCO_mag_0.Delay_Cell_mag_2.OUTB.n18 VCO_mag_0.Delay_Cell_mag_2.OUTB.n11 0.329196
R49 VDD_VCO.n375 VDD_VCO.t84 335.682
R50 VDD_VCO.n323 VDD_VCO.t138 335.682
R51 VDD_VCO.n167 VDD_VCO.t114 179.427
R52 VDD_VCO.n596 VDD_VCO.t175 179.427
R53 VDD_VCO.n178 VDD_VCO.t117 112.441
R54 VDD_VCO.n602 VDD_VCO.t195 112.441
R55 VDD_VCO.n180 VDD_VCO.t107 52.6321
R56 VDD_VCO.n600 VDD_VCO.t178 52.6321
R57 VDD_VCO.n305 VDD_VCO.t12 46.3367
R58 VDD_VCO.n358 VDD_VCO.t152 46.3367
R59 VDD_VCO.n439 VDD_VCO.t50 42.1692
R60 VDD_VCO.n549 VDD_VCO.t8 42.1692
R61 VDD_VCO.n617 VDD_VCO.t70 42.1692
R62 VDD_VCO.n61 VDD_VCO.t77 42.1692
R63 VDD_VCO.n380 VDD_VCO.t162 39.8225
R64 VDD_VCO.n328 VDD_VCO.t141 39.8225
R65 VDD_VCO.n436 VDD_VCO.t46 35.5427
R66 VDD_VCO.n552 VDD_VCO.t3 35.5427
R67 VDD_VCO.n620 VDD_VCO.t61 35.5427
R68 VDD_VCO.n58 VDD_VCO.t82 35.5427
R69 VDD_VCO.n308 VDD_VCO.t17 32.3281
R70 VDD_VCO.n361 VDD_VCO.t149 32.3281
R71 VDD_VCO.n406 VDD_VCO.t129 30.7234
R72 VDD_VCO.n582 VDD_VCO.t88 30.7234
R73 VDD_VCO.n650 VDD_VCO.t104 30.7234
R74 VDD_VCO.n28 VDD_VCO.t33 30.7234
R75 VDD_VCO.n433 VDD_VCO.t43 28.9162
R76 VDD_VCO.n555 VDD_VCO.t6 28.9162
R77 VDD_VCO.n623 VDD_VCO.t63 28.9162
R78 VDD_VCO.n55 VDD_VCO.t58 28.9162
R79 VDD_VCO.n409 VDD_VCO.t135 24.0969
R80 VDD_VCO.n579 VDD_VCO.t40 24.0969
R81 VDD_VCO.n647 VDD_VCO.t110 24.0969
R82 VDD_VCO.n31 VDD_VCO.t24 24.0969
R83 VDD_VCO.n171 VDD_VCO.t96 23.9239
R84 VDD_VCO.n608 VDD_VCO.t193 23.9239
R85 VDD_VCO.n430 VDD_VCO.t48 22.2897
R86 VDD_VCO.n558 VDD_VCO.t0 22.2897
R87 VDD_VCO.n626 VDD_VCO.t67 22.2897
R88 VDD_VCO.n52 VDD_VCO.t80 22.2897
R89 VDD_VCO.n412 VDD_VCO.t131 17.4704
R90 VDD_VCO.n576 VDD_VCO.t86 17.4704
R91 VDD_VCO.n644 VDD_VCO.t98 17.4704
R92 VDD_VCO.n34 VDD_VCO.t28 17.4704
R93 VDD_VCO.n292 VDD_VCO.t10 16.8707
R94 VDD_VCO.n345 VDD_VCO.t154 16.8707
R95 VDD_VCO.n298 VDD_VCO.t14 16.1643
R96 VDD_VCO.n351 VDD_VCO.t146 16.1643
R97 VDD_VCO.n427 VDD_VCO.t140 15.6632
R98 VDD_VCO.n561 VDD_VCO.t95 15.6632
R99 VDD_VCO.n629 VDD_VCO.t100 15.6632
R100 VDD_VCO.n49 VDD_VCO.t25 15.6632
R101 VDD_VCO.n415 VDD_VCO.t126 10.8439
R102 VDD_VCO.n573 VDD_VCO.t90 10.8439
R103 VDD_VCO.n641 VDD_VCO.t101 10.8439
R104 VDD_VCO.n37 VDD_VCO.t32 10.8439
R105 VDD_VCO.n380 VDD_VCO.n379 9.93878
R106 VDD_VCO.n328 VDD_VCO.n327 9.93878
R107 VDD_VCO.n386 VDD_VCO.t164 9.6712
R108 VDD_VCO.n334 VDD_VCO.t143 9.6712
R109 VDD_VCO.n424 VDD_VCO.t133 9.03664
R110 VDD_VCO.n564 VDD_VCO.t93 9.03664
R111 VDD_VCO.n632 VDD_VCO.t113 9.03664
R112 VDD_VCO.n46 VDD_VCO.t22 9.03664
R113 VDD_VCO.n181 VDD_VCO.n179 8.70445
R114 VDD_VCO.n603 VDD_VCO.n601 8.70445
R115 VDD_VCO.n373 VDD_VCO.t85 8.26313
R116 VDD_VCO.n321 VDD_VCO.t139 8.26313
R117 VDD_VCO.n299 VDD_VCO.n297 8.15819
R118 VDD_VCO.n352 VDD_VCO.n350 8.15819
R119 VDD_VCO.n706 VDD_VCO.n705 7.10822
R120 VDD_VCO.n598 VDD_VCO.n595 6.66125
R121 VDD_VCO.n173 VDD_VCO.t97 6.58259
R122 VDD_VCO.n184 VDD_VCO.n166 6.49073
R123 VDD_VCO.n611 VDD_VCO.t194 6.48786
R124 VDD_VCO.n313 VDD_VCO.n312 6.3005
R125 VDD_VCO.n312 VDD_VCO.n311 6.3005
R126 VDD_VCO.n592 VDD_VCO.n184 6.07717
R127 VDD_VCO.n317 VDD_VCO.n316 5.38954
R128 VDD_VCO.n447 VDD_VCO.n446 4.85019
R129 VDD_VCO VDD_VCO.n736 4.55945
R130 VDD_VCO.n400 VDD_VCO.n399 4.5005
R131 VDD_VCO.n445 VDD_VCO.n266 4.5005
R132 VDD_VCO.n189 VDD_VCO.n188 4.5005
R133 VDD_VCO.n613 VDD_VCO.n612 4.46272
R134 VDD_VCO.n379 VDD_VCO.t163 4.3192
R135 VDD_VCO.n390 VDD_VCO.n378 4.3192
R136 VDD_VCO.n327 VDD_VCO.t142 4.3192
R137 VDD_VCO.n338 VDD_VCO.n326 4.3192
R138 VDD_VCO.n377 VDD_VCO.n376 4.29708
R139 VDD_VCO.n325 VDD_VCO.n324 4.29333
R140 VDD_VCO.n418 VDD_VCO.t134 4.21737
R141 VDD_VCO.n570 VDD_VCO.t94 4.21737
R142 VDD_VCO.n638 VDD_VCO.t109 4.21737
R143 VDD_VCO.n40 VDD_VCO.t20 4.21737
R144 VDD_VCO.n367 VDD_VCO.n366 3.94094
R145 VDD_VCO.n291 VDD_VCO.t11 3.92746
R146 VDD_VCO.n318 VDD_VCO.n288 3.92746
R147 VDD_VCO.n344 VDD_VCO.t155 3.92746
R148 VDD_VCO.n211 VDD_VCO.n210 3.9192
R149 VDD_VCO.n521 VDD_VCO.n520 3.9192
R150 VDD_VCO.n140 VDD_VCO.n139 3.9192
R151 VDD_VCO.n23 VDD_VCO.n22 3.9192
R152 VDD_VCO.n192 VDD_VCO.t130 3.80738
R153 VDD_VCO.n502 VDD_VCO.t89 3.80738
R154 VDD_VCO.n121 VDD_VCO.t105 3.80738
R155 VDD_VCO.n4 VDD_VCO.t182 3.80738
R156 VDD_VCO.n170 VDD_VCO.t108 3.6405
R157 VDD_VCO.n170 VDD_VCO.n169 3.6405
R158 VDD_VCO.n594 VDD_VCO.t179 3.6405
R159 VDD_VCO.n594 VDD_VCO.n593 3.6405
R160 VDD_VCO.n301 VDD_VCO.n290 3.27746
R161 VDD_VCO.n354 VDD_VCO.n343 3.27746
R162 VDD_VCO.n374 VDD_VCO.n373 3.19668
R163 VDD_VCO.n322 VDD_VCO.n321 3.19668
R164 VDD_VCO.n183 VDD_VCO.n168 3.1505
R165 VDD_VCO.n168 VDD_VCO.n167 3.1505
R166 VDD_VCO.n173 VDD_VCO.n172 3.1505
R167 VDD_VCO.n172 VDD_VCO.n171 3.1505
R168 VDD_VCO.n182 VDD_VCO.n181 3.1505
R169 VDD_VCO.n181 VDD_VCO.n180 3.1505
R170 VDD_VCO.n179 VDD_VCO.n177 3.1505
R171 VDD_VCO.n179 VDD_VCO.n178 3.1505
R172 VDD_VCO.n176 VDD_VCO.n175 3.1505
R173 VDD_VCO.n175 VDD_VCO.n174 3.1505
R174 VDD_VCO.n601 VDD_VCO.n599 3.1505
R175 VDD_VCO.n601 VDD_VCO.n600 3.1505
R176 VDD_VCO.n610 VDD_VCO.n609 3.1505
R177 VDD_VCO.n609 VDD_VCO.n608 3.1505
R178 VDD_VCO.n607 VDD_VCO.n606 3.1505
R179 VDD_VCO.n606 VDD_VCO.n605 3.1505
R180 VDD_VCO.n604 VDD_VCO.n603 3.1505
R181 VDD_VCO.n603 VDD_VCO.n602 3.1505
R182 VDD_VCO.n598 VDD_VCO.n597 3.1505
R183 VDD_VCO.n597 VDD_VCO.n596 3.1505
R184 VDD_VCO.n372 VDD_VCO.n371 3.1505
R185 VDD_VCO.n375 VDD_VCO.n374 3.1505
R186 VDD_VCO.n385 VDD_VCO.n384 3.1505
R187 VDD_VCO.n384 VDD_VCO.n383 3.1505
R188 VDD_VCO.n382 VDD_VCO.n381 3.1505
R189 VDD_VCO.n388 VDD_VCO.n387 3.1505
R190 VDD_VCO.n310 VDD_VCO.n309 3.1505
R191 VDD_VCO.n309 VDD_VCO.n308 3.1505
R192 VDD_VCO.n307 VDD_VCO.n306 3.1505
R193 VDD_VCO.n306 VDD_VCO.n305 3.1505
R194 VDD_VCO.n304 VDD_VCO.n303 3.1505
R195 VDD_VCO.n303 VDD_VCO.n302 3.1505
R196 VDD_VCO.n300 VDD_VCO.n299 3.1505
R197 VDD_VCO.n299 VDD_VCO.n298 3.1505
R198 VDD_VCO.n297 VDD_VCO.n295 3.1505
R199 VDD_VCO.n297 VDD_VCO.n296 3.1505
R200 VDD_VCO.n294 VDD_VCO.n293 3.1505
R201 VDD_VCO.n363 VDD_VCO.n362 3.1505
R202 VDD_VCO.n362 VDD_VCO.n361 3.1505
R203 VDD_VCO.n360 VDD_VCO.n359 3.1505
R204 VDD_VCO.n359 VDD_VCO.n358 3.1505
R205 VDD_VCO.n357 VDD_VCO.n356 3.1505
R206 VDD_VCO.n356 VDD_VCO.n355 3.1505
R207 VDD_VCO.n353 VDD_VCO.n352 3.1505
R208 VDD_VCO.n352 VDD_VCO.n351 3.1505
R209 VDD_VCO.n350 VDD_VCO.n348 3.1505
R210 VDD_VCO.n350 VDD_VCO.n349 3.1505
R211 VDD_VCO.n347 VDD_VCO.n346 3.1505
R212 VDD_VCO.n333 VDD_VCO.n332 3.1505
R213 VDD_VCO.n332 VDD_VCO.n331 3.1505
R214 VDD_VCO.n330 VDD_VCO.n329 3.1505
R215 VDD_VCO.n336 VDD_VCO.n335 3.1505
R216 VDD_VCO.n323 VDD_VCO.n322 3.1505
R217 VDD_VCO.n320 VDD_VCO.n319 3.1505
R218 VDD_VCO.n442 VDD_VCO.n268 3.1505
R219 VDD_VCO.n268 VDD_VCO.n267 3.1505
R220 VDD_VCO.n441 VDD_VCO.n440 3.1505
R221 VDD_VCO.n440 VDD_VCO.n439 3.1505
R222 VDD_VCO.n438 VDD_VCO.n437 3.1505
R223 VDD_VCO.n437 VDD_VCO.n436 3.1505
R224 VDD_VCO.n435 VDD_VCO.n434 3.1505
R225 VDD_VCO.n434 VDD_VCO.n433 3.1505
R226 VDD_VCO.n432 VDD_VCO.n431 3.1505
R227 VDD_VCO.n431 VDD_VCO.n430 3.1505
R228 VDD_VCO.n429 VDD_VCO.n428 3.1505
R229 VDD_VCO.n428 VDD_VCO.n427 3.1505
R230 VDD_VCO.n426 VDD_VCO.n425 3.1505
R231 VDD_VCO.n425 VDD_VCO.n424 3.1505
R232 VDD_VCO.n423 VDD_VCO.n422 3.1505
R233 VDD_VCO.n422 VDD_VCO.n421 3.1505
R234 VDD_VCO.n420 VDD_VCO.n419 3.1505
R235 VDD_VCO.n419 VDD_VCO.n418 3.1505
R236 VDD_VCO.n417 VDD_VCO.n416 3.1505
R237 VDD_VCO.n416 VDD_VCO.n415 3.1505
R238 VDD_VCO.n414 VDD_VCO.n413 3.1505
R239 VDD_VCO.n413 VDD_VCO.n412 3.1505
R240 VDD_VCO.n411 VDD_VCO.n410 3.1505
R241 VDD_VCO.n410 VDD_VCO.n409 3.1505
R242 VDD_VCO.n408 VDD_VCO.n407 3.1505
R243 VDD_VCO.n407 VDD_VCO.n406 3.1505
R244 VDD_VCO.n405 VDD_VCO.n404 3.1505
R245 VDD_VCO.n404 VDD_VCO.n403 3.1505
R246 VDD_VCO.n270 VDD_VCO.n269 3.1505
R247 VDD_VCO.n273 VDD_VCO.n272 3.1505
R248 VDD_VCO.n275 VDD_VCO.n274 3.1505
R249 VDD_VCO.n278 VDD_VCO.n277 3.1505
R250 VDD_VCO.n280 VDD_VCO.n279 3.1505
R251 VDD_VCO.n283 VDD_VCO.n282 3.1505
R252 VDD_VCO.n287 VDD_VCO.n286 3.1505
R253 VDD_VCO.n240 VDD_VCO.n239 3.1505
R254 VDD_VCO.n238 VDD_VCO.n237 3.1505
R255 VDD_VCO.n236 VDD_VCO.n235 3.1505
R256 VDD_VCO.n234 VDD_VCO.n233 3.1505
R257 VDD_VCO.n232 VDD_VCO.n231 3.1505
R258 VDD_VCO.n230 VDD_VCO.n229 3.1505
R259 VDD_VCO.n228 VDD_VCO.n227 3.1505
R260 VDD_VCO.n226 VDD_VCO.n225 3.1505
R261 VDD_VCO.n224 VDD_VCO.n223 3.1505
R262 VDD_VCO.n222 VDD_VCO.n221 3.1505
R263 VDD_VCO.n220 VDD_VCO.n219 3.1505
R264 VDD_VCO.n218 VDD_VCO.n217 3.1505
R265 VDD_VCO.n216 VDD_VCO.n215 3.1505
R266 VDD_VCO.n214 VDD_VCO.n213 3.1505
R267 VDD_VCO.n258 VDD_VCO.n257 3.1505
R268 VDD_VCO.n255 VDD_VCO.n254 3.1505
R269 VDD_VCO.n251 VDD_VCO.n250 3.1505
R270 VDD_VCO.n248 VDD_VCO.n247 3.1505
R271 VDD_VCO.n245 VDD_VCO.n244 3.1505
R272 VDD_VCO.n262 VDD_VCO.n261 3.1505
R273 VDD_VCO.n243 VDD_VCO.n242 3.1505
R274 VDD_VCO.n449 VDD_VCO.n448 3.1505
R275 VDD_VCO.n451 VDD_VCO.n450 3.1505
R276 VDD_VCO.n453 VDD_VCO.n452 3.1505
R277 VDD_VCO.n455 VDD_VCO.n454 3.1505
R278 VDD_VCO.n457 VDD_VCO.n456 3.1505
R279 VDD_VCO.n459 VDD_VCO.n458 3.1505
R280 VDD_VCO.n461 VDD_VCO.n460 3.1505
R281 VDD_VCO.n463 VDD_VCO.n462 3.1505
R282 VDD_VCO.n465 VDD_VCO.n464 3.1505
R283 VDD_VCO.n467 VDD_VCO.n466 3.1505
R284 VDD_VCO.n469 VDD_VCO.n468 3.1505
R285 VDD_VCO.n471 VDD_VCO.n470 3.1505
R286 VDD_VCO.n473 VDD_VCO.n472 3.1505
R287 VDD_VCO.n475 VDD_VCO.n474 3.1505
R288 VDD_VCO.n539 VDD_VCO.n538 3.1505
R289 VDD_VCO.n536 VDD_VCO.n535 3.1505
R290 VDD_VCO.n532 VDD_VCO.n531 3.1505
R291 VDD_VCO.n529 VDD_VCO.n528 3.1505
R292 VDD_VCO.n527 VDD_VCO.n526 3.1505
R293 VDD_VCO.n541 VDD_VCO.n540 3.1505
R294 VDD_VCO.n545 VDD_VCO.n544 3.1505
R295 VDD_VCO.n547 VDD_VCO.n546 3.1505
R296 VDD_VCO.n548 VDD_VCO.n547 3.1505
R297 VDD_VCO.n551 VDD_VCO.n550 3.1505
R298 VDD_VCO.n550 VDD_VCO.n549 3.1505
R299 VDD_VCO.n554 VDD_VCO.n553 3.1505
R300 VDD_VCO.n553 VDD_VCO.n552 3.1505
R301 VDD_VCO.n557 VDD_VCO.n556 3.1505
R302 VDD_VCO.n556 VDD_VCO.n555 3.1505
R303 VDD_VCO.n560 VDD_VCO.n559 3.1505
R304 VDD_VCO.n559 VDD_VCO.n558 3.1505
R305 VDD_VCO.n563 VDD_VCO.n562 3.1505
R306 VDD_VCO.n562 VDD_VCO.n561 3.1505
R307 VDD_VCO.n566 VDD_VCO.n565 3.1505
R308 VDD_VCO.n565 VDD_VCO.n564 3.1505
R309 VDD_VCO.n569 VDD_VCO.n568 3.1505
R310 VDD_VCO.n568 VDD_VCO.n567 3.1505
R311 VDD_VCO.n572 VDD_VCO.n571 3.1505
R312 VDD_VCO.n571 VDD_VCO.n570 3.1505
R313 VDD_VCO.n575 VDD_VCO.n574 3.1505
R314 VDD_VCO.n574 VDD_VCO.n573 3.1505
R315 VDD_VCO.n578 VDD_VCO.n577 3.1505
R316 VDD_VCO.n577 VDD_VCO.n576 3.1505
R317 VDD_VCO.n581 VDD_VCO.n580 3.1505
R318 VDD_VCO.n580 VDD_VCO.n579 3.1505
R319 VDD_VCO.n584 VDD_VCO.n583 3.1505
R320 VDD_VCO.n583 VDD_VCO.n582 3.1505
R321 VDD_VCO.n587 VDD_VCO.n586 3.1505
R322 VDD_VCO.n586 VDD_VCO.n585 3.1505
R323 VDD_VCO.n478 VDD_VCO.n477 3.1505
R324 VDD_VCO.n480 VDD_VCO.n479 3.1505
R325 VDD_VCO.n483 VDD_VCO.n482 3.1505
R326 VDD_VCO.n485 VDD_VCO.n484 3.1505
R327 VDD_VCO.n488 VDD_VCO.n487 3.1505
R328 VDD_VCO.n490 VDD_VCO.n489 3.1505
R329 VDD_VCO.n494 VDD_VCO.n493 3.1505
R330 VDD_VCO.n685 VDD_VCO.n656 3.1505
R331 VDD_VCO.n700 VDD_VCO.n699 3.1505
R332 VDD_VCO.n698 VDD_VCO.n697 3.1505
R333 VDD_VCO.n695 VDD_VCO.n694 3.1505
R334 VDD_VCO.n693 VDD_VCO.n692 3.1505
R335 VDD_VCO.n690 VDD_VCO.n689 3.1505
R336 VDD_VCO.n688 VDD_VCO.n687 3.1505
R337 VDD_VCO.n704 VDD_VCO.n703 3.1505
R338 VDD_VCO.n658 VDD_VCO.n657 3.1505
R339 VDD_VCO.n660 VDD_VCO.n659 3.1505
R340 VDD_VCO.n662 VDD_VCO.n661 3.1505
R341 VDD_VCO.n664 VDD_VCO.n663 3.1505
R342 VDD_VCO.n666 VDD_VCO.n665 3.1505
R343 VDD_VCO.n668 VDD_VCO.n667 3.1505
R344 VDD_VCO.n670 VDD_VCO.n669 3.1505
R345 VDD_VCO.n672 VDD_VCO.n671 3.1505
R346 VDD_VCO.n674 VDD_VCO.n673 3.1505
R347 VDD_VCO.n676 VDD_VCO.n675 3.1505
R348 VDD_VCO.n678 VDD_VCO.n677 3.1505
R349 VDD_VCO.n680 VDD_VCO.n679 3.1505
R350 VDD_VCO.n682 VDD_VCO.n681 3.1505
R351 VDD_VCO.n684 VDD_VCO.n683 3.1505
R352 VDD_VCO.n146 VDD_VCO.n145 3.1505
R353 VDD_VCO.n148 VDD_VCO.n147 3.1505
R354 VDD_VCO.n151 VDD_VCO.n150 3.1505
R355 VDD_VCO.n155 VDD_VCO.n154 3.1505
R356 VDD_VCO.n158 VDD_VCO.n157 3.1505
R357 VDD_VCO.n161 VDD_VCO.n160 3.1505
R358 VDD_VCO.n143 VDD_VCO.n142 3.1505
R359 VDD_VCO.n165 VDD_VCO.n164 3.1505
R360 VDD_VCO.n616 VDD_VCO.n615 3.1505
R361 VDD_VCO.n615 VDD_VCO.n614 3.1505
R362 VDD_VCO.n619 VDD_VCO.n618 3.1505
R363 VDD_VCO.n618 VDD_VCO.n617 3.1505
R364 VDD_VCO.n622 VDD_VCO.n621 3.1505
R365 VDD_VCO.n621 VDD_VCO.n620 3.1505
R366 VDD_VCO.n625 VDD_VCO.n624 3.1505
R367 VDD_VCO.n624 VDD_VCO.n623 3.1505
R368 VDD_VCO.n628 VDD_VCO.n627 3.1505
R369 VDD_VCO.n627 VDD_VCO.n626 3.1505
R370 VDD_VCO.n631 VDD_VCO.n630 3.1505
R371 VDD_VCO.n630 VDD_VCO.n629 3.1505
R372 VDD_VCO.n634 VDD_VCO.n633 3.1505
R373 VDD_VCO.n633 VDD_VCO.n632 3.1505
R374 VDD_VCO.n637 VDD_VCO.n636 3.1505
R375 VDD_VCO.n636 VDD_VCO.n635 3.1505
R376 VDD_VCO.n640 VDD_VCO.n639 3.1505
R377 VDD_VCO.n639 VDD_VCO.n638 3.1505
R378 VDD_VCO.n643 VDD_VCO.n642 3.1505
R379 VDD_VCO.n642 VDD_VCO.n641 3.1505
R380 VDD_VCO.n646 VDD_VCO.n645 3.1505
R381 VDD_VCO.n645 VDD_VCO.n644 3.1505
R382 VDD_VCO.n649 VDD_VCO.n648 3.1505
R383 VDD_VCO.n648 VDD_VCO.n647 3.1505
R384 VDD_VCO.n652 VDD_VCO.n651 3.1505
R385 VDD_VCO.n651 VDD_VCO.n650 3.1505
R386 VDD_VCO.n655 VDD_VCO.n654 3.1505
R387 VDD_VCO.n654 VDD_VCO.n653 3.1505
R388 VDD_VCO.n27 VDD_VCO.n26 3.1505
R389 VDD_VCO.n26 VDD_VCO.n25 3.1505
R390 VDD_VCO.n30 VDD_VCO.n29 3.1505
R391 VDD_VCO.n29 VDD_VCO.n28 3.1505
R392 VDD_VCO.n33 VDD_VCO.n32 3.1505
R393 VDD_VCO.n32 VDD_VCO.n31 3.1505
R394 VDD_VCO.n36 VDD_VCO.n35 3.1505
R395 VDD_VCO.n35 VDD_VCO.n34 3.1505
R396 VDD_VCO.n39 VDD_VCO.n38 3.1505
R397 VDD_VCO.n38 VDD_VCO.n37 3.1505
R398 VDD_VCO.n42 VDD_VCO.n41 3.1505
R399 VDD_VCO.n41 VDD_VCO.n40 3.1505
R400 VDD_VCO.n45 VDD_VCO.n44 3.1505
R401 VDD_VCO.n44 VDD_VCO.n43 3.1505
R402 VDD_VCO.n48 VDD_VCO.n47 3.1505
R403 VDD_VCO.n47 VDD_VCO.n46 3.1505
R404 VDD_VCO.n51 VDD_VCO.n50 3.1505
R405 VDD_VCO.n50 VDD_VCO.n49 3.1505
R406 VDD_VCO.n54 VDD_VCO.n53 3.1505
R407 VDD_VCO.n53 VDD_VCO.n52 3.1505
R408 VDD_VCO.n57 VDD_VCO.n56 3.1505
R409 VDD_VCO.n56 VDD_VCO.n55 3.1505
R410 VDD_VCO.n60 VDD_VCO.n59 3.1505
R411 VDD_VCO.n59 VDD_VCO.n58 3.1505
R412 VDD_VCO.n63 VDD_VCO.n62 3.1505
R413 VDD_VCO.n62 VDD_VCO.n61 3.1505
R414 VDD_VCO.n65 VDD_VCO.n64 3.1505
R415 VDD_VCO.n87 VDD_VCO.n86 3.1505
R416 VDD_VCO.n83 VDD_VCO.n82 3.1505
R417 VDD_VCO.n80 VDD_VCO.n79 3.1505
R418 VDD_VCO.n76 VDD_VCO.n75 3.1505
R419 VDD_VCO.n73 VDD_VCO.n72 3.1505
R420 VDD_VCO.n70 VDD_VCO.n69 3.1505
R421 VDD_VCO.n89 VDD_VCO.n88 3.1505
R422 VDD_VCO.n68 VDD_VCO.n67 3.1505
R423 VDD_VCO.n92 VDD_VCO.n91 3.1505
R424 VDD_VCO.n91 VDD_VCO.n90 3.1505
R425 VDD_VCO.n94 VDD_VCO.n93 3.1505
R426 VDD_VCO.n96 VDD_VCO.n95 3.1505
R427 VDD_VCO.n98 VDD_VCO.n97 3.1505
R428 VDD_VCO.n100 VDD_VCO.n99 3.1505
R429 VDD_VCO.n102 VDD_VCO.n101 3.1505
R430 VDD_VCO.n104 VDD_VCO.n103 3.1505
R431 VDD_VCO.n106 VDD_VCO.n105 3.1505
R432 VDD_VCO.n108 VDD_VCO.n107 3.1505
R433 VDD_VCO.n110 VDD_VCO.n109 3.1505
R434 VDD_VCO.n112 VDD_VCO.n111 3.1505
R435 VDD_VCO.n114 VDD_VCO.n113 3.1505
R436 VDD_VCO.n116 VDD_VCO.n115 3.1505
R437 VDD_VCO.n118 VDD_VCO.n117 3.1505
R438 VDD_VCO.n722 VDD_VCO.n721 3.1505
R439 VDD_VCO.n718 VDD_VCO.n717 3.1505
R440 VDD_VCO.n715 VDD_VCO.n714 3.1505
R441 VDD_VCO.n713 VDD_VCO.n712 3.1505
R442 VDD_VCO.n710 VDD_VCO.n709 3.1505
R443 VDD_VCO.n724 VDD_VCO.n723 3.1505
R444 VDD_VCO.n708 VDD_VCO.n707 3.1505
R445 VDD_VCO.n728 VDD_VCO.n727 3.10174
R446 VDD_VCO.n729 VDD_VCO.n728 3.081
R447 VDD_VCO.n211 VDD_VCO.n208 3.07111
R448 VDD_VCO.n521 VDD_VCO.n518 3.07111
R449 VDD_VCO.n140 VDD_VCO.n137 3.07111
R450 VDD_VCO.n23 VDD_VCO.n20 3.07111
R451 VDD_VCO.n247 VDD_VCO.n246 3.001
R452 VDD_VCO.n250 VDD_VCO.n249 3.001
R453 VDD_VCO.n254 VDD_VCO.n253 3.001
R454 VDD_VCO.n531 VDD_VCO.n530 3.001
R455 VDD_VCO.n535 VDD_VCO.n534 3.001
R456 VDD_VCO.n160 VDD_VCO.n159 3.001
R457 VDD_VCO.n157 VDD_VCO.n156 3.001
R458 VDD_VCO.n154 VDD_VCO.n153 3.001
R459 VDD_VCO.n150 VDD_VCO.n149 3.001
R460 VDD_VCO.n72 VDD_VCO.n71 3.001
R461 VDD_VCO.n75 VDD_VCO.n74 3.001
R462 VDD_VCO.n79 VDD_VCO.n78 3.001
R463 VDD_VCO.n82 VDD_VCO.n81 3.001
R464 VDD_VCO.n369 VDD_VCO.n368 2.96108
R465 VDD_VCO.n592 VDD_VCO.n591 2.86102
R466 VDD_VCO VDD_VCO.n170 2.82941
R467 VDD_VCO VDD_VCO.n594 2.82941
R468 VDD_VCO.n206 VDD_VCO.n205 2.64616
R469 VDD_VCO.n516 VDD_VCO.n515 2.64616
R470 VDD_VCO.n135 VDD_VCO.n134 2.64616
R471 VDD_VCO.n18 VDD_VCO.n17 2.64616
R472 VDD_VCO.n590 VDD_VCO.n499 2.6255
R473 VDD_VCO.n393 VDD_VCO.n377 2.46744
R474 VDD_VCO.n421 VDD_VCO.t125 2.41014
R475 VDD_VCO.n567 VDD_VCO.t39 2.41014
R476 VDD_VCO.n635 VDD_VCO.t106 2.41014
R477 VDD_VCO.n43 VDD_VCO.t29 2.41014
R478 VDD_VCO.n612 VDD_VCO.n611 2.25606
R479 VDD_VCO.n732 VDD_VCO.n731 2.2505
R480 VDD_VCO.n717 VDD_VCO.n716 2.03394
R481 VDD_VCO.n712 VDD_VCO.n711 2.03394
R482 VDD_VCO.n272 VDD_VCO.n271 2.03336
R483 VDD_VCO.n544 VDD_VCO.n543 2.03336
R484 VDD_VCO.n277 VDD_VCO.n276 2.03326
R485 VDD_VCO.n282 VDD_VCO.n281 2.03326
R486 VDD_VCO.n487 VDD_VCO.n486 2.03326
R487 VDD_VCO.n493 VDD_VCO.n492 2.03326
R488 VDD_VCO.n703 VDD_VCO.n702 2.03326
R489 VDD_VCO.n697 VDD_VCO.n696 2.03326
R490 VDD_VCO.n692 VDD_VCO.n691 2.03326
R491 VDD_VCO.n687 VDD_VCO.n686 2.03326
R492 VDD_VCO.n341 VDD_VCO.n325 2.02931
R493 VDD_VCO.n261 VDD_VCO.n260 1.88586
R494 VDD_VCO.n286 VDD_VCO.n285 1.87058
R495 VDD_VCO.n365 VDD_VCO.n364 1.85344
R496 VDD_VCO.n208 VDD_VCO.t56 1.8205
R497 VDD_VCO.n208 VDD_VCO.n207 1.8205
R498 VDD_VCO.n210 VDD_VCO.t55 1.8205
R499 VDD_VCO.n210 VDD_VCO.n209 1.8205
R500 VDD_VCO.n191 VDD_VCO.t132 1.8205
R501 VDD_VCO.n191 VDD_VCO.n190 1.8205
R502 VDD_VCO.n194 VDD_VCO.t171 1.8205
R503 VDD_VCO.n194 VDD_VCO.n193 1.8205
R504 VDD_VCO.n197 VDD_VCO.t172 1.8205
R505 VDD_VCO.n197 VDD_VCO.n196 1.8205
R506 VDD_VCO.n200 VDD_VCO.t49 1.8205
R507 VDD_VCO.n200 VDD_VCO.n199 1.8205
R508 VDD_VCO.n203 VDD_VCO.t47 1.8205
R509 VDD_VCO.n203 VDD_VCO.n202 1.8205
R510 VDD_VCO.n518 VDD_VCO.t9 1.8205
R511 VDD_VCO.n518 VDD_VCO.n517 1.8205
R512 VDD_VCO.n520 VDD_VCO.t7 1.8205
R513 VDD_VCO.n520 VDD_VCO.n519 1.8205
R514 VDD_VCO.n501 VDD_VCO.t87 1.8205
R515 VDD_VCO.n501 VDD_VCO.n500 1.8205
R516 VDD_VCO.n504 VDD_VCO.t159 1.8205
R517 VDD_VCO.n504 VDD_VCO.n503 1.8205
R518 VDD_VCO.n507 VDD_VCO.t158 1.8205
R519 VDD_VCO.n507 VDD_VCO.n506 1.8205
R520 VDD_VCO.n510 VDD_VCO.t57 1.8205
R521 VDD_VCO.n510 VDD_VCO.n509 1.8205
R522 VDD_VCO.n513 VDD_VCO.t38 1.8205
R523 VDD_VCO.n513 VDD_VCO.n512 1.8205
R524 VDD_VCO.n137 VDD_VCO.t71 1.8205
R525 VDD_VCO.n137 VDD_VCO.n136 1.8205
R526 VDD_VCO.n139 VDD_VCO.t64 1.8205
R527 VDD_VCO.n139 VDD_VCO.n138 1.8205
R528 VDD_VCO.n120 VDD_VCO.t99 1.8205
R529 VDD_VCO.n120 VDD_VCO.n119 1.8205
R530 VDD_VCO.n123 VDD_VCO.t190 1.8205
R531 VDD_VCO.n123 VDD_VCO.n122 1.8205
R532 VDD_VCO.n126 VDD_VCO.t189 1.8205
R533 VDD_VCO.n126 VDD_VCO.n125 1.8205
R534 VDD_VCO.n129 VDD_VCO.t76 1.8205
R535 VDD_VCO.n129 VDD_VCO.n128 1.8205
R536 VDD_VCO.n132 VDD_VCO.t62 1.8205
R537 VDD_VCO.n132 VDD_VCO.n131 1.8205
R538 VDD_VCO.n20 VDD_VCO.t188 1.8205
R539 VDD_VCO.n20 VDD_VCO.n19 1.8205
R540 VDD_VCO.n22 VDD_VCO.t183 1.8205
R541 VDD_VCO.n22 VDD_VCO.n21 1.8205
R542 VDD_VCO.n3 VDD_VCO.t122 1.8205
R543 VDD_VCO.n3 VDD_VCO.n2 1.8205
R544 VDD_VCO.n6 VDD_VCO.t21 1.8205
R545 VDD_VCO.n6 VDD_VCO.n5 1.8205
R546 VDD_VCO.n9 VDD_VCO.t23 1.8205
R547 VDD_VCO.n9 VDD_VCO.n8 1.8205
R548 VDD_VCO.n12 VDD_VCO.t81 1.8205
R549 VDD_VCO.n12 VDD_VCO.n11 1.8205
R550 VDD_VCO.n15 VDD_VCO.t83 1.8205
R551 VDD_VCO.n15 VDD_VCO.n14 1.8205
R552 VDD_VCO.n242 VDD_VCO.n241 1.72716
R553 VDD_VCO.n526 VDD_VCO.n525 1.72716
R554 VDD_VCO.n164 VDD_VCO.n163 1.72716
R555 VDD_VCO.n67 VDD_VCO.n66 1.72716
R556 VDD_VCO.n257 VDD_VCO.n256 1.72703
R557 VDD_VCO.n477 VDD_VCO.n476 1.72703
R558 VDD_VCO.n482 VDD_VCO.n481 1.72703
R559 VDD_VCO.n538 VDD_VCO.n537 1.72703
R560 VDD_VCO.n145 VDD_VCO.n144 1.72703
R561 VDD_VCO.n721 VDD_VCO.n720 1.72703
R562 VDD_VCO.n86 VDD_VCO.n85 1.72703
R563 VDD_VCO.n395 VDD_VCO.n394 1.60323
R564 VDD_VCO.n370 VDD_VCO.n318 1.52757
R565 VDD_VCO.n368 VDD_VCO.n367 1.43172
R566 VDD_VCO.n192 VDD_VCO.n191 1.42427
R567 VDD_VCO.n195 VDD_VCO.n194 1.42427
R568 VDD_VCO.n198 VDD_VCO.n197 1.42427
R569 VDD_VCO.n201 VDD_VCO.n200 1.42427
R570 VDD_VCO.n204 VDD_VCO.n203 1.42427
R571 VDD_VCO.n502 VDD_VCO.n501 1.42427
R572 VDD_VCO.n505 VDD_VCO.n504 1.42427
R573 VDD_VCO.n508 VDD_VCO.n507 1.42427
R574 VDD_VCO.n511 VDD_VCO.n510 1.42427
R575 VDD_VCO.n514 VDD_VCO.n513 1.42427
R576 VDD_VCO.n121 VDD_VCO.n120 1.42427
R577 VDD_VCO.n124 VDD_VCO.n123 1.42427
R578 VDD_VCO.n127 VDD_VCO.n126 1.42427
R579 VDD_VCO.n130 VDD_VCO.n129 1.42427
R580 VDD_VCO.n133 VDD_VCO.n132 1.42427
R581 VDD_VCO.n4 VDD_VCO.n3 1.42427
R582 VDD_VCO.n7 VDD_VCO.n6 1.42427
R583 VDD_VCO.n10 VDD_VCO.n9 1.42427
R584 VDD_VCO.n13 VDD_VCO.n12 1.42427
R585 VDD_VCO.n16 VDD_VCO.n15 1.42427
R586 VDD_VCO.n368 VDD_VCO.n341 1.34003
R587 VDD_VCO.n499 VDD_VCO.n497 1.31777
R588 VDD_VCO.n394 VDD_VCO.n370 1.30655
R589 VDD_VCO.n499 VDD_VCO.n498 1.27368
R590 VDD_VCO.n612 VDD_VCO.n592 1.18161
R591 VDD_VCO.n206 VDD_VCO.n204 1.16194
R592 VDD_VCO.n516 VDD_VCO.n514 1.16194
R593 VDD_VCO.n135 VDD_VCO.n133 1.16194
R594 VDD_VCO.n18 VDD_VCO.n16 1.16194
R595 VDD_VCO.n264 VDD_VCO.n263 1.08868
R596 VDD_VCO.n163 VDD_VCO.n162 0.950516
R597 VDD_VCO.n85 VDD_VCO.n84 0.950315
R598 VDD_VCO.n720 VDD_VCO.n719 0.950315
R599 VDD_VCO.n734 VDD_VCO.n733 0.941249
R600 VDD_VCO.n188 VDD_VCO.n187 0.916864
R601 VDD_VCO.n736 VDD_VCO.n735 0.899828
R602 VDD_VCO.n392 VDD_VCO.n391 0.898937
R603 VDD_VCO.n340 VDD_VCO.n339 0.898718
R604 VDD_VCO.n397 VDD_VCO.n396 0.859591
R605 VDD_VCO.n285 VDD_VCO.n284 0.754483
R606 VDD_VCO.n260 VDD_VCO.n259 0.745201
R607 VDD_VCO.n728 VDD_VCO.n726 0.718169
R608 VDD_VCO.n290 VDD_VCO.t13 0.6505
R609 VDD_VCO.n290 VDD_VCO.n289 0.6505
R610 VDD_VCO.n343 VDD_VCO.t153 0.6505
R611 VDD_VCO.n343 VDD_VCO.n342 0.6505
R612 VDD_VCO.n195 VDD_VCO.n192 0.562605
R613 VDD_VCO.n198 VDD_VCO.n195 0.562605
R614 VDD_VCO.n201 VDD_VCO.n198 0.562605
R615 VDD_VCO.n204 VDD_VCO.n201 0.562605
R616 VDD_VCO.n505 VDD_VCO.n502 0.562605
R617 VDD_VCO.n508 VDD_VCO.n505 0.562605
R618 VDD_VCO.n511 VDD_VCO.n508 0.562605
R619 VDD_VCO.n514 VDD_VCO.n511 0.562605
R620 VDD_VCO.n124 VDD_VCO.n121 0.562605
R621 VDD_VCO.n127 VDD_VCO.n124 0.562605
R622 VDD_VCO.n130 VDD_VCO.n127 0.562605
R623 VDD_VCO.n133 VDD_VCO.n130 0.562605
R624 VDD_VCO.n7 VDD_VCO.n4 0.562605
R625 VDD_VCO.n10 VDD_VCO.n7 0.562605
R626 VDD_VCO.n13 VDD_VCO.n10 0.562605
R627 VDD_VCO.n16 VDD_VCO.n13 0.562605
R628 VDD_VCO.n543 VDD_VCO.n542 0.560113
R629 VDD_VCO.n492 VDD_VCO.n491 0.559871
R630 VDD_VCO.n702 VDD_VCO.n701 0.559871
R631 VDD_VCO.n376 VDD_VCO.n375 0.526923
R632 VDD_VCO.n324 VDD_VCO.n323 0.526923
R633 VDD_VCO.n212 VDD_VCO.n211 0.418343
R634 VDD_VCO.n522 VDD_VCO.n521 0.418343
R635 VDD_VCO.n141 VDD_VCO.n140 0.418343
R636 VDD_VCO.n24 VDD_VCO.n23 0.418343
R637 VDD_VCO.n212 VDD_VCO.n206 0.41547
R638 VDD_VCO.n522 VDD_VCO.n516 0.41547
R639 VDD_VCO.n141 VDD_VCO.n135 0.41547
R640 VDD_VCO.n24 VDD_VCO.n18 0.41547
R641 VDD_VCO.n726 VDD_VCO.n725 0.412906
R642 VDD_VCO.n735 VDD_VCO.n734 0.367012
R643 VDD_VCO.n393 VDD_VCO.n392 0.348354
R644 VDD_VCO.n399 VDD_VCO.n398 0.286864
R645 VDD_VCO.n341 VDD_VCO.n340 0.272998
R646 VDD_VCO.n316 VDD_VCO.n315 0.2719
R647 VDD_VCO.n398 VDD_VCO.n397 0.229591
R648 VDD_VCO.n265 VDD_VCO.n264 0.229591
R649 VDD_VCO.n186 VDD_VCO.n185 0.222053
R650 VDD_VCO.n187 VDD_VCO.n186 0.222053
R651 VDD_VCO.n293 VDD_VCO.n292 0.209658
R652 VDD_VCO.n346 VDD_VCO.n345 0.209419
R653 VDD_VCO.n442 VDD_VCO.n441 0.185
R654 VDD_VCO.n441 VDD_VCO.n438 0.185
R655 VDD_VCO.n438 VDD_VCO.n435 0.185
R656 VDD_VCO.n435 VDD_VCO.n432 0.185
R657 VDD_VCO.n432 VDD_VCO.n429 0.185
R658 VDD_VCO.n429 VDD_VCO.n426 0.185
R659 VDD_VCO.n426 VDD_VCO.n423 0.185
R660 VDD_VCO.n423 VDD_VCO.n420 0.185
R661 VDD_VCO.n420 VDD_VCO.n417 0.185
R662 VDD_VCO.n417 VDD_VCO.n414 0.185
R663 VDD_VCO.n414 VDD_VCO.n411 0.185
R664 VDD_VCO.n411 VDD_VCO.n408 0.185
R665 VDD_VCO.n408 VDD_VCO.n405 0.185
R666 VDD_VCO.n240 VDD_VCO.n238 0.185
R667 VDD_VCO.n238 VDD_VCO.n236 0.185
R668 VDD_VCO.n236 VDD_VCO.n234 0.185
R669 VDD_VCO.n234 VDD_VCO.n232 0.185
R670 VDD_VCO.n232 VDD_VCO.n230 0.185
R671 VDD_VCO.n230 VDD_VCO.n228 0.185
R672 VDD_VCO.n228 VDD_VCO.n226 0.185
R673 VDD_VCO.n226 VDD_VCO.n224 0.185
R674 VDD_VCO.n224 VDD_VCO.n222 0.185
R675 VDD_VCO.n222 VDD_VCO.n220 0.185
R676 VDD_VCO.n220 VDD_VCO.n218 0.185
R677 VDD_VCO.n218 VDD_VCO.n216 0.185
R678 VDD_VCO.n216 VDD_VCO.n214 0.185
R679 VDD_VCO.n451 VDD_VCO.n449 0.185
R680 VDD_VCO.n453 VDD_VCO.n451 0.185
R681 VDD_VCO.n455 VDD_VCO.n453 0.185
R682 VDD_VCO.n457 VDD_VCO.n455 0.185
R683 VDD_VCO.n459 VDD_VCO.n457 0.185
R684 VDD_VCO.n461 VDD_VCO.n459 0.185
R685 VDD_VCO.n463 VDD_VCO.n461 0.185
R686 VDD_VCO.n465 VDD_VCO.n463 0.185
R687 VDD_VCO.n467 VDD_VCO.n465 0.185
R688 VDD_VCO.n469 VDD_VCO.n467 0.185
R689 VDD_VCO.n471 VDD_VCO.n469 0.185
R690 VDD_VCO.n473 VDD_VCO.n471 0.185
R691 VDD_VCO.n475 VDD_VCO.n473 0.185
R692 VDD_VCO.n551 VDD_VCO.n548 0.185
R693 VDD_VCO.n554 VDD_VCO.n551 0.185
R694 VDD_VCO.n557 VDD_VCO.n554 0.185
R695 VDD_VCO.n560 VDD_VCO.n557 0.185
R696 VDD_VCO.n563 VDD_VCO.n560 0.185
R697 VDD_VCO.n566 VDD_VCO.n563 0.185
R698 VDD_VCO.n569 VDD_VCO.n566 0.185
R699 VDD_VCO.n572 VDD_VCO.n569 0.185
R700 VDD_VCO.n575 VDD_VCO.n572 0.185
R701 VDD_VCO.n578 VDD_VCO.n575 0.185
R702 VDD_VCO.n581 VDD_VCO.n578 0.185
R703 VDD_VCO.n584 VDD_VCO.n581 0.185
R704 VDD_VCO.n587 VDD_VCO.n584 0.185
R705 VDD_VCO.n660 VDD_VCO.n658 0.185
R706 VDD_VCO.n662 VDD_VCO.n660 0.185
R707 VDD_VCO.n664 VDD_VCO.n662 0.185
R708 VDD_VCO.n666 VDD_VCO.n664 0.185
R709 VDD_VCO.n668 VDD_VCO.n666 0.185
R710 VDD_VCO.n670 VDD_VCO.n668 0.185
R711 VDD_VCO.n672 VDD_VCO.n670 0.185
R712 VDD_VCO.n674 VDD_VCO.n672 0.185
R713 VDD_VCO.n676 VDD_VCO.n674 0.185
R714 VDD_VCO.n678 VDD_VCO.n676 0.185
R715 VDD_VCO.n680 VDD_VCO.n678 0.185
R716 VDD_VCO.n682 VDD_VCO.n680 0.185
R717 VDD_VCO.n684 VDD_VCO.n682 0.185
R718 VDD_VCO.n619 VDD_VCO.n616 0.185
R719 VDD_VCO.n622 VDD_VCO.n619 0.185
R720 VDD_VCO.n625 VDD_VCO.n622 0.185
R721 VDD_VCO.n628 VDD_VCO.n625 0.185
R722 VDD_VCO.n631 VDD_VCO.n628 0.185
R723 VDD_VCO.n634 VDD_VCO.n631 0.185
R724 VDD_VCO.n637 VDD_VCO.n634 0.185
R725 VDD_VCO.n640 VDD_VCO.n637 0.185
R726 VDD_VCO.n643 VDD_VCO.n640 0.185
R727 VDD_VCO.n646 VDD_VCO.n643 0.185
R728 VDD_VCO.n649 VDD_VCO.n646 0.185
R729 VDD_VCO.n652 VDD_VCO.n649 0.185
R730 VDD_VCO.n655 VDD_VCO.n652 0.185
R731 VDD_VCO.n63 VDD_VCO.n60 0.185
R732 VDD_VCO.n60 VDD_VCO.n57 0.185
R733 VDD_VCO.n57 VDD_VCO.n54 0.185
R734 VDD_VCO.n54 VDD_VCO.n51 0.185
R735 VDD_VCO.n51 VDD_VCO.n48 0.185
R736 VDD_VCO.n48 VDD_VCO.n45 0.185
R737 VDD_VCO.n45 VDD_VCO.n42 0.185
R738 VDD_VCO.n42 VDD_VCO.n39 0.185
R739 VDD_VCO.n39 VDD_VCO.n36 0.185
R740 VDD_VCO.n36 VDD_VCO.n33 0.185
R741 VDD_VCO.n33 VDD_VCO.n30 0.185
R742 VDD_VCO.n30 VDD_VCO.n27 0.185
R743 VDD_VCO.n94 VDD_VCO.n92 0.185
R744 VDD_VCO.n96 VDD_VCO.n94 0.185
R745 VDD_VCO.n98 VDD_VCO.n96 0.185
R746 VDD_VCO.n100 VDD_VCO.n98 0.185
R747 VDD_VCO.n102 VDD_VCO.n100 0.185
R748 VDD_VCO.n104 VDD_VCO.n102 0.185
R749 VDD_VCO.n106 VDD_VCO.n104 0.185
R750 VDD_VCO.n108 VDD_VCO.n106 0.185
R751 VDD_VCO.n110 VDD_VCO.n108 0.185
R752 VDD_VCO.n112 VDD_VCO.n110 0.185
R753 VDD_VCO.n114 VDD_VCO.n112 0.185
R754 VDD_VCO.n116 VDD_VCO.n114 0.185
R755 VDD_VCO.n118 VDD_VCO.n116 0.185
R756 VDD_VCO.n478 VDD_VCO.n475 0.172236
R757 VDD_VCO.n184 VDD_VCO.n183 0.171026
R758 VDD_VCO.n273 VDD_VCO.n270 0.164136
R759 VDD_VCO.n275 VDD_VCO.n273 0.164136
R760 VDD_VCO.n278 VDD_VCO.n275 0.164136
R761 VDD_VCO.n280 VDD_VCO.n278 0.164136
R762 VDD_VCO.n283 VDD_VCO.n280 0.164136
R763 VDD_VCO.n287 VDD_VCO.n283 0.164136
R764 VDD_VCO.n245 VDD_VCO.n243 0.164136
R765 VDD_VCO.n248 VDD_VCO.n245 0.164136
R766 VDD_VCO.n251 VDD_VCO.n248 0.164136
R767 VDD_VCO.n258 VDD_VCO.n255 0.164136
R768 VDD_VCO.n262 VDD_VCO.n258 0.164136
R769 VDD_VCO.n529 VDD_VCO.n527 0.164136
R770 VDD_VCO.n532 VDD_VCO.n529 0.164136
R771 VDD_VCO.n539 VDD_VCO.n536 0.164136
R772 VDD_VCO.n541 VDD_VCO.n539 0.164136
R773 VDD_VCO.n545 VDD_VCO.n541 0.164136
R774 VDD_VCO.n480 VDD_VCO.n478 0.164136
R775 VDD_VCO.n483 VDD_VCO.n480 0.164136
R776 VDD_VCO.n485 VDD_VCO.n483 0.164136
R777 VDD_VCO.n488 VDD_VCO.n485 0.164136
R778 VDD_VCO.n490 VDD_VCO.n488 0.164136
R779 VDD_VCO.n494 VDD_VCO.n490 0.164136
R780 VDD_VCO.n704 VDD_VCO.n700 0.164136
R781 VDD_VCO.n700 VDD_VCO.n698 0.164136
R782 VDD_VCO.n698 VDD_VCO.n695 0.164136
R783 VDD_VCO.n695 VDD_VCO.n693 0.164136
R784 VDD_VCO.n693 VDD_VCO.n690 0.164136
R785 VDD_VCO.n690 VDD_VCO.n688 0.164136
R786 VDD_VCO.n688 VDD_VCO.n685 0.164136
R787 VDD_VCO.n165 VDD_VCO.n161 0.164136
R788 VDD_VCO.n161 VDD_VCO.n158 0.164136
R789 VDD_VCO.n158 VDD_VCO.n155 0.164136
R790 VDD_VCO.n151 VDD_VCO.n148 0.164136
R791 VDD_VCO.n148 VDD_VCO.n146 0.164136
R792 VDD_VCO.n146 VDD_VCO.n143 0.164136
R793 VDD_VCO.n70 VDD_VCO.n68 0.164136
R794 VDD_VCO.n73 VDD_VCO.n70 0.164136
R795 VDD_VCO.n76 VDD_VCO.n73 0.164136
R796 VDD_VCO.n83 VDD_VCO.n80 0.164136
R797 VDD_VCO.n87 VDD_VCO.n83 0.164136
R798 VDD_VCO.n89 VDD_VCO.n87 0.164136
R799 VDD_VCO.n724 VDD_VCO.n722 0.164136
R800 VDD_VCO.n722 VDD_VCO.n718 0.164136
R801 VDD_VCO.n718 VDD_VCO.n715 0.164136
R802 VDD_VCO.n715 VDD_VCO.n713 0.164136
R803 VDD_VCO.n713 VDD_VCO.n710 0.164136
R804 VDD_VCO.n710 VDD_VCO.n708 0.164136
R805 VDD_VCO.n255 VDD_VCO.n252 0.161682
R806 VDD_VCO.n536 VDD_VCO.n533 0.161682
R807 VDD_VCO.n152 VDD_VCO.n151 0.161682
R808 VDD_VCO.n80 VDD_VCO.n77 0.161682
R809 VDD_VCO.n446 VDD_VCO.n262 0.159829
R810 VDD_VCO.n527 VDD_VCO.n524 0.157591
R811 VDD_VCO.n395 VDD_VCO.n287 0.155743
R812 VDD_VCO.n243 VDD_VCO.n240 0.151536
R813 VDD_VCO.n68 VDD_VCO.n65 0.151536
R814 VDD_VCO.n730 VDD_VCO.n724 0.149409
R815 VDD_VCO.n183 VDD_VCO.n182 0.143789
R816 VDD_VCO.n599 VDD_VCO.n598 0.143789
R817 VDD_VCO.n325 VDD_VCO.n320 0.140912
R818 VDD_VCO.n27 VDD_VCO.n1 0.140679
R819 VDD_VCO.n685 VDD_VCO.n684 0.137873
R820 VDD_VCO.n588 VDD_VCO.n587 0.137055
R821 VDD_VCO.n591 VDD_VCO.n494 0.136132
R822 VDD_VCO.n405 VDD_VCO.n402 0.1346
R823 VDD_VCO.n377 VDD_VCO.n372 0.134192
R824 VDD_VCO.n252 VDD_VCO 0.130885
R825 VDD_VCO.n533 VDD_VCO 0.130885
R826 VDD_VCO.n152 VDD_VCO 0.130885
R827 VDD_VCO.n77 VDD_VCO 0.130885
R828 VDD_VCO.n449 VDD_VCO.n447 0.130485
R829 VDD_VCO.n177 VDD_VCO.n176 0.127211
R830 VDD_VCO.n607 VDD_VCO.n604 0.127211
R831 VDD_VCO.n387 VDD_VCO.n386 0.12598
R832 VDD_VCO.n335 VDD_VCO.n334 0.12598
R833 VDD_VCO.n381 VDD_VCO.n380 0.125861
R834 VDD_VCO.n329 VDD_VCO.n328 0.125861
R835 VDD_VCO.n176 VDD_VCO.n173 0.123658
R836 VDD_VCO.n610 VDD_VCO.n607 0.123658
R837 VDD_VCO.n548 VDD_VCO.n545 0.117173
R838 VDD_VCO.n92 VDD_VCO.n89 0.117173
R839 VDD_VCO.n310 VDD_VCO.n307 0.117038
R840 VDD_VCO.n307 VDD_VCO.n304 0.117038
R841 VDD_VCO.n295 VDD_VCO.n294 0.117038
R842 VDD_VCO.n365 VDD_VCO.n363 0.117038
R843 VDD_VCO.n363 VDD_VCO.n360 0.117038
R844 VDD_VCO.n360 VDD_VCO.n357 0.117038
R845 VDD_VCO.n348 VDD_VCO.n347 0.117038
R846 VDD_VCO.n443 VDD_VCO.n442 0.1139
R847 VDD_VCO.n313 VDD_VCO.n310 0.1055
R848 VDD_VCO.n388 VDD_VCO.n385 0.102773
R849 VDD_VCO.n385 VDD_VCO.n382 0.102773
R850 VDD_VCO.n336 VDD_VCO.n333 0.102773
R851 VDD_VCO.n333 VDD_VCO.n330 0.102773
R852 VDD_VCO VDD_VCO.n63 0.0968
R853 VDD_VCO.n611 VDD_VCO.n610 0.0952368
R854 VDD_VCO.n705 VDD_VCO.n704 0.0921364
R855 VDD_VCO.n65 VDD_VCO 0.0887
R856 VDD_VCO.n294 VDD_VCO.n291 0.0858846
R857 VDD_VCO.n347 VDD_VCO.n344 0.0858846
R858 VDD_VCO.n301 VDD_VCO.n300 0.0835769
R859 VDD_VCO.n354 VDD_VCO.n353 0.0835769
R860 VDD_VCO.n616 VDD_VCO.n613 0.0815
R861 VDD_VCO.n705 VDD_VCO.n655 0.0806
R862 VDD_VCO.n706 VDD_VCO.n118 0.0788
R863 VDD_VCO.n337 VDD_VCO.n336 0.0782273
R864 VDD_VCO.n182 VDD_VCO 0.0774737
R865 VDD_VCO.n599 VDD_VCO 0.0774737
R866 VDD_VCO.n389 VDD_VCO.n388 0.0772045
R867 VDD_VCO VDD_VCO.n372 0.0715526
R868 VDD_VCO VDD_VCO.n320 0.0715526
R869 VDD_VCO.n300 VDD_VCO 0.0708846
R870 VDD_VCO.n353 VDD_VCO 0.0708846
R871 VDD_VCO.n613 VDD_VCO.n165 0.0705364
R872 VDD_VCO.n708 VDD_VCO.n706 0.0595727
R873 VDD_VCO.n266 VDD_VCO.n265 0.0577727
R874 VDD_VCO.n382 VDD_VCO 0.0526591
R875 VDD_VCO.n330 VDD_VCO 0.0526591
R876 VDD_VCO.n177 VDD_VCO 0.0478684
R877 VDD_VCO.n604 VDD_VCO 0.0478684
R878 VDD_VCO.n295 VDD_VCO 0.0466538
R879 VDD_VCO.n348 VDD_VCO 0.0466538
R880 VDD_VCO.n394 VDD_VCO.n393 0.0423605
R881 VDD_VCO VDD_VCO.n212 0.0374231
R882 VDD_VCO VDD_VCO.n522 0.0374231
R883 VDD_VCO VDD_VCO.n141 0.0374231
R884 VDD_VCO VDD_VCO.n24 0.0374231
R885 VDD_VCO.n304 VDD_VCO.n301 0.0339615
R886 VDD_VCO.n357 VDD_VCO.n354 0.0339615
R887 VDD_VCO.n496 VDD_VCO.n495 0.0295068
R888 VDD_VCO.n497 VDD_VCO.n496 0.0295068
R889 VDD_VCO.n373 VDD_VCO 0.0253684
R890 VDD_VCO.n321 VDD_VCO 0.0253684
R891 VDD_VCO.n732 VDD_VCO.n0 0.0240501
R892 VDD_VCO.n731 VDD_VCO.n1 0.0210263
R893 VDD_VCO.n590 VDD_VCO.n589 0.0193182
R894 VDD_VCO.n391 VDD_VCO.n390 0.0178864
R895 VDD_VCO.n339 VDD_VCO.n338 0.0178864
R896 VDD_VCO.n317 VDD_VCO.n314 0.0178077
R897 VDD_VCO.n379 VDD_VCO 0.0148182
R898 VDD_VCO.n327 VDD_VCO 0.0148182
R899 VDD_VCO.n731 VDD_VCO.n730 0.0123421
R900 VDD_VCO.n314 VDD_VCO.n313 0.0120385
R901 VDD_VCO.n591 VDD_VCO.n590 0.011585
R902 VDD_VCO VDD_VCO.n735 0.010631
R903 VDD_VCO.n447 VDD_VCO.n189 0.0103779
R904 VDD_VCO.n370 VDD_VCO.n369 0.0099186
R905 VDD_VCO.n390 VDD_VCO.n389 0.00868182
R906 VDD_VCO.n733 VDD_VCO.n732 0.00787217
R907 VDD_VCO.n338 VDD_VCO.n337 0.00765909
R908 VDD_VCO.n367 VDD_VCO.n365 0.00742767
R909 VDD_VCO.n524 VDD_VCO.n523 0.00704545
R910 VDD_VCO.n400 VDD_VCO.n395 0.00672312
R911 VDD_VCO.n446 VDD_VCO.n445 0.00590945
R912 VDD_VCO.n401 VDD_VCO.n400 0.00459091
R913 VDD_VCO.n402 VDD_VCO.n401 0.00377273
R914 VDD_VCO.n444 VDD_VCO.n443 0.00377273
R915 VDD_VCO.n252 VDD_VCO.n251 0.00295455
R916 VDD_VCO.n533 VDD_VCO.n532 0.00295455
R917 VDD_VCO.n155 VDD_VCO.n152 0.00295455
R918 VDD_VCO.n77 VDD_VCO.n76 0.00295455
R919 VDD_VCO.n318 VDD_VCO.n317 0.00165385
R920 VDD_VCO.n445 VDD_VCO.n444 0.00131818
R921 VDD_VCO.n589 VDD_VCO.n588 0.00131818
R922 VDD_VCO.n730 VDD_VCO.n729 0.00128947
R923 VDD.t486 VDD.n412 57397.6
R924 VDD.t477 VDD.n451 57397.6
R925 VDD.t474 VDD.n270 57397.6
R926 VDD.n604 VDD.n603 37257.5
R927 VDD.t48 VDD.t203 9544.02
R928 VDD.n56 VDD.t549 2529.02
R929 VDD.n62 VDD 2301.38
R930 VDD.n563 VDD 2301.38
R931 VDD.n63 VDD.n62 1842.37
R932 VDD.n564 VDD.n563 1842.37
R933 VDD.n66 VDD.t368 1403.56
R934 VDD.n68 VDD.t637 1242.86
R935 VDD.n301 VDD.t509 1105.93
R936 VDD.n59 VDD.t505 1105.93
R937 VDD.t516 VDD.n53 1011.51
R938 VDD.t221 VDD.t339 961.905
R939 VDD.t667 VDD.t547 961.905
R940 VDD.t6 VDD.t511 961.905
R941 VDD.t321 VDD.t373 961.905
R942 VDD.t284 VDD.t653 961.905
R943 VDD.t436 VDD.t147 961.905
R944 VDD.n412 VDD.t423 864.287
R945 VDD.n451 VDD.t24 864.287
R946 VDD.n270 VDD.t461 864.287
R947 VDD.t513 VDD.n39 857.144
R948 VDD.t610 VDD.n43 857.144
R949 VDD.n62 VDD.t591 812.681
R950 VDD.n563 VDD.t621 812.681
R951 VDD.t98 VDD.n606 768.971
R952 VDD.t588 VDD.t156 765.152
R953 VDD.t331 VDD.t387 765.152
R954 VDD.t309 VDD.t414 765.152
R955 VDD.t160 VDD.t79 765.152
R956 VDD.t534 VDD.t686 765.152
R957 VDD.t457 VDD.t514 765.152
R958 VDD.t611 VDD.t281 765.152
R959 VDD.t463 VDD.t246 765.152
R960 VDD.t106 VDD.t239 765.152
R961 VDD.t3 VDD.t131 765.152
R962 VDD.t81 VDD.t21 765.152
R963 VDD.t290 VDD.t646 765.152
R964 VDD.t507 VDD.t218 765.152
R965 VDD.t425 VDD.t539 765.152
R966 VDD.t619 VDD.t635 765.152
R967 VDD.t545 VDD.t563 765.152
R968 VDD.t213 VDD.t337 765.152
R969 VDD.t346 VDD.t140 765.152
R970 VDD.t560 VDD.t149 765.152
R971 VDD.t335 VDD.t211 765.152
R972 VDD.t268 VDD.t623 765.152
R973 VDD.t163 VDD.t154 765.152
R974 VDD.t684 VDD.t537 765.152
R975 VDD.t520 VDD.t42 765.152
R976 VDD.t119 VDD.t642 765.152
R977 VDD.t103 VDD.t65 765.152
R978 VDD.t197 VDD.t593 765.152
R979 VDD.t385 VDD.t499 765.152
R980 VDD.t187 VDD.t613 765.152
R981 VDD.t192 VDD.t113 765.152
R982 VDD.t502 VDD.t471 765.152
R983 VDD.t615 VDD.t190 765.152
R984 VDD.t366 VDD.t551 765.152
R985 VDD.t639 VDD.t571 765.152
R986 VDD.t63 VDD.t101 765.152
R987 VDD.t226 VDD.t569 765.152
R988 VDD.t585 VDD.t216 765.152
R989 VDD.t333 VDD.t390 765.152
R990 VDD.t292 VDD.t38 765.152
R991 VDD.n298 VDD.t497 747.159
R992 VDD.n606 VDD.t153 677.782
R993 VDD.t311 VDD.t573 642.843
R994 VDD.n60 VDD.t543 581.375
R995 VDD VDD.n60 572.967
R996 VDD.n612 VDD.n611 555.557
R997 VDD VDD.t121 551.043
R998 VDD.n531 VDD.t40 480.199
R999 VDD.t368 VDD.t399 461.096
R1000 VDD.t368 VDD.t344 461.096
R1001 VDD.t341 VDD.t224 461.096
R1002 VDD.t522 VDD.t228 461.096
R1003 VDD.n31 VDD.t301 443.07
R1004 VDD.n603 VDD.n599 438.12
R1005 VDD.n597 VDD.t349 436.957
R1006 VDD VDD.n201 429.187
R1007 VDD VDD.n169 429.187
R1008 VDD VDD.n186 429.187
R1009 VDD VDD.n515 426.699
R1010 VDD VDD.n488 426.699
R1011 VDD VDD.n441 426.699
R1012 VDD VDD.n401 426.699
R1013 VDD.n313 VDD 424.618
R1014 VDD VDD.n307 424.618
R1015 VDD VDD.n302 422.557
R1016 VDD.n524 VDD.n523 421.611
R1017 VDD.n53 VDD.t625 420.793
R1018 VDD.n604 VDD.n598 417.5
R1019 VDD.n599 VDD.n598 413.366
R1020 VDD.t558 VDD.t98 387.098
R1021 VDD.t93 VDD.t95 387.098
R1022 VDD.t153 VDD.t152 386.404
R1023 VDD.n201 VDD.t169 386.365
R1024 VDD.n232 VDD.t580 386.365
R1025 VDD.n515 VDD.t495 386.365
R1026 VDD.n488 VDD.t630 386.365
R1027 VDD.n441 VDD.t483 386.365
R1028 VDD.n401 VDD.t567 386.365
R1029 VDD.n313 VDD.t659 386.365
R1030 VDD.n307 VDD.t443 386.365
R1031 VDD.n186 VDD.t392 386.365
R1032 VDD.n169 VDD.t117 386.365
R1033 VDD.t541 VDD.t607 380.952
R1034 VDD.t326 VDD.t667 380.952
R1035 VDD.t83 VDD.t675 380.952
R1036 VDD.t431 VDD.t321 380.952
R1037 VDD.t248 VDD.t681 380.952
R1038 VDD.t126 VDD.t436 380.952
R1039 VDD.t661 VDD.n313 378.788
R1040 VDD.n307 VDD.t313 378.788
R1041 VDD.n302 VDD.t669 378.788
R1042 VDD.t232 VDD.n236 375
R1043 VDD.n233 VDD.n232 368.159
R1044 VDD.t657 VDD.n683 354.539
R1045 VDD.t9 VDD.n730 354.539
R1046 VDD.n62 VDD.t341 351.586
R1047 VDD.n563 VDD.t522 351.586
R1048 VDD.t350 VDD.t352 347.827
R1049 VDD.t356 VDD.t350 347.827
R1050 VDD.t353 VDD.t356 347.827
R1051 VDD.t348 VDD.t353 347.827
R1052 VDD.t354 VDD.t348 347.827
R1053 VDD.t351 VDD.t354 347.827
R1054 VDD.t357 VDD.t351 347.827
R1055 VDD.t355 VDD.t357 347.827
R1056 VDD.t349 VDD.t355 347.827
R1057 VDD.n236 VDD.n234 343.137
R1058 VDD.t26 VDD.n524 306.118
R1059 VDD.t73 VDD.t309 303.031
R1060 VDD.t577 VDD.t457 303.031
R1061 VDD.t239 VDD.t123 303.031
R1062 VDD.t438 VDD.t290 303.031
R1063 VDD.t635 VDD.t323 303.031
R1064 VDD.t140 VDD.t445 303.031
R1065 VDD.t598 VDD.t335 303.031
R1066 VDD.t448 VDD.t268 303.031
R1067 VDD.t604 VDD.t684 303.031
R1068 VDD.t76 VDD.t520 303.031
R1069 VDD.t593 VDD.t67 303.031
R1070 VDD.t113 VDD.t411 303.031
R1071 VDD.t672 VDD.t615 303.031
R1072 VDD.t70 VDD.t366 303.031
R1073 VDD.t678 VDD.t63 303.031
R1074 VDD.t408 VDD.t226 303.031
R1075 VDD.t601 VDD.t333 303.031
R1076 VDD.t401 VDD.t292 303.031
R1077 VDD.n527 VDD.n239 298.536
R1078 VDD.n619 VDD.t19 289.017
R1079 VDD.n730 VDD 288.426
R1080 VDD.n531 VDD.n239 288
R1081 VDD.n683 VDD 285.887
R1082 VDD.n683 VDD.t138 280.245
R1083 VDD.n730 VDD.t556 280.245
R1084 VDD.n619 VDD.t50 265.897
R1085 VDD.n610 VDD.t558 261.649
R1086 VDD.n404 VDD.t664 242.857
R1087 VDD.n406 VDD.t221 242.857
R1088 VDD.t607 VDD.n409 242.857
R1089 VDD.n413 VDD.t326 242.857
R1090 VDD.n443 VDD.t318 242.857
R1091 VDD.n445 VDD.t6 242.857
R1092 VDD.t675 VDD.n448 242.857
R1093 VDD.n452 VDD.t431 242.857
R1094 VDD.n262 VDD.t428 242.857
R1095 VDD.n264 VDD.t284 242.857
R1096 VDD.t681 VDD.n267 242.857
R1097 VDD.n271 VDD.t126 242.857
R1098 VDD.n603 VDD.n602 242.417
R1099 VDD.n7 VDD.t194 232.809
R1100 VDD.n669 VDD.t451 232.809
R1101 VDD.n10 VDD.t145 232.803
R1102 VDD.n672 VDD.t529 232.803
R1103 VDD.t14 VDD.t16 231.214
R1104 VDD.t11 VDD.t14 231.214
R1105 VDD.t19 VDD.t11 231.214
R1106 VDD.t50 VDD.t61 231.214
R1107 VDD.t61 VDD.t55 231.214
R1108 VDD.t55 VDD.t53 231.214
R1109 VDD.n681 VDD.t135 230.548
R1110 VDD.n681 VDD.t277 230.548
R1111 VDD.n15 VDD.t553 230.548
R1112 VDD.n15 VDD.t419 230.548
R1113 VDD.n8 VDD.t467 227.667
R1114 VDD.n9 VDD.t58 227.667
R1115 VDD.n671 VDD.t176 227.667
R1116 VDD.n670 VDD.t89 227.667
R1117 VDD.n611 VDD.t93 213.262
R1118 VDD.n41 VDD.n40 199.562
R1119 VDD.n45 VDD.n44 199.562
R1120 VDD.n192 VDD.t306 193.183
R1121 VDD.n193 VDD.t588 193.183
R1122 VDD.n199 VDD.t387 193.183
R1123 VDD.n200 VDD.t73 193.183
R1124 VDD.n224 VDD.t454 193.183
R1125 VDD.n226 VDD.t160 193.183
R1126 VDD.n228 VDD.t534 193.183
R1127 VDD.n231 VDD.t577 193.183
R1128 VDD.n237 VDD.t232 193.183
R1129 VDD.n497 VDD.t241 193.183
R1130 VDD.n503 VDD.t281 193.183
R1131 VDD.n504 VDD.t463 193.183
R1132 VDD.n514 VDD.t123 193.183
R1133 VDD.n475 VDD.t287 193.183
R1134 VDD.n476 VDD.t3 193.183
R1135 VDD.n486 VDD.t21 193.183
R1136 VDD.n487 VDD.t438 193.183
R1137 VDD.n427 VDD.t632 193.183
R1138 VDD.n433 VDD.t218 193.183
R1139 VDD.n434 VDD.t425 193.183
R1140 VDD.n440 VDD.t323 193.183
R1141 VDD.n388 VDD.t627 193.183
R1142 VDD.n394 VDD.t563 193.183
R1143 VDD.n395 VDD.t213 193.183
R1144 VDD.n400 VDD.t445 193.183
R1145 VDD.n333 VDD.t271 193.183
R1146 VDD.n335 VDD.t560 193.183
R1147 VDD.n338 VDD.t598 193.183
R1148 VDD.n341 VDD.t448 193.183
R1149 VDD.n314 VDD.t661 193.183
R1150 VDD.n312 VDD.t313 193.183
R1151 VDD.n306 VDD.t669 193.183
R1152 VDD.n203 VDD.t517 193.183
R1153 VDD.n205 VDD.t163 193.183
R1154 VDD.n208 VDD.t604 193.183
R1155 VDD.n211 VDD.t76 193.183
R1156 VDD.n173 VDD.t595 193.183
R1157 VDD.n179 VDD.t642 193.183
R1158 VDD.n180 VDD.t103 193.183
R1159 VDD.n185 VDD.t67 193.183
R1160 VDD.n156 VDD.t110 193.183
R1161 VDD.n162 VDD.t499 193.183
R1162 VDD.n163 VDD.t187 193.183
R1163 VDD.n168 VDD.t411 193.183
R1164 VDD.n135 VDD.t361 193.183
R1165 VDD.n137 VDD.t502 193.183
R1166 VDD.n140 VDD.t672 193.183
R1167 VDD.n143 VDD.t70 193.183
R1168 VDD.n107 VDD.t235 193.183
R1169 VDD.n109 VDD.t639 193.183
R1170 VDD.n112 VDD.t678 193.183
R1171 VDD.n115 VDD.t408 193.183
R1172 VDD.n79 VDD.t296 193.183
R1173 VDD.n81 VDD.t585 193.183
R1174 VDD.n84 VDD.t601 193.183
R1175 VDD.n87 VDD.t401 193.183
R1176 VDD.n715 VDD.t142 193.183
R1177 VDD.n25 VDD.t250 193.183
R1178 VDD.n23 VDD.t254 193.183
R1179 VDD.n21 VDD.t260 193.183
R1180 VDD.n690 VDD.t257 193.183
R1181 VDD.n693 VDD.t263 193.183
R1182 VDD.n700 VDD.t531 193.183
R1183 VDD.n575 VDD.t303 193.183
R1184 VDD.n526 VDD.t294 191.288
R1185 VDD.n641 VDD.t48 191.288
R1186 VDD.t655 VDD.t270 175.631
R1187 VDD.t466 VDD.t516 175.631
R1188 VDD.t173 VDD.n660 175.573
R1189 VDD.n40 VDD.t513 170.577
R1190 VDD.n40 VDD.t371 170.577
R1191 VDD.n44 VDD.t610 170.577
R1192 VDD.n44 VDD.t459 170.577
R1193 VDD.t33 VDD.t36 165.977
R1194 VDD.t201 VDD.t383 164.123
R1195 VDD.t497 VDD.n297 153.678
R1196 VDD.t549 VDD.n55 153.678
R1197 VDD.t185 VDD.t173 152.673
R1198 VDD.t294 VDD.t358 151.516
R1199 VDD.n598 VDD.t87 150
R1200 VDD.t179 VDD.t28 146.947
R1201 VDD.n681 VDD.t274 143.345
R1202 VDD.n15 VDD.t416 143.345
R1203 VDD.t339 VDD.n404 138.095
R1204 VDD.t423 VDD.n406 138.095
R1205 VDD.t547 VDD.n409 138.095
R1206 VDD.n413 VDD.t486 138.095
R1207 VDD.t511 VDD.n443 138.095
R1208 VDD.t24 VDD.n445 138.095
R1209 VDD.t373 VDD.n448 138.095
R1210 VDD.n452 VDD.t477 138.095
R1211 VDD.t653 VDD.n262 138.095
R1212 VDD.t461 VDD.n264 138.095
R1213 VDD.t147 VDD.n267 138.095
R1214 VDD.n271 VDD.t474 138.095
R1215 VDD.t199 VDD.t378 137.405
R1216 VDD.n236 VDD.t133 132.353
R1217 VDD.t95 VDD.n610 125.448
R1218 VDD.n247 VDD.t266 124.511
R1219 VDD.t203 VDD.t375 124.046
R1220 VDD.n527 VDD.n526 117.216
R1221 VDD.n234 VDD.n233 112.746
R1222 VDD.n641 VDD.t182 111.743
R1223 VDD.t156 VDD.n192 109.849
R1224 VDD.n193 VDD.t331 109.849
R1225 VDD.t414 VDD.n199 109.849
R1226 VDD.t169 VDD.n200 109.849
R1227 VDD.t79 VDD.n224 109.849
R1228 VDD.t686 VDD.n226 109.849
R1229 VDD.t514 VDD.n228 109.849
R1230 VDD.t580 VDD.n231 109.849
R1231 VDD.n237 VDD.t364 109.849
R1232 VDD.n497 VDD.t611 109.849
R1233 VDD.t246 VDD.n503 109.849
R1234 VDD.n504 VDD.t106 109.849
R1235 VDD.t495 VDD.n514 109.849
R1236 VDD.t131 VDD.n475 109.849
R1237 VDD.n476 VDD.t81 109.849
R1238 VDD.t646 VDD.n486 109.849
R1239 VDD.t630 VDD.n487 109.849
R1240 VDD.n427 VDD.t507 109.849
R1241 VDD.t539 VDD.n433 109.849
R1242 VDD.n434 VDD.t619 109.849
R1243 VDD.t483 VDD.n440 109.849
R1244 VDD.n388 VDD.t545 109.849
R1245 VDD.t337 VDD.n394 109.849
R1246 VDD.n395 VDD.t346 109.849
R1247 VDD.t567 VDD.n400 109.849
R1248 VDD.t149 VDD.n333 109.849
R1249 VDD.t211 VDD.n335 109.849
R1250 VDD.t623 VDD.n338 109.849
R1251 VDD.n341 VDD.t489 109.849
R1252 VDD.n314 VDD.t316 109.849
R1253 VDD.t659 VDD.n312 109.849
R1254 VDD.t443 VDD.n306 109.849
R1255 VDD.t154 VDD.n203 109.849
R1256 VDD.t537 VDD.n205 109.849
R1257 VDD.t42 VDD.n208 109.849
R1258 VDD.n211 VDD.t582 109.849
R1259 VDD.n173 VDD.t119 109.849
R1260 VDD.t65 VDD.n179 109.849
R1261 VDD.n180 VDD.t197 109.849
R1262 VDD.t392 VDD.n185 109.849
R1263 VDD.n156 VDD.t385 109.849
R1264 VDD.t613 VDD.n162 109.849
R1265 VDD.n163 VDD.t192 109.849
R1266 VDD.t117 VDD.n168 109.849
R1267 VDD.t471 VDD.n135 109.849
R1268 VDD.t190 VDD.n137 109.849
R1269 VDD.t551 VDD.n140 109.849
R1270 VDD.n143 VDD.t115 109.849
R1271 VDD.t571 VDD.n107 109.849
R1272 VDD.t101 VDD.n109 109.849
R1273 VDD.t569 VDD.n112 109.849
R1274 VDD.n115 VDD.t394 109.849
R1275 VDD.t216 VDD.n79 109.849
R1276 VDD.t390 VDD.n81 109.849
R1277 VDD.t38 VDD.n84 109.849
R1278 VDD.n87 VDD.t651 109.849
R1279 VDD.n715 VDD.t492 109.849
R1280 VDD.n25 VDD.t469 109.849
R1281 VDD.n23 VDD.t44 109.849
R1282 VDD.n21 VDD.t209 109.849
R1283 VDD.n690 VDD.t244 109.849
R1284 VDD.n693 VDD.t279 109.849
R1285 VDD.n700 VDD.t480 109.849
R1286 VDD.n575 VDD.t91 109.849
R1287 VDD.n598 VDD.n597 99.0104
R1288 VDD.n412 VDD.t541 97.6195
R1289 VDD.n451 VDD.t83 97.6195
R1290 VDD.n270 VDD.t248 97.6195
R1291 VDD.t358 VDD.n246 96.5914
R1292 VDD.n640 VDD.t380 92.5578
R1293 VDD.n684 VDD.t657 92.1507
R1294 VDD.n731 VDD.t9 92.1507
R1295 VDD.n602 VDD.t2 91.7103
R1296 VDD.n525 VDD.n247 90.2261
R1297 VDD.t27 VDD.t645 87.2098
R1298 VDD.t253 VDD.t27 87.2098
R1299 VDD.t151 VDD.t253 87.2098
R1300 VDD.t566 VDD.t151 87.2098
R1301 VDD.t584 VDD.t650 87.2098
R1302 VDD.t650 VDD.t396 87.2098
R1303 VDD.t396 VDD.t168 87.2098
R1304 VDD.t168 VDD.t656 87.2098
R1305 VDD.n60 VDD.t421 80.0005
R1306 VDD.n32 VDD.n31 76.7332
R1307 VDD.n525 VDD.t26 76.2337
R1308 VDD.n661 VDD.t31 73.4738
R1309 VDD.t637 VDD 68.2053
R1310 VDD.n750 VDD.t584 66.4976
R1311 VDD.n53 VDD 65.7064
R1312 VDD.n515 VDD.t129 62.1896
R1313 VDD.n488 VDD.t441 62.1896
R1314 VDD.n441 VDD.t329 62.1896
R1315 VDD.n401 VDD.t434 62.1896
R1316 VDD.n68 VDD.t299 61.9053
R1317 VDD.n313 VDD.t108 61.8817
R1318 VDD.n307 VDD.t617 61.8817
R1319 VDD.n302 VDD.t311 61.5769
R1320 VDD VDD.n233 61.0269
R1321 VDD.n661 VDD.t171 60.115
R1322 VDD.n201 VDD.t404 59.702
R1323 VDD.n232 VDD.t575 59.702
R1324 VDD.n186 VDD.t397 59.702
R1325 VDD.n169 VDD.t406 59.702
R1326 VDD.n524 VDD.t158 59.4064
R1327 VDD.n673 VDD.n672 59.3792
R1328 VDD.n739 VDD.n10 59.3792
R1329 VDD.t206 VDD.n640 58.2066
R1330 VDD.n669 VDD.n668 56.5869
R1331 VDD.n740 VDD.n7 56.5869
R1332 VDD.n298 VDD.t509 55.0852
R1333 VDD.t573 VDD.n301 55.0852
R1334 VDD.n56 VDD.t505 55.0852
R1335 VDD.t543 VDD.n59 55.0852
R1336 VDD.n246 VDD.t230 54.9247
R1337 VDD.n597 VDD.t527 49.5054
R1338 VDD.t171 VDD.t33 32.4432
R1339 VDD.n371 VDD.t488 30.9379
R1340 VDD.n343 VDD.t476 30.9379
R1341 VDD.n570 VDD.t491 30.9379
R1342 VDD.n571 VDD.t479 30.9379
R1343 VDD.n362 VDD.t482 30.7203
R1344 VDD.n349 VDD.t494 30.7203
R1345 VDD.n682 VDD.n681 30.7172
R1346 VDD.n16 VDD.n15 30.7172
R1347 VDD.n367 VDD.t485 30.2877
R1348 VDD.n355 VDD.t473 29.1661
R1349 VDD.t375 VDD.t199 28.6265
R1350 VDD.n33 VDD.n32 28.1049
R1351 VDD.n660 VDD.t383 26.7181
R1352 VDD.n367 VDD.t690 24.9141
R1353 VDD.n371 VDD.t688 24.5101
R1354 VDD.n357 VDD.t695 24.5101
R1355 VDD.n343 VDD.t692 24.5101
R1356 VDD.n349 VDD.t689 24.4814
R1357 VDD.n362 VDD.t693 24.4814
R1358 VDD.n297 VDD.t655 21.9544
R1359 VDD.n55 VDD.t466 21.9544
R1360 VDD.n570 VDD.t691 21.6422
R1361 VDD.n571 VDD.t694 21.6422
R1362 VDD.n750 VDD.t566 20.7127
R1363 VDD.n526 VDD.n525 20.147
R1364 VDD.t31 VDD.t179 19.0845
R1365 VDD.n567 VDD.n566 18.577
R1366 VDD.n719 VDD.n712 17.9105
R1367 VDD.t378 VDD.t206 15.2677
R1368 VDD.n51 VDD.t544 14.0055
R1369 VDD.n54 VDD.t550 13.2223
R1370 VDD.n659 VDD.n589 12.9385
R1371 VDD.n299 VDD.t510 12.3869
R1372 VDD.n57 VDD.t506 12.3869
R1373 VDD.n46 VDD.t638 12.3869
R1374 VDD.n666 VDD.n665 11.1336
R1375 VDD.n638 VDD.n637 10.918
R1376 VDD.n51 VDD.t422 10.1341
R1377 VDD.n529 VDD.n528 9.64171
R1378 VDD.n696 VDD.n695 8.95925
R1379 VDD.t2 VDD.t85 8.90522
R1380 VDD.n357 VDD.n356 8.0005
R1381 VDD.n355 VDD.n354 8.0005
R1382 VDD.n698 VDD.n577 7.3805
R1383 VDD.n523 VDD.n522 7.01458
R1384 VDD.n684 VDD.n682 6.82644
R1385 VDD.n731 VDD.n16 6.82644
R1386 VDD.n530 VDD.n529 6.69176
R1387 VDD.n4 VDD.n3 6.5905
R1388 VDD.n624 VDD.t20 6.5805
R1389 VDD.n633 VDD.t94 6.51327
R1390 VDD.n636 VDD.n607 6.51327
R1391 VDD.n645 VDD.n594 6.45726
R1392 VDD.n657 VDD.t384 6.45726
R1393 VDD.n655 VDD.n651 6.45726
R1394 VDD.n665 VDD.t37 6.45726
R1395 VDD.n572 VDD.t92 6.45146
R1396 VDD.n678 VDD.t278 6.44246
R1397 VDD.n372 VDD.n370 6.39748
R1398 VDD.n602 VDD 6.30798
R1399 VDD.n297 VDD 6.30126
R1400 VDD VDD.n531 6.3005
R1401 VDD.n533 VDD.n239 6.3005
R1402 VDD VDD.n527 6.3005
R1403 VDD.n385 VDD.n333 6.3005
R1404 VDD.n382 VDD.n335 6.3005
R1405 VDD.n379 VDD.n338 6.3005
R1406 VDD.n376 VDD.n341 6.3005
R1407 VDD.n389 VDD.n388 6.3005
R1408 VDD.n394 VDD.n393 6.3005
R1409 VDD.n396 VDD.n395 6.3005
R1410 VDD.n400 VDD.n399 6.3005
R1411 VDD.n423 VDD.n404 6.3005
R1412 VDD.n420 VDD.n406 6.3005
R1413 VDD.n417 VDD.n409 6.3005
R1414 VDD.n414 VDD.n413 6.3005
R1415 VDD.n428 VDD.n427 6.3005
R1416 VDD.n433 VDD.n432 6.3005
R1417 VDD.n435 VDD.n434 6.3005
R1418 VDD VDD.n298 6.3005
R1419 VDD.n301 VDD.n300 6.3005
R1420 VDD.n306 VDD.n305 6.3005
R1421 VDD.n312 VDD.n311 6.3005
R1422 VDD.n315 VDD.n314 6.3005
R1423 VDD.n440 VDD.n439 6.3005
R1424 VDD.n462 VDD.n443 6.3005
R1425 VDD.n459 VDD.n445 6.3005
R1426 VDD.n456 VDD.n448 6.3005
R1427 VDD.n453 VDD.n452 6.3005
R1428 VDD.n475 VDD.n474 6.3005
R1429 VDD.n477 VDD.n476 6.3005
R1430 VDD.n486 VDD.n485 6.3005
R1431 VDD.n487 VDD.n284 6.3005
R1432 VDD.n281 VDD.n262 6.3005
R1433 VDD.n278 VDD.n264 6.3005
R1434 VDD.n275 VDD.n267 6.3005
R1435 VDD.n272 VDD.n271 6.3005
R1436 VDD.n498 VDD.n497 6.3005
R1437 VDD.n503 VDD.n502 6.3005
R1438 VDD.n505 VDD.n504 6.3005
R1439 VDD.n514 VDD.n513 6.3005
R1440 VDD.n536 VDD.n237 6.3005
R1441 VDD VDD.n234 6.3005
R1442 VDD.n212 VDD.n211 6.3005
R1443 VDD.n215 VDD.n208 6.3005
R1444 VDD.n218 VDD.n205 6.3005
R1445 VDD.n221 VDD.n203 6.3005
R1446 VDD.n550 VDD.n224 6.3005
R1447 VDD.n547 VDD.n226 6.3005
R1448 VDD.n544 VDD.n228 6.3005
R1449 VDD.n541 VDD.n231 6.3005
R1450 VDD.n144 VDD.n143 6.3005
R1451 VDD.n147 VDD.n140 6.3005
R1452 VDD.n150 VDD.n137 6.3005
R1453 VDD.n153 VDD.n135 6.3005
R1454 VDD.n157 VDD.n156 6.3005
R1455 VDD.n162 VDD.n161 6.3005
R1456 VDD.n164 VDD.n163 6.3005
R1457 VDD.n168 VDD.n167 6.3005
R1458 VDD.n116 VDD.n115 6.3005
R1459 VDD.n119 VDD.n112 6.3005
R1460 VDD.n122 VDD.n109 6.3005
R1461 VDD.n125 VDD.n107 6.3005
R1462 VDD.n174 VDD.n173 6.3005
R1463 VDD.n179 VDD.n178 6.3005
R1464 VDD.n181 VDD.n180 6.3005
R1465 VDD.n185 VDD.n184 6.3005
R1466 VDD.n88 VDD.n87 6.3005
R1467 VDD.n91 VDD.n84 6.3005
R1468 VDD.n94 VDD.n81 6.3005
R1469 VDD.n97 VDD.n79 6.3005
R1470 VDD.n192 VDD.n191 6.3005
R1471 VDD.n194 VDD.n193 6.3005
R1472 VDD.n199 VDD.n198 6.3005
R1473 VDD.n555 VDD.n200 6.3005
R1474 VDD.n55 VDD.n54 6.3005
R1475 VDD.n59 VDD.n58 6.3005
R1476 VDD VDD.n56 6.3005
R1477 VDD.n69 VDD.n68 6.3005
R1478 VDD.n39 VDD 6.3005
R1479 VDD.n43 VDD 6.3005
R1480 VDD.n30 VDD.n29 6.3005
R1481 VDD.n29 VDD.n28 6.3005
R1482 VDD VDD.n599 6.3005
R1483 VDD VDD.n604 6.3005
R1484 VDD.n576 VDD.n575 6.3005
R1485 VDD.n701 VDD.n700 6.3005
R1486 VDD.n694 VDD.n693 6.3005
R1487 VDD.n691 VDD.n690 6.3005
R1488 VDD.n662 VDD.n661 6.3005
R1489 VDD.n642 VDD.n641 6.3005
R1490 VDD.n637 VDD.n606 6.3005
R1491 VDD VDD.n612 6.3005
R1492 VDD.n634 VDD.n610 6.3005
R1493 VDD.n632 VDD.n611 6.3005
R1494 VDD.n623 VDD.n619 6.3005
R1495 VDD.n22 VDD.n21 6.3005
R1496 VDD.n724 VDD.n23 6.3005
R1497 VDD.n721 VDD.n25 6.3005
R1498 VDD.n717 VDD.n715 6.3005
R1499 VDD.n751 VDD.n750 6.3005
R1500 VDD.n749 VDD.n748 6.11967
R1501 VDD.n61 VDD.t592 5.85907
R1502 VDD.n706 VDD.n705 5.84038
R1503 VDD.n704 VDD.n703 5.78069
R1504 VDD.t28 VDD.t185 5.72569
R1505 VDD.n557 VDD.n556 5.69603
R1506 VDD.n9 VDD.n8 5.60274
R1507 VDD.n671 VDD.n670 5.60274
R1508 VDD.n692 VDD.n580 5.43849
R1509 VDD.n627 VDD.n613 5.41564
R1510 VDD.n621 VDD.n1 5.35178
R1511 VDD.n626 VDD.n625 5.35178
R1512 VDD.n628 VDD.n627 5.35178
R1513 VDD.n745 VDD.n744 5.333
R1514 VDD.n360 VDD.n359 5.30733
R1515 VDD.n688 VDD.t139 5.26584
R1516 VDD VDD.t122 5.22218
R1517 VDD.n22 VDD.t210 5.21805
R1518 VDD.n701 VDD.t481 5.21701
R1519 VDD.n727 VDD.n20 5.21429
R1520 VDD.n414 VDD.t487 5.213
R1521 VDD.n453 VDD.t478 5.213
R1522 VDD.n272 VDD.t475 5.213
R1523 VDD.n212 VDD.t583 5.213
R1524 VDD.n144 VDD.t116 5.213
R1525 VDD.n116 VDD.t395 5.213
R1526 VDD.n88 VDD.t652 5.213
R1527 VDD.n718 VDD.n714 5.20057
R1528 VDD.n699 VDD.n574 5.18056
R1529 VDD.n30 VDD.t302 5.17584
R1530 VDD.n601 VDD.t528 5.17584
R1531 VDD.n600 VDD.t86 5.17584
R1532 VDD.n729 VDD.t557 5.17584
R1533 VDD.n605 VDD.t88 5.17411
R1534 VDD.n436 VDD.t620 5.16792
R1535 VDD.n631 VDD.t649 5.16718
R1536 VDD.n716 VDD.t493 5.16674
R1537 VDD.n535 VDD.t365 5.15377
R1538 VDD.n723 VDD.t45 5.13746
R1539 VDD.n579 VDD.t245 5.13746
R1540 VDD.n695 VDD.t280 5.13746
R1541 VDD.n17 VDD.t420 5.13746
R1542 VDD.n26 VDD.t470 5.13746
R1543 VDD.n667 VDD.n585 5.13586
R1544 VDD.n674 VDD.t90 5.13586
R1545 VDD.n738 VDD.t468 5.13586
R1546 VDD.n741 VDD.n6 5.13586
R1547 VDD.n537 VDD.n235 5.13287
R1548 VDD.n243 VDD.n242 5.13287
R1549 VDD.n244 VDD.t238 5.13287
R1550 VDD.n244 VDD.t231 5.13287
R1551 VDD.n386 VDD.n332 5.13287
R1552 VDD.n384 VDD.t150 5.13287
R1553 VDD.n383 VDD.n334 5.13287
R1554 VDD.n381 VDD.t212 5.13287
R1555 VDD.n378 VDD.t624 5.13287
R1556 VDD.n387 VDD.n331 5.13287
R1557 VDD.n390 VDD.t546 5.13287
R1558 VDD.n391 VDD.n330 5.13287
R1559 VDD.n392 VDD.t338 5.13287
R1560 VDD.n329 VDD.n328 5.13287
R1561 VDD.n397 VDD.t347 5.13287
R1562 VDD.n325 VDD.t568 5.13287
R1563 VDD.n424 VDD.n403 5.13287
R1564 VDD.n422 VDD.t340 5.13287
R1565 VDD.n421 VDD.n405 5.13287
R1566 VDD.n419 VDD.t424 5.13287
R1567 VDD.n416 VDD.t548 5.13287
R1568 VDD.n426 VDD.n324 5.13287
R1569 VDD.n429 VDD.t508 5.13287
R1570 VDD.n430 VDD.n323 5.13287
R1571 VDD.n431 VDD.t540 5.13287
R1572 VDD.n322 VDD.n321 5.13287
R1573 VDD.n318 VDD.t484 5.13287
R1574 VDD.n304 VDD.n294 5.13287
R1575 VDD.n293 VDD.t444 5.13287
R1576 VDD.n309 VDD.n292 5.13287
R1577 VDD.n310 VDD.t660 5.13287
R1578 VDD.n290 VDD.n289 5.13287
R1579 VDD.n316 VDD.t317 5.13287
R1580 VDD.n463 VDD.n442 5.13287
R1581 VDD.n461 VDD.t512 5.13287
R1582 VDD.n460 VDD.n444 5.13287
R1583 VDD.n458 VDD.t25 5.13287
R1584 VDD.n455 VDD.t374 5.13287
R1585 VDD.n288 VDD.n287 5.13287
R1586 VDD.n473 VDD.t132 5.13287
R1587 VDD.n472 VDD.n471 5.13287
R1588 VDD.n478 VDD.t82 5.13287
R1589 VDD.n479 VDD.n285 5.13287
R1590 VDD.n483 VDD.t647 5.13287
R1591 VDD.n490 VDD.t631 5.13287
R1592 VDD.n282 VDD.n261 5.13287
R1593 VDD.n280 VDD.t654 5.13287
R1594 VDD.n279 VDD.n263 5.13287
R1595 VDD.n277 VDD.t462 5.13287
R1596 VDD.n274 VDD.t148 5.13287
R1597 VDD.n496 VDD.n260 5.13287
R1598 VDD.n499 VDD.t612 5.13287
R1599 VDD.n501 VDD.n259 5.13287
R1600 VDD.n257 VDD.t247 5.13287
R1601 VDD.n506 VDD.n258 5.13287
R1602 VDD.n255 VDD.t107 5.13287
R1603 VDD.n252 VDD.t496 5.13287
R1604 VDD.n540 VDD.t581 5.13287
R1605 VDD.n543 VDD.t515 5.13287
R1606 VDD.n545 VDD.n227 5.13287
R1607 VDD.n546 VDD.t687 5.13287
R1608 VDD.n548 VDD.n225 5.13287
R1609 VDD.n549 VDD.t80 5.13287
R1610 VDD.n551 VDD.n223 5.13287
R1611 VDD.n214 VDD.t43 5.13287
R1612 VDD.n217 VDD.t538 5.13287
R1613 VDD.n219 VDD.n204 5.13287
R1614 VDD.n220 VDD.t155 5.13287
R1615 VDD.n222 VDD.n202 5.13287
R1616 VDD.n127 VDD.t118 5.13287
R1617 VDD.n165 VDD.t193 5.13287
R1618 VDD.n131 VDD.n130 5.13287
R1619 VDD.n160 VDD.t614 5.13287
R1620 VDD.n159 VDD.n132 5.13287
R1621 VDD.n158 VDD.t386 5.13287
R1622 VDD.n155 VDD.n133 5.13287
R1623 VDD.n146 VDD.t552 5.13287
R1624 VDD.n149 VDD.t191 5.13287
R1625 VDD.n151 VDD.n136 5.13287
R1626 VDD.n152 VDD.t472 5.13287
R1627 VDD.n154 VDD.n134 5.13287
R1628 VDD.n118 VDD.t570 5.13287
R1629 VDD.n121 VDD.t102 5.13287
R1630 VDD.n123 VDD.n108 5.13287
R1631 VDD.n124 VDD.t572 5.13287
R1632 VDD.n126 VDD.n106 5.13287
R1633 VDD.n99 VDD.t393 5.13287
R1634 VDD.n182 VDD.t198 5.13287
R1635 VDD.n103 VDD.n102 5.13287
R1636 VDD.n177 VDD.t66 5.13287
R1637 VDD.n176 VDD.n104 5.13287
R1638 VDD.n175 VDD.t120 5.13287
R1639 VDD.n172 VDD.n105 5.13287
R1640 VDD.n554 VDD.t170 5.13287
R1641 VDD.n197 VDD.t415 5.13287
R1642 VDD.n196 VDD.n74 5.13287
R1643 VDD.n195 VDD.t332 5.13287
R1644 VDD.n76 VDD.n75 5.13287
R1645 VDD.n190 VDD.t157 5.13287
R1646 VDD.n189 VDD.n77 5.13287
R1647 VDD.n90 VDD.t39 5.13287
R1648 VDD.n93 VDD.t391 5.13287
R1649 VDD.n95 VDD.n80 5.13287
R1650 VDD.n96 VDD.t217 5.13287
R1651 VDD.n98 VDD.n78 5.13287
R1652 VDD.n64 VDD.t225 5.13287
R1653 VDD.n50 VDD.n49 5.13287
R1654 VDD.n67 VDD.t345 5.13287
R1655 VDD.n565 VDD.t229 5.13287
R1656 VDD.n561 VDD.n560 5.13287
R1657 VDD.n19 VDD.n18 5.13287
R1658 VDD.n689 VDD.n581 5.13287
R1659 VDD.n697 VDD.n578 5.13287
R1660 VDD.n583 VDD.n582 5.13287
R1661 VDD.n735 VDD.n12 5.13287
R1662 VDD.n722 VDD.n24 5.13287
R1663 VDD.n675 VDD.t530 5.13129
R1664 VDD.n666 VDD.n586 5.13129
R1665 VDD.n742 VDD.n5 5.13129
R1666 VDD.n737 VDD.t146 5.13129
R1667 VDD.n687 VDD.t658 5.10854
R1668 VDD.n14 VDD.t10 5.10854
R1669 VDD.n677 VDD.n584 5.10445
R1670 VDD.n736 VDD.n11 5.10445
R1671 VDD VDD.t626 5.10424
R1672 VDD.n295 VDD.t574 5.09836
R1673 VDD.n528 VDD.t267 5.09407
R1674 VDD.n530 VDD.t41 5.09407
R1675 VDD.n402 VDD.t435 5.09407
R1676 VDD.n303 VDD.t312 5.09407
R1677 VDD.n308 VDD.t618 5.09407
R1678 VDD.n291 VDD.t109 5.09407
R1679 VDD.n465 VDD.t330 5.09407
R1680 VDD.n489 VDD.t442 5.09407
R1681 VDD.n250 VDD.t130 5.09407
R1682 VDD.n248 VDD.t159 5.09407
R1683 VDD.n538 VDD.t134 5.09407
R1684 VDD.n539 VDD.t576 5.09407
R1685 VDD.n553 VDD.t405 5.09407
R1686 VDD.n170 VDD.t407 5.09407
R1687 VDD.n187 VDD.t398 5.09407
R1688 VDD.n562 VDD.t622 5.09407
R1689 VDD.n38 VDD.t47 5.09407
R1690 VDD.n42 VDD.t167 5.09407
R1691 VDD.n639 VDD.n596 5.09246
R1692 VDD.n643 VDD.t49 5.08866
R1693 VDD.n500 VDD.n256 5.0055
R1694 VDD.n484 VDD.n283 5.0055
R1695 VDD.n517 VDD.n516 5.0005
R1696 VDD.n512 VDD.n251 5.0005
R1697 VDD.n510 VDD.n509 5.0005
R1698 VDD.n468 VDD.n286 4.9955
R1699 VDD.n508 VDD.n507 4.9905
R1700 VDD.n494 VDD.n493 4.9905
R1701 VDD.n470 VDD.n469 4.9905
R1702 VDD.n492 VDD.n491 4.9855
R1703 VDD.n467 VDD.n466 4.9805
R1704 VDD.n70 VDD.t300 4.9655
R1705 VDD.n523 VDD 4.91611
R1706 VDD.n737 VDD.n736 4.88931
R1707 VDD.n375 VDD.t490 4.8755
R1708 VDD.n676 VDD.n675 4.86034
R1709 VDD.n370 VDD.n360 4.84121
R1710 VDD.n519 VDD.n518 4.7947
R1711 VDD.n615 VDD.n614 4.76177
R1712 VDD.n743 VDD.t54 4.7565
R1713 VDD.n622 VDD.n620 4.7565
R1714 VDD.n664 VDD.t172 4.713
R1715 VDD.n656 VDD.n650 4.713
R1716 VDD.n649 VDD.t202 4.713
R1717 VDD.n644 VDD.n595 4.713
R1718 VDD.n698 VDD.n697 4.69819
R1719 VDD.n618 VDD.n617 4.6705
R1720 VDD.n711 VDD.n710 4.56932
R1721 VDD.n350 VDD.n348 4.5005
R1722 VDD.n351 VDD.n348 4.5005
R1723 VDD.n344 VDD.n342 4.5005
R1724 VDD.n345 VDD.n342 4.5005
R1725 VDD.n363 VDD.n361 4.5005
R1726 VDD.n364 VDD.n361 4.5005
R1727 VDD.n520 VDD.n238 4.5005
R1728 VDD.n519 VDD.n249 4.5005
R1729 VDD.n37 VDD.n36 4.5005
R1730 VDD.n36 VDD.n35 4.5005
R1731 VDD.n41 VDD.t372 4.40826
R1732 VDD.n45 VDD.t460 4.3915
R1733 VDD.n696 VDD.n579 4.34898
R1734 VDD.n39 VDD.t46 4.26489
R1735 VDD.n43 VDD.t166 4.26489
R1736 VDD.n729 VDD.n728 4.21364
R1737 VDD.n532 VDD.t1 4.11379
R1738 VDD VDD.n570 4.005
R1739 VDD VDD.n571 4.005
R1740 VDD.n296 VDD.t498 3.94862
R1741 VDD.n171 VDD.n126 3.90405
R1742 VDD.n743 VDD.n742 3.78851
R1743 VDD VDD.n296 3.6765
R1744 VDD.n591 VDD.t379 3.6405
R1745 VDD.n591 VDD.n590 3.6405
R1746 VDD.n588 VDD.t32 3.6405
R1747 VDD.n588 VDD.n587 3.6405
R1748 VDD.n609 VDD.t559 3.6405
R1749 VDD.n609 VDD.n608 3.6405
R1750 VDD.n612 VDD.t648 3.58471
R1751 VDD.n699 VDD.n698 3.24518
R1752 VDD.n246 VDD.n245 3.1505
R1753 VDD.n34 VDD 3.1505
R1754 VDD.n686 VDD.n685 3.1505
R1755 VDD.n685 VDD.n684 3.1505
R1756 VDD.n680 VDD.n679 3.1505
R1757 VDD.n682 VDD.n680 3.1505
R1758 VDD.n659 VDD.n658 3.1505
R1759 VDD.n660 VDD.n659 3.1505
R1760 VDD.n647 VDD.n589 3.1505
R1761 VDD.n640 VDD.n589 3.1505
R1762 VDD.n734 VDD.n13 3.1505
R1763 VDD.n16 VDD.n13 3.1505
R1764 VDD.n733 VDD.n732 3.1505
R1765 VDD.n732 VDD.n731 3.1505
R1766 VDD.n708 VDD.n707 3.13856
R1767 VDD.n639 VDD.n638 2.9013
R1768 VDD.n654 VDD.n653 2.893
R1769 VDD.n646 VDD.n593 2.893
R1770 VDD.n372 VDD.n371 2.88182
R1771 VDD.n358 VDD.n357 2.88074
R1772 VDD.n635 VDD.n609 2.87327
R1773 VDD.n243 VDD.n241 2.85787
R1774 VDD.n380 VDD.n337 2.85787
R1775 VDD.n377 VDD.n340 2.85787
R1776 VDD.n398 VDD.n327 2.85787
R1777 VDD.n418 VDD.n408 2.85787
R1778 VDD.n415 VDD.n411 2.85787
R1779 VDD.n438 VDD.n320 2.85787
R1780 VDD.n457 VDD.n447 2.85787
R1781 VDD.n454 VDD.n450 2.85787
R1782 VDD.n482 VDD.n481 2.85787
R1783 VDD.n276 VDD.n266 2.85787
R1784 VDD.n273 VDD.n269 2.85787
R1785 VDD.n511 VDD.n254 2.85787
R1786 VDD.n542 VDD.n230 2.85787
R1787 VDD.n213 VDD.n210 2.85787
R1788 VDD.n216 VDD.n207 2.85787
R1789 VDD.n166 VDD.n129 2.85787
R1790 VDD.n145 VDD.n142 2.85787
R1791 VDD.n148 VDD.n139 2.85787
R1792 VDD.n117 VDD.n114 2.85787
R1793 VDD.n120 VDD.n111 2.85787
R1794 VDD.n183 VDD.n101 2.85787
R1795 VDD.n73 VDD.n72 2.85787
R1796 VDD.n89 VDD.n86 2.85787
R1797 VDD.n92 VDD.n83 2.85787
R1798 VDD.n65 VDD.n48 2.85787
R1799 VDD.n648 VDD.n591 2.81726
R1800 VDD.n663 VDD.n588 2.81726
R1801 VDD.n728 VDD.n727 2.72534
R1802 VDD.n638 VDD.n605 2.679
R1803 VDD.n518 VDD.n517 2.65128
R1804 VDD.n567 VDD.n37 2.64581
R1805 VDD.n241 VDD.t295 2.2755
R1806 VDD.n241 VDD.n240 2.2755
R1807 VDD.n337 VDD.t336 2.2755
R1808 VDD.n337 VDD.n336 2.2755
R1809 VDD.n340 VDD.t269 2.2755
R1810 VDD.n340 VDD.n339 2.2755
R1811 VDD.n327 VDD.t141 2.2755
R1812 VDD.n327 VDD.n326 2.2755
R1813 VDD.n408 VDD.t542 2.2755
R1814 VDD.n408 VDD.n407 2.2755
R1815 VDD.n411 VDD.t668 2.2755
R1816 VDD.n411 VDD.n410 2.2755
R1817 VDD.n320 VDD.t636 2.2755
R1818 VDD.n320 VDD.n319 2.2755
R1819 VDD.n447 VDD.t84 2.2755
R1820 VDD.n447 VDD.n446 2.2755
R1821 VDD.n450 VDD.t322 2.2755
R1822 VDD.n450 VDD.n449 2.2755
R1823 VDD.n481 VDD.t291 2.2755
R1824 VDD.n481 VDD.n480 2.2755
R1825 VDD.n266 VDD.t249 2.2755
R1826 VDD.n266 VDD.n265 2.2755
R1827 VDD.n269 VDD.t437 2.2755
R1828 VDD.n269 VDD.n268 2.2755
R1829 VDD.n254 VDD.t240 2.2755
R1830 VDD.n254 VDD.n253 2.2755
R1831 VDD.n230 VDD.t458 2.2755
R1832 VDD.n230 VDD.n229 2.2755
R1833 VDD.n210 VDD.t521 2.2755
R1834 VDD.n210 VDD.n209 2.2755
R1835 VDD.n207 VDD.t685 2.2755
R1836 VDD.n207 VDD.n206 2.2755
R1837 VDD.n129 VDD.t114 2.2755
R1838 VDD.n129 VDD.n128 2.2755
R1839 VDD.n142 VDD.t367 2.2755
R1840 VDD.n142 VDD.n141 2.2755
R1841 VDD.n139 VDD.t616 2.2755
R1842 VDD.n139 VDD.n138 2.2755
R1843 VDD.n114 VDD.t227 2.2755
R1844 VDD.n114 VDD.n113 2.2755
R1845 VDD.n111 VDD.t64 2.2755
R1846 VDD.n111 VDD.n110 2.2755
R1847 VDD.n101 VDD.t594 2.2755
R1848 VDD.n101 VDD.n100 2.2755
R1849 VDD.n72 VDD.t310 2.2755
R1850 VDD.n72 VDD.n71 2.2755
R1851 VDD.n86 VDD.t293 2.2755
R1852 VDD.n86 VDD.n85 2.2755
R1853 VDD.n83 VDD.t334 2.2755
R1854 VDD.n83 VDD.n82 2.2755
R1855 VDD.n48 VDD.t400 2.2755
R1856 VDD.n48 VDD.n47 2.2755
R1857 VDD.n540 VDD 2.25904
R1858 VDD.n709 VDD.n708 2.2505
R1859 VDD.n748 VDD.n747 2.2505
R1860 VDD.n353 VDD.n352 2.2439
R1861 VDD.n366 VDD.n365 2.2439
R1862 VDD.n347 VDD.n346 2.24362
R1863 VDD.n344 VDD.n343 2.12277
R1864 VDD.t380 VDD.t201 1.9089
R1865 VDD.n368 VDD.n367 1.82213
R1866 VDD.n3 VDD.t62 1.8205
R1867 VDD.n3 VDD.n2 1.8205
R1868 VDD.n617 VDD.t15 1.8205
R1869 VDD.n617 VDD.n616 1.8205
R1870 VDD.n653 VDD.t186 1.8205
R1871 VDD.n653 VDD.n652 1.8205
R1872 VDD.n593 VDD.t200 1.8205
R1873 VDD.n593 VDD.n592 1.8205
R1874 VDD VDD.n325 1.81785
R1875 VDD.n357 VDD.n355 1.77234
R1876 VDD.n749 VDD 1.6722
R1877 VDD.n36 VDD.n34 1.67038
R1878 VDD.n359 VDD.n353 1.6239
R1879 VDD.n369 VDD.n366 1.6239
R1880 VDD.n678 VDD.n583 1.5845
R1881 VDD.n521 VDD.n520 1.50339
R1882 VDD.n363 VDD.n362 1.39846
R1883 VDD.n350 VDD.n349 1.39728
R1884 VDD.n728 VDD.n19 1.39383
R1885 VDD.n708 VDD.n569 1.20737
R1886 VDD.n387 VDD.n386 1.16167
R1887 VDD.n359 VDD.n358 1.12314
R1888 VDD.n369 VDD.n368 1.12224
R1889 VDD.n425 VDD.n424 1.07428
R1890 VDD.n552 VDD.n222 1.02928
R1891 VDD.n188 VDD.n98 1.02928
R1892 VDD.n464 VDD.n463 1.01882
R1893 VDD.n495 VDD.n282 1.01882
R1894 VDD.n676 VDD.n583 0.920186
R1895 VDD.n155 VDD.n154 0.881662
R1896 VDD.n631 VDD.n630 0.829892
R1897 VDD VDD.n67 0.819742
R1898 VDD.n247 VDD.t0 0.783764
R1899 VDD.n751 VDD.n749 0.754
R1900 VDD.n573 VDD.n572 0.7205
R1901 VDD.n559 VDD.n38 0.66512
R1902 VDD.n718 VDD.n713 0.636929
R1903 VDD.n558 VDD.n42 0.634017
R1904 VDD VDD.n17 0.57316
R1905 VDD.n705 VDD 0.56151
R1906 VDD.n706 VDD 0.550028
R1907 VDD.n370 VDD.n369 0.52356
R1908 VDD.n629 VDD.n615 0.500134
R1909 VDD.n360 VDD.n347 0.497812
R1910 VDD.n747 VDD 0.445652
R1911 VDD VDD.n745 0.372092
R1912 VDD.n376 VDD.n375 0.337997
R1913 VDD.n703 VDD.n702 0.336214
R1914 VDD.n375 VDD.n374 0.333658
R1915 VDD VDD.n557 0.281196
R1916 VDD.n695 VDD.n694 0.257375
R1917 VDD.n437 VDD.n317 0.25039
R1918 VDD.n689 VDD.n688 0.245004
R1919 VDD.n697 VDD.n696 0.238698
R1920 VDD.n381 VDD.n380 0.233919
R1921 VDD.n378 VDD.n377 0.233919
R1922 VDD.n419 VDD.n418 0.233919
R1923 VDD.n416 VDD.n415 0.233919
R1924 VDD.n458 VDD.n457 0.233919
R1925 VDD.n455 VDD.n454 0.233919
R1926 VDD.n277 VDD.n276 0.233919
R1927 VDD.n274 VDD.n273 0.233919
R1928 VDD.n217 VDD.n216 0.233919
R1929 VDD.n214 VDD.n213 0.233919
R1930 VDD.n149 VDD.n148 0.233919
R1931 VDD.n146 VDD.n145 0.233919
R1932 VDD.n121 VDD.n120 0.233919
R1933 VDD.n118 VDD.n117 0.233919
R1934 VDD.n93 VDD.n92 0.233919
R1935 VDD.n90 VDD.n89 0.233919
R1936 VDD.n534 VDD.n533 0.224447
R1937 VDD.n539 VDD 0.205357
R1938 VDD.n566 VDD.n565 0.203989
R1939 VDD.n535 VDD.n534 0.202146
R1940 VDD.n492 VDD.n283 0.201676
R1941 VDD.n748 VDD.n0 0.201567
R1942 VDD.n467 VDD.n317 0.200832
R1943 VDD.n634 VDD.n633 0.196412
R1944 VDD.n468 VDD.n283 0.183147
R1945 VDD.n518 VDD.n250 0.182938
R1946 VDD.n469 VDD.n467 0.1805
R1947 VDD.n469 VDD.n468 0.177853
R1948 VDD.n720 VDD.n711 0.171929
R1949 VDD.n562 VDD.n561 0.170231
R1950 VDD.n553 VDD.n552 0.167533
R1951 VDD.n493 VDD.n256 0.167265
R1952 VDD VDD.n296 0.16613
R1953 VDD.n493 VDD.n492 0.161971
R1954 VDD VDD.n99 0.160716
R1955 VDD.n554 VDD 0.158984
R1956 VDD VDD.n127 0.157289
R1957 VDD.n188 VDD.n187 0.155496
R1958 VDD.n632 VDD 0.154644
R1959 VDD.n171 VDD.n170 0.154581
R1960 VDD.n508 VDD.n256 0.151382
R1961 VDD.n703 VDD 0.15032
R1962 VDD.n723 VDD.n722 0.149994
R1963 VDD VDD.n52 0.149922
R1964 VDD.n688 VDD.n687 0.149577
R1965 VDD.n509 VDD.n251 0.148735
R1966 VDD.n509 VDD.n508 0.146088
R1967 VDD.n426 VDD.n425 0.144547
R1968 VDD.n559 VDD.n558 0.142342
R1969 VDD.n384 VDD.n383 0.141016
R1970 VDD.n391 VDD.n390 0.141016
R1971 VDD.n392 VDD.n329 0.141016
R1972 VDD.n422 VDD.n421 0.141016
R1973 VDD.n430 VDD.n429 0.141016
R1974 VDD.n431 VDD.n322 0.141016
R1975 VDD.n461 VDD.n460 0.141016
R1976 VDD.n280 VDD.n279 0.141016
R1977 VDD.n220 VDD.n219 0.141016
R1978 VDD.n152 VDD.n151 0.141016
R1979 VDD.n124 VDD.n123 0.141016
R1980 VDD.n96 VDD.n95 0.141016
R1981 VDD.n425 VDD.n402 0.138896
R1982 VDD.n685 VDD.n680 0.138205
R1983 VDD.n732 VDD.n13 0.138205
R1984 VDD.n172 VDD.n171 0.131861
R1985 VDD.n538 VDD.n537 0.130567
R1986 VDD.n744 VDD.n4 0.128315
R1987 VDD.n549 VDD.n548 0.123551
R1988 VDD.n546 VDD.n545 0.123551
R1989 VDD.n176 VDD.n175 0.123551
R1990 VDD.n177 VDD.n103 0.123551
R1991 VDD.n703 VDD.n573 0.122835
R1992 VDD VDD.n397 0.122435
R1993 VDD.n517 VDD.n251 0.122265
R1994 VDD.n190 VDD.n76 0.122176
R1995 VDD.n196 VDD.n195 0.122176
R1996 VDD.n747 VDD.n746 0.121062
R1997 VDD.n159 VDD.n158 0.120831
R1998 VDD.n160 VDD.n131 0.120831
R1999 VDD.n625 VDD.n618 0.119239
R2000 VDD.n10 VDD.n9 0.117546
R2001 VDD.n672 VDD.n671 0.117546
R2002 VDD.n710 VDD 0.117041
R2003 VDD.n552 VDD.n551 0.116432
R2004 VDD.n636 VDD 0.115362
R2005 VDD.n189 VDD.n188 0.115137
R2006 VDD.n398 VDD 0.111984
R2007 VDD.n8 VDD.n7 0.111412
R2008 VDD.n670 VDD.n669 0.111412
R2009 VDD.n368 VDD 0.110941
R2010 VDD VDD.n52 0.107354
R2011 VDD.n386 VDD.n385 0.107339
R2012 VDD.n383 VDD.n382 0.107339
R2013 VDD.n389 VDD.n387 0.107339
R2014 VDD.n393 VDD.n391 0.107339
R2015 VDD.n396 VDD.n329 0.107339
R2016 VDD.n424 VDD.n423 0.107339
R2017 VDD.n421 VDD.n420 0.107339
R2018 VDD.n428 VDD.n426 0.107339
R2019 VDD.n432 VDD.n430 0.107339
R2020 VDD.n435 VDD.n322 0.107339
R2021 VDD.n463 VDD.n462 0.107339
R2022 VDD.n460 VDD.n459 0.107339
R2023 VDD.n282 VDD.n281 0.107339
R2024 VDD.n279 VDD.n278 0.107339
R2025 VDD.n537 VDD.n536 0.107339
R2026 VDD.n222 VDD.n221 0.107339
R2027 VDD.n219 VDD.n218 0.107339
R2028 VDD.n154 VDD.n153 0.107339
R2029 VDD.n151 VDD.n150 0.107339
R2030 VDD.n126 VDD.n125 0.107339
R2031 VDD.n123 VDD.n122 0.107339
R2032 VDD.n98 VDD.n97 0.107339
R2033 VDD.n95 VDD.n94 0.107339
R2034 VDD.n564 VDD.n561 0.107339
R2035 VDD.n543 VDD 0.10728
R2036 VDD VDD.n182 0.10728
R2037 VDD.n380 VDD 0.106177
R2038 VDD.n377 VDD 0.106177
R2039 VDD VDD.n398 0.106177
R2040 VDD.n418 VDD 0.106177
R2041 VDD.n415 VDD 0.106177
R2042 VDD.n457 VDD 0.106177
R2043 VDD.n454 VDD 0.106177
R2044 VDD.n276 VDD 0.106177
R2045 VDD.n273 VDD 0.106177
R2046 VDD.n216 VDD 0.106177
R2047 VDD.n213 VDD 0.106177
R2048 VDD.n148 VDD 0.106177
R2049 VDD.n145 VDD 0.106177
R2050 VDD.n120 VDD 0.106177
R2051 VDD.n117 VDD 0.106177
R2052 VDD.n92 VDD 0.106177
R2053 VDD.n89 VDD 0.106177
R2054 VDD.n197 VDD 0.106087
R2055 VDD VDD.n165 0.10492
R2056 VDD VDD.n635 0.100445
R2057 VDD.n626 VDD.n1 0.0999848
R2058 VDD VDD.n542 0.0981271
R2059 VDD.n183 VDD 0.0981271
R2060 VDD.n637 VDD.n636 0.0974613
R2061 VDD VDD.n73 0.0970363
R2062 VDD.n559 VDD.n41 0.096125
R2063 VDD.n166 VDD 0.0959696
R2064 VDD.n61 VDD 0.0956733
R2065 VDD.n551 VDD.n550 0.0940593
R2066 VDD.n548 VDD.n547 0.0940593
R2067 VDD.n545 VDD.n544 0.0940593
R2068 VDD.n174 VDD.n172 0.0940593
R2069 VDD.n178 VDD.n176 0.0940593
R2070 VDD.n181 VDD.n103 0.0940593
R2071 VDD.n542 VDD 0.0930424
R2072 VDD VDD.n183 0.0930424
R2073 VDD.n191 VDD.n189 0.093014
R2074 VDD.n194 VDD.n76 0.093014
R2075 VDD.n198 VDD.n196 0.093014
R2076 VDD.n157 VDD.n155 0.0919917
R2077 VDD.n161 VDD.n159 0.0919917
R2078 VDD.n164 VDD.n131 0.0919917
R2079 VDD VDD.n166 0.0909972
R2080 VDD.n558 VDD.n45 0.0905
R2081 VDD.n720 VDD.n719 0.0905
R2082 VDD.n629 VDD.n628 0.0897437
R2083 VDD.n709 VDD.n27 0.0869056
R2084 VDD VDD.n293 0.084523
R2085 VDD.n310 VDD 0.084523
R2086 VDD VDD.n295 0.0842767
R2087 VDD.n356 VDD 0.0839415
R2088 VDD.n678 VDD.n677 0.0835769
R2089 VDD.n718 VDD 0.0830688
R2090 VDD.n569 VDD.n568 0.0828897
R2091 VDD.n317 VDD.n316 0.0826283
R2092 VDD.n566 VDD 0.0823094
R2093 VDD.n534 VDD.n238 0.0819374
R2094 VDD.n622 VDD.n621 0.0818025
R2095 VDD.n65 VDD.n64 0.0817097
R2096 VDD.n351 VDD 0.0816915
R2097 VDD.n516 VDD.n252 0.0816286
R2098 VDD.n379 VDD.n378 0.080629
R2099 VDD.n399 VDD.n325 0.080629
R2100 VDD.n417 VDD.n416 0.080629
R2101 VDD.n456 VDD.n455 0.080629
R2102 VDD.n275 VDD.n274 0.080629
R2103 VDD.n215 VDD.n214 0.080629
R2104 VDD.n147 VDD.n146 0.080629
R2105 VDD.n119 VDD.n118 0.080629
R2106 VDD.n91 VDD.n90 0.080629
R2107 VDD.n364 VDD 0.0805665
R2108 VDD.n717 VDD.n716 0.079766
R2109 VDD VDD.n384 0.0794677
R2110 VDD VDD.n381 0.0794677
R2111 VDD.n390 VDD 0.0794677
R2112 VDD VDD.n392 0.0794677
R2113 VDD.n397 VDD 0.0794677
R2114 VDD VDD.n422 0.0794677
R2115 VDD VDD.n419 0.0794677
R2116 VDD.n429 VDD 0.0794677
R2117 VDD VDD.n431 0.0794677
R2118 VDD VDD.n461 0.0794677
R2119 VDD VDD.n458 0.0794677
R2120 VDD VDD.n280 0.0794677
R2121 VDD VDD.n277 0.0794677
R2122 VDD VDD.n220 0.0794677
R2123 VDD VDD.n217 0.0794677
R2124 VDD VDD.n152 0.0794677
R2125 VDD VDD.n149 0.0794677
R2126 VDD VDD.n124 0.0794677
R2127 VDD VDD.n121 0.0794677
R2128 VDD VDD.n96 0.0794677
R2129 VDD VDD.n93 0.0794677
R2130 VDD.n745 VDD.n1 0.0789075
R2131 VDD.n735 VDD 0.0786463
R2132 VDD.n436 VDD 0.0765085
R2133 VDD.n565 VDD 0.0759839
R2134 VDD.n345 VDD 0.0738165
R2135 VDD.n374 VDD.n372 0.0725
R2136 VDD.n577 VDD 0.0721766
R2137 VDD.n665 VDD.n664 0.0716397
R2138 VDD.n528 VDD 0.0709717
R2139 VDD.n402 VDD 0.0709717
R2140 VDD.n248 VDD 0.0709717
R2141 VDD VDD.n539 0.0709717
R2142 VDD VDD.n562 0.0709717
R2143 VDD VDD.n38 0.0709717
R2144 VDD VDD.n42 0.0709717
R2145 VDD.n541 VDD.n540 0.0706695
R2146 VDD.n184 VDD.n99 0.0706695
R2147 VDD.n722 VDD 0.0699068
R2148 VDD.n555 VDD.n554 0.0698855
R2149 VDD VDD.n549 0.0696525
R2150 VDD VDD.n546 0.0696525
R2151 VDD VDD.n543 0.0696525
R2152 VDD.n175 VDD 0.0696525
R2153 VDD VDD.n177 0.0696525
R2154 VDD.n182 VDD 0.0696525
R2155 VDD.n167 VDD.n127 0.0691188
R2156 VDD.n627 VDD.n626 0.0690012
R2157 VDD VDD.n190 0.0688799
R2158 VDD.n195 VDD 0.0688799
R2159 VDD VDD.n197 0.0688799
R2160 VDD.n158 VDD 0.0681243
R2161 VDD VDD.n160 0.0681243
R2162 VDD.n165 VDD 0.0681243
R2163 VDD.n373 VDD 0.0659545
R2164 VDD.n646 VDD.n645 0.0653529
R2165 VDD.n473 VDD.n472 0.0647478
R2166 VDD.n479 VDD.n478 0.0647478
R2167 VDD.n687 VDD.n686 0.0618846
R2168 VDD.n304 VDD.n303 0.0618169
R2169 VDD.n309 VDD.n308 0.0618169
R2170 VDD.n291 VDD.n290 0.0618169
R2171 VDD.n725 VDD.n19 0.0612407
R2172 VDD.n615 VDD.n613 0.0612211
R2173 VDD.n643 VDD 0.0610515
R2174 VDD.n464 VDD.n288 0.0607039
R2175 VDD.n496 VDD.n495 0.0607039
R2176 VDD.n300 VDD.n299 0.0599607
R2177 VDD.n507 VDD.n506 0.0597035
R2178 VDD.n733 VDD.n14 0.0588902
R2179 VDD.n501 VDD.n500 0.0586416
R2180 VDD.n702 VDD 0.0585645
R2181 VDD.n649 VDD.n648 0.0574118
R2182 VDD.n654 VDD 0.0570809
R2183 VDD.n483 VDD 0.0562522
R2184 VDD VDD.n51 0.0559424
R2185 VDD VDD.n532 0.0555633
R2186 VDD VDD.n535 0.0550806
R2187 VDD.n465 VDD.n464 0.0536232
R2188 VDD.n655 VDD.n654 0.0534412
R2189 VDD VDD.n243 0.0533387
R2190 VDD.n556 VDD.n73 0.0532933
R2191 VDD.n656 VDD.n655 0.0531103
R2192 VDD VDD.n510 0.0522699
R2193 VDD.n299 VDD 0.0518708
R2194 VDD.n624 VDD 0.0515504
R2195 VDD.n438 VDD 0.0514734
R2196 VDD VDD.n482 0.0514734
R2197 VDD.n511 VDD 0.0514734
R2198 VDD.n724 VDD.n723 0.0512407
R2199 VDD.n485 VDD.n479 0.0493496
R2200 VDD.n498 VDD.n496 0.0493496
R2201 VDD.n502 VDD.n501 0.0493496
R2202 VDD.n506 VDD.n505 0.0493496
R2203 VDD VDD.n438 0.0488186
R2204 VDD.n474 VDD.n470 0.0488186
R2205 VDD.n482 VDD 0.0488186
R2206 VDD.n305 VDD.n304 0.0487799
R2207 VDD.n311 VDD.n309 0.0487799
R2208 VDD.n315 VDD.n290 0.0487799
R2209 VDD.n710 VDD.n26 0.0481695
R2210 VDD.n466 VDD.n318 0.046557
R2211 VDD.n642 VDD.n639 0.0461618
R2212 VDD.n605 VDD 0.0456836
R2213 VDD.n374 VDD.n373 0.0455
R2214 VDD.n664 VDD.n663 0.0455
R2215 VDD VDD.n646 0.0451691
R2216 VDD.n58 VDD.n57 0.0446736
R2217 VDD VDD.n50 0.0444695
R2218 VDD.n512 VDD.n511 0.0437743
R2219 VDD VDD.n538 0.043431
R2220 VDD VDD.n631 0.0432624
R2221 VDD.n645 VDD.n644 0.0411985
R2222 VDD.n623 VDD.n622 0.0409622
R2223 VDD.n668 VDD.n667 0.040956
R2224 VDD.n741 VDD.n740 0.040956
R2225 VDD.n674 VDD.n673 0.0406629
R2226 VDD.n739 VDD.n738 0.0406629
R2227 VDD.n187 VDD 0.0404465
R2228 VDD VDD.n553 0.0400238
R2229 VDD.n170 VDD 0.0396099
R2230 VDD.n466 VDD 0.0394398
R2231 VDD.n576 VDD.n573 0.0393024
R2232 VDD.n556 VDD 0.0392151
R2233 VDD.n489 VDD 0.039182
R2234 VDD.n57 VDD 0.0386636
R2235 VDD.n692 VDD.n689 0.0383228
R2236 VDD VDD.n244 0.0382419
R2237 VDD VDD.n649 0.0382206
R2238 VDD VDD.n709 0.0380335
R2239 VDD.n716 VDD.n713 0.0379096
R2240 VDD.n490 VDD 0.0377891
R2241 VDD.n644 VDD.n643 0.0372279
R2242 VDD.n437 VDD.n436 0.0371957
R2243 VDD.n439 VDD.n318 0.0371372
R2244 VDD.n513 VDD.n252 0.0371372
R2245 VDD VDD.n473 0.0366062
R2246 VDD.n478 VDD 0.0366062
R2247 VDD.n499 VDD 0.0366062
R2248 VDD VDD.n257 0.0366062
R2249 VDD VDD.n255 0.0366062
R2250 VDD VDD.n692 0.036125
R2251 VDD VDD.n295 0.0350843
R2252 VDD VDD.n293 0.0346108
R2253 VDD VDD.n310 0.0346108
R2254 VDD.n316 VDD 0.0346108
R2255 VDD.n529 VDD.n243 0.0344677
R2256 VDD VDD.n27 0.0341842
R2257 VDD.n37 VDD.n30 0.0341842
R2258 VDD.n522 VDD.n248 0.0327642
R2259 VDD VDD.n530 0.032019
R2260 VDD.n69 VDD.n46 0.0319625
R2261 VDD.n691 VDD.n579 0.0317152
R2262 VDD.n677 VDD.n676 0.0309615
R2263 VDD.n472 VDD.n286 0.0291726
R2264 VDD.n720 VDD.n26 0.0291017
R2265 VDD.n34 VDD.n33 0.028942
R2266 VDD VDD.n729 0.0284422
R2267 VDD VDD.n46 0.0276819
R2268 VDD.n352 VDD.n351 0.0275
R2269 VDD.n356 VDD.n354 0.0275
R2270 VDD.n484 VDD.n483 0.0265177
R2271 VDD.n365 VDD.n364 0.026375
R2272 VDD.n63 VDD.n50 0.0257824
R2273 VDD.n353 VDD.n348 0.025705
R2274 VDD.n366 VDD.n361 0.025705
R2275 VDD VDD.n65 0.0256227
R2276 VDD.n721 VDD.n720 0.0241441
R2277 VDD.n491 VDD.n284 0.0233319
R2278 VDD.n705 VDD.n704 0.023
R2279 VDD.n249 VDD.n238 0.0225755
R2280 VDD VDD.n465 0.021904
R2281 VDD VDD.n489 0.021904
R2282 VDD VDD.n250 0.021904
R2283 VDD.n303 VDD 0.0216615
R2284 VDD.n308 VDD 0.0216615
R2285 VDD VDD.n291 0.0216615
R2286 VDD VDD.n437 0.0214735
R2287 VDD.n346 VDD.n345 0.02075
R2288 VDD.n477 VDD.n286 0.020677
R2289 VDD.n744 VDD.n743 0.0201639
R2290 VDD.n707 VDD.n706 0.0200181
R2291 VDD.n67 VDD.n66 0.0195491
R2292 VDD.n520 VDD.n519 0.0193811
R2293 VDD.n70 VDD 0.0184587
R2294 VDD.n635 VDD.n634 0.0184006
R2295 VDD.n64 VDD 0.0183626
R2296 VDD.n347 VDD.n342 0.0169383
R2297 VDD VDD.n601 0.0163291
R2298 VDD.n657 VDD.n656 0.0157206
R2299 VDD.n727 VDD.n726 0.0151468
R2300 VDD.n558 VDD 0.0147612
R2301 VDD.n491 VDD.n490 0.0143053
R2302 VDD VDD.n657 0.0140662
R2303 VDD.n557 VDD.n70 0.0137976
R2304 VDD.n621 VDD.n4 0.0133571
R2305 VDD VDD.n52 0.0127264
R2306 VDD.n495 VDD.n494 0.0126203
R2307 VDD.n37 VDD 0.0120789
R2308 VDD VDD.n484 0.0105885
R2309 VDD.n726 VDD 0.00991177
R2310 VDD.n346 VDD.n344 0.0095
R2311 VDD.n630 VDD.n629 0.00881933
R2312 VDD.n373 VDD 0.00868182
R2313 VDD.n704 VDD 0.00844118
R2314 VDD.n713 VDD.n712 0.00809036
R2315 VDD.n725 VDD 0.00716667
R2316 VDD.n658 VDD 0.00711765
R2317 VDD.n707 VDD 0.00700602
R2318 VDD.n500 VDD.n499 0.00660619
R2319 VDD VDD.n559 0.00608887
R2320 VDD.n633 VDD.n632 0.00596961
R2321 VDD.n507 VDD.n257 0.00554425
R2322 VDD VDD.n512 0.00554425
R2323 VDD.n532 VDD 0.00543671
R2324 VDD.n712 VDD.n711 0.00537952
R2325 VDD.n536 VDD 0.00514516
R2326 VDD VDD.n564 0.00514516
R2327 VDD.n688 VDD 0.00489024
R2328 VDD VDD.n51 0.00485726
R2329 VDD.n628 VDD.n618 0.00465966
R2330 VDD.n625 VDD.n624 0.00465966
R2331 VDD.n510 VDD.n255 0.0044823
R2332 VDD.n516 VDD 0.00436819
R2333 VDD.n694 VDD 0.00425
R2334 VDD.n692 VDD 0.00414557
R2335 VDD.n365 VDD.n363 0.003875
R2336 VDD.n719 VDD.n718 0.00371429
R2337 VDD.n648 VDD.n647 0.00347794
R2338 VDD.n663 VDD.n662 0.00347794
R2339 VDD.n533 VDD 0.00315823
R2340 VDD.n675 VDD.n674 0.00284528
R2341 VDD.n738 VDD.n737 0.00284528
R2342 VDD.n245 VDD 0.00282258
R2343 VDD.n494 VDD 0.00282092
R2344 VDD.n352 VDD.n350 0.00275
R2345 VDD.n305 VDD 0.00259913
R2346 VDD.n311 VDD 0.00259913
R2347 VDD VDD.n315 0.00259913
R2348 VDD.n667 VDD.n666 0.00255212
R2349 VDD.n742 VDD.n741 0.00255212
R2350 VDD.n726 VDD.n725 0.00241489
R2351 VDD.n736 VDD.n735 0.0022561
R2352 VDD.n17 VDD.n14 0.0022561
R2353 VDD VDD.n717 0.00215138
R2354 VDD VDD.n623 0.00201261
R2355 VDD.n600 VDD 0.00185678
R2356 VDD.n647 VDD 0.00182353
R2357 VDD.n658 VDD 0.00182353
R2358 VDD.n662 VDD 0.00182353
R2359 VDD.n358 VDD.n354 0.00171994
R2360 VDD VDD.n22 0.00167647
R2361 VDD.n385 VDD 0.00166129
R2362 VDD.n382 VDD 0.00166129
R2363 VDD VDD.n379 0.00166129
R2364 VDD VDD.n376 0.00166129
R2365 VDD VDD.n389 0.00166129
R2366 VDD.n393 VDD 0.00166129
R2367 VDD VDD.n396 0.00166129
R2368 VDD.n399 VDD 0.00166129
R2369 VDD.n423 VDD 0.00166129
R2370 VDD.n420 VDD 0.00166129
R2371 VDD VDD.n417 0.00166129
R2372 VDD VDD.n414 0.00166129
R2373 VDD VDD.n428 0.00166129
R2374 VDD.n432 VDD 0.00166129
R2375 VDD VDD.n435 0.00166129
R2376 VDD.n462 VDD 0.00166129
R2377 VDD.n459 VDD 0.00166129
R2378 VDD VDD.n456 0.00166129
R2379 VDD VDD.n453 0.00166129
R2380 VDD.n281 VDD 0.00166129
R2381 VDD.n278 VDD 0.00166129
R2382 VDD VDD.n275 0.00166129
R2383 VDD VDD.n272 0.00166129
R2384 VDD.n221 VDD 0.00166129
R2385 VDD.n218 VDD 0.00166129
R2386 VDD VDD.n215 0.00166129
R2387 VDD VDD.n212 0.00166129
R2388 VDD.n153 VDD 0.00166129
R2389 VDD.n150 VDD 0.00166129
R2390 VDD VDD.n147 0.00166129
R2391 VDD VDD.n144 0.00166129
R2392 VDD.n125 VDD 0.00166129
R2393 VDD.n122 VDD 0.00166129
R2394 VDD VDD.n119 0.00166129
R2395 VDD VDD.n116 0.00166129
R2396 VDD.n97 VDD 0.00166129
R2397 VDD.n94 VDD 0.00166129
R2398 VDD VDD.n91 0.00166129
R2399 VDD VDD.n88 0.00166129
R2400 VDD VDD.n701 0.00166129
R2401 VDD VDD.n63 0.00159924
R2402 VDD VDD.n576 0.00157784
R2403 VDD.n522 VDD.n521 0.00156548
R2404 VDD.n550 VDD 0.00151695
R2405 VDD.n547 VDD 0.00151695
R2406 VDD.n544 VDD 0.00151695
R2407 VDD VDD.n541 0.00151695
R2408 VDD VDD.n174 0.00151695
R2409 VDD.n178 VDD 0.00151695
R2410 VDD VDD.n181 0.00151695
R2411 VDD.n184 VDD 0.00151695
R2412 VDD.n191 VDD 0.00150559
R2413 VDD VDD.n194 0.00150559
R2414 VDD.n198 VDD 0.00150559
R2415 VDD VDD.n555 0.00150559
R2416 VDD VDD.n751 0.0015
R2417 VDD VDD.n157 0.00149448
R2418 VDD.n161 VDD 0.00149448
R2419 VDD VDD.n164 0.00149448
R2420 VDD.n167 VDD 0.00149448
R2421 VDD VDD.n678 0.00142308
R2422 VDD.n679 VDD 0.00142308
R2423 VDD.n679 VDD 0.00142308
R2424 VDD.n686 VDD 0.00142308
R2425 VDD VDD.n734 0.00137805
R2426 VDD.n734 VDD 0.00137805
R2427 VDD VDD.n733 0.00137805
R2428 VDD.n521 VDD.n249 0.00128347
R2429 VDD VDD.n721 0.00126271
R2430 VDD VDD.n724 0.00124074
R2431 VDD.n568 VDD.n567 0.00116176
R2432 VDD.n673 VDD 0.00108632
R2433 VDD VDD.n739 0.00108632
R2434 VDD.n245 VDD 0.00108064
R2435 VDD.n702 VDD.n699 0.00106301
R2436 VDD.n439 VDD 0.00103097
R2437 VDD.n470 VDD.n288 0.00103097
R2438 VDD.n474 VDD 0.00103097
R2439 VDD VDD.n477 0.00103097
R2440 VDD.n485 VDD 0.00103097
R2441 VDD VDD.n284 0.00103097
R2442 VDD VDD.n498 0.00103097
R2443 VDD.n502 VDD 0.00103097
R2444 VDD.n505 VDD 0.00103097
R2445 VDD.n513 VDD 0.00103097
R2446 VDD.n54 VDD 0.00100943
R2447 VDD.n630 VDD.n613 0.000997238
R2448 VDD VDD.n691 0.000955696
R2449 VDD.n300 VDD 0.000904494
R2450 VDD VDD.n642 0.000830882
R2451 VDD.n569 VDD.n0 0.000830882
R2452 VDD.n58 VDD 0.000800501
R2453 VDD.n668 VDD 0.00079316
R2454 VDD.n740 VDD 0.00079316
R2455 VDD.n66 VDD 0.000776074
R2456 VDD VDD.n61 0.000774809
R2457 VDD.n601 VDD.n600 0.000726131
R2458 VDD VDD.n69 0.000714031
R2459 VSS.n1755 VSS.n1754 1.24442e+07
R2460 VSS.n277 VSS.t241 2.77509e+06
R2461 VSS.n1100 VSS.n1098 326625
R2462 VSS.n278 VSS.n277 291662
R2463 VSS.n1150 VSS.t516 69136.7
R2464 VSS.t335 VSS.n579 68883.1
R2465 VSS.n1432 VSS.n1431 51936
R2466 VSS.n278 VSS.n275 46337.6
R2467 VSS.n561 VSS.n560 32848.9
R2468 VSS.n1101 VSS.n1100 32388.1
R2469 VSS.n1100 VSS.n1099 27173.2
R2470 VSS.t275 VSS.n847 17548.9
R2471 VSS.t80 VSS.n2154 17230
R2472 VSS.t564 VSS.t50 16169.8
R2473 VSS.n275 VSS.n274 15482
R2474 VSS.n2366 VSS.t271 15334.5
R2475 VSS.n279 VSS.n278 14833.1
R2476 VSS.n1154 VSS.n1153 12018.1
R2477 VSS.n126 VSS.t454 10467.5
R2478 VSS.n2369 VSS.n2368 10113
R2479 VSS.n1432 VSS.n1430 9805.53
R2480 VSS.n2216 VSS.n2215 9589.42
R2481 VSS.n106 VSS.n105 9415.54
R2482 VSS.n2369 VSS.n2 9049.5
R2483 VSS.n1429 VSS.n1428 8817.76
R2484 VSS.n2276 VSS.n2275 7059.24
R2485 VSS.n51 VSS.t502 7006.49
R2486 VSS.n856 VSS.n855 6477.06
R2487 VSS.n2270 VSS.n2 6109.02
R2488 VSS.n559 VSS.n557 5720.33
R2489 VSS.n49 VSS.n8 5573.78
R2490 VSS.n180 VSS.n179 5552.94
R2491 VSS.n2365 VSS.n2364 5437.96
R2492 VSS.n1079 VSS.n1078 5431.91
R2493 VSS.t363 VSS.n1101 5106.06
R2494 VSS.n1118 VSS.n1117 5047.28
R2495 VSS.n388 VSS.t177 4775.5
R2496 VSS.n2363 VSS.n8 4690.81
R2497 VSS.n2364 VSS.n2363 4646.68
R2498 VSS.n2162 VSS.n2161 4516.79
R2499 VSS.n2236 VSS.n2183 3893.61
R2500 VSS.n1117 VSS.n1116 3620.01
R2501 VSS.n1120 VSS.n1119 3526.41
R2502 VSS.n1150 VSS.n1149 3506.18
R2503 VSS.n1152 VSS.n1151 3502.33
R2504 VSS.n2293 VSS.n2292 3472.05
R2505 VSS.n1430 VSS.n1429 3339.89
R2506 VSS.n92 VSS.n91 3262.63
R2507 VSS.n562 VSS.n561 3238.68
R2508 VSS.n1428 VSS.n1427 3205.07
R2509 VSS.n2195 VSS.t482 3112.87
R2510 VSS.n91 VSS.n90 3004.05
R2511 VSS.n2368 VSS.n2367 2891.55
R2512 VSS.n2150 VSS.n2149 2682.86
R2513 VSS.n126 VSS.n125 2588.5
R2514 VSS.n2296 VSS.n2295 2416.67
R2515 VSS.t135 VSS.t624 2307.56
R2516 VSS.t77 VSS.t110 2307.56
R2517 VSS.t571 VSS.t169 2307.56
R2518 VSS.t315 VSS.t347 2307.56
R2519 VSS.t294 VSS.t358 2307.56
R2520 VSS.t484 VSS.t345 2307.56
R2521 VSS.t602 VSS.t213 2307.56
R2522 VSS.t214 VSS.t129 2307.56
R2523 VSS.t488 VSS.t237 2307.56
R2524 VSS.t367 VSS.t526 2307.56
R2525 VSS.t470 VSS.t311 2307.56
R2526 VSS.t144 VSS.t3 2307.56
R2527 VSS.t16 VSS.t89 2307.56
R2528 VSS.t281 VSS.t625 2307.56
R2529 VSS.t87 VSS.t173 2307.56
R2530 VSS.t667 VSS.t523 2307.56
R2531 VSS.t496 VSS.t447 2307.56
R2532 VSS.t599 VSS.t278 2307.56
R2533 VSS.t451 VSS.t254 2307.56
R2534 VSS.t113 VSS.t250 2307.56
R2535 VSS.n2297 VSS.n2296 2213.34
R2536 VSS.n125 VSS.t535 2166.67
R2537 VSS.n50 VSS.n49 2138.2
R2538 VSS.n1093 VSS.n1091 2111.77
R2539 VSS.n1420 VSS.n1419 2052.63
R2540 VSS.n2287 VSS.t450 2050.53
R2541 VSS.n1811 VSS.n1810 2050.44
R2542 VSS.n2276 VSS.t559 1984.24
R2543 VSS.t556 VSS.n2184 1878.69
R2544 VSS.n2257 VSS.t155 1862.04
R2545 VSS.n1058 VSS.n1057 1819.72
R2546 VSS.n1433 VSS.n1432 1782.85
R2547 VSS.t46 VSS.n588 1739.89
R2548 VSS.n105 VSS.t598 1731.96
R2549 VSS.t619 VSS.n2216 1713.53
R2550 VSS.t280 VSS.n2237 1713.53
R2551 VSS.t251 VSS.n2299 1713.53
R2552 VSS.n561 VSS.n559 1637.58
R2553 VSS.n131 VSS.t575 1635.55
R2554 VSS.n2237 VSS.n2236 1565.03
R2555 VSS.n576 VSS.n575 1524.83
R2556 VSS.n2312 VSS.t141 1439.29
R2557 VSS.n181 VSS.n180 1425.15
R2558 VSS.n51 VSS.n50 1310.77
R2559 VSS.n53 VSS.t561 1272.1
R2560 VSS.n105 VSS.n92 1249.34
R2561 VSS.n2157 VSS.t353 1199.47
R2562 VSS.n66 VSS.t131 1199.47
R2563 VSS.n2311 VSS.t478 1199.47
R2564 VSS.n1079 VSS.t266 1166.91
R2565 VSS.n2367 VSS.n2366 1156.81
R2566 VSS.t293 VSS.n2162 1153.78
R2567 VSS.t130 VSS.n8 1153.78
R2568 VSS.n2365 VSS.t638 1150.77
R2569 VSS.t621 VSS.n2148 1143.48
R2570 VSS.n128 VSS.n127 1139.06
R2571 VSS.t509 VSS.t507 1132.9
R2572 VSS.t507 VSS.t511 1132.9
R2573 VSS.n373 VSS.n372 1127.25
R2574 VSS.n2289 VSS.n2288 1119.51
R2575 VSS.n575 VSS.n572 1115.8
R2576 VSS.t361 VSS.n1079 1113.16
R2577 VSS.n2363 VSS.t327 1093.68
R2578 VSS.t201 VSS.n576 1093.54
R2579 VSS.n947 VSS.t260 1075.7
R2580 VSS.n4 VSS.n3 1062.21
R2581 VSS.t243 VSS.t563 1058.09
R2582 VSS.n373 VSS.n371 988.177
R2583 VSS.n1102 VSS.t363 968.703
R2584 VSS.t138 VSS.n1093 963.861
R2585 VSS.t96 VSS.n1058 955.883
R2586 VSS.t162 VSS.t485 952.793
R2587 VSS.t614 VSS.t328 952.793
R2588 VSS.n109 VSS.t616 927.716
R2589 VSS.t82 VSS.t577 913.885
R2590 VSS.t85 VSS.t294 913.885
R2591 VSS.t129 VSS.t558 913.885
R2592 VSS.t310 VSS.t620 913.885
R2593 VSS.t437 VSS.t281 913.885
R2594 VSS.t447 VSS.t560 913.885
R2595 VSS.t250 VSS.t143 913.885
R2596 VSS.n2299 VSS.n2298 902.461
R2597 VSS.n1149 VSS.n1148 870.861
R2598 VSS.n1153 VSS.n1152 868.078
R2599 VSS.n1151 VSS.t229 857.508
R2600 VSS.n2298 VSS.n2297 839.713
R2601 VSS.n2214 VSS.t605 838.187
R2602 VSS.n126 VSS.n106 791.109
R2603 VSS.t157 VSS.n1076 765.686
R2604 VSS.n2297 VSS.n2257 756.466
R2605 VSS.n1116 VSS.t138 750.745
R2606 VSS.n2156 VSS.t80 730.073
R2607 VSS.n1091 VSS.n1090 707.154
R2608 VSS.n1076 VSS.n1075 690.782
R2609 VSS.n585 VSS.t343 688.312
R2610 VSS.n2183 VSS.t355 680.952
R2611 VSS.n2194 VSS.t638 671.942
R2612 VSS.n1812 VSS.n1811 666.105
R2613 VSS.n366 VSS.t283 663.793
R2614 VSS.n2292 VSS.n2291 650.433
R2615 VSS.t236 VSS.t554 635.715
R2616 VSS.t651 VSS.t552 635.715
R2617 VSS.n2270 VSS.t564 631.266
R2618 VSS.t457 VSS.t150 623.288
R2619 VSS.n1707 VSS.n1706 602.758
R2620 VSS.t284 VSS.n2147 595.653
R2621 VSS.n127 VSS.t324 578.554
R2622 VSS.n579 VSS.t62 567.638
R2623 VSS.n2161 VSS.t313 564.287
R2624 VSS.n372 VSS.t448 555.885
R2625 VSS.t598 VSS.n104 548.331
R2626 VSS.t624 VSS.n103 548.331
R2627 VSS.t110 VSS.n102 548.331
R2628 VSS.n97 VSS.t82 548.331
R2629 VSS.n2165 VSS.t293 548.331
R2630 VSS.n2166 VSS.t571 548.331
R2631 VSS.n2171 VSS.t347 548.331
R2632 VSS.n2172 VSS.t85 548.331
R2633 VSS.n56 VSS.t130 548.331
R2634 VSS.n57 VSS.t484 548.331
R2635 VSS.n65 VSS.t558 548.331
R2636 VSS.n2217 VSS.t619 548.331
R2637 VSS.n2222 VSS.t237 548.331
R2638 VSS.n2223 VSS.t367 548.331
R2639 VSS.n2226 VSS.t310 548.331
R2640 VSS.n2238 VSS.t280 548.331
R2641 VSS.n2243 VSS.t3 548.331
R2642 VSS.n2244 VSS.t16 548.331
R2643 VSS.n2247 VSS.t437 548.331
R2644 VSS.t450 VSS.n2286 548.331
R2645 VSS.t173 VSS.n2285 548.331
R2646 VSS.t523 VSS.n2284 548.331
R2647 VSS.t560 VSS.n2283 548.331
R2648 VSS.n2300 VSS.t251 548.331
R2649 VSS.n2305 VSS.t278 548.331
R2650 VSS.n2306 VSS.t451 548.331
R2651 VSS.n2310 VSS.t143 548.331
R2652 VSS.n2291 VSS.n2290 545.501
R2653 VSS.t9 VSS.t11 519.481
R2654 VSS.t504 VSS.n562 495.966
R2655 VSS.n848 VSS.t153 491.512
R2656 VSS.t482 VSS.n2194 479.959
R2657 VSS.n81 VSS.t480 470.426
R2658 VSS.t14 VSS.t340 457.793
R2659 VSS.t636 VSS.t498 457.144
R2660 VSS.n2288 VSS.n2287 453.219
R2661 VSS.t63 VSS.n585 451.3
R2662 VSS.n2216 VSS.n6 451.231
R2663 VSS.n2257 VSS.t440 445.519
R2664 VSS.t74 VSS.t38 431.818
R2665 VSS.n1708 VSS.n1707 431.416
R2666 VSS.n92 VSS.n66 426.769
R2667 VSS.t2 VSS.t234 405.356
R2668 VSS.t348 VSS.t91 405.356
R2669 VSS.t314 VSS.t48 405.356
R2670 VSS.n347 VSS.t330 404.658
R2671 VSS.t6 VSS.n580 399.351
R2672 VSS.t443 VSS.t295 398.623
R2673 VSS.t322 VSS.n2150 396.058
R2674 VSS.n5 VSS.n4 383.952
R2675 VSS.t439 VSS.t314 381.512
R2676 VSS.t442 VSS.t140 380.952
R2677 VSS.t559 VSS.t500 380.952
R2678 VSS.n90 VSS.t653 373.81
R2679 VSS.t654 VSS.t318 370.132
R2680 VSS.n104 VSS.t135 365.555
R2681 VSS.n103 VSS.t77 365.555
R2682 VSS.n102 VSS.t217 365.555
R2683 VSS.n97 VSS.t353 365.555
R2684 VSS.t169 VSS.n2165 365.555
R2685 VSS.n2166 VSS.t315 365.555
R2686 VSS.t358 VSS.n2171 365.555
R2687 VSS.n2172 VSS.t189 365.555
R2688 VSS.t345 VSS.n56 365.555
R2689 VSS.n57 VSS.t602 365.555
R2690 VSS.n60 VSS.t214 365.555
R2691 VSS.t131 VSS.n65 365.555
R2692 VSS.n2217 VSS.t488 365.555
R2693 VSS.t526 VSS.n2222 365.555
R2694 VSS.n2223 VSS.t607 365.555
R2695 VSS.n2226 VSS.t470 365.555
R2696 VSS.n2238 VSS.t144 365.555
R2697 VSS.t89 VSS.n2243 365.555
R2698 VSS.n2247 VSS.t155 365.555
R2699 VSS.n2286 VSS.t87 365.555
R2700 VSS.n2285 VSS.t667 365.555
R2701 VSS.n2284 VSS.t496 365.555
R2702 VSS.n2283 VSS.t566 365.555
R2703 VSS.n2300 VSS.t599 365.555
R2704 VSS.t254 VSS.n2305 365.555
R2705 VSS.n2306 VSS.t113 365.555
R2706 VSS.t478 VSS.n2310 365.555
R2707 VSS.n570 VSS.t148 353.382
R2708 VSS.n127 VSS.n126 345.394
R2709 VSS.t43 VSS.t66 340.909
R2710 VSS.t76 VSS.t528 326.19
R2711 VSS.t249 VSS.t651 326.19
R2712 VSS.t246 VSS.t146 312.255
R2713 VSS.n559 VSS.n558 309.524
R2714 VSS.n106 VSS.n51 297.363
R2715 VSS.n2295 VSS.n2294 287.072
R2716 VSS.n589 VSS.t71 282.469
R2717 VSS.n48 VSS.t365 281.091
R2718 VSS.n857 VSS.n854 275.611
R2719 VSS.n570 VSS.t457 269.906
R2720 VSS.n346 VSS.t578 269.688
R2721 VSS.n1710 VSS.n1709 269.413
R2722 VSS.t62 VSS.n577 267.123
R2723 VSS.t506 VSS.t510 262.361
R2724 VSS.n361 VSS.t501 255.748
R2725 VSS.t238 VSS.t512 245.964
R2726 VSS.n563 VSS.t505 241.044
R2727 VSS.t158 VSS.n1147 240.087
R2728 VSS.n1192 VSS.n1191 239.475
R2729 VSS.n2185 VSS.t443 231.852
R2730 VSS.n952 VSS.t545 230.024
R2731 VSS.n34 VSS.t286 228.907
R2732 VSS.n37 VSS.t2 228.907
R2733 VSS.n36 VSS.t572 228.907
R2734 VSS.n41 VSS.t595 228.907
R2735 VSS.n46 VSS.t357 228.907
R2736 VSS.t313 VSS.n2160 228.796
R2737 VSS.t653 VSS.n89 228.571
R2738 VSS.n84 VSS.t236 228.571
R2739 VSS.n27 VSS.t594 228.571
R2740 VSS.n2229 VSS.t307 228.571
R2741 VSS.t498 VSS.n2176 228.571
R2742 VSS.n2258 VSS.t279 228.571
R2743 VSS.n2177 VSS.t174 228.571
R2744 VSS.n2180 VSS.t655 228.571
R2745 VSS.n2272 VSS.t596 228.571
R2746 VSS.t140 VSS.n2181 228.571
R2747 VSS.n948 VSS.n947 226.314
R2748 VSS.n1084 VSS.t264 225.036
R2749 VSS.n568 VSS.t515 225.013
R2750 VSS.t66 VSS.t46 224.026
R2751 VSS.n1209 VSS.t287 218.702
R2752 VSS.t269 VSS.n2362 217.304
R2753 VSS.t543 VSS.n10 217.304
R2754 VSS.n15 VSS.t656 217.304
R2755 VSS.n20 VSS.t436 217.304
R2756 VSS.n997 VSS.t103 215.216
R2757 VSS.t308 VSS.t127 211.208
R2758 VSS.n2364 VSS.n5 206.661
R2759 VSS.n2295 VSS.t175 202.679
R2760 VSS.n1077 VSS.t517 197.663
R2761 VSS.n1081 VSS.t541 197.663
R2762 VSS.n2215 VSS.n2184 195.244
R2763 VSS.t448 VSS.n346 192.633
R2764 VSS.t332 VSS.n2151 186.381
R2765 VSS.t224 VSS.t221 186.113
R2766 VSS.n1709 VSS.n1708 185.804
R2767 VSS.t267 VSS.t0 184.518
R2768 VSS.n348 VSS.t246 181.619
R2769 VSS.t71 VSS.t43 178.571
R2770 VSS.n577 VSS.t201 178.083
R2771 VSS.t563 VSS.n2152 176.673
R2772 VSS.t317 VSS.t597 176.45
R2773 VSS.t282 VSS.t439 176.45
R2774 VSS.t320 VSS.n23 173.81
R2775 VSS.n706 VSS.n705 172.927
R2776 VSS.n997 VSS.t92 171.69
R2777 VSS.n1294 VSS.t518 167.84
R2778 VSS.t438 VSS.n2293 166.667
R2779 VSS.n90 VSS.n83 164.286
R2780 VSS.t247 VSS.n276 163.793
R2781 VSS.n1146 VSS.t468 159.215
R2782 VSS.n988 VSS.t95 154.762
R2783 VSS.n2160 VSS.t492 152.606
R2784 VSS.t234 VSS.n34 152.606
R2785 VSS.n37 VSS.t17 152.606
R2786 VSS.n36 VSS.t348 152.606
R2787 VSS.n42 VSS.t333 152.606
R2788 VSS.t48 VSS.n41 152.606
R2789 VSS.n2250 VSS.t472 152.606
R2790 VSS.t175 VSS.n46 152.606
R2791 VSS.t554 VSS.n23 152.381
R2792 VSS.n24 VSS.t111 152.381
R2793 VSS.t552 VSS.n26 152.381
R2794 VSS.t355 VSS.n31 152.381
R2795 VSS.n2262 VSS.t636 152.381
R2796 VSS.t167 VSS.n2176 152.381
R2797 VSS.n2258 VSS.t452 152.381
R2798 VSS.n2177 VSS.t524 152.381
R2799 VSS.n2180 VSS.t160 152.381
R2800 VSS.n2272 VSS.t52 152.381
R2801 VSS.t466 VSS.n2181 152.381
R2802 VSS.n2195 VSS.t490 150.845
R2803 VSS.n2198 VSS.t556 150.845
R2804 VSS.n1085 VSS.t252 149.236
R2805 VSS.n2364 VSS.n6 142.794
R2806 VSS.n1161 VSS.t276 141.113
R2807 VSS.t37 VSS.t504 141.019
R2808 VSS.n2188 VSS.t464 140.889
R2809 VSS.n11 VSS.t211 140.889
R2810 VSS.n16 VSS.t537 140.889
R2811 VSS.t133 VSS.n80 140.889
R2812 VSS.t94 VSS.n1653 140.849
R2813 VSS.n1127 VSS.t108 140.446
R2814 VSS.n437 VSS.n436 134.505
R2815 VSS.n1162 VSS.t265 134.499
R2816 VSS.n2152 VSS.t332 133.962
R2817 VSS.t41 VSS.t74 133.118
R2818 VSS.n696 VSS.t289 132.238
R2819 VSS.n1074 VSS.t68 131.083
R2820 VSS.n1080 VSS.t273 131.083
R2821 VSS.t633 VSS.n571 130.78
R2822 VSS.n2153 VSS.t243 124.254
R2823 VSS.n2151 VSS.t322 124.254
R2824 VSS.t279 VSS.t167 123.811
R2825 VSS.t524 VSS.t256 123.811
R2826 VSS.t52 VSS.t442 123.811
R2827 VSS.n2213 VSS.t308 122.846
R2828 VSS.t512 VSS.t37 121.343
R2829 VSS.n2236 VSS.n2235 119.948
R2830 VSS.t233 VSS.t434 113.144
R2831 VSS.t548 VSS.n565 113.144
R2832 VSS.n774 VSS.n773 112.609
R2833 VSS.t153 VSS.t275 110.341
R2834 VSS.t343 VSS.t14 107.144
R2835 VSS.n1000 VSS.t101 106.4
R2836 VSS.n1413 VSS.n1412 105.803
R2837 VSS.n580 VSS.t338 103.897
R2838 VSS.n589 VSS.t41 103.897
R2839 VSS.t515 VSS.t548 102.752
R2840 VSS.n243 VSS.n242 99.4576
R2841 VSS.n2154 VSS.t324 99.0148
R2842 VSS.n1119 VSS.n1118 98.0801
R2843 VSS.n89 VSS.t245 97.6195
R2844 VSS.n84 VSS.t623 97.6195
R2845 VSS.n27 VSS.t657 97.6195
R2846 VSS.n2229 VSS.t79 97.6195
R2847 VSS.n1435 VSS.t460 95.3545
R2848 VSS.t171 VSS.n2369 94.4338
R2849 VSS.n397 VSS.t630 93.7031
R2850 VSS.n218 VSS.t664 93.7031
R2851 VSS.n879 VSS.t292 89.9735
R2852 VSS.t330 VSS.t60 89.2162
R2853 VSS.t38 VSS.t63 87.6628
R2854 VSS.n2154 VSS.n2153 87.3661
R2855 VSS.n1176 VSS.t446 81.0285
R2856 VSS.t221 VSS.n1753 79.0986
R2857 VSS.n1162 VSS.n1161 77.1715
R2858 VSS.n493 VSS.n492 76.2916
R2859 VSS.t160 VSS.t666 76.191
R2860 VSS.t500 VSS.t466 76.191
R2861 VSS.t216 VSS.n1433 75.3151
R2862 VSS.n374 VSS.n373 73.2848
R2863 VSS.n1319 VSS.n1318 73.1516
R2864 VSS.n1174 VSS.t106 71.0388
R2865 VSS.t106 VSS.n1173 71.0388
R2866 VSS.n1155 VSS.n1154 70.2233
R2867 VSS.n1175 VSS.n1174 68.8188
R2868 VSS.n1075 VSS.t152 64.9263
R2869 VSS.n1057 VSS.t513 63.726
R2870 VSS.n1059 VSS.t96 63.726
R2871 VSS.n994 VSS.t100 62.8725
R2872 VSS.n2293 VSS.n2262 61.9053
R2873 VSS.t340 VSS.t6 61.6888
R2874 VSS.n198 VSS.n197 60.5636
R2875 VSS.n972 VSS.t198 59.3241
R2876 VSS.t539 VSS.t4 59.0031
R2877 VSS.n83 VSS.n82 57.1434
R2878 VSS.t245 VSS.t320 54.7624
R2879 VSS.t623 VSS.t368 54.7624
R2880 VSS.t594 VSS.t76 54.7624
R2881 VSS.t657 VSS.t533 54.7624
R2882 VSS.t307 VSS.t249 54.7624
R2883 VSS.t79 VSS.t476 54.7624
R2884 VSS.n42 VSS.t317 52.4583
R2885 VSS.n2250 VSS.t282 52.4583
R2886 VSS.n427 VSS.t573 51.6126
R2887 VSS.n1666 VSS.t123 51.5878
R2888 VSS.t263 VSS.n1439 49.63
R2889 VSS.n1711 VSS.n1710 49.5445
R2890 VSS.n175 VSS.t570 48.4151
R2891 VSS.n1439 VSS.n1437 48.2204
R2892 VSS.n2149 VSS.t621 47.8266
R2893 VSS.n2148 VSS.t284 47.8266
R2894 VSS.n1811 VSS.n1809 47.1019
R2895 VSS.n2021 VSS.n2020 46.8512
R2896 VSS.n182 VSS.n181 46.7394
R2897 VSS.n1954 VSS.n1953 46.1999
R2898 VSS.n991 VSS.t104 45.9454
R2899 VSS.n2376 VSS.t19 45.8147
R2900 VSS.t105 VSS.t94 45.4352
R2901 VSS.n783 VSS.t574 45.3566
R2902 VSS.n1593 VSS.t159 45.3348
R2903 VSS.n307 VSS.t297 45.1394
R2904 VSS.n1857 VSS.t530 44.9166
R2905 VSS.n2380 VSS.t499 44.8088
R2906 VSS.n2135 VSS.n2134 44.7339
R2907 VSS.n66 VSS.n53 41.0359
R2908 VSS.t54 VSS.n1441 40.9633
R2909 VSS.n1441 VSS.t262 40.8071
R2910 VSS.n7 VSS.t445 40.409
R2911 VSS.n165 VSS.n164 39.3991
R2912 VSS.n1860 VSS.t35 37.8583
R2913 VSS.t446 VSS.n1175 37.7396
R2914 VSS.n2312 VSS.n2311 37.1434
R2915 VSS.n928 VSS.t206 36.0599
R2916 VSS.n502 VSS.t521 35.603
R2917 VSS.n389 VSS.n388 35.0237
R2918 VSS.n424 VSS.t121 34.4086
R2919 VSS.n1669 VSS.t351 34.392
R2920 VSS.n2235 VSS.t311 34.2711
R2921 VSS.t440 VSS.n2256 34.2711
R2922 VSS.t0 VSS.n2376 32.7249
R2923 VSS.n185 VSS.t609 31.5986
R2924 VSS.n2277 VSS.n2276 30.9563
R2925 VSS.n1863 VSS.t33 30.8001
R2926 VSS.t219 VSS.n1712 30.4891
R2927 VSS.n2380 VSS.t239 29.8727
R2928 VSS.n400 VSS.t662 29.5908
R2929 VSS.n215 VSS.t627 29.5908
R2930 VSS.t11 VSS.t335 29.2213
R2931 VSS.n156 VSS.t102 28.6811
R2932 VSS.n786 VSS.t258 28.1526
R2933 VSS.n1590 VSS.t36 28.139
R2934 VSS.n2294 VSS.t438 25.9531
R2935 VSS.n532 VSS.n531 25.5911
R2936 VSS.t445 VSS.t233 25.4001
R2937 VSS.n572 VSS.t633 25.0433
R2938 VSS.t191 VSS.n279 25.0252
R2939 VSS.n188 VSS.t618 24.3574
R2940 VSS.n857 VSS.n856 24.2542
R2941 VSS.n1866 VSS.t32 23.7419
R2942 VSS.n2157 VSS.n2156 23.5512
R2943 VSS.n795 VSS.t193 23.4606
R2944 VSS.n1581 VSS.t164 23.4493
R2945 VSS.n2290 VSS.t83 22.8476
R2946 VSS.n978 VSS.t195 22.1014
R2947 VSS.n925 VSS.n924 22.1014
R2948 VSS.n1427 VSS.n1426 22.1014
R2949 VSS.n2215 VSS.n2214 21.6311
R2950 VSS.n563 VSS.t508 21.3174
R2951 VSS.n565 VSS.t506 21.3174
R2952 VSS.n245 VSS.n244 21.1752
R2953 VSS.n292 VSS.t25 20.5182
R2954 VSS.n1318 VSS.n1317 20.3448
R2955 VSS.n1756 VSS.n1755 20.3365
R2956 VSS.t501 VSS.t326 20.1154
R2957 VSS.t241 VSS.t247 20.1154
R2958 VSS.n569 VSS.t509 19.8143
R2959 VSS.n1050 VSS.t98 19.3457
R2960 VSS.n1813 VSS.n1812 18.6512
R2961 VSS.n975 VSS.t204 18.6118
R2962 VSS.n267 VSS.t531 18.6086
R2963 VSS.n1749 VSS.t227 18.209
R2964 VSS.n1723 VSS.t219 17.3621
R2965 VSS.n1766 VSS.t27 17.3238
R2966 VSS.n366 VSS.t612 17.2419
R2967 VSS.n421 VSS.t542 17.2045
R2968 VSS.n1876 VSS.t547 17.2045
R2969 VSS.n1672 VSS.t350 17.1963
R2970 VSS.n1677 VSS.t352 17.1963
R2971 VSS.n191 VSS.t583 17.1162
R2972 VSS.n1977 VSS.t34 16.6836
R2973 VSS.t177 VSS.n387 16.5119
R2974 VSS.t508 VSS.t238 16.3981
R2975 VSS.n82 VSS.n81 16.3322
R2976 VSS.n2215 VSS.n2185 16.2708
R2977 VSS.t338 VSS.t9 16.2343
R2978 VSS.n1654 VSS.t105 14.4828
R2979 VSS.n2010 VSS.t185 14.4161
R2980 VSS.n1434 VSS.t216 14.1297
R2981 VSS.n1436 VSS.t360 14.1258
R2982 VSS.n1442 VSS.t263 14.0965
R2983 VSS.t262 VSS.n1440 14.092
R2984 VSS.n2021 VSS.t179 13.6953
R2985 VSS.n2138 VSS.t569 13.656
R2986 VSS.n182 VSS.n178 13.1664
R2987 VSS.n178 VSS.t117 13.1543
R2988 VSS.t360 VSS.n1435 12.9487
R2989 VSS.t327 VSS.t269 11.9402
R2990 VSS.t464 VSS.t162 11.9402
R2991 VSS.t485 VSS.t543 11.9402
R2992 VSS.t211 VSS.t231 11.9402
R2993 VSS.t318 VSS.t601 11.9402
R2994 VSS.t656 VSS.t654 11.9402
R2995 VSS.t537 VSS.t614 11.9402
R2996 VSS.t328 VSS.t270 11.9402
R2997 VSS.t436 VSS.t86 11.9402
R2998 VSS.t480 VSS.t133 11.9402
R2999 VSS.n1964 VSS.t635 11.5504
R3000 VSS.n2459 VSS.n2383 11.445
R3001 VSS.n569 VSS.n568 11.4425
R3002 VSS.n2290 VSS.n2289 11.424
R3003 VSS.n1760 VSS.t22 11.2983
R3004 VSS.n789 VSS.t259 10.9485
R3005 VSS.n1587 VSS.t166 10.9433
R3006 VSS.n849 VSS.n848 10.0314
R3007 VSS.n194 VSS.t58 9.87492
R3008 VSS.n1871 VSS.t589 9.62538
R3009 VSS.n1465 VSS.t634 9.5108
R3010 VSS.n2162 VSS.n2157 9.42079
R3011 VSS.t460 VSS.n1434 9.41994
R3012 VSS.t4 VSS.n1436 9.41738
R3013 VSS.n140 VSS.t285 9.40866
R3014 VSS.n1442 VSS.t54 9.39781
R3015 VSS.n1440 VSS.t462 9.39484
R3016 VSS.n2192 VSS.t483 9.37686
R3017 VSS.n67 VSS.t435 9.3736
R3018 VSS.n52 VSS.t562 9.3736
R3019 VSS.n2263 VSS.t84 9.3736
R3020 VSS.n2155 VSS.t81 9.3736
R3021 VSS.n2271 VSS.t565 9.3736
R3022 VSS.n2313 VSS.t142 9.3736
R3023 VSS.n2255 VSS.t441 9.3736
R3024 VSS.n2234 VSS.t312 9.3736
R3025 VSS.n1061 VSS.t97 9.36804
R3026 VSS.n1055 VSS.t514 9.36804
R3027 VSS.n1087 VSS.t364 9.36804
R3028 VSS.n1135 VSS.t139 9.36804
R3029 VSS.n1443 VSS.t540 9.36804
R3030 VSS.n1053 VSS.t99 9.36804
R3031 VSS.n1169 VSS.t154 9.36804
R3032 VSS.n380 VSS.t61 9.3645
R3033 VSS.n384 VSS.n345 9.3221
R3034 VSS.n382 VSS.t449 9.3221
R3035 VSS.n378 VSS.n351 9.3221
R3036 VSS.n357 VSS.t331 9.3221
R3037 VSS.n385 VSS.t178 9.30652
R3038 VSS.n350 VSS.t147 9.30652
R3039 VSS.n365 VSS.t613 9.30652
R3040 VSS.n2379 VSS.t268 9.30652
R3041 VSS.n115 VSS.t529 9.30652
R3042 VSS.n133 VSS.t576 9.30652
R3043 VSS.n2211 VSS.t128 9.30652
R3044 VSS.n2206 VSS.t606 9.30652
R3045 VSS.n2202 VSS.t296 9.30652
R3046 VSS.n111 VSS.t617 9.30652
R3047 VSS.n360 VSS.t51 9.30652
R3048 VSS.n117 VSS.t487 9.30518
R3049 VSS.n130 VSS.t366 9.30518
R3050 VSS.n2197 VSS.t491 9.30518
R3051 VSS.n123 VSS.t536 9.30323
R3052 VSS.n2372 VSS.t172 9.3025
R3053 VSS.n2373 VSS.n1 9.30189
R3054 VSS.n2374 VSS.t1 9.30189
R3055 VSS.n139 VSS.t622 9.29981
R3056 VSS.n2200 VSS.t557 9.25414
R3057 VSS.n576 VSS.n574 9.05343
R3058 VSS.n1472 VSS.n564 8.84542
R3059 VSS.n1468 VSS.t149 8.84542
R3060 VSS.n1475 VSS.n1473 8.84448
R3061 VSS.t108 VSS.n1126 8.77835
R3062 VSS.n2215 VSS.n2213 8.62119
R3063 VSS.n2141 VSS.t59 8.4763
R3064 VSS.n1799 VSS.n1798 8.13028
R3065 VSS.n2147 VSS.n2146 8.00543
R3066 VSS.n854 VSS.n853 7.52365
R3067 VSS.n370 VSS.n369 7.39136
R3068 VSS VSS.t309 7.30633
R3069 VSS.n1170 VSS.t641 7.19156
R3070 VSS.n1445 VSS.t5 7.19156
R3071 VSS.n1083 VSS.t253 7.19156
R3072 VSS.n1086 VSS.t230 7.19156
R3073 VSS.n1464 VSS.n573 7.19156
R3074 VSS.n356 VSS.t329 7.19156
R3075 VSS.n2308 VSS.t114 7.19156
R3076 VSS.n2303 VSS.t255 7.19156
R3077 VSS.n2302 VSS.t600 7.19156
R3078 VSS.n2179 VSS.t453 7.19156
R3079 VSS.n2260 VSS.t637 7.19156
R3080 VSS.n2246 VSS.t626 7.19156
R3081 VSS.n2241 VSS.t90 7.19156
R3082 VSS.n2240 VSS.t145 7.19156
R3083 VSS.n39 VSS.t18 7.19156
R3084 VSS.n2158 VSS.t493 7.19156
R3085 VSS.n2225 VSS.t608 7.19156
R3086 VSS.n2220 VSS.t527 7.19156
R3087 VSS.n2219 VSS.t489 7.19156
R3088 VSS.n85 VSS.t369 7.19156
R3089 VSS.n87 VSS.t321 7.19156
R3090 VSS.n13 VSS.t232 7.19156
R3091 VSS.n2189 VSS.t163 7.19156
R3092 VSS.n73 VSS.t325 7.19156
R3093 VSS.n71 VSS.t319 7.19156
R3094 VSS.n69 VSS.t532 7.19156
R3095 VSS.n1082 VSS.t274 7.18989
R3096 VSS.n1072 VSS.n883 7.18989
R3097 VSS.n595 VSS.n594 7.18989
R3098 VSS.n882 VSS.t362 7.18989
R3099 VSS VSS.t463 7.18966
R3100 VSS.n2347 VSS.t555 7.17323
R3101 VSS.n2345 VSS.t112 7.17323
R3102 VSS.n2322 VSS.t168 7.17323
R3103 VSS.n2178 VSS.t525 7.17323
R3104 VSS.n135 VSS.t244 7.17156
R3105 VSS.n2334 VSS.t235 7.16989
R3106 VSS.n2332 VSS.t349 7.16989
R3107 VSS.n2360 VSS.t465 7.16656
R3108 VSS.n2357 VSS.t212 7.16656
R3109 VSS.n2461 VSS.t242 7.16085
R3110 VSS.n2382 VSS.t240 7.15156
R3111 VSS.n94 VSS.t136 7.13489
R3112 VSS.n96 VSS.t78 7.13489
R3113 VSS.n100 VSS.t218 7.13489
R3114 VSS.n2265 VSS.t88 7.13323
R3115 VSS.n2267 VSS.t668 7.13323
R3116 VSS.n2269 VSS.t497 7.13323
R3117 VSS.n2163 VSS.t170 7.13156
R3118 VSS.n2168 VSS.t316 7.13156
R3119 VSS.n2169 VSS.t359 7.13156
R3120 VSS.n122 VSS.n121 7.1285
R3121 VSS.n54 VSS.t346 7.12823
R3122 VSS.n59 VSS.t603 7.12823
R3123 VSS.n62 VSS.t215 7.12823
R3124 VSS.n1438 VSS.t55 7.12323
R3125 VSS.n1128 VSS.t109 7.12323
R3126 VSS.n1145 VSS.t475 7.12156
R3127 VSS.n1088 VSS.t469 7.11989
R3128 VSS.n1105 VSS.t277 7.11156
R3129 VSS.n1446 VSS.t461 7.03656
R3130 VSS.n1172 VSS.t107 7.02489
R3131 VSS.n2204 VSS.t444 6.88656
R3132 VSS.n2207 VSS.t652 6.88656
R3133 VSS.n1104 VSS.n1103 6.84992
R3134 VSS.n1461 VSS.n578 6.64949
R3135 VSS.n892 VSS.n891 6.61132
R3136 VSS.n895 VSS.t222 6.61132
R3137 VSS.n987 VSS.n886 6.61132
R3138 VSS.n1069 VSS.t207 6.61132
R3139 VSS.n1457 VSS.t15 6.59043
R3140 VSS.n1454 VSS.n586 6.59043
R3141 VSS.n1449 VSS.t67 6.59043
R3142 VSS.n1072 VSS.n1071 6.46225
R3143 VSS.n1447 VSS 6.32556
R3144 VSS.n792 VSS.t257 6.25652
R3145 VSS.n1584 VSS.t165 6.25351
R3146 VSS.n1812 VSS.t302 6.21739
R3147 VSS VSS.t248 6.02876
R3148 VSS.n2187 VSS.n2186 6.01414
R3149 VSS.n2187 VSS.t272 6.01414
R3150 VSS.n108 VSS.n107 6.01414
R3151 VSS.n108 VSS.t503 6.01414
R3152 VSS.n2049 VSS.n2048 5.99763
R3153 VSS.n1935 VSS.n1934 5.99763
R3154 VSS.n757 VSS.n756 5.99763
R3155 VSS.n552 VSS.n551 5.99763
R3156 VSS.n1062 VSS.n1061 5.94887
R3157 VSS.n2182 VSS.t479 5.91399
R3158 VSS.n2315 VSS.t467 5.91399
R3159 VSS.n2317 VSS.t161 5.91399
R3160 VSS.n2249 VSS.t156 5.91399
R3161 VSS.n2252 VSS.t473 5.91399
R3162 VSS.n44 VSS.t334 5.91399
R3163 VSS.n2228 VSS.t471 5.91399
R3164 VSS.n2231 VSS.t477 5.91399
R3165 VSS.n29 VSS.t534 5.91399
R3166 VSS.n78 VSS.t481 5.91399
R3167 VSS.n18 VSS.t615 5.91399
R3168 VSS.n75 VSS.t551 5.91399
R3169 VSS.n137 VSS.t323 5.89898
R3170 VSS.n2342 VSS.t553 5.89565
R3171 VSS.n2339 VSS.t356 5.89565
R3172 VSS.n2274 VSS.t53 5.89565
R3173 VSS.n2278 VSS.t568 5.89565
R3174 VSS.n2329 VSS.t49 5.89232
R3175 VSS.n2326 VSS.t176 5.89232
R3176 VSS.n2354 VSS.t538 5.88898
R3177 VSS.n2351 VSS.t134 5.88898
R3178 VSS.n98 VSS.t354 5.85732
R3179 VSS.n2281 VSS.t567 5.85565
R3180 VSS.n2174 VSS.t190 5.85398
R3181 VSS.n63 VSS.t132 5.85065
R3182 VSS.n984 VSS.n983 5.81653
R3183 VSS.n1303 VSS.t522 5.80213
R3184 VSS.n1208 VSS.t288 5.80213
R3185 VSS.n1293 VSS.n1251 5.80209
R3186 VSS.n1218 VSS.n1181 5.80209
R3187 VSS VSS.t261 5.6909
R3188 VSS VSS.t546 5.6909
R3189 VSS.n567 VSS.n566 5.4005
R3190 VSS.n567 VSS.t151 5.4005
R3191 VSS.n1132 VSS.n1131 5.37891
R3192 VSS.n2461 VSS.n2460 5.37816
R3193 VSS.n1754 VSS.t224 5.27799
R3194 VSS.n1821 VSS.n1820 5.26095
R3195 VSS.n2289 VSS 5.20137
R3196 VSS.n104 VSS.n93 5.2005
R3197 VSS.n103 VSS.n95 5.2005
R3198 VSS.n102 VSS.n101 5.2005
R3199 VSS.n99 VSS.n97 5.2005
R3200 VSS VSS.n1442 5.2005
R3201 VSS.n1440 VSS 5.2005
R3202 VSS.n1134 VSS.n1133 5.2005
R3203 VSS.n1097 VSS.n1096 5.2005
R3204 VSS.n1095 VSS.n1094 5.2005
R3205 VSS.n1084 VSS 5.2005
R3206 VSS.n1147 VSS 5.2005
R3207 VSS.n1146 VSS 5.2005
R3208 VSS VSS.n1085 5.2005
R3209 VSS.n1471 VSS.n565 5.2005
R3210 VSS.n1473 VSS.n563 5.2005
R3211 VSS.n986 VSS.n985 5.2005
R3212 VSS.n985 VSS.n984 5.2005
R3213 VSS.n904 VSS.n902 5.2005
R3214 VSS.n904 VSS.n903 5.2005
R3215 VSS.n1052 VSS.n1051 5.2005
R3216 VSS VSS.n1127 5.2005
R3217 VSS.n1161 VSS 5.2005
R3218 VSS.n387 VSS.n386 5.2005
R3219 VSS.n383 VSS.n346 5.2005
R3220 VSS.n367 VSS.n366 5.2005
R3221 VSS.n2376 VSS.n2375 5.2005
R3222 VSS.n2371 VSS.n2370 5.2005
R3223 VSS.n2381 VSS.n2380 5.2005
R3224 VSS.n2378 VSS.n2377 5.2005
R3225 VSS VSS.n848 5.2005
R3226 VSS.n850 VSS.n849 5.2005
R3227 VSS.n1080 VSS 5.2005
R3228 VSS VSS.n1077 5.2005
R3229 VSS VSS.n1081 5.2005
R3230 VSS.n1074 VSS 5.2005
R3231 VSS VSS.n1436 5.2005
R3232 VSS.n1444 VSS.n1437 5.2005
R3233 VSS VSS.n1434 5.2005
R3234 VSS.n1174 VSS 5.2005
R3235 VSS.n354 VSS.n353 5.2005
R3236 VSS.n349 VSS.n348 5.2005
R3237 VSS.n381 VSS.n347 5.2005
R3238 VSS.n132 VSS.n131 5.2005
R3239 VSS.n2148 VSS.n140 5.2005
R3240 VSS.n2149 VSS.n138 5.2005
R3241 VSS.n2151 VSS.n136 5.2005
R3242 VSS.n2153 VSS.n134 5.2005
R3243 VSS.n2156 VSS.n2155 5.2005
R3244 VSS.n2165 VSS.n2164 5.2005
R3245 VSS.n2167 VSS.n2166 5.2005
R3246 VSS.n2171 VSS.n2170 5.2005
R3247 VSS.n2173 VSS.n2172 5.2005
R3248 VSS.n2336 VSS.n34 5.2005
R3249 VSS.n2333 VSS.n36 5.2005
R3250 VSS.n2330 VSS.n41 5.2005
R3251 VSS.n2327 VSS.n46 5.2005
R3252 VSS.n2251 VSS.n2250 5.2005
R3253 VSS.n43 VSS.n42 5.2005
R3254 VSS.n38 VSS.n37 5.2005
R3255 VSS.n2160 VSS.n2159 5.2005
R3256 VSS.n74 VSS.n5 5.2005
R3257 VSS.n72 VSS.n5 5.2005
R3258 VSS.n70 VSS.n5 5.2005
R3259 VSS.n68 VSS.n5 5.2005
R3260 VSS.n67 VSS.n7 5.2005
R3261 VSS.n53 VSS.n52 5.2005
R3262 VSS.n56 VSS.n55 5.2005
R3263 VSS.n58 VSS.n57 5.2005
R3264 VSS.n61 VSS.n60 5.2005
R3265 VSS.n65 VSS.n64 5.2005
R3266 VSS.n2352 VSS.n20 5.2005
R3267 VSS.n2355 VSS.n15 5.2005
R3268 VSS.n2358 VSS.n10 5.2005
R3269 VSS.n2362 VSS.n2361 5.2005
R3270 VSS.n80 VSS.n79 5.2005
R3271 VSS.n17 VSS.n16 5.2005
R3272 VSS.n12 VSS.n11 5.2005
R3273 VSS.n2190 VSS.n2188 5.2005
R3274 VSS.n2194 VSS.n2193 5.2005
R3275 VSS.n2199 VSS.n2198 5.2005
R3276 VSS.n2196 VSS.n2195 5.2005
R3277 VSS.n2201 VSS.n2185 5.2005
R3278 VSS.n2209 VSS.n2208 5.2005
R3279 VSS.n2210 VSS.n2209 5.2005
R3280 VSS.n2213 VSS.n2212 5.2005
R3281 VSS.n2248 VSS.n2247 5.2005
R3282 VSS.n2245 VSS.n2244 5.2005
R3283 VSS.n2243 VSS.n2242 5.2005
R3284 VSS.n2239 VSS.n2238 5.2005
R3285 VSS.n2256 VSS.n2255 5.2005
R3286 VSS.n2227 VSS.n2226 5.2005
R3287 VSS.n2224 VSS.n2223 5.2005
R3288 VSS.n2222 VSS.n2221 5.2005
R3289 VSS.n2218 VSS.n2217 5.2005
R3290 VSS.n2235 VSS.n2234 5.2005
R3291 VSS.n2340 VSS.n31 5.2005
R3292 VSS.n2343 VSS.n26 5.2005
R3293 VSS.n2346 VSS.n24 5.2005
R3294 VSS.n2348 VSS.n23 5.2005
R3295 VSS.n2230 VSS.n2229 5.2005
R3296 VSS.n28 VSS.n27 5.2005
R3297 VSS.n86 VSS.n84 5.2005
R3298 VSS.n89 VSS.n88 5.2005
R3299 VSS.n110 VSS.n109 5.2005
R3300 VSS.n125 VSS.n124 5.2005
R3301 VSS.n129 VSS.n128 5.2005
R3302 VSS.n120 VSS.n119 5.2005
R3303 VSS.n116 VSS.n48 5.2005
R3304 VSS.n1452 VSS.n589 5.2005
R3305 VSS.n1455 VSS.n585 5.2005
R3306 VSS.n1460 VSS.n580 5.2005
R3307 VSS.n1466 VSS.n572 5.2005
R3308 VSS.n1467 VSS.n571 5.2005
R3309 VSS.n1469 VSS.n570 5.2005
R3310 VSS VSS.n577 5.2005
R3311 VSS.n1057 VSS.n1056 5.2005
R3312 VSS.n1060 VSS.n1059 5.2005
R3313 VSS.n2286 VSS.n2264 5.2005
R3314 VSS.n2285 VSS.n2266 5.2005
R3315 VSS.n2284 VSS.n2268 5.2005
R3316 VSS.n2283 VSS.n2282 5.2005
R3317 VSS.n2313 VSS.n2312 5.2005
R3318 VSS.n2273 VSS.n2272 5.2005
R3319 VSS.n2321 VSS.n2177 5.2005
R3320 VSS.n2323 VSS.n2176 5.2005
R3321 VSS.n2316 VSS.n2181 5.2005
R3322 VSS.n2318 VSS.n2180 5.2005
R3323 VSS.n2259 VSS.n2258 5.2005
R3324 VSS.n2262 VSS.n2261 5.2005
R3325 VSS.n2310 VSS.n2309 5.2005
R3326 VSS.n2307 VSS.n2306 5.2005
R3327 VSS.n2305 VSS.n2304 5.2005
R3328 VSS.n2301 VSS.n2300 5.2005
R3329 VSS.n2271 VSS.n2270 5.2005
R3330 VSS.n359 VSS.n358 5.2005
R3331 VSS.n362 VSS.n361 5.2005
R3332 VSS.n276 VSS.n0 5.2005
R3333 VSS.n2024 VSS.n201 5.15437
R3334 VSS.n396 VSS.n330 5.15437
R3335 VSS.n244 VSS.n243 5.13377
R3336 VSS VSS.t186 5.11524
R3337 VSS VSS.t665 5.11524
R3338 VSS.n1070 VSS.n1069 5.10136
R3339 VSS.n2051 VSS.t588 5.0898
R3340 VSS.n1937 VSS.t590 5.0898
R3341 VSS.n759 VSS.t194 5.0898
R3342 VSS.n554 VSS.t593 5.0898
R3343 VSS.n1067 VSS.n1066 5.07824
R3344 VSS.n1463 VSS.n1462 5.06621
R3345 VSS.n1456 VSS.t344 5.04745
R3346 VSS.n2013 VSS.t182 5.04596
R3347 VSS.n1453 VSS.n587 5.02656
R3348 VSS.n1448 VSS.t47 4.99985
R3349 VSS.n1759 VSS.n546 4.79593
R3350 VSS.n1779 VSS.t26 4.79593
R3351 VSS.n1794 VSS.n452 4.79593
R3352 VSS.n1819 VSS.t303 4.79593
R3353 VSS.n2364 VSS.n7 4.61862
R3354 VSS.n2451 VSS.n2384 4.53825
R3355 VSS.n2456 VSS.n2386 4.52915
R3356 VSS.n2457 VSS.n2384 4.52872
R3357 VSS VSS.n2386 4.52418
R3358 VSS.n2455 VSS.n2454 4.5005
R3359 VSS.n2457 VSS.n2385 4.5005
R3360 VSS.n1093 VSS.n1092 4.5005
R3361 VSS.n888 VSS.n887 4.5005
R3362 VSS.n369 VSS.n368 4.5005
R3363 VSS.n1967 VSS.t192 4.49211
R3364 VSS.n1353 VSS.n1352 4.44039
R3365 VSS.n2383 VSS.t137 4.37478
R3366 VSS.n2017 VSS.t187 4.32518
R3367 VSS VSS.n2457 4.32389
R3368 VSS.n368 VSS 4.12455
R3369 VSS.n1465 VSS.n1464 3.90454
R3370 VSS.n1130 VSS.n1129 3.69451
R3371 VSS.t365 VSS.t486 3.67489
R3372 VSS.n128 VSS.n48 3.67489
R3373 VSS VSS.n545 3.60246
R3374 VSS VSS.n451 3.60246
R3375 VSS.n2016 VSS.n203 3.51637
R3376 VSS.n403 VSS.n329 3.51637
R3377 VSS.n2049 VSS.n2047 3.51441
R3378 VSS.n2050 VSS.n2045 3.51441
R3379 VSS.n1935 VSS.n1933 3.51441
R3380 VSS.n1936 VSS.n1931 3.51441
R3381 VSS.n757 VSS.n755 3.51441
R3382 VSS.n758 VSS.n753 3.51441
R3383 VSS.n552 VSS.n550 3.51441
R3384 VSS.n553 VSS.n548 3.51441
R3385 VSS.n1470 VSS.n567 3.44542
R3386 VSS.n1450 VSS.n593 3.37758
R3387 VSS.n1458 VSS.n584 3.37758
R3388 VSS.n2191 VSS.n2187 3.36323
R3389 VSS.n893 VSS.n890 3.33532
R3390 VSS.n1068 VSS.n885 3.33532
R3391 VSS.n1459 VSS.n582 3.31443
R3392 VSS.n1451 VSS.n591 3.31443
R3393 VSS.n2146 VSS.t56 3.29665
R3394 VSS.n113 VSS.n108 3.28959
R3395 VSS.n582 VSS.t10 3.2765
R3396 VSS.n582 VSS.n581 3.2765
R3397 VSS.n591 VSS.t75 3.2765
R3398 VSS.n591 VSS.n590 3.2765
R3399 VSS.n890 VSS.t228 3.2765
R3400 VSS.n890 VSS.n889 3.2765
R3401 VSS.n885 VSS.t205 3.2765
R3402 VSS.n885 VSS.n884 3.2765
R3403 VSS.n2408 VSS.t392 3.26618
R3404 VSS.n2401 VSS.t390 3.26618
R3405 VSS.n2394 VSS.t413 3.26618
R3406 VSS.n2387 VSS.t384 3.26618
R3407 VSS.n2418 VSS.t396 3.26618
R3408 VSS.n2425 VSS.t389 3.26618
R3409 VSS.n2432 VSS.t406 3.26618
R3410 VSS.n2439 VSS.t394 3.26618
R3411 VSS.n121 VSS.n120 3.03722
R3412 VSS.n316 VSS.n315 3.00849
R3413 VSS.n319 VSS.n318 3.00849
R3414 VSS.n322 VSS.n321 3.00849
R3415 VSS.n2036 VSS.n2035 3.00849
R3416 VSS.n1144 VSS.n1143 2.85704
R3417 VSS.n2370 VSS.t171 2.80545
R3418 VSS.n2377 VSS.t267 2.80102
R3419 VSS.n1142 VSS.n1089 2.69391
R3420 VSS.n1143 VSS.n1087 2.66505
R3421 VSS.n198 VSS.t57 2.63368
R3422 VSS.n1151 VSS.n1150 2.61336
R3423 VSS.n440 VSS.n420 2.60693
R3424 VSS.n865 VSS.n861 2.60693
R3425 VSS.n1483 VSS.n1482 2.60693
R3426 VSS.n1656 VSS.n1655 2.60693
R3427 VSS.n163 VSS.n162 2.60371
R3428 VSS.n1556 VSS.n1555 2.60371
R3429 VSS.n822 VSS.n751 2.60371
R3430 VSS.n1357 VSS.n1177 2.60343
R3431 VSS.n1335 VSS.n1247 2.60343
R3432 VSS.n259 VSS.n258 2.60243
R3433 VSS.n772 VSS.n771 2.60243
R3434 VSS.n1848 VSS.n289 2.60179
R3435 VSS.n1500 VSS.n1480 2.60179
R3436 VSS.n842 VSS.n619 2.60179
R3437 VSS.n2069 VSS.n2068 2.60179
R3438 VSS.n1310 VSS.n1309 2.60148
R3439 VSS.n1204 VSS.n1203 2.60148
R3440 VSS.n395 VSS.n394 2.6005
R3441 VSS.n394 VSS.n393 2.6005
R3442 VSS.n399 VSS.n398 2.6005
R3443 VSS.n398 VSS.n397 2.6005
R3444 VSS.n402 VSS.n401 2.6005
R3445 VSS.n401 VSS.n400 2.6005
R3446 VSS.n406 VSS.n405 2.6005
R3447 VSS.n405 VSS.n404 2.6005
R3448 VSS.n409 VSS.n408 2.6005
R3449 VSS.n408 VSS.n407 2.6005
R3450 VSS.n413 VSS.n412 2.6005
R3451 VSS.n412 VSS.n411 2.6005
R3452 VSS.n177 VSS.n176 2.6005
R3453 VSS.n176 VSS.n175 2.6005
R3454 VSS.n168 VSS.n167 2.6005
R3455 VSS.n167 VSS.n166 2.6005
R3456 VSS.n171 VSS.n170 2.6005
R3457 VSS.n170 VSS.n169 2.6005
R3458 VSS.n174 VSS.n173 2.6005
R3459 VSS.n173 VSS.n172 2.6005
R3460 VSS.n1351 VSS.n1350 2.6005
R3461 VSS.n1345 VSS.n1344 2.6005
R3462 VSS.n1347 VSS.n1346 2.6005
R3463 VSS.n1387 VSS.n1386 2.6005
R3464 VSS.n1380 VSS.n1379 2.6005
R3465 VSS.n1384 VSS.n1383 2.6005
R3466 VSS.n612 VSS.n611 2.6005
R3467 VSS.n611 VSS.n610 2.6005
R3468 VSS.n609 VSS.n608 2.6005
R3469 VSS.n608 VSS.n607 2.6005
R3470 VSS.n606 VSS.n605 2.6005
R3471 VSS.n605 VSS.n604 2.6005
R3472 VSS.n1338 VSS.n1337 2.6005
R3473 VSS.n1342 VSS.n1341 2.6005
R3474 VSS.n1258 VSS.n1257 2.6005
R3475 VSS.n1256 VSS.n1255 2.6005
R3476 VSS.n1253 VSS.n1252 2.6005
R3477 VSS.n1250 VSS.n1249 2.6005
R3478 VSS.n603 VSS.n602 2.6005
R3479 VSS.n602 VSS.n601 2.6005
R3480 VSS.n600 VSS.n599 2.6005
R3481 VSS.n599 VSS.n598 2.6005
R3482 VSS.n1378 VSS.n1377 2.6005
R3483 VSS.n597 VSS.n596 2.6005
R3484 VSS.n1245 VSS.n1244 2.6005
R3485 VSS.n1244 VSS.n1243 2.6005
R3486 VSS.n1242 VSS.n1241 2.6005
R3487 VSS.n1241 VSS.n1240 2.6005
R3488 VSS.n1239 VSS.n1238 2.6005
R3489 VSS.n1238 VSS.n1237 2.6005
R3490 VSS.n1236 VSS.n1235 2.6005
R3491 VSS.n1235 VSS.n1234 2.6005
R3492 VSS.n1233 VSS.n1232 2.6005
R3493 VSS.n1232 VSS.n1231 2.6005
R3494 VSS.n1330 VSS.n1329 2.6005
R3495 VSS.n1329 VSS.n1328 2.6005
R3496 VSS.n1327 VSS.n1326 2.6005
R3497 VSS.n1326 VSS.n1325 2.6005
R3498 VSS.n1324 VSS.n1323 2.6005
R3499 VSS.n1323 VSS.n1322 2.6005
R3500 VSS.n1321 VSS.n1320 2.6005
R3501 VSS.n1320 VSS.n1319 2.6005
R3502 VSS.n1333 VSS.n1332 2.6005
R3503 VSS.n1332 VSS.n1331 2.6005
R3504 VSS.n1230 VSS.n1229 2.6005
R3505 VSS.n1226 VSS.n1225 2.6005
R3506 VSS.n1221 VSS.n1220 2.6005
R3507 VSS.n1220 VSS.n1219 2.6005
R3508 VSS.n1217 VSS.n1216 2.6005
R3509 VSS.n1216 VSS.n1215 2.6005
R3510 VSS.n1214 VSS.n1213 2.6005
R3511 VSS.n1213 VSS.n1212 2.6005
R3512 VSS.n1211 VSS.n1210 2.6005
R3513 VSS.n1210 VSS.n1209 2.6005
R3514 VSS.n1207 VSS.n1206 2.6005
R3515 VSS.n1206 VSS.n1205 2.6005
R3516 VSS.n1224 VSS.n1223 2.6005
R3517 VSS.n1316 VSS.n1315 2.6005
R3518 VSS.n1312 VSS.n1311 2.6005
R3519 VSS.n1292 VSS.n1291 2.6005
R3520 VSS.n1291 VSS.n1290 2.6005
R3521 VSS.n1296 VSS.n1295 2.6005
R3522 VSS.n1295 VSS.n1294 2.6005
R3523 VSS.n1299 VSS.n1298 2.6005
R3524 VSS.n1298 VSS.n1297 2.6005
R3525 VSS.n1302 VSS.n1301 2.6005
R3526 VSS.n1301 VSS.n1300 2.6005
R3527 VSS.n1306 VSS.n1305 2.6005
R3528 VSS.n1305 VSS.n1304 2.6005
R3529 VSS.n1309 VSS.n1308 2.6005
R3530 VSS.n507 VSS.n506 2.6005
R3531 VSS.n506 VSS.n505 2.6005
R3532 VSS.n511 VSS.n510 2.6005
R3533 VSS.n510 VSS.n509 2.6005
R3534 VSS.n495 VSS.n494 2.6005
R3535 VSS.n494 VSS.n493 2.6005
R3536 VSS.n498 VSS.n497 2.6005
R3537 VSS.n497 VSS.n496 2.6005
R3538 VSS.n501 VSS.n500 2.6005
R3539 VSS.n500 VSS.n499 2.6005
R3540 VSS.n504 VSS.n503 2.6005
R3541 VSS.n503 VSS.n502 2.6005
R3542 VSS.n1268 VSS.n1267 2.6005
R3543 VSS.n1267 VSS.n1266 2.6005
R3544 VSS.n1271 VSS.n1270 2.6005
R3545 VSS.n1270 VSS.n1269 2.6005
R3546 VSS.n1274 VSS.n1273 2.6005
R3547 VSS.n1273 VSS.n1272 2.6005
R3548 VSS.n1277 VSS.n1276 2.6005
R3549 VSS.n1276 VSS.n1275 2.6005
R3550 VSS.n1280 VSS.n1279 2.6005
R3551 VSS.n1279 VSS.n1278 2.6005
R3552 VSS.n1283 VSS.n1282 2.6005
R3553 VSS.n1282 VSS.n1281 2.6005
R3554 VSS.n1286 VSS.n1285 2.6005
R3555 VSS.n1285 VSS.n1284 2.6005
R3556 VSS.n1289 VSS.n1288 2.6005
R3557 VSS.n1288 VSS.n1287 2.6005
R3558 VSS.n485 VSS.n484 2.6005
R3559 VSS.n489 VSS.n488 2.6005
R3560 VSS.n491 VSS.n490 2.6005
R3561 VSS.n1264 VSS.n1263 2.6005
R3562 VSS.n1262 VSS.n1261 2.6005
R3563 VSS.n927 VSS.n926 2.6005
R3564 VSS.n926 VSS.n925 2.6005
R3565 VSS.n1425 VSS.n1424 2.6005
R3566 VSS.n1426 VSS.n1425 2.6005
R3567 VSS.n1423 VSS.n1422 2.6005
R3568 VSS.n1422 VSS.n1421 2.6005
R3569 VSS.n967 VSS.n929 2.6005
R3570 VSS.n929 VSS.n928 2.6005
R3571 VSS.n963 VSS.n962 2.6005
R3572 VSS.n962 VSS.n961 2.6005
R3573 VSS.n960 VSS.n959 2.6005
R3574 VSS.n959 VSS.n958 2.6005
R3575 VSS.n957 VSS.n956 2.6005
R3576 VSS.n956 VSS.n955 2.6005
R3577 VSS.n954 VSS.n953 2.6005
R3578 VSS.n953 VSS.n952 2.6005
R3579 VSS.n966 VSS.n965 2.6005
R3580 VSS.n965 VSS.n964 2.6005
R3581 VSS.n951 VSS.n950 2.6005
R3582 VSS.n935 VSS.n934 2.6005
R3583 VSS.n938 VSS.n937 2.6005
R3584 VSS.n940 VSS.n939 2.6005
R3585 VSS.n944 VSS.n943 2.6005
R3586 VSS.n946 VSS.n945 2.6005
R3587 VSS.n919 VSS.n918 2.6005
R3588 VSS.n918 VSS.n917 2.6005
R3589 VSS.n916 VSS.n915 2.6005
R3590 VSS.n915 VSS.n914 2.6005
R3591 VSS.n913 VSS.n912 2.6005
R3592 VSS.n912 VSS.n911 2.6005
R3593 VSS.n910 VSS.n909 2.6005
R3594 VSS.n909 VSS.n908 2.6005
R3595 VSS.n907 VSS.n906 2.6005
R3596 VSS.n906 VSS.n905 2.6005
R3597 VSS.n931 VSS.n930 2.6005
R3598 VSS.n922 VSS.n921 2.6005
R3599 VSS.n921 VSS.n920 2.6005
R3600 VSS.n982 VSS.n981 2.6005
R3601 VSS.n983 VSS.n982 2.6005
R3602 VSS.n980 VSS.n979 2.6005
R3603 VSS.n979 VSS.n978 2.6005
R3604 VSS.n977 VSS.n976 2.6005
R3605 VSS.n976 VSS.n975 2.6005
R3606 VSS.n974 VSS.n973 2.6005
R3607 VSS.n973 VSS.n972 2.6005
R3608 VSS.n971 VSS.n970 2.6005
R3609 VSS.n970 VSS.n969 2.6005
R3610 VSS.n1047 VSS.n1046 2.6005
R3611 VSS.n1045 VSS.n1044 2.6005
R3612 VSS.n990 VSS.n989 2.6005
R3613 VSS.n989 VSS.n988 2.6005
R3614 VSS.n993 VSS.n992 2.6005
R3615 VSS.n992 VSS.n991 2.6005
R3616 VSS.n996 VSS.n995 2.6005
R3617 VSS.n995 VSS.n994 2.6005
R3618 VSS.n999 VSS.n998 2.6005
R3619 VSS.n998 VSS.n997 2.6005
R3620 VSS.n1002 VSS.n1001 2.6005
R3621 VSS.n1001 VSS.n1000 2.6005
R3622 VSS.n1005 VSS.n1004 2.6005
R3623 VSS.n1004 VSS.n1003 2.6005
R3624 VSS.n1008 VSS.n1007 2.6005
R3625 VSS.n1007 VSS.n1006 2.6005
R3626 VSS.n1049 VSS.n1048 2.6005
R3627 VSS.n1050 VSS.n1049 2.6005
R3628 VSS.n852 VSS.n851 2.6005
R3629 VSS.n858 VSS.n857 2.6005
R3630 VSS.n1164 VSS.n1163 2.6005
R3631 VSS.n1163 VSS.n1162 2.6005
R3632 VSS.n1160 VSS.n1159 2.6005
R3633 VSS.n1159 VSS.n1158 2.6005
R3634 VSS.n1157 VSS.n1156 2.6005
R3635 VSS.n1156 VSS.n1155 2.6005
R3636 VSS.n881 VSS.n880 2.6005
R3637 VSS.n880 VSS.n879 2.6005
R3638 VSS.n1125 VSS.n1124 2.6005
R3639 VSS.n1126 VSS.n1125 2.6005
R3640 VSS.n1123 VSS.n1122 2.6005
R3641 VSS.n1115 VSS.n1114 2.6005
R3642 VSS.n1113 VSS.n1112 2.6005
R3643 VSS.n1110 VSS.n1109 2.6005
R3644 VSS.n776 VSS.n775 2.6005
R3645 VSS.n689 VSS.n688 2.6005
R3646 VSS.n687 VSS.n686 2.6005
R3647 VSS.n685 VSS.n684 2.6005
R3648 VSS.n683 VSS.n682 2.6005
R3649 VSS.n681 VSS.n680 2.6005
R3650 VSS.n679 VSS.n678 2.6005
R3651 VSS.n677 VSS.n676 2.6005
R3652 VSS.n675 VSS.n674 2.6005
R3653 VSS.n673 VSS.n672 2.6005
R3654 VSS.n671 VSS.n670 2.6005
R3655 VSS.n669 VSS.n668 2.6005
R3656 VSS.n667 VSS.n666 2.6005
R3657 VSS.n665 VSS.n664 2.6005
R3658 VSS.n663 VSS.n662 2.6005
R3659 VSS.n661 VSS.n660 2.6005
R3660 VSS.n659 VSS.n658 2.6005
R3661 VSS.n821 VSS.n820 2.6005
R3662 VSS.n820 VSS.n819 2.6005
R3663 VSS.n818 VSS.n817 2.6005
R3664 VSS.n817 VSS.n816 2.6005
R3665 VSS.n815 VSS.n814 2.6005
R3666 VSS.n814 VSS.n813 2.6005
R3667 VSS.n812 VSS.n811 2.6005
R3668 VSS.n811 VSS.n810 2.6005
R3669 VSS.n809 VSS.n808 2.6005
R3670 VSS.n808 VSS.n807 2.6005
R3671 VSS.n806 VSS.n805 2.6005
R3672 VSS.n805 VSS.n804 2.6005
R3673 VSS.n803 VSS.n802 2.6005
R3674 VSS.n802 VSS.n801 2.6005
R3675 VSS.n800 VSS.n799 2.6005
R3676 VSS.n799 VSS.n798 2.6005
R3677 VSS.n797 VSS.n796 2.6005
R3678 VSS.n796 VSS.n795 2.6005
R3679 VSS.n794 VSS.n793 2.6005
R3680 VSS.n793 VSS.n792 2.6005
R3681 VSS.n791 VSS.n790 2.6005
R3682 VSS.n790 VSS.n789 2.6005
R3683 VSS.n788 VSS.n787 2.6005
R3684 VSS.n787 VSS.n786 2.6005
R3685 VSS.n785 VSS.n784 2.6005
R3686 VSS.n784 VSS.n783 2.6005
R3687 VSS.n782 VSS.n781 2.6005
R3688 VSS.n781 VSS.n780 2.6005
R3689 VSS.n779 VSS.n778 2.6005
R3690 VSS.n778 VSS.n777 2.6005
R3691 VSS.n775 VSS.n774 2.6005
R3692 VSS.n439 VSS.n438 2.6005
R3693 VSS.n438 VSS.n437 2.6005
R3694 VSS.n435 VSS.n434 2.6005
R3695 VSS.n434 VSS.n433 2.6005
R3696 VSS.n432 VSS.n431 2.6005
R3697 VSS.n431 VSS.n430 2.6005
R3698 VSS.n429 VSS.n428 2.6005
R3699 VSS.n428 VSS.n427 2.6005
R3700 VSS.n426 VSS.n425 2.6005
R3701 VSS.n425 VSS.n424 2.6005
R3702 VSS.n423 VSS.n422 2.6005
R3703 VSS.n422 VSS.n421 2.6005
R3704 VSS.n1875 VSS.n1874 2.6005
R3705 VSS.n1874 VSS.t544 2.6005
R3706 VSS.n1878 VSS.n1877 2.6005
R3707 VSS.n1877 VSS.n1876 2.6005
R3708 VSS.n1881 VSS.n1880 2.6005
R3709 VSS.n1880 VSS.n1879 2.6005
R3710 VSS.n1884 VSS.n1883 2.6005
R3711 VSS.n1883 VSS.n1882 2.6005
R3712 VSS.n1887 VSS.n1886 2.6005
R3713 VSS.n1886 VSS.n1885 2.6005
R3714 VSS.n1890 VSS.n1889 2.6005
R3715 VSS.n1889 VSS.n1888 2.6005
R3716 VSS.n1893 VSS.n1892 2.6005
R3717 VSS.n1892 VSS.n1891 2.6005
R3718 VSS.n1896 VSS.n1895 2.6005
R3719 VSS.n1895 VSS.n1894 2.6005
R3720 VSS.n1899 VSS.n1898 2.6005
R3721 VSS.n1898 VSS.n1897 2.6005
R3722 VSS.n1902 VSS.n1901 2.6005
R3723 VSS.n1901 VSS.n1900 2.6005
R3724 VSS.n625 VSS.n624 2.6005
R3725 VSS.n624 VSS.n623 2.6005
R3726 VSS.n628 VSS.n627 2.6005
R3727 VSS.n627 VSS.n626 2.6005
R3728 VSS.n631 VSS.n630 2.6005
R3729 VSS.n630 VSS.n629 2.6005
R3730 VSS.n634 VSS.n633 2.6005
R3731 VSS.n633 VSS.n632 2.6005
R3732 VSS.n637 VSS.n636 2.6005
R3733 VSS.n636 VSS.n635 2.6005
R3734 VSS.n640 VSS.n639 2.6005
R3735 VSS.n639 VSS.n638 2.6005
R3736 VSS.n643 VSS.n642 2.6005
R3737 VSS.n642 VSS.n641 2.6005
R3738 VSS.n622 VSS.n621 2.6005
R3739 VSS.n621 VSS.n620 2.6005
R3740 VSS.n1108 VSS.n1107 2.6005
R3741 VSS.n1107 VSS.n1106 2.6005
R3742 VSS.n657 VSS.n656 2.6005
R3743 VSS.n656 VSS.n655 2.6005
R3744 VSS.n652 VSS.n651 2.6005
R3745 VSS.n651 VSS.n650 2.6005
R3746 VSS.n649 VSS.n648 2.6005
R3747 VSS.n648 VSS.n647 2.6005
R3748 VSS.n646 VSS.n645 2.6005
R3749 VSS.n645 VSS.n644 2.6005
R3750 VSS.n763 VSS.n762 2.6005
R3751 VSS.n762 VSS.n761 2.6005
R3752 VSS.n766 VSS.n765 2.6005
R3753 VSS.n765 VSS.n764 2.6005
R3754 VSS.n769 VSS.n768 2.6005
R3755 VSS.n768 VSS.n767 2.6005
R3756 VSS.n771 VSS.n770 2.6005
R3757 VSS.n1905 VSS.n1904 2.6005
R3758 VSS.n1904 VSS.n1903 2.6005
R3759 VSS.n1908 VSS.n1907 2.6005
R3760 VSS.n1907 VSS.n1906 2.6005
R3761 VSS.n1911 VSS.n1910 2.6005
R3762 VSS.n1910 VSS.n1909 2.6005
R3763 VSS.n1914 VSS.n1913 2.6005
R3764 VSS.n1913 VSS.n1912 2.6005
R3765 VSS.n1917 VSS.n1916 2.6005
R3766 VSS.n1916 VSS.n1915 2.6005
R3767 VSS.n1920 VSS.n1919 2.6005
R3768 VSS.n1919 VSS.n1918 2.6005
R3769 VSS.n1923 VSS.n1922 2.6005
R3770 VSS.n1922 VSS.n1921 2.6005
R3771 VSS.n1926 VSS.n1925 2.6005
R3772 VSS.n1925 VSS.n1924 2.6005
R3773 VSS.n1929 VSS.n1928 2.6005
R3774 VSS.n1928 VSS.n1927 2.6005
R3775 VSS.n1952 VSS.n1951 2.6005
R3776 VSS.n1951 VSS.n1950 2.6005
R3777 VSS.n1947 VSS.n1946 2.6005
R3778 VSS.n1946 VSS.n1945 2.6005
R3779 VSS.n1944 VSS.n1943 2.6005
R3780 VSS.n1943 VSS.n1942 2.6005
R3781 VSS.n1941 VSS.n1940 2.6005
R3782 VSS.n1940 VSS.n1939 2.6005
R3783 VSS.n250 VSS.n249 2.6005
R3784 VSS.n249 VSS.n248 2.6005
R3785 VSS.n253 VSS.n252 2.6005
R3786 VSS.n252 VSS.n251 2.6005
R3787 VSS.n256 VSS.n255 2.6005
R3788 VSS.n255 VSS.n254 2.6005
R3789 VSS.n258 VSS.n257 2.6005
R3790 VSS.n282 VSS.n281 2.6005
R3791 VSS.n284 VSS.n283 2.6005
R3792 VSS.n287 VSS.n286 2.6005
R3793 VSS.n1851 VSS.n1850 2.6005
R3794 VSS.n1850 VSS.n1849 2.6005
R3795 VSS.n1853 VSS.n1852 2.6005
R3796 VSS.n1856 VSS.n1855 2.6005
R3797 VSS.n1855 VSS.n1854 2.6005
R3798 VSS.n1859 VSS.n1858 2.6005
R3799 VSS.n1858 VSS.n1857 2.6005
R3800 VSS.n1862 VSS.n1861 2.6005
R3801 VSS.n1861 VSS.n1860 2.6005
R3802 VSS.n1865 VSS.n1864 2.6005
R3803 VSS.n1864 VSS.n1863 2.6005
R3804 VSS.n1868 VSS.n1867 2.6005
R3805 VSS.n1867 VSS.n1866 2.6005
R3806 VSS.n1870 VSS.n1869 2.6005
R3807 VSS.n1873 VSS.n1872 2.6005
R3808 VSS.n1872 VSS.n1871 2.6005
R3809 VSS.n1971 VSS.n1970 2.6005
R3810 VSS.n1972 VSS.n1971 2.6005
R3811 VSS.n1969 VSS.n1968 2.6005
R3812 VSS.n1968 VSS.n1967 2.6005
R3813 VSS.n1966 VSS.n1965 2.6005
R3814 VSS.n1965 VSS.n1964 2.6005
R3815 VSS.n1963 VSS.n1962 2.6005
R3816 VSS.n1961 VSS.n1960 2.6005
R3817 VSS.n1959 VSS.n1958 2.6005
R3818 VSS.n1958 VSS.n1957 2.6005
R3819 VSS.n1956 VSS.n1955 2.6005
R3820 VSS.n1955 VSS.n1954 2.6005
R3821 VSS.n240 VSS.n239 2.6005
R3822 VSS.n2001 VSS.n2000 2.6005
R3823 VSS.n261 VSS.n260 2.6005
R3824 VSS.n263 VSS.n262 2.6005
R3825 VSS.n266 VSS.n265 2.6005
R3826 VSS.n265 VSS.n264 2.6005
R3827 VSS.n269 VSS.n268 2.6005
R3828 VSS.n268 VSS.n267 2.6005
R3829 VSS.n271 VSS.n270 2.6005
R3830 VSS.n273 VSS.n272 2.6005
R3831 VSS.n1974 VSS.n1973 2.6005
R3832 VSS.n1973 VSS.n1972 2.6005
R3833 VSS.n1976 VSS.n1975 2.6005
R3834 VSS.n1979 VSS.n1978 2.6005
R3835 VSS.n1978 VSS.n1977 2.6005
R3836 VSS.n1981 VSS.n1980 2.6005
R3837 VSS.n1983 VSS.n1982 2.6005
R3838 VSS.n1985 VSS.n1984 2.6005
R3839 VSS.n1987 VSS.n1986 2.6005
R3840 VSS.n1989 VSS.n1988 2.6005
R3841 VSS.n1992 VSS.n1991 2.6005
R3842 VSS.n1991 VSS.n1990 2.6005
R3843 VSS.n1994 VSS.n1993 2.6005
R3844 VSS.n247 VSS.n246 2.6005
R3845 VSS.n246 VSS.n245 2.6005
R3846 VSS.n1999 VSS.n1998 2.6005
R3847 VSS.n835 VSS.n834 2.6005
R3848 VSS.n834 VSS.n833 2.6005
R3849 VSS.n838 VSS.n837 2.6005
R3850 VSS.n837 VSS.n836 2.6005
R3851 VSS.n841 VSS.n840 2.6005
R3852 VSS.n840 VSS.n839 2.6005
R3853 VSS.n864 VSS.n863 2.6005
R3854 VSS.n863 VSS.n862 2.6005
R3855 VSS.n616 VSS.n615 2.6005
R3856 VSS.n615 VSS.n614 2.6005
R3857 VSS.n1364 VSS.n1363 2.6005
R3858 VSS.n1363 VSS.n1362 2.6005
R3859 VSS.n1367 VSS.n1366 2.6005
R3860 VSS.n1366 VSS.n1365 2.6005
R3861 VSS.n1370 VSS.n1369 2.6005
R3862 VSS.n1369 VSS.n1368 2.6005
R3863 VSS.n1373 VSS.n1372 2.6005
R3864 VSS.n1372 VSS.n1371 2.6005
R3865 VSS.n1361 VSS.n1360 2.6005
R3866 VSS.n1360 VSS.n1359 2.6005
R3867 VSS.n845 VSS.n844 2.6005
R3868 VSS.n844 VSS.n843 2.6005
R3869 VSS.n619 VSS.n618 2.6005
R3870 VSS.n832 VSS.n831 2.6005
R3871 VSS.n831 VSS.n830 2.6005
R3872 VSS.n828 VSS.n827 2.6005
R3873 VSS.n827 VSS.n826 2.6005
R3874 VSS.n825 VSS.n824 2.6005
R3875 VSS.n824 VSS.n823 2.6005
R3876 VSS.n751 VSS.n750 2.6005
R3877 VSS.n443 VSS.n442 2.6005
R3878 VSS.n442 VSS.n441 2.6005
R3879 VSS.n420 VSS.n419 2.6005
R3880 VSS.n446 VSS.n445 2.6005
R3881 VSS.n445 VSS.n444 2.6005
R3882 VSS.n1843 VSS.n1842 2.6005
R3883 VSS.n1842 VSS.n1841 2.6005
R3884 VSS.n1840 VSS.n1839 2.6005
R3885 VSS.n1839 VSS.n1838 2.6005
R3886 VSS.n1837 VSS.n1836 2.6005
R3887 VSS.n1836 VSS.n1835 2.6005
R3888 VSS.n1834 VSS.n1833 2.6005
R3889 VSS.n1833 VSS.n1832 2.6005
R3890 VSS.n1831 VSS.n1830 2.6005
R3891 VSS.n1830 VSS.n1829 2.6005
R3892 VSS.n1846 VSS.n1845 2.6005
R3893 VSS.n1845 VSS.n1844 2.6005
R3894 VSS.n867 VSS.n866 2.6005
R3895 VSS.n871 VSS.n870 2.6005
R3896 VSS.n873 VSS.n872 2.6005
R3897 VSS.n876 VSS.n875 2.6005
R3898 VSS.n878 VSS.n877 2.6005
R3899 VSS.n1418 VSS.n1417 2.6005
R3900 VSS.n1416 VSS.n1415 2.6005
R3901 VSS.n1411 VSS.n1410 2.6005
R3902 VSS.n1389 VSS.n1388 2.6005
R3903 VSS.n1355 VSS.n1354 2.6005
R3904 VSS.n1354 VSS.n1353 2.6005
R3905 VSS.n1177 VSS.n1176 2.6005
R3906 VSS.n1402 VSS.n1401 2.6005
R3907 VSS.n1399 VSS.n1398 2.6005
R3908 VSS.n1396 VSS.n1395 2.6005
R3909 VSS.n1394 VSS.n1393 2.6005
R3910 VSS.n1404 VSS.n1403 2.6005
R3911 VSS.n1408 VSS.n1407 2.6005
R3912 VSS.n1392 VSS.n1391 2.6005
R3913 VSS.n1391 VSS.n1390 2.6005
R3914 VSS.n1184 VSS.n1183 2.6005
R3915 VSS.n1183 VSS.n1182 2.6005
R3916 VSS.n1187 VSS.n1186 2.6005
R3917 VSS.n1186 VSS.n1185 2.6005
R3918 VSS.n1190 VSS.n1189 2.6005
R3919 VSS.n1189 VSS.n1188 2.6005
R3920 VSS.n1194 VSS.n1193 2.6005
R3921 VSS.n1193 VSS.n1192 2.6005
R3922 VSS.n1197 VSS.n1196 2.6005
R3923 VSS.n1196 VSS.n1195 2.6005
R3924 VSS.n1200 VSS.n1199 2.6005
R3925 VSS.n1199 VSS.n1198 2.6005
R3926 VSS.n1180 VSS.n1179 2.6005
R3927 VSS.n1179 VSS.n1178 2.6005
R3928 VSS.n1203 VSS.n1202 2.6005
R3929 VSS.n376 VSS.n375 2.6005
R3930 VSS.n375 VSS.n374 2.6005
R3931 VSS.n327 VSS.n326 2.6005
R3932 VSS.n323 VSS.n322 2.6005
R3933 VSS.n320 VSS.n319 2.6005
R3934 VSS.n317 VSS.n316 2.6005
R3935 VSS.n314 VSS.n313 2.6005
R3936 VSS.n312 VSS.n311 2.6005
R3937 VSS.n416 VSS.n415 2.6005
R3938 VSS.n415 VSS.n414 2.6005
R3939 VSS.n238 VSS.n237 2.6005
R3940 VSS.n228 VSS.n227 2.6005
R3941 VSS.n230 VSS.n229 2.6005
R3942 VSS.n233 VSS.n232 2.6005
R3943 VSS.n235 VSS.n234 2.6005
R3944 VSS.n2027 VSS.n2026 2.6005
R3945 VSS.n2026 VSS.n2025 2.6005
R3946 VSS.n2023 VSS.n2022 2.6005
R3947 VSS.n2022 VSS.n2021 2.6005
R3948 VSS.n2019 VSS.n2018 2.6005
R3949 VSS.n2018 VSS.n2017 2.6005
R3950 VSS.n2015 VSS.n2014 2.6005
R3951 VSS.n2014 VSS.n2013 2.6005
R3952 VSS.n2012 VSS.n2011 2.6005
R3953 VSS.n2011 VSS.n2010 2.6005
R3954 VSS.n2008 VSS.n2007 2.6005
R3955 VSS.n2007 VSS.n2006 2.6005
R3956 VSS.n2005 VSS.n2004 2.6005
R3957 VSS.n208 VSS.n207 2.6005
R3958 VSS.n207 VSS.n206 2.6005
R3959 VSS.n211 VSS.n210 2.6005
R3960 VSS.n210 VSS.n209 2.6005
R3961 VSS.n214 VSS.n213 2.6005
R3962 VSS.n213 VSS.n212 2.6005
R3963 VSS.n217 VSS.n216 2.6005
R3964 VSS.n216 VSS.n215 2.6005
R3965 VSS.n220 VSS.n219 2.6005
R3966 VSS.n219 VSS.n218 2.6005
R3967 VSS.n223 VSS.n222 2.6005
R3968 VSS.n222 VSS.n221 2.6005
R3969 VSS.n225 VSS.n224 2.6005
R3970 VSS.n205 VSS.n204 2.6005
R3971 VSS.n2040 VSS.n2039 2.6005
R3972 VSS.n2037 VSS.n2036 2.6005
R3973 VSS.n2034 VSS.n2033 2.6005
R3974 VSS.n2032 VSS.n2031 2.6005
R3975 VSS.n2042 VSS.n2041 2.6005
R3976 VSS.n2029 VSS.n2028 2.6005
R3977 VSS.n291 VSS.n290 2.6005
R3978 VSS.n333 VSS.n332 2.6005
R3979 VSS.n335 VSS.n334 2.6005
R3980 VSS.n338 VSS.n337 2.6005
R3981 VSS.n340 VSS.n339 2.6005
R3982 VSS.n344 VSS.n343 2.6005
R3983 VSS.n392 VSS.n391 2.6005
R3984 VSS.n391 VSS.n390 2.6005
R3985 VSS.n537 VSS.n536 2.6005
R3986 VSS.n539 VSS.n538 2.6005
R3987 VSS.n543 VSS.n542 2.6005
R3988 VSS.n294 VSS.n293 2.6005
R3989 VSS.n293 VSS.n292 2.6005
R3990 VSS.n297 VSS.n296 2.6005
R3991 VSS.n296 VSS.n295 2.6005
R3992 VSS.n300 VSS.n299 2.6005
R3993 VSS.n299 VSS.n298 2.6005
R3994 VSS.n303 VSS.n302 2.6005
R3995 VSS.n302 VSS.n301 2.6005
R3996 VSS.n306 VSS.n305 2.6005
R3997 VSS.n305 VSS.n304 2.6005
R3998 VSS.n309 VSS.n308 2.6005
R3999 VSS.n308 VSS.n307 2.6005
R4000 VSS.n518 VSS.n517 2.6005
R4001 VSS.n517 VSS.n516 2.6005
R4002 VSS.n521 VSS.n520 2.6005
R4003 VSS.n520 VSS.n519 2.6005
R4004 VSS.n524 VSS.n523 2.6005
R4005 VSS.n523 VSS.n522 2.6005
R4006 VSS.n527 VSS.n526 2.6005
R4007 VSS.n526 VSS.n525 2.6005
R4008 VSS.n530 VSS.n529 2.6005
R4009 VSS.n529 VSS.n528 2.6005
R4010 VSS.n534 VSS.n533 2.6005
R4011 VSS.n533 VSS.n532 2.6005
R4012 VSS.n515 VSS.n514 2.6005
R4013 VSS.n514 VSS.n513 2.6005
R4014 VSS.n456 VSS.n455 2.6005
R4015 VSS.n455 VSS.n454 2.6005
R4016 VSS.n479 VSS.n478 2.6005
R4017 VSS.n476 VSS.n475 2.6005
R4018 VSS.n474 VSS.n473 2.6005
R4019 VSS.n473 VSS.n472 2.6005
R4020 VSS.n471 VSS.n470 2.6005
R4021 VSS.n470 VSS.n469 2.6005
R4022 VSS.n468 VSS.n467 2.6005
R4023 VSS.n467 VSS.n466 2.6005
R4024 VSS.n465 VSS.n464 2.6005
R4025 VSS.n464 VSS.n463 2.6005
R4026 VSS.n462 VSS.n461 2.6005
R4027 VSS.n461 VSS.n460 2.6005
R4028 VSS.n459 VSS.n458 2.6005
R4029 VSS.n458 VSS.n457 2.6005
R4030 VSS.n481 VSS.n480 2.6005
R4031 VSS.n748 VSS.n747 2.6005
R4032 VSS.n747 VSS.n746 2.6005
R4033 VSS.n692 VSS.n691 2.6005
R4034 VSS.n691 VSS.n690 2.6005
R4035 VSS.n695 VSS.n694 2.6005
R4036 VSS.n694 VSS.n693 2.6005
R4037 VSS.n698 VSS.n697 2.6005
R4038 VSS.n697 VSS.n696 2.6005
R4039 VSS.n701 VSS.n700 2.6005
R4040 VSS.n700 VSS.n699 2.6005
R4041 VSS.n704 VSS.n703 2.6005
R4042 VSS.n703 VSS.n702 2.6005
R4043 VSS.n708 VSS.n707 2.6005
R4044 VSS.n707 VSS.n706 2.6005
R4045 VSS.n710 VSS.n709 2.6005
R4046 VSS.n714 VSS.n713 2.6005
R4047 VSS.n716 VSS.n715 2.6005
R4048 VSS.n740 VSS.n739 2.6005
R4049 VSS.n739 VSS.n738 2.6005
R4050 VSS.n737 VSS.n736 2.6005
R4051 VSS.n736 VSS.n735 2.6005
R4052 VSS.n734 VSS.n733 2.6005
R4053 VSS.n733 VSS.n732 2.6005
R4054 VSS.n731 VSS.n730 2.6005
R4055 VSS.n730 VSS.n729 2.6005
R4056 VSS.n728 VSS.n727 2.6005
R4057 VSS.n727 VSS.n726 2.6005
R4058 VSS.n725 VSS.n724 2.6005
R4059 VSS.n724 VSS.n723 2.6005
R4060 VSS.n722 VSS.n721 2.6005
R4061 VSS.n721 VSS.n720 2.6005
R4062 VSS.n719 VSS.n718 2.6005
R4063 VSS.n718 VSS.n717 2.6005
R4064 VSS.n449 VSS.n448 2.6005
R4065 VSS.n448 VSS.n447 2.6005
R4066 VSS.n743 VSS.n742 2.6005
R4067 VSS.n742 VSS.n741 2.6005
R4068 VSS.n1790 VSS.n1789 2.6005
R4069 VSS.n1758 VSS.n1757 2.6005
R4070 VSS.n1757 VSS.n1756 2.6005
R4071 VSS.n1762 VSS.n1761 2.6005
R4072 VSS.n1761 VSS.n1760 2.6005
R4073 VSS.n1765 VSS.n1764 2.6005
R4074 VSS.n1764 VSS.n1763 2.6005
R4075 VSS.n1768 VSS.n1767 2.6005
R4076 VSS.n1767 VSS.n1766 2.6005
R4077 VSS.n1772 VSS.n1771 2.6005
R4078 VSS.n1771 VSS.n1770 2.6005
R4079 VSS.n1775 VSS.n1774 2.6005
R4080 VSS.n1774 VSS.n1773 2.6005
R4081 VSS.n1778 VSS.n1777 2.6005
R4082 VSS.n1777 VSS.n1776 2.6005
R4083 VSS.n1782 VSS.n1781 2.6005
R4084 VSS.n1781 VSS.n1780 2.6005
R4085 VSS.n1785 VSS.n1784 2.6005
R4086 VSS.n1784 VSS.n1783 2.6005
R4087 VSS.n1793 VSS.n1792 2.6005
R4088 VSS.n1792 VSS.n1791 2.6005
R4089 VSS.n1797 VSS.n1796 2.6005
R4090 VSS.n1796 VSS.n1795 2.6005
R4091 VSS.n1801 VSS.n1800 2.6005
R4092 VSS.n1800 VSS.n1799 2.6005
R4093 VSS.n1804 VSS.n1803 2.6005
R4094 VSS.n1803 VSS.n1802 2.6005
R4095 VSS.n1808 VSS.n1807 2.6005
R4096 VSS.n1807 VSS.n1806 2.6005
R4097 VSS.n1815 VSS.n1814 2.6005
R4098 VSS.n1814 VSS.n1813 2.6005
R4099 VSS.n1818 VSS.n1817 2.6005
R4100 VSS.n1817 VSS.n1816 2.6005
R4101 VSS.n1823 VSS.n1822 2.6005
R4102 VSS.n1822 VSS.n1821 2.6005
R4103 VSS.n1826 VSS.n1825 2.6005
R4104 VSS.n1825 VSS.n1824 2.6005
R4105 VSS.n2071 VSS.n2070 2.6005
R4106 VSS.n2073 VSS.n2072 2.6005
R4107 VSS.n2075 VSS.n2074 2.6005
R4108 VSS.n2077 VSS.n2076 2.6005
R4109 VSS.n2079 VSS.n2078 2.6005
R4110 VSS.n2081 VSS.n2080 2.6005
R4111 VSS.n2083 VSS.n2082 2.6005
R4112 VSS.n2085 VSS.n2084 2.6005
R4113 VSS.n2087 VSS.n2086 2.6005
R4114 VSS.n2089 VSS.n2088 2.6005
R4115 VSS.n184 VSS.n183 2.6005
R4116 VSS.n183 VSS.n182 2.6005
R4117 VSS.n187 VSS.n186 2.6005
R4118 VSS.n186 VSS.n185 2.6005
R4119 VSS.n190 VSS.n189 2.6005
R4120 VSS.n189 VSS.n188 2.6005
R4121 VSS.n193 VSS.n192 2.6005
R4122 VSS.n192 VSS.n191 2.6005
R4123 VSS.n196 VSS.n195 2.6005
R4124 VSS.n195 VSS.n194 2.6005
R4125 VSS.n200 VSS.n199 2.6005
R4126 VSS.n199 VSS.n198 2.6005
R4127 VSS.n2064 VSS.n2063 2.6005
R4128 VSS.n2061 VSS.n2060 2.6005
R4129 VSS.n1639 VSS.n1638 2.6005
R4130 VSS.n1642 VSS.n1641 2.6005
R4131 VSS.n1645 VSS.n1644 2.6005
R4132 VSS.n1648 VSS.n1647 2.6005
R4133 VSS.n1651 VSS.n1650 2.6005
R4134 VSS.n1655 VSS.n1654 2.6005
R4135 VSS.n2066 VSS.n2065 2.6005
R4136 VSS.n2058 VSS.n2057 2.6005
R4137 VSS.n2055 VSS.n2054 2.6005
R4138 VSS.n2053 VSS.n2052 2.6005
R4139 VSS.n143 VSS.n142 2.6005
R4140 VSS.n145 VSS.n144 2.6005
R4141 VSS.n159 VSS.n158 2.6005
R4142 VSS.n162 VSS.n161 2.6005
R4143 VSS.n1497 VSS.n1496 2.6005
R4144 VSS.n1495 VSS.n1494 2.6005
R4145 VSS.n1493 VSS.n1492 2.6005
R4146 VSS.n1491 VSS.n1490 2.6005
R4147 VSS.n1489 VSS.n1488 2.6005
R4148 VSS.n1487 VSS.n1486 2.6005
R4149 VSS.n1485 VSS.n1484 2.6005
R4150 VSS.n1499 VSS.n1498 2.6005
R4151 VSS.n1478 VSS.n1477 2.6005
R4152 VSS.n1475 VSS.n1474 2.6005
R4153 VSS.n1547 VSS.n1546 2.6005
R4154 VSS.n1549 VSS.n1548 2.6005
R4155 VSS.n1551 VSS.n1550 2.6005
R4156 VSS.n1553 VSS.n1552 2.6005
R4157 VSS.n1042 VSS.n1041 2.6005
R4158 VSS.n1040 VSS.n1039 2.6005
R4159 VSS.n1037 VSS.n1036 2.6005
R4160 VSS.n1035 VSS.n1034 2.6005
R4161 VSS.n1031 VSS.n1030 2.6005
R4162 VSS.n1029 VSS.n1028 2.6005
R4163 VSS.n1659 VSS.n1658 2.6005
R4164 VSS.n1658 VSS.n1657 2.6005
R4165 VSS.n1662 VSS.n1661 2.6005
R4166 VSS.n1661 VSS.n1660 2.6005
R4167 VSS.n1665 VSS.n1664 2.6005
R4168 VSS.n1664 VSS.n1663 2.6005
R4169 VSS.n1668 VSS.n1667 2.6005
R4170 VSS.n1667 VSS.n1666 2.6005
R4171 VSS.n1671 VSS.n1670 2.6005
R4172 VSS.n1670 VSS.n1669 2.6005
R4173 VSS.n1674 VSS.n1673 2.6005
R4174 VSS.n1673 VSS.n1672 2.6005
R4175 VSS.n1676 VSS.n1675 2.6005
R4176 VSS.n1675 VSS.t119 2.6005
R4177 VSS.n1679 VSS.n1678 2.6005
R4178 VSS.n1678 VSS.n1677 2.6005
R4179 VSS.n1682 VSS.n1681 2.6005
R4180 VSS.n1681 VSS.n1680 2.6005
R4181 VSS.n1685 VSS.n1684 2.6005
R4182 VSS.n1684 VSS.n1683 2.6005
R4183 VSS.n1688 VSS.n1687 2.6005
R4184 VSS.n1687 VSS.n1686 2.6005
R4185 VSS.n1691 VSS.n1690 2.6005
R4186 VSS.n1690 VSS.n1689 2.6005
R4187 VSS.n1694 VSS.n1693 2.6005
R4188 VSS.n1693 VSS.n1692 2.6005
R4189 VSS.n1697 VSS.n1696 2.6005
R4190 VSS.n1696 VSS.n1695 2.6005
R4191 VSS.n1700 VSS.n1699 2.6005
R4192 VSS.n1699 VSS.n1698 2.6005
R4193 VSS.n1703 VSS.n1702 2.6005
R4194 VSS.n1702 VSS.n1701 2.6005
R4195 VSS.n1502 VSS.n1501 2.6005
R4196 VSS.n1504 VSS.n1503 2.6005
R4197 VSS.n1506 VSS.n1505 2.6005
R4198 VSS.n1508 VSS.n1507 2.6005
R4199 VSS.n1510 VSS.n1509 2.6005
R4200 VSS.n1512 VSS.n1511 2.6005
R4201 VSS.n1514 VSS.n1513 2.6005
R4202 VSS.n1516 VSS.n1515 2.6005
R4203 VSS.n1518 VSS.n1517 2.6005
R4204 VSS.n1520 VSS.n1519 2.6005
R4205 VSS.n1522 VSS.n1521 2.6005
R4206 VSS.n1524 VSS.n1523 2.6005
R4207 VSS.n1526 VSS.n1525 2.6005
R4208 VSS.n1528 VSS.n1527 2.6005
R4209 VSS.n1530 VSS.n1529 2.6005
R4210 VSS.n1532 VSS.n1531 2.6005
R4211 VSS.n1559 VSS.n1558 2.6005
R4212 VSS.n1558 VSS.n1557 2.6005
R4213 VSS.n1562 VSS.n1561 2.6005
R4214 VSS.n1561 VSS.n1560 2.6005
R4215 VSS.n1565 VSS.n1564 2.6005
R4216 VSS.n1564 VSS.n1563 2.6005
R4217 VSS.n1568 VSS.n1567 2.6005
R4218 VSS.n1567 VSS.n1566 2.6005
R4219 VSS.n1571 VSS.n1570 2.6005
R4220 VSS.n1570 VSS.n1569 2.6005
R4221 VSS.n1574 VSS.n1573 2.6005
R4222 VSS.n1573 VSS.n1572 2.6005
R4223 VSS.n1577 VSS.n1576 2.6005
R4224 VSS.n1576 VSS.n1575 2.6005
R4225 VSS.n1580 VSS.n1579 2.6005
R4226 VSS.n1579 VSS.n1578 2.6005
R4227 VSS.n1583 VSS.n1582 2.6005
R4228 VSS.n1582 VSS.n1581 2.6005
R4229 VSS.n1586 VSS.n1585 2.6005
R4230 VSS.n1585 VSS.n1584 2.6005
R4231 VSS.n1589 VSS.n1588 2.6005
R4232 VSS.n1588 VSS.n1587 2.6005
R4233 VSS.n1592 VSS.n1591 2.6005
R4234 VSS.n1591 VSS.n1590 2.6005
R4235 VSS.n1595 VSS.n1594 2.6005
R4236 VSS.n1594 VSS.n1593 2.6005
R4237 VSS.n1598 VSS.n1597 2.6005
R4238 VSS.n1597 VSS.n1596 2.6005
R4239 VSS.n1601 VSS.n1600 2.6005
R4240 VSS.n1600 VSS.n1599 2.6005
R4241 VSS.n1604 VSS.n1603 2.6005
R4242 VSS.n1603 VSS.n1602 2.6005
R4243 VSS.n1540 VSS.n1539 2.6005
R4244 VSS.n1542 VSS.n1541 2.6005
R4245 VSS.n1545 VSS.n1544 2.6005
R4246 VSS.n1752 VSS.n1751 2.6005
R4247 VSS.n483 VSS.n482 2.6005
R4248 VSS.n1615 VSS.n1614 2.6005
R4249 VSS.n1617 VSS.n1616 2.6005
R4250 VSS.n1620 VSS.n1619 2.6005
R4251 VSS.n1622 VSS.n1621 2.6005
R4252 VSS.n1625 VSS.n1624 2.6005
R4253 VSS.n1627 VSS.n1626 2.6005
R4254 VSS.n1630 VSS.n1629 2.6005
R4255 VSS.n1632 VSS.n1631 2.6005
R4256 VSS.n1635 VSS.n1634 2.6005
R4257 VSS.n1637 VSS.n1636 2.6005
R4258 VSS.n1732 VSS.n1731 2.6005
R4259 VSS.n1734 VSS.n1733 2.6005
R4260 VSS.n1737 VSS.n1736 2.6005
R4261 VSS.n1740 VSS.n1739 2.6005
R4262 VSS.n1743 VSS.n1742 2.6005
R4263 VSS.n1746 VSS.n1745 2.6005
R4264 VSS.n1705 VSS.n1704 2.6005
R4265 VSS.n1726 VSS.n1725 2.6005
R4266 VSS.n1729 VSS.n1728 2.6005
R4267 VSS.n1610 VSS.n1609 2.6005
R4268 VSS.n1608 VSS.n1607 2.6005
R4269 VSS.n1538 VSS.n1537 2.6005
R4270 VSS.n1535 VSS.n1534 2.6005
R4271 VSS.n556 VSS.n555 2.6005
R4272 VSS.n1011 VSS.n1010 2.6005
R4273 VSS.n1013 VSS.n1012 2.6005
R4274 VSS.n1015 VSS.n1014 2.6005
R4275 VSS.n1017 VSS.n1016 2.6005
R4276 VSS.n1019 VSS.n1018 2.6005
R4277 VSS.n1026 VSS.n1025 2.6005
R4278 VSS.n1024 VSS.n1023 2.6005
R4279 VSS.n1022 VSS.n1021 2.6005
R4280 VSS.n1606 VSS.n1605 2.6005
R4281 VSS.n2110 VSS.n2109 2.6005
R4282 VSS.n2112 VSS.n2111 2.6005
R4283 VSS.n2117 VSS.n2116 2.6005
R4284 VSS.n2121 VSS.n2120 2.6005
R4285 VSS.n2123 VSS.n2122 2.6005
R4286 VSS.n2107 VSS.n2106 2.6005
R4287 VSS.n2091 VSS.n2090 2.6005
R4288 VSS.n2093 VSS.n2092 2.6005
R4289 VSS.n2095 VSS.n2094 2.6005
R4290 VSS.n2097 VSS.n2096 2.6005
R4291 VSS.n2099 VSS.n2098 2.6005
R4292 VSS.n2101 VSS.n2100 2.6005
R4293 VSS.n2104 VSS.n2103 2.6005
R4294 VSS.n2145 VSS.n2144 2.6005
R4295 VSS.n2146 VSS.n2145 2.6005
R4296 VSS.n2143 VSS.n2142 2.6005
R4297 VSS.n2142 VSS.n2141 2.6005
R4298 VSS.n2140 VSS.n2139 2.6005
R4299 VSS.n2139 VSS.n2138 2.6005
R4300 VSS.n2137 VSS.n2136 2.6005
R4301 VSS.n2136 VSS.n2135 2.6005
R4302 VSS.n2133 VSS.n2132 2.6005
R4303 VSS.n2132 VSS.n2131 2.6005
R4304 VSS.n2130 VSS.n2129 2.6005
R4305 VSS.n2129 VSS.n2128 2.6005
R4306 VSS.n2127 VSS.n2126 2.6005
R4307 VSS.n2126 VSS.n2125 2.6005
R4308 VSS.n2060 VSS.n2059 2.58211
R4309 VSS.n1647 VSS.n1646 2.58211
R4310 VSS.n1644 VSS.n1643 2.58211
R4311 VSS.n1641 VSS.n1640 2.58211
R4312 VSS.n1745 VSS.n1744 2.58211
R4313 VSS.n1742 VSS.n1741 2.58211
R4314 VSS.n1739 VSS.n1738 2.58211
R4315 VSS.n1736 VSS.n1735 2.58211
R4316 VSS.n1972 VSS.t191 2.56713
R4317 VSS.t102 VSS.n146 2.54175
R4318 VSS.t516 VSS.t158 2.52772
R4319 VSS.n1147 VSS.n1146 2.52772
R4320 VSS.t468 VSS.t474 2.52772
R4321 VSS.n1132 VSS.n1093 2.51205
R4322 VSS.n1003 VSS.t93 2.41865
R4323 VSS.n1051 VSS.n1050 2.41865
R4324 VSS.n2191 VSS 2.40845
R4325 VSS.n1131 VSS.n1130 2.37524
R4326 VSS.t266 VSS.t264 2.3693
R4327 VSS.n1085 VSS.n1084 2.3693
R4328 VSS.t252 VSS.t229 2.3693
R4329 VSS.n1421 VSS.n1420 2.32691
R4330 VSS.n2408 VSS.t383 2.25486
R4331 VSS.n2409 VSS.t403 2.25486
R4332 VSS.n2410 VSS.t410 2.25486
R4333 VSS.n2411 VSS.t433 2.25486
R4334 VSS.n2412 VSS.t378 2.25486
R4335 VSS.n2413 VSS.t418 2.25486
R4336 VSS.n2414 VSS.t409 2.25486
R4337 VSS.n2401 VSS.t382 2.25486
R4338 VSS.n2402 VSS.t402 2.25486
R4339 VSS.n2403 VSS.t405 2.25486
R4340 VSS.n2404 VSS.t432 2.25486
R4341 VSS.n2405 VSS.t377 2.25486
R4342 VSS.n2406 VSS.t371 2.25486
R4343 VSS.n2407 VSS.t424 2.25486
R4344 VSS.n2394 VSS.t399 2.25486
R4345 VSS.n2395 VSS.t423 2.25486
R4346 VSS.n2396 VSS.t430 2.25486
R4347 VSS.n2397 VSS.t388 2.25486
R4348 VSS.n2398 VSS.t393 2.25486
R4349 VSS.n2399 VSS.t414 2.25486
R4350 VSS.n2400 VSS.t401 2.25486
R4351 VSS.n2387 VSS.t370 2.25486
R4352 VSS.n2388 VSS.t395 2.25486
R4353 VSS.n2389 VSS.t398 2.25486
R4354 VSS.n2390 VSS.t421 2.25486
R4355 VSS.n2391 VSS.t429 2.25486
R4356 VSS.n2392 VSS.t373 2.25486
R4357 VSS.n2393 VSS.t428 2.25486
R4358 VSS.n2418 VSS.t386 2.25486
R4359 VSS.n2419 VSS.t408 2.25486
R4360 VSS.n2420 VSS.t416 2.25486
R4361 VSS.n2421 VSS.t375 2.25486
R4362 VSS.n2422 VSS.t381 2.25486
R4363 VSS.n2423 VSS.t372 2.25486
R4364 VSS.n2424 VSS.t425 2.25486
R4365 VSS.n2425 VSS.t379 2.25486
R4366 VSS.n2426 VSS.t400 2.25486
R4367 VSS.n2427 VSS.t404 2.25486
R4368 VSS.n2428 VSS.t431 2.25486
R4369 VSS.n2429 VSS.t376 2.25486
R4370 VSS.n2430 VSS.t419 2.25486
R4371 VSS.n2431 VSS.t411 2.25486
R4372 VSS.n2432 VSS.t397 2.25486
R4373 VSS.n2433 VSS.t422 2.25486
R4374 VSS.n2434 VSS.t427 2.25486
R4375 VSS.n2435 VSS.t387 2.25486
R4376 VSS.n2436 VSS.t391 2.25486
R4377 VSS.n2437 VSS.t420 2.25486
R4378 VSS.n2438 VSS.t412 2.25486
R4379 VSS.n2439 VSS.t385 2.25486
R4380 VSS.n2440 VSS.t407 2.25486
R4381 VSS.n2441 VSS.t415 2.25486
R4382 VSS.n2442 VSS.t374 2.25486
R4383 VSS.n2443 VSS.t380 2.25486
R4384 VSS.n2444 VSS.t426 2.25486
R4385 VSS.n2445 VSS.t417 2.25486
R4386 VSS.n1140 VSS.n1139 2.24529
R4387 VSS.n1138 VSS.n1137 2.24398
R4388 VSS.n123 VSS.n122 2.13762
R4389 VSS.t68 VSS.t208 2.08117
R4390 VSS.n1077 VSS.n1074 2.08117
R4391 VSS.t517 VSS.t157 2.08117
R4392 VSS.t152 VSS.t541 2.08117
R4393 VSS.n1081 VSS.n1080 2.08117
R4394 VSS.t273 VSS.t361 2.08117
R4395 VSS.n112 VSS 2.03762
R4396 VSS.n1170 VSS.n1169 1.9795
R4397 VSS.n232 VSS.n231 1.90645
R4398 VSS.n343 VSS.n342 1.90327
R4399 VSS.n237 VSS.n236 1.90327
R4400 VSS.n1130 VSS.n1104 1.80706
R4401 VSS.n1398 VSS.n1397 1.79328
R4402 VSS.n1415 VSS.n1414 1.7776
R4403 VSS.n1383 VSS.n1382 1.77751
R4404 VSS.n227 VSS.n226 1.74691
R4405 VSS.n1315 VSS.n1314 1.72783
R4406 VSS.n859 VSS.n852 1.7266
R4407 VSS.n1122 VSS.n1121 1.7266
R4408 VSS.n1112 VSS.n1111 1.7266
R4409 VSS.n2057 VSS.n2056 1.7266
R4410 VSS.n2109 VSS.n2108 1.7266
R4411 VSS.n2120 VSS.n2119 1.7266
R4412 VSS.n1044 VSS.n1043 1.72602
R4413 VSS.n859 VSS.n858 1.72602
R4414 VSS.n142 VSS.n141 1.72602
R4415 VSS.n158 VSS.n157 1.72602
R4416 VSS.n1039 VSS.n1038 1.72602
R4417 VSS.n1034 VSS.n1033 1.72602
R4418 VSS.n1028 VSS.n1027 1.72602
R4419 VSS.n2116 VSS.n2115 1.72602
R4420 VSS.n1998 VSS.n1997 1.72592
R4421 VSS.n870 VSS.n869 1.72592
R4422 VSS.n875 VSS.n874 1.72592
R4423 VSS.n1341 VSS.n1340 1.69507
R4424 VSS.n1255 VSS.n1254 1.69507
R4425 VSS.n1261 VSS.n1260 1.69507
R4426 VSS.n1249 VSS.n1248 1.69497
R4427 VSS.n2031 VSS.n2030 1.68203
R4428 VSS.n332 VSS.n331 1.68193
R4429 VSS.n337 VSS.n336 1.68193
R4430 VSS.n2039 VSS.n2038 1.68193
R4431 VSS.n326 VSS.n325 1.67823
R4432 VSS.n2047 VSS.t118 1.6385
R4433 VSS.n2047 VSS.n2046 1.6385
R4434 VSS.n2045 VSS.t646 1.6385
R4435 VSS.n2045 VSS.n2044 1.6385
R4436 VSS.n203 VSS.t188 1.6385
R4437 VSS.n203 VSS.n202 1.6385
R4438 VSS.n329 VSS.t663 1.6385
R4439 VSS.n329 VSS.n328 1.6385
R4440 VSS.n1933 VSS.t642 1.6385
R4441 VSS.n1933 VSS.n1932 1.6385
R4442 VSS.n1931 VSS.t126 1.6385
R4443 VSS.n1931 VSS.n1930 1.6385
R4444 VSS.n755 VSS.t122 1.6385
R4445 VSS.n755 VSS.n754 1.6385
R4446 VSS.n753 VSS.t645 1.6385
R4447 VSS.n753 VSS.n752 1.6385
R4448 VSS.n550 VSS.t604 1.6385
R4449 VSS.n550 VSS.n549 1.6385
R4450 VSS.n548 VSS.t120 1.6385
R4451 VSS.n548 VSS.n547 1.6385
R4452 VSS.n593 VSS.t42 1.6385
R4453 VSS.n593 VSS.n592 1.6385
R4454 VSS.n584 VSS.t339 1.6385
R4455 VSS.n584 VSS.n583 1.6385
R4456 VSS.n2415 VSS.n2414 1.63171
R4457 VSS.n2446 VSS.n2445 1.6308
R4458 VSS.n478 VSS.n477 1.62689
R4459 VSS.n1624 VSS.n1623 1.62622
R4460 VSS.n1629 VSS.n1628 1.62622
R4461 VSS.n1634 VSS.n1633 1.62622
R4462 VSS.n950 VSS.n949 1.55471
R4463 VSS.n1407 VSS.n1406 1.55166
R4464 VSS.n1401 VSS.n1400 1.55155
R4465 VSS.n488 VSS.n487 1.53476
R4466 VSS.n713 VSS.n712 1.53476
R4467 VSS.n937 VSS.n936 1.53464
R4468 VSS.n943 VSS.n942 1.53464
R4469 VSS.n1725 VSS.n1724 1.53235
R4470 VSS.t208 VSS.n1073 1.51003
R4471 VSS.n900 VSS.n899 1.50472
R4472 VSS.n311 VSS.n310 1.50072
R4473 VSS.n2453 VSS.n2452 1.5005
R4474 VSS.n1229 VSS.n1228 1.4928
R4475 VSS.n985 VSS.n904 1.48535
R4476 VSS.n286 VSS.n285 1.47758
R4477 VSS.n1650 VSS.n1649 1.47758
R4478 VSS.n1728 VSS.n1727 1.47758
R4479 VSS.n281 VSS.n280 1.47745
R4480 VSS.n1731 VSS.n1730 1.47745
R4481 VSS.n2063 VSS.n2062 1.47745
R4482 VSS VSS.n2051 1.46704
R4483 VSS VSS.n1937 1.46704
R4484 VSS VSS.n759 1.46704
R4485 VSS VSS.n554 1.46704
R4486 VSS.n1377 VSS.n1376 1.45083
R4487 VSS.n934 VSS.n933 1.45083
R4488 VSS.n1344 VSS.n1343 1.44361
R4489 VSS.n1350 VSS.n1349 1.44361
R4490 VSS.n1806 VSS.t304 1.43517
R4491 VSS.t150 VSS.n569 1.41853
R4492 VSS.n904 VSS.n888 1.37929
R4493 VSS.n536 VSS.n535 1.36965
R4494 VSS.n542 VSS.n541 1.36965
R4495 VSS.n1614 VSS.n1613 1.36965
R4496 VSS.n1619 VSS.n1618 1.36965
R4497 VSS.n1437 VSS.t539 1.32475
R4498 VSS.n156 VSS.n151 1.31044
R4499 VSS.n156 VSS.n152 1.31044
R4500 VSS.n156 VSS.n153 1.31044
R4501 VSS.n156 VSS.n154 1.31044
R4502 VSS.n1723 VSS.n1717 1.31044
R4503 VSS.n1723 VSS.n1718 1.31044
R4504 VSS.n1723 VSS.n1719 1.31044
R4505 VSS.n1723 VSS.n1720 1.31044
R4506 VSS.n1751 VSS.n1750 1.28563
R4507 VSS.n1789 VSS.n1788 1.28498
R4508 VSS.n1223 VSS.n1222 1.25894
R4509 VSS.n545 VSS.t28 1.1705
R4510 VSS.n545 VSS.n544 1.1705
R4511 VSS.n451 VSS.t301 1.1705
R4512 VSS.n451 VSS.n450 1.1705
R4513 VSS.n1103 VSS.n1102 1.15416
R4514 VSS.n1770 VSS.t29 1.13028
R4515 VSS.n2457 VSS.n2456 1.1247
R4516 VSS.n382 VSS 1.09141
R4517 VSS.n2417 VSS.n2416 1.07514
R4518 VSS.n2448 VSS.n2447 1.07514
R4519 VSS.n2416 VSS.n2415 1.07476
R4520 VSS.n2447 VSS.n2446 1.07438
R4521 VSS.n2315 VSS.n2314 1.03389
R4522 VSS.n2124 VSS 1.03013
R4523 VSS.n2458 VSS 1.0234
R4524 VSS.n2409 VSS.n2408 1.01182
R4525 VSS.n2410 VSS.n2409 1.01182
R4526 VSS.n2411 VSS.n2410 1.01182
R4527 VSS.n2412 VSS.n2411 1.01182
R4528 VSS.n2413 VSS.n2412 1.01182
R4529 VSS.n2414 VSS.n2413 1.01182
R4530 VSS.n2402 VSS.n2401 1.01182
R4531 VSS.n2403 VSS.n2402 1.01182
R4532 VSS.n2404 VSS.n2403 1.01182
R4533 VSS.n2405 VSS.n2404 1.01182
R4534 VSS.n2406 VSS.n2405 1.01182
R4535 VSS.n2407 VSS.n2406 1.01182
R4536 VSS.n2395 VSS.n2394 1.01182
R4537 VSS.n2396 VSS.n2395 1.01182
R4538 VSS.n2397 VSS.n2396 1.01182
R4539 VSS.n2398 VSS.n2397 1.01182
R4540 VSS.n2399 VSS.n2398 1.01182
R4541 VSS.n2400 VSS.n2399 1.01182
R4542 VSS.n2388 VSS.n2387 1.01182
R4543 VSS.n2389 VSS.n2388 1.01182
R4544 VSS.n2390 VSS.n2389 1.01182
R4545 VSS.n2391 VSS.n2390 1.01182
R4546 VSS.n2392 VSS.n2391 1.01182
R4547 VSS.n2393 VSS.n2392 1.01182
R4548 VSS.n2419 VSS.n2418 1.01182
R4549 VSS.n2420 VSS.n2419 1.01182
R4550 VSS.n2421 VSS.n2420 1.01182
R4551 VSS.n2422 VSS.n2421 1.01182
R4552 VSS.n2423 VSS.n2422 1.01182
R4553 VSS.n2424 VSS.n2423 1.01182
R4554 VSS.n2426 VSS.n2425 1.01182
R4555 VSS.n2427 VSS.n2426 1.01182
R4556 VSS.n2428 VSS.n2427 1.01182
R4557 VSS.n2429 VSS.n2428 1.01182
R4558 VSS.n2430 VSS.n2429 1.01182
R4559 VSS.n2431 VSS.n2430 1.01182
R4560 VSS.n2433 VSS.n2432 1.01182
R4561 VSS.n2434 VSS.n2433 1.01182
R4562 VSS.n2435 VSS.n2434 1.01182
R4563 VSS.n2436 VSS.n2435 1.01182
R4564 VSS.n2437 VSS.n2436 1.01182
R4565 VSS.n2438 VSS.n2437 1.01182
R4566 VSS.n2440 VSS.n2439 1.01182
R4567 VSS.n2441 VSS.n2440 1.01182
R4568 VSS.n2442 VSS.n2441 1.01182
R4569 VSS.n2443 VSS.n2442 1.01182
R4570 VSS.n2444 VSS.n2443 1.01182
R4571 VSS.n2445 VSS.n2444 1.01182
R4572 VSS.n121 VSS.n48 1.00481
R4573 VSS.n324 VSS.t300 0.956945
R4574 VSS.n2381 VSS.n2379 0.939556
R4575 VSS.n2118 VSS.n2043 0.938847
R4576 VSS.n2279 VSS 0.930989
R4577 VSS.n1847 VSS.n417 0.929805
R4578 VSS.n2003 VSS.n2002 0.91886
R4579 VSS.n2451 VSS.n2450 0.898925
R4580 VSS.t271 VSS.n2365 0.878785
R4581 VSS.n1723 VSS.n1711 0.847406
R4582 VSS.n1749 VSS.n1748 0.847406
R4583 VSS.n2254 VSS.n2253 0.846463
R4584 VSS.n2233 VSS.n2232 0.846463
R4585 VSS.n77 VSS.n76 0.846463
R4586 VSS.n2050 VSS.n2049 0.845717
R4587 VSS.n1936 VSS.n1935 0.845717
R4588 VSS.n758 VSS.n757 0.845717
R4589 VSS.n553 VSS.n552 0.845717
R4590 VSS.n2350 VSS.n21 0.843955
R4591 VSS VSS.n882 0.841511
R4592 VSS VSS.n1082 0.840934
R4593 VSS.n2051 VSS.n2050 0.827256
R4594 VSS.n1937 VSS.n1936 0.827256
R4595 VSS.n759 VSS.n758 0.827256
R4596 VSS.n554 VSS.n553 0.827256
R4597 VSS.n541 VSS.n540 0.8219
R4598 VSS.n1349 VSS.n1348 0.772592
R4599 VSS.n247 VSS 0.765857
R4600 VSS.n2459 VSS.n2458 0.75996
R4601 VSS.n156 VSS.n155 0.750234
R4602 VSS.n1723 VSS.n1721 0.750234
R4603 VSS.n156 VSS.n150 0.75003
R4604 VSS.n1723 VSS.n1716 0.75003
R4605 VSS.n1228 VSS.n1227 0.739798
R4606 VSS.n2337 VSS.n33 0.73944
R4607 VSS.n2450 VSS.n2449 0.71213
R4608 VSS.n1406 VSS.n1405 0.700841
R4609 VSS VSS.n130 0.676801
R4610 VSS.n1750 VSS.n1749 0.659244
R4611 VSS.n1788 VSS.n1787 0.65901
R4612 VSS.n2460 VSS.n2382 0.649205
R4613 VSS.n2458 VSS 0.647475
R4614 VSS.n2280 VSS.n2279 0.645242
R4615 VSS.n112 VSS.n111 0.616742
R4616 VSS.n325 VSS.n324 0.616183
R4617 VSS.n1409 VSS.n1374 0.606056
R4618 VSS.n2324 VSS.n2175 0.605183
R4619 VSS.n1376 VSS.n1375 0.576657
R4620 VSS.n933 VSS.n932 0.576657
R4621 VSS.n2415 VSS.n2407 0.556878
R4622 VSS.n2416 VSS.n2400 0.556878
R4623 VSS.n2417 VSS.n2393 0.556878
R4624 VSS.n2448 VSS.n2424 0.556878
R4625 VSS.n2447 VSS.n2431 0.556878
R4626 VSS.n2446 VSS.n2438 0.556878
R4627 VSS.n1083 VSS 0.545498
R4628 VSS VSS.n1086 0.545498
R4629 VSS.n2449 VSS.n2417 0.539639
R4630 VSS.n1724 VSS.n1723 0.535627
R4631 VSS.n1723 VSS.n1722 0.535627
R4632 VSS.n2449 VSS.n2448 0.53562
R4633 VSS.n487 VSS.n486 0.53442
R4634 VSS.n712 VSS.n711 0.53442
R4635 VSS.n949 VSS.n948 0.52472
R4636 VSS.n1358 VSS.n1357 0.5185
R4637 VSS.n420 VSS.n418 0.5005
R4638 VSS.n1655 VSS.n1652 0.5005
R4639 VSS.n861 VSS.n860 0.5005
R4640 VSS.n1482 VSS.n1481 0.5005
R4641 VSS.n120 VSS.n114 0.486611
R4642 VSS.n2317 VSS.n2316 0.480225
R4643 VSS.n1062 VSS.n1053 0.467323
R4644 VSS.n1340 VSS.n1339 0.454258
R4645 VSS.n1260 VSS.n1259 0.454258
R4646 VSS.n136 VSS.n135 0.439554
R4647 VSS VSS.n32 0.43894
R4648 VSS.n1166 VSS.n859 0.438783
R4649 VSS.n1121 VSS.n1120 0.438783
R4650 VSS.n157 VSS.n156 0.438783
R4651 VSS.n1033 VSS.n1032 0.438783
R4652 VSS.n1723 VSS.n1714 0.438783
R4653 VSS.n1723 VSS.n1713 0.438783
R4654 VSS.n1723 VSS.n1715 0.438783
R4655 VSS.n2115 VSS.n2114 0.438783
R4656 VSS.n1997 VSS.n1996 0.43854
R4657 VSS.n869 VSS.n868 0.43854
R4658 VSS.n156 VSS.n149 0.43854
R4659 VSS.n156 VSS.n148 0.43854
R4660 VSS.n156 VSS.n147 0.43854
R4661 VSS.n1314 VSS.n1313 0.438169
R4662 VSS.n1414 VSS.n1413 0.412988
R4663 VSS.n1382 VSS.n1381 0.412744
R4664 VSS.n2211 VSS.n2210 0.395692
R4665 VSS.n2208 VSS.n2206 0.395692
R4666 VSS.n2203 VSS.n2202 0.395692
R4667 VSS.n370 VSS.n355 0.382171
R4668 VSS.n2192 VSS 0.378121
R4669 VSS.n390 VSS.n389 0.377093
R4670 VSS.n77 VSS.n22 0.35472
R4671 VSS.n342 VSS.n341 0.349863
R4672 VSS.n1143 VSS.n1142 0.349591
R4673 VSS.n79 VSS.n19 0.348115
R4674 VSS VSS.n2302 0.343161
R4675 VSS.n2303 VSS 0.343161
R4676 VSS VSS.n2240 0.343161
R4677 VSS.n2241 VSS 0.343161
R4678 VSS VSS.n2219 0.343161
R4679 VSS.n2220 VSS 0.343161
R4680 VSS.n87 VSS 0.343161
R4681 VSS.n2260 VSS 0.343161
R4682 VSS VSS.n69 0.343161
R4683 VSS VSS.n71 0.343161
R4684 VSS.n363 VSS.n360 0.338437
R4685 VSS.n1142 VSS.n1141 0.325955
R4686 VSS.n17 VSS.n14 0.325821
R4687 VSS.n134 VSS.n133 0.316175
R4688 VSS.n28 VSS.n25 0.313436
R4689 VSS VSS.n137 0.311851
R4690 VSS VSS.n2197 0.310668
R4691 VSS.n1247 VSS.n1246 0.304848
R4692 VSS.n1177 VSS.n846 0.304848
R4693 VSS.n2319 VSS.n2318 0.294445
R4694 VSS.n2309 VSS 0.289491
R4695 VSS.n2248 VSS 0.289491
R4696 VSS.n2227 VSS 0.289491
R4697 VSS.n74 VSS 0.289491
R4698 VSS.n2273 VSS.n2178 0.286539
R4699 VSS.n2207 VSS 0.27984
R4700 VSS VSS.n2204 0.27984
R4701 VSS.n1446 VSS 0.278241
R4702 VSS.n364 VSS.n0 0.277931
R4703 VSS.n363 VSS.n362 0.272151
R4704 VSS.n2230 VSS.n30 0.268849
R4705 VSS.n2279 VSS.n2278 0.262771
R4706 VSS VSS.n94 0.261689
R4707 VSS VSS.n96 0.261689
R4708 VSS VSS.n2265 0.259875
R4709 VSS VSS.n2267 0.259875
R4710 VSS.n2460 VSS.n2459 0.258628
R4711 VSS.n2163 VSS 0.258086
R4712 VSS VSS.n2168 0.258086
R4713 VSS.n1443 VSS 0.256849
R4714 VSS.n1063 VSS.n1062 0.255428
R4715 VSS.n54 VSS 0.254582
R4716 VSS VSS.n59 0.254582
R4717 VSS.n2251 VSS.n45 0.252335
R4718 VSS.n40 VSS.n39 0.250683
R4719 VSS.n246 VSS.n241 0.2505
R4720 VSS.n162 VSS.n160 0.2505
R4721 VSS.n751 VSS.n749 0.2505
R4722 VSS.n1555 VSS.n1554 0.2505
R4723 VSS VSS.n2200 0.250123
R4724 VSS.n2200 VSS.n2199 0.247195
R4725 VSS VSS.n2207 0.243604
R4726 VSS.n2204 VSS 0.243604
R4727 VSS VSS.n9 0.240775
R4728 VSS VSS.n35 0.23417
R4729 VSS.n43 VSS.n40 0.230041
R4730 VSS.n45 VSS.n44 0.22839
R4731 VSS.n2113 VSS 0.224346
R4732 VSS.n1938 VSS 0.224346
R4733 VSS.n760 VSS 0.224346
R4734 VSS.n1543 VSS 0.224346
R4735 VSS VSS.n139 0.223676
R4736 VSS VSS.n99 0.22078
R4737 VSS VSS.n1438 0.22033
R4738 VSS.n2282 VSS 0.21925
R4739 VSS.n2173 VSS 0.217741
R4740 VSS.n64 VSS 0.214786
R4741 VSS.n30 VSS.n29 0.211876
R4742 VSS.n1447 VSS.n595 0.206733
R4743 VSS.n2253 VSS.n47 0.201142
R4744 VSS.n2337 VSS 0.192251
R4745 VSS VSS.n2308 0.191234
R4746 VSS VSS.n2246 0.191234
R4747 VSS VSS.n2225 0.191234
R4748 VSS VSS.n73 0.191234
R4749 VSS.n78 VSS.n77 0.187931
R4750 VSS.n2232 VSS.n2231 0.187931
R4751 VSS.n2253 VSS.n2252 0.187931
R4752 VSS.n379 VSS.n350 0.187704
R4753 VSS.n2319 VSS.n2179 0.18628
R4754 VSS.n1169 VSS.n1168 0.185
R4755 VSS.n385 VSS.n384 0.184546
R4756 VSS.n335 VSS.n333 0.183918
R4757 VSS.n338 VSS.n335 0.183918
R4758 VSS.n340 VSS.n338 0.183918
R4759 VSS.n317 VSS.n314 0.183918
R4760 VSS.n320 VSS.n317 0.183918
R4761 VSS.n323 VSS.n320 0.183918
R4762 VSS.n230 VSS.n228 0.183918
R4763 VSS.n233 VSS.n230 0.183918
R4764 VSS.n235 VSS.n233 0.183918
R4765 VSS.n2034 VSS.n2032 0.183918
R4766 VSS.n2037 VSS.n2034 0.183918
R4767 VSS.n2040 VSS.n2037 0.183918
R4768 VSS.n344 VSS.n340 0.182778
R4769 VSS.n327 VSS.n323 0.182778
R4770 VSS.n238 VSS.n235 0.182778
R4771 VSS.n2042 VSS.n2040 0.182778
R4772 VSS.n117 VSS 0.182492
R4773 VSS.n113 VSS.n112 0.180913
R4774 VSS.n1133 VSS.n1132 0.178908
R4775 VSS.n294 VSS.n291 0.177207
R4776 VSS.n297 VSS.n294 0.177207
R4777 VSS.n300 VSS.n297 0.177207
R4778 VSS.n303 VSS.n300 0.177207
R4779 VSS.n306 VSS.n303 0.177207
R4780 VSS.n309 VSS.n306 0.177207
R4781 VSS.n312 VSS.n309 0.177207
R4782 VSS.n395 VSS.n392 0.177207
R4783 VSS.n402 VSS.n399 0.177207
R4784 VSS.n409 VSS.n406 0.177207
R4785 VSS.n416 VSS.n413 0.177207
R4786 VSS.n2029 VSS.n2027 0.177207
R4787 VSS.n2023 VSS.n2019 0.177207
R4788 VSS.n2015 VSS.n2012 0.177207
R4789 VSS.n2008 VSS.n2005 0.177207
R4790 VSS.n208 VSS.n205 0.177207
R4791 VSS.n211 VSS.n208 0.177207
R4792 VSS.n214 VSS.n211 0.177207
R4793 VSS.n217 VSS.n214 0.177207
R4794 VSS.n220 VSS.n217 0.177207
R4795 VSS.n223 VSS.n220 0.177207
R4796 VSS.n225 VSS.n223 0.177207
R4797 VSS.n85 VSS.n25 0.167289
R4798 VSS.n1129 VSS.n1128 0.165962
R4799 VSS VSS.n22 0.165638
R4800 VSS.n1069 VSS.n1068 0.161394
R4801 VSS.n893 VSS.n892 0.160891
R4802 VSS.n1058 VSS.n1054 0.160039
R4803 VSS.n1067 VSS.n987 0.158377
R4804 VSS VSS.n2461 0.158206
R4805 VSS.n2277 VSS.n2274 0.156125
R4806 VSS.n1394 VSS.n1392 0.155256
R4807 VSS.n954 VSS.n951 0.155256
R4808 VSS.n14 VSS.n13 0.154904
R4809 VSS.n1172 VSS 0.154423
R4810 VSS.n2197 VSS.n2196 0.152211
R4811 VSS.n612 VSS.n609 0.1505
R4812 VSS.n609 VSS.n606 0.1505
R4813 VSS.n606 VSS.n603 0.1505
R4814 VSS.n603 VSS.n600 0.1505
R4815 VSS.n600 VSS.n597 0.1505
R4816 VSS.n919 VSS.n916 0.1505
R4817 VSS.n916 VSS.n913 0.1505
R4818 VSS.n913 VSS.n910 0.1505
R4819 VSS.n910 VSS.n907 0.1505
R4820 VSS.n168 VSS.n163 0.149643
R4821 VSS.n1995 VSS.n1994 0.149643
R4822 VSS.n1851 VSS.n1848 0.149643
R4823 VSS.n1559 VSS.n1556 0.149643
R4824 VSS.n1502 VSS.n1500 0.149643
R4825 VSS.n842 VSS.n689 0.149643
R4826 VSS.n822 VSS.n821 0.149643
R4827 VSS.n2071 VSS.n2069 0.149643
R4828 VSS.n1408 VSS.n1404 0.148671
R4829 VSS.n1404 VSS.n1402 0.148671
R4830 VSS.n1402 VSS.n1399 0.148671
R4831 VSS.n1399 VSS.n1396 0.148671
R4832 VSS.n1396 VSS.n1394 0.148671
R4833 VSS.n967 VSS.n966 0.148671
R4834 VSS.n966 VSS.n963 0.148671
R4835 VSS.n963 VSS.n960 0.148671
R4836 VSS.n960 VSS.n957 0.148671
R4837 VSS.n957 VSS.n954 0.148671
R4838 VSS.n1905 VSS.n1902 0.147071
R4839 VSS.n1029 VSS.n1026 0.147071
R4840 VSS.n1110 VSS.n1108 0.147071
R4841 VSS.n1705 VSS.n1703 0.147071
R4842 VSS.n100 VSS 0.145885
R4843 VSS VSS.n2269 0.144875
R4844 VSS.n1380 VSS.n1378 0.144731
R4845 VSS.n1384 VSS.n1380 0.144731
R4846 VSS.n1389 VSS.n1387 0.144731
R4847 VSS.n938 VSS.n935 0.144731
R4848 VSS.n940 VSS.n938 0.144731
R4849 VSS.n946 VSS.n944 0.144731
R4850 VSS.n2328 VSS.n2327 0.144447
R4851 VSS.n2169 VSS 0.143879
R4852 VSS VSS.n62 0.141929
R4853 VSS.n1424 VSS.n1423 0.139389
R4854 VSS.n1423 VSS.n1418 0.139389
R4855 VSS.n1418 VSS.n1416 0.139389
R4856 VSS.n1416 VSS.n1411 0.139389
R4857 VSS.n981 VSS.n980 0.139389
R4858 VSS.n980 VSS.n977 0.139389
R4859 VSS.n977 VSS.n974 0.139389
R4860 VSS.n974 VSS.n971 0.139389
R4861 VSS.n2193 VSS.n2191 0.138903
R4862 VSS.n2344 VSS.n2343 0.138304
R4863 VSS.n1424 VSS.n613 0.138278
R4864 VSS.n981 VSS.n923 0.138278
R4865 VSS.n1167 VSS.n1166 0.137808
R4866 VSS.n1458 VSS.n1457 0.137706
R4867 VSS.n2331 VSS.n2330 0.137236
R4868 VSS.n314 VSS.n312 0.137167
R4869 VSS.n228 VSS.n225 0.137167
R4870 VSS.n76 VSS 0.137136
R4871 VSS.n2314 VSS 0.137136
R4872 VSS VSS.n2254 0.137136
R4873 VSS VSS.n2233 0.137136
R4874 VSS.n895 VSS.n894 0.136757
R4875 VSS.n384 VSS.n383 0.136634
R4876 VSS.n1271 VSS.n1268 0.1355
R4877 VSS.n1274 VSS.n1271 0.1355
R4878 VSS.n1277 VSS.n1274 0.1355
R4879 VSS.n1280 VSS.n1277 0.1355
R4880 VSS.n1283 VSS.n1280 0.1355
R4881 VSS.n1286 VSS.n1283 0.1355
R4882 VSS.n1245 VSS.n1242 0.1355
R4883 VSS.n1242 VSS.n1239 0.1355
R4884 VSS.n1239 VSS.n1236 0.1355
R4885 VSS.n1236 VSS.n1233 0.1355
R4886 VSS.n1233 VSS.n1230 0.1355
R4887 VSS.n1230 VSS.n1226 0.1355
R4888 VSS.n1473 VSS.n1472 0.135039
R4889 VSS VSS.n1105 0.132962
R4890 VSS.n1752 VSS.n1747 0.132808
R4891 VSS.n19 VSS.n18 0.13261
R4892 VSS.n1333 VSS.n1330 0.132565
R4893 VSS.n1330 VSS.n1327 0.132565
R4894 VSS.n1327 VSS.n1324 0.132565
R4895 VSS.n1324 VSS.n1321 0.132565
R4896 VSS.n1321 VSS.n1316 0.132565
R4897 VSS.n1316 VSS.n1312 0.132565
R4898 VSS.n1184 VSS.n1180 0.132565
R4899 VSS.n1187 VSS.n1184 0.132565
R4900 VSS.n1190 VSS.n1187 0.132565
R4901 VSS.n1194 VSS.n1190 0.132565
R4902 VSS.n1197 VSS.n1194 0.132565
R4903 VSS.n1200 VSS.n1197 0.132565
R4904 VSS.n1612 VSS.n1611 0.132449
R4905 VSS.n2058 VSS.n2055 0.132286
R4906 VSS.n2055 VSS.n2053 0.132286
R4907 VSS.n145 VSS.n143 0.132286
R4908 VSS.n159 VSS.n145 0.132286
R4909 VSS.n171 VSS.n168 0.132286
R4910 VSS.n174 VSS.n171 0.132286
R4911 VSS.n177 VSS.n174 0.132286
R4912 VSS.n184 VSS.n177 0.132286
R4913 VSS.n187 VSS.n184 0.132286
R4914 VSS.n190 VSS.n187 0.132286
R4915 VSS.n193 VSS.n190 0.132286
R4916 VSS.n196 VSS.n193 0.132286
R4917 VSS.n200 VSS.n196 0.132286
R4918 VSS.n2144 VSS.n200 0.132286
R4919 VSS.n2144 VSS.n2143 0.132286
R4920 VSS.n2143 VSS.n2140 0.132286
R4921 VSS.n2140 VSS.n2137 0.132286
R4922 VSS.n2137 VSS.n2133 0.132286
R4923 VSS.n2133 VSS.n2130 0.132286
R4924 VSS.n287 VSS.n284 0.132286
R4925 VSS.n284 VSS.n282 0.132286
R4926 VSS.n2001 VSS.n1999 0.132286
R4927 VSS.n1994 VSS.n1992 0.132286
R4928 VSS.n1992 VSS.n1989 0.132286
R4929 VSS.n1989 VSS.n1987 0.132286
R4930 VSS.n1987 VSS.n1985 0.132286
R4931 VSS.n1985 VSS.n1983 0.132286
R4932 VSS.n1983 VSS.n1981 0.132286
R4933 VSS.n1981 VSS.n1979 0.132286
R4934 VSS.n1979 VSS.n1976 0.132286
R4935 VSS.n1976 VSS.n1974 0.132286
R4936 VSS.n1974 VSS.n273 0.132286
R4937 VSS.n273 VSS.n271 0.132286
R4938 VSS.n271 VSS.n269 0.132286
R4939 VSS.n269 VSS.n266 0.132286
R4940 VSS.n266 VSS.n263 0.132286
R4941 VSS.n263 VSS.n261 0.132286
R4942 VSS.n1911 VSS.n1908 0.132286
R4943 VSS.n1914 VSS.n1911 0.132286
R4944 VSS.n1917 VSS.n1914 0.132286
R4945 VSS.n1920 VSS.n1917 0.132286
R4946 VSS.n1923 VSS.n1920 0.132286
R4947 VSS.n1926 VSS.n1923 0.132286
R4948 VSS.n1929 VSS.n1926 0.132286
R4949 VSS.n1947 VSS.n1944 0.132286
R4950 VSS.n1944 VSS.n1941 0.132286
R4951 VSS.n253 VSS.n250 0.132286
R4952 VSS.n256 VSS.n253 0.132286
R4953 VSS.n1853 VSS.n1851 0.132286
R4954 VSS.n1856 VSS.n1853 0.132286
R4955 VSS.n1859 VSS.n1856 0.132286
R4956 VSS.n1862 VSS.n1859 0.132286
R4957 VSS.n1865 VSS.n1862 0.132286
R4958 VSS.n1868 VSS.n1865 0.132286
R4959 VSS.n1870 VSS.n1868 0.132286
R4960 VSS.n1873 VSS.n1870 0.132286
R4961 VSS.n1970 VSS.n1873 0.132286
R4962 VSS.n1970 VSS.n1969 0.132286
R4963 VSS.n1969 VSS.n1966 0.132286
R4964 VSS.n1966 VSS.n1963 0.132286
R4965 VSS.n1963 VSS.n1961 0.132286
R4966 VSS.n1961 VSS.n1959 0.132286
R4967 VSS.n1959 VSS.n1956 0.132286
R4968 VSS.n446 VSS.n443 0.132286
R4969 VSS.n1834 VSS.n1831 0.132286
R4970 VSS.n1837 VSS.n1834 0.132286
R4971 VSS.n1840 VSS.n1837 0.132286
R4972 VSS.n1843 VSS.n1840 0.132286
R4973 VSS.n1846 VSS.n1843 0.132286
R4974 VSS.n439 VSS.n435 0.132286
R4975 VSS.n435 VSS.n432 0.132286
R4976 VSS.n432 VSS.n429 0.132286
R4977 VSS.n429 VSS.n426 0.132286
R4978 VSS.n426 VSS.n423 0.132286
R4979 VSS.n1878 VSS.n1875 0.132286
R4980 VSS.n1881 VSS.n1878 0.132286
R4981 VSS.n1884 VSS.n1881 0.132286
R4982 VSS.n1887 VSS.n1884 0.132286
R4983 VSS.n1890 VSS.n1887 0.132286
R4984 VSS.n1893 VSS.n1890 0.132286
R4985 VSS.n1896 VSS.n1893 0.132286
R4986 VSS.n1899 VSS.n1896 0.132286
R4987 VSS.n1902 VSS.n1899 0.132286
R4988 VSS.n1549 VSS.n1547 0.132286
R4989 VSS.n1551 VSS.n1549 0.132286
R4990 VSS.n1553 VSS.n1551 0.132286
R4991 VSS.n1562 VSS.n1559 0.132286
R4992 VSS.n1565 VSS.n1562 0.132286
R4993 VSS.n1568 VSS.n1565 0.132286
R4994 VSS.n1571 VSS.n1568 0.132286
R4995 VSS.n1574 VSS.n1571 0.132286
R4996 VSS.n1577 VSS.n1574 0.132286
R4997 VSS.n1580 VSS.n1577 0.132286
R4998 VSS.n1583 VSS.n1580 0.132286
R4999 VSS.n1586 VSS.n1583 0.132286
R5000 VSS.n1589 VSS.n1586 0.132286
R5001 VSS.n1592 VSS.n1589 0.132286
R5002 VSS.n1595 VSS.n1592 0.132286
R5003 VSS.n1598 VSS.n1595 0.132286
R5004 VSS.n1601 VSS.n1598 0.132286
R5005 VSS.n1604 VSS.n1601 0.132286
R5006 VSS.n871 VSS.n867 0.132286
R5007 VSS.n873 VSS.n871 0.132286
R5008 VSS.n876 VSS.n873 0.132286
R5009 VSS.n878 VSS.n876 0.132286
R5010 VSS.n864 VSS.n616 0.132286
R5011 VSS.n1373 VSS.n1370 0.132286
R5012 VSS.n1370 VSS.n1367 0.132286
R5013 VSS.n1367 VSS.n1364 0.132286
R5014 VSS.n1364 VSS.n1361 0.132286
R5015 VSS.n1024 VSS.n1022 0.132286
R5016 VSS.n1019 VSS.n1017 0.132286
R5017 VSS.n1017 VSS.n1015 0.132286
R5018 VSS.n1015 VSS.n1013 0.132286
R5019 VSS.n1013 VSS.n1011 0.132286
R5020 VSS.n1540 VSS.n1538 0.132286
R5021 VSS.n1542 VSS.n1540 0.132286
R5022 VSS.n1610 VSS.n1608 0.132286
R5023 VSS.n1504 VSS.n1502 0.132286
R5024 VSS.n1506 VSS.n1504 0.132286
R5025 VSS.n1508 VSS.n1506 0.132286
R5026 VSS.n1510 VSS.n1508 0.132286
R5027 VSS.n1512 VSS.n1510 0.132286
R5028 VSS.n1514 VSS.n1512 0.132286
R5029 VSS.n1516 VSS.n1514 0.132286
R5030 VSS.n1518 VSS.n1516 0.132286
R5031 VSS.n1520 VSS.n1518 0.132286
R5032 VSS.n1522 VSS.n1520 0.132286
R5033 VSS.n1524 VSS.n1522 0.132286
R5034 VSS.n1526 VSS.n1524 0.132286
R5035 VSS.n1528 VSS.n1526 0.132286
R5036 VSS.n1530 VSS.n1528 0.132286
R5037 VSS.n1532 VSS.n1530 0.132286
R5038 VSS.n1487 VSS.n1485 0.132286
R5039 VSS.n1489 VSS.n1487 0.132286
R5040 VSS.n1491 VSS.n1489 0.132286
R5041 VSS.n1493 VSS.n1491 0.132286
R5042 VSS.n1495 VSS.n1493 0.132286
R5043 VSS.n1497 VSS.n1495 0.132286
R5044 VSS.n1499 VSS.n1497 0.132286
R5045 VSS.n993 VSS.n990 0.132286
R5046 VSS.n996 VSS.n993 0.132286
R5047 VSS.n999 VSS.n996 0.132286
R5048 VSS.n1002 VSS.n999 0.132286
R5049 VSS.n1005 VSS.n1002 0.132286
R5050 VSS.n1008 VSS.n1005 0.132286
R5051 VSS.n1048 VSS.n1008 0.132286
R5052 VSS.n1048 VSS.n1047 0.132286
R5053 VSS.n1047 VSS.n1045 0.132286
R5054 VSS.n1045 VSS.n1042 0.132286
R5055 VSS.n1042 VSS.n1040 0.132286
R5056 VSS.n1040 VSS.n1037 0.132286
R5057 VSS.n1037 VSS.n1035 0.132286
R5058 VSS.n1035 VSS.n1031 0.132286
R5059 VSS.n1031 VSS.n1029 0.132286
R5060 VSS.n1164 VSS.n1160 0.132286
R5061 VSS.n1160 VSS.n1157 0.132286
R5062 VSS.n1157 VSS.n881 0.132286
R5063 VSS.n1124 VSS.n881 0.132286
R5064 VSS.n1124 VSS.n1123 0.132286
R5065 VSS.n1123 VSS.n1115 0.132286
R5066 VSS.n1115 VSS.n1113 0.132286
R5067 VSS.n1113 VSS.n1110 0.132286
R5068 VSS.n625 VSS.n622 0.132286
R5069 VSS.n628 VSS.n625 0.132286
R5070 VSS.n631 VSS.n628 0.132286
R5071 VSS.n634 VSS.n631 0.132286
R5072 VSS.n637 VSS.n634 0.132286
R5073 VSS.n640 VSS.n637 0.132286
R5074 VSS.n643 VSS.n640 0.132286
R5075 VSS.n652 VSS.n649 0.132286
R5076 VSS.n649 VSS.n646 0.132286
R5077 VSS.n766 VSS.n763 0.132286
R5078 VSS.n769 VSS.n766 0.132286
R5079 VSS.n689 VSS.n687 0.132286
R5080 VSS.n687 VSS.n685 0.132286
R5081 VSS.n685 VSS.n683 0.132286
R5082 VSS.n683 VSS.n681 0.132286
R5083 VSS.n681 VSS.n679 0.132286
R5084 VSS.n679 VSS.n677 0.132286
R5085 VSS.n677 VSS.n675 0.132286
R5086 VSS.n675 VSS.n673 0.132286
R5087 VSS.n673 VSS.n671 0.132286
R5088 VSS.n671 VSS.n669 0.132286
R5089 VSS.n669 VSS.n667 0.132286
R5090 VSS.n667 VSS.n665 0.132286
R5091 VSS.n665 VSS.n663 0.132286
R5092 VSS.n663 VSS.n661 0.132286
R5093 VSS.n661 VSS.n659 0.132286
R5094 VSS.n841 VSS.n838 0.132286
R5095 VSS.n838 VSS.n835 0.132286
R5096 VSS.n835 VSS.n832 0.132286
R5097 VSS.n828 VSS.n825 0.132286
R5098 VSS.n821 VSS.n818 0.132286
R5099 VSS.n818 VSS.n815 0.132286
R5100 VSS.n815 VSS.n812 0.132286
R5101 VSS.n812 VSS.n809 0.132286
R5102 VSS.n809 VSS.n806 0.132286
R5103 VSS.n806 VSS.n803 0.132286
R5104 VSS.n803 VSS.n800 0.132286
R5105 VSS.n800 VSS.n797 0.132286
R5106 VSS.n797 VSS.n794 0.132286
R5107 VSS.n794 VSS.n791 0.132286
R5108 VSS.n791 VSS.n788 0.132286
R5109 VSS.n788 VSS.n785 0.132286
R5110 VSS.n785 VSS.n782 0.132286
R5111 VSS.n782 VSS.n779 0.132286
R5112 VSS.n779 VSS.n776 0.132286
R5113 VSS.n1651 VSS.n1648 0.132286
R5114 VSS.n1648 VSS.n1645 0.132286
R5115 VSS.n1645 VSS.n1642 0.132286
R5116 VSS.n1642 VSS.n1639 0.132286
R5117 VSS.n2064 VSS.n2061 0.132286
R5118 VSS.n2066 VSS.n2064 0.132286
R5119 VSS.n1662 VSS.n1659 0.132286
R5120 VSS.n1665 VSS.n1662 0.132286
R5121 VSS.n1668 VSS.n1665 0.132286
R5122 VSS.n1671 VSS.n1668 0.132286
R5123 VSS.n1674 VSS.n1671 0.132286
R5124 VSS.n1676 VSS.n1674 0.132286
R5125 VSS.n1679 VSS.n1676 0.132286
R5126 VSS.n1682 VSS.n1679 0.132286
R5127 VSS.n1685 VSS.n1682 0.132286
R5128 VSS.n1688 VSS.n1685 0.132286
R5129 VSS.n1691 VSS.n1688 0.132286
R5130 VSS.n1694 VSS.n1691 0.132286
R5131 VSS.n1697 VSS.n1694 0.132286
R5132 VSS.n1700 VSS.n1697 0.132286
R5133 VSS.n1703 VSS.n1700 0.132286
R5134 VSS.n1729 VSS.n1726 0.132286
R5135 VSS.n1746 VSS.n1743 0.132286
R5136 VSS.n1743 VSS.n1740 0.132286
R5137 VSS.n1740 VSS.n1737 0.132286
R5138 VSS.n1737 VSS.n1734 0.132286
R5139 VSS.n1734 VSS.n1732 0.132286
R5140 VSS.n2110 VSS.n2107 0.132286
R5141 VSS.n2112 VSS.n2110 0.132286
R5142 VSS.n2123 VSS.n2121 0.132286
R5143 VSS.n2073 VSS.n2071 0.132286
R5144 VSS.n2075 VSS.n2073 0.132286
R5145 VSS.n2077 VSS.n2075 0.132286
R5146 VSS.n2079 VSS.n2077 0.132286
R5147 VSS.n2081 VSS.n2079 0.132286
R5148 VSS.n2083 VSS.n2081 0.132286
R5149 VSS.n2085 VSS.n2083 0.132286
R5150 VSS.n2087 VSS.n2085 0.132286
R5151 VSS.n2089 VSS.n2087 0.132286
R5152 VSS.n2091 VSS.n2089 0.132286
R5153 VSS.n2093 VSS.n2091 0.132286
R5154 VSS.n2095 VSS.n2093 0.132286
R5155 VSS.n2097 VSS.n2095 0.132286
R5156 VSS.n2099 VSS.n2097 0.132286
R5157 VSS.n2101 VSS.n2099 0.132286
R5158 VSS.n1171 VSS.n1170 0.1305
R5159 VSS.n1334 VSS.n1333 0.128652
R5160 VSS.n1356 VSS.n1180 0.128652
R5161 VSS.n2280 VSS 0.127807
R5162 VSS.n515 VSS.n512 0.127656
R5163 VSS.n744 VSS.n743 0.127656
R5164 VSS.n1790 VSS.n1786 0.127423
R5165 VSS VSS.n21 0.127258
R5166 VSS.n440 VSS.n439 0.125857
R5167 VSS.n867 VSS.n865 0.125857
R5168 VSS.n1659 VSS.n1656 0.125857
R5169 VSS.n1453 VSS 0.125794
R5170 VSS.n365 VSS.n364 0.12579
R5171 VSS.n1292 VSS.n1289 0.1255
R5172 VSS.n1299 VSS.n1296 0.1255
R5173 VSS.n1224 VSS.n1221 0.1255
R5174 VSS.n1217 VSS.n1214 0.1255
R5175 VSS.n259 VSS.n256 0.124571
R5176 VSS.n772 VSS.n769 0.124571
R5177 VSS.n1264 VSS.n1262 0.124126
R5178 VSS.n1262 VSS.n1258 0.124126
R5179 VSS.n1258 VSS.n1256 0.124126
R5180 VSS.n1256 VSS.n1253 0.124126
R5181 VSS.n1253 VSS.n1250 0.124126
R5182 VSS.n1342 VSS.n1338 0.124126
R5183 VSS.n1345 VSS.n1342 0.124126
R5184 VSS.n1347 VSS.n1345 0.124126
R5185 VSS.n1351 VSS.n1347 0.124126
R5186 VSS.n1355 VSS.n1351 0.124126
R5187 VSS.n1545 VSS.n1543 0.123929
R5188 VSS.n763 VSS.n760 0.123929
R5189 VSS.n2117 VSS.n2113 0.123929
R5190 VSS.n2341 VSS.n2340 0.123883
R5191 VSS.n1956 VSS.n1952 0.123286
R5192 VSS.n1535 VSS.n1532 0.123286
R5193 VSS.n659 VSS.n657 0.123286
R5194 VSS.n2104 VSS.n2101 0.123286
R5195 VSS.n2130 VSS.n2127 0.122
R5196 VSS.n1606 VSS.n1604 0.122
R5197 VSS.n1450 VSS.n1449 0.121824
R5198 VSS.n1615 VSS.n1612 0.12105
R5199 VSS.n456 VSS.n453 0.12105
R5200 VSS.n510 VSS.n508 0.120158
R5201 VSS.n747 VSS.n745 0.120158
R5202 VSS.n1758 VSS.n1752 0.119731
R5203 VSS.n1793 VSS.n1790 0.119731
R5204 VSS.n1828 VSS.n1827 0.118962
R5205 VSS VSS.n1083 0.118573
R5206 VSS.n1086 VSS 0.118573
R5207 VSS.n2302 VSS.n2301 0.118573
R5208 VSS.n2304 VSS.n2303 0.118573
R5209 VSS.n2308 VSS.n2307 0.118573
R5210 VSS.n2240 VSS.n2239 0.118573
R5211 VSS.n2242 VSS.n2241 0.118573
R5212 VSS.n2246 VSS.n2245 0.118573
R5213 VSS.n2219 VSS.n2218 0.118573
R5214 VSS.n2221 VSS.n2220 0.118573
R5215 VSS.n2225 VSS.n2224 0.118573
R5216 VSS.n2190 VSS.n2189 0.118573
R5217 VSS.n13 VSS.n12 0.118573
R5218 VSS.n88 VSS.n87 0.118573
R5219 VSS.n86 VSS.n85 0.118573
R5220 VSS.n2159 VSS.n2158 0.118573
R5221 VSS.n39 VSS.n38 0.118573
R5222 VSS.n2261 VSS.n2260 0.118573
R5223 VSS.n2259 VSS.n2179 0.118573
R5224 VSS.n69 VSS.n68 0.118573
R5225 VSS.n71 VSS.n70 0.118573
R5226 VSS.n73 VSS.n72 0.118573
R5227 VSS VSS.n1463 0.118373
R5228 VSS.n512 VSS.n507 0.117958
R5229 VSS.n744 VSS.n716 0.117958
R5230 VSS.n410 VSS.n409 0.117939
R5231 VSS.n2012 VSS.n2009 0.117939
R5232 VSS.n1385 VSS 0.117309
R5233 VSS.n941 VSS 0.117309
R5234 VSS.n829 VSS.n748 0.117084
R5235 VSS.n399 VSS.n396 0.116841
R5236 VSS.n2024 VSS.n2023 0.116841
R5237 VSS.n2350 VSS.n2349 0.116405
R5238 VSS VSS.n382 0.115458
R5239 VSS VSS.n2182 0.115271
R5240 VSS.n2249 VSS 0.115271
R5241 VSS.n2228 VSS 0.115271
R5242 VSS.n18 VSS 0.115271
R5243 VSS VSS.n78 0.115271
R5244 VSS.n29 VSS 0.115271
R5245 VSS.n2231 VSS 0.115271
R5246 VSS.n44 VSS 0.115271
R5247 VSS.n2252 VSS 0.115271
R5248 VSS VSS.n2317 0.115271
R5249 VSS VSS.n2315 0.115271
R5250 VSS.n75 VSS 0.115271
R5251 VSS.n613 VSS.n612 0.114944
R5252 VSS.n1445 VSS 0.114176
R5253 VSS VSS.n2192 0.113945
R5254 VSS.n923 VSS.n919 0.113833
R5255 VSS.n1385 VSS.n1384 0.112423
R5256 VSS.n941 VSS.n940 0.112423
R5257 VSS.n518 VSS.n515 0.111968
R5258 VSS.n521 VSS.n518 0.111968
R5259 VSS.n524 VSS.n521 0.111968
R5260 VSS.n527 VSS.n524 0.111968
R5261 VSS.n530 VSS.n527 0.111968
R5262 VSS.n534 VSS.n530 0.111968
R5263 VSS.n537 VSS.n534 0.111968
R5264 VSS.n539 VSS.n537 0.111968
R5265 VSS.n543 VSS.n539 0.111968
R5266 VSS.n1617 VSS.n1615 0.111968
R5267 VSS.n1620 VSS.n1617 0.111968
R5268 VSS.n1622 VSS.n1620 0.111968
R5269 VSS.n1625 VSS.n1622 0.111968
R5270 VSS.n1627 VSS.n1625 0.111968
R5271 VSS.n1630 VSS.n1627 0.111968
R5272 VSS.n1632 VSS.n1630 0.111968
R5273 VSS.n1635 VSS.n1632 0.111968
R5274 VSS.n1637 VSS.n1635 0.111968
R5275 VSS.n459 VSS.n456 0.111968
R5276 VSS.n462 VSS.n459 0.111968
R5277 VSS.n465 VSS.n462 0.111968
R5278 VSS.n468 VSS.n465 0.111968
R5279 VSS.n471 VSS.n468 0.111968
R5280 VSS.n474 VSS.n471 0.111968
R5281 VSS.n476 VSS.n474 0.111968
R5282 VSS.n479 VSS.n476 0.111968
R5283 VSS.n481 VSS.n479 0.111968
R5284 VSS.n743 VSS.n740 0.111968
R5285 VSS.n740 VSS.n737 0.111968
R5286 VSS.n737 VSS.n734 0.111968
R5287 VSS.n734 VSS.n731 0.111968
R5288 VSS.n731 VSS.n728 0.111968
R5289 VSS.n728 VSS.n725 0.111968
R5290 VSS.n725 VSS.n722 0.111968
R5291 VSS.n722 VSS.n719 0.111968
R5292 VSS.n719 VSS.n449 0.111968
R5293 VSS.n2353 VSS.n2352 0.111598
R5294 VSS.n2347 VSS 0.111331
R5295 VSS.n2334 VSS 0.111331
R5296 VSS.n1461 VSS 0.110913
R5297 VSS.n115 VSS 0.109909
R5298 VSS.n2158 VSS.n35 0.109491
R5299 VSS.n139 VSS.n138 0.109351
R5300 VSS.n968 VSS.n927 0.107167
R5301 VSS VSS.n33 0.106575
R5302 VSS.n1828 VSS.n446 0.105286
R5303 VSS.n1747 VSS.n1729 0.105286
R5304 VSS.n2356 VSS.n2355 0.104387
R5305 VSS.n2189 VSS.n9 0.102885
R5306 VSS.n1948 VSS.n1929 0.102071
R5307 VSS.n845 VSS.n842 0.102071
R5308 VSS.n1536 VSS.n556 0.102071
R5309 VSS.n1500 VSS.n1499 0.102071
R5310 VSS.n653 VSS.n643 0.102071
R5311 VSS.n2069 VSS.n2066 0.102071
R5312 VSS.n2314 VSS.n2182 0.10206
R5313 VSS.n2254 VSS.n2249 0.10206
R5314 VSS.n2233 VSS.n2228 0.10206
R5315 VSS.n76 VSS.n75 0.10206
R5316 VSS.n1336 VSS.n1335 0.101005
R5317 VSS.n1165 VSS.n1164 0.100786
R5318 VSS.n289 VSS.n288 0.1005
R5319 VSS.n1951 VSS.n1949 0.1005
R5320 VSS.n2068 VSS.n2067 0.1005
R5321 VSS.n2103 VSS.n2102 0.1005
R5322 VSS.n619 VSS.n617 0.1005
R5323 VSS.n656 VSS.n654 0.1005
R5324 VSS.n1480 VSS.n1479 0.1005
R5325 VSS.n1534 VSS.n1533 0.1005
R5326 VSS.n1392 VSS.n1389 0.0996745
R5327 VSS.n951 VSS.n946 0.0996745
R5328 VSS.n1066 VSS.n1065 0.0983462
R5329 VSS.n1312 VSS.n1310 0.0983261
R5330 VSS.n1204 VSS.n1200 0.0983261
R5331 VSS.n1071 VSS.n1070 0.0976538
R5332 VSS.n1765 VSS.n1762 0.0966538
R5333 VSS.n1768 VSS.n1765 0.0966538
R5334 VSS.n1775 VSS.n1772 0.0966538
R5335 VSS.n1778 VSS.n1775 0.0966538
R5336 VSS.n1785 VSS.n1782 0.0966538
R5337 VSS.n1801 VSS.n1797 0.0966538
R5338 VSS.n1804 VSS.n1801 0.0966538
R5339 VSS.n1815 VSS.n1808 0.0966538
R5340 VSS.n1818 VSS.n1815 0.0966538
R5341 VSS.n1826 VSS.n1823 0.0966538
R5342 VSS.n1908 VSS.n1905 0.0962857
R5343 VSS.n1026 VSS.n1024 0.0962857
R5344 VSS.n1726 VSS.n1705 0.0962857
R5345 VSS.n485 VSS.n483 0.095839
R5346 VSS.n489 VSS.n485 0.095839
R5347 VSS.n491 VSS.n489 0.095839
R5348 VSS.n495 VSS.n491 0.095839
R5349 VSS.n498 VSS.n495 0.095839
R5350 VSS.n501 VSS.n498 0.095839
R5351 VSS.n504 VSS.n501 0.095839
R5352 VSS.n507 VSS.n504 0.095839
R5353 VSS.n695 VSS.n692 0.095839
R5354 VSS.n698 VSS.n695 0.095839
R5355 VSS.n701 VSS.n698 0.095839
R5356 VSS.n704 VSS.n701 0.095839
R5357 VSS.n708 VSS.n704 0.095839
R5358 VSS.n710 VSS.n708 0.095839
R5359 VSS.n714 VSS.n710 0.095839
R5360 VSS.n716 VSS.n714 0.095839
R5361 VSS.n1022 VSS.n1020 0.0956429
R5362 VSS.n443 VSS.n440 0.095
R5363 VSS.n865 VSS.n864 0.095
R5364 VSS.n1374 VSS.n616 0.095
R5365 VSS.n1485 VSS.n1483 0.095
R5366 VSS.n1656 VSS.n1651 0.095
R5367 VSS.n1289 VSS.n1286 0.0945
R5368 VSS.n1226 VSS.n1224 0.0945
R5369 VSS.n2374 VSS 0.0924934
R5370 VSS.n94 VSS.n93 0.0905
R5371 VSS.n96 VSS.n95 0.0905
R5372 VSS.n101 VSS.n100 0.0905
R5373 VSS.n1104 VSS 0.0905
R5374 VSS.n2349 VSS 0.0905
R5375 VSS.n2265 VSS.n2264 0.089875
R5376 VSS.n2267 VSS.n2266 0.089875
R5377 VSS.n2269 VSS.n2268 0.089875
R5378 VSS.n1065 VSS.n1064 0.0895769
R5379 VSS.n1167 VSS 0.0895769
R5380 VSS.n116 VSS.n115 0.0895055
R5381 VSS.n403 VSS.n402 0.0894024
R5382 VSS.n2019 VSS.n2016 0.0894024
R5383 VSS.n2164 VSS.n2163 0.0892586
R5384 VSS.n2168 VSS.n2167 0.0892586
R5385 VSS.n2170 VSS.n2169 0.0892586
R5386 VSS.n1064 VSS.n1063 0.0886538
R5387 VSS.n406 VSS.n403 0.0883049
R5388 VSS.n2016 VSS.n2015 0.0883049
R5389 VSS.n1449 VSS.n1448 0.0881535
R5390 VSS.n55 VSS.n54 0.088051
R5391 VSS.n59 VSS.n58 0.088051
R5392 VSS.n62 VSS.n61 0.088051
R5393 VSS VSS.n98 0.0879825
R5394 VSS.n2382 VSS 0.0879825
R5395 VSS VSS.n1072 0.0874595
R5396 VSS.n1082 VSS 0.0874595
R5397 VSS VSS.n595 0.0874595
R5398 VSS VSS.n882 0.0874595
R5399 VSS VSS.n2281 0.087375
R5400 VSS.n118 VSS.n117 0.0869264
R5401 VSS.n2174 VSS 0.0867759
R5402 VSS.n1471 VSS 0.0861997
R5403 VSS.n1782 VSS.n1779 0.0858846
R5404 VSS.n1823 VSS.n1819 0.0858846
R5405 VSS VSS.n1145 0.0857318
R5406 VSS.n1088 VSS 0.0856259
R5407 VSS VSS.n63 0.085602
R5408 VSS.n135 VSS 0.085027
R5409 VSS.n137 VSS 0.085027
R5410 VSS.n2325 VSS.n47 0.0847202
R5411 VSS.n2328 VSS.n45 0.0847202
R5412 VSS.n2331 VSS.n40 0.0847202
R5413 VSS.n2335 VSS.n35 0.0847202
R5414 VSS.n2338 VSS.n32 0.0847202
R5415 VSS.n2341 VSS.n30 0.0847202
R5416 VSS.n2344 VSS.n25 0.0847202
R5417 VSS.n2349 VSS.n22 0.0847202
R5418 VSS.n2353 VSS.n19 0.0847202
R5419 VSS.n2356 VSS.n14 0.0847202
R5420 VSS.n2359 VSS.n9 0.0847202
R5421 VSS.n2320 VSS.n2319 0.0847202
R5422 VSS.n935 VSS.n931 0.084688
R5423 VSS.n1478 VSS.n1476 0.0834286
R5424 VSS.n1848 VSS.n1847 0.0827857
R5425 VSS.n1171 VSS 0.0826538
R5426 VSS.n1608 VSS.n1606 0.0821429
R5427 VSS.n1411 VSS.n1409 0.0816111
R5428 VSS.n971 VSS.n968 0.0816111
R5429 VSS.n1306 VSS.n1303 0.0815
R5430 VSS.n1208 VSS.n1207 0.0815
R5431 VSS.n2232 VSS.n32 0.0814174
R5432 VSS.n1334 VSS.n1250 0.0806099
R5433 VSS.n1356 VSS.n1355 0.0806099
R5434 VSS.n1310 VSS.n1306 0.0805
R5435 VSS.n1207 VSS.n1204 0.0805
R5436 VSS.n163 VSS.n159 0.0795714
R5437 VSS.n2002 VSS.n2001 0.0795714
R5438 VSS.n1999 VSS.n1995 0.0795714
R5439 VSS.n261 VSS.n259 0.0795714
R5440 VSS.n1556 VSS.n1553 0.0795714
R5441 VSS.n825 VSS.n822 0.0795714
R5442 VSS.n776 VSS.n772 0.0795714
R5443 VSS.n2121 VSS.n2118 0.0795714
R5444 VSS.n2124 VSS.n2123 0.0795714
R5445 VSS.n98 VSS.n33 0.0779126
R5446 VSS.n364 VSS.n363 0.0777727
R5447 VSS.n2281 VSS.n2280 0.077375
R5448 VSS.n2359 VSS 0.0768798
R5449 VSS.n2175 VSS.n2174 0.0768448
R5450 VSS.n1309 VSS.n1307 0.076587
R5451 VSS.n1203 VSS.n1201 0.076587
R5452 VSS.n1055 VSS 0.0765345
R5453 VSS.n2324 VSS 0.0760786
R5454 VSS.n124 VSS.n113 0.0760505
R5455 VSS.n63 VSS.n21 0.0758061
R5456 VSS.n829 VSS.n828 0.0757143
R5457 VSS.n1611 VSS.n1610 0.0750714
R5458 VSS.n1469 VSS.n1468 0.0742201
R5459 VSS.n2263 VSS.n2175 0.0727596
R5460 VSS.n2069 VSS.n2058 0.0725
R5461 VSS.n1848 VSS.n287 0.0725
R5462 VSS.n1948 VSS.n1947 0.0725
R5463 VSS.n1500 VSS.n1478 0.0725
R5464 VSS.n1293 VSS.n1292 0.0725
R5465 VSS.n1221 VSS.n1218 0.0725
R5466 VSS.n1538 VSS.n1536 0.0725
R5467 VSS.n653 VSS.n652 0.0725
R5468 VSS.n842 VSS.n841 0.0725
R5469 VSS.n2107 VSS.n2105 0.0725
R5470 VSS.n375 VSS.n370 0.071566
R5471 VSS.n378 VSS.n377 0.0706762
R5472 VSS.n1358 VSS.n845 0.0692857
R5473 VSS.n122 VSS 0.0691188
R5474 VSS.n2373 VSS.n2372 0.0689718
R5475 VSS.n392 VSS.n344 0.0687711
R5476 VSS.n1009 VSS.n556 0.0686429
R5477 VSS.n386 VSS.n385 0.0675755
R5478 VSS.n350 VSS.n349 0.0675755
R5479 VSS.n367 VSS.n365 0.0675755
R5480 VSS.n133 VSS.n132 0.0675755
R5481 VSS.n2212 VSS.n2211 0.0675755
R5482 VSS.n2206 VSS.n2205 0.0675755
R5483 VSS.n2202 VSS.n2201 0.0675755
R5484 VSS.n111 VSS.n110 0.0675755
R5485 VSS.n360 VSS.n359 0.0675755
R5486 VSS.n2274 VSS 0.0666607
R5487 VSS.n417 VSS.n327 0.066576
R5488 VSS.n2003 VSS.n238 0.066576
R5489 VSS.n2043 VSS.n2042 0.066576
R5490 VSS.n1752 VSS.n1637 0.0657294
R5491 VSS.n1790 VSS.n481 0.0657294
R5492 VSS.n1302 VSS 0.0655
R5493 VSS VSS.n1211 0.0655
R5494 VSS.n1772 VSS.n1769 0.0651154
R5495 VSS.n1808 VSS.n1805 0.0651154
R5496 VSS.n1135 VSS.n1134 0.0644474
R5497 VSS.n1470 VSS.n1469 0.0643908
R5498 VSS.n1011 VSS.n1009 0.0641429
R5499 VSS.n1468 VSS.n1467 0.0640001
R5500 VSS.n1095 VSS.n1087 0.0636579
R5501 VSS.n2326 VSS.n2325 0.0635267
R5502 VSS.n1361 VSS.n1358 0.0635
R5503 VSS.n1061 VSS.n1060 0.0633448
R5504 VSS VSS.n123 0.0624266
R5505 VSS.n2351 VSS.n2350 0.0611231
R5506 VSS.n396 VSS.n395 0.0608659
R5507 VSS.n2027 VSS.n2024 0.0608659
R5508 VSS VSS.n1299 0.0605
R5509 VSS.n1214 VSS 0.0605
R5510 VSS.n413 VSS.n410 0.0597683
R5511 VSS.n2009 VSS.n2008 0.0597683
R5512 VSS.n1786 VSS.n543 0.0591239
R5513 VSS.n1827 VSS.n449 0.0591239
R5514 VSS.n1168 VSS.n1167 0.0591154
R5515 VSS.n1611 VSS.n1545 0.0577143
R5516 VSS.n832 VSS.n829 0.0570714
R5517 VSS.n1053 VSS 0.0565526
R5518 VSS VSS.n1055 0.0555862
R5519 VSS VSS.n1446 0.055266
R5520 VSS VSS.n1438 0.055266
R5521 VSS.n356 VSS 0.0548172
R5522 VSS.n2375 VSS.n2373 0.0543206
R5523 VSS.n1296 VSS.n1293 0.0535
R5524 VSS.n1218 VSS.n1217 0.0535
R5525 VSS.n1071 VSS 0.0533462
R5526 VSS.n2002 VSS.n240 0.0532143
R5527 VSS.n2118 VSS.n2117 0.0532143
R5528 VSS.n1448 VSS.n1447 0.0530664
R5529 VSS.n1759 VSS.n1758 0.0528077
R5530 VSS.n1794 VSS.n1793 0.0528077
R5531 VSS.n1268 VSS.n1265 0.0525
R5532 VSS.n1336 VSS.n1245 0.0525
R5533 VSS.n2357 VSS.n2356 0.051776
R5534 VSS.n2339 VSS.n2338 0.0507077
R5535 VSS VSS.n1445 0.05
R5536 VSS.n1145 VSS.n1144 0.0499702
R5537 VSS.n1089 VSS.n1088 0.0496447
R5538 VSS.n1464 VSS 0.0485224
R5539 VSS VSS.n2374 0.0459485
R5540 VSS.n379 VSS.n378 0.0449053
R5541 VSS.n1165 VSS.n878 0.0448571
R5542 VSS.n2354 VSS.n2353 0.0445653
R5543 VSS.n1303 VSS.n1302 0.0445
R5544 VSS.n1211 VSS.n1208 0.0445
R5545 VSS.n1762 VSS.n1759 0.0443462
R5546 VSS.n1797 VSS.n1794 0.0443462
R5547 VSS.n896 VSS.n895 0.044243
R5548 VSS.n130 VSS.n129 0.04
R5549 VSS.n2009 VSS 0.0396304
R5550 VSS.n410 VSS 0.0396304
R5551 VSS VSS.n1470 0.0395102
R5552 VSS.n2361 VSS.n2360 0.0386899
R5553 VSS.n2358 VSS.n2357 0.0386899
R5554 VSS.n2348 VSS.n2347 0.0386899
R5555 VSS.n2346 VSS.n2345 0.0386899
R5556 VSS.n2333 VSS.n2332 0.0386899
R5557 VSS.n2323 VSS.n2322 0.0386899
R5558 VSS.n1374 VSS.n1373 0.0377857
R5559 VSS.n2278 VSS 0.0377321
R5560 VSS VSS.n2354 0.0376217
R5561 VSS VSS.n2351 0.0376217
R5562 VSS VSS.n2342 0.0376217
R5563 VSS VSS.n2339 0.0376217
R5564 VSS VSS.n2329 0.0376217
R5565 VSS VSS.n2326 0.0376217
R5566 VSS.n1020 VSS.n1019 0.0371429
R5567 VSS VSS.n1455 0.0362353
R5568 VSS.n375 VSS.n354 0.036033
R5569 VSS.n2454 VSS.n2386 0.0357703
R5570 VSS.n1463 VSS.n1461 0.0356813
R5571 VSS.n2360 VSS.n2359 0.034951
R5572 VSS.n2320 VSS.n2178 0.0344169
R5573 VSS VSS.n1172 0.0335
R5574 VSS.n1105 VSS 0.0335
R5575 VSS.n1128 VSS 0.0335
R5576 VSS.n1387 VSS.n1385 0.0328077
R5577 VSS.n944 VSS.n941 0.0328077
R5578 VSS.n2342 VSS.n2341 0.0322804
R5579 VSS.n1769 VSS.n1768 0.0320385
R5580 VSS.n1805 VSS.n1804 0.0320385
R5581 VSS.n899 VSS.n898 0.0315345
R5582 VSS.n1141 VSS.n1140 0.0295909
R5583 VSS.n1168 VSS.n850 0.0286538
R5584 VSS.n1444 VSS.n1443 0.0283244
R5585 VSS.n2335 VSS.n2334 0.0277404
R5586 VSS.n1831 VSS.n1828 0.0275
R5587 VSS VSS.n1171 0.0275
R5588 VSS.n1747 VSS.n1746 0.0275
R5589 VSS.n2452 VSS.n2384 0.0267703
R5590 VSS.n381 VSS.n380 0.0263107
R5591 VSS.n1136 VSS.n1135 0.0257632
R5592 VSS.n894 VSS.n893 0.0251369
R5593 VSS.n2372 VSS.n2371 0.0241213
R5594 VSS.n1769 VSS 0.0239783
R5595 VSS.n1805 VSS 0.0239783
R5596 VSS VSS.n1454 0.0238824
R5597 VSS.n2379 VSS.n2378 0.0235097
R5598 VSS.n368 VSS.n357 0.0211167
R5599 VSS.n1460 VSS.n1459 0.0203529
R5600 VSS.n1456 VSS 0.0203529
R5601 VSS.n1451 VSS.n1450 0.0203529
R5602 VSS.n1847 VSS.n1846 0.0197857
R5603 VSS.n2332 VSS.n2331 0.0189273
R5604 VSS.n166 VSS.n165 0.0181879
R5605 VSS.n2345 VSS.n2344 0.017859
R5606 VSS.n987 VSS.n986 0.017595
R5607 VSS.n1457 VSS.n1456 0.0168235
R5608 VSS VSS.n47 0.0161881
R5609 VSS.n2322 VSS 0.0154555
R5610 VSS.n897 VSS.n896 0.0145782
R5611 VSS.n1139 VSS.n1138 0.0135995
R5612 VSS.n1139 VSS.n1136 0.0135929
R5613 VSS.n902 VSS.n901 0.0135726
R5614 VSS.n1472 VSS.n1471 0.013401
R5615 VSS.n2338 VSS.n2337 0.0130519
R5616 VSS.n2329 VSS.n2328 0.0117166
R5617 VSS.n2336 VSS.n2335 0.0114496
R5618 VSS.n1779 VSS.n1778 0.0112692
R5619 VSS.n1819 VSS.n1818 0.0112692
R5620 VSS.n1467 VSS 0.0112609
R5621 VSS.n1466 VSS.n1465 0.010087
R5622 VSS.n986 VSS 0.0100531
R5623 VSS.n380 VSS.n379 0.00961702
R5624 VSS.n1941 VSS.n1938 0.00885714
R5625 VSS.n1543 VSS.n1542 0.00885714
R5626 VSS.n2113 VSS.n2112 0.00885714
R5627 VSS.n2453 VSS.n2451 0.008809
R5628 VSS VSS.n1052 0.00839474
R5629 VSS.n901 VSS.n900 0.00834709
R5630 VSS.n1056 VSS 0.00825862
R5631 VSS.n2456 VSS.n2455 0.00798833
R5632 VSS.n1454 VSS.n1453 0.00711765
R5633 VSS.n357 VSS.n356 0.00644714
R5634 VSS.n2301 VSS 0.00545413
R5635 VSS.n2304 VSS 0.00545413
R5636 VSS.n2307 VSS 0.00545413
R5637 VSS.n2239 VSS 0.00545413
R5638 VSS.n2242 VSS 0.00545413
R5639 VSS.n2245 VSS 0.00545413
R5640 VSS.n2218 VSS 0.00545413
R5641 VSS.n2221 VSS 0.00545413
R5642 VSS.n2224 VSS 0.00545413
R5643 VSS VSS.n2190 0.00545413
R5644 VSS.n12 VSS 0.00545413
R5645 VSS.n88 VSS 0.00545413
R5646 VSS VSS.n86 0.00545413
R5647 VSS.n2159 VSS 0.00545413
R5648 VSS.n38 VSS 0.00545413
R5649 VSS.n2261 VSS 0.00545413
R5650 VSS VSS.n2259 0.00545413
R5651 VSS.n68 VSS 0.00545413
R5652 VSS.n70 VSS 0.00545413
R5653 VSS.n72 VSS 0.00545413
R5654 VSS VSS.n1460 0.00535294
R5655 VSS VSS.n1452 0.00535294
R5656 VSS.n902 VSS 0.00502514
R5657 VSS.n2321 VSS.n2320 0.004773
R5658 VSS.n900 VSS.n897 0.0046963
R5659 VSS.n2454 VSS.n2453 0.00463514
R5660 VSS.n1459 VSS.n1458 0.00447059
R5661 VSS.n1455 VSS 0.00447059
R5662 VSS.n1452 VSS.n1451 0.00447059
R5663 VSS.n1265 VSS.n1264 0.00445604
R5664 VSS.n1338 VSS.n1336 0.00445604
R5665 VSS.n93 VSS 0.00427622
R5666 VSS.n95 VSS 0.00427622
R5667 VSS.n101 VSS 0.00427622
R5668 VSS.n2264 VSS 0.00425
R5669 VSS.n2266 VSS 0.00425
R5670 VSS.n2268 VSS 0.00425
R5671 VSS.n2164 VSS 0.00422414
R5672 VSS.n2167 VSS 0.00422414
R5673 VSS.n2170 VSS 0.00422414
R5674 VSS.n55 VSS 0.00417347
R5675 VSS.n58 VSS 0.00417347
R5676 VSS.n61 VSS 0.00417347
R5677 VSS.n2325 VSS.n2324 0.00397181
R5678 VSS.n2309 VSS 0.00380275
R5679 VSS VSS.n2248 0.00380275
R5680 VSS VSS.n2227 0.00380275
R5681 VSS.n2210 VSS 0.00380275
R5682 VSS.n2208 VSS 0.00380275
R5683 VSS VSS.n2203 0.00380275
R5684 VSS VSS.n17 0.00380275
R5685 VSS.n79 VSS 0.00380275
R5686 VSS VSS.n28 0.00380275
R5687 VSS VSS.n2230 0.00380275
R5688 VSS VSS.n43 0.00380275
R5689 VSS VSS.n2251 0.00380275
R5690 VSS.n2318 VSS 0.00380275
R5691 VSS.n2316 VSS 0.00380275
R5692 VSS VSS.n74 0.00380275
R5693 VSS.n362 VSS 0.00380275
R5694 VSS VSS.n0 0.00380275
R5695 VSS.n1995 VSS.n247 0.00371429
R5696 VSS.n383 VSS 0.00352521
R5697 VSS.n2193 VSS 0.00352521
R5698 VSS VSS.n2273 0.0035
R5699 VSS.n2127 VSS.n2124 0.00307143
R5700 VSS.n99 VSS 0.00301748
R5701 VSS VSS.n2381 0.00301748
R5702 VSS.n1068 VSS.n1067 0.00301397
R5703 VSS.n2282 VSS 0.003
R5704 VSS.n119 VSS.n118 0.00298619
R5705 VSS VSS.n2173 0.00298276
R5706 VSS.n64 VSS 0.00294898
R5707 VSS VSS.n134 0.00293243
R5708 VSS VSS.n136 0.00293243
R5709 VSS.n1131 VSS 0.00286842
R5710 VSS.n417 VSS.n416 0.00269512
R5711 VSS.n1409 VSS.n1408 0.00269512
R5712 VSS.n2043 VSS.n2029 0.00269512
R5713 VSS.n2005 VSS.n2003 0.00269512
R5714 VSS.n2455 VSS.n2385 0.00268919
R5715 VSS.n2452 VSS.n2385 0.00244595
R5716 VSS VSS.n67 0.00219811
R5717 VSS.n52 VSS 0.00219811
R5718 VSS.n2155 VSS 0.00219811
R5719 VSS.n386 VSS 0.00219811
R5720 VSS.n349 VSS 0.00219811
R5721 VSS VSS.n367 0.00219811
R5722 VSS VSS.n2271 0.00219811
R5723 VSS.n132 VSS 0.00219811
R5724 VSS VSS.n2313 0.00219811
R5725 VSS.n2255 VSS 0.00219811
R5726 VSS.n2234 VSS 0.00219811
R5727 VSS.n2212 VSS 0.00219811
R5728 VSS.n2205 VSS 0.00219811
R5729 VSS.n2201 VSS 0.00219811
R5730 VSS.n2199 VSS 0.00219811
R5731 VSS.n2196 VSS 0.00219811
R5732 VSS.n110 VSS 0.00219811
R5733 VSS.n359 VSS 0.00219811
R5734 VSS.n124 VSS 0.00215138
R5735 VSS.n2361 VSS 0.00210237
R5736 VSS VSS.n2358 0.00210237
R5737 VSS VSS.n2348 0.00210237
R5738 VSS VSS.n2346 0.00210237
R5739 VSS VSS.n2336 0.00210237
R5740 VSS VSS.n2333 0.00210237
R5741 VSS VSS.n2323 0.00210237
R5742 VSS VSS.n2321 0.00210237
R5743 VSS.n512 VSS.n511 0.00202542
R5744 VSS.n748 VSS.n744 0.00202542
R5745 VSS.n1952 VSS.n1948 0.00178571
R5746 VSS.n1536 VSS.n1535 0.00178571
R5747 VSS.n657 VSS.n653 0.00178571
R5748 VSS.n2105 VSS.n2104 0.00178571
R5749 VSS.n138 VSS 0.00171622
R5750 VSS.n140 VSS 0.00171622
R5751 VSS.n2375 VSS 0.00169601
R5752 VSS.n1476 VSS.n1475 0.00168421
R5753 VSS.n927 VSS.n613 0.00161111
R5754 VSS.n923 VSS.n922 0.00161111
R5755 VSS.n968 VSS.n967 0.00159756
R5756 VSS VSS.n2277 0.00157143
R5757 VSS.n2355 VSS 0.00156825
R5758 VSS.n2352 VSS 0.00156825
R5759 VSS.n2343 VSS 0.00156825
R5760 VSS.n2340 VSS 0.00156825
R5761 VSS.n2330 VSS 0.00156825
R5762 VSS.n2327 VSS 0.00156825
R5763 VSS.n129 VSS 0.0015
R5764 VSS.n119 VSS 0.00149448
R5765 VSS VSS.n116 0.00149448
R5766 VSS.n1335 VSS.n1334 0.00147826
R5767 VSS.n1357 VSS.n1356 0.00147826
R5768 VSS VSS.n2263 0.00136539
R5769 VSS VSS.n381 0.0013
R5770 VSS.n376 VSS.n352 0.00129295
R5771 VSS VSS.n352 0.00129295
R5772 VSS VSS.n1097 0.00128947
R5773 VSS.n1097 VSS.n1095 0.00128947
R5774 VSS.n1134 VSS 0.00128947
R5775 VSS.n1052 VSS 0.00128947
R5776 VSS.n1056 VSS 0.00127586
R5777 VSS.n1060 VSS 0.00127586
R5778 VSS.n1786 VSS.n1785 0.00126923
R5779 VSS.n1827 VSS.n1826 0.00126923
R5780 VSS.n2371 VSS 0.00109801
R5781 VSS.n2378 VSS 0.00108252
R5782 VSS.n1166 VSS.n1165 0.000961538
R5783 VSS.n2450 VSS 0.000932432
R5784 VSS.n377 VSS.n376 0.000896476
R5785 VSS VSS.n1444 0.000843511
R5786 VSS.n850 VSS 0.000730769
R5787 VSS VSS.n1466 0.000695652
R5788 VSS.n2383 VSS 0.000613314
R5789 VCO_op.n9 VCO_op.t30 36.935
R5790 VCO_op.n3 VCO_op.t28 36.935
R5791 VCO_op.n23 VCO_op.t24 36.935
R5792 VCO_op.n17 VCO_op.t13 36.935
R5793 VCO_op.n41 VCO_op.t27 36.935
R5794 VCO_op.n35 VCO_op.t25 36.935
R5795 VCO_op.n65 VCO_op.t19 36.935
R5796 VCO_op.n59 VCO_op.t16 36.935
R5797 VCO_op.n52 VCO_op.t32 36.935
R5798 VCO_op.n28 VCO_op.t11 25.5364
R5799 VCO_op.n46 VCO_op.t12 25.5364
R5800 VCO_op.n70 VCO_op.t8 25.5361
R5801 VCO_op.n77 VCO_op.t26 25.5361
R5802 VCO_op.n9 VCO_op.t29 18.1962
R5803 VCO_op.n3 VCO_op.t23 18.1962
R5804 VCO_op.n23 VCO_op.t22 18.1962
R5805 VCO_op.n17 VCO_op.t10 18.1962
R5806 VCO_op.n41 VCO_op.t15 18.1962
R5807 VCO_op.n35 VCO_op.t20 18.1962
R5808 VCO_op.n65 VCO_op.t18 18.1962
R5809 VCO_op.n59 VCO_op.t14 18.1962
R5810 VCO_op.n52 VCO_op.t9 18.1962
R5811 VCO_op.n28 VCO_op.t21 14.0749
R5812 VCO_op.n46 VCO_op.t31 14.0749
R5813 VCO_op.n70 VCO_op.t17 14.0734
R5814 VCO_op.n77 VCO_op.t33 14.0734
R5815 VCO_op VCO_op.n92 13.2272
R5816 VCO_op.n75 VCO_op 5.77906
R5817 VCO_op.n79 VCO_op.n76 5.11659
R5818 VCO_op.n5 VCO_op.n2 4.5005
R5819 VCO_op.n5 VCO_op.n4 4.5005
R5820 VCO_op.n8 VCO_op.n7 4.5005
R5821 VCO_op.n10 VCO_op.n7 4.5005
R5822 VCO_op.n19 VCO_op.n16 4.5005
R5823 VCO_op.n19 VCO_op.n18 4.5005
R5824 VCO_op.n22 VCO_op.n21 4.5005
R5825 VCO_op.n24 VCO_op.n21 4.5005
R5826 VCO_op.n31 VCO_op.n30 4.5005
R5827 VCO_op.n30 VCO_op.n29 4.5005
R5828 VCO_op.n37 VCO_op.n34 4.5005
R5829 VCO_op.n37 VCO_op.n36 4.5005
R5830 VCO_op.n40 VCO_op.n39 4.5005
R5831 VCO_op.n42 VCO_op.n39 4.5005
R5832 VCO_op.n49 VCO_op.n48 4.5005
R5833 VCO_op.n48 VCO_op.n47 4.5005
R5834 VCO_op.n61 VCO_op.n58 4.5005
R5835 VCO_op.n61 VCO_op.n60 4.5005
R5836 VCO_op.n64 VCO_op.n63 4.5005
R5837 VCO_op.n66 VCO_op.n63 4.5005
R5838 VCO_op.n73 VCO_op.n72 4.5005
R5839 VCO_op.n72 VCO_op.n71 4.5005
R5840 VCO_op.n53 VCO_op.n50 4.5005
R5841 VCO_op.n80 VCO_op.n79 4.5005
R5842 VCO_op.n79 VCO_op.n78 4.5005
R5843 VCO_op.n76 VCO_op 4.43149
R5844 VCO_op.n81 VCO_op 4.16645
R5845 VCO_op.n74 VCO_op.n55 4.05348
R5846 VCO_op.n91 VCO_op.n85 3.58485
R5847 VCO_op.n90 VCO_op.n89 3.58485
R5848 VCO_op.n75 VCO_op.n74 3.5258
R5849 VCO_op.n91 VCO_op.n83 3.32833
R5850 VCO_op.n90 VCO_op.n87 3.32833
R5851 VCO_op.n74 VCO_op 2.3355
R5852 VCO_op VCO_op.n81 2.26961
R5853 VCO_op.n12 VCO_op.n11 2.25107
R5854 VCO_op.n26 VCO_op.n25 2.25107
R5855 VCO_op.n44 VCO_op.n43 2.25107
R5856 VCO_op.n68 VCO_op.n67 2.25107
R5857 VCO_op.n51 VCO_op.n50 2.24763
R5858 VCO_op.n55 VCO_op.n54 2.2455
R5859 VCO_op.n27 VCO_op.n14 2.24235
R5860 VCO_op.n45 VCO_op.n32 2.24235
R5861 VCO_op.n69 VCO_op.n56 2.24235
R5862 VCO_op.n13 VCO_op.n0 2.24235
R5863 VCO_op.n53 VCO_op.n52 2.12226
R5864 VCO_op.n4 VCO_op.n3 2.12175
R5865 VCO_op.n18 VCO_op.n17 2.12175
R5866 VCO_op.n36 VCO_op.n35 2.12175
R5867 VCO_op.n60 VCO_op.n59 2.12175
R5868 VCO_op.n10 VCO_op.n9 2.12075
R5869 VCO_op.n24 VCO_op.n23 2.12075
R5870 VCO_op.n42 VCO_op.n41 2.12075
R5871 VCO_op.n66 VCO_op.n65 2.12075
R5872 VCO_op.n7 VCO_op.n6 1.74297
R5873 VCO_op.n21 VCO_op.n20 1.74297
R5874 VCO_op.n39 VCO_op.n38 1.74297
R5875 VCO_op.n63 VCO_op.n62 1.74297
R5876 VCO_op.n76 VCO_op.n75 1.62556
R5877 VCO_op.n6 VCO_op.n1 1.49778
R5878 VCO_op.n20 VCO_op.n15 1.49778
R5879 VCO_op.n38 VCO_op.n33 1.49778
R5880 VCO_op.n62 VCO_op.n57 1.49778
R5881 VCO_op.n71 VCO_op.n70 1.42775
R5882 VCO_op.n78 VCO_op.n77 1.42775
R5883 VCO_op.n29 VCO_op.n28 1.42706
R5884 VCO_op.n47 VCO_op.n46 1.42706
R5885 VCO_op.n85 VCO_op.t0 1.1705
R5886 VCO_op.n85 VCO_op.n84 1.1705
R5887 VCO_op.n89 VCO_op.t3 1.1705
R5888 VCO_op.n89 VCO_op.n88 1.1705
R5889 VCO_op.n13 VCO_op.n12 0.97145
R5890 VCO_op.n27 VCO_op.n26 0.97145
R5891 VCO_op.n45 VCO_op.n44 0.97145
R5892 VCO_op.n69 VCO_op.n68 0.97145
R5893 VCO_op.n91 VCO_op.n90 0.68137
R5894 VCO_op.n83 VCO_op.t7 0.6505
R5895 VCO_op.n83 VCO_op.n82 0.6505
R5896 VCO_op.n87 VCO_op.t6 0.6505
R5897 VCO_op.n87 VCO_op.n86 0.6505
R5898 VCO_op VCO_op.n91 0.297891
R5899 VCO_op VCO_op.n31 0.1605
R5900 VCO_op VCO_op.n49 0.1605
R5901 VCO_op VCO_op.n73 0.1605
R5902 VCO_op VCO_op.n80 0.1605
R5903 VCO_op.n92 VCO_op 0.13958
R5904 VCO_op.n51 VCO_op 0.052998
R5905 VCO_op.n8 VCO_op 0.0473512
R5906 VCO_op.n2 VCO_op 0.0473512
R5907 VCO_op.n22 VCO_op 0.0473512
R5908 VCO_op.n16 VCO_op 0.0473512
R5909 VCO_op.n40 VCO_op 0.0473512
R5910 VCO_op.n34 VCO_op 0.0473512
R5911 VCO_op.n64 VCO_op 0.0473512
R5912 VCO_op.n58 VCO_op 0.0473512
R5913 VCO_op.n11 VCO_op.n8 0.0361897
R5914 VCO_op.n2 VCO_op.n1 0.0361897
R5915 VCO_op.n25 VCO_op.n22 0.0361897
R5916 VCO_op.n16 VCO_op.n15 0.0361897
R5917 VCO_op.n43 VCO_op.n40 0.0361897
R5918 VCO_op.n34 VCO_op.n33 0.0361897
R5919 VCO_op.n67 VCO_op.n64 0.0361897
R5920 VCO_op.n58 VCO_op.n57 0.0361897
R5921 VCO_op.n31 VCO_op.n14 0.03175
R5922 VCO_op.n49 VCO_op.n32 0.03175
R5923 VCO_op.n73 VCO_op.n56 0.03175
R5924 VCO_op.n80 VCO_op.n0 0.03175
R5925 VCO_op.n30 VCO_op.n27 0.0246174
R5926 VCO_op.n48 VCO_op.n45 0.0246174
R5927 VCO_op.n72 VCO_op.n69 0.0246174
R5928 VCO_op.n79 VCO_op.n13 0.0246174
R5929 VCO_op.n54 VCO_op.n53 0.0210263
R5930 VCO_op.n54 VCO_op.n51 0.0183424
R5931 VCO_op.n92 VCO_op 0.0161522
R5932 VCO_op.n6 VCO_op.n5 0.0131772
R5933 VCO_op.n20 VCO_op.n19 0.0131772
R5934 VCO_op.n38 VCO_op.n37 0.0131772
R5935 VCO_op.n62 VCO_op.n61 0.0131772
R5936 VCO_op.n55 VCO_op.n50 0.0128848
R5937 VCO_op.n12 VCO_op.n7 0.0122182
R5938 VCO_op.n26 VCO_op.n21 0.0122182
R5939 VCO_op.n44 VCO_op.n39 0.0122182
R5940 VCO_op.n68 VCO_op.n63 0.0122182
R5941 VCO_op.n81 VCO_op 0.00567241
R5942 VCO_op.n11 VCO_op.n10 0.00515517
R5943 VCO_op.n4 VCO_op.n1 0.00515517
R5944 VCO_op.n25 VCO_op.n24 0.00515517
R5945 VCO_op.n18 VCO_op.n15 0.00515517
R5946 VCO_op.n43 VCO_op.n42 0.00515517
R5947 VCO_op.n36 VCO_op.n33 0.00515517
R5948 VCO_op.n67 VCO_op.n66 0.00515517
R5949 VCO_op.n60 VCO_op.n57 0.00515517
R5950 VCO_op.n29 VCO_op.n14 0.00175
R5951 VCO_op.n47 VCO_op.n32 0.00175
R5952 VCO_op.n71 VCO_op.n56 0.00175
R5953 VCO_op.n78 VCO_op.n0 0.00175
R5954 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 37.1981
R5955 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 31.528
R5956 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 30.5752
R5957 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 24.6493
R5958 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 17.6611
R5959 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 17.0533
R5960 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 15.3826
R5961 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 7.62758
R5962 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 3.28711
R5963 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 2.99416
R5964 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.81128
R5965 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.66613
R5966 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t2 2.2755
R5967 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 2.2755
R5968 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 2.2505
R5969 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 1.80834
R5970 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 1.43706
R5971 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 0.281955
R5972 VCO_mag_0.VCONT.n45 VCO_mag_0.VCONT.t56 21.8873
R5973 VCO_mag_0.VCONT.n41 VCO_mag_0.VCONT.t51 21.8873
R5974 VCO_mag_0.VCONT.n38 VCO_mag_0.VCONT.t59 21.8873
R5975 VCO_mag_0.VCONT.n35 VCO_mag_0.VCONT.t50 21.8873
R5976 VCO_mag_0.VCONT.n46 VCO_mag_0.VCONT.n45 12.5576
R5977 VCO_mag_0.VCONT.n42 VCO_mag_0.VCONT.n41 12.5576
R5978 VCO_mag_0.VCONT.n39 VCO_mag_0.VCONT.n38 12.5576
R5979 VCO_mag_0.VCONT.n36 VCO_mag_0.VCONT.n35 12.5576
R5980 VCO_mag_0.VCONT.n47 VCO_mag_0.VCONT.t58 12.1889
R5981 VCO_mag_0.VCONT.n43 VCO_mag_0.VCONT.t52 12.1889
R5982 VCO_mag_0.VCONT.n40 VCO_mag_0.VCONT.t53 12.1889
R5983 VCO_mag_0.VCONT.n37 VCO_mag_0.VCONT.t47 12.1889
R5984 VCO_mag_0.VCONT.n47 VCO_mag_0.VCONT.n46 9.69888
R5985 VCO_mag_0.VCONT.n43 VCO_mag_0.VCONT.n42 9.69888
R5986 VCO_mag_0.VCONT.n40 VCO_mag_0.VCONT.n39 9.69888
R5987 VCO_mag_0.VCONT.n37 VCO_mag_0.VCONT.n36 9.69888
R5988 VCO_mag_0.VCONT.n49 VCO_mag_0.VCONT 9.06976
R5989 VCO_mag_0.VCONT.n44 VCO_mag_0.VCONT 8.99233
R5990 VCO_mag_0.VCONT.n50 VCO_mag_0.VCONT 6.57545
R5991 VCO_mag_0.VCONT.n45 VCO_mag_0.VCONT.t46 6.51836
R5992 VCO_mag_0.VCONT.n46 VCO_mag_0.VCONT.t44 6.51836
R5993 VCO_mag_0.VCONT.n41 VCO_mag_0.VCONT.t45 6.51836
R5994 VCO_mag_0.VCONT.n42 VCO_mag_0.VCONT.t55 6.51836
R5995 VCO_mag_0.VCONT.n38 VCO_mag_0.VCONT.t54 6.51836
R5996 VCO_mag_0.VCONT.n39 VCO_mag_0.VCONT.t48 6.51836
R5997 VCO_mag_0.VCONT.n35 VCO_mag_0.VCONT.t49 6.51836
R5998 VCO_mag_0.VCONT.n36 VCO_mag_0.VCONT.t57 6.51836
R5999 VCO_mag_0.VCONT.n31 VCO_mag_0.VCONT.n30 5.4005
R6000 VCO_mag_0.VCONT.n31 VCO_mag_0.VCONT.t10 5.4005
R6001 VCO_mag_0.VCONT.n50 VCO_mag_0.VCONT.n49 4.79502
R6002 VCO_mag_0.VCONT.n44 VCO_mag_0.VCONT 4.75244
R6003 VCO_mag_0.VCONT VCO_mag_0.VCONT.n47 4.63297
R6004 VCO_mag_0.VCONT VCO_mag_0.VCONT.n43 4.63297
R6005 VCO_mag_0.VCONT VCO_mag_0.VCONT.n40 4.63297
R6006 VCO_mag_0.VCONT VCO_mag_0.VCONT.n37 4.63297
R6007 VCO_mag_0.VCONT.n49 VCO_mag_0.VCONT.n48 4.50173
R6008 VCO_mag_0.VCONT.n34 VCO_mag_0.VCONT.n31 3.71064
R6009 VCO_mag_0.VCONT.n33 VCO_mag_0.VCONT.t21 3.6405
R6010 VCO_mag_0.VCONT.n33 VCO_mag_0.VCONT.n32 3.6405
R6011 VCO_mag_0.VCONT.n19 VCO_mag_0.VCONT.n18 3.16355
R6012 VCO_mag_0.VCONT.n75 VCO_mag_0.VCONT.n74 3.16355
R6013 VCO_mag_0.VCONT.n14 VCO_mag_0.VCONT.n13 3.15771
R6014 VCO_mag_0.VCONT.n9 VCO_mag_0.VCONT.n8 3.15771
R6015 VCO_mag_0.VCONT.n4 VCO_mag_0.VCONT.n3 3.15771
R6016 VCO_mag_0.VCONT.n60 VCO_mag_0.VCONT.n57 3.15771
R6017 VCO_mag_0.VCONT.n65 VCO_mag_0.VCONT.n62 3.15771
R6018 VCO_mag_0.VCONT.n70 VCO_mag_0.VCONT.n67 3.15771
R6019 VCO_mag_0.VCONT.n19 VCO_mag_0.VCONT.n16 3.15264
R6020 VCO_mag_0.VCONT.n75 VCO_mag_0.VCONT.n72 3.15264
R6021 VCO_mag_0.VCONT.n14 VCO_mag_0.VCONT.n11 3.1505
R6022 VCO_mag_0.VCONT.n9 VCO_mag_0.VCONT.n6 3.1505
R6023 VCO_mag_0.VCONT.n4 VCO_mag_0.VCONT.n1 3.1505
R6024 VCO_mag_0.VCONT.n25 VCO_mag_0.VCONT.n24 3.1505
R6025 VCO_mag_0.VCONT.n60 VCO_mag_0.VCONT.n59 3.1505
R6026 VCO_mag_0.VCONT.n65 VCO_mag_0.VCONT.n64 3.1505
R6027 VCO_mag_0.VCONT.n70 VCO_mag_0.VCONT.n69 3.1505
R6028 VCO_mag_0.VCONT.n79 VCO_mag_0.VCONT.n55 3.1505
R6029 VCO_mag_0.VCONT.n80 VCO_mag_0.VCONT.n53 2.93535
R6030 VCO_mag_0.VCONT.n28 VCO_mag_0.VCONT.n27 2.93403
R6031 VCO_mag_0.VCONT VCO_mag_0.VCONT.n50 2.64399
R6032 VCO_mag_0.VCONT.n81 VCO_mag_0.VCONT.n80 2.54229
R6033 VCO_mag_0.VCONT.n29 VCO_mag_0.VCONT.n28 2.54091
R6034 VCO_mag_0.VCONT.n51 VCO_mag_0.VCONT 2.36677
R6035 VCO_mag_0.VCONT.n49 VCO_mag_0.VCONT.n44 2.29048
R6036 VCO_mag_0.VCONT.n27 VCO_mag_0.VCONT.t26 1.8205
R6037 VCO_mag_0.VCONT.n27 VCO_mag_0.VCONT.n26 1.8205
R6038 VCO_mag_0.VCONT.n18 VCO_mag_0.VCONT.t27 1.8205
R6039 VCO_mag_0.VCONT.n18 VCO_mag_0.VCONT.n17 1.8205
R6040 VCO_mag_0.VCONT.n13 VCO_mag_0.VCONT.t25 1.8205
R6041 VCO_mag_0.VCONT.n13 VCO_mag_0.VCONT.n12 1.8205
R6042 VCO_mag_0.VCONT.n8 VCO_mag_0.VCONT.t24 1.8205
R6043 VCO_mag_0.VCONT.n8 VCO_mag_0.VCONT.n7 1.8205
R6044 VCO_mag_0.VCONT.n3 VCO_mag_0.VCONT.t28 1.8205
R6045 VCO_mag_0.VCONT.n3 VCO_mag_0.VCONT.n2 1.8205
R6046 VCO_mag_0.VCONT.n57 VCO_mag_0.VCONT.t6 1.8205
R6047 VCO_mag_0.VCONT.n57 VCO_mag_0.VCONT.n56 1.8205
R6048 VCO_mag_0.VCONT.n62 VCO_mag_0.VCONT.t7 1.8205
R6049 VCO_mag_0.VCONT.n62 VCO_mag_0.VCONT.n61 1.8205
R6050 VCO_mag_0.VCONT.n67 VCO_mag_0.VCONT.t8 1.8205
R6051 VCO_mag_0.VCONT.n67 VCO_mag_0.VCONT.n66 1.8205
R6052 VCO_mag_0.VCONT.n74 VCO_mag_0.VCONT.t5 1.8205
R6053 VCO_mag_0.VCONT.n74 VCO_mag_0.VCONT.n73 1.8205
R6054 VCO_mag_0.VCONT.n53 VCO_mag_0.VCONT.t9 1.8205
R6055 VCO_mag_0.VCONT.n53 VCO_mag_0.VCONT.n52 1.8205
R6056 VCO_mag_0.VCONT.n34 VCO_mag_0.VCONT.n33 1.6852
R6057 VCO_mag_0.VCONT.n24 VCO_mag_0.VCONT.t34 1.6385
R6058 VCO_mag_0.VCONT.n24 VCO_mag_0.VCONT.n23 1.6385
R6059 VCO_mag_0.VCONT.n16 VCO_mag_0.VCONT.t35 1.6385
R6060 VCO_mag_0.VCONT.n16 VCO_mag_0.VCONT.n15 1.6385
R6061 VCO_mag_0.VCONT.n11 VCO_mag_0.VCONT.t38 1.6385
R6062 VCO_mag_0.VCONT.n11 VCO_mag_0.VCONT.n10 1.6385
R6063 VCO_mag_0.VCONT.n6 VCO_mag_0.VCONT.t37 1.6385
R6064 VCO_mag_0.VCONT.n6 VCO_mag_0.VCONT.n5 1.6385
R6065 VCO_mag_0.VCONT.n1 VCO_mag_0.VCONT.t36 1.6385
R6066 VCO_mag_0.VCONT.n1 VCO_mag_0.VCONT.n0 1.6385
R6067 VCO_mag_0.VCONT.n55 VCO_mag_0.VCONT.t17 1.6385
R6068 VCO_mag_0.VCONT.n55 VCO_mag_0.VCONT.n54 1.6385
R6069 VCO_mag_0.VCONT.n59 VCO_mag_0.VCONT.t19 1.6385
R6070 VCO_mag_0.VCONT.n59 VCO_mag_0.VCONT.n58 1.6385
R6071 VCO_mag_0.VCONT.n64 VCO_mag_0.VCONT.t20 1.6385
R6072 VCO_mag_0.VCONT.n64 VCO_mag_0.VCONT.n63 1.6385
R6073 VCO_mag_0.VCONT.n69 VCO_mag_0.VCONT.t16 1.6385
R6074 VCO_mag_0.VCONT.n69 VCO_mag_0.VCONT.n68 1.6385
R6075 VCO_mag_0.VCONT.n72 VCO_mag_0.VCONT.t18 1.6385
R6076 VCO_mag_0.VCONT.n72 VCO_mag_0.VCONT.n71 1.6385
R6077 VCO_mag_0.VCONT VCO_mag_0.VCONT.n34 1.33738
R6078 VCO_mag_0.VCONT.n81 VCO_mag_0.VCONT.n51 0.773
R6079 VCO_mag_0.VCONT.n51 VCO_mag_0.VCONT.n29 0.74925
R6080 VCO_mag_0.VCONT.n25 VCO_mag_0.VCONT.n22 0.690059
R6081 VCO_mag_0.VCONT.n79 VCO_mag_0.VCONT.n78 0.690059
R6082 VCO_mag_0.VCONT.n20 VCO_mag_0.VCONT.n19 0.686845
R6083 VCO_mag_0.VCONT.n76 VCO_mag_0.VCONT.n75 0.686845
R6084 VCO_mag_0.VCONT.n21 VCO_mag_0.VCONT.n20 0.424029
R6085 VCO_mag_0.VCONT.n77 VCO_mag_0.VCONT.n76 0.424029
R6086 VCO_mag_0.VCONT.n22 VCO_mag_0.VCONT.n21 0.422706
R6087 VCO_mag_0.VCONT.n78 VCO_mag_0.VCONT.n77 0.422706
R6088 VCO_mag_0.VCONT.n20 VCO_mag_0.VCONT.n14 0.263882
R6089 VCO_mag_0.VCONT.n21 VCO_mag_0.VCONT.n9 0.263882
R6090 VCO_mag_0.VCONT.n22 VCO_mag_0.VCONT.n4 0.263882
R6091 VCO_mag_0.VCONT.n78 VCO_mag_0.VCONT.n60 0.263882
R6092 VCO_mag_0.VCONT.n77 VCO_mag_0.VCONT.n65 0.263882
R6093 VCO_mag_0.VCONT.n76 VCO_mag_0.VCONT.n70 0.263882
R6094 VCO_mag_0.VCONT.n48 VCO_mag_0.VCONT 0.244813
R6095 VCO_mag_0.VCONT.n28 VCO_mag_0.VCONT.n25 0.224176
R6096 VCO_mag_0.VCONT.n80 VCO_mag_0.VCONT.n79 0.222853
R6097 VCO_mag_0.VCONT.n29 VCO_mag_0.VCONT 0.0946163
R6098 VCO_mag_0.VCONT VCO_mag_0.VCONT.n81 0.093312
R6099 VCO_mag_0.VCONT.n48 VCO_mag_0.VCONT 0.0469095
R6100 a_67077_18370.t10 a_67077_18370.n5 22.8782
R6101 a_67077_18370.n6 a_67077_18370.t10 22.4219
R6102 a_67077_18370.n3 a_67077_18370.t17 22.2916
R6103 a_67077_18370.n5 a_67077_18370.n4 14.0791
R6104 a_67077_18370.n4 a_67077_18370.n3 14.0791
R6105 a_67077_18370.n7 a_67077_18370.n6 14.0791
R6106 a_67077_18370.n2 a_67077_18370.t8 11.3416
R6107 a_67077_18370.n6 a_67077_18370.t6 8.34336
R6108 a_67077_18370.n7 a_67077_18370.t4 8.34336
R6109 a_67077_18370.n5 a_67077_18370.t16 8.213
R6110 a_67077_18370.n4 a_67077_18370.t13 8.213
R6111 a_67077_18370.n3 a_67077_18370.t15 8.213
R6112 a_67077_18370.n0 a_67077_18370.n7 8.17193
R6113 a_67077_18370.n1 a_67077_18370.n2 4.0005
R6114 a_67077_18370.n0 a_67077_18370.n9 3.63045
R6115 a_67077_18370.n17 a_67077_18370.n1 2.89398
R6116 a_67077_18370.n14 a_67077_18370.n11 2.26392
R6117 a_67077_18370.n9 a_67077_18370.t11 1.8205
R6118 a_67077_18370.n9 a_67077_18370.n8 1.8205
R6119 a_67077_18370.n17 a_67077_18370.t5 1.8205
R6120 a_67077_18370.n18 a_67077_18370.n17 1.8205
R6121 a_67077_18370.n11 a_67077_18370.t2 1.6385
R6122 a_67077_18370.n11 a_67077_18370.n10 1.6385
R6123 a_67077_18370.n13 a_67077_18370.t0 1.6385
R6124 a_67077_18370.n13 a_67077_18370.n12 1.6385
R6125 a_67077_18370.n2 a_67077_18370.n16 1.62996
R6126 a_67077_18370.n14 a_67077_18370.n13 1.4936
R6127 a_67077_18370.n1 a_67077_18370.n15 1.22554
R6128 a_67077_18370.n15 a_67077_18370.n14 1.18673
R6129 a_67077_18370.n1 a_67077_18370.n0 0.1505
R6130 VCO_op_bar.n6 VCO_op_bar 12.4956
R6131 VCO_op_bar.n9 VCO_op_bar.n8 3.59137
R6132 VCO_op_bar.n10 VCO_op_bar.n3 3.58485
R6133 VCO_op_bar.n10 VCO_op_bar.n1 3.32833
R6134 VCO_op_bar.n6 VCO_op_bar.n5 3.28266
R6135 VCO_op_bar.n3 VCO_op_bar.t0 1.1705
R6136 VCO_op_bar.n3 VCO_op_bar.n2 1.1705
R6137 VCO_op_bar.n8 VCO_op_bar.t3 1.1705
R6138 VCO_op_bar.n8 VCO_op_bar.n7 1.1705
R6139 VCO_op_bar.n1 VCO_op_bar.t5 0.6505
R6140 VCO_op_bar.n1 VCO_op_bar.n0 0.6505
R6141 VCO_op_bar.n5 VCO_op_bar.t4 0.6505
R6142 VCO_op_bar.n5 VCO_op_bar.n4 0.6505
R6143 VCO_op_bar.n10 VCO_op_bar.n9 0.544413
R6144 VCO_op_bar VCO_op_bar.n10 0.297728
R6145 VCO_op_bar.n9 VCO_op_bar.n6 0.0142143
R6146 a_67077_14631.t2 a_67077_14631.n5 22.8782
R6147 a_67077_14631.n6 a_67077_14631.t2 22.4219
R6148 a_67077_14631.n3 a_67077_14631.t12 22.2916
R6149 a_67077_14631.n5 a_67077_14631.n4 14.0791
R6150 a_67077_14631.n4 a_67077_14631.n3 14.0791
R6151 a_67077_14631.n7 a_67077_14631.n6 14.0791
R6152 a_67077_14631.n1 a_67077_14631.t0 11.3416
R6153 a_67077_14631.n6 a_67077_14631.t6 8.34336
R6154 a_67077_14631.n7 a_67077_14631.t4 8.34336
R6155 a_67077_14631.n5 a_67077_14631.t17 8.213
R6156 a_67077_14631.n4 a_67077_14631.t14 8.213
R6157 a_67077_14631.n3 a_67077_14631.t15 8.213
R6158 a_67077_14631.n2 a_67077_14631.n7 8.17193
R6159 a_67077_14631.n0 a_67077_14631.n1 4.0005
R6160 a_67077_14631.n17 a_67077_14631.n2 3.63045
R6161 a_67077_14631.n0 a_67077_14631.n9 2.89398
R6162 a_67077_14631.n14 a_67077_14631.n11 2.26392
R6163 a_67077_14631.n9 a_67077_14631.t5 1.8205
R6164 a_67077_14631.n9 a_67077_14631.n8 1.8205
R6165 a_67077_14631.n17 a_67077_14631.t3 1.8205
R6166 a_67077_14631.n18 a_67077_14631.n17 1.8205
R6167 a_67077_14631.n11 a_67077_14631.t11 1.6385
R6168 a_67077_14631.n11 a_67077_14631.n10 1.6385
R6169 a_67077_14631.n13 a_67077_14631.t9 1.6385
R6170 a_67077_14631.n13 a_67077_14631.n12 1.6385
R6171 a_67077_14631.n1 a_67077_14631.n16 1.62996
R6172 a_67077_14631.n14 a_67077_14631.n13 1.4936
R6173 a_67077_14631.n0 a_67077_14631.n15 1.22554
R6174 a_67077_14631.n15 a_67077_14631.n14 1.18673
R6175 a_67077_14631.n2 a_67077_14631.n0 0.1505
R6176 RST_DIV.n4 RST_DIV.t9 36.935
R6177 RST_DIV.n57 RST_DIV.t15 36.935
R6178 RST_DIV.n14 RST_DIV.t3 36.935
R6179 RST_DIV.n47 RST_DIV.t5 36.935
R6180 RST_DIV.n33 RST_DIV.t12 36.935
R6181 RST_DIV.n31 RST_DIV.t2 36.935
R6182 RST_DIV.n27 RST_DIV.t6 36.935
R6183 RST_DIV.n37 RST_DIV.t11 36.935
R6184 RST_DIV.n4 RST_DIV.t8 18.1962
R6185 RST_DIV.n57 RST_DIV.t13 18.1962
R6186 RST_DIV.n14 RST_DIV.t1 18.1962
R6187 RST_DIV.n47 RST_DIV.t4 18.1962
R6188 RST_DIV.n33 RST_DIV.t0 18.1962
R6189 RST_DIV.n31 RST_DIV.t7 18.1962
R6190 RST_DIV.n37 RST_DIV.t14 18.1962
R6191 RST_DIV.n28 RST_DIV.t10 16.3712
R6192 RST_DIV.n29 RST_DIV.n28 8.0005
R6193 RST_DIV.n65 RST_DIV.n64 6.42884
R6194 RST_DIV.n35 RST_DIV.n34 5.39866
R6195 RST_DIV.n66 RST_DIV.n0 4.52907
R6196 RST_DIV.n21 RST_DIV.n20 4.51211
R6197 RST_DIV.n16 RST_DIV.n13 4.5005
R6198 RST_DIV.n16 RST_DIV.n15 4.5005
R6199 RST_DIV.n19 RST_DIV.n17 4.5005
R6200 RST_DIV.n23 RST_DIV.n22 4.5005
R6201 RST_DIV.n30 RST_DIV.n24 4.5005
R6202 RST_DIV.n30 RST_DIV.n29 4.5005
R6203 RST_DIV.n19 RST_DIV.n18 4.5005
R6204 RST_DIV.n36 RST_DIV.n35 3.52872
R6205 RST_DIV RST_DIV.n36 3.47469
R6206 RST_DIV.n7 RST_DIV.n6 2.2505
R6207 RST_DIV.n55 RST_DIV.n21 2.24707
R6208 RST_DIV.n34 RST_DIV.n33 2.13714
R6209 RST_DIV.n32 RST_DIV.n31 2.13714
R6210 RST_DIV.n38 RST_DIV.n37 2.1359
R6211 RST_DIV.n58 RST_DIV.n57 2.12318
R6212 RST_DIV.n15 RST_DIV.n14 2.12318
R6213 RST_DIV.n48 RST_DIV.n47 2.1224
R6214 RST_DIV.n5 RST_DIV.n4 2.12188
R6215 RST_DIV.n27 RST_DIV.n26 2.12075
R6216 RST_DIV.n62 RST_DIV.n56 1.88263
R6217 RST_DIV.n35 RST_DIV.n32 1.8704
R6218 RST_DIV.n54 RST_DIV.n53 1.86678
R6219 RST_DIV.n40 RST_DIV 1.83526
R6220 RST_DIV.n28 RST_DIV.n27 1.8255
R6221 RST_DIV.n39 RST_DIV.n38 1.76243
R6222 RST_DIV.n25 RST_DIV.n22 1.51223
R6223 RST_DIV.n50 RST_DIV.n49 1.5005
R6224 RST_DIV.n52 RST_DIV.n51 1.5005
R6225 RST_DIV.n10 RST_DIV.n9 1.5005
R6226 RST_DIV.n65 RST_DIV.n1 1.49919
R6227 RST_DIV.n64 RST_DIV.n63 1.18935
R6228 RST_DIV.n62 RST_DIV.n61 1.13307
R6229 RST_DIV.n36 RST_DIV.n30 1.1235
R6230 RST_DIV.n60 RST_DIV.n59 0.898107
R6231 RST_DIV.n41 RST_DIV.n40 0.839477
R6232 RST_DIV.n64 RST_DIV.n11 0.711378
R6233 RST_DIV.n42 RST_DIV.n41 0.627203
R6234 RST_DIV.n40 RST_DIV.n39 0.388998
R6235 RST_DIV.n38 RST_DIV 0.0687763
R6236 RST_DIV.n32 RST_DIV 0.0675415
R6237 RST_DIV.n34 RST_DIV 0.0675409
R6238 RST_DIV.n39 RST_DIV 0.0544779
R6239 RST_DIV.n59 RST_DIV 0.0518307
R6240 RST_DIV.n23 RST_DIV 0.0394837
R6241 RST_DIV.n25 RST_DIV.n24 0.0367013
R6242 RST_DIV.n46 RST_DIV 0.0363802
R6243 RST_DIV.n6 RST_DIV.n3 0.0361897
R6244 RST_DIV.n49 RST_DIV.n46 0.0346379
R6245 RST_DIV.n3 RST_DIV 0.031725
R6246 RST_DIV.n59 RST_DIV.n58 0.0249551
R6247 RST_DIV.n17 RST_DIV 0.0239664
R6248 RST_DIV.n16 RST_DIV.n12 0.0236959
R6249 RST_DIV.n11 RST_DIV.n10 0.0205676
R6250 RST_DIV.n53 RST_DIV.n52 0.0193514
R6251 RST_DIV.n51 RST_DIV.n44 0.0181289
R6252 RST_DIV.n55 RST_DIV.n54 0.0144865
R6253 RST_DIV.n21 RST_DIV.n19 0.0130264
R6254 RST_DIV.n6 RST_DIV.n5 0.0129138
R6255 RST_DIV.n63 RST_DIV.n62 0.0117735
R6256 RST_DIV.n7 RST_DIV.n2 0.0116103
R6257 RST_DIV.n66 RST_DIV.n65 0.00944245
R6258 RST_DIV.n49 RST_DIV.n48 0.00825862
R6259 RST_DIV.n56 RST_DIV.n55 0.0077973
R6260 RST_DIV.n26 RST_DIV.n25 0.00540913
R6261 RST_DIV.n9 RST_DIV.n8 0.00513918
R6262 RST_DIV.n50 RST_DIV.n45 0.00513918
R6263 RST_DIV.n1 RST_DIV.n0 0.00407143
R6264 RST_DIV.n30 RST_DIV.n22 0.003875
R6265 RST_DIV.n9 RST_DIV.n7 0.00328351
R6266 RST_DIV.n61 RST_DIV.n60 0.00328351
R6267 RST_DIV.n51 RST_DIV.n50 0.00328351
R6268 RST_DIV RST_DIV.n66 0.00253008
R6269 RST_DIV.n52 RST_DIV.n43 0.00232432
R6270 RST_DIV.n43 RST_DIV.n42 0.00232432
R6271 RST_DIV.n24 RST_DIV.n23 0.00205172
R6272 RST_DIV.n29 RST_DIV.n26 0.00173095
R6273 RST_DIV.n19 RST_DIV.n16 0.00142783
R6274 RST_DIV.n41 RST_DIV 0.00104041
R6275 EN EN.n1 60.8984
R6276 EN EN.n2 60.8974
R6277 EN EN.n0 60.897
R6278 EN EN.n5 60.8619
R6279 EN.n5 EN.t0 22.6826
R6280 EN.n0 EN.t2 22.6826
R6281 EN.n1 EN.t5 22.6826
R6282 EN.n2 EN.t1 22.6826
R6283 EN.n3 EN 9.24918
R6284 EN.n4 EN 9.00634
R6285 EN.n5 EN.t7 8.60407
R6286 EN.n0 EN.t6 8.60407
R6287 EN.n1 EN.t4 8.60407
R6288 EN.n2 EN.t3 8.60407
R6289 EN.n3 EN 4.52738
R6290 EN.n11 EN.n10 4.5243
R6291 EN.n7 EN.n6 4.5043
R6292 EN.n4 EN.n3 2.26677
R6293 EN.n9 EN.n8 1.12302
R6294 EN.n8 EN.n7 0.603745
R6295 EN.n7 EN.n4 0.173528
R6296 EN.n6 EN 0.1555
R6297 EN.n6 EN 0.0196667
R6298 EN.n11 EN.n8 0.00847126
R6299 EN.n10 EN.n9 0.00266346
R6300 EN EN.n11 0.00183663
R6301 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 37.1986
R6302 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 31.528
R6303 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 30.6344
R6304 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 27.3855
R6305 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 17.6614
R6306 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 15.3826
R6307 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 7.62751
R6308 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.09789
R6309 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 2.8877
R6310 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.67866
R6311 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 2.2505
R6312 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 1.43709
R6313 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.4325
R6314 LP_ext.n2 LP_ext.t17 5.34571
R6315 LP_ext.n28 LP_ext.n0 5.13526
R6316 LP_ext.n27 LP_ext.n1 4.4205
R6317 LP_ext.n2 LP_ext.t1 4.4205
R6318 LP_ext.n7 LP_ext.n4 3.70771
R6319 LP_ext.n13 LP_ext.n10 3.70771
R6320 LP_ext.n19 LP_ext.n16 3.70771
R6321 LP_ext.n25 LP_ext.n22 3.70771
R6322 LP_ext.n7 LP_ext.n6 2.6005
R6323 LP_ext.n13 LP_ext.n12 2.6005
R6324 LP_ext.n19 LP_ext.n18 2.6005
R6325 LP_ext.n25 LP_ext.n24 2.6005
R6326 LP_ext.n6 LP_ext.t9 1.8205
R6327 LP_ext.n6 LP_ext.n5 1.8205
R6328 LP_ext.n12 LP_ext.t6 1.8205
R6329 LP_ext.n12 LP_ext.n11 1.8205
R6330 LP_ext.n18 LP_ext.t5 1.8205
R6331 LP_ext.n18 LP_ext.n17 1.8205
R6332 LP_ext.n24 LP_ext.t2 1.8205
R6333 LP_ext.n24 LP_ext.n23 1.8205
R6334 LP_ext.n4 LP_ext.t15 1.6385
R6335 LP_ext.n4 LP_ext.n3 1.6385
R6336 LP_ext.n10 LP_ext.t12 1.6385
R6337 LP_ext.n10 LP_ext.n9 1.6385
R6338 LP_ext.n16 LP_ext.t11 1.6385
R6339 LP_ext.n16 LP_ext.n15 1.6385
R6340 LP_ext.n22 LP_ext.t18 1.6385
R6341 LP_ext.n22 LP_ext.n21 1.6385
R6342 LP_ext.n8 LP_ext.n2 0.600059
R6343 LP_ext.n27 LP_ext.n26 0.600059
R6344 LP_ext.n14 LP_ext.n8 0.361929
R6345 LP_ext.n26 LP_ext.n20 0.361929
R6346 LP_ext.n20 LP_ext.n14 0.359071
R6347 LP_ext LP_ext.n28 0.26819
R6348 LP_ext.n8 LP_ext.n7 0.240059
R6349 LP_ext.n14 LP_ext.n13 0.240059
R6350 LP_ext.n20 LP_ext.n19 0.240059
R6351 LP_ext.n26 LP_ext.n25 0.240059
R6352 LP_ext.n28 LP_ext.n27 0.120941
R6353 VCO_mag_0.Delay_Cell_mag_2.OUT.n13 VCO_mag_0.Delay_Cell_mag_2.OUT.t23 22.3568
R6354 VCO_mag_0.Delay_Cell_mag_2.OUT.n2 VCO_mag_0.Delay_Cell_mag_2.OUT.t8 22.096
R6355 VCO_mag_0.Delay_Cell_mag_2.OUT.n12 VCO_mag_0.Delay_Cell_mag_2.OUT.t18 19.4889
R6356 VCO_mag_0.Delay_Cell_mag_2.OUT.n25 VCO_mag_0.Delay_Cell_mag_2.OUT.t27 19.1891
R6357 VCO_mag_0.Delay_Cell_mag_2.OUT.n26 VCO_mag_0.Delay_Cell_mag_2.OUT.t16 19.1891
R6358 VCO_mag_0.Delay_Cell_mag_2.OUT.n27 VCO_mag_0.Delay_Cell_mag_2.OUT.t26 19.1891
R6359 VCO_mag_0.Delay_Cell_mag_2.OUT.n28 VCO_mag_0.Delay_Cell_mag_2.OUT.t22 18.6676
R6360 VCO_mag_0.Delay_Cell_mag_2.OUT.n26 VCO_mag_0.Delay_Cell_mag_2.OUT.n25 16.9365
R6361 VCO_mag_0.Delay_Cell_mag_2.OUT.n27 VCO_mag_0.Delay_Cell_mag_2.OUT.n26 16.9365
R6362 VCO_mag_0.Delay_Cell_mag_2.OUT.n28 VCO_mag_0.Delay_Cell_mag_2.OUT.n27 16.6457
R6363 VCO_mag_0.Delay_Cell_mag_2.OUT.n3 VCO_mag_0.Delay_Cell_mag_2.OUT.n2 14.0791
R6364 VCO_mag_0.Delay_Cell_mag_2.OUT.n4 VCO_mag_0.Delay_Cell_mag_2.OUT.n3 14.0791
R6365 VCO_mag_0.Delay_Cell_mag_2.OUT.n25 VCO_mag_0.Delay_Cell_mag_2.OUT.t24 11.6805
R6366 VCO_mag_0.Delay_Cell_mag_2.OUT.n26 VCO_mag_0.Delay_Cell_mag_2.OUT.t28 11.6805
R6367 VCO_mag_0.Delay_Cell_mag_2.OUT.n27 VCO_mag_0.Delay_Cell_mag_2.OUT.t21 11.6805
R6368 VCO_mag_0.Delay_Cell_mag_2.OUT.n28 VCO_mag_0.Delay_Cell_mag_2.OUT.t20 11.4719
R6369 VCO_mag_0.Delay_Cell_mag_2.OUT.n14 VCO_mag_0.Delay_Cell_mag_2.OUT.n13 9.33211
R6370 VCO_mag_0.Delay_Cell_mag_2.OUT.n13 VCO_mag_0.Delay_Cell_mag_2.OUT.t17 8.27818
R6371 VCO_mag_0.Delay_Cell_mag_2.OUT.n11 VCO_mag_0.Delay_Cell_mag_2.OUT.t19 8.27818
R6372 VCO_mag_0.Delay_Cell_mag_2.OUT.n2 VCO_mag_0.Delay_Cell_mag_2.OUT.t6 8.01746
R6373 VCO_mag_0.Delay_Cell_mag_2.OUT.n3 VCO_mag_0.Delay_Cell_mag_2.OUT.t12 8.01746
R6374 VCO_mag_0.Delay_Cell_mag_2.OUT.n4 VCO_mag_0.Delay_Cell_mag_2.OUT.t10 8.01746
R6375 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.OUT.n28 7.18457
R6376 VCO_mag_0.Delay_Cell_mag_2.OUT.n0 VCO_mag_0.Delay_Cell_mag_2.OUT 5.23607
R6377 VCO_mag_0.Delay_Cell_mag_2.OUT.n19 VCO_mag_0.Delay_Cell_mag_2.OUT.n18 4.67659
R6378 VCO_mag_0.Delay_Cell_mag_2.OUT.n1 VCO_mag_0.Delay_Cell_mag_2.OUT.n19 3.51328
R6379 VCO_mag_0.Delay_Cell_mag_2.OUT.n24 VCO_mag_0.Delay_Cell_mag_2.OUT.n23 3.20507
R6380 VCO_mag_0.Delay_Cell_mag_2.OUT.n19 VCO_mag_0.Delay_Cell_mag_2.OUT.n16 3.1505
R6381 VCO_mag_0.Delay_Cell_mag_2.OUT.n21 VCO_mag_0.Delay_Cell_mag_2.OUT.n8 3.02311
R6382 VCO_mag_0.Delay_Cell_mag_2.OUT.n24 VCO_mag_0.Delay_Cell_mag_2.OUT.n6 2.98985
R6383 VCO_mag_0.Delay_Cell_mag_2.OUT.n12 VCO_mag_0.Delay_Cell_mag_2.OUT.n11 2.86836
R6384 VCO_mag_0.Delay_Cell_mag_2.OUT.n0 VCO_mag_0.Delay_Cell_mag_2.OUT.n4 2.6373
R6385 VCO_mag_0.Delay_Cell_mag_2.OUT.n20 VCO_mag_0.Delay_Cell_mag_2.OUT.n10 2.6005
R6386 VCO_mag_0.Delay_Cell_mag_2.OUT.n1 VCO_mag_0.Delay_Cell_mag_2.OUT.n12 2.11815
R6387 VCO_mag_0.Delay_Cell_mag_2.OUT.n6 VCO_mag_0.Delay_Cell_mag_2.OUT.t13 1.8205
R6388 VCO_mag_0.Delay_Cell_mag_2.OUT.n6 VCO_mag_0.Delay_Cell_mag_2.OUT.n5 1.8205
R6389 VCO_mag_0.Delay_Cell_mag_2.OUT.n10 VCO_mag_0.Delay_Cell_mag_2.OUT.t1 1.8205
R6390 VCO_mag_0.Delay_Cell_mag_2.OUT.n10 VCO_mag_0.Delay_Cell_mag_2.OUT.n9 1.8205
R6391 VCO_mag_0.Delay_Cell_mag_2.OUT.n8 VCO_mag_0.Delay_Cell_mag_2.OUT.t9 1.8205
R6392 VCO_mag_0.Delay_Cell_mag_2.OUT.n8 VCO_mag_0.Delay_Cell_mag_2.OUT.n7 1.8205
R6393 VCO_mag_0.Delay_Cell_mag_2.OUT.n23 VCO_mag_0.Delay_Cell_mag_2.OUT.t3 1.8205
R6394 VCO_mag_0.Delay_Cell_mag_2.OUT.n23 VCO_mag_0.Delay_Cell_mag_2.OUT.n22 1.8205
R6395 VCO_mag_0.Delay_Cell_mag_2.OUT.n16 VCO_mag_0.Delay_Cell_mag_2.OUT.t15 1.6385
R6396 VCO_mag_0.Delay_Cell_mag_2.OUT.n16 VCO_mag_0.Delay_Cell_mag_2.OUT.n15 1.6385
R6397 VCO_mag_0.Delay_Cell_mag_2.OUT.n18 VCO_mag_0.Delay_Cell_mag_2.OUT.t5 1.6385
R6398 VCO_mag_0.Delay_Cell_mag_2.OUT.n18 VCO_mag_0.Delay_Cell_mag_2.OUT.n17 1.6385
R6399 VCO_mag_0.Delay_Cell_mag_2.OUT.n1 VCO_mag_0.Delay_Cell_mag_2.OUT.n14 1.50108
R6400 VCO_mag_0.Delay_Cell_mag_2.OUT.n20 VCO_mag_0.Delay_Cell_mag_2.OUT.n1 1.32596
R6401 VCO_mag_0.Delay_Cell_mag_2.OUT.n24 VCO_mag_0.Delay_Cell_mag_2.OUT.n21 0.826273
R6402 VCO_mag_0.Delay_Cell_mag_2.OUT.n21 VCO_mag_0.Delay_Cell_mag_2.OUT.n20 0.640283
R6403 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.OUT.n0 0.156737
R6404 VCO_mag_0.Delay_Cell_mag_2.OUT.n0 VCO_mag_0.Delay_Cell_mag_2.OUT.n24 0.128582
R6405 VCO_mag_0.Delay_Cell_mag_0.OUTB.n23 VCO_mag_0.Delay_Cell_mag_0.OUTB.t22 22.2916
R6406 VCO_mag_0.Delay_Cell_mag_0.OUTB.n9 VCO_mag_0.Delay_Cell_mag_0.OUTB.t6 22.1612
R6407 VCO_mag_0.Delay_Cell_mag_0.OUTB.n0 VCO_mag_0.Delay_Cell_mag_0.OUTB.t17 21.774
R6408 VCO_mag_0.Delay_Cell_mag_0.OUTB.t22 VCO_mag_0.Delay_Cell_mag_0.OUTB.n22 17.311
R6409 VCO_mag_0.Delay_Cell_mag_0.OUTB.n11 VCO_mag_0.Delay_Cell_mag_0.OUTB.t8 15.1219
R6410 VCO_mag_0.Delay_Cell_mag_0.OUTB.n10 VCO_mag_0.Delay_Cell_mag_0.OUTB.n9 14.0791
R6411 VCO_mag_0.Delay_Cell_mag_0.OUTB.n24 VCO_mag_0.Delay_Cell_mag_0.OUTB.n23 14.0791
R6412 VCO_mag_0.Delay_Cell_mag_0.OUTB.n25 VCO_mag_0.Delay_Cell_mag_0.OUTB.n24 14.0791
R6413 VCO_mag_0.Delay_Cell_mag_0.OUTB.n1 VCO_mag_0.Delay_Cell_mag_0.OUTB.n0 12.7222
R6414 VCO_mag_0.Delay_Cell_mag_0.OUTB.n2 VCO_mag_0.Delay_Cell_mag_0.OUTB.t19 11.6444
R6415 VCO_mag_0.Delay_Cell_mag_0.OUTB.n2 VCO_mag_0.Delay_Cell_mag_0.OUTB.n1 10.0261
R6416 VCO_mag_0.Delay_Cell_mag_0.OUTB.n23 VCO_mag_0.Delay_Cell_mag_0.OUTB.t18 8.213
R6417 VCO_mag_0.Delay_Cell_mag_0.OUTB.n24 VCO_mag_0.Delay_Cell_mag_0.OUTB.t16 8.213
R6418 VCO_mag_0.Delay_Cell_mag_0.OUTB.n25 VCO_mag_0.Delay_Cell_mag_0.OUTB.t20 8.213
R6419 VCO_mag_0.Delay_Cell_mag_0.OUTB.n10 VCO_mag_0.Delay_Cell_mag_0.OUTB.t4 8.08264
R6420 VCO_mag_0.Delay_Cell_mag_0.OUTB.n9 VCO_mag_0.Delay_Cell_mag_0.OUTB.t10 8.08264
R6421 VCO_mag_0.Delay_Cell_mag_0.OUTB.n11 VCO_mag_0.Delay_Cell_mag_0.OUTB.n10 7.03979
R6422 VCO_mag_0.Delay_Cell_mag_0.OUTB.n0 VCO_mag_0.Delay_Cell_mag_0.OUTB.t25 6.51836
R6423 VCO_mag_0.Delay_Cell_mag_0.OUTB.n1 VCO_mag_0.Delay_Cell_mag_0.OUTB.t24 6.51836
R6424 VCO_mag_0.Delay_Cell_mag_0.OUTB.n17 VCO_mag_0.Delay_Cell_mag_0.OUTB.n16 4.70398
R6425 VCO_mag_0.Delay_Cell_mag_0.OUTB.n20 VCO_mag_0.Delay_Cell_mag_0.OUTB.n17 4.4843
R6426 VCO_mag_0.Delay_Cell_mag_0.OUTB.n12 VCO_mag_0.Delay_Cell_mag_0.OUTB.n11 4.0005
R6427 VCO_mag_0.Delay_Cell_mag_0.OUTB.n22 VCO_mag_0.Delay_Cell_mag_0.OUTB.n4 3.3342
R6428 VCO_mag_0.Delay_Cell_mag_0.OUTB.n17 VCO_mag_0.Delay_Cell_mag_0.OUTB.n14 3.1505
R6429 VCO_mag_0.Delay_Cell_mag_0.OUTB.n12 VCO_mag_0.Delay_Cell_mag_0.OUTB.n8 2.94411
R6430 VCO_mag_0.Delay_Cell_mag_0.OUTB.n22 VCO_mag_0.Delay_Cell_mag_0.OUTB.n6 2.9292
R6431 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.OUTB.n25 2.70614
R6432 VCO_mag_0.Delay_Cell_mag_0.OUTB.n20 VCO_mag_0.Delay_Cell_mag_0.OUTB.n19 2.6005
R6433 VCO_mag_0.Delay_Cell_mag_0.OUTB.n8 VCO_mag_0.Delay_Cell_mag_0.OUTB.t9 1.8205
R6434 VCO_mag_0.Delay_Cell_mag_0.OUTB.n8 VCO_mag_0.Delay_Cell_mag_0.OUTB.n7 1.8205
R6435 VCO_mag_0.Delay_Cell_mag_0.OUTB.n6 VCO_mag_0.Delay_Cell_mag_0.OUTB.t0 1.8205
R6436 VCO_mag_0.Delay_Cell_mag_0.OUTB.n6 VCO_mag_0.Delay_Cell_mag_0.OUTB.n5 1.8205
R6437 VCO_mag_0.Delay_Cell_mag_0.OUTB.n4 VCO_mag_0.Delay_Cell_mag_0.OUTB.t11 1.8205
R6438 VCO_mag_0.Delay_Cell_mag_0.OUTB.n4 VCO_mag_0.Delay_Cell_mag_0.OUTB.n3 1.8205
R6439 VCO_mag_0.Delay_Cell_mag_0.OUTB.n19 VCO_mag_0.Delay_Cell_mag_0.OUTB.t3 1.8205
R6440 VCO_mag_0.Delay_Cell_mag_0.OUTB.n19 VCO_mag_0.Delay_Cell_mag_0.OUTB.n18 1.8205
R6441 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.OUTB.n2 1.77023
R6442 VCO_mag_0.Delay_Cell_mag_0.OUTB.n14 VCO_mag_0.Delay_Cell_mag_0.OUTB.t13 1.6385
R6443 VCO_mag_0.Delay_Cell_mag_0.OUTB.n14 VCO_mag_0.Delay_Cell_mag_0.OUTB.n13 1.6385
R6444 VCO_mag_0.Delay_Cell_mag_0.OUTB.n16 VCO_mag_0.Delay_Cell_mag_0.OUTB.t12 1.6385
R6445 VCO_mag_0.Delay_Cell_mag_0.OUTB.n16 VCO_mag_0.Delay_Cell_mag_0.OUTB.n15 1.6385
R6446 VCO_mag_0.Delay_Cell_mag_0.OUTB.n22 VCO_mag_0.Delay_Cell_mag_0.OUTB.n21 0.845717
R6447 VCO_mag_0.Delay_Cell_mag_0.OUTB.n21 VCO_mag_0.Delay_Cell_mag_0.OUTB.n12 0.335065
R6448 VCO_mag_0.Delay_Cell_mag_0.OUTB.n21 VCO_mag_0.Delay_Cell_mag_0.OUTB.n20 0.329196
R6449 pd.n0 pd.t8 18.5164
R6450 pd.n11 pd.n0 5.96897
R6451 pd.n0 pd.t9 4.95003
R6452 pd.n5 pd.n4 3.416
R6453 pd.n10 pd.n9 3.416
R6454 pd.n4 pd.t2 3.2765
R6455 pd.n4 pd.n3 3.2765
R6456 pd.n9 pd.t0 3.2765
R6457 pd.n9 pd.n8 3.2765
R6458 pd.n5 pd.n2 3.013
R6459 pd.n10 pd.n7 3.013
R6460 pd.n11 pd 2.83268
R6461 pd.n2 pd.t7 1.8205
R6462 pd.n2 pd.n1 1.8205
R6463 pd.n7 pd.t6 1.8205
R6464 pd.n7 pd.n6 1.8205
R6465 pd.n10 pd.n5 0.445308
R6466 pd pd.n10 0.310308
R6467 pd pd.n11 0.0166053
R6468 LF_mag_0.VCNTL LF_mag_0.VCNTL.n0 17.1693
R6469 LF_mag_0.VCNTL.n0 LF_mag_0.VCNTL 9.27059
R6470 LF_mag_0.VCNTL LF_mag_0.VCNTL.t20 7.13043
R6471 LF_mag_0.VCNTL.n7 LF_mag_0.VCNTL.t11 5.34571
R6472 LF_mag_0.VCNTL.n29 LF_mag_0.VCNTL.n1 5.13526
R6473 LF_mag_0.VCNTL.n28 LF_mag_0.VCNTL.n27 4.4205
R6474 LF_mag_0.VCNTL.n7 LF_mag_0.VCNTL.t7 4.4205
R6475 LF_mag_0.VCNTL.n6 LF_mag_0.VCNTL.n5 3.70771
R6476 LF_mag_0.VCNTL.n12 LF_mag_0.VCNTL.n11 3.70771
R6477 LF_mag_0.VCNTL.n18 LF_mag_0.VCNTL.n17 3.70771
R6478 LF_mag_0.VCNTL.n24 LF_mag_0.VCNTL.n21 3.70771
R6479 LF_mag_0.VCNTL.n6 LF_mag_0.VCNTL.n3 2.6005
R6480 LF_mag_0.VCNTL.n12 LF_mag_0.VCNTL.n9 2.6005
R6481 LF_mag_0.VCNTL.n18 LF_mag_0.VCNTL.n15 2.6005
R6482 LF_mag_0.VCNTL.n24 LF_mag_0.VCNTL.n23 2.6005
R6483 LF_mag_0.VCNTL LF_mag_0.VCNTL.t21 2.35318
R6484 LF_mag_0.VCNTL.n3 LF_mag_0.VCNTL.t5 1.8205
R6485 LF_mag_0.VCNTL.n3 LF_mag_0.VCNTL.n2 1.8205
R6486 LF_mag_0.VCNTL.n9 LF_mag_0.VCNTL.t3 1.8205
R6487 LF_mag_0.VCNTL.n9 LF_mag_0.VCNTL.n8 1.8205
R6488 LF_mag_0.VCNTL.n15 LF_mag_0.VCNTL.t0 1.8205
R6489 LF_mag_0.VCNTL.n15 LF_mag_0.VCNTL.n14 1.8205
R6490 LF_mag_0.VCNTL.n23 LF_mag_0.VCNTL.t9 1.8205
R6491 LF_mag_0.VCNTL.n23 LF_mag_0.VCNTL.n22 1.8205
R6492 LF_mag_0.VCNTL.n21 LF_mag_0.VCNTL.t13 1.6385
R6493 LF_mag_0.VCNTL.n21 LF_mag_0.VCNTL.n20 1.6385
R6494 LF_mag_0.VCNTL.n5 LF_mag_0.VCNTL.t19 1.6385
R6495 LF_mag_0.VCNTL.n5 LF_mag_0.VCNTL.n4 1.6385
R6496 LF_mag_0.VCNTL.n11 LF_mag_0.VCNTL.t17 1.6385
R6497 LF_mag_0.VCNTL.n11 LF_mag_0.VCNTL.n10 1.6385
R6498 LF_mag_0.VCNTL.n17 LF_mag_0.VCNTL.t14 1.6385
R6499 LF_mag_0.VCNTL.n17 LF_mag_0.VCNTL.n16 1.6385
R6500 LF_mag_0.VCNTL.n28 LF_mag_0.VCNTL.n26 0.598735
R6501 LF_mag_0.VCNTL.n13 LF_mag_0.VCNTL.n7 0.598735
R6502 LF_mag_0.VCNTL.n19 LF_mag_0.VCNTL.n13 0.361929
R6503 LF_mag_0.VCNTL.n26 LF_mag_0.VCNTL.n25 0.361929
R6504 LF_mag_0.VCNTL.n25 LF_mag_0.VCNTL.n19 0.359071
R6505 LF_mag_0.VCNTL LF_mag_0.VCNTL.n29 0.296971
R6506 LF_mag_0.VCNTL.n26 LF_mag_0.VCNTL.n6 0.238735
R6507 LF_mag_0.VCNTL.n13 LF_mag_0.VCNTL.n12 0.238735
R6508 LF_mag_0.VCNTL.n19 LF_mag_0.VCNTL.n18 0.238735
R6509 LF_mag_0.VCNTL.n25 LF_mag_0.VCNTL.n24 0.238735
R6510 LF_mag_0.VCNTL.n0 LF_mag_0.VCNTL 0.222567
R6511 LF_mag_0.VCNTL.n29 LF_mag_0.VCNTL.n28 0.120941
R6512 IPD+.n2 IPD+.t6 19.4169
R6513 IPD+.n3 IPD+.n2 14.623
R6514 IPD+.n4 IPD+.t0 11.2885
R6515 IPD+.n4 IPD+.n3 6.54523
R6516 IPD+.n1 IPD+.n0 5.4005
R6517 IPD+.n1 IPD+.t3 5.4005
R6518 IPD+.n5 IPD+.n4 4.10208
R6519 IPD+.n6 IPD+ 2.28854
R6520 IPD+.n5 IPD+.n1 1.84943
R6521 IPD+.n6 IPD+.n5 1.84768
R6522 IPD+.n2 IPD+.t4 1.8255
R6523 IPD+.n3 IPD+.t2 1.8255
R6524 IPD+ IPD+.n6 0.022768
R6525 VCO_mag_0.Delay_Cell_mag_1.INB.n13 VCO_mag_0.Delay_Cell_mag_1.INB.t20 22.3568
R6526 VCO_mag_0.Delay_Cell_mag_1.INB.n2 VCO_mag_0.Delay_Cell_mag_1.INB.t2 22.096
R6527 VCO_mag_0.Delay_Cell_mag_1.INB.n25 VCO_mag_0.Delay_Cell_mag_1.INB.t26 21.8182
R6528 VCO_mag_0.Delay_Cell_mag_1.INB.n12 VCO_mag_0.Delay_Cell_mag_1.INB.t24 19.4889
R6529 VCO_mag_0.Delay_Cell_mag_1.INB.n28 VCO_mag_0.Delay_Cell_mag_1.INB.t23 17.2487
R6530 VCO_mag_0.Delay_Cell_mag_1.INB.n3 VCO_mag_0.Delay_Cell_mag_1.INB.n2 14.0791
R6531 VCO_mag_0.Delay_Cell_mag_1.INB.n4 VCO_mag_0.Delay_Cell_mag_1.INB.n3 14.0791
R6532 VCO_mag_0.Delay_Cell_mag_1.INB.n26 VCO_mag_0.Delay_Cell_mag_1.INB.n25 12.6801
R6533 VCO_mag_0.Delay_Cell_mag_1.INB.n28 VCO_mag_0.Delay_Cell_mag_1.INB.t27 12.2493
R6534 VCO_mag_0.Delay_Cell_mag_1.INB.n27 VCO_mag_0.Delay_Cell_mag_1.INB.t22 12.0585
R6535 VCO_mag_0.Delay_Cell_mag_1.INB.n27 VCO_mag_0.Delay_Cell_mag_1.INB.n26 9.76014
R6536 VCO_mag_0.Delay_Cell_mag_1.INB.n14 VCO_mag_0.Delay_Cell_mag_1.INB.n13 9.33211
R6537 VCO_mag_0.Delay_Cell_mag_1.INB.n13 VCO_mag_0.Delay_Cell_mag_1.INB.t25 8.27818
R6538 VCO_mag_0.Delay_Cell_mag_1.INB.n11 VCO_mag_0.Delay_Cell_mag_1.INB.t18 8.27818
R6539 VCO_mag_0.Delay_Cell_mag_1.INB.n2 VCO_mag_0.Delay_Cell_mag_1.INB.t6 8.01746
R6540 VCO_mag_0.Delay_Cell_mag_1.INB.n3 VCO_mag_0.Delay_Cell_mag_1.INB.t0 8.01746
R6541 VCO_mag_0.Delay_Cell_mag_1.INB.n4 VCO_mag_0.Delay_Cell_mag_1.INB.t4 8.01746
R6542 VCO_mag_0.Delay_Cell_mag_1.INB.n25 VCO_mag_0.Delay_Cell_mag_1.INB.t19 6.51836
R6543 VCO_mag_0.Delay_Cell_mag_1.INB.n26 VCO_mag_0.Delay_Cell_mag_1.INB.t16 6.51836
R6544 VCO_mag_0.Delay_Cell_mag_1.INB.n19 VCO_mag_0.Delay_Cell_mag_1.INB.n18 4.67659
R6545 VCO_mag_0.Delay_Cell_mag_1.INB.n29 VCO_mag_0.Delay_Cell_mag_1.INB 4.34457
R6546 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_1.INB.n28 4.1467
R6547 VCO_mag_0.Delay_Cell_mag_1.INB.n29 VCO_mag_0.Delay_Cell_mag_1.INB 4.06926
R6548 VCO_mag_0.Delay_Cell_mag_1.INB.n0 VCO_mag_0.Delay_Cell_mag_1.INB.n19 3.51328
R6549 VCO_mag_0.Delay_Cell_mag_1.INB.n24 VCO_mag_0.Delay_Cell_mag_1.INB.n8 3.20507
R6550 VCO_mag_0.Delay_Cell_mag_1.INB.n19 VCO_mag_0.Delay_Cell_mag_1.INB.n16 3.1505
R6551 VCO_mag_0.Delay_Cell_mag_1.INB.n23 VCO_mag_0.Delay_Cell_mag_1.INB.n22 3.02311
R6552 VCO_mag_0.Delay_Cell_mag_1.INB.n24 VCO_mag_0.Delay_Cell_mag_1.INB.n6 2.98985
R6553 VCO_mag_0.Delay_Cell_mag_1.INB.n12 VCO_mag_0.Delay_Cell_mag_1.INB.n11 2.86836
R6554 VCO_mag_0.Delay_Cell_mag_1.INB.n1 VCO_mag_0.Delay_Cell_mag_1.INB.n4 2.63789
R6555 VCO_mag_0.Delay_Cell_mag_1.INB.n20 VCO_mag_0.Delay_Cell_mag_1.INB.n10 2.6005
R6556 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_1.INB.n27 2.55586
R6557 VCO_mag_0.Delay_Cell_mag_1.INB.n1 VCO_mag_0.Delay_Cell_mag_1.INB.n29 2.17974
R6558 VCO_mag_0.Delay_Cell_mag_1.INB.n0 VCO_mag_0.Delay_Cell_mag_1.INB.n12 2.11815
R6559 VCO_mag_0.Delay_Cell_mag_1.INB.n10 VCO_mag_0.Delay_Cell_mag_1.INB.t8 1.8205
R6560 VCO_mag_0.Delay_Cell_mag_1.INB.n10 VCO_mag_0.Delay_Cell_mag_1.INB.n9 1.8205
R6561 VCO_mag_0.Delay_Cell_mag_1.INB.n8 VCO_mag_0.Delay_Cell_mag_1.INB.t11 1.8205
R6562 VCO_mag_0.Delay_Cell_mag_1.INB.n8 VCO_mag_0.Delay_Cell_mag_1.INB.n7 1.8205
R6563 VCO_mag_0.Delay_Cell_mag_1.INB.n6 VCO_mag_0.Delay_Cell_mag_1.INB.t1 1.8205
R6564 VCO_mag_0.Delay_Cell_mag_1.INB.n6 VCO_mag_0.Delay_Cell_mag_1.INB.n5 1.8205
R6565 VCO_mag_0.Delay_Cell_mag_1.INB.n22 VCO_mag_0.Delay_Cell_mag_1.INB.t3 1.8205
R6566 VCO_mag_0.Delay_Cell_mag_1.INB.n22 VCO_mag_0.Delay_Cell_mag_1.INB.n21 1.8205
R6567 VCO_mag_0.Delay_Cell_mag_1.INB.n16 VCO_mag_0.Delay_Cell_mag_1.INB.t14 1.6385
R6568 VCO_mag_0.Delay_Cell_mag_1.INB.n16 VCO_mag_0.Delay_Cell_mag_1.INB.n15 1.6385
R6569 VCO_mag_0.Delay_Cell_mag_1.INB.n18 VCO_mag_0.Delay_Cell_mag_1.INB.t12 1.6385
R6570 VCO_mag_0.Delay_Cell_mag_1.INB.n18 VCO_mag_0.Delay_Cell_mag_1.INB.n17 1.6385
R6571 VCO_mag_0.Delay_Cell_mag_1.INB.n0 VCO_mag_0.Delay_Cell_mag_1.INB.n14 1.50108
R6572 VCO_mag_0.Delay_Cell_mag_1.INB.n20 VCO_mag_0.Delay_Cell_mag_1.INB.n0 1.32596
R6573 VCO_mag_0.Delay_Cell_mag_1.INB.n24 VCO_mag_0.Delay_Cell_mag_1.INB.n23 0.826273
R6574 VCO_mag_0.Delay_Cell_mag_1.INB.n23 VCO_mag_0.Delay_Cell_mag_1.INB.n20 0.640283
R6575 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_1.INB.n1 0.16328
R6576 VCO_mag_0.Delay_Cell_mag_1.INB.n1 VCO_mag_0.Delay_Cell_mag_1.INB.n24 0.123037
R6577 VCO_mag_0.Delay_Cell_mag_2.IN.n20 VCO_mag_0.Delay_Cell_mag_2.IN.t20 22.2916
R6578 VCO_mag_0.Delay_Cell_mag_2.IN.n4 VCO_mag_0.Delay_Cell_mag_2.IN.t10 22.1612
R6579 VCO_mag_0.Delay_Cell_mag_2.IN.n23 VCO_mag_0.Delay_Cell_mag_2.IN.t17 21.774
R6580 VCO_mag_0.Delay_Cell_mag_2.IN.t20 VCO_mag_0.Delay_Cell_mag_2.IN.n19 17.311
R6581 VCO_mag_0.Delay_Cell_mag_2.IN.n6 VCO_mag_0.Delay_Cell_mag_2.IN.t14 15.1219
R6582 VCO_mag_0.Delay_Cell_mag_2.IN.n21 VCO_mag_0.Delay_Cell_mag_2.IN.n20 14.0791
R6583 VCO_mag_0.Delay_Cell_mag_2.IN.n22 VCO_mag_0.Delay_Cell_mag_2.IN.n21 14.0791
R6584 VCO_mag_0.Delay_Cell_mag_2.IN.n5 VCO_mag_0.Delay_Cell_mag_2.IN.n4 14.0791
R6585 VCO_mag_0.Delay_Cell_mag_2.IN.n24 VCO_mag_0.Delay_Cell_mag_2.IN.n23 12.7222
R6586 VCO_mag_0.Delay_Cell_mag_2.IN.n25 VCO_mag_0.Delay_Cell_mag_2.IN.t18 11.9934
R6587 VCO_mag_0.Delay_Cell_mag_2.IN.n25 VCO_mag_0.Delay_Cell_mag_2.IN.n24 9.78115
R6588 VCO_mag_0.Delay_Cell_mag_2.IN.n20 VCO_mag_0.Delay_Cell_mag_2.IN.t23 8.213
R6589 VCO_mag_0.Delay_Cell_mag_2.IN.n21 VCO_mag_0.Delay_Cell_mag_2.IN.t16 8.213
R6590 VCO_mag_0.Delay_Cell_mag_2.IN.n22 VCO_mag_0.Delay_Cell_mag_2.IN.t19 8.213
R6591 VCO_mag_0.Delay_Cell_mag_2.IN.n5 VCO_mag_0.Delay_Cell_mag_2.IN.t12 8.08264
R6592 VCO_mag_0.Delay_Cell_mag_2.IN.n4 VCO_mag_0.Delay_Cell_mag_2.IN.t8 8.08264
R6593 VCO_mag_0.Delay_Cell_mag_2.IN.n6 VCO_mag_0.Delay_Cell_mag_2.IN.n5 7.03979
R6594 VCO_mag_0.Delay_Cell_mag_2.IN.n23 VCO_mag_0.Delay_Cell_mag_2.IN.t25 6.51836
R6595 VCO_mag_0.Delay_Cell_mag_2.IN.n24 VCO_mag_0.Delay_Cell_mag_2.IN.t21 6.51836
R6596 VCO_mag_0.Delay_Cell_mag_2.IN.n14 VCO_mag_0.Delay_Cell_mag_2.IN.n13 4.70398
R6597 VCO_mag_0.Delay_Cell_mag_2.IN.n15 VCO_mag_0.Delay_Cell_mag_2.IN.n14 4.4843
R6598 VCO_mag_0.Delay_Cell_mag_2.IN.n7 VCO_mag_0.Delay_Cell_mag_2.IN.n6 4.0005
R6599 VCO_mag_0.Delay_Cell_mag_2.IN.n19 VCO_mag_0.Delay_Cell_mag_2.IN.n1 3.3342
R6600 VCO_mag_0.Delay_Cell_mag_2.IN.n14 VCO_mag_0.Delay_Cell_mag_2.IN.n11 3.1505
R6601 VCO_mag_0.Delay_Cell_mag_2.IN.n7 VCO_mag_0.Delay_Cell_mag_2.IN.n3 2.94411
R6602 VCO_mag_0.Delay_Cell_mag_2.IN.n19 VCO_mag_0.Delay_Cell_mag_2.IN.n18 2.9292
R6603 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_2.IN.n22 2.69696
R6604 VCO_mag_0.Delay_Cell_mag_2.IN.n15 VCO_mag_0.Delay_Cell_mag_2.IN.n9 2.6005
R6605 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_2.IN.n25 2.10481
R6606 VCO_mag_0.Delay_Cell_mag_2.IN.n1 VCO_mag_0.Delay_Cell_mag_2.IN.t9 1.8205
R6607 VCO_mag_0.Delay_Cell_mag_2.IN.n1 VCO_mag_0.Delay_Cell_mag_2.IN.n0 1.8205
R6608 VCO_mag_0.Delay_Cell_mag_2.IN.n9 VCO_mag_0.Delay_Cell_mag_2.IN.t2 1.8205
R6609 VCO_mag_0.Delay_Cell_mag_2.IN.n9 VCO_mag_0.Delay_Cell_mag_2.IN.n8 1.8205
R6610 VCO_mag_0.Delay_Cell_mag_2.IN.n3 VCO_mag_0.Delay_Cell_mag_2.IN.t15 1.8205
R6611 VCO_mag_0.Delay_Cell_mag_2.IN.n3 VCO_mag_0.Delay_Cell_mag_2.IN.n2 1.8205
R6612 VCO_mag_0.Delay_Cell_mag_2.IN.n18 VCO_mag_0.Delay_Cell_mag_2.IN.t3 1.8205
R6613 VCO_mag_0.Delay_Cell_mag_2.IN.n18 VCO_mag_0.Delay_Cell_mag_2.IN.n17 1.8205
R6614 VCO_mag_0.Delay_Cell_mag_2.IN.n11 VCO_mag_0.Delay_Cell_mag_2.IN.t6 1.6385
R6615 VCO_mag_0.Delay_Cell_mag_2.IN.n11 VCO_mag_0.Delay_Cell_mag_2.IN.n10 1.6385
R6616 VCO_mag_0.Delay_Cell_mag_2.IN.n13 VCO_mag_0.Delay_Cell_mag_2.IN.t5 1.6385
R6617 VCO_mag_0.Delay_Cell_mag_2.IN.n13 VCO_mag_0.Delay_Cell_mag_2.IN.n12 1.6385
R6618 VCO_mag_0.Delay_Cell_mag_2.IN.n19 VCO_mag_0.Delay_Cell_mag_2.IN.n16 0.845717
R6619 VCO_mag_0.Delay_Cell_mag_2.IN.n16 VCO_mag_0.Delay_Cell_mag_2.IN.n7 0.335065
R6620 VCO_mag_0.Delay_Cell_mag_2.IN.n16 VCO_mag_0.Delay_Cell_mag_2.IN.n15 0.329196
R6621 a_60634_14631.t6 a_60634_14631.n5 22.8782
R6622 a_60634_14631.n6 a_60634_14631.t6 22.4219
R6623 a_60634_14631.n3 a_60634_14631.t16 22.2916
R6624 a_60634_14631.n5 a_60634_14631.n4 14.0791
R6625 a_60634_14631.n4 a_60634_14631.n3 14.0791
R6626 a_60634_14631.n7 a_60634_14631.n6 14.0791
R6627 a_60634_14631.n1 a_60634_14631.t8 11.3416
R6628 a_60634_14631.n6 a_60634_14631.t10 8.34336
R6629 a_60634_14631.n7 a_60634_14631.t4 8.34336
R6630 a_60634_14631.n5 a_60634_14631.t17 8.213
R6631 a_60634_14631.n4 a_60634_14631.t15 8.213
R6632 a_60634_14631.n3 a_60634_14631.t12 8.213
R6633 a_60634_14631.n2 a_60634_14631.n7 8.17193
R6634 a_60634_14631.n0 a_60634_14631.n1 4.0005
R6635 a_60634_14631.n17 a_60634_14631.n2 3.63045
R6636 a_60634_14631.n0 a_60634_14631.n9 2.89398
R6637 a_60634_14631.n14 a_60634_14631.n11 2.26392
R6638 a_60634_14631.n9 a_60634_14631.t5 1.8205
R6639 a_60634_14631.n9 a_60634_14631.n8 1.8205
R6640 a_60634_14631.n17 a_60634_14631.t7 1.8205
R6641 a_60634_14631.n18 a_60634_14631.n17 1.8205
R6642 a_60634_14631.n11 a_60634_14631.t1 1.6385
R6643 a_60634_14631.n11 a_60634_14631.n10 1.6385
R6644 a_60634_14631.n13 a_60634_14631.t2 1.6385
R6645 a_60634_14631.n13 a_60634_14631.n12 1.6385
R6646 a_60634_14631.n1 a_60634_14631.n16 1.62996
R6647 a_60634_14631.n14 a_60634_14631.n13 1.4936
R6648 a_60634_14631.n0 a_60634_14631.n15 1.22554
R6649 a_60634_14631.n15 a_60634_14631.n14 1.18673
R6650 a_60634_14631.n2 a_60634_14631.n0 0.1505
R6651 pu.n0 pu.t8 25.4398
R6652 pu.n0 pu.t9 17.6975
R6653 pu pu.n0 4.24451
R6654 pu.n5 pu.n4 3.416
R6655 pu.n10 pu.n9 3.416
R6656 pu.n4 pu.t0 3.2765
R6657 pu.n4 pu.n3 3.2765
R6658 pu.n9 pu.t2 3.2765
R6659 pu.n9 pu.n8 3.2765
R6660 pu.n5 pu.n2 3.013
R6661 pu.n10 pu.n7 3.013
R6662 pu.n2 pu.t4 1.8205
R6663 pu.n2 pu.n1 1.8205
R6664 pu.n7 pu.t6 1.8205
R6665 pu.n7 pu.n6 1.8205
R6666 pu.n10 pu.n5 0.445308
R6667 pu pu.n10 0.310308
R6668 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.t2 30.9379
R6669 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.t4 30.664
R6670 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.t5 24.5385
R6671 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.t3 24.5101
R6672 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n2 7.46763
R6673 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n3 5.28703
R6674 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n1 4.09208
R6675 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT 3.12156
R6676 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT 1.86016
R6677 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.OUT.n0 1.4252
R6678 IPD_.n0 IPD_.t4 16.5741
R6679 IPD_.n2 IPD_.t0 11.4186
R6680 IPD_.n1 IPD_.n0 10.5125
R6681 IPD_.n0 IPD_.t5 6.06211
R6682 IPD_.n1 IPD_.t2 6.06211
R6683 IPD_.n2 IPD_.n1 5.27348
R6684 IPD_.n5 IPD_.n2 4.21062
R6685 IPD_.n4 IPD_.t3 3.6405
R6686 IPD_.n4 IPD_.n3 3.6405
R6687 IPD_.n6 IPD_ 2.29359
R6688 IPD_.n6 IPD_.n5 1.93868
R6689 IPD_.n5 IPD_.n4 1.64004
R6690 IPD_ IPD_.n6 0.00720213
R6691 a_60634_18369.t6 a_60634_18369.n16 22.8782
R6692 a_60634_18369.n17 a_60634_18369.t6 22.4219
R6693 a_60634_18369.n14 a_60634_18369.t16 22.2916
R6694 a_60634_18369.n16 a_60634_18369.n15 14.0791
R6695 a_60634_18369.n15 a_60634_18369.n14 14.0791
R6696 a_60634_18369.n18 a_60634_18369.n17 14.0791
R6697 a_60634_18369.n12 a_60634_18369.t8 11.3416
R6698 a_60634_18369.n17 a_60634_18369.t10 8.34336
R6699 a_60634_18369.n18 a_60634_18369.t4 8.34336
R6700 a_60634_18369.n16 a_60634_18369.t17 8.213
R6701 a_60634_18369.n15 a_60634_18369.t15 8.213
R6702 a_60634_18369.n14 a_60634_18369.t14 8.213
R6703 a_60634_18369.n2 a_60634_18369.n13 4.0005
R6704 a_60634_18369.n1 a_60634_18369.n21 4.0005
R6705 a_60634_18369.n23 a_60634_18369.n1 3.63045
R6706 a_60634_18369.n0 a_60634_18369.n4 2.89398
R6707 a_60634_18369.n19 a_60634_18369.n18 2.60764
R6708 a_60634_18369.n9 a_60634_18369.n6 2.26392
R6709 a_60634_18369.n4 a_60634_18369.t5 1.8205
R6710 a_60634_18369.n4 a_60634_18369.n3 1.8205
R6711 a_60634_18369.t7 a_60634_18369.n23 1.8205
R6712 a_60634_18369.n23 a_60634_18369.n22 1.8205
R6713 a_60634_18369.n6 a_60634_18369.t2 1.6385
R6714 a_60634_18369.n6 a_60634_18369.n5 1.6385
R6715 a_60634_18369.n8 a_60634_18369.t3 1.6385
R6716 a_60634_18369.n8 a_60634_18369.n7 1.6385
R6717 a_60634_18369.n21 a_60634_18369.n19 1.56479
R6718 a_60634_18369.n13 a_60634_18369.n11 1.56479
R6719 a_60634_18369.n9 a_60634_18369.n8 1.4936
R6720 a_60634_18369.n2 a_60634_18369.n10 1.22554
R6721 a_60634_18369.n10 a_60634_18369.n9 1.18673
R6722 a_60634_18369.n1 a_60634_18369.n0 0.0789615
R6723 a_60634_18369.n0 a_60634_18369.n2 0.0720385
R6724 a_60634_18369.n21 a_60634_18369.n20 0.0656786
R6725 a_60634_18369.n13 a_60634_18369.n12 0.0656786
R6726 Vref.n0 Vref.t0 25.4398
R6727 Vref.n0 Vref.t1 17.6975
R6728 Vref Vref.n0 4.24656
C0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0951f
C1 VCO_mag_0.Delay_Cell_mag_0.OUTB a_65581_14091# 0.4f
C2 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 VDD 1.03f
C3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0013f
C4 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_69304_5529# 0.0202f
C5 a_69173_7501# VDD 2.21e-19
C6 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 3.14e-20
C7 a_63430_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C8 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00675f
C9 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 RST_DIV 0.138f
C10 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.79e-20
C11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_63270_5529# 0.00117f
C12 a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT VCO_mag_0.Delay_Cell_mag_1.IN 2.03e-21
C13 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.36e-19
C14 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.103f
C15 PFD_layout_0.VDIV VDD 1.74f
C16 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_66059_7499# 2.69e-19
C17 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD 0.651f
C18 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 4.36e-20
C19 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VCO_op 0.275f
C20 VDD IPD_ 1.06f
C21 IPD_ pd 9.43e-19
C22 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 a_72152_3335# 0.00138f
C23 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C24 PFD_layout_0.DFF__1.QB PFD_layout_0.nand2_0.IN1 0.618f
C25 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__1.inv_0.OUT 0.00685f
C26 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.00264f
C27 a_66213_6402# RST_DIV 0.00257f
C28 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00115f
C29 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C30 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VDD 5.47f
C31 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.0312f
C32 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_66287_5529# 1.04e-19
C33 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C34 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_67011_5529# 1.04e-19
C35 a_58943_16333# EN 0.0879f
C36 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C37 a_66783_7543# VCO_op 3.81e-19
C38 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 9.25e-19
C39 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 RST_DIV 0.00368f
C40 a_63270_5529# a_63430_5529# 0.0504f
C41 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.nand2_1.IN1 0.176f
C42 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_67735_5529# 0.00859f
C43 a_70188_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00696f
C44 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_64930_6448# 0.0157f
C45 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 1.5e-20
C46 a_66059_7499# a_66219_7499# 0.0504f
C47 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT RST_DIV 0.0915f
C48 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K RST_DIV 1.55e-19
C49 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD 0.916f
C50 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 2.11e-19
C51 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 VCO_op 0.0585f
C52 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.937f
C53 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 3.61e-20
C54 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 3.18e-19
C55 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_2.OUT 6.54e-20
C56 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD 1f
C57 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.57f
C58 a_67911_7543# VDD 3.56e-19
C59 VCO_mag_0.GF_INV16_2.IN VCO_mag_0.Delay_Cell_mag_2.OUT 3.48e-19
C60 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST_DIV 0.256f
C61 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.397f
C62 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_72487_4432# 2.06e-19
C63 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.0127f
C64 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0143f
C65 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT 0.026f
C66 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VCO_op 0.527f
C67 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C68 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT RST_DIV 5.45e-20
C69 PFD_layout_0.DFF__0.inv_0.OUT a_61538_21913# 0.00372f
C70 PFD_layout_0.VDIV VDD_VCO 0.0612f
C71 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 5.55e-19
C72 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C73 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.IN 0.0384f
C74 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 1.23e-19
C75 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.21e-20
C76 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C77 LF_mag_0.VCNTL PFD_layout_0.DFF__0.nand2_2.IN2 0.0599f
C78 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_63084_7501# 3.43e-19
C79 VCO_mag_0.GF_INV16_1.IN VCO_mag_0.GF_INV16_2.IN 0.0054f
C80 PFD_layout_0.DFF__1.QB a_62433_26095# 0.00619f
C81 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.GF_INV16_1.IN 5.46e-19
C82 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 2.34f
C83 VCO_mag_0.GF_INV1_1.OUT VCO_mag_0.Delay_Cell_mag_1.INB 0.00154f
C84 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C85 a_71248_9766# a_71408_9766# 0.186f
C86 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.GF_INV1_0.OUT 0.00842f
C87 a_66053_6402# RST_DIV 0.00257f
C88 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C89 a_69167_6404# VDD 2.76e-19
C90 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 9.87e-20
C91 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_60140_9217# 0.00572f
C92 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_73205_5529# 8.64e-19
C93 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 RST_DIV 0.0225f
C94 PFD_layout_0.DFF__1.nand2_1.IN1 PFD_layout_0.DFF__1.nand2_5.OUT 0.176f
C95 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C96 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_66213_6402# 0.00193f
C97 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 7.32e-20
C98 a_63430_5529# VCO_op 4.62e-19
C99 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0432f
C100 VCO_mag_0.Delay_Cell_mag_2.INB VCO_op 0.455f
C101 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.00442f
C102 a_66219_7499# VCO_op 0.0105f
C103 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.652f
C104 PFD_layout_0.DFF__0.nand2_5.OUT a_60305_23482# 3.83e-19
C105 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C106 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_70752_5529# 0.00378f
C107 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_64366_6448# 0.00859f
C108 a_70028_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00695f
C109 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.001f
C110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 0.132f
C111 a_66777_6402# a_66937_6402# 0.0504f
C112 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_0.INB 0.159f
C113 a_57637_42026# a_58117_42026# 0.0759f
C114 a_68299_5529# VDD 0.00152f
C115 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 2.03e-20
C116 a_64154_5529# VDD 0.00101f
C117 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_66783_7543# 0.00378f
C118 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.783f
C119 VCO_mag_0.Delay_Cell_mag_1.INB a_65581_17830# 0.487f
C120 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00262f
C121 VCO_mag_0.GF_INV16_2.IN a_65581_17830# 7.82e-20
C122 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.36f
C123 PFD_layout_0.DFF__1.nand2_2.IN1 Vref 3.73e-19
C124 a_67347_7543# VDD 3.14e-19
C125 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C126 a_73205_5529# RST_DIV 0.00146f
C127 a_58357_44128# VDD 0.248f
C128 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_72327_4432# 2.94e-19
C129 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 6.37e-19
C130 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.065f
C131 PFD_layout_0.DFF__1.CLK PFD_layout_0.DFF__0.nand2_5.OUT 6.57e-19
C132 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00367f
C133 VDD RST_DIV 2.81f
C134 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C135 PFD_layout_0.DFF__0.inv_0.OUT a_60302_21847# 1.29e-20
C136 LF_mag_0.VCNTL VCO_mag_0.Delay_Cell_mag_2.IN 0.0205f
C137 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.63e-19
C138 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2.18e-21
C139 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_62924_7501# 4.47e-19
C140 LF_mag_0.VCNTL PFD_layout_0.DFF__0.nand2_3.OUT 0.00837f
C141 PFD_layout_0.DFF__0.nand2_1.IN1 PFD_layout_0.DFF__0.nand2_2.IN2 0.459f
C142 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0622f
C143 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_63648_7545# 0.00378f
C144 VCO_mag_0.Delay_Cell_mag_1.INB a_59138_17829# 0.37f
C145 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 4.44e-20
C146 a_64930_6448# RST_DIV 0.00154f
C147 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 1.84e-19
C148 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 5.45e-20
C149 a_68065_6446# VDD 3.14e-19
C150 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_69470_4432# 9.32e-19
C151 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD 0.647f
C152 a_63270_5529# VCO_op 4.62e-19
C153 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_66053_6402# 0.00193f
C154 a_72487_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C155 PFD_layout_0.DFF__1.nand2_1.IN1 PFD_layout_0.nand2_0.IN1 0.0119f
C156 a_66059_7499# VCO_op 0.0114f
C157 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0582f
C158 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.48e-19
C159 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_63802_6404# 0.0101f
C160 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.654f
C161 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VCO_op 1.48e-19
C162 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_72492_7497# 1.19e-20
C163 a_67735_5529# VDD 0.00152f
C164 VCO_mag_0.Delay_Cell_mag_2.OUTB EN 0.43f
C165 a_61544_9654# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.132f
C166 a_63994_5529# VDD 0.00123f
C167 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00188f
C168 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_66219_7499# 0.0732f
C169 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 1.99f
C170 VCO_mag_0.Delay_Cell_mag_1.INB a_65386_20072# 0.566f
C171 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.36e-19
C172 a_66783_7543# VDD 3.14e-19
C173 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.CLK 0.0318f
C174 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0905f
C175 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.INB 3.11f
C176 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.28f
C177 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VCO_op 0.307f
C178 a_58117_42026# VDD 0.358f
C179 a_73045_5529# RST_DIV 0.00195f
C180 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.322f
C181 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_74380_2641# 3.02e-19
C182 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C183 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.294f
C184 a2x1mux_mag_0.Transmission_gate_mag_0.CLK IPD+ 0.00707f
C185 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00111f
C186 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_66937_6402# 2.88e-20
C187 a_58943_16333# VCO_op_bar 0.0232f
C188 a_60305_23482# PFD_layout_0.DFF__0.nand2_2.IN2 2.82e-20
C189 VCO_mag_0.Delay_Cell_mag_0.OUTB a_65386_16333# 0.455f
C190 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.65e-20
C191 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 VDD 4.24f
C192 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 9.8e-19
C193 PFD_layout_0.DFF__0.nand2_1.IN1 PFD_layout_0.DFF__0.nand2_3.OUT 0.39f
C194 a_60301_26043# PFD_layout_0.DFF__1.nand2_3.OUT 0.069f
C195 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_63084_7501# 0.0732f
C196 PFD_layout_0.DFF__0.inv_0.OUT VDD 0.346f
C197 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 1.17e-19
C198 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 1.59e-20
C199 a_61552_8823# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 3.01e-20
C200 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VCO_op 0.553f
C201 a_64366_6448# RST_DIV 0.00184f
C202 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD 1.17f
C203 PFD_layout_0.DFF__0.QB VCO_mag_0.Delay_Cell_mag_1.INB 0.0261f
C204 a_67501_6446# VDD 3.14e-19
C205 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 2.39e-20
C206 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_69310_4432# 0.00111f
C207 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.44e-20
C208 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN 0.389f
C209 PFD_layout_0.DFF__1.nand2_1.IN1 a_62433_26095# 1.63e-20
C210 a_64776_7545# VCO_op 9.34e-19
C211 a_72327_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C212 VCO_mag_0.Delay_Cell_mag_2.IN a_58943_16333# 0.0324f
C213 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C214 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0161f
C215 PFD_layout_0.DFF__0.CLK PFD_layout_0.VDIV 0.122f
C216 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C217 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VCO_op 1.96e-19
C218 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_61544_9654# 0.00718f
C219 a_66287_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.81e-19
C220 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_63642_6404# 0.0102f
C221 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0346f
C222 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 0.0409f
C223 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_72332_7497# 1.52e-20
C224 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 7.24e-20
C225 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN 1.2e-19
C226 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C227 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C228 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.316f
C229 a_70034_4432# RST_DIV 1.23e-20
C230 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_66059_7499# 0.0203f
C231 a_63430_5529# VDD 0.00892f
C232 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_74220_2641# 9.21e-20
C233 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_70216_3335# 2.36e-22
C234 a_72481_5529# RST_DIV 0.00247f
C235 a_58943_20071# VCO_mag_0.Delay_Cell_mag_1.INB 0.0406f
C236 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_70216_3335# 0.00929f
C237 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT a_69897_7545# 1.39e-19
C238 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.122f
C239 a_66213_6402# VCO_op 0.00164f
C240 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_73051_4432# 6.43e-21
C241 VDD IPD+ 0.0135f
C242 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_66777_6402# 9.1e-19
C243 IPD+ pd 0.493f
C244 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.2e-19
C245 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.98e-19
C246 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.06e-20
C247 VCO_mag_0.Delay_Cell_mag_2.OUT EN 0.3f
C248 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 1.76e-20
C249 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT RST_DIV 0.00539f
C250 a_71408_9766# VDD 0.0418f
C251 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.54e-20
C252 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.31f
C253 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 RST_DIV 0.00237f
C254 a_59584_26036# PFD_layout_0.DFF__1.nand2_3.OUT 1.26e-20
C255 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_62924_7501# 0.0203f
C256 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.32e-21
C257 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 1.47e-20
C258 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VCO_op 0.00637f
C259 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 3.4e-19
C260 PFD_layout_0.DFF__0.inv_0.OUT VDD_VCO 2.41e-19
C261 a_63802_6404# RST_DIV 0.00349f
C262 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT a_61552_8823# 1.78e-20
C263 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C264 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_68145_4432# 7.4e-19
C265 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_op 0.441f
C266 PFD_layout_0.nand2_0.IN1 PFD_layout_0.buffer_loading_mag_1.IN 0.28f
C267 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VCO_op 0.26f
C268 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.391f
C269 VCO_mag_0.GF_INV16_1.IN EN 0.183f
C270 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_0.IN 0.253f
C271 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C272 PFD_layout_0.buffer_mag_0.OUT a_60304_24408# 0.00519f
C273 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 0.00243f
C274 a_64212_7545# VCO_op 9.23e-19
C275 VCO_mag_0.GF_INV1_1.OUT EN 0.0419f
C276 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 7.1e-22
C277 a_72327_4432# a_72487_4432# 0.0504f
C278 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.93e-20
C279 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.93e-20
C280 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_63078_6404# 0.0152f
C281 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 7.89e-20
C282 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VCO_op 0.275f
C283 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_71025_7545# 0.0114f
C284 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0685f
C285 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 3.38e-19
C286 a_56677_42026# LF_mag_0.res_48k_mag_0.B 1.73e-19
C287 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0432f
C288 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_61552_8823# 0.0205f
C289 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C290 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0854f
C291 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0626f
C292 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_67806_9704# 0.0121f
C293 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD 0.648f
C294 a_67806_9704# VCO_op 0.00487f
C295 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.768f
C296 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0352f
C297 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN 1.61e-19
C298 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.54e-21
C299 a_62434_21795# VDD 3.15e-19
C300 a_63270_5529# VDD 0.0132f
C301 a_66059_7499# VDD 2.21e-19
C302 PFD_layout_0.DFF__1.nand2_2.IN2 a_61537_25977# 0.0769f
C303 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.nand2_2.IN1 0.492f
C304 a_72321_5529# RST_DIV 0.00247f
C305 VCO_mag_0.Delay_Cell_mag_2.INB VDD_VCO 3.18f
C306 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_70752_5529# 0.0036f
C307 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VDD 0.408f
C308 a_66053_6402# VCO_op 0.00117f
C309 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT a_69333_7501# 8.21e-19
C310 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_72481_5529# 0.0024f
C311 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.11f
C312 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_66213_6402# 0.0731f
C313 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__0.nand2_5.OUT 4.96e-19
C314 a_65581_17830# EN 0.202f
C315 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VCO_op 3.99e-20
C316 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 3.44e-20
C317 PFD_layout_0.DFF__1.nand2_3.OUT VDD 0.887f
C318 a_71248_9766# VDD 0.235f
C319 a_63436_4432# RST_DIV 7.81e-19
C320 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_71179_6448# 0.0811f
C321 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C322 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.17e-19
C323 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD 0.904f
C324 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 1.32e-19
C325 a_63642_6404# RST_DIV 0.00207f
C326 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C327 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT RST_DIV 0.28f
C328 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_67581_4432# 7.4e-19
C329 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 2.57e-19
C330 a_66777_6402# VDD 2.21e-19
C331 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 6.71e-19
C332 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_71184_3335# 1.29e-22
C333 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.INB 0.266f
C334 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_op_bar 0.0208f
C335 VCO_mag_0.Delay_Cell_mag_2.OUTB a_59138_14091# 0.4f
C336 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_66453_4432# 0.00939f
C337 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 1.83e-19
C338 a_59138_17829# EN 0.497f
C339 PFD_layout_0.buffer_mag_0.OUT a_59418_24365# 8.75e-20
C340 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.00178f
C341 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.1e-22
C342 PFD_layout_0.DFF__0.nand2_5.OUT a_62430_23292# 0.00454f
C343 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C344 a_63648_7545# VCO_op 3.8e-19
C345 a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT IPD+ 5.77e-19
C346 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0854f
C347 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_72327_4432# 8.64e-19
C348 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_62918_6404# 0.0124f
C349 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_70461_7545# 2.96e-19
C350 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 5.51e-20
C351 a_66053_6402# a_66213_6402# 0.0504f
C352 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD 3.83f
C353 VDD VCO_op 6.07f
C354 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C355 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.144f
C356 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C357 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.00174f
C358 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_0.IN 1.85e-19
C359 PFD_layout_0.DFF__1.nand2_1.IN1 Vref 1.13e-20
C360 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_67646_9704# 0.00747f
C361 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_69470_4432# 0.00119f
C362 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_70188_5529# 0.0101f
C363 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_70188_5529# 8.64e-19
C364 a_61538_21913# VDD 3.22e-19
C365 a_64776_7545# VDD 3.56e-19
C366 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_2.OUTB 0.269f
C367 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD 4.16f
C368 PFD_layout_0.DFF__0.nand2_5.OUT a_59419_23525# 0.00432f
C369 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.0266f
C370 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00109f
C371 a_57877_44128# VDD 0.248f
C372 a_61544_9654# VDD 0.165f
C373 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.nand2_2.IN1 0.0753f
C374 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT a_69173_7501# 0.00598f
C375 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_60147_7030# 0.069f
C376 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_72321_5529# 0.0024f
C377 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_66053_6402# 0.0202f
C378 PFD_layout_0.nand2_0.IN1 PFD_layout_0.buffer_mag_0.IN 0.44f
C379 a_65386_20072# EN 8.31e-20
C380 a_60301_26043# VDD 3.56e-19
C381 a_68511_9745# VDD 3.14e-19
C382 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00154f
C383 VCO_mag_0.Delay_Cell_mag_1.IN EN 0.267f
C384 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0275f
C385 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_70615_6448# 0.00964f
C386 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 0.0163f
C387 a_63276_4432# RST_DIV 9.37e-19
C388 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.198f
C389 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C390 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00586f
C391 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00776f
C392 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VCO_op 6.86e-20
C393 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0894f
C394 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00233f
C395 a_63078_6404# RST_DIV 9.47e-19
C396 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_63436_4432# 0.00939f
C397 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_67017_4432# 3.12e-19
C398 a_66213_6402# VDD 1.04e-19
C399 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 1.1e-19
C400 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_66293_4432# 0.0101f
C401 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.19e-19
C402 PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.DFF__0.nand2_2.IN2 0.0753f
C403 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 0.0683f
C404 a_63084_7501# VCO_op 0.0105f
C405 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_66453_4432# 0.00119f
C406 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 3.61e-21
C407 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD 0.397f
C408 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00917f
C409 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.04e-20
C410 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_69897_7545# 3.08e-19
C411 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 7.16e-20
C412 PFD_layout_0.DFF__1.QB PFD_layout_0.DFF__0.nand2_5.OUT 1.73e-20
C413 a_67611_25266# pu 1.66e-20
C414 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.02e-20
C415 VCO_mag_0.Delay_Cell_mag_2.OUT a_59138_14091# 0.487f
C416 VDD_VCO VCO_op 1.39f
C417 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_op_bar 0.0238f
C418 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_68511_9745# 3.04e-20
C419 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 7.55e-19
C420 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD 0.642f
C421 a_72327_4432# VDD 2.21e-19
C422 a_60140_9217# VCO_op 1.81e-19
C423 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_70028_5529# 0.0102f
C424 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 9.5e-19
C425 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VDD 0.496f
C426 a_73205_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C427 a_60302_21847# VDD 3.14e-19
C428 a_64212_7545# VDD 3.14e-19
C429 a_57637_42026# VDD 0.358f
C430 a2x1mux_mag_0.Transmission_gate_mag_0.CLK pd 0.033f
C431 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00397f
C432 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.994f
C433 a2x1mux_mag_0.Transmission_gate_mag_0.CLK VDD 0.483f
C434 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C435 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT 0.209f
C436 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.648f
C437 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT a_67911_7543# 8.11e-19
C438 a_67611_25266# VCO_mag_0.VCONT 0.219f
C439 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.59e-21
C440 PFD_layout_0.buffer_loading_mag_1.IN VCO_mag_0.Delay_Cell_mag_1.INB 0.00393f
C441 VCO_mag_0.GF_INV1_1.OUT VCO_op_bar 2.64e-19
C442 VCO_mag_0.GF_INV16_1.IN VCO_op_bar 0.46f
C443 PFD_layout_0.DFF__1.inv_0.OUT a_61537_25977# 0.00372f
C444 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.QB 0.581f
C445 a_58943_20071# EN 4.97e-19
C446 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.25f
C447 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_70051_6404# 0.00696f
C448 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_72152_3335# 0.0027f
C449 a_59584_26036# VDD 5.14e-19
C450 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN VDD 0.572f
C451 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_2.OUT 0.379f
C452 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C453 a_67646_9704# a_67806_9704# 0.0504f
C454 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_67171_5529# 2.88e-20
C455 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_71316_5529# 0.00372f
C456 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_63436_4432# 0.00119f
C457 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_63276_4432# 0.0101f
C458 a_62918_6404# RST_DIV 8.14e-19
C459 a_67618_24851# pu 2.15e-19
C460 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.442f
C461 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00165f
C462 a_66053_6402# VDD 2.21e-19
C463 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.395f
C464 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_65128_4432# 0.069f
C465 PFD_layout_0.buffer_mag_0.OUT a_61533_24598# 0.00168f
C466 a_59419_23525# PFD_layout_0.DFF__0.nand2_2.IN2 1.16e-20
C467 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-20
C468 a_62924_7501# VCO_op 0.0114f
C469 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.nand2_2.OUT 1.33e-19
C470 PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.DFF__0.nand2_3.OUT 0.0185f
C471 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 RST_DIV 2.96e-19
C472 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT a_69167_6404# 8.64e-19
C473 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.GF_INV16_1.IN 7.74e-23
C474 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_69464_5529# 3.66e-20
C475 a_72481_5529# VCO_op 1.84e-20
C476 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.QB 0.147f
C477 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_70034_4432# 1.25e-20
C478 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_69333_7501# 0.00392f
C479 a_57397_44128# a_57877_44128# 0.0759f
C480 a_72152_3335# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C481 VCO_mag_0.VCONT a_67618_24851# 0.151f
C482 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C483 CP_mag_0.inv_0.OUT pu 0.127f
C484 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_67806_9704# 8.5e-20
C485 VCO_mag_0.Delay_Cell_mag_0.OUT VDD_VCO 3.34f
C486 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_61106_7416# 1.14e-19
C487 a_71162_4432# VDD 3.56e-19
C488 a_59585_21854# VDD 3.14e-19
C489 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT 0.00935f
C490 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_69464_5529# 0.00789f
C491 a_63648_7545# VDD 3.14e-19
C492 a_73045_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C493 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.71e-20
C494 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 9e-20
C495 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.47e-20
C496 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT a_67347_7543# 3.47e-19
C497 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_72487_4432# 0.00119f
C498 CP_mag_0.inv_0.OUT VCO_mag_0.VCONT 0.283f
C499 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2f
C500 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00157f
C501 a_63016_9651# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.132f
C502 VDD pd 1.18f
C503 a_59138_17829# VCO_op_bar 0.0347f
C504 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0209f
C505 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C506 a_67646_9704# VDD 5.08e-19
C507 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 1.03e-19
C508 PFD_layout_0.DFF__0.nand2_5.OUT a_61534_23292# 0.0703f
C509 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT RST_DIV 0.0789f
C510 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_69891_6404# 0.00695f
C511 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.116f
C512 a_64154_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00696f
C513 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__1.inv_0.OUT 4.23e-20
C514 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.111f
C515 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_74179_4432# 0.069f
C516 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_67011_5529# 9.1e-19
C517 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_70752_5529# 0.069f
C518 PFD_layout_0.DFF__0.nand2_2.IN2 VCO_mag_0.Delay_Cell_mag_1.IN 2.01e-19
C519 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB RST_DIV 0.253f
C520 a_64930_6448# VDD 3.14e-19
C521 a_72152_3335# VDD 3.14e-19
C522 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 6.24e-20
C523 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_64564_4432# 6.06e-21
C524 a2x1mux_mag_0.Transmission_gate_mag_0.CLK a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT 0.247f
C525 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C526 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.88e-21
C527 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__0.inv_0.OUT 8.72e-22
C528 a_67911_7543# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C529 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C530 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 2.01e-19
C531 VCO_mag_0.Delay_Cell_mag_2.IN a_59138_17829# 0.404f
C532 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.92e-20
C533 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 RST_DIV 0.188f
C534 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.48e-19
C535 a_67611_25266# a_67618_24851# 0.279f
C536 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD 0.523f
C537 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C538 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 2.47e-19
C539 PFD_layout_0.DFF__0.QB PFD_layout_0.DFF__0.nand2_2.IN2 0.147f
C540 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT 0.127f
C541 a_65581_17830# a_65386_16333# 0.00414f
C542 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_67646_9704# 1.32e-19
C543 VCO_mag_0.Delay_Cell_mag_1.IN VCO_op_bar 0.496f
C544 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_mag_0.Delay_Cell_mag_0.INB 0.0121f
C545 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0385f
C546 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_69304_5529# 0.00335f
C547 a_70598_4432# VDD 3.14e-19
C548 PFD_layout_0.DFF__1.nand2_2.OUT PFD_layout_0.DFF__1.nand2_3.OUT 0.106f
C549 a_72481_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C550 a_73045_5529# a_73205_5529# 0.0504f
C551 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 9.94e-21
C552 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 4.88e-19
C553 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0384f
C554 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_67017_4432# 0.00378f
C555 a_73045_5529# VDD 2.21e-19
C556 a_63642_6404# VCO_op 6.8e-19
C557 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0836f
C558 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VCO_op 0.0854f
C559 PFD_layout_0.DFF__0.nand2_2.IN2 PFD_layout_0.DFF__0.nand2_2.OUT 0.159f
C560 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_74333_5529# 0.0157f
C561 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C562 PFD_layout_0.DFF__1.nand2_1.IN1 PFD_layout_0.DFF__0.nand2_5.OUT 1.69e-19
C563 CP_mag_0.inv_0.OUT a_67611_25266# 0.183f
C564 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0631f
C565 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.77e-20
C566 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C567 VDD VDD_VCO 0.217f
C568 a_63994_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00695f
C569 a_60140_9217# VDD 3.14e-19
C570 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_64718_5529# 0.00378f
C571 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.53e-20
C572 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_66447_5529# 0.0731f
C573 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_1.IN 0.0362f
C574 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C575 LF_mag_0.VCNTL VCO_mag_0.VCONT 4.11f
C576 PFD_layout_0.DFF__0.nand2_2.IN2 a_58943_20071# 0.0133f
C577 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.0262f
C578 PFD_layout_0.DFF__1.CLK a_60304_24408# 0.00347f
C579 a_65282_5529# RST_DIV 0.00138f
C580 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.35e-20
C581 a_64366_6448# VDD 3.14e-19
C582 a_63452_24694# PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN 0.002f
C583 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.103f
C584 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0707f
C585 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.307f
C586 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 0.00132f
C587 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 1.19f
C588 a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT VDD 1.33f
C589 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C590 a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT pd 1.55e-20
C591 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_69327_6404# 4.66e-19
C592 PFD_layout_0.VDIV Vref 3.36e-19
C593 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00213f
C594 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 RST_DIV 0.0298f
C595 CP_mag_0.inv_0.OUT a_67618_24851# 0.211f
C596 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_0.OUTB 0.214f
C597 a_57157_42026# a_57637_42026# 0.0759f
C598 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 3.7f
C599 PFD_layout_0.DFF__0.nand2_3.OUT PFD_layout_0.DFF__0.QB 0.0138f
C600 a_70034_4432# VDD 3.14e-19
C601 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_67347_7543# 4.52e-20
C602 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 7.07e-19
C603 a_72321_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C604 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.nand2_1.IN1 0.459f
C605 PFD_layout_0.DFF__1.nand2_2.OUT a_60301_26043# 0.00364f
C606 a_62924_7501# VDD 2.21e-19
C607 PFD_layout_0.DFF__1.QB PFD_layout_0.DFF__1.inv_0.OUT 0.00316f
C608 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 1.17e-19
C609 a_70615_6448# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.81e-20
C610 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00125f
C611 a_57397_44128# VDD 0.248f
C612 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT RST_DIV 0.286f
C613 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 2.46e-20
C614 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 3.98e-20
C615 a_72481_5529# VDD 0.00299f
C616 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_73769_5529# 0.00859f
C617 LF_mag_0.VCNTL PFD_layout_0.buffer_mag_0.OUT 0.00424f
C618 a_63078_6404# VCO_op 0.00253f
C619 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_68065_6446# 0.00372f
C620 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.23e-20
C621 PFD_layout_0.DFF__0.nand2_3.OUT PFD_layout_0.DFF__0.nand2_2.OUT 0.106f
C622 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_0.INB 0.256f
C623 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_67911_7543# 0.069f
C624 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_64212_7545# 4.52e-20
C625 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.109f
C626 VCO_mag_0.Delay_Cell_mag_2.IN a_58943_20071# 0.454f
C627 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0281f
C628 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.745f
C629 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_66287_5529# 0.0202f
C630 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.14f
C631 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C632 PFD_layout_0.DFF__0.nand2_3.OUT a_58943_20071# 2.71e-21
C633 a_64718_5529# RST_DIV 0.0015f
C634 PFD_layout_0.DFF__1.CLK a_59418_24365# 9.59e-19
C635 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C636 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.125f
C637 a_71184_3335# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C638 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.DFF__1.nand2_5.OUT 0.42f
C639 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.28f
C640 a_60307_8532# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 0.0732f
C641 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_69167_6404# 6.02e-19
C642 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.74e-19
C643 a_62924_7501# a_63084_7501# 0.0504f
C644 VCO_mag_0.VCONT a_58943_16333# 7.78e-19
C645 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 7.33e-20
C646 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.54e-20
C647 PFD_layout_0.DFF__0.nand2_3.OUT a_61534_23292# 0.00594f
C648 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_66783_7543# 0.0195f
C649 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN a_63591_22645# 8.3e-19
C650 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 RST_DIV 0.446f
C651 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 6.03e-20
C652 PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.nand2_5.OUT 0.0652f
C653 a_57157_42026# VDD 0.358f
C654 PFD_layout_0.DFF__1.nand2_2.OUT a_59584_26036# 0.069f
C655 a_72321_5529# VDD 0.00727f
C656 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_67501_6446# 0.069f
C657 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.nand2_1.IN1 0.487f
C658 a_62918_6404# VCO_op 0.00224f
C659 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C660 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.88e-19
C661 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 0.133f
C662 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT 0.00574f
C663 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C664 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 6.46e-20
C665 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_63648_7545# 0.0195f
C666 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 1.93e-20
C667 a_63436_4432# VDD 2.66e-19
C668 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 RST_DIV 0.166f
C669 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 5.49e-19
C670 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C671 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 6.36e-19
C672 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_67501_6446# 0.00378f
C673 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1e-19
C674 PFD_layout_0.DFF__0.CLK a_59585_21854# 1.27e-19
C675 a_63642_6404# VDD 2.21e-19
C676 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.994f
C677 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C678 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 4.69e-20
C679 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.nand2_0.IN1 2.23e-19
C680 a_60147_8532# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 0.0202f
C681 PFD_layout_0.DFF__0.CLK VDD 1f
C682 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_68065_6446# 0.0157f
C683 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 8.93e-19
C684 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.92f
C685 PFD_layout_0.DFF__1.nand2_2.OUT VDD 0.396f
C686 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT VCO_op 0.925f
C687 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 1.76f
C688 PFD_layout_0.buffer_loading_mag_1.IN a_65208_24138# 0.00403f
C689 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.299f
C690 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C691 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 4.31e-20
C692 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 RST_DIV 0.0697f
C693 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 2.51e-19
C694 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.0159f
C695 PFD_layout_0.buffer_mag_0.OUT a_60305_23482# 0.00519f
C696 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VCO_op 1.61e-19
C697 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C698 PFD_layout_0.DFF__1.inv_0.OUT PFD_layout_0.DFF__1.nand2_1.IN1 0.0551f
C699 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.306f
C700 a_72481_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C701 a_63276_4432# VDD 0.00752f
C702 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.00656f
C703 PFD_layout_0.VDIV EN 0.0787f
C704 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_66937_6402# 0.0733f
C705 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VCO_op 0.0844f
C706 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 6.91e-20
C707 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT a_68511_9745# 2.5e-19
C708 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_71184_3335# 1.45e-20
C709 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C710 a_63452_24694# pu 0.334f
C711 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.253f
C712 a_74179_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 1.54e-19
C713 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C714 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__1.CLK 0.0528f
C715 a_59584_26036# PFD_layout_0.DFF__1.nand2_5.OUT 1.99e-20
C716 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.19e-19
C717 PFD_layout_0.DFF__1.nand2_3.OUT a_62433_26095# 9.07e-21
C718 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.105f
C719 PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.nand2_2.IN2 0.117f
C720 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_64718_5529# 0.0036f
C721 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.2e-19
C722 a_60147_8532# a_60307_8532# 0.0504f
C723 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 2.49e-20
C724 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_67501_6446# 0.00859f
C725 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT a_72332_7497# 0.00472f
C726 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C727 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 6.91e-20
C728 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN 0.00134f
C729 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_64366_6448# 0.00378f
C730 IPD+ LP_ext 4.42e-20
C731 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 6.87e-20
C732 a_72321_5529# a_72481_5529# 0.0504f
C733 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_1.INB 0.00447f
C734 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_71408_9766# 1.9e-19
C735 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 1.89e-19
C736 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C737 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_74380_2641# 5.39e-20
C738 a2x1mux_mag_0.Transmission_gate_mag_0.CLK a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT 0.00208f
C739 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_2.OUTB 0.167f
C740 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT a_72326_6400# 8.64e-19
C741 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 1.82e-19
C742 VCO_mag_0.GF_INV1_0.OUT VCO_op 2.76e-19
C743 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_67347_7543# 0.0059f
C744 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_66219_7499# 2.79e-20
C745 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 RST_DIV 0.00434f
C746 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0838f
C747 VCO_mag_0.VCONT a2x1mux_mag_0.SEL 0.501f
C748 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2e-19
C749 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.105f
C750 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT 0.0128f
C751 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 RST_DIV 0.187f
C752 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT VCO_op 0.00322f
C753 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_66777_6402# 0.0203f
C754 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.24e-20
C755 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 4.85e-20
C756 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C757 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C758 a_62918_6404# VDD 2.21e-19
C759 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 1.65e-21
C760 PFD_layout_0.DFF__1.nand2_5.OUT VDD 0.802f
C761 a_63436_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C762 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VCO_op 0.00995f
C763 PFD_layout_0.DFF__1.nand2_2.IN1 a_59418_24365# 0.069f
C764 LF_mag_0.VCNTL PFD_layout_0.DFF__0.nand2_1.IN1 0.00437f
C765 PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.nand2_3.OUT 2.23e-19
C766 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 RST_DIV 0.301f
C767 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_64212_7545# 0.0059f
C768 PFD_layout_0.buffer_mag_0.IN a_65208_24138# 0.0691f
C769 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C770 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_70188_5529# 3.66e-20
C771 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.0116f
C772 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_66937_6402# 0.0101f
C773 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.92e-19
C774 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VCO_op 0.0834f
C775 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 8.56e-20
C776 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C777 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 0.0693f
C778 a_63642_6404# a_63802_6404# 0.0504f
C779 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_63802_6404# 0.0733f
C780 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C781 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C782 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 9.22e-20
C783 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C784 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.198f
C785 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 2.44e-20
C786 a_62434_21795# VCO_mag_0.Delay_Cell_mag_1.INB 2.94e-19
C787 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.342f
C788 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 3.69e-19
C789 a_56917_44128# VDD 0.248f
C790 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.038f
C791 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_74220_2641# 9.16e-20
C792 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_73056_7541# 0.00378f
C793 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD 0.396f
C794 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 3.61e-20
C795 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT a_71179_6448# 2.75e-21
C796 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_66783_7543# 0.0697f
C797 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0766f
C798 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT VDD 0.866f
C799 a_71316_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0811f
C800 a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT VDD 1.33f
C801 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.129f
C802 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 6.01e-19
C803 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_66213_6402# 1.5e-20
C804 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 4.69e-20
C805 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 1.82e-19
C806 a_67171_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0733f
C807 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 2.12e-19
C808 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 5.62e-19
C809 a_63276_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C810 PFD_layout_0.nand2_0.IN1 pd 0.00108f
C811 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_2.OUT 0.0362f
C812 PFD_layout_0.VDIV PFD_layout_0.DFF__0.nand2_2.IN2 0.00816f
C813 PFD_layout_0.nand2_0.IN1 VDD 1.99f
C814 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.5e-20
C815 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD 0.92f
C816 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_63648_7545# 0.0697f
C817 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C818 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K RST_DIV 3.04f
C819 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 4.75f
C820 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 VCO_op 0.748f
C821 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT RST_DIV 0.268f
C822 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_66777_6402# 0.0102f
C823 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00157f
C824 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.00774f
C825 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C826 VCO_mag_0.GF_INV16_2.IN VCO_op 0.282f
C827 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_63642_6404# 0.0203f
C828 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.651f
C829 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C830 VCO_mag_0.VCONT VCO_mag_0.GF_INV1_1.OUT 0.146f
C831 VCO_mag_0.Delay_Cell_mag_1.INB VCO_op 0.00408f
C832 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.129f
C833 VCO_mag_0.VCONT VCO_mag_0.GF_INV16_1.IN 0.0252f
C834 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_65282_5529# 0.00372f
C835 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 4.04e-19
C836 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00311f
C837 PFD_layout_0.VDIV a_59138_14091# 1.73e-19
C838 PFD_layout_0.VDIV VCO_op_bar 0.0161f
C839 a_56677_42026# VDD 0.368f
C840 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C841 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_72492_7497# 0.0732f
C842 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 0.888f
C843 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VCO_op 1.48f
C844 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_70051_6404# 2.88e-20
C845 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C846 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT a_70615_6448# 5.58e-22
C847 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0248f
C848 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_61544_9654# 0.00186f
C849 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_73615_4432# 0.0059f
C850 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 9.64e-20
C851 a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT VDD_VCO 4e-19
C852 a_70752_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00964f
C853 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.768f
C854 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_66053_6402# 1.17e-20
C855 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C856 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 RST_DIV 1.36e-19
C857 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 3.98e-20
C858 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0715f
C859 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_66219_7499# 1.24e-20
C860 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C861 PFD_layout_0.VDIV VCO_mag_0.Delay_Cell_mag_2.IN 6.82e-19
C862 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.nand2_2.IN1 0.0963f
C863 VCO_mag_0.VCONT a_65581_17830# 0.155f
C864 a_67011_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0203f
C865 a_65282_5529# VDD 0.00152f
C866 a_63276_4432# a_63436_4432# 0.0504f
C867 a_62433_26095# VDD 3.15e-19
C868 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_67911_7543# 0.00118f
C869 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 4.42e-19
C870 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0598f
C871 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0615f
C872 a_60305_23482# PFD_layout_0.DFF__0.nand2_1.IN1 0.069f
C873 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.buffer_mag_0.OUT 0.0963f
C874 a_71179_6448# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.81e-20
C875 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_66213_6402# 0.00789f
C876 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT VDD 0.434f
C877 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.0108f
C878 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C879 a_70188_5529# RST_DIV 0.00211f
C880 a2x1mux_mag_0.Transmission_gate_mag_0.CLK LP_ext 0.223f
C881 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_66937_6402# 8.64e-19
C882 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.52e-20
C883 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 6.22e-20
C884 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.002f
C885 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J 9.69e-19
C886 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VCO_op 0.519f
C887 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 1.01e-19
C888 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_63078_6404# 1.5e-20
C889 a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT 0.176f
C890 a_56917_44128# a_57397_44128# 0.0759f
C891 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 2.48e-19
C892 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.392f
C893 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 6.32e-22
C894 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_0.OUT 0.00336f
C895 VCO_mag_0.VCONT a_59138_17829# 0.035f
C896 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C897 VCO_mag_0.GF_INV16_2.IN VCO_mag_0.Delay_Cell_mag_0.OUT 1.68e-19
C898 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 6.18e-19
C899 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_64776_7545# 0.00118f
C900 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_64718_5529# 0.069f
C901 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C902 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.18e-19
C903 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C904 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_72332_7497# 0.0203f
C905 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN RST_DIV 4.25e-20
C906 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_68145_4432# 0.00372f
C907 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 1.74e-19
C908 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD 0.995f
C909 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 1.72e-19
C910 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_69891_6404# 9.1e-19
C911 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN 1.2e-19
C912 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C913 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_69470_4432# 0.00392f
C914 PFD_layout_0.DFF__1.QB a_62429_24598# 0.0692f
C915 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.inv_0.OUT 1.02e-21
C916 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_63016_9651# 0.015f
C917 VCO_mag_0.Delay_Cell_mag_2.INB EN 0.368f
C918 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_67171_5529# 8.64e-19
C919 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_73051_4432# 0.0697f
C920 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 4.39e-19
C921 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 9.75e-19
C922 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_66059_7499# 1.59e-20
C923 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 0.00252f
C924 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 0.117f
C925 PFD_layout_0.buffer_mag_0.OUT a_59419_23525# 8.75e-20
C926 PFD_layout_0.DFF__1.nand2_1.IN1 a_60304_24408# 0.069f
C927 a_64718_5529# VDD 0.00152f
C928 LF_mag_0.VCNTL a2x1mux_mag_0.SEL 0.295f
C929 VCO_mag_0.VCONT a_65386_20072# 0.00592f
C930 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_67347_7543# 0.011f
C931 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00388f
C932 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.03e-20
C933 a_67011_5529# a_67171_5529# 0.0504f
C934 a_66447_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.5e-20
C935 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_1.IN 0.359f
C936 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.329f
C937 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.103f
C938 VCO_mag_0.GF_INV1_0.OUT VDD_VCO 1.16f
C939 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C940 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.98e-19
C941 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 RST_DIV 0.0705f
C942 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C943 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C944 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.49e-19
C945 a_70028_5529# RST_DIV 0.00198f
C946 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_66053_6402# 0.00335f
C947 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.48e-19
C948 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00158f
C949 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00165f
C950 a_73051_4432# RST_DIV 2.78e-19
C951 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.159f
C952 VDD LP_ext 0.308f
C953 pd LP_ext 0.00207f
C954 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_62918_6404# 1.17e-20
C955 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_71248_9766# 8.09e-22
C956 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_64212_7545# 0.011f
C957 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_66453_4432# 0.00392f
C958 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 VDD 9.71f
C959 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.2e-20
C960 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 3.53e-19
C961 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VCO_op 0.0843f
C962 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__0.CLK 6.58e-19
C963 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_67581_4432# 0.069f
C964 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_69327_6404# 0.0731f
C965 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_63802_6404# 8.64e-19
C966 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C967 PFD_layout_0.DFF__1.nand2_2.OUT PFD_layout_0.DFF__1.nand2_5.OUT 1.33e-19
C968 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT RST_DIV 3.84e-20
C969 VCO_mag_0.Delay_Cell_mag_1.INB VDD 0.0069f
C970 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 2.52e-20
C971 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0485f
C972 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VCO_op 0.64f
C973 PFD_layout_0.DFF__1.QB PFD_layout_0.buffer_mag_0.OUT 1.19e-19
C974 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_loading_mag_1.IN 0.0224f
C975 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VCO_op 0.32f
C976 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD 2.82f
C977 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 0.00115f
C978 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C979 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 0.242f
C980 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C981 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_60307_8532# 1.75e-19
C982 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_64776_7545# 0.0114f
C983 a_66287_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.17e-20
C984 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_66783_7543# 1.43e-19
C985 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C986 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.107f
C987 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VCO_op 0.00323f
C988 VCO_mag_0.VCONT a_58943_20071# 7.89e-19
C989 a_61544_9654# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.69e-22
C990 LF_mag_0.VCNTL a_63591_22645# 0.00439f
C991 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.74e-19
C992 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 2.33e-19
C993 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_71184_3335# 0.0112f
C994 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_63436_4432# 0.00392f
C995 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_70216_3335# 0.0105f
C996 a_69464_5529# RST_DIV 0.00247f
C997 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.QB 9.68e-20
C998 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C999 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_67011_5529# 3.6e-22
C1000 a_62918_6404# a_63078_6404# 0.0504f
C1001 PFD_layout_0.DFF__0.inv_0.OUT PFD_layout_0.DFF__0.nand2_2.IN2 0.155f
C1002 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 3.38e-20
C1003 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.85e-19
C1004 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 1.83e-19
C1005 VDD Vref 0.217f
C1006 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_68511_9745# 2.05e-19
C1007 a_56677_42026# a_57157_42026# 0.0759f
C1008 VCO_mag_0.Delay_Cell_mag_2.OUTB a_58943_16333# 0.422f
C1009 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C1010 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_63648_7545# 1.43e-19
C1011 LF_mag_0.VCNTL PFD_layout_0.DFF__0.nand2_2.IN1 0.00414f
C1012 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 8.64e-20
C1013 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.101f
C1014 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_67501_6446# 0.0036f
C1015 a_69470_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0732f
C1016 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 RST_DIV 0.0555f
C1017 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 0.106f
C1018 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.nand2_2.OUT 0.0494f
C1019 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_69167_6404# 0.0202f
C1020 EN VCO_op 0.114f
C1021 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00156f
C1022 LF_mag_0.VCNTL VCO_mag_0.GF_INV1_1.OUT 0.00165f
C1023 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.15f
C1024 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C1025 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.DFF__0.nand2_5.OUT 1.35e-19
C1026 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 0.076f
C1027 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_0.OUTB 3.07e-20
C1028 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C1029 VCO_mag_0.GF_INV16_2.IN VDD_VCO 1.89f
C1030 VCO_mag_0.Delay_Cell_mag_1.INB VDD_VCO 4.09f
C1031 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 8.75e-20
C1032 a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT LP_ext 0.591f
C1033 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K VCO_op 8.07e-21
C1034 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.31e-19
C1035 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.71e-21
C1036 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_72487_4432# 0.00486f
C1037 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 7.36e-21
C1038 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VCO_op 3.15e-20
C1039 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C1040 PFD_layout_0.DFF__0.nand2_2.IN2 VCO_mag_0.Delay_Cell_mag_2.INB 0.00104f
C1041 a_65581_14091# VCO_op 0.0155f
C1042 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_60147_8532# 0.00369f
C1043 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_64212_7545# 2.96e-19
C1044 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_66219_7499# 0.00119f
C1045 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.96f
C1046 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0378f
C1047 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0871f
C1048 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_61552_8823# 0.00379f
C1049 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C1050 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C1051 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C1052 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2.62e-20
C1053 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C1054 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_66447_5529# 0.00166f
C1055 a_69304_5529# RST_DIV 0.00247f
C1056 PFD_layout_0.buffer_mag_0.OUT a_61534_23292# 0.00168f
C1057 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT RST_DIV 0.0914f
C1058 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0894f
C1059 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.458f
C1060 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 1.29e-19
C1061 PFD_layout_0.DFF__0.nand2_3.OUT PFD_layout_0.DFF__0.inv_0.OUT 0.142f
C1062 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 a_67911_7543# 0.00372f
C1063 VCO_mag_0.Delay_Cell_mag_2.INB VCO_op_bar 0.0736f
C1064 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_67806_9704# 0.0731f
C1065 VCO_mag_0.Delay_Cell_mag_2.INB a_59138_14091# 0.347f
C1066 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN 0.131f
C1067 PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.DFF__0.nand2_1.IN1 0.00714f
C1068 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_63084_7501# 0.00119f
C1069 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.nand2_3.OUT 0.0986f
C1070 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00101f
C1071 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.buffer_mag_0.IN 0.393f
C1072 a_69310_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0203f
C1073 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C1074 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.25e-19
C1075 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.13e-20
C1076 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VCO_op 0.00637f
C1077 VCO_mag_0.Delay_Cell_mag_0.OUT EN 0.0613f
C1078 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.57e-19
C1079 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 1.18e-19
C1080 VCO_mag_0.Delay_Cell_mag_2.OUT a_58943_16333# 1.31f
C1081 a_65581_17830# VCO_mag_0.Delay_Cell_mag_0.OUTB 0.584f
C1082 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 a_64776_7545# 0.00372f
C1083 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_67581_4432# 4.52e-20
C1084 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 9.45e-20
C1085 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.401f
C1086 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_71316_5529# 5.02e-20
C1087 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.37e-21
C1088 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.IN 3.03f
C1089 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_72327_4432# 0.00111f
C1090 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0156f
C1091 PFD_layout_0.DFF__0.nand2_2.IN2 a_62434_21795# 0.00411f
C1092 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C1093 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_64366_6448# 0.0036f
C1094 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.651f
C1095 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_63648_7545# 3.33e-19
C1096 PFD_layout_0.DFF__1.nand2_1.IN1 a_61533_24598# 0.00376f
C1097 VCO_mag_0.Delay_Cell_mag_0.OUT a_65581_14091# 0.487f
C1098 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.251f
C1099 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_71316_5529# 0.0157f
C1100 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_73051_4432# 0.00378f
C1101 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__1.nand2_1.IN1 0.487f
C1102 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD 1.32f
C1103 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_66287_5529# 0.001f
C1104 LF_mag_0.VCNTL a_65386_20072# 0.0112f
C1105 VCO_mag_0.Delay_Cell_mag_0.IN VCO_op 0.0227f
C1106 LF_mag_0.VCNTL VCO_mag_0.Delay_Cell_mag_1.IN 0.0719f
C1107 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 7.14e-19
C1108 a_66447_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.46e-19
C1109 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD 1.19f
C1110 PFD_layout_0.nand2_0.IN1 PFD_layout_0.DFF__1.nand2_5.OUT 0.0678f
C1111 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.424f
C1112 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 a_67347_7543# 0.069f
C1113 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT RST_DIV 0.346f
C1114 a_70216_3335# VDD 6e-19
C1115 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_67646_9704# 0.0202f
C1116 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00262f
C1117 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.103f
C1118 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_64930_6448# 0.0811f
C1119 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 9.73e-19
C1120 PFD_layout_0.DFF__1.nand2_2.IN2 a_60301_26043# 0.0144f
C1121 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 RST_DIV 1.38e-19
C1122 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 8.51e-22
C1123 a_69310_4432# a_69470_4432# 0.0504f
C1124 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C1125 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_64564_4432# 4.52e-20
C1126 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.54e-19
C1127 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C1128 LF_mag_0.VCNTL PFD_layout_0.DFF__0.QB 0.0129f
C1129 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 a_64212_7545# 0.069f
C1130 a_65128_4432# RST_DIV 6.14e-19
C1131 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 8.64e-20
C1132 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_67017_4432# 0.0202f
C1133 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_0.OUTB 0.04f
C1134 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 7.17e-19
C1135 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VCO_op 0.519f
C1136 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00125f
C1137 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.122f
C1138 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.25e-19
C1139 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0187f
C1140 PFD_layout_0.DFF__0.nand2_2.IN2 a_61538_21913# 0.0769f
C1141 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_71162_4432# 7.4e-19
C1142 PFD_layout_0.DFF__1.CLK PFD_layout_0.DFF__0.nand2_2.IN1 4.28e-19
C1143 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_63084_7501# 0.00392f
C1144 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_68145_4432# 9.26e-19
C1145 PFD_layout_0.buffer_loading_mag_1.IN pu 5.72e-19
C1146 VDD EN 0.00619f
C1147 PFD_layout_0.DFF__0.nand2_3.OUT a_62434_21795# 9.07e-21
C1148 LF_mag_0.VCNTL PFD_layout_0.DFF__0.nand2_2.OUT 0.00686f
C1149 a_66287_5529# a_66447_5529# 0.0504f
C1150 a_73205_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00696f
C1151 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_70752_5529# 0.00859f
C1152 a_59138_17829# a_58943_16333# 0.0277f
C1153 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 1.7e-20
C1154 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_70028_5529# 3.6e-22
C1155 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__1.CLK 0.146f
C1156 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K VDD 1.66f
C1157 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.DFF__0.nand2_3.OUT 5.53e-19
C1158 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_73615_4432# 4.52e-20
C1159 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.05e-19
C1160 VCO_op_bar VCO_op 0.0013f
C1161 a_59138_14091# VCO_op 0.0156f
C1162 LF_mag_0.VCNTL a_58943_20071# 0.0272f
C1163 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD 1f
C1164 a_74179_4432# VDD 3.56e-19
C1165 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 0.622f
C1166 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.IN 0.314f
C1167 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C1168 PFD_layout_0.DFF__0.nand2_5.OUT a_59585_21854# 1.99e-20
C1169 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 2.08e-20
C1170 a_61552_8823# VDD 3.85e-19
C1171 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_64366_6448# 0.00964f
C1172 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 2.01e-19
C1173 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.0212f
C1174 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 0.00243f
C1175 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_64000_4432# 0.0202f
C1176 PFD_layout_0.DFF__1.nand2_2.IN2 a_59584_26036# 0.0175f
C1177 PFD_layout_0.DFF__0.nand2_5.OUT VDD 0.803f
C1178 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_67581_4432# 0.0059f
C1179 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_66213_6402# 1.46e-19
C1180 a_74220_2641# a_74380_2641# 0.186f
C1181 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C1182 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_60147_7030# 0.00347f
C1183 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0129f
C1184 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 2.85e-20
C1185 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C1186 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 2.03e-20
C1187 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_69333_7501# 1.16e-20
C1188 a_64564_4432# RST_DIV 6.14e-19
C1189 VCO_mag_0.Delay_Cell_mag_2.IN VCO_op 0.00281f
C1190 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.DFF__1.inv_0.OUT 0.142f
C1191 VCO_mag_0.Delay_Cell_mag_1.IN a_58943_16333# 0.0923f
C1192 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT RST_DIV 0.0792f
C1193 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 2.29e-19
C1194 PFD_layout_0.DFF__0.nand2_1.IN1 PFD_layout_0.DFF__0.QB 0.273f
C1195 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 RST_DIV 0.0189f
C1196 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_70598_4432# 7.4e-19
C1197 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_69470_4432# 2.79e-20
C1198 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C1199 PFD_layout_0.DFF__1.CLK a_59419_23525# 1.82e-19
C1200 PFD_layout_0.DFF__0.nand2_2.IN2 a_60302_21847# 0.0144f
C1201 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.397f
C1202 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 0.124f
C1203 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_70598_4432# 4.52e-20
C1204 PFD_layout_0.DFF__0.nand2_3.OUT a_61538_21913# 2.09e-19
C1205 a_63591_22645# a2x1mux_mag_0.SEL 9.45e-19
C1206 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C1207 a_61106_7416# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C1208 VDD_VCO EN 1.18f
C1209 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.buffer_loading_mag_1.IN 0.0112f
C1210 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_73769_5529# 0.00378f
C1211 a_73045_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00695f
C1212 a_71025_7545# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C1213 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_73774_6444# 0.00378f
C1214 VCO_mag_0.Delay_Cell_mag_2.OUT VCO_mag_0.Delay_Cell_mag_2.OUTB 2.47f
C1215 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_68145_4432# 0.00118f
C1216 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_69464_5529# 0.00166f
C1217 a_74333_5529# VDD 3.14e-19
C1218 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VCO_op 7.51e-20
C1219 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C1220 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.96e-20
C1221 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_73051_4432# 0.0202f
C1222 a_65386_16333# VCO_op 0.0268f
C1223 a_70188_5529# VDD 0.00101f
C1224 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_64564_4432# 0.0059f
C1225 a_73615_4432# VDD 3.14e-19
C1226 a_65581_14091# VDD_VCO 0.0541f
C1227 a_69891_6404# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.49e-20
C1228 a_65282_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0811f
C1229 VCO_mag_0.GF_INV16_1.IN VCO_mag_0.Delay_Cell_mag_2.OUTB 0.00108f
C1230 a_62433_26095# PFD_layout_0.nand2_0.IN1 0.069f
C1231 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 7.47e-19
C1232 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C1233 PFD_layout_0.DFF__1.nand2_2.IN2 VDD 0.837f
C1234 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VCO_op 5.56e-19
C1235 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_63802_6404# 0.00696f
C1236 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.00115f
C1237 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_73620_7541# 4.52e-20
C1238 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 4.67e-22
C1239 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 8.33e-20
C1240 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VCO_op 5.73e-19
C1241 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_67017_4432# 0.0697f
C1242 a_65208_24138# VDD 3.26e-19
C1243 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_71179_6448# 0.00372f
C1244 a_65208_24138# pd 6.49e-19
C1245 PFD_layout_0.buffer_mag_0.IN pu 5.63e-19
C1246 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_66453_4432# 2.79e-20
C1247 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN VDD 0.582f
C1248 a_64000_4432# RST_DIV 2.66e-19
C1249 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_69173_7501# 1.49e-20
C1250 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C1251 PFD_layout_0.DFF__0.nand2_1.IN1 a_61534_23292# 0.00376f
C1252 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.72e-19
C1253 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.124f
C1254 a_60301_26043# PFD_layout_0.DFF__1.inv_0.OUT 1.29e-20
C1255 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C1256 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_65128_4432# 0.00118f
C1257 a_60302_21847# VCO_mag_0.Delay_Cell_mag_2.IN 1.82e-20
C1258 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C1259 a_69304_5529# VCO_op 3.76e-20
C1260 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 2.59e-19
C1261 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_70034_4432# 3.12e-19
C1262 a_72152_3335# CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 2.94e-20
C1263 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C1264 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VCO_op 0.26f
C1265 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_63078_6404# 8.66e-20
C1266 PFD_layout_0.DFF__0.nand2_2.IN2 a_59585_21854# 0.0175f
C1267 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 2.48e-19
C1268 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_68511_9745# 0.069f
C1269 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_67017_4432# 6.43e-21
C1270 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_70034_4432# 0.0202f
C1271 PFD_layout_0.DFF__0.nand2_3.OUT a_60302_21847# 0.069f
C1272 pu IPD_ 0.0891f
C1273 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_73210_6400# 0.0733f
C1274 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_67581_4432# 0.011f
C1275 PFD_layout_0.DFF__0.nand2_2.IN2 VDD 0.71f
C1276 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.76e-20
C1277 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_69304_5529# 0.00119f
C1278 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.146f
C1279 a_73769_5529# VDD 3.14e-19
C1280 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 1.83e-20
C1281 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 6.03e-19
C1282 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 9.05e-22
C1283 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.18f
C1284 a_70028_5529# VDD 0.00123f
C1285 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_64000_4432# 0.0697f
C1286 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 1.41e-20
C1287 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 1.84e-21
C1288 VCO_mag_0.Delay_Cell_mag_0.OUT a_65386_16333# 0.699f
C1289 VCO_mag_0.VCONT IPD_ 0.00567f
C1290 a_73051_4432# VDD 3.14e-19
C1291 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.283f
C1292 a_59138_17829# VCO_mag_0.Delay_Cell_mag_2.OUTB 5.63e-19
C1293 a_64718_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00964f
C1294 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 6.91e-20
C1295 a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT LP_ext 0.0331f
C1296 a_72486_6400# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 7.56e-21
C1297 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT 0.203f
C1298 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_63642_6404# 0.00695f
C1299 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C1300 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_73056_7541# 0.0195f
C1301 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_74179_4432# 0.00118f
C1302 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_70615_6448# 0.069f
C1303 PFD_layout_0.DFF__1.nand2_1.IN1 PFD_layout_0.DFF__0.nand2_1.IN1 8.9e-19
C1304 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 6.93e-19
C1305 VCO_mag_0.Delay_Cell_mag_0.IN VDD_VCO 0.513f
C1306 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 0.161f
C1307 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.buffer_mag_0.IN 0.00294f
C1308 VCO_mag_0.GF_INV16_1.IN VCO_mag_0.Delay_Cell_mag_2.OUT 0.00213f
C1309 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT RST_DIV 0.0157f
C1310 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_67911_7543# 0.0114f
C1311 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD 0.649f
C1312 PFD_layout_0.DFF__1.QB a_63452_24694# 0.00174f
C1313 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_64000_4432# 6.43e-21
C1314 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_64564_4432# 0.011f
C1315 PFD_layout_0.DFF__0.nand2_3.OUT a_59585_21854# 1.26e-20
C1316 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_67806_9704# 4.43e-21
C1317 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__0.nand2_2.IN1 0.00935f
C1318 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C1319 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 1.34e-19
C1320 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.84e-20
C1321 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN 1.48e-19
C1322 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_73050_6400# 0.0203f
C1323 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 9.88e-20
C1324 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 2.42f
C1325 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT VCO_op 0.578f
C1326 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 0.291f
C1327 a_66937_6402# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 1.04e-19
C1328 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_2.OUTB 0.00793f
C1329 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_67017_4432# 1.43e-19
C1330 VCO_mag_0.GF_INV1_1.OUT VCO_mag_0.GF_INV16_1.IN 0.219f
C1331 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 6.57e-19
C1332 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C1333 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 6.35e-19
C1334 a2x1mux_mag_0.SEL a_65386_20072# 2.86e-19
C1335 PFD_layout_0.DFF__0.nand2_3.OUT VDD 0.886f
C1336 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VCO_op 0.00639f
C1337 PFD_layout_0.DFF__0.nand2_2.IN2 VDD_VCO 0.023f
C1338 a2x1mux_mag_0.SEL VCO_mag_0.Delay_Cell_mag_1.IN 5.56e-19
C1339 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00545f
C1340 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C1341 LF_mag_0.VCNTL LF_mag_0.res_48k_mag_0.B 0.436f
C1342 a_69464_5529# VDD 0.00891f
C1343 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_71162_4432# 0.00118f
C1344 a_67611_25266# IPD_ 0.111f
C1345 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT 0.139f
C1346 LF_mag_0.VCNTL PFD_layout_0.buffer_loading_mag_1.IN 0.00905f
C1347 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J 0.133f
C1348 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_73615_4432# 0.011f
C1349 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 1.12e-19
C1350 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 1.37e-20
C1351 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C1352 VCO_mag_0.Delay_Cell_mag_0.INB VCO_op 0.55f
C1353 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.08f
C1354 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C1355 VDD_VCO VCO_op_bar 1.29f
C1356 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.149f
C1357 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.0758f
C1358 PFD_layout_0.DFF__1.inv_0.OUT VDD 0.347f
C1359 a_59138_14091# VDD_VCO 0.054f
C1360 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.29e-19
C1361 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_67347_7543# 2.96e-19
C1362 a_59138_17829# VCO_mag_0.Delay_Cell_mag_2.OUT 0.00237f
C1363 a_59419_23525# PFD_layout_0.DFF__0.nand2_2.IN1 0.069f
C1364 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00808f
C1365 a_66453_4432# VDD 2.66e-19
C1366 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.434f
C1367 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 0.00718f
C1368 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_64000_4432# 1.43e-19
C1369 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD 0.424f
C1370 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 2.18e-21
C1371 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1.74e-19
C1372 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB RST_DIV 0.295f
C1373 a_67618_24851# IPD_ 0.00945f
C1374 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 7.16e-20
C1375 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_67646_9704# 3.44e-21
C1376 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.777f
C1377 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.83e-19
C1378 PFD_layout_0.DFF__1.nand2_1.IN1 PFD_layout_0.DFF__1.CLK 0.114f
C1379 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT RST_DIV 0.0784f
C1380 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_72486_6400# 1.5e-20
C1381 VCO_mag_0.Delay_Cell_mag_2.IN VDD_VCO 4.54f
C1382 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.GF_INV1_0.OUT 0.156f
C1383 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.CLK 0.115f
C1384 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.012f
C1385 VCO_mag_0.GF_INV1_0.OUT VCO_mag_0.GF_INV16_2.IN 0.228f
C1386 a_59138_17829# VCO_mag_0.GF_INV16_1.IN 4.81e-20
C1387 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_68065_6446# 0.0811f
C1388 PFD_layout_0.DFF__0.nand2_3.OUT VDD_VCO 2.74e-19
C1389 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 3.6e-21
C1390 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 0.00154f
C1391 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_70598_4432# 0.011f
C1392 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1393 CP_mag_0.inv_0.OUT IPD_ 0.27f
C1394 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1395 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_69897_7545# 0.00378f
C1396 a_69304_5529# VDD 0.0132f
C1397 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD 0.642f
C1398 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C1399 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_68145_4432# 4.52e-20
C1400 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_73769_5529# 0.0036f
C1401 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 8.26e-20
C1402 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_2.OUT 0.00529f
C1403 a_73050_6400# a_73210_6400# 0.0504f
C1404 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 7.11e-19
C1405 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 1.05e-20
C1406 PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.nand2_1.IN1 0.0119f
C1407 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT 0.0599f
C1408 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VCO_op 3.39e-20
C1409 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_73051_4432# 1.43e-19
C1410 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 1.89e-19
C1411 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C1412 a_67806_9704# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 4.33e-21
C1413 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C1414 VCO_mag_0.Delay_Cell_mag_0.OUT VCO_mag_0.Delay_Cell_mag_0.INB 0.00336f
C1415 a_65386_16333# VDD_VCO 1.13f
C1416 a_71184_3335# CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.00138f
C1417 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_74380_2641# 0.019f
C1418 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_66783_7543# 3.12e-19
C1419 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.GF_INV1_1.OUT 0.348f
C1420 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.GF_INV16_1.IN 0.252f
C1421 a_66293_4432# VDD 3.78e-19
C1422 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_73620_7541# 0.00605f
C1423 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0345f
C1424 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 1.39e-19
C1425 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00119f
C1426 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00254f
C1427 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_72326_6400# 1.17e-20
C1428 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_72486_6400# 4.28e-19
C1429 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 2.76e-19
C1430 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 5.48e-20
C1431 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 2.59e-19
C1432 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.nand2_2.OUT 0.159f
C1433 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C1434 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_65128_4432# 4.52e-20
C1435 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C1436 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_60307_8532# 6.63e-20
C1437 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_67501_6446# 0.00964f
C1438 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 2.27e-20
C1439 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J RST_DIV 0.00458f
C1440 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_69333_7501# 0.0732f
C1441 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 1.93f
C1442 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_70034_4432# 1.43e-19
C1443 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_73210_6400# 8.64e-19
C1444 PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.DFF__0.nand2_2.OUT 0.451f
C1445 LF_mag_0.VCNTL PFD_layout_0.VDIV 0.108f
C1446 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 1.32e-19
C1447 VCO_mag_0.Delay_Cell_mag_1.IN a_65581_17830# 0.4f
C1448 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT VDD 0.829f
C1449 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 4e-19
C1450 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 1.33e-20
C1451 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00253f
C1452 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.397f
C1453 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0934f
C1454 PFD_layout_0.DFF__0.CLK PFD_layout_0.DFF__0.nand2_2.IN2 0.0318f
C1455 PFD_layout_0.DFF__0.QB a_62430_23292# 0.0692f
C1456 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 RST_DIV 9.24e-20
C1457 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.199f
C1458 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN 3.11e-19
C1459 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_66219_7499# 0.00392f
C1460 a_65128_4432# VDD 3.56e-19
C1461 VCO_mag_0.Delay_Cell_mag_1.IN a_59138_17829# 0.337f
C1462 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 3.27e-20
C1463 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.GF_INV16_2.IN 3.07e-19
C1464 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.109f
C1465 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0379f
C1466 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.119f
C1467 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_73056_7541# 0.0697f
C1468 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_74179_4432# 4.52e-20
C1469 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C1470 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__0.nand2_5.OUT 1.45f
C1471 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 4.8e-20
C1472 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C1473 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 9.58e-19
C1474 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 3.09e-19
C1475 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.342f
C1476 pu IPD+ 0.0687f
C1477 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_2.INB 0.0215f
C1478 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_74179_4432# 0.00372f
C1479 PFD_layout_0.DFF__1.nand2_1.IN1 a_61537_25977# 0.00384f
C1480 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_72326_6400# 5.5e-19
C1481 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.inv_0.OUT 0.00685f
C1482 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_60147_8532# 4.15e-19
C1483 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 3.39e-20
C1484 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_66937_6402# 0.00696f
C1485 VCO_mag_0.VCONT IPD+ 3.29e-19
C1486 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.88e-20
C1487 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_69173_7501# 0.0203f
C1488 a_74179_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 2.1e-20
C1489 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J 5.85e-19
C1490 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00123f
C1491 PFD_layout_0.DFF__0.nand2_1.IN1 PFD_layout_0.VDIV 4.13e-21
C1492 VCO_mag_0.Delay_Cell_mag_1.IN a_65386_20072# 0.454f
C1493 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VCO_op 0.267f
C1494 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C1495 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0306f
C1496 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.59e-21
C1497 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.14e-19
C1498 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 9.83e-19
C1499 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_73210_6400# 2.88e-20
C1500 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.25f
C1501 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_71162_4432# 4.52e-20
C1502 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_71025_7545# 0.069f
C1503 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_74333_5529# 0.00372f
C1504 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.nand2_5.OUT 0.0065f
C1505 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00136f
C1506 a_64564_4432# VDD 3.14e-19
C1507 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD 0.748f
C1508 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C1509 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C1510 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 1.36e-20
C1511 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00952f
C1512 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN VDD 1f
C1513 PFD_layout_0.DFF__0.QB VCO_mag_0.Delay_Cell_mag_1.IN 1.13e-19
C1514 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN pd 0.00115f
C1515 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.395f
C1516 VCO_mag_0.Delay_Cell_mag_0.INB VDD_VCO 0.795f
C1517 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_73615_4432# 0.069f
C1518 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.01e-19
C1519 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__1.nand2_1.IN1 0.00714f
C1520 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_71179_6448# 0.0157f
C1521 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_74184_7541# 0.00118f
C1522 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_66777_6402# 0.00695f
C1523 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 RST_DIV 0.03f
C1524 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C1525 a_67611_25266# IPD+ 3.09e-19
C1526 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 4.07e-19
C1527 VCO_mag_0.GF_INV1_0.OUT EN 0.0349f
C1528 a_72332_7497# a_72492_7497# 0.0504f
C1529 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0346f
C1530 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_73050_6400# 9.1e-19
C1531 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00121f
C1532 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VCO_op 0.484f
C1533 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C1534 a_67171_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00696f
C1535 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 8.64e-20
C1536 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_73774_6444# 0.0036f
C1537 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 3.97e-19
C1538 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 4.26e-19
C1539 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_73769_5529# 0.069f
C1540 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VCO_op 8.88e-20
C1541 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 7.34e-20
C1542 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.nand2_0.IN1 0.117f
C1543 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 6.51e-19
C1544 a_64000_4432# VDD 3.14e-19
C1545 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB RST_DIV 0.182f
C1546 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.026f
C1547 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.22e-20
C1548 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT RST_DIV 0.268f
C1549 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.349f
C1550 a_67618_24851# IPD+ 0.0463f
C1551 a_60304_24408# VDD 4.86e-19
C1552 PFD_layout_0.nand2_0.IN1 a_65208_24138# 0.00348f
C1553 VCO_mag_0.VCONT VCO_op 0.086f
C1554 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C1555 PFD_layout_0.DFF__1.nand2_3.OUT a_61533_24598# 0.00594f
C1556 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.211f
C1557 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT a_60147_7030# 4.44e-20
C1558 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 1.85e-19
C1559 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.61e-21
C1560 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 4.78e-20
C1561 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__1.nand2_3.OUT 0.889f
C1562 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_70615_6448# 0.00859f
C1563 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_73620_7541# 0.011f
C1564 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00391f
C1565 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00126f
C1566 PFD_layout_0.DFF__0.nand2_2.OUT a_58943_20071# 6.28e-20
C1567 CP_mag_0.inv_0.OUT IPD+ 0.127f
C1568 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C1569 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.77e-19
C1570 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0072f
C1571 PFD_layout_0.buffer_loading_mag_1.IN a_63591_22645# 0.453f
C1572 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0106f
C1573 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VCO_op 5.45e-20
C1574 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 1.12e-19
C1575 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0661f
C1576 a_72326_6400# a_72486_6400# 0.0504f
C1577 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00156f
C1578 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0378f
C1579 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT RST_DIV 5.36e-20
C1580 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__0.nand2_3.OUT 1.36e-19
C1581 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_72486_6400# 0.0731f
C1582 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C1583 a_63452_24694# PFD_layout_0.buffer_mag_0.IN 0.0158f
C1584 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 1.89e-20
C1585 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN a_63016_9651# 2.4e-20
C1586 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.0549f
C1587 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C1588 a_67011_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00695f
C1589 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_67735_5529# 0.00378f
C1590 LF_mag_0.VCNTL PFD_layout_0.DFF__0.inv_0.OUT 0.00546f
C1591 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 5.2e-20
C1592 PFD_layout_0.DFF__1.QB PFD_layout_0.DFF__1.nand2_1.IN1 0.273f
C1593 PFD_layout_0.DFF__1.nand2_2.IN2 a_62433_26095# 0.00411f
C1594 a_71316_5529# RST_DIV 0.00122f
C1595 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.348f
C1596 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD 0.647f
C1597 a2x1mux_mag_0.Transmission_gate_mag_0.CLK pu 1.27e-20
C1598 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.113f
C1599 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C1600 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0497f
C1601 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.342f
C1602 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN 0.00296f
C1603 a_67171_5529# RST_DIV 0.00211f
C1604 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_60147_7030# 0.0111f
C1605 a_59418_24365# VDD 0.00503f
C1606 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C1607 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_0.OUT 0.222f
C1608 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 a_74380_2641# 0.00894f
C1609 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J VCO_op 0.779f
C1610 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.71e-21
C1611 VCO_mag_0.Delay_Cell_mag_1.INB EN 0.209f
C1612 PFD_layout_0.DFF__1.inv_0.OUT PFD_layout_0.DFF__1.nand2_5.OUT 1.02e-21
C1613 VCO_mag_0.GF_INV16_2.IN EN 0.178f
C1614 a_63452_24694# IPD_ 1.01e-19
C1615 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 2.48e-19
C1616 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 3.54e-20
C1617 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.31e-20
C1618 PFD_layout_0.buffer_mag_0.OUT a_60301_26043# 0.00348f
C1619 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_70051_6404# 0.0101f
C1620 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.289f
C1621 PFD_layout_0.VDIV a_74380_2641# 0.198f
C1622 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C1623 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.25e-20
C1624 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.CLK 0.499f
C1625 PFD_layout_0.VDIV VCO_mag_0.Delay_Cell_mag_2.OUTB 3.01e-19
C1626 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_73056_7541# 1.43e-19
C1627 LF_mag_0.VCNTL VCO_mag_0.Delay_Cell_mag_2.INB 0.022f
C1628 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.209f
C1629 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_69470_4432# 1.41e-20
C1630 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_63016_9651# 0.00589f
C1631 PFD_layout_0.buffer_loading_mag_1.IN a_62430_23292# 0.00347f
C1632 a_63016_9651# VCO_op 1.64e-20
C1633 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 6.12e-21
C1634 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_72326_6400# 0.0202f
C1635 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C1636 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.38e-19
C1637 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C1638 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT RST_DIV 0.0596f
C1639 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 2.17e-21
C1640 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 0.305f
C1641 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN VCO_op 7e-19
C1642 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT RST_DIV 3.84e-20
C1643 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_69333_7501# 2.79e-20
C1644 PFD_layout_0.DFF__0.nand2_1.IN1 PFD_layout_0.DFF__0.inv_0.OUT 0.0551f
C1645 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 1.51e-19
C1646 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 RST_DIV 0.178f
C1647 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 4.22e-20
C1648 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0899f
C1649 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 6.23e-19
C1650 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C1651 PFD_layout_0.buffer_mag_0.OUT a_60302_21847# 0.00348f
C1652 a_70752_5529# RST_DIV 0.00119f
C1653 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT a_61106_7416# 0.0177f
C1654 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 a_74220_2641# 0.0294f
C1655 a_67011_5529# RST_DIV 0.00195f
C1656 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C1657 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_64000_4432# 0.00378f
C1658 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD 0.904f
C1659 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_64154_5529# 0.0101f
C1660 a_62429_24598# VDD 3.15e-19
C1661 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.28f
C1662 pu pd 0.0986f
C1663 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 0.00118f
C1664 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C1665 a_70216_3335# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C1666 VDD pu 0.921f
C1667 PFD_layout_0.buffer_mag_0.IN a_63591_22645# 0.0088f
C1668 PFD_layout_0.DFF__1.inv_0.OUT PFD_layout_0.nand2_0.IN1 5.29e-19
C1669 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD 0.768f
C1670 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_66453_4432# 1.41e-20
C1671 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 RST_DIV 0.237f
C1672 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_69891_6404# 0.0102f
C1673 a_67611_25266# a2x1mux_mag_0.Transmission_gate_mag_0.CLK 1.21e-19
C1674 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C1675 PFD_layout_0.VDIV a_74220_2641# 0.0133f
C1676 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN 0.0121f
C1677 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_72492_7497# 0.00119f
C1678 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 6.62e-20
C1679 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT 0.00103f
C1680 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD 0.517f
C1681 VCO_mag_0.VCONT pd 0.0409f
C1682 LF_mag_0.VCNTL a_62434_21795# 9.16e-19
C1683 VCO_mag_0.VCONT VDD 2.89f
C1684 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_69310_4432# 1.86e-20
C1685 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.299f
C1686 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 a_74184_7541# 0.00372f
C1687 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.105f
C1688 PFD_layout_0.VDIV VCO_mag_0.Delay_Cell_mag_2.OUT 2.74e-19
C1689 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 0.104f
C1690 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C1691 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.24f
C1692 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_60307_8532# 0.0177f
C1693 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C1694 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.125f
C1695 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C1696 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_72486_6400# 1.46e-19
C1697 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 8.24e-19
C1698 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.179f
C1699 PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.VDIV 2.43e-19
C1700 VCO_mag_0.Delay_Cell_mag_2.INB a_58943_16333# 7.46e-19
C1701 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.0145f
C1702 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VDD 0.41f
C1703 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_71184_3335# 0.0084f
C1704 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00403f
C1705 a_67618_24851# a2x1mux_mag_0.Transmission_gate_mag_0.CLK 5.79e-19
C1706 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.71e-21
C1707 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 3.21e-20
C1708 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C1709 a_66447_5529# RST_DIV 0.00247f
C1710 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_63994_5529# 0.0102f
C1711 a_61533_24598# VDD 3.14e-19
C1712 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.71e-21
C1713 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VCO_op 0.01f
C1714 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 5.7e-20
C1715 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 7.99e-19
C1716 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 2.89e-20
C1717 PFD_layout_0.buffer_mag_0.OUT VDD 1.9f
C1718 PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.QB 0.62f
C1719 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0231f
C1720 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_66293_4432# 1.86e-20
C1721 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_70752_5529# 5.02e-20
C1722 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 1.83f
C1723 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_69327_6404# 0.00789f
C1724 PFD_layout_0.DFF__0.nand2_2.IN2 VCO_mag_0.Delay_Cell_mag_1.INB 0.0104f
C1725 CP_mag_0.inv_0.OUT a2x1mux_mag_0.Transmission_gate_mag_0.CLK 1.28e-19
C1726 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 0.104f
C1727 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 RST_DIV 0.0573f
C1728 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VCO_op 0.0765f
C1729 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.11e-20
C1730 a_67611_25266# pd 0.00441f
C1731 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 0.158f
C1732 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J VDD 0.623f
C1733 PFD_layout_0.DFF__0.nand2_1.IN1 a_62434_21795# 1.63e-20
C1734 VCO_mag_0.VCONT VDD_VCO 2.16f
C1735 LF_mag_0.VCNTL a_61538_21913# 7.5e-19
C1736 a_67611_25266# VDD 0.771f
C1737 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.86e-19
C1738 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_68145_4432# 0.0114f
C1739 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.126f
C1740 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 5.55e-21
C1741 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 a_73620_7541# 0.069f
C1742 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0274f
C1743 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.DFF__0.nand2_1.IN1 4.77e-22
C1744 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_op 0.153f
C1745 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_72487_4432# 1.41e-20
C1746 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 0.195f
C1747 VCO_mag_0.GF_INV16_2.IN VCO_op_bar 0.00206f
C1748 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_60147_8532# 0.00765f
C1749 a_60147_8532# VCO_op 3.18e-19
C1750 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_68511_9745# 0.00476f
C1751 VCO_mag_0.Delay_Cell_mag_1.INB VCO_op_bar 0.0404f
C1752 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT RST_DIV 0.269f
C1753 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.311f
C1754 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0052f
C1755 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD 0.399f
C1756 a_63016_9651# VDD 0.165f
C1757 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C1758 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT 0.173f
C1759 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C1760 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C1761 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 3.89e-20
C1762 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_70216_3335# 3.38e-20
C1763 a_67618_24851# pd 0.144f
C1764 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_63430_5529# 0.00789f
C1765 a_66287_5529# RST_DIV 0.00247f
C1766 PFD_layout_0.VDIV a_59138_17829# 1.73e-19
C1767 a_67618_24851# VDD 0.018f
C1768 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_67735_5529# 0.0036f
C1769 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.432f
C1770 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN VDD 0.664f
C1771 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 8.28e-20
C1772 PFD_layout_0.buffer_mag_0.OUT VDD_VCO 2.66e-19
C1773 a_61552_8823# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C1774 VCO_mag_0.Delay_Cell_mag_2.IN VCO_mag_0.Delay_Cell_mag_1.INB 0.266f
C1775 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_65128_4432# 0.0114f
C1776 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_69167_6404# 0.00335f
C1777 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 3.4e-19
C1778 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VCO_op 0.276f
C1779 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C1780 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN 1.23e-19
C1781 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN 0.163f
C1782 LF_mag_0.VCNTL a_60302_21847# 3.1e-19
C1783 CP_mag_0.inv_0.OUT VDD 0.568f
C1784 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_72152_3335# 5.1e-20
C1785 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_70461_7545# 4.52e-20
C1786 CP_mag_0.inv_0.OUT pd 0.164f
C1787 PFD_layout_0.DFF__0.nand2_1.IN1 a_61538_21913# 0.00384f
C1788 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_67581_4432# 2.96e-19
C1789 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.57e-19
C1790 LF_mag_0.VCNTL a2x1mux_mag_0.Transmission_gate_mag_0.CLK 0.00135f
C1791 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 7.22e-20
C1792 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0593f
C1793 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00943f
C1794 a_59418_24365# PFD_layout_0.DFF__0.CLK 1.82e-19
C1795 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.0022f
C1796 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 5.7e-19
C1797 a_65581_14091# EN 0.201f
C1798 a_73620_7541# RST_DIV 1.31e-19
C1799 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_72327_4432# 1.86e-20
C1800 VCO_mag_0.Delay_Cell_mag_0.OUTB VCO_mag_0.Delay_Cell_mag_0.OUT 1.6f
C1801 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 4.08e-20
C1802 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_67806_9704# 0.00107f
C1803 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 5.73e-20
C1804 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0334f
C1805 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN 0.00147f
C1806 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 RST_DIV 0.182f
C1807 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_70615_6448# 0.00378f
C1808 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_67171_5529# 0.0101f
C1809 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00157f
C1810 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_74179_4432# 0.0114f
C1811 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C1812 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 1.9e-19
C1813 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_63270_5529# 0.00335f
C1814 a_71184_3335# VDD 3.14e-19
C1815 a_63452_24694# IPD+ 9.68e-20
C1816 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 RST_DIV 0.178f
C1817 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 RST_DIV 0.11f
C1818 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.0609f
C1819 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J a_62924_7501# 0.00472f
C1820 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.OUTB 0.263f
C1821 a_73210_6400# RST_DIV 0.0017f
C1822 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C1823 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_64564_4432# 2.96e-19
C1824 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C1825 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.198f
C1826 PFD_layout_0.DFF__1.nand2_5.OUT a_60304_24408# 3.83e-19
C1827 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C1828 LF_mag_0.VCNTL a_59585_21854# 3.72e-19
C1829 PFD_layout_0.nand2_0.IN1 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN 0.292f
C1830 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT RST_DIV 0.0779f
C1831 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD 0.392f
C1832 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VCO_op 0.271f
C1833 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_69897_7545# 0.0195f
C1834 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_67017_4432# 3.25e-19
C1835 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 9.58e-20
C1836 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VCO_op 7.37e-20
C1837 a2x1mux_mag_0.SEL IPD+ 2.52e-20
C1838 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C1839 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C1840 LF_mag_0.VCNTL pd 0.00248f
C1841 LF_mag_0.VCNTL VDD 6.19f
C1842 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_74338_6444# 0.00372f
C1843 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C1844 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 4.01e-20
C1845 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VDD 0.797f
C1846 PFD_layout_0.VDIV a_58943_20071# 5.72e-19
C1847 a_73056_7541# RST_DIV 4.54e-19
C1848 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_71162_4432# 0.0114f
C1849 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C1850 a_74333_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0811f
C1851 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_67646_9704# 0.00271f
C1852 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 5.42e-20
C1853 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_67011_5529# 0.0102f
C1854 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_70051_6404# 0.0733f
C1855 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VCO_op 0.00187f
C1856 a_70188_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0733f
C1857 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_73615_4432# 2.96e-19
C1858 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 0.191f
C1859 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD 0.913f
C1860 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_72487_4432# 0.00939f
C1861 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN 0.257f
C1862 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.25f
C1863 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C1864 VCO_mag_0.Delay_Cell_mag_0.IN EN 0.279f
C1865 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD 1f
C1866 a_60147_8532# VDD 2.21e-19
C1867 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 2.6e-20
C1868 PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.DFF__0.inv_0.OUT 4.23e-20
C1869 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 1.16f
C1870 a_74184_7541# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C1871 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.124f
C1872 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0309f
C1873 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C1874 a_73050_6400# RST_DIV 0.00199f
C1875 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_64000_4432# 3.33e-19
C1876 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 3.3e-19
C1877 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.61e-19
C1878 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.111f
C1879 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_64154_5529# 2.88e-20
C1880 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_68299_5529# 0.00372f
C1881 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 0.507f
C1882 VCO_mag_0.Delay_Cell_mag_0.IN a_65581_14091# 0.61f
C1883 PFD_layout_0.DFF__1.nand2_5.OUT a_59418_24365# 0.00432f
C1884 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00137f
C1885 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.252f
C1886 a_60147_7030# VCO_op 1.79e-19
C1887 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 5.24e-20
C1888 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.029f
C1889 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_74338_6444# 0.0811f
C1890 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 6.18e-19
C1891 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT RST_DIV 0.0979f
C1892 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_2.OUT 0.00326f
C1893 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0032f
C1894 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_73774_6444# 0.069f
C1895 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD 0.647f
C1896 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 RST_DIV 0.0189f
C1897 LF_mag_0.VCNTL VDD_VCO 0.408f
C1898 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00122f
C1899 PFD_layout_0.DFF__0.nand2_1.IN1 VDD 1.3f
C1900 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_69470_4432# 0.00939f
C1901 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_70598_4432# 2.96e-19
C1902 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.CLK 0.0528f
C1903 a_72492_7497# RST_DIV 0.002f
C1904 PFD_layout_0.DFF__0.nand2_2.IN1 VCO_mag_0.Delay_Cell_mag_2.INB 4.19e-19
C1905 a_67017_4432# RST_DIV 1.23e-20
C1906 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 4.54f
C1907 a_73769_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00964f
C1908 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 3.79e-20
C1909 PFD_layout_0.DFF__1.nand2_2.OUT PFD_layout_0.buffer_mag_0.OUT 0.0494f
C1910 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_69891_6404# 0.0203f
C1911 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_74338_6444# 0.0157f
C1912 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C1913 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_66447_5529# 0.00789f
C1914 a_70028_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0203f
C1915 a_71316_5529# VDD 0.00152f
C1916 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_74184_7541# 0.0114f
C1917 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 2.87e-19
C1918 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_73051_4432# 3.25e-19
C1919 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VCO_op 7.06e-20
C1920 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.487f
C1921 EN VCO_op_bar 0.325f
C1922 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_72327_4432# 0.0101f
C1923 a_59138_14091# EN 0.405f
C1924 a_67171_5529# VDD 0.00101f
C1925 VCO_mag_0.Delay_Cell_mag_2.OUTB VCO_op 0.0312f
C1926 VCO_mag_0.Delay_Cell_mag_0.OUTB VDD_VCO 3.63f
C1927 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.nand2_2.IN2 0.0065f
C1928 LF_mag_0.VCNTL a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT 0.0388f
C1929 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00164f
C1930 VCO_mag_0.GF_INV16_2.IN VCO_mag_0.Delay_Cell_mag_0.INB 8.2e-19
C1931 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.249f
C1932 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 RST_DIV 0.164f
C1933 PFD_layout_0.DFF__1.nand2_3.OUT a_61537_25977# 2.09e-19
C1934 a_59584_26036# PFD_layout_0.DFF__1.CLK 1.27e-19
C1935 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 6.36e-20
C1936 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C1937 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00127f
C1938 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VCO_op 0.00127f
C1939 a_72486_6400# RST_DIV 0.00256f
C1940 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C1941 PFD_layout_0.DFF__1.nand2_5.OUT a_62429_24598# 0.00454f
C1942 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_63994_5529# 9.1e-19
C1943 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_67735_5529# 0.069f
C1944 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C1945 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_74184_7541# 0.069f
C1946 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.205f
C1947 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_73774_6444# 0.00964f
C1948 VCO_mag_0.Delay_Cell_mag_2.IN EN 0.375f
C1949 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VCO_op 6.64e-19
C1950 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00544f
C1951 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C1952 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0349f
C1953 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.048f
C1954 a_60305_23482# VDD 4.85e-19
C1955 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C1956 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.236f
C1957 PFD_layout_0.DFF__0.nand2_1.IN1 VDD_VCO 2.05e-19
C1958 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C1959 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_69310_4432# 0.0101f
C1960 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_70461_7545# 0.0059f
C1961 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_70034_4432# 3.25e-19
C1962 a_72332_7497# RST_DIV 0.00274f
C1963 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 0.0224f
C1964 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN RST_DIV 0.0454f
C1965 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 2.48e-19
C1966 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD 0.642f
C1967 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0365f
C1968 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.74e-19
C1969 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD 0.741f
C1970 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD 0.653f
C1971 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VCO_op 1.84e-19
C1972 VCO_mag_0.Delay_Cell_mag_2.INB a_59138_17829# 0.499f
C1973 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_69327_6404# 1.5e-20
C1974 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_72492_7497# 1.88e-19
C1975 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.00525f
C1976 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_66287_5529# 0.00335f
C1977 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.27e-19
C1978 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00393f
C1979 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_73774_6444# 0.00859f
C1980 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_73620_7541# 2.96e-19
C1981 a_70752_5529# VDD 0.00152f
C1982 a_69464_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.5e-20
C1983 a_70028_5529# a_70188_5529# 0.0504f
C1984 a_65386_16333# EN 8.31e-20
C1985 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_71162_4432# 9.45e-19
C1986 PFD_layout_0.DFF__1.CLK VDD 1.12f
C1987 a_67011_5529# VDD 0.00123f
C1988 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.42e-19
C1989 a_58943_16333# VDD_VCO 0.846f
C1990 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN a_61544_9654# 2.7e-20
C1991 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN RST_DIV 0.00399f
C1992 PFD_layout_0.DFF__0.nand2_5.OUT PFD_layout_0.DFF__0.nand2_3.OUT 0.42f
C1993 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 1.87e-19
C1994 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0501f
C1995 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C1996 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 1.76e-21
C1997 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C1998 a_72326_6400# RST_DIV 0.00256f
C1999 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_61106_7416# 3.17e-19
C2000 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__1.nand2_3.OUT 0.0185f
C2001 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00916f
C2002 a_61106_7416# VCO_op 2.02e-20
C2003 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.159f
C2004 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT 0.205f
C2005 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT RST_DIV 0.102f
C2006 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 6.94e-19
C2007 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD 5.32f
C2008 PFD_layout_0.DFF__1.nand2_5.OUT a_61533_24598# 0.0703f
C2009 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.11f
C2010 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_63430_5529# 0.0731f
C2011 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_66453_4432# 9.32e-19
C2012 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_72486_6400# 0.00194f
C2013 PFD_layout_0.nand2_0.IN1 a_62429_24598# 0.00351f
C2014 a_73051_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN 5.94e-20
C2015 PFD_layout_0.DFF__0.QB PFD_layout_0.DFF__0.inv_0.OUT 0.00316f
C2016 PFD_layout_0.nand2_0.IN1 pu 0.00662f
C2017 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 RST_DIV 0.0409f
C2018 a2x1mux_mag_0.Transmission_gate_mag_0.CLK a2x1mux_mag_0.SEL 0.177f
C2019 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_73210_6400# 0.00696f
C2020 VCO_mag_0.VCONT a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT 0.166f
C2021 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__1.nand2_5.OUT 0.391f
C2022 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT a_61544_9654# 0.0202f
C2023 PFD_layout_0.buffer_mag_0.IN PFD_layout_0.buffer_loading_mag_1.IN 0.137f
C2024 a_69891_6404# a_70051_6404# 0.0504f
C2025 VCO_mag_0.Delay_Cell_mag_2.INB VCO_mag_0.Delay_Cell_mag_1.IN 0.245f
C2026 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 3.23f
C2027 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VCO_op 0.581f
C2028 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C2029 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_72152_3335# 0.01f
C2030 PFD_layout_0.DFF__1.inv_0.OUT PFD_layout_0.DFF__0.nand2_5.OUT 8.72e-22
C2031 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_68145_4432# 0.069f
C2032 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.57e-20
C2033 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_69897_7545# 0.0697f
C2034 a_71025_7545# RST_DIV 5.35e-19
C2035 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J a_62918_6404# 8.64e-19
C2036 a_60147_7030# VDD 3.14e-19
C2037 VCO_mag_0.GF_INV16_1.IN VCO_op 4.93e-19
C2038 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00125f
C2039 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 9.86e-19
C2040 a_69470_4432# VDD 2.66e-19
C2041 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 8.26e-20
C2042 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VCO_op 8.66e-20
C2043 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VCO_op 2.51e-20
C2044 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_72332_7497# 2.7e-19
C2045 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_61544_9654# 0.0186f
C2046 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_73210_6400# 0.0101f
C2047 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C2048 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.123f
C2049 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_69167_6404# 1.17e-20
C2050 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.88e-20
C2051 a_69304_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.17e-20
C2052 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_70598_4432# 6.06e-21
C2053 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C2054 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_73056_7541# 3.33e-19
C2055 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 1.08f
C2056 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.00584f
C2057 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 0.98f
C2058 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_68511_9745# 0.015f
C2059 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00152f
C2060 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_65128_4432# 0.00372f
C2061 a_63452_24694# pd 7.76e-19
C2062 a_66447_5529# VDD 0.00863f
C2063 a_63452_24694# VDD 1.2f
C2064 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 5.36e-20
C2065 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 0.00452f
C2066 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VCO_op 1.52e-20
C2067 LF_mag_0.VCNTL PFD_layout_0.DFF__0.CLK 3.38e-20
C2068 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_70051_6404# 8.64e-19
C2069 PFD_layout_0.DFF__1.nand2_2.IN1 a_60301_26043# 9.39e-21
C2070 a_71179_6448# RST_DIV 0.0013f
C2071 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 1.71e-21
C2072 a_74338_6444# VDD 3.14e-19
C2073 PFD_layout_0.DFF__0.nand2_2.OUT VCO_mag_0.Delay_Cell_mag_2.INB 5.75e-21
C2074 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_63270_5529# 0.0202f
C2075 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C2076 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_66293_4432# 0.00876f
C2077 a_74380_2641# VDD 0.0407f
C2078 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_72326_6400# 0.00194f
C2079 a_73056_7541# VCO_op 6.43e-21
C2080 a_65581_17830# VCO_op 0.0271f
C2081 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD 1.03f
C2082 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 2.22e-20
C2083 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT RST_DIV 0.00693f
C2084 a2x1mux_mag_0.Transmission_gate_mag_0.CLK a_63591_22645# 5.39e-20
C2085 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00265f
C2086 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_73050_6400# 0.00695f
C2087 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 5.2e-20
C2088 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.11f
C2089 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.nand2_0.IN1 0.375f
C2090 a2x1mux_mag_0.SEL VDD 0.725f
C2091 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J 2.21e-19
C2092 a2x1mux_mag_0.SEL pd 0.00306f
C2093 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT RST_DIV 0.285f
C2094 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.DFF__1.inv_0.OUT 0.155f
C2095 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_70034_4432# 0.00378f
C2096 a_69173_7501# a_69333_7501# 0.0504f
C2097 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.313f
C2098 VCO_mag_0.Delay_Cell_mag_2.INB a_58943_20071# 0.542f
C2099 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VDD 0.497f
C2100 PFD_layout_0.DFF__0.nand2_2.IN2 VCO_mag_0.Delay_Cell_mag_2.IN 9.39e-19
C2101 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_67581_4432# 6.06e-21
C2102 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_74220_2641# 2.85e-20
C2103 PFD_layout_0.DFF__0.nand2_3.OUT PFD_layout_0.DFF__0.nand2_2.IN2 0.0984f
C2104 PFD_layout_0.DFF__0.nand2_2.IN1 a_60302_21847# 9.39e-21
C2105 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C2106 a_70461_7545# RST_DIV 2.53e-19
C2107 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 2.67e-20
C2108 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.161f
C2109 VCO_mag_0.VCONT VCO_mag_0.GF_INV1_0.OUT 0.107f
C2110 a_74184_7541# VDD 3.56e-19
C2111 a_69310_4432# VDD 0.00746f
C2112 PFD_layout_0.DFF__1.QB PFD_layout_0.DFF__1.nand2_3.OUT 0.0138f
C2113 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_73050_6400# 0.0102f
C2114 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN a_71408_9766# 0.198f
C2115 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD 0.994f
C2116 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 1.17e-19
C2117 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_72327_4432# 6.36e-19
C2118 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.289f
C2119 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C2120 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_72492_7497# 0.00392f
C2121 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_71025_7545# 0.00118f
C2122 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_64564_4432# 0.069f
C2123 PFD_layout_0.DFF__0.QB a_62434_21795# 0.00619f
C2124 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.11e-21
C2125 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_67806_9704# 5.19e-20
C2126 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.45e-22
C2127 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN 3.09e-19
C2128 a_61537_25977# VDD 3.22e-19
C2129 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_63802_6404# 2.88e-20
C2130 a_66287_5529# VDD 0.0123f
C2131 VCO_mag_0.Delay_Cell_mag_2.IN a_59138_14091# 0.679f
C2132 VCO_mag_0.Delay_Cell_mag_2.IN VCO_op_bar 0.0635f
C2133 PFD_layout_0.DFF__0.CLK PFD_layout_0.DFF__0.nand2_1.IN1 0.114f
C2134 PFD_layout_0.DFF__1.nand2_2.IN1 a_59584_26036# 0.00348f
C2135 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_72481_5529# 0.00164f
C2136 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VCO_op 8.16e-19
C2137 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN a_71408_9766# 2.31e-19
C2138 a_70615_6448# RST_DIV 0.00129f
C2139 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.423f
C2140 a_73774_6444# VDD 3.14e-19
C2141 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_63084_7501# 1.03e-20
C2142 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C2143 a_74220_2641# VDD 0.234f
C2144 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0404f
C2145 VCO_mag_0.Delay_Cell_mag_0.INB EN 0.11f
C2146 a_65581_17830# VCO_mag_0.Delay_Cell_mag_0.OUT 0.324f
C2147 a_72492_7497# VCO_op 0.00939f
C2148 VCO_mag_0.Delay_Cell_mag_1.IN VCO_op 0.00695f
C2149 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C2150 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_72492_7497# 2.79e-20
C2151 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C2152 VCO_mag_0.Delay_Cell_mag_2.OUTB VDD_VCO 5.03f
C2153 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 RST_DIV 0.0784f
C2154 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.305f
C2155 a_63591_22645# pd 0.332f
C2156 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C2157 a_63591_22645# VDD 1.22f
C2158 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.136f
C2159 a_61106_7416# VDD 0.173f
C2160 a2x1mux_mag_0.SEL VDD_VCO 0.00895f
C2161 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT VDD 0.339f
C2162 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT 8.02e-19
C2163 a_58357_44128# LF_mag_0.res_48k_mag_0.B 0.113f
C2164 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 RST_DIV 0.0316f
C2165 VCO_mag_0.Delay_Cell_mag_0.INB a_65581_14091# 0.354f
C2166 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 1.87e-19
C2167 a_69897_7545# RST_DIV 3.68e-20
C2168 PFD_layout_0.DFF__0.nand2_2.IN1 a_59585_21854# 0.00348f
C2169 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 RST_DIV 9.24e-20
C2170 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 8.28e-20
C2171 a_73620_7541# VDD 3.14e-19
C2172 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C2173 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 2.27e-20
C2174 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VCO_op 9.85e-20
C2175 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00209f
C2176 a_68145_4432# VDD 3.56e-19
C2177 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00425f
C2178 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN a_71248_9766# 0.0135f
C2179 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_71162_4432# 0.069f
C2180 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_72486_6400# 0.00789f
C2181 a_72486_6400# VCO_op 0.00164f
C2182 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT 3.41e-19
C2183 a_66453_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0732f
C2184 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD 3.46f
C2185 PFD_layout_0.DFF__0.nand2_2.IN1 VDD 0.918f
C2186 VCO_mag_0.VCONT LP_ext 3.96f
C2187 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_70461_7545# 0.011f
C2188 a2x1mux_mag_0.SEL a2x1mux_mag_0.Transmission_gate_mag_0.inv_my_mag_0.OUT 0.00848f
C2189 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 3.8e-20
C2190 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_67646_9704# 3.35e-20
C2191 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_63642_6404# 9.1e-19
C2192 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C2193 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD 0.653f
C2194 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_72321_5529# 0.00117f
C2195 PFD_layout_0.DFF__0.CLK a_60305_23482# 0.00347f
C2196 PFD_layout_0.DFF__1.nand2_2.IN1 VDD 0.942f
C2197 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C2198 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VDD 2.86f
C2199 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN a_71248_9766# 3.59e-19
C2200 a_70051_6404# RST_DIV 0.00216f
C2201 a_69464_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.46e-19
C2202 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 1.97f
C2203 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN a_60140_9217# 0.069f
C2204 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0286f
C2205 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_62924_7501# 1.29e-20
C2206 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_73205_5529# 2.88e-20
C2207 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_63436_4432# 2.79e-20
C2208 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_1.INB 0.317f
C2209 LF_mag_0.VCNTL a_56917_44128# 0.0767f
C2210 a_72332_7497# VCO_op 0.0101f
C2211 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT RST_DIV 0.00758f
C2212 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN 6.99e-20
C2213 VCO_mag_0.VCONT VCO_mag_0.GF_INV16_2.IN 0.0245f
C2214 VCO_mag_0.Delay_Cell_mag_1.IN VCO_mag_0.Delay_Cell_mag_0.OUT 0.257f
C2215 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD 0.792f
C2216 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00586f
C2217 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_70615_6448# 0.0036f
C2218 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_72152_3335# 0.0096f
C2219 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT a_71408_9766# 2.84e-20
C2220 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 2.84e-20
C2221 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C2222 a_62430_23292# VDD 4.2e-19
C2223 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C2224 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 7.38e-19
C2225 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 1.86e-19
C2226 PFD_layout_0.DFF__1.CLK PFD_layout_0.DFF__0.CLK 0.00128f
C2227 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT 0.00125f
C2228 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 7.16e-20
C2229 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.211f
C2230 LF_mag_0.VCNTL a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT 0.61f
C2231 VCO_mag_0.Delay_Cell_mag_2.OUT VDD_VCO 4.23f
C2232 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.61e-19
C2233 a_73056_7541# VDD 3.14e-19
C2234 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 1.77e-19
C2235 PFD_layout_0.DFF__1.nand2_2.OUT PFD_layout_0.DFF__1.CLK 0.00375f
C2236 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 0.00441f
C2237 a_67581_4432# VDD 3.14e-19
C2238 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 3.21e-20
C2239 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_72326_6400# 0.00335f
C2240 PFD_layout_0.buffer_mag_0.gf_inv_mag_1.IN PFD_layout_0.DFF__0.nand2_5.OUT 3.54e-19
C2241 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_70598_4432# 0.0059f
C2242 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__0.nand2_1.IN1 2.09e-19
C2243 a_72326_6400# VCO_op 0.00117f
C2244 a_59419_23525# VDD 0.00503f
C2245 PFD_layout_0.DFF__0.nand2_2.IN1 VDD_VCO 2.44e-19
C2246 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 8.64e-20
C2247 a_69304_5529# a_69464_5529# 0.0504f
C2248 a_66293_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0203f
C2249 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C2250 VCO_mag_0.Delay_Cell_mag_0.INB VCO_mag_0.Delay_Cell_mag_0.IN 0.899f
C2251 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_69897_7545# 1.43e-19
C2252 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VCO_op 0.235f
C2253 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_73045_5529# 3.6e-22
C2254 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-20
C2255 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_63078_6404# 0.0731f
C2256 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_60140_9217# 0.00544f
C2257 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.57e-20
C2258 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00301f
C2259 PFD_layout_0.buffer_loading_mag_1.IN PFD_layout_0.DFF__0.inv_0.OUT 5.29e-19
C2260 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0515f
C2261 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 6.69e-19
C2262 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.00274f
C2263 PFD_layout_0.DFF__1.nand2_3.OUT PFD_layout_0.DFF__1.nand2_1.IN1 0.39f
C2264 VCO_mag_0.GF_INV1_1.OUT VDD_VCO 0.888f
C2265 VCO_mag_0.GF_INV16_1.IN VDD_VCO 1.58f
C2266 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_72487_4432# 2.79e-20
C2267 a_69891_6404# RST_DIV 0.00199f
C2268 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C2269 PFD_layout_0.DFF__0.nand2_2.OUT a_60302_21847# 0.00364f
C2270 a_73050_6400# VDD 2.21e-19
C2271 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_73045_5529# 9.1e-19
C2272 a_71025_7545# VCO_op 9.36e-19
C2273 LF_mag_0.VCNTL a_56677_42026# 0.0161f
C2274 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD 0.769f
C2275 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT a_71248_9766# 9.09e-19
C2276 a_69167_6404# a_69327_6404# 0.0504f
C2277 a_58117_42026# a_58597_42026# 0.0754f
C2278 a_67618_24851# LP_ext 6.98e-20
C2279 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J 0.0579f
C2280 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00359f
C2281 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_63016_9651# 0.0131f
C2282 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD 0.395f
C2283 a_65386_20072# VDD 0.171f
C2284 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0998f
C2285 a_65581_17830# VDD_VCO 0.0996f
C2286 PFD_layout_0.DFF__1.QB VDD 1.14f
C2287 VCO_mag_0.Delay_Cell_mag_1.IN VDD 0.00731f
C2288 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 7.97e-19
C2289 a_67017_4432# VDD 3.14e-19
C2290 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00117f
C2291 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 RST_DIV 0.187f
C2292 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C2293 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_69333_7501# 1.87e-19
C2294 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_70034_4432# 0.0697f
C2295 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_69333_7501# 0.00119f
C2296 LF_mag_0.VCNTL VCO_mag_0.GF_INV1_0.OUT 0.00161f
C2297 a_66293_4432# a_66453_4432# 0.0504f
C2298 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_72481_5529# 1.86e-20
C2299 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 1.32e-19
C2300 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_62918_6404# 0.0202f
C2301 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_63016_9651# 0.0115f
C2302 a_59138_17829# VDD_VCO 0.152f
C2303 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 RST_DIV 0.179f
C2304 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VCO_op 0.0833f
C2305 a_69327_6404# RST_DIV 0.00257f
C2306 PFD_layout_0.DFF__0.QB VDD 1.11f
C2307 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD 0.66f
C2308 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 3.94e-19
C2309 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0377f
C2310 a_68299_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0811f
C2311 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.116f
C2312 PFD_layout_0.DFF__0.nand2_2.OUT a_59585_21854# 0.069f
C2313 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 a_71025_7545# 0.00372f
C2314 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 0.306f
C2315 PFD_layout_0.DFF__1.CLK PFD_layout_0.DFF__1.nand2_5.OUT 0.115f
C2316 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0569f
C2317 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C2318 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0502f
C2319 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_72481_5529# 0.0731f
C2320 a_70461_7545# VCO_op 9.24e-19
C2321 PFD_layout_0.DFF__0.nand2_2.OUT VDD 0.39f
C2322 a_64154_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C2323 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 2.25e-21
C2324 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB RST_DIV 0.182f
C2325 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_71408_9766# 8.64e-19
C2326 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00107f
C2327 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 9.75e-21
C2328 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C2329 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST_DIV 0.288f
C2330 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C2331 PFD_layout_0.buffer_loading_mag_1.IN a_62434_21795# 0.069f
C2332 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT 4.11e-19
C2333 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.7e-19
C2334 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.61e-20
C2335 a_72332_7497# VDD 2.21e-19
C2336 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 RST_DIV 3.32e-19
C2337 PFD_layout_0.DFF__1.nand2_2.IN2 a_60304_24408# 2.82e-20
C2338 a_65386_20072# VDD_VCO 1.13f
C2339 VCO_mag_0.Delay_Cell_mag_1.IN VDD_VCO 4.34f
C2340 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_2.IN VDD 0.345f
C2341 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_69173_7501# 2.69e-19
C2342 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C2343 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C2344 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 3.79e-19
C2345 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.89e-20
C2346 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 5.6e-19
C2347 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 5.63e-21
C2348 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_72321_5529# 2.55e-20
C2349 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0399f
C2350 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VCO_op 0.416f
C2351 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C2352 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C2353 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD 0.516f
C2354 a_61534_23292# VDD 3.14e-19
C2355 LF_mag_0.VCNTL LP_ext 0.253f
C2356 a_69167_6404# RST_DIV 0.00257f
C2357 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C2358 a_72326_6400# VDD 2.21e-19
C2359 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.768f
C2360 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 0.341f
C2361 a_67735_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00964f
C2362 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 a_70461_7545# 0.069f
C2363 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_60307_8532# 8.95e-19
C2364 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VCO_op 0.01f
C2365 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD 0.642f
C2366 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0432f
C2367 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00158f
C2368 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 RST_DIV 0.152f
C2369 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_69327_6404# 0.00192f
C2370 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_73205_5529# 0.0101f
C2371 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_72321_5529# 0.0202f
C2372 a_69897_7545# VCO_op 3.8e-19
C2373 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 VDD 1.18f
C2374 a_63994_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C2375 a_64776_7545# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C2376 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.11e-19
C2377 PFD_layout_0.DFF__0.nand2_2.IN1 PFD_layout_0.DFF__0.CLK 0.145f
C2378 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_69327_6404# 1.46e-19
C2379 PFD_layout_0.DFF__0.nand2_2.OUT VDD_VCO 3.19e-19
C2380 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 1.96f
C2381 a_68299_5529# RST_DIV 0.00122f
C2382 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C2383 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT 1.5e-20
C2384 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_71248_9766# 0.0105f
C2385 VCO_mag_0.VCONT EN 1.24f
C2386 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0151f
C2387 LF_mag_0.VCNTL VCO_mag_0.Delay_Cell_mag_1.INB 0.321f
C2388 PFD_layout_0.VDIV VCO_mag_0.Delay_Cell_mag_2.INB 0.0612f
C2389 a_64154_5529# RST_DIV 0.00283f
C2390 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C2391 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__0.CLK 4.55e-19
C2392 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C2393 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.71e-21
C2394 PFD_layout_0.DFF__1.nand2_2.IN2 a_59418_24365# 1.16e-20
C2395 PFD_layout_0.buffer_loading_mag_1.IN a_61538_21913# 1.06e-19
C2396 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C2397 a_71025_7545# VDD 3.56e-19
C2398 a_58943_20071# VDD_VCO 1.12f
C2399 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.12e-19
C2400 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 2.97e-20
C2401 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J 2.8e-19
C2402 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C2403 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__1.nand2_2.OUT 0.451f
C2404 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 9.82e-21
C2405 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 0.00392f
C2406 VCO_mag_0.VCONT a_65581_14091# 0.0688f
C2407 IPD_ IPD+ 0.145f
C2408 PFD_layout_0.DFF__1.nand2_1.IN1 VDD 1.3f
C2409 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.J 4.68e-20
C2410 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_0.OUTB 0.316f
C2411 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00187f
C2412 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT VCO_op 0.00104f
C2413 VCO_mag_0.GF_INV16_2.IN VCO_mag_0.Delay_Cell_mag_0.OUTB 0.0157f
C2414 a_68065_6446# RST_DIV 0.00129f
C2415 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_74380_2641# 2.44e-20
C2416 a_71179_6448# VDD 3.14e-19
C2417 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.07e-20
C2418 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 5.98e-20
C2419 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_64154_5529# 8.64e-19
C2420 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_71408_9766# 0.0504f
C2421 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_73045_5529# 0.0102f
C2422 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 8.26e-20
C2423 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 8.94e-19
C2424 PFD_layout_0.nand2_0.IN1 a_63452_24694# 0.365f
C2425 a_69333_7501# VCO_op 0.0105f
C2426 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_69167_6404# 0.00192f
C2427 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_63016_9651# 8.64e-19
C2428 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C2429 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.OUT VDD 0.515f
C2430 a_63994_5529# a_64154_5529# 0.0504f
C2431 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 RST_DIV 0.192f
C2432 a_63430_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C2433 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 7e-19
C2434 a_59419_23525# PFD_layout_0.DFF__0.CLK 9.59e-19
C2435 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_68511_9745# 6.43e-19
C2436 a_67735_5529# RST_DIV 0.00119f
C2437 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD 0.995f
C2438 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_65282_5529# 0.0157f
C2439 a_63994_5529# RST_DIV 0.00283f
C2440 a2x1mux_mag_0.SEL a2x1mux_mag_0.Transmission_gate_mag_1.inv_my_mag_0.OUT 0.234f
C2441 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.08e-20
C2442 a_66783_7543# RST_DIV 3.08e-20
C2443 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_71184_3335# 5.1e-20
C2444 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_70188_5529# 2.88e-20
C2445 a_70461_7545# VDD 3.14e-19
C2446 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.IN 4.36e-19
C2447 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 5.25e-20
C2448 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C2449 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 3.32e-20
C2450 a_73615_4432# CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 5.94e-20
C2451 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.nand2_5.OUT 0.389f
C2452 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 RST_DIV 0.56f
C2453 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT 0.0444f
C2454 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT VCO_op 2.39e-19
C2455 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 3.83e-19
C2456 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 1.03e-19
C2457 VCO_mag_0.Delay_Cell_mag_1.INB a_58943_16333# 1.77e-19
C2458 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 1.4e-20
C2459 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C2460 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 RST_DIV 0.072f
C2461 a_67501_6446# RST_DIV 0.00129f
C2462 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__0.nand2_2.IN1 4.94e-19
C2463 a_70615_6448# VDD 3.14e-19
C2464 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C2465 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_0.IN 0.0304f
C2466 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_74220_2641# 9.02e-19
C2467 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_71248_9766# 0.0186f
C2468 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C2469 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_72481_5529# 0.00789f
C2470 PFD_layout_0.nand2_0.IN1 a_61537_25977# 1.06e-19
C2471 a_69173_7501# VCO_op 0.0114f
C2472 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 1.64e-20
C2473 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 6.04e-21
C2474 PFD_layout_0.DFF__1.nand2_2.IN1 PFD_layout_0.DFF__1.nand2_5.OUT 0.492f
C2475 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_71162_4432# 0.00372f
C2476 a_63270_5529# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C2477 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.16f
C2478 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.0529f
C2479 PFD_layout_0.VDIV VCO_op 1.51f
C2480 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 3.56e-19
C2481 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VCO_op 0.0846f
C2482 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C2483 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 3.25e-19
C2484 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_64718_5529# 0.00859f
C2485 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN 0.00982f
C2486 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0263f
C2487 a_63430_5529# RST_DIV 0.0037f
C2488 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C2489 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 5.68e-19
C2490 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_70028_5529# 9.1e-19
C2491 a_69897_7545# VDD 3.14e-19
C2492 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 2.75e-19
C2493 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.397f
C2494 LF_mag_0.res_48k_mag_0.B VDD 0.812f
C2495 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VCO_op 1.45f
C2496 PFD_layout_0.DFF__1.nand2_2.IN2 PFD_layout_0.buffer_mag_0.OUT 0.0259f
C2497 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.128f
C2498 a_69327_6404# VCO_op 0.00164f
C2499 PFD_layout_0.nand2_0.IN1 a_63591_22645# 5.62e-19
C2500 PFD_layout_0.buffer_loading_mag_1.IN VDD 2.88f
C2501 PFD_layout_0.buffer_loading_mag_1.IN pd 0.0708f
C2502 a_71408_9766# RST_DIV 0.00416f
C2503 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 RST_DIV 0.0717f
C2504 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C2505 PFD_layout_0.DFF__0.CLK PFD_layout_0.DFF__0.nand2_2.OUT 0.00375f
C2506 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 8.58e-20
C2507 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_64776_7545# 0.069f
C2508 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_64930_6448# 0.00372f
C2509 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.221f
C2510 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.OUT 1.93f
C2511 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 7.94e-20
C2512 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C2513 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 3.87e-19
C2514 a_66937_6402# RST_DIV 0.00216f
C2515 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.407f
C2516 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 2.04e-19
C2517 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 RST_DIV 0.00146f
C2518 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 1.85e-19
C2519 VCO_mag_0.VCONT a_59138_14091# 0.0346f
C2520 VCO_mag_0.VCONT VCO_op_bar 0.00171f
C2521 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_72321_5529# 0.00335f
C2522 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VCO_op 9.92e-20
C2523 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 0.0659f
C2524 a_67911_7543# VCO_op 9.33e-19
C2525 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VCO_op 1.48e-20
C2526 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C2527 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.11f
C2528 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_70598_4432# 0.069f
C2529 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 1.96f
C2530 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 2.6e-19
C2531 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT VDD 0.304f
C2532 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_66213_6402# 4.52e-19
C2533 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 3.38e-19
C2534 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 1.86e-19
C2535 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C2536 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.nand2_2.IN2 0.0259f
C2537 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.94e-20
C2538 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT RST_DIV 0.00229f
C2539 a_63270_5529# RST_DIV 0.00334f
C2540 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C2541 PFD_layout_0.DFF__1.CLK Vref 0.123f
C2542 VCO_mag_0.VCONT VCO_mag_0.Delay_Cell_mag_2.IN 0.0301f
C2543 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_69464_5529# 0.0731f
C2544 a_58597_42026# VDD 0.379f
C2545 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_63430_5529# 0.00164f
C2546 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 a_66219_7499# 1.88e-19
C2547 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.77e-20
C2548 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 3.26e-20
C2549 a_69167_6404# VCO_op 0.00117f
C2550 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.06e-19
C2551 a_71248_9766# RST_DIV 0.00402f
C2552 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C2553 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_64366_6448# 0.069f
C2554 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C2555 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.15e-20
C2556 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT a_61106_7416# 0.0178f
C2557 PFD_layout_0.DFF__1.QB PFD_layout_0.DFF__1.nand2_5.OUT 0.581f
C2558 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB RST_DIV 0.147f
C2559 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.415f
C2560 a2x1mux_mag_0.SEL LP_ext 0.00419f
C2561 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 8.71e-20
C2562 PFD_layout_0.VDIV CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.74e-19
C2563 a_66777_6402# RST_DIV 0.00199f
C2564 a_69891_6404# VDD 2.21e-19
C2565 VCO_mag_0.VCONT a_65386_16333# 0.104f
C2566 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 1.19e-19
C2567 VCO_mag_0.Delay_Cell_mag_0.OUTB EN 0.0652f
C2568 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.IN 0.0238f
C2569 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_0.OUT VDD 0.69f
C2570 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Vdiv11 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 1.79e-19
C2571 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0835f
C2572 a_67347_7543# VCO_op 9.25e-19
C2573 VCO_mag_0.GF_INV1_0.OUT VCO_mag_0.GF_INV16_1.IN 0.00101f
C2574 LF_mag_0.VCNTL PFD_layout_0.DFF__0.nand2_5.OUT 2.83e-19
C2575 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.OUT 3.8e-20
C2576 VCO_mag_0.Delay_Cell_mag_1.INB VCO_mag_0.Delay_Cell_mag_2.OUTB 0.00334f
C2577 VCO_mag_0.GF_INV1_1.OUT VCO_mag_0.GF_INV1_0.OUT 0.00589f
C2578 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_68299_5529# 0.0157f
C2579 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.25f
C2580 PFD_layout_0.buffer_mag_0.OUT VCO_mag_0.Delay_Cell_mag_2.IN 2.48e-19
C2581 PFD_layout_0.DFF__1.nand2_5.OUT PFD_layout_0.DFF__0.QB 1.82e-20
C2582 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_66053_6402# 5.83e-19
C2583 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0334f
C2584 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 RST_DIV 0.119f
C2585 VCO_op RST_DIV 3.82f
C2586 PFD_layout_0.buffer_mag_0.OUT PFD_layout_0.DFF__0.nand2_3.OUT 0.889f
C2587 PFD_layout_0.buffer_mag_0.IN pd 0.0044f
C2588 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 7.43e-20
C2589 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.49e-20
C2590 PFD_layout_0.buffer_mag_0.IN VDD 0.838f
C2591 a_57877_44128# a_58357_44128# 0.0759f
.ends

