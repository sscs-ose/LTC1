magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2357 -2097 2357 2097
<< psubdiff >>
rect -357 75 357 97
rect -357 29 -335 75
rect -289 29 -231 75
rect -185 29 -127 75
rect -81 29 -23 75
rect 23 29 81 75
rect 127 29 185 75
rect 231 29 289 75
rect 335 29 357 75
rect -357 -29 357 29
rect -357 -75 -335 -29
rect -289 -75 -231 -29
rect -185 -75 -127 -29
rect -81 -75 -23 -29
rect 23 -75 81 -29
rect 127 -75 185 -29
rect 231 -75 289 -29
rect 335 -75 357 -29
rect -357 -97 357 -75
<< psubdiffcont >>
rect -335 29 -289 75
rect -231 29 -185 75
rect -127 29 -81 75
rect -23 29 23 75
rect 81 29 127 75
rect 185 29 231 75
rect 289 29 335 75
rect -335 -75 -289 -29
rect -231 -75 -185 -29
rect -127 -75 -81 -29
rect -23 -75 23 -29
rect 81 -75 127 -29
rect 185 -75 231 -29
rect 289 -75 335 -29
<< metal1 >>
rect -346 75 346 86
rect -346 29 -335 75
rect -289 29 -231 75
rect -185 29 -127 75
rect -81 29 -23 75
rect 23 29 81 75
rect 127 29 185 75
rect 231 29 289 75
rect 335 29 346 75
rect -346 -29 346 29
rect -346 -75 -335 -29
rect -289 -75 -231 -29
rect -185 -75 -127 -29
rect -81 -75 -23 -29
rect 23 -75 81 -29
rect 127 -75 185 -29
rect 231 -75 289 -29
rect 335 -75 346 -29
rect -346 -86 346 -75
<< end >>
