* NGSPICE file created from CM_MSB_flat.ext - technology: gf180mcuC

.subckt CM_MSB_flat IM_T IM VSS OUT SD
X0 SD IM.t0 VSS.t127 VSS.t77 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X1 VSS IM.t1 SD.t79 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X2 SD IM_T.t0 OUT.t63 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X3 OUT IM_T.t1 SD.t81 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X4 VSS IM.t2 SD.t78 VSS.t59 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X5 OUT IM_T.t2 SD.t11 VSS.t10 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1.2u
X6 SD IM.t3 VSS.t122 VSS.t3 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X7 OUT IM_T.t3 SD.t104 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X8 SD IM.t4 VSS.t121 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=1.2u
X9 VSS IM.t5 SD.t75 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X10 VSS IM.t6 SD.t74 VSS.t75 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X11 SD IM_T.t4 OUT.t59 VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X12 OUT IM_T.t5 SD.t88 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X13 OUT IM_T.t6 SD.t92 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X14 VSS IM.t7 SD.t73 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X15 SD IM_T.t7 OUT.t56 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=1.2u
X16 SD IM.t8 VSS.t114 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X17 SD IM_T.t8 OUT.t55 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X18 SD IM_T.t9 OUT.t54 VSS.t77 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X19 SD IM_T.t10 OUT.t53 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X20 OUT IM_T.t11 SD.t93 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X21 SD IM_T.t12 OUT.t51 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X22 VSS IM.t9 SD.t71 VSS.t62 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X23 VSS IM.t10 SD.t70 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X24 VSS IM.t11 SD.t69 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X25 SD IM_T.t13 OUT.t50 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X26 SD IM_T.t14 OUT.t49 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X27 OUT IM_T.t15 SD.t122 VSS.t27 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X28 OUT IM_T.t16 SD.t115 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X29 VSS IM.t12 SD.t68 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X30 OUT IM_T.t17 SD.t125 VSS.t75 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X31 SD IM_T.t18 OUT.t45 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X32 VSS IM.t13 SD.t67 VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X33 OUT IM_T.t19 SD.t97 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X34 SD IM.t14 VSS.t103 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X35 SD IM_T.t20 OUT.t43 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X36 VSS IM.t15 SD.t65 VSS.t10 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1.2u
X37 VSS IM.t16 SD.t64 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X38 SD IM_T.t21 OUT.t42 VSS.t14 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X39 SD IM.t17 VSS.t90 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X40 SD IM_T.t22 OUT.t41 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X41 VSS IM.t18 SD.t62 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X42 OUT IM_T.t23 SD.t113 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X43 VSS IM.t19 SD.t61 VSS.t10 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1.2u
X44 OUT IM_T.t24 SD.t96 VSS.t59 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X45 SD IM.t20 VSS.t89 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X46 VSS IM.t21 SD.t59 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X47 OUT IM_T.t25 SD.t118 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X48 VSS IM.t22 SD.t58 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X49 SD IM_T.t26 OUT.t37 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X50 OUT IM_T.t27 SD.t4 VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X51 SD IM.t23 VSS.t86 VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X52 SD IM.t24 VSS.t85 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=1.2u
X53 SD IM_T.t28 OUT.t35 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X54 SD IM.t25 VSS.t84 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X55 OUT IM_T.t29 SD.t8 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X56 SD IM_T.t30 OUT.t33 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X57 SD IM.t26 VSS.t78 VSS.t77 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X58 SD IM.t27 VSS.t83 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X59 VSS IM.t28 SD.t52 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X60 SD IM_T.t31 OUT.t32 VSS.t3 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X61 OUT IM_T.t32 SD.t82 VSS.t62 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X62 SD IM.t29 VSS.t80 VSS.t3 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X63 OUT IM_T.t33 SD.t103 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X64 VSS IM.t30 SD.t50 VSS.t75 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X65 SD IM_T.t34 OUT.t29 VSS.t14 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X66 VSS IM.t31 SD.t49 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X67 OUT IM_T.t35 SD.t0 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X68 VSS IM.t32 SD.t48 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X69 OUT IM_T.t36 SD.t1 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X70 SD IM_T.t37 OUT.t26 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X71 SD IM_T.t38 OUT.t25 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X72 SD IM.t33 VSS.t70 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X73 SD IM_T.t39 OUT.t24 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X74 SD IM.t34 VSS.t69 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X75 OUT IM_T.t40 SD.t99 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X76 SD IM_T.t41 OUT.t22 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X77 SD IM.t35 VSS.t68 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X78 SD IM.t36 VSS.t67 VSS.t14 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X79 OUT IM_T.t42 SD.t121 VSS.t59 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X80 SD IM_T.t43 OUT.t20 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X81 SD IM.t37 VSS.t66 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X82 SD IM.t38 VSS.t65 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X83 OUT IM_T.t44 SD.t85 VSS.t27 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X84 SD IM_T.t45 OUT.t18 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X85 VSS IM.t39 SD.t41 VSS.t62 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X86 OUT IM_T.t46 SD.t102 VSS.t10 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1.2u
X87 OUT IM_T.t47 SD.t13 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X88 VSS IM.t40 SD.t40 VSS.t59 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X89 OUT IM_T.t48 SD.t98 VSS.t87 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X90 VSS IM.t41 SD.t39 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X91 VSS IM.t42 SD.t38 VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X92 VSS IM.t43 SD.t37 VSS.t12 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X93 SD IM.t44 VSS.t50 VSS.t8 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X94 SD IM_T.t49 OUT.t14 VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=1.2u
X95 VSS IM.t45 SD.t35 VSS.t27 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X96 SD IM_T.t50 OUT.t13 VSS.t77 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X97 SD IM.t46 VSS.t23 VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X98 VSS IM.t47 SD.t33 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X99 OUT IM_T.t51 SD.t101 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X100 SD IM_T.t52 OUT.t11 VSS.t3 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X101 OUT IM_T.t53 SD.t84 VSS.t75 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X102 VSS IM.t48 SD.t32 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X103 OUT IM_T.t54 SD.t108 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X104 VSS IM.t49 SD.t31 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X105 SD IM.t50 VSS.t36 VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X106 SD IM.t51 VSS.t42 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X107 SD IM_T.t55 OUT.t8 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X108 SD IM.t52 VSS.t40 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X109 SD IM.t53 VSS.t39 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X110 SD IM.t54 VSS.t34 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X111 VSS IM.t55 SD.t25 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X112 OUT IM_T.t56 SD.t90 VSS.t62 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X113 SD IM_T.t57 OUT.t6 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X114 SD IM.t56 VSS.t30 VSS.t29 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X115 VSS IM.t57 SD.t23 VSS.t27 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X116 OUT IM_T.t58 SD.t6 VSS.t6 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X117 SD IM.t58 VSS.t26 VSS.t25 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X118 OUT IM_T.t59 SD.t7 VSS.t1 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X119 VSS IM.t59 SD.t21 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X120 SD IM.t60 VSS.t19 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X121 OUT IM_T.t60 SD.t16 VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X122 SD IM_T.t61 OUT.t2 VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X123 SD IM.t61 VSS.t18 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X124 SD IM_T.t62 OUT.t1 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X125 SD IM.t62 VSS.t17 VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X126 SD IM_T.t63 OUT.t0 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
X127 SD IM.t63 VSS.t15 VSS.t14 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1.2u
R0 IM.n64 IM.n30 42.4777
R1 IM.n63 IM.n61 41.09
R2 IM.n0 IM.t19 33.0683
R3 IM.n31 IM.t15 33.0683
R4 IM.n3 IM.n2 32.0551
R5 IM.n7 IM.n6 32.0551
R6 IM.n11 IM.n10 32.0551
R7 IM.n15 IM.n14 32.0551
R8 IM.n19 IM.n18 32.0551
R9 IM.n23 IM.n22 32.0551
R10 IM.n27 IM.n26 32.0551
R11 IM.n34 IM.n33 32.0551
R12 IM.n38 IM.n37 32.0551
R13 IM.n42 IM.n41 32.0551
R14 IM.n46 IM.n45 32.0551
R15 IM.n50 IM.n49 32.0551
R16 IM.n54 IM.n53 32.0551
R17 IM.n58 IM.n57 32.0551
R18 IM.n4 IM.n3 31.2433
R19 IM.n8 IM.n7 31.2433
R20 IM.n12 IM.n11 31.2433
R21 IM.n16 IM.n15 31.2433
R22 IM.n20 IM.n19 31.2433
R23 IM.n24 IM.n23 31.2433
R24 IM.n28 IM.n27 31.2433
R25 IM.n35 IM.n34 31.2433
R26 IM.n39 IM.n38 31.2433
R27 IM.n43 IM.n42 31.2433
R28 IM.n47 IM.n46 31.2433
R29 IM.n51 IM.n50 31.2433
R30 IM.n55 IM.n54 31.2433
R31 IM.n59 IM.n58 31.2433
R32 IM.n2 IM.n1 31.2433
R33 IM.n6 IM.n5 31.2433
R34 IM.n10 IM.n9 31.2433
R35 IM.n14 IM.n13 31.2433
R36 IM.n18 IM.n17 31.2433
R37 IM.n22 IM.n21 31.2433
R38 IM.n26 IM.n25 31.2433
R39 IM.n30 IM.n29 31.2433
R40 IM.n33 IM.n32 31.2433
R41 IM.n37 IM.n36 31.2433
R42 IM.n41 IM.n40 31.2433
R43 IM.n45 IM.n44 31.2433
R44 IM.n49 IM.n48 31.2433
R45 IM.n53 IM.n52 31.2433
R46 IM.n57 IM.n56 31.2433
R47 IM.n61 IM.n60 31.2433
R48 IM.n1 IM.n0 30.4315
R49 IM.n5 IM.n4 30.4315
R50 IM.n9 IM.n8 30.4315
R51 IM.n13 IM.n12 30.4315
R52 IM.n17 IM.n16 30.4315
R53 IM.n21 IM.n20 30.4315
R54 IM.n25 IM.n24 30.4315
R55 IM.n29 IM.n28 30.4315
R56 IM.n32 IM.n31 30.4315
R57 IM.n36 IM.n35 30.4315
R58 IM.n40 IM.n39 30.4315
R59 IM.n44 IM.n43 30.4315
R60 IM.n48 IM.n47 30.4315
R61 IM.n52 IM.n51 30.4315
R62 IM.n56 IM.n55 30.4315
R63 IM.n60 IM.n59 30.4315
R64 IM.n64 IM.n63 2.2505
R65 IM.n0 IM.t63 1.8255
R66 IM.n1 IM.t59 1.8255
R67 IM.n2 IM.t52 1.8255
R68 IM.n3 IM.t48 1.8255
R69 IM.n4 IM.t26 1.8255
R70 IM.n5 IM.t2 1.8255
R71 IM.n6 IM.t14 1.8255
R72 IM.n7 IM.t12 1.8255
R73 IM.n8 IM.t50 1.8255
R74 IM.n9 IM.t30 1.8255
R75 IM.n10 IM.t46 1.8255
R76 IM.n11 IM.t18 1.8255
R77 IM.n12 IM.t61 1.8255
R78 IM.n13 IM.t55 1.8255
R79 IM.n14 IM.t51 1.8255
R80 IM.n15 IM.t1 1.8255
R81 IM.n16 IM.t29 1.8255
R82 IM.n17 IM.t42 1.8255
R83 IM.n18 IM.t56 1.8255
R84 IM.n19 IM.t9 1.8255
R85 IM.n20 IM.t53 1.8255
R86 IM.n21 IM.t10 1.8255
R87 IM.n22 IM.t17 1.8255
R88 IM.n23 IM.t21 1.8255
R89 IM.n24 IM.t8 1.8255
R90 IM.n25 IM.t31 1.8255
R91 IM.n26 IM.t54 1.8255
R92 IM.n27 IM.t57 1.8255
R93 IM.n28 IM.t62 1.8255
R94 IM.n29 IM.t5 1.8255
R95 IM.n30 IM.t24 1.8255
R96 IM.n31 IM.t36 1.8255
R97 IM.n32 IM.t32 1.8255
R98 IM.n33 IM.t60 1.8255
R99 IM.n34 IM.t11 1.8255
R100 IM.n35 IM.t0 1.8255
R101 IM.n36 IM.t40 1.8255
R102 IM.n37 IM.t34 1.8255
R103 IM.n38 IM.t49 1.8255
R104 IM.n39 IM.t23 1.8255
R105 IM.n40 IM.t6 1.8255
R106 IM.n41 IM.t27 1.8255
R107 IM.n42 IM.t43 1.8255
R108 IM.n43 IM.t35 1.8255
R109 IM.n44 IM.t28 1.8255
R110 IM.n45 IM.t20 1.8255
R111 IM.n46 IM.t16 1.8255
R112 IM.n47 IM.t3 1.8255
R113 IM.n48 IM.t13 1.8255
R114 IM.n49 IM.t38 1.8255
R115 IM.n50 IM.t39 1.8255
R116 IM.n51 IM.t25 1.8255
R117 IM.n52 IM.t47 1.8255
R118 IM.n53 IM.t33 1.8255
R119 IM.n54 IM.t22 1.8255
R120 IM.n55 IM.t44 1.8255
R121 IM.n56 IM.t7 1.8255
R122 IM.n57 IM.t58 1.8255
R123 IM.n58 IM.t45 1.8255
R124 IM.n59 IM.t37 1.8255
R125 IM.n60 IM.t41 1.8255
R126 IM.n61 IM.t4 1.8255
R127 IM IM.n64 0.005
R128 IM.n63 IM.n62 0.00360345
R129 VSS.n162 VSS.t27 135.689
R130 VSS.n268 VSS.t2 133.079
R131 VSS.n147 VSS.t62 133.079
R132 VSS.n132 VSS.t12 130.47
R133 VSS.n292 VSS.t41 130.47
R134 VSS.n117 VSS.t0 127.861
R135 VSS.n316 VSS.t5 127.861
R136 VSS.n341 VSS.t11 125.251
R137 VSS.n253 VSS.t20 93.9387
R138 VSS.n156 VSS.t8 93.9387
R139 VSS.n277 VSS.t75 91.3293
R140 VSS.n141 VSS.t3 91.3293
R141 VSS.n126 VSS.t35 88.7199
R142 VSS.n301 VSS.t4 88.7199
R143 VSS.n111 VSS.t14 86.1105
R144 VSS.n325 VSS.t6 86.1105
R145 VSS.n165 VSS.t51 54.7978
R146 VSS.n261 VSS.t77 52.1884
R147 VSS.n150 VSS.t7 52.1884
R148 VSS.n285 VSS.t9 49.579
R149 VSS.n135 VSS.t32 49.579
R150 VSS.n120 VSS.t59 46.9696
R151 VSS.n309 VSS.t38 46.9696
R152 VSS.n336 VSS.t16 44.3602
R153 VSS.n243 VSS.t10 13.0475
R154 VSS.n159 VSS.t25 13.0475
R155 VSS.n270 VSS.t1 10.4381
R156 VSS.n144 VSS.t29 10.4381
R157 VSS.n129 VSS.t22 7.82868
R158 VSS.n294 VSS.t91 7.82868
R159 VSS.n353 VSS.t85 6.37407
R160 VSS.n167 VSS.t121 6.36851
R161 VSS.n24 VSS.n23 6.35417
R162 VSS.n108 VSS.n107 6.35325
R163 VSS.n342 VSS.n341 5.28001
R164 VSS.n114 VSS.t13 5.21929
R165 VSS.n318 VSS.t87 5.21929
R166 VSS.n360 VSS.n359 5.2005
R167 VSS.n333 VSS.n332 5.2005
R168 VSS.n102 VSS.n101 5.2005
R169 VSS.n221 VSS.n218 5.2005
R170 VSS.n168 VSS.n166 5.2005
R171 VSS.n169 VSS.n165 5.2005
R172 VSS.n170 VSS.n164 5.2005
R173 VSS.n171 VSS.n163 5.2005
R174 VSS.n172 VSS.n162 5.2005
R175 VSS.n174 VSS.n159 5.2005
R176 VSS.n175 VSS.n158 5.2005
R177 VSS.n176 VSS.n157 5.2005
R178 VSS.n177 VSS.n156 5.2005
R179 VSS.n178 VSS.n155 5.2005
R180 VSS.n180 VSS.n152 5.2005
R181 VSS.n181 VSS.n151 5.2005
R182 VSS.n182 VSS.n150 5.2005
R183 VSS.n183 VSS.n149 5.2005
R184 VSS.n184 VSS.n148 5.2005
R185 VSS.n185 VSS.n147 5.2005
R186 VSS.n187 VSS.n144 5.2005
R187 VSS.n188 VSS.n143 5.2005
R188 VSS.n189 VSS.n142 5.2005
R189 VSS.n190 VSS.n141 5.2005
R190 VSS.n191 VSS.n140 5.2005
R191 VSS.n193 VSS.n137 5.2005
R192 VSS.n194 VSS.n136 5.2005
R193 VSS.n195 VSS.n135 5.2005
R194 VSS.n196 VSS.n134 5.2005
R195 VSS.n197 VSS.n133 5.2005
R196 VSS.n198 VSS.n132 5.2005
R197 VSS.n200 VSS.n129 5.2005
R198 VSS.n201 VSS.n128 5.2005
R199 VSS.n202 VSS.n127 5.2005
R200 VSS.n203 VSS.n126 5.2005
R201 VSS.n204 VSS.n125 5.2005
R202 VSS.n206 VSS.n122 5.2005
R203 VSS.n207 VSS.n121 5.2005
R204 VSS.n208 VSS.n120 5.2005
R205 VSS.n209 VSS.n119 5.2005
R206 VSS.n210 VSS.n118 5.2005
R207 VSS.n211 VSS.n117 5.2005
R208 VSS.n213 VSS.n114 5.2005
R209 VSS.n214 VSS.n113 5.2005
R210 VSS.n215 VSS.n112 5.2005
R211 VSS.n216 VSS.n111 5.2005
R212 VSS.n246 VSS.n242 5.2005
R213 VSS.n17 VSS.n15 5.2005
R214 VSS.n246 VSS.n241 5.2005
R215 VSS.n246 VSS.n245 5.2005
R216 VSS.n249 VSS.n248 5.2005
R217 VSS.n251 VSS.n250 5.2005
R218 VSS.n254 VSS.n253 5.2005
R219 VSS.n256 VSS.n255 5.2005
R220 VSS.n258 VSS.n257 5.2005
R221 VSS.n260 VSS.n259 5.2005
R222 VSS.n262 VSS.n261 5.2005
R223 VSS.n265 VSS.n264 5.2005
R224 VSS.n267 VSS.n266 5.2005
R225 VSS.n269 VSS.n268 5.2005
R226 VSS.n271 VSS.n270 5.2005
R227 VSS.n273 VSS.n272 5.2005
R228 VSS.n275 VSS.n274 5.2005
R229 VSS.n278 VSS.n277 5.2005
R230 VSS.n280 VSS.n279 5.2005
R231 VSS.n282 VSS.n281 5.2005
R232 VSS.n284 VSS.n283 5.2005
R233 VSS.n286 VSS.n285 5.2005
R234 VSS.n289 VSS.n288 5.2005
R235 VSS.n291 VSS.n290 5.2005
R236 VSS.n293 VSS.n292 5.2005
R237 VSS.n295 VSS.n294 5.2005
R238 VSS.n297 VSS.n296 5.2005
R239 VSS.n299 VSS.n298 5.2005
R240 VSS.n302 VSS.n301 5.2005
R241 VSS.n304 VSS.n303 5.2005
R242 VSS.n306 VSS.n305 5.2005
R243 VSS.n308 VSS.n307 5.2005
R244 VSS.n310 VSS.n309 5.2005
R245 VSS.n313 VSS.n312 5.2005
R246 VSS.n315 VSS.n314 5.2005
R247 VSS.n317 VSS.n316 5.2005
R248 VSS.n319 VSS.n318 5.2005
R249 VSS.n321 VSS.n320 5.2005
R250 VSS.n323 VSS.n322 5.2005
R251 VSS.n326 VSS.n325 5.2005
R252 VSS.n334 VSS.n333 5.2005
R253 VSS.n346 VSS.n335 5.2005
R254 VSS.n345 VSS.n336 5.2005
R255 VSS.n343 VSS.n339 5.2005
R256 VSS.n342 VSS.n340 5.2005
R257 VSS.n221 VSS.n220 4.5005
R258 VSS.n240 VSS.n17 4.5005
R259 VSS.n17 VSS.n16 4.5005
R260 VSS.n240 VSS.n239 4.5005
R261 VSS.n94 VSS.n33 3.62007
R262 VSS.n86 VSS.n37 3.62007
R263 VSS.n79 VSS.n41 3.62007
R264 VSS.n71 VSS.n45 3.62007
R265 VSS.n64 VSS.n49 3.62007
R266 VSS.n56 VSS.n53 3.62007
R267 VSS.n350 VSS.n349 3.62007
R268 VSS.n212 VSS.n116 3.62007
R269 VSS.n205 VSS.n124 3.62007
R270 VSS.n199 VSS.n131 3.62007
R271 VSS.n192 VSS.n139 3.62007
R272 VSS.n186 VSS.n146 3.62007
R273 VSS.n179 VSS.n154 3.62007
R274 VSS.n173 VSS.n161 3.62007
R275 VSS.n356 VSS.n352 3.56724
R276 VSS.n330 VSS.n328 3.56724
R277 VSS.n60 VSS.n51 3.56724
R278 VSS.n67 VSS.n47 3.56724
R279 VSS.n75 VSS.n43 3.56724
R280 VSS.n82 VSS.n39 3.56724
R281 VSS.n90 VSS.n35 3.56724
R282 VSS.n97 VSS.n31 3.56724
R283 VSS.n344 VSS.n338 3.56724
R284 VSS.n324 VSS.n1 3.56724
R285 VSS.n311 VSS.n3 3.56724
R286 VSS.n300 VSS.n5 3.56724
R287 VSS.n287 VSS.n7 3.56724
R288 VSS.n276 VSS.n9 3.56724
R289 VSS.n263 VSS.n11 3.56724
R290 VSS.n252 VSS.n13 3.56724
R291 VSS.n33 VSS.t40 2.7305
R292 VSS.n33 VSS.n32 2.7305
R293 VSS.n37 VSS.t103 2.7305
R294 VSS.n37 VSS.n36 2.7305
R295 VSS.n41 VSS.t23 2.7305
R296 VSS.n41 VSS.n40 2.7305
R297 VSS.n45 VSS.t42 2.7305
R298 VSS.n45 VSS.n44 2.7305
R299 VSS.n49 VSS.t30 2.7305
R300 VSS.n49 VSS.n48 2.7305
R301 VSS.n53 VSS.t90 2.7305
R302 VSS.n53 VSS.n52 2.7305
R303 VSS.n349 VSS.t34 2.7305
R304 VSS.n349 VSS.n348 2.7305
R305 VSS.n352 VSS.t66 2.7305
R306 VSS.n352 VSS.n351 2.7305
R307 VSS.n328 VSS.t50 2.7305
R308 VSS.n328 VSS.n327 2.7305
R309 VSS.n51 VSS.t84 2.7305
R310 VSS.n51 VSS.n50 2.7305
R311 VSS.n47 VSS.t122 2.7305
R312 VSS.n47 VSS.n46 2.7305
R313 VSS.n43 VSS.t68 2.7305
R314 VSS.n43 VSS.n42 2.7305
R315 VSS.n39 VSS.t86 2.7305
R316 VSS.n39 VSS.n38 2.7305
R317 VSS.n35 VSS.t127 2.7305
R318 VSS.n35 VSS.n34 2.7305
R319 VSS.n31 VSS.t67 2.7305
R320 VSS.n31 VSS.n30 2.7305
R321 VSS.n116 VSS.t19 2.7305
R322 VSS.n116 VSS.n115 2.7305
R323 VSS.n124 VSS.t69 2.7305
R324 VSS.n124 VSS.n123 2.7305
R325 VSS.n131 VSS.t83 2.7305
R326 VSS.n131 VSS.n130 2.7305
R327 VSS.n139 VSS.t89 2.7305
R328 VSS.n139 VSS.n138 2.7305
R329 VSS.n146 VSS.t65 2.7305
R330 VSS.n146 VSS.n145 2.7305
R331 VSS.n154 VSS.t70 2.7305
R332 VSS.n154 VSS.n153 2.7305
R333 VSS.n161 VSS.t26 2.7305
R334 VSS.n161 VSS.n160 2.7305
R335 VSS.n338 VSS.t17 2.7305
R336 VSS.n338 VSS.n337 2.7305
R337 VSS.n1 VSS.t114 2.7305
R338 VSS.n1 VSS.n0 2.7305
R339 VSS.n3 VSS.t39 2.7305
R340 VSS.n3 VSS.n2 2.7305
R341 VSS.n5 VSS.t80 2.7305
R342 VSS.n5 VSS.n4 2.7305
R343 VSS.n7 VSS.t18 2.7305
R344 VSS.n7 VSS.n6 2.7305
R345 VSS.n9 VSS.t36 2.7305
R346 VSS.n9 VSS.n8 2.7305
R347 VSS.n11 VSS.t78 2.7305
R348 VSS.n11 VSS.n10 2.7305
R349 VSS.n13 VSS.t15 2.7305
R350 VSS.n13 VSS.n12 2.7305
R351 VSS.n223 VSS.n222 2.60175
R352 VSS.n362 VSS.n361 2.6005
R353 VSS.n361 VSS.n360 2.6005
R354 VSS.n244 VSS.n243 2.39249
R355 VSS.n102 VSS.n29 2.39249
R356 VSS.n228 VSS.n108 2.2505
R357 VSS.n227 VSS.n226 2.2505
R358 VSS.n234 VSS.n24 2.2505
R359 VSS.n238 VSS.n237 2.25028
R360 VSS.n236 VSS.n235 2.2497
R361 VSS.n233 VSS.n106 2.24958
R362 VSS.n221 VSS.n219 1.92278
R363 VSS.n361 VSS.n347 1.63262
R364 VSS.n26 VSS.n25 1.56009
R365 VSS.n15 VSS.n14 1.3052
R366 VSS.n28 VSS.n27 1.23366
R367 VSS.n229 VSS.n228 1.01937
R368 VSS.n235 VSS.n234 0.514333
R369 VSS.n222 VSS.n221 0.424592
R370 VSS.n245 VSS.n244 0.41801
R371 VSS.n29 VSS.n28 0.41801
R372 VSS.n29 VSS.n26 0.41801
R373 VSS.n216 VSS.n215 0.0800053
R374 VSS.n215 VSS.n214 0.0800053
R375 VSS.n214 VSS.n213 0.0800053
R376 VSS.n211 VSS.n210 0.0800053
R377 VSS.n210 VSS.n209 0.0800053
R378 VSS.n209 VSS.n208 0.0800053
R379 VSS.n208 VSS.n207 0.0800053
R380 VSS.n207 VSS.n206 0.0800053
R381 VSS.n204 VSS.n203 0.0800053
R382 VSS.n203 VSS.n202 0.0800053
R383 VSS.n202 VSS.n201 0.0800053
R384 VSS.n201 VSS.n200 0.0800053
R385 VSS.n198 VSS.n197 0.0800053
R386 VSS.n197 VSS.n196 0.0800053
R387 VSS.n196 VSS.n195 0.0800053
R388 VSS.n195 VSS.n194 0.0800053
R389 VSS.n194 VSS.n193 0.0800053
R390 VSS.n191 VSS.n190 0.0800053
R391 VSS.n190 VSS.n189 0.0800053
R392 VSS.n189 VSS.n188 0.0800053
R393 VSS.n188 VSS.n187 0.0800053
R394 VSS.n185 VSS.n184 0.0800053
R395 VSS.n184 VSS.n183 0.0800053
R396 VSS.n183 VSS.n182 0.0800053
R397 VSS.n182 VSS.n181 0.0800053
R398 VSS.n181 VSS.n180 0.0800053
R399 VSS.n178 VSS.n177 0.0800053
R400 VSS.n177 VSS.n176 0.0800053
R401 VSS.n176 VSS.n175 0.0800053
R402 VSS.n175 VSS.n174 0.0800053
R403 VSS.n172 VSS.n171 0.0800053
R404 VSS.n171 VSS.n170 0.0800053
R405 VSS.n170 VSS.n169 0.0800053
R406 VSS.n169 VSS.n168 0.0800053
R407 VSS.n168 VSS.n167 0.0800053
R408 VSS.n251 VSS.n249 0.0800053
R409 VSS.n256 VSS.n254 0.0800053
R410 VSS.n258 VSS.n256 0.0800053
R411 VSS.n260 VSS.n258 0.0800053
R412 VSS.n262 VSS.n260 0.0800053
R413 VSS.n267 VSS.n265 0.0800053
R414 VSS.n269 VSS.n267 0.0800053
R415 VSS.n271 VSS.n269 0.0800053
R416 VSS.n273 VSS.n271 0.0800053
R417 VSS.n275 VSS.n273 0.0800053
R418 VSS.n280 VSS.n278 0.0800053
R419 VSS.n282 VSS.n280 0.0800053
R420 VSS.n284 VSS.n282 0.0800053
R421 VSS.n286 VSS.n284 0.0800053
R422 VSS.n291 VSS.n289 0.0800053
R423 VSS.n293 VSS.n291 0.0800053
R424 VSS.n295 VSS.n293 0.0800053
R425 VSS.n297 VSS.n295 0.0800053
R426 VSS.n299 VSS.n297 0.0800053
R427 VSS.n304 VSS.n302 0.0800053
R428 VSS.n306 VSS.n304 0.0800053
R429 VSS.n308 VSS.n306 0.0800053
R430 VSS.n310 VSS.n308 0.0800053
R431 VSS.n315 VSS.n313 0.0800053
R432 VSS.n317 VSS.n315 0.0800053
R433 VSS.n319 VSS.n317 0.0800053
R434 VSS.n321 VSS.n319 0.0800053
R435 VSS.n323 VSS.n321 0.0800053
R436 VSS.n334 VSS.n326 0.0800053
R437 VSS.n362 VSS.n346 0.0800053
R438 VSS.n346 VSS.n345 0.0800053
R439 VSS.n343 VSS.n342 0.0800053
R440 VSS.n99 VSS.n98 0.0794474
R441 VSS.n96 VSS.n95 0.0794474
R442 VSS.n93 VSS.n92 0.0794474
R443 VSS.n92 VSS.n91 0.0794474
R444 VSS.n89 VSS.n88 0.0794474
R445 VSS.n88 VSS.n87 0.0794474
R446 VSS.n85 VSS.n84 0.0794474
R447 VSS.n84 VSS.n83 0.0794474
R448 VSS.n81 VSS.n80 0.0794474
R449 VSS.n78 VSS.n77 0.0794474
R450 VSS.n77 VSS.n76 0.0794474
R451 VSS.n74 VSS.n73 0.0794474
R452 VSS.n73 VSS.n72 0.0794474
R453 VSS.n70 VSS.n69 0.0794474
R454 VSS.n69 VSS.n68 0.0794474
R455 VSS.n66 VSS.n65 0.0794474
R456 VSS.n63 VSS.n62 0.0794474
R457 VSS.n62 VSS.n61 0.0794474
R458 VSS.n59 VSS.n58 0.0794474
R459 VSS.n58 VSS.n57 0.0794474
R460 VSS.n55 VSS.n54 0.0794474
R461 VSS.n332 VSS.n331 0.0794474
R462 VSS.n359 VSS.n358 0.0794474
R463 VSS.n358 VSS.n357 0.0794474
R464 VSS.n355 VSS.n354 0.0794474
R465 VSS.n354 VSS.n353 0.0794474
R466 VSS.n254 VSS.n252 0.0780972
R467 VSS.n97 VSS.n96 0.0775526
R468 VSS.n278 VSS.n276 0.0774611
R469 VSS.n217 VSS.n216 0.0771431
R470 VSS.n82 VSS.n81 0.0769211
R471 VSS.n302 VSS.n300 0.0768251
R472 VSS.n67 VSS.n66 0.0762895
R473 VSS.n326 VSS.n324 0.076189
R474 VSS.n331 VSS.n330 0.0756579
R475 VSS.n249 VSS.n247 0.0739629
R476 VSS.n100 VSS.n99 0.0734474
R477 VSS VSS.n334 0.0711007
R478 VSS.n205 VSS.n204 0.0634682
R479 VSS.n65 VSS.n64 0.0630263
R480 VSS.n192 VSS.n191 0.0628322
R481 VSS.n80 VSS.n79 0.0623947
R482 VSS.n179 VSS.n178 0.0621961
R483 VSS.n95 VSS.n94 0.0617632
R484 VSS.n174 VSS.n173 0.0583799
R485 VSS.n187 VSS.n186 0.0577438
R486 VSS.n86 VSS.n85 0.0573421
R487 VSS.n200 VSS.n199 0.0571078
R488 VSS.n71 VSS.n70 0.0567105
R489 VSS.n213 VSS.n212 0.0564717
R490 VSS.n56 VSS.n55 0.056079
R491 VSS.n227 VSS.n110 0.0517376
R492 VSS.n345 VSS.n344 0.0443869
R493 VSS.n357 VSS.n356 0.0440789
R494 VSS.n311 VSS.n310 0.0437509
R495 VSS.n61 VSS.n60 0.0434474
R496 VSS.n287 VSS.n286 0.0431148
R497 VSS.n76 VSS.n75 0.0428158
R498 VSS.n263 VSS.n262 0.0424788
R499 VSS.n91 VSS.n90 0.0421842
R500 VSS.n265 VSS.n263 0.0380265
R501 VSS.n90 VSS.n89 0.0377632
R502 VSS.n289 VSS.n287 0.0373905
R503 VSS.n75 VSS.n74 0.0371316
R504 VSS.n313 VSS.n311 0.0367544
R505 VSS.n60 VSS.n59 0.0365
R506 VSS.n344 VSS.n343 0.0361184
R507 VSS.n356 VSS.n355 0.0358684
R508 VSS.n19 VSS.n18 0.0284859
R509 VSS.n232 VSS.n231 0.0249038
R510 VSS.n233 VSS.n232 0.0249038
R511 VSS.n212 VSS.n211 0.0240336
R512 VSS.n57 VSS.n56 0.0238684
R513 VSS.n199 VSS.n198 0.0233975
R514 VSS.n72 VSS.n71 0.0232368
R515 VSS.n186 VSS.n185 0.0227615
R516 VSS.n87 VSS.n86 0.0226053
R517 VSS.n173 VSS.n172 0.0221254
R518 VSS.n224 VSS.n223 0.0205353
R519 VSS.n180 VSS.n179 0.0183092
R520 VSS.n94 VSS.n93 0.0181842
R521 VSS.n193 VSS.n192 0.0176731
R522 VSS.n79 VSS.n78 0.0175526
R523 VSS.n246 VSS.n240 0.0173551
R524 VSS.n103 VSS.n102 0.0172368
R525 VSS.n206 VSS.n205 0.0170371
R526 VSS.n64 VSS.n63 0.0169211
R527 VSS.n359 VSS.n350 0.0162895
R528 VSS VSS.n362 0.00940459
R529 VSS.n226 VSS.n224 0.00686042
R530 VSS.n22 VSS.n21 0.00662565
R531 VSS.n231 VSS.n230 0.00662565
R532 VSS.n247 VSS.n246 0.0065424
R533 VSS.n102 VSS.n100 0.0065
R534 VSS.n236 VSS.n20 0.00622438
R535 VSS.n235 VSS.n22 0.00547495
R536 VSS.n230 VSS.n229 0.00547495
R537 VSS.n324 VSS.n323 0.00431625
R538 VSS.n330 VSS.n329 0.00428947
R539 VSS.n106 VSS.n105 0.0041561
R540 VSS.n106 VSS.n104 0.00384031
R541 VSS.n300 VSS.n299 0.00368021
R542 VSS.n68 VSS.n67 0.00365789
R543 VSS.n223 VSS.n217 0.00336219
R544 VSS.n104 VSS.n103 0.00334211
R545 VSS.n276 VSS.n275 0.00304417
R546 VSS.n83 VSS.n82 0.00302632
R547 VSS.n238 VSS.n236 0.00243064
R548 VSS.n240 VSS.n238 0.00243064
R549 VSS.n252 VSS.n251 0.00240813
R550 VSS.n98 VSS.n97 0.00239474
R551 VSS.n110 VSS.n109 0.00228218
R552 VSS.n226 VSS.n225 0.00227173
R553 VSS.n234 VSS.n233 0.000971204
R554 VSS.n228 VSS.n227 0.000945545
R555 VSS.n20 VSS.n19 0.000818021
R556 SD.n281 SD.n20 3.42994
R557 SD.n209 SD.n160 3.4191
R558 SD.n196 SD.n167 3.41548
R559 SD.n181 SD.n180 3.41548
R560 SD.n289 SD.n1 3.00983
R561 SD.n202 SD.n165 3.00364
R562 SD.n223 SD.n127 3.00306
R563 SD.n231 SD.n122 2.99802
R564 SD.n243 SD.n96 2.997
R565 SD.n217 SD.n129 2.99431
R566 SD.n193 SD.n172 2.99196
R567 SD.n254 SD.n86 2.99039
R568 SD.n251 SD.n91 2.99018
R569 SD.n278 SD.n32 2.98846
R570 SD.n260 SD.n84 2.98001
R571 SD.n267 SD.n55 2.97893
R572 SD.n30 SD.n29 2.93962
R573 SD.n158 SD.n157 2.93841
R574 SD.n170 SD.n169 2.93801
R575 SD.n178 SD.n177 2.93801
R576 SD.n283 SD.n282 2.90232
R577 SD.n24 SD.n23 2.90232
R578 SD.n184 SD.n183 2.90222
R579 SD.n137 SD.n136 2.90222
R580 SD.n274 SD.n273 2.90218
R581 SD.n38 SD.n37 2.90218
R582 SD.n263 SD.n262 2.90214
R583 SD.n84 SD.n83 2.90214
R584 SD.n46 SD.n45 2.90214
R585 SD.n81 SD.n80 2.90214
R586 SD.n55 SD.n54 2.87834
R587 SD.n52 SD.n51 2.87834
R588 SD.n270 SD.n269 2.87832
R589 SD.n34 SD.n33 2.87832
R590 SD.n32 SD.n31 2.85397
R591 SD.n43 SD.n42 2.85397
R592 SD.n86 SD.t90 2.7305
R593 SD.n86 SD.n85 2.7305
R594 SD.n256 SD.t71 2.7305
R595 SD.n256 SD.n255 2.7305
R596 SD.n91 SD.t38 2.7305
R597 SD.n91 SD.n90 2.7305
R598 SD.n248 SD.t16 2.7305
R599 SD.n248 SD.n247 2.7305
R600 SD.n240 SD.t79 2.7305
R601 SD.n240 SD.n239 2.7305
R602 SD.n234 SD.t93 2.7305
R603 SD.n234 SD.n233 2.7305
R604 SD.n129 SD.t50 2.7305
R605 SD.n129 SD.n128 2.7305
R606 SD.n219 SD.t84 2.7305
R607 SD.n219 SD.n218 2.7305
R608 SD.n213 SD.t68 2.7305
R609 SD.n213 SD.n212 2.7305
R610 SD.n205 SD.t96 2.7305
R611 SD.n205 SD.n204 2.7305
R612 SD.n167 SD.t0 2.7305
R613 SD.n167 SD.n166 2.7305
R614 SD.n198 SD.t32 2.7305
R615 SD.n198 SD.n197 2.7305
R616 SD.n172 SD.t21 2.7305
R617 SD.n172 SD.n171 2.7305
R618 SD.n190 SD.t115 2.7305
R619 SD.n190 SD.n189 2.7305
R620 SD.n227 SD.t62 2.7305
R621 SD.n227 SD.n226 2.7305
R622 SD.n20 SD.t85 2.7305
R623 SD.n20 SD.n19 2.7305
R624 SD.n180 SD.t11 2.7305
R625 SD.n180 SD.n179 2.7305
R626 SD.n165 SD.t78 2.7305
R627 SD.n165 SD.n164 2.7305
R628 SD.n160 SD.t7 2.7305
R629 SD.n160 SD.n159 2.7305
R630 SD.n127 SD.t81 2.7305
R631 SD.n127 SD.n126 2.7305
R632 SD.n122 SD.t25 2.7305
R633 SD.n122 SD.n121 2.7305
R634 SD.n96 SD.t101 2.7305
R635 SD.n96 SD.n95 2.7305
R636 SD.n1 SD.t75 2.7305
R637 SD.n1 SD.n0 2.7305
R638 SD.n8 SD.t39 2.7305
R639 SD.n8 SD.n7 2.7305
R640 SD.n88 SD.t82 2.7305
R641 SD.n88 SD.n87 2.7305
R642 SD.n75 SD.t41 2.7305
R643 SD.n75 SD.n74 2.7305
R644 SD.n93 SD.t67 2.7305
R645 SD.n93 SD.n92 2.7305
R646 SD.n57 SD.t4 2.7305
R647 SD.n57 SD.n56 2.7305
R648 SD.n60 SD.t64 2.7305
R649 SD.n60 SD.n59 2.7305
R650 SD.n63 SD.t88 2.7305
R651 SD.n63 SD.n62 2.7305
R652 SD.n131 SD.t74 2.7305
R653 SD.n131 SD.n130 2.7305
R654 SD.n112 SD.t125 2.7305
R655 SD.n112 SD.n111 2.7305
R656 SD.n106 SD.t31 2.7305
R657 SD.n106 SD.n105 2.7305
R658 SD.n151 SD.t121 2.7305
R659 SD.n151 SD.n150 2.7305
R660 SD.n169 SD.t92 2.7305
R661 SD.n169 SD.n168 2.7305
R662 SD.n145 SD.t69 2.7305
R663 SD.n145 SD.n144 2.7305
R664 SD.n174 SD.t48 2.7305
R665 SD.n174 SD.n173 2.7305
R666 SD.n134 SD.t103 2.7305
R667 SD.n134 SD.n133 2.7305
R668 SD.n103 SD.t37 2.7305
R669 SD.n103 SD.n102 2.7305
R670 SD.n29 SD.t122 2.7305
R671 SD.n29 SD.n28 2.7305
R672 SD.n12 SD.t97 2.7305
R673 SD.n12 SD.n11 2.7305
R674 SD.n177 SD.t102 2.7305
R675 SD.n177 SD.n176 2.7305
R676 SD.n162 SD.t40 2.7305
R677 SD.n162 SD.n161 2.7305
R678 SD.n157 SD.t1 2.7305
R679 SD.n157 SD.n156 2.7305
R680 SD.n124 SD.t13 2.7305
R681 SD.n124 SD.n123 2.7305
R682 SD.n101 SD.t52 2.7305
R683 SD.n101 SD.n100 2.7305
R684 SD.n98 SD.t113 2.7305
R685 SD.n98 SD.n97 2.7305
R686 SD.n4 SD.t118 2.7305
R687 SD.n4 SD.n3 2.7305
R688 SD.n17 SD.n8 2.56388
R689 SD.n163 SD.n162 2.5636
R690 SD.n89 SD.n88 2.5632
R691 SD.n94 SD.n93 2.5632
R692 SD.n125 SD.n124 2.56319
R693 SD.n120 SD.n101 2.56301
R694 SD.n175 SD.n174 2.56295
R695 SD.n99 SD.n98 2.5627
R696 SD.n132 SD.n131 2.56252
R697 SD.n82 SD.n81 2.51058
R698 SD.n53 SD.n52 2.50789
R699 SD.n44 SD.n43 2.50617
R700 SD.n138 SD.n137 2.50572
R701 SD.n32 SD.t49 2.46898
R702 SD.n43 SD.t73 2.46898
R703 SD.n270 SD.t59 2.4382
R704 SD.n34 SD.t58 2.4382
R705 SD.n55 SD.t104 2.43819
R706 SD.n52 SD.t98 2.43819
R707 SD.n263 SD.t8 2.40702
R708 SD.n84 SD.t70 2.40702
R709 SD.n46 SD.t99 2.40702
R710 SD.n81 SD.t33 2.40702
R711 SD.n274 SD.t108 2.40698
R712 SD.n38 SD.t6 2.40698
R713 SD.n184 SD.t61 2.40695
R714 SD.n137 SD.t65 2.40695
R715 SD.n283 SD.t23 2.40687
R716 SD.n24 SD.t35 2.40687
R717 SD.n14 SD.n13 2.25075
R718 SD.n250 SD.n249 2.25075
R719 SD.n288 SD.n6 2.25075
R720 SD.n192 SD.n191 2.25049
R721 SD.n242 SD.n241 2.25049
R722 SD.n40 SD.n39 2.24974
R723 SD.n276 SD.n275 2.24974
R724 SD.n26 SD.n25 2.24545
R725 SD.n36 SD.n35 2.24545
R726 SD.n285 SD.n284 2.24545
R727 SD.n272 SD.n271 2.24545
R728 SD.n48 SD.n47 2.2452
R729 SD.n186 SD.n185 2.2452
R730 SD.n265 SD.n264 2.2452
R731 SD.n153 SD.n152 2.24495
R732 SD.n65 SD.n64 2.24495
R733 SD.n207 SD.n206 2.24495
R734 SD.n236 SD.n235 2.24495
R735 SD.n229 SD.n228 2.2447
R736 SD.n215 SD.n214 2.2447
R737 SD.n117 SD.n104 1.49529
R738 SD.n147 SD.n146 1.49529
R739 SD.n69 SD.n58 1.49529
R740 SD.n200 SD.n199 1.49529
R741 SD.n139 SD.n135 1.49529
R742 SD.n66 SD.n61 1.49529
R743 SD.n114 SD.n113 1.49518
R744 SD.n77 SD.n76 1.49518
R745 SD.n221 SD.n220 1.49518
R746 SD.n258 SD.n257 1.49518
R747 SD.n108 SD.n107 1.49507
R748 SD.n13 SD.n12 1.4398
R749 SD.n5 SD.n4 1.43954
R750 SD.n191 SD.n190 1.439
R751 SD.n228 SD.n227 1.439
R752 SD.n135 SD.n134 1.439
R753 SD.n104 SD.n103 1.439
R754 SD.n220 SD.n219 1.43841
R755 SD.n113 SD.n112 1.43841
R756 SD.n206 SD.n205 1.43819
R757 SD.n199 SD.n198 1.43819
R758 SD.n152 SD.n151 1.43819
R759 SD.n146 SD.n145 1.43819
R760 SD.n241 SD.n240 1.43801
R761 SD.n61 SD.n60 1.43801
R762 SD.n257 SD.n256 1.43752
R763 SD.n249 SD.n248 1.43752
R764 SD.n235 SD.n234 1.43752
R765 SD.n76 SD.n75 1.43752
R766 SD.n58 SD.n57 1.43752
R767 SD.n64 SD.n63 1.43752
R768 SD.n214 SD.n213 1.43734
R769 SD.n107 SD.n106 1.43734
R770 SD.n225 SD.n125 1.20162
R771 SD.n188 SD.n175 1.1255
R772 SD.n254 SD.n89 1.12404
R773 SD.n246 SD.n94 1.12404
R774 SD.n268 SD.n53 1.12287
R775 SD.n261 SD.n82 1.12272
R776 SD.n217 SD.n132 1.12097
R777 SD.n238 SD.n99 1.11849
R778 SD.n182 SD.n178 1.11776
R779 SD.n196 SD.n170 1.11732
R780 SD.n232 SD.n120 1.116
R781 SD.n18 SD.n17 1.11279
R782 SD.n203 SD.n163 1.1125
R783 SD.n211 SD.n158 1.11235
R784 SD.n277 SD.n44 1.11206
R785 SD.n281 SD.n30 1.10709
R786 SD.n25 SD.n24 1.01162
R787 SD.n284 SD.n283 1.01162
R788 SD.n185 SD.n184 1.01104
R789 SD.n39 SD.n38 1.0108
R790 SD.n275 SD.n274 1.0108
R791 SD.n47 SD.n46 1.01058
R792 SD.n264 SD.n263 1.01058
R793 SD.n271 SD.n270 1.00825
R794 SD.n35 SD.n34 1.00825
R795 SD.n78 SD.n77 0.68891
R796 SD.n259 SD.n258 0.68891
R797 SD.n40 SD.n36 0.681527
R798 SD.n276 SD.n272 0.681527
R799 SD.n49 SD.n48 0.681026
R800 SD.n266 SD.n265 0.681026
R801 SD.n148 SD.n147 0.677238
R802 SD.n201 SD.n200 0.677238
R803 SD.n118 SD.n117 0.676563
R804 SD.n139 SD.n138 0.676193
R805 SD.n66 SD.n65 0.672859
R806 SD.n230 SD.n229 0.671376
R807 SD.n22 SD.n21 0.667916
R808 SD.n280 SD.n279 0.667916
R809 SD.n115 SD.n114 0.662617
R810 SD.n222 SD.n221 0.662617
R811 SD.n69 SD.n68 0.662613
R812 SD.n109 SD.n108 0.662274
R813 SD.n154 SD.n153 0.657259
R814 SD.n208 SD.n207 0.657259
R815 SD.n216 SD.n215 0.656751
R816 SD.n237 SD.n236 0.655237
R817 SD.n286 SD.n285 0.65322
R818 SD.n187 SD.n186 0.652712
R819 SD.n72 SD.n71 0.645669
R820 SD.n253 SD.n252 0.645669
R821 SD.n142 SD.n141 0.644657
R822 SD.n195 SD.n194 0.644657
R823 SD.n245 SD.n244 0.644657
R824 SD.n287 SD.n18 0.6305
R825 SD.n30 SD.n27 0.490825
R826 SD.n17 SD.n16 0.484396
R827 SD.n44 SD.n41 0.482789
R828 SD.n158 SD.n155 0.481182
R829 SD.n120 SD.n119 0.477968
R830 SD.n53 SD.n50 0.471539
R831 SD.n82 SD.n79 0.469932
R832 SD.n141 SD.n140 0.0257809
R833 SD.n143 SD.n142 0.0257809
R834 SD.n110 SD.n109 0.0257809
R835 SD.n71 SD.n70 0.0257809
R836 SD.n73 SD.n72 0.0257809
R837 SD.n194 SD.n193 0.0257809
R838 SD.n196 SD.n195 0.0257809
R839 SD.n217 SD.n216 0.0257809
R840 SD.n246 SD.n245 0.0257809
R841 SD.n252 SD.n251 0.0257809
R842 SD.n254 SD.n253 0.0257809
R843 SD.n68 SD.n67 0.0247697
R844 SD.n188 SD.n187 0.0247697
R845 SD.n238 SD.n237 0.0247697
R846 SD.n244 SD.n243 0.0247697
R847 SD.n155 SD.n154 0.0237584
R848 SD.n10 SD.n9 0.0237584
R849 SD.n209 SD.n208 0.0237584
R850 SD.n287 SD.n286 0.0237584
R851 SD.n116 SD.n115 0.021736
R852 SD.n16 SD.n15 0.021736
R853 SD.n223 SD.n222 0.021736
R854 SD.n279 SD.n278 0.021736
R855 SD.n149 SD.n148 0.0151247
R856 SD.n202 SD.n201 0.0151247
R857 SD.n117 SD.n116 0.0144442
R858 SD.n153 SD.n149 0.0141134
R859 SD.n119 SD.n118 0.0141134
R860 SD.n231 SD.n230 0.0141134
R861 SD.n215 SD.n211 0.013605
R862 SD.n229 SD.n225 0.013605
R863 SD.n207 SD.n203 0.0131022
R864 SD.n236 SD.n232 0.0131022
R865 SD SD.n290 0.0126348
R866 SD.n186 SD.n182 0.0125992
R867 SD.n265 SD.n261 0.0125992
R868 SD.n27 SD.n26 0.0120962
R869 SD.n272 SD.n268 0.0120962
R870 SD.n285 SD.n281 0.0120962
R871 SD.n67 SD.n66 0.0120831
R872 SD.n140 SD.n139 0.0110719
R873 SD.n147 SD.n143 0.0107344
R874 SD.n70 SD.n69 0.0107344
R875 SD.n200 SD.n196 0.0107344
R876 SD.n114 SD.n110 0.00973004
R877 SD.n77 SD.n73 0.00973004
R878 SD.n221 SD.n217 0.00973004
R879 SD.n258 SD.n254 0.00973004
R880 SD SD.n289 0.00960112
R881 SD.n27 SD.n22 0.00656742
R882 SD.n281 SD.n280 0.00656742
R883 SD.n16 SD.n14 0.0055505
R884 SD.n289 SD.n288 0.0055505
R885 SD.n41 SD.n40 0.00554914
R886 SD.n5 SD.n2 0.00461062
R887 SD.n79 SD.n78 0.00454494
R888 SD.n50 SD.n49 0.00454494
R889 SD.n182 SD.n181 0.00454494
R890 SD.n224 SD.n223 0.00454494
R891 SD.n260 SD.n259 0.00454494
R892 SD.n267 SD.n266 0.00454494
R893 SD.n14 SD.n10 0.00352803
R894 SD.n288 SD.n287 0.00352803
R895 SD.n277 SD.n276 0.00352667
R896 SD.n243 SD.n242 0.00302224
R897 SD.n211 SD.n210 0.00252247
R898 SD.n232 SD.n231 0.00252247
R899 SD.n268 SD.n267 0.00252247
R900 SD.n278 SD.n277 0.00252247
R901 SD.n6 SD.n5 0.00206204
R902 SD.n192 SD.n188 0.00201101
R903 SD.n242 SD.n238 0.00201101
R904 SD.n193 SD.n192 0.00201101
R905 SD.n203 SD.n202 0.00151124
R906 SD.n210 SD.n209 0.00151124
R907 SD.n225 SD.n224 0.00151124
R908 SD.n261 SD.n260 0.00151124
R909 SD.n250 SD.n246 0.00150556
R910 SD.n251 SD.n250 0.00150556
R911 IM_T.n52 IM_T.n51 156.624
R912 IM_T.n54 IM_T.n53 156.624
R913 IM_T.n56 IM_T.n55 156.624
R914 IM_T.n58 IM_T.n57 156.624
R915 IM_T.n60 IM_T.n59 156.624
R916 IM_T.n62 IM_T.n61 156.624
R917 IM_T.n64 IM_T.n63 156.624
R918 IM_T.n17 IM_T.n16 156.624
R919 IM_T.n19 IM_T.n18 156.624
R920 IM_T.n21 IM_T.n20 156.624
R921 IM_T.n23 IM_T.n22 156.624
R922 IM_T.n25 IM_T.n24 156.624
R923 IM_T.n27 IM_T.n26 156.624
R924 IM_T.n29 IM_T.n28 156.624
R925 IM_T.n50 IM_T.t2 156.208
R926 IM_T.n15 IM_T.t46 156.208
R927 IM_T.n1 IM_T.n0 156.143
R928 IM_T.n3 IM_T.n2 156.143
R929 IM_T.n5 IM_T.n4 156.143
R930 IM_T.n7 IM_T.n6 156.143
R931 IM_T.n9 IM_T.n8 156.143
R932 IM_T.n11 IM_T.n10 156.143
R933 IM_T.n13 IM_T.n12 156.143
R934 IM_T.n31 IM_T.n30 156.143
R935 IM_T.n33 IM_T.n32 156.143
R936 IM_T.n35 IM_T.n34 156.143
R937 IM_T.n37 IM_T.n36 156.143
R938 IM_T.n39 IM_T.n38 156.143
R939 IM_T.n41 IM_T.n40 156.143
R940 IM_T.n43 IM_T.n42 156.143
R941 IM_T.n45 IM_T.n44 110.537
R942 IM_T.n46 IM_T.n14 109.225
R943 IM_T.n45 IM_T.n29 42.8895
R944 IM_T.n65 IM_T.n64 33.8925
R945 IM_T.n51 IM_T.n50 31.0633
R946 IM_T.n53 IM_T.n52 31.0633
R947 IM_T.n55 IM_T.n54 31.0633
R948 IM_T.n57 IM_T.n56 31.0633
R949 IM_T.n59 IM_T.n58 31.0633
R950 IM_T.n61 IM_T.n60 31.0633
R951 IM_T.n63 IM_T.n62 31.0633
R952 IM_T.n16 IM_T.n15 31.0633
R953 IM_T.n18 IM_T.n17 31.0633
R954 IM_T.n20 IM_T.n19 31.0633
R955 IM_T.n22 IM_T.n21 31.0633
R956 IM_T.n24 IM_T.n23 31.0633
R957 IM_T.n26 IM_T.n25 31.0633
R958 IM_T.n28 IM_T.n27 31.0633
R959 IM_T.n0 IM_T.t21 30.5914
R960 IM_T.n30 IM_T.t34 30.5914
R961 IM_T.n2 IM_T.n1 30.5831
R962 IM_T.n4 IM_T.n3 30.5831
R963 IM_T.n6 IM_T.n5 30.5831
R964 IM_T.n8 IM_T.n7 30.5831
R965 IM_T.n10 IM_T.n9 30.5831
R966 IM_T.n12 IM_T.n11 30.5831
R967 IM_T.n14 IM_T.n13 30.5831
R968 IM_T.n32 IM_T.n31 30.5831
R969 IM_T.n34 IM_T.n33 30.5831
R970 IM_T.n36 IM_T.n35 30.5831
R971 IM_T.n38 IM_T.n37 30.5831
R972 IM_T.n40 IM_T.n39 30.5831
R973 IM_T.n42 IM_T.n41 30.5831
R974 IM_T.n44 IM_T.n43 30.5831
R975 IM_T.n66 IM_T.n49 4.52761
R976 IM_T.n66 IM_T.n65 2.25833
R977 IM_T.n48 IM_T.n47 2.24388
R978 IM_T.n50 IM_T.t38 1.8255
R979 IM_T.n51 IM_T.t35 1.8255
R980 IM_T.n52 IM_T.t62 1.8255
R981 IM_T.n53 IM_T.t59 1.8255
R982 IM_T.n54 IM_T.t30 1.8255
R983 IM_T.n55 IM_T.t1 1.8255
R984 IM_T.n56 IM_T.t37 1.8255
R985 IM_T.n57 IM_T.t51 1.8255
R986 IM_T.n58 IM_T.t45 1.8255
R987 IM_T.n59 IM_T.t56 1.8255
R988 IM_T.n60 IM_T.t63 1.8255
R989 IM_T.n61 IM_T.t3 1.8255
R990 IM_T.n62 IM_T.t39 1.8255
R991 IM_T.n63 IM_T.t44 1.8255
R992 IM_T.n64 IM_T.t7 1.8255
R993 IM_T.n0 IM_T.t16 1.8255
R994 IM_T.n1 IM_T.t50 1.8255
R995 IM_T.n2 IM_T.t24 1.8255
R996 IM_T.n3 IM_T.t4 1.8255
R997 IM_T.n4 IM_T.t53 1.8255
R998 IM_T.n5 IM_T.t20 1.8255
R999 IM_T.n6 IM_T.t11 1.8255
R1000 IM_T.n7 IM_T.t52 1.8255
R1001 IM_T.n8 IM_T.t60 1.8255
R1002 IM_T.n9 IM_T.t8 1.8255
R1003 IM_T.n10 IM_T.t29 1.8255
R1004 IM_T.n11 IM_T.t28 1.8255
R1005 IM_T.n12 IM_T.t54 1.8255
R1006 IM_T.n13 IM_T.t22 1.8255
R1007 IM_T.n14 IM_T.t25 1.8255
R1008 IM_T.n15 IM_T.t12 1.8255
R1009 IM_T.n16 IM_T.t6 1.8255
R1010 IM_T.n17 IM_T.t41 1.8255
R1011 IM_T.n18 IM_T.t36 1.8255
R1012 IM_T.n19 IM_T.t0 1.8255
R1013 IM_T.n20 IM_T.t47 1.8255
R1014 IM_T.n21 IM_T.t10 1.8255
R1015 IM_T.n22 IM_T.t23 1.8255
R1016 IM_T.n23 IM_T.t14 1.8255
R1017 IM_T.n24 IM_T.t32 1.8255
R1018 IM_T.n25 IM_T.t43 1.8255
R1019 IM_T.n26 IM_T.t48 1.8255
R1020 IM_T.n27 IM_T.t13 1.8255
R1021 IM_T.n28 IM_T.t15 1.8255
R1022 IM_T.n29 IM_T.t49 1.8255
R1023 IM_T.n30 IM_T.t33 1.8255
R1024 IM_T.n31 IM_T.t9 1.8255
R1025 IM_T.n32 IM_T.t42 1.8255
R1026 IM_T.n33 IM_T.t61 1.8255
R1027 IM_T.n34 IM_T.t17 1.8255
R1028 IM_T.n35 IM_T.t57 1.8255
R1029 IM_T.n36 IM_T.t5 1.8255
R1030 IM_T.n37 IM_T.t31 1.8255
R1031 IM_T.n38 IM_T.t27 1.8255
R1032 IM_T.n39 IM_T.t55 1.8255
R1033 IM_T.n40 IM_T.t40 1.8255
R1034 IM_T.n41 IM_T.t26 1.8255
R1035 IM_T.n42 IM_T.t58 1.8255
R1036 IM_T.n43 IM_T.t18 1.8255
R1037 IM_T.n44 IM_T.t19 1.8255
R1038 IM_T.n47 IM_T.n46 1.09765
R1039 IM_T.n46 IM_T.n45 0.566812
R1040 IM_T.n66 IM_T.n47 0.0163077
R1041 IM_T IM_T.n66 0.00685294
R1042 IM_T.n49 IM_T.n48 0.00483735
R1043 OUT.n78 OUT.t14 6.89543
R1044 OUT.n31 OUT.t56 6.89543
R1045 OUT.n93 OUT.n47 6.10159
R1046 OUT.n46 OUT.n0 6.10159
R1047 OUT.n78 OUT.n77 3.49485
R1048 OUT.n80 OUT.n73 3.49485
R1049 OUT.n82 OUT.n69 3.49485
R1050 OUT.n84 OUT.n65 3.49485
R1051 OUT.n86 OUT.n61 3.49485
R1052 OUT.n88 OUT.n57 3.49485
R1053 OUT.n90 OUT.n53 3.49485
R1054 OUT.n92 OUT.n49 3.49485
R1055 OUT.n31 OUT.n30 3.49485
R1056 OUT.n33 OUT.n26 3.49485
R1057 OUT.n35 OUT.n22 3.49485
R1058 OUT.n37 OUT.n18 3.49485
R1059 OUT.n39 OUT.n14 3.49485
R1060 OUT.n41 OUT.n10 3.49485
R1061 OUT.n43 OUT.n6 3.49485
R1062 OUT.n45 OUT.n2 3.49485
R1063 OUT.n91 OUT.n51 3.37159
R1064 OUT.n89 OUT.n55 3.37159
R1065 OUT.n87 OUT.n59 3.37159
R1066 OUT.n85 OUT.n63 3.37159
R1067 OUT.n83 OUT.n67 3.37159
R1068 OUT.n81 OUT.n71 3.37159
R1069 OUT.n79 OUT.n75 3.37159
R1070 OUT.n44 OUT.n4 3.37159
R1071 OUT.n42 OUT.n8 3.37159
R1072 OUT.n40 OUT.n12 3.37159
R1073 OUT.n38 OUT.n16 3.37159
R1074 OUT.n36 OUT.n20 3.37159
R1075 OUT.n34 OUT.n24 3.37159
R1076 OUT.n32 OUT.n28 3.37159
R1077 OUT.n51 OUT.t51 2.7305
R1078 OUT.n51 OUT.n50 2.7305
R1079 OUT.n55 OUT.t22 2.7305
R1080 OUT.n55 OUT.n54 2.7305
R1081 OUT.n59 OUT.t63 2.7305
R1082 OUT.n59 OUT.n58 2.7305
R1083 OUT.n63 OUT.t53 2.7305
R1084 OUT.n63 OUT.n62 2.7305
R1085 OUT.n67 OUT.t49 2.7305
R1086 OUT.n67 OUT.n66 2.7305
R1087 OUT.n71 OUT.t20 2.7305
R1088 OUT.n71 OUT.n70 2.7305
R1089 OUT.n75 OUT.t50 2.7305
R1090 OUT.n75 OUT.n74 2.7305
R1091 OUT.n77 OUT.t45 2.7305
R1092 OUT.n77 OUT.n76 2.7305
R1093 OUT.n73 OUT.t37 2.7305
R1094 OUT.n73 OUT.n72 2.7305
R1095 OUT.n69 OUT.t8 2.7305
R1096 OUT.n69 OUT.n68 2.7305
R1097 OUT.n65 OUT.t32 2.7305
R1098 OUT.n65 OUT.n64 2.7305
R1099 OUT.n61 OUT.t6 2.7305
R1100 OUT.n61 OUT.n60 2.7305
R1101 OUT.n57 OUT.t2 2.7305
R1102 OUT.n57 OUT.n56 2.7305
R1103 OUT.n53 OUT.t54 2.7305
R1104 OUT.n53 OUT.n52 2.7305
R1105 OUT.n49 OUT.t29 2.7305
R1106 OUT.n49 OUT.n48 2.7305
R1107 OUT.n4 OUT.t25 2.7305
R1108 OUT.n4 OUT.n3 2.7305
R1109 OUT.n8 OUT.t1 2.7305
R1110 OUT.n8 OUT.n7 2.7305
R1111 OUT.n12 OUT.t33 2.7305
R1112 OUT.n12 OUT.n11 2.7305
R1113 OUT.n16 OUT.t26 2.7305
R1114 OUT.n16 OUT.n15 2.7305
R1115 OUT.n20 OUT.t18 2.7305
R1116 OUT.n20 OUT.n19 2.7305
R1117 OUT.n24 OUT.t0 2.7305
R1118 OUT.n24 OUT.n23 2.7305
R1119 OUT.n28 OUT.t24 2.7305
R1120 OUT.n28 OUT.n27 2.7305
R1121 OUT.n30 OUT.t41 2.7305
R1122 OUT.n30 OUT.n29 2.7305
R1123 OUT.n26 OUT.t35 2.7305
R1124 OUT.n26 OUT.n25 2.7305
R1125 OUT.n22 OUT.t55 2.7305
R1126 OUT.n22 OUT.n21 2.7305
R1127 OUT.n18 OUT.t11 2.7305
R1128 OUT.n18 OUT.n17 2.7305
R1129 OUT.n14 OUT.t43 2.7305
R1130 OUT.n14 OUT.n13 2.7305
R1131 OUT.n10 OUT.t59 2.7305
R1132 OUT.n10 OUT.n9 2.7305
R1133 OUT.n6 OUT.t13 2.7305
R1134 OUT.n6 OUT.n5 2.7305
R1135 OUT.n2 OUT.t42 2.7305
R1136 OUT.n2 OUT.n1 2.7305
R1137 OUT.n93 OUT.n92 0.794346
R1138 OUT.n92 OUT.n91 0.794346
R1139 OUT.n91 OUT.n90 0.794346
R1140 OUT.n90 OUT.n89 0.794346
R1141 OUT.n89 OUT.n88 0.794346
R1142 OUT.n88 OUT.n87 0.794346
R1143 OUT.n87 OUT.n86 0.794346
R1144 OUT.n86 OUT.n85 0.794346
R1145 OUT.n85 OUT.n84 0.794346
R1146 OUT.n84 OUT.n83 0.794346
R1147 OUT.n83 OUT.n82 0.794346
R1148 OUT.n82 OUT.n81 0.794346
R1149 OUT.n81 OUT.n80 0.794346
R1150 OUT.n80 OUT.n79 0.794346
R1151 OUT.n79 OUT.n78 0.794346
R1152 OUT.n46 OUT.n45 0.794346
R1153 OUT.n45 OUT.n44 0.794346
R1154 OUT.n44 OUT.n43 0.794346
R1155 OUT.n43 OUT.n42 0.794346
R1156 OUT.n42 OUT.n41 0.794346
R1157 OUT.n41 OUT.n40 0.794346
R1158 OUT.n40 OUT.n39 0.794346
R1159 OUT.n39 OUT.n38 0.794346
R1160 OUT.n38 OUT.n37 0.794346
R1161 OUT.n37 OUT.n36 0.794346
R1162 OUT.n36 OUT.n35 0.794346
R1163 OUT.n35 OUT.n34 0.794346
R1164 OUT.n34 OUT.n33 0.794346
R1165 OUT.n33 OUT.n32 0.794346
R1166 OUT.n32 OUT.n31 0.794346
R1167 OUT OUT.n46 0.568215
R1168 OUT OUT.n93 0.48286
C0 OUT IM 4.31f
C1 SD IM_T 3.58f
C2 IM_T IM 8.25f
C3 OUT IM_T 2.97f
C4 SD IM 2.93f
C5 OUT SD 7.2f
.ends

