magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -3261 -1019 3261 1019
<< metal1 >>
rect -2261 13 2261 19
rect -2261 -13 -2255 13
rect -2229 -13 -2179 13
rect -2153 -13 -2103 13
rect -2077 -13 -2027 13
rect -2001 -13 -1951 13
rect -1925 -13 -1875 13
rect -1849 -13 -1799 13
rect -1773 -13 -1723 13
rect -1697 -13 -1647 13
rect -1621 -13 -1571 13
rect -1545 -13 -1495 13
rect -1469 -13 -1419 13
rect -1393 -13 -1343 13
rect -1317 -13 -1267 13
rect -1241 -13 -1191 13
rect -1165 -13 -1115 13
rect -1089 -13 -1039 13
rect -1013 -13 -963 13
rect -937 -13 -887 13
rect -861 -13 -811 13
rect -785 -13 -735 13
rect -709 -13 -659 13
rect -633 -13 -583 13
rect -557 -13 -507 13
rect -481 -13 -431 13
rect -405 -13 -355 13
rect -329 -13 -279 13
rect -253 -13 -203 13
rect -177 -13 -127 13
rect -101 -13 -51 13
rect -25 -13 25 13
rect 51 -13 101 13
rect 127 -13 177 13
rect 203 -13 253 13
rect 279 -13 329 13
rect 355 -13 405 13
rect 431 -13 481 13
rect 507 -13 557 13
rect 583 -13 633 13
rect 659 -13 709 13
rect 735 -13 785 13
rect 811 -13 861 13
rect 887 -13 937 13
rect 963 -13 1013 13
rect 1039 -13 1089 13
rect 1115 -13 1165 13
rect 1191 -13 1241 13
rect 1267 -13 1317 13
rect 1343 -13 1393 13
rect 1419 -13 1469 13
rect 1495 -13 1545 13
rect 1571 -13 1621 13
rect 1647 -13 1697 13
rect 1723 -13 1773 13
rect 1799 -13 1849 13
rect 1875 -13 1925 13
rect 1951 -13 2001 13
rect 2027 -13 2077 13
rect 2103 -13 2153 13
rect 2179 -13 2229 13
rect 2255 -13 2261 13
rect -2261 -19 2261 -13
<< via1 >>
rect -2255 -13 -2229 13
rect -2179 -13 -2153 13
rect -2103 -13 -2077 13
rect -2027 -13 -2001 13
rect -1951 -13 -1925 13
rect -1875 -13 -1849 13
rect -1799 -13 -1773 13
rect -1723 -13 -1697 13
rect -1647 -13 -1621 13
rect -1571 -13 -1545 13
rect -1495 -13 -1469 13
rect -1419 -13 -1393 13
rect -1343 -13 -1317 13
rect -1267 -13 -1241 13
rect -1191 -13 -1165 13
rect -1115 -13 -1089 13
rect -1039 -13 -1013 13
rect -963 -13 -937 13
rect -887 -13 -861 13
rect -811 -13 -785 13
rect -735 -13 -709 13
rect -659 -13 -633 13
rect -583 -13 -557 13
rect -507 -13 -481 13
rect -431 -13 -405 13
rect -355 -13 -329 13
rect -279 -13 -253 13
rect -203 -13 -177 13
rect -127 -13 -101 13
rect -51 -13 -25 13
rect 25 -13 51 13
rect 101 -13 127 13
rect 177 -13 203 13
rect 253 -13 279 13
rect 329 -13 355 13
rect 405 -13 431 13
rect 481 -13 507 13
rect 557 -13 583 13
rect 633 -13 659 13
rect 709 -13 735 13
rect 785 -13 811 13
rect 861 -13 887 13
rect 937 -13 963 13
rect 1013 -13 1039 13
rect 1089 -13 1115 13
rect 1165 -13 1191 13
rect 1241 -13 1267 13
rect 1317 -13 1343 13
rect 1393 -13 1419 13
rect 1469 -13 1495 13
rect 1545 -13 1571 13
rect 1621 -13 1647 13
rect 1697 -13 1723 13
rect 1773 -13 1799 13
rect 1849 -13 1875 13
rect 1925 -13 1951 13
rect 2001 -13 2027 13
rect 2077 -13 2103 13
rect 2153 -13 2179 13
rect 2229 -13 2255 13
<< metal2 >>
rect -2261 13 2261 19
rect -2261 -13 -2255 13
rect -2229 -13 -2179 13
rect -2153 -13 -2103 13
rect -2077 -13 -2027 13
rect -2001 -13 -1951 13
rect -1925 -13 -1875 13
rect -1849 -13 -1799 13
rect -1773 -13 -1723 13
rect -1697 -13 -1647 13
rect -1621 -13 -1571 13
rect -1545 -13 -1495 13
rect -1469 -13 -1419 13
rect -1393 -13 -1343 13
rect -1317 -13 -1267 13
rect -1241 -13 -1191 13
rect -1165 -13 -1115 13
rect -1089 -13 -1039 13
rect -1013 -13 -963 13
rect -937 -13 -887 13
rect -861 -13 -811 13
rect -785 -13 -735 13
rect -709 -13 -659 13
rect -633 -13 -583 13
rect -557 -13 -507 13
rect -481 -13 -431 13
rect -405 -13 -355 13
rect -329 -13 -279 13
rect -253 -13 -203 13
rect -177 -13 -127 13
rect -101 -13 -51 13
rect -25 -13 25 13
rect 51 -13 101 13
rect 127 -13 177 13
rect 203 -13 253 13
rect 279 -13 329 13
rect 355 -13 405 13
rect 431 -13 481 13
rect 507 -13 557 13
rect 583 -13 633 13
rect 659 -13 709 13
rect 735 -13 785 13
rect 811 -13 861 13
rect 887 -13 937 13
rect 963 -13 1013 13
rect 1039 -13 1089 13
rect 1115 -13 1165 13
rect 1191 -13 1241 13
rect 1267 -13 1317 13
rect 1343 -13 1393 13
rect 1419 -13 1469 13
rect 1495 -13 1545 13
rect 1571 -13 1621 13
rect 1647 -13 1697 13
rect 1723 -13 1773 13
rect 1799 -13 1849 13
rect 1875 -13 1925 13
rect 1951 -13 2001 13
rect 2027 -13 2077 13
rect 2103 -13 2153 13
rect 2179 -13 2229 13
rect 2255 -13 2261 13
rect -2261 -19 2261 -13
<< end >>
