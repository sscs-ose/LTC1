magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1071 -1019 1071 1019
<< metal1 >>
rect -71 13 71 19
rect -71 -13 -65 13
rect 65 -13 71 13
rect -71 -19 71 -13
<< via1 >>
rect -65 -13 65 13
<< metal2 >>
rect -71 13 71 19
rect -71 -13 -65 13
rect 65 -13 71 13
rect -71 -19 71 -13
<< end >>
