magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2000 -2000 17064 59297
<< isosubstrate >>
rect 294 20724 14770 56850
rect 1350 15369 13714 20724
<< psubdiff >>
rect 3116 19749 11948 19993
rect 3116 19267 3360 19749
rect 11704 19267 11948 19749
rect 3116 18869 11948 19267
rect 3116 18395 3360 18869
rect 11704 18395 11948 18869
rect 3116 17997 11948 18395
rect 3116 17523 3360 17997
rect 11704 17523 11948 17997
rect 3116 17125 11948 17523
rect 3116 16643 3360 17125
rect 11704 16643 11948 17125
rect 3116 16399 11948 16643
<< metal1 >>
rect 0 20368 122 57254
rect 388 56398 14676 56756
rect 388 52450 14676 53098
rect 388 48502 14676 49150
rect 388 44554 14676 45202
rect 388 40606 14676 41254
rect 388 36658 14676 37306
rect 388 32710 14676 33358
rect 388 28762 14676 29410
rect 388 24814 14676 25462
rect 388 21156 14676 21514
rect 0 19368 300 20368
rect 2862 20262 2948 20630
rect 12116 20262 12202 20630
rect 14942 20368 15064 57254
rect 3127 19760 11937 19982
rect 0 19168 122 19368
rect 3127 19256 3349 19760
rect 11715 19256 11937 19760
rect 14764 19368 15064 20368
rect 0 18168 300 19168
rect 3127 18880 11937 19256
rect 14942 19168 15064 19368
rect 3127 18384 3349 18880
rect 11715 18384 11937 18880
rect 0 17968 122 18168
rect 3127 18008 11937 18384
rect 14764 18168 15064 19168
rect 0 16968 300 17968
rect 3127 17512 3349 18008
rect 11715 17512 11937 18008
rect 14942 17968 15064 18168
rect 3127 17136 11937 17512
rect 0 16768 122 16968
rect 0 15768 300 16768
rect 3127 16632 3349 17136
rect 11715 16632 11937 17136
rect 14764 16968 15064 17968
rect 14942 16768 15064 16968
rect 3127 16410 11937 16632
rect 0 15568 122 15768
rect 2862 15762 2948 16130
rect 12116 15762 12202 16130
rect 14764 15768 15064 16768
rect 14942 15568 15064 15768
rect 0 14568 300 15568
rect 14764 14568 15064 15568
rect 0 14368 122 14568
rect 14942 14368 15064 14568
rect 0 13368 300 14368
rect 14764 13368 15064 14368
rect 0 13168 122 13368
rect 14942 13168 15064 13368
rect 0 12168 300 13168
rect 14764 12168 15064 13168
rect 0 11968 122 12168
rect 14942 11968 15064 12168
rect 0 10968 300 11968
rect 14764 10968 15064 11968
rect 0 10768 122 10968
rect 14942 10768 15064 10968
rect 0 9768 300 10768
rect 14764 9768 15064 10768
rect 0 9100 122 9768
rect 14942 9100 15064 9768
rect 0 8100 300 9100
rect 14764 8100 15064 9100
rect 0 7900 122 8100
rect 14942 7900 15064 8100
rect 0 6900 300 7900
rect 14764 6900 15064 7900
rect 0 6700 122 6900
rect 14942 6700 15064 6900
rect 0 5700 300 6700
rect 14764 5700 15064 6700
rect 0 5500 122 5700
rect 14942 5500 15064 5700
rect 0 4500 300 5500
rect 14764 4500 15064 5500
rect 0 4300 122 4500
rect 14942 4300 15064 4500
rect 0 3300 300 4300
rect 14764 3300 15064 4300
rect 0 3100 122 3300
rect 14942 3100 15064 3300
rect 0 2100 300 3100
rect 14764 2100 15064 3100
rect 0 1900 122 2100
rect 14942 1900 15064 2100
rect 0 900 300 1900
rect 14764 900 15064 1900
rect 0 405 122 900
rect 14942 405 15064 900
<< metal2 >>
rect 32 50897 122 52297
rect 32 36497 122 37897
rect 260 900 768 56975
rect 828 38097 1028 50697
rect 1136 900 1336 53160
rect 1396 15762 1904 56975
rect 1964 15762 2472 56975
rect 2532 15762 3040 56975
rect 3668 15762 4176 56975
rect 4804 15762 5312 56975
rect 5940 15762 6448 56975
rect 7076 15762 7502 56975
rect 7562 15762 7988 56975
rect 8616 15762 9124 56975
rect 9752 15762 10260 56975
rect 10888 15762 11396 56975
rect 12024 15762 12532 56975
rect 12592 15762 13100 56975
rect 13160 52427 13668 56975
rect 13160 36497 13360 52297
rect 13468 36260 13668 52427
rect 13160 15762 13668 36260
rect 13728 900 14236 56975
rect 14296 900 14804 56975
rect 14942 50897 15032 52297
rect 14942 36497 15032 37897
use comp018green_esd_hbm  comp018green_esd_hbm_0
timestamp 1713338890
transform 1 0 1401 0 1 857
box -51 -857 12313 56440
use M1_NWELL_CDNS_40661953145380  M1_NWELL_CDNS_40661953145380_0
timestamp 1713338890
transform 1 0 2678 0 1 18196
box -278 -2528 278 2528
use M1_NWELL_CDNS_40661953145380  M1_NWELL_CDNS_40661953145380_1
timestamp 1713338890
transform 1 0 12386 0 1 18196
box -278 -2528 278 2528
use M1_NWELL_CDNS_40661953145384  M1_NWELL_CDNS_40661953145384_0
timestamp 1713338890
transform 1 0 7532 0 1 15946
box -4678 -278 4678 278
use M1_NWELL_CDNS_40661953145384  M1_NWELL_CDNS_40661953145384_1
timestamp 1713338890
transform 1 0 7532 0 1 20446
box -4678 -278 4678 278
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_0
timestamp 1713338890
transform 1 0 7532 0 1 16598
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_1
timestamp 1713338890
transform 1 0 7532 0 1 17478
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_2
timestamp 1713338890
transform 1 0 7532 0 1 17170
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_3
timestamp 1713338890
transform 1 0 7532 0 1 18042
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_4
timestamp 1713338890
transform 1 0 7532 0 1 18350
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_5
timestamp 1713338890
transform 1 0 7532 0 1 19222
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_6
timestamp 1713338890
transform 1 0 7532 0 1 18914
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316521  M1_PSUB_CDNS_6903358316521_7
timestamp 1713338890
transform 1 0 7532 0 1 19794
box -4087 -45 4087 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_0
timestamp 1713338890
transform 1 0 7532 0 1 21190
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_1
timestamp 1713338890
transform 1 0 7532 0 1 25138
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_2
timestamp 1713338890
transform 1 0 7532 0 1 29086
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_3
timestamp 1713338890
transform 1 0 7532 0 1 33034
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_4
timestamp 1713338890
transform 1 0 7532 0 1 36982
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_5
timestamp 1713338890
transform 1 0 7532 0 1 40930
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_6
timestamp 1713338890
transform 1 0 7532 0 1 44878
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_7
timestamp 1713338890
transform 1 0 7532 0 1 48826
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_8
timestamp 1713338890
transform 1 0 7532 0 1 52774
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316522  M1_PSUB_CDNS_6903358316522_9
timestamp 1713338890
transform 1 0 7532 0 1 56722
box -7001 -45 7001 45
use M1_PSUB_CDNS_6903358316525  M1_PSUB_CDNS_6903358316525_0
timestamp 1713338890
transform 1 0 422 0 1 38956
box -45 -17811 45 17811
use M1_PSUB_CDNS_6903358316525  M1_PSUB_CDNS_6903358316525_1
timestamp 1713338890
transform 1 0 14642 0 1 38956
box -45 -17811 45 17811
use M1_PSUB_CDNS_6903358316526  M1_PSUB_CDNS_6903358316526_0
timestamp 1713338890
transform 1 0 7532 0 1 17324
box -4228 -45 4228 45
use M1_PSUB_CDNS_6903358316526  M1_PSUB_CDNS_6903358316526_1
timestamp 1713338890
transform 1 0 7532 0 1 18196
box -4228 -45 4228 45
use M1_PSUB_CDNS_6903358316526  M1_PSUB_CDNS_6903358316526_2
timestamp 1713338890
transform 1 0 7532 0 1 19068
box -4228 -45 4228 45
use M1_PSUB_CDNS_6903358316527  M1_PSUB_CDNS_6903358316527_0
timestamp 1713338890
transform 1 0 7532 0 1 16444
box -4416 -45 4416 45
use M1_PSUB_CDNS_6903358316527  M1_PSUB_CDNS_6903358316527_1
timestamp 1713338890
transform 1 0 7532 0 1 19948
box -4416 -45 4416 45
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_0
timestamp 1713338890
transform 1 0 3315 0 1 16888
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_1
timestamp 1713338890
transform 1 0 11749 0 1 16888
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_2
timestamp 1713338890
transform 1 0 3315 0 1 17760
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_3
timestamp 1713338890
transform 1 0 11749 0 1 17760
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_4
timestamp 1713338890
transform 1 0 3315 0 1 18632
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_5
timestamp 1713338890
transform 1 0 11749 0 1 18632
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_6
timestamp 1713338890
transform 1 0 3315 0 1 19504
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_7
timestamp 1713338890
transform 1 0 11749 0 1 19504
box -45 -327 45 327
use M1_PSUB_CDNS_6903358316548  M1_PSUB_CDNS_6903358316548_0
timestamp 1713338890
transform 1 0 3161 0 1 18196
box -45 -1643 45 1643
use M1_PSUB_CDNS_6903358316548  M1_PSUB_CDNS_6903358316548_1
timestamp 1713338890
transform 1 0 11903 0 1 18196
box -45 -1643 45 1643
use M1_PSUB_CDNS_6903358316549  M1_PSUB_CDNS_6903358316549_0
timestamp 1713338890
transform 1 0 684 0 1 10634
box -395 -9745 395 9745
use M1_PSUB_CDNS_6903358316549  M1_PSUB_CDNS_6903358316549_1
timestamp 1713338890
transform -1 0 14380 0 1 10634
box -395 -9745 395 9745
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_0
timestamp 1713338890
transform 1 0 1128 0 1 23164
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_1
timestamp 1713338890
transform -1 0 13936 0 1 23164
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_2
timestamp 1713338890
transform 1 0 1128 0 1 27112
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_3
timestamp 1713338890
transform -1 0 13936 0 1 27112
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_4
timestamp 1713338890
transform 1 0 1128 0 1 31060
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_5
timestamp 1713338890
transform -1 0 13936 0 1 31060
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_6
timestamp 1713338890
transform 1 0 1128 0 1 35008
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_7
timestamp 1713338890
transform -1 0 13936 0 1 35008
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_8
timestamp 1713338890
transform -1 0 13936 0 1 38956
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_9
timestamp 1713338890
transform -1 0 13936 0 1 42904
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_10
timestamp 1713338890
transform -1 0 13936 0 1 46852
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_11
timestamp 1713338890
transform -1 0 13936 0 1 50800
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_12
timestamp 1713338890
transform 1 0 1128 0 1 54748
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316523  M2_M1_CDNS_6903358316523_13
timestamp 1713338890
transform -1 0 13936 0 1 54748
box -162 -1588 162 1588
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_0
timestamp 1713338890
transform 1 0 3755 0 1 23164
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_1
timestamp 1713338890
transform 1 0 6361 0 1 23164
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_2
timestamp 1713338890
transform -1 0 8703 0 1 23164
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_3
timestamp 1713338890
transform -1 0 11309 0 1 23164
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_4
timestamp 1713338890
transform 1 0 3755 0 1 27112
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_5
timestamp 1713338890
transform 1 0 6361 0 1 27112
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_6
timestamp 1713338890
transform -1 0 8703 0 1 27112
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_7
timestamp 1713338890
transform -1 0 11309 0 1 27112
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_8
timestamp 1713338890
transform 1 0 3755 0 1 31060
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_9
timestamp 1713338890
transform 1 0 6361 0 1 31060
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_10
timestamp 1713338890
transform -1 0 8703 0 1 31060
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_11
timestamp 1713338890
transform -1 0 11309 0 1 31060
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_12
timestamp 1713338890
transform 1 0 3755 0 1 35008
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_13
timestamp 1713338890
transform 1 0 6361 0 1 35008
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_14
timestamp 1713338890
transform -1 0 8703 0 1 35008
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_15
timestamp 1713338890
transform -1 0 11309 0 1 35008
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_16
timestamp 1713338890
transform 1 0 3755 0 1 38956
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_17
timestamp 1713338890
transform 1 0 6361 0 1 38956
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_18
timestamp 1713338890
transform -1 0 8703 0 1 38956
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_19
timestamp 1713338890
transform -1 0 11309 0 1 38956
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_20
timestamp 1713338890
transform 1 0 3755 0 1 42904
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_21
timestamp 1713338890
transform 1 0 6361 0 1 42904
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_22
timestamp 1713338890
transform -1 0 8703 0 1 42904
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_23
timestamp 1713338890
transform -1 0 11309 0 1 42904
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_24
timestamp 1713338890
transform 1 0 3755 0 1 46852
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_25
timestamp 1713338890
transform 1 0 6361 0 1 46852
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_26
timestamp 1713338890
transform -1 0 8703 0 1 46852
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_27
timestamp 1713338890
transform -1 0 11309 0 1 46852
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_28
timestamp 1713338890
transform 1 0 3755 0 1 50800
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_29
timestamp 1713338890
transform 1 0 6361 0 1 50800
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_30
timestamp 1713338890
transform -1 0 8703 0 1 50800
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_31
timestamp 1713338890
transform -1 0 11309 0 1 50800
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_32
timestamp 1713338890
transform 1 0 3755 0 1 54748
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_33
timestamp 1713338890
transform 1 0 6361 0 1 54748
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_34
timestamp 1713338890
transform -1 0 8703 0 1 54748
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316524  M2_M1_CDNS_6903358316524_35
timestamp 1713338890
transform -1 0 11309 0 1 54748
box -38 -1550 38 1550
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_0
timestamp 1713338890
transform 1 0 7414 0 1 23164
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_1
timestamp 1713338890
transform -1 0 7650 0 1 23164
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_2
timestamp 1713338890
transform 1 0 7414 0 1 27112
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_3
timestamp 1713338890
transform -1 0 7650 0 1 27112
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_4
timestamp 1713338890
transform 1 0 7414 0 1 31060
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_5
timestamp 1713338890
transform -1 0 7650 0 1 31060
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_6
timestamp 1713338890
transform 1 0 7414 0 1 35008
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_7
timestamp 1713338890
transform -1 0 7650 0 1 35008
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_8
timestamp 1713338890
transform 1 0 7414 0 1 38956
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_9
timestamp 1713338890
transform -1 0 7650 0 1 38956
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_10
timestamp 1713338890
transform 1 0 7414 0 1 42904
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_11
timestamp 1713338890
transform -1 0 7650 0 1 42904
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_12
timestamp 1713338890
transform 1 0 7414 0 1 46852
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_13
timestamp 1713338890
transform -1 0 7650 0 1 46852
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_14
timestamp 1713338890
transform 1 0 7414 0 1 50800
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_15
timestamp 1713338890
transform -1 0 7650 0 1 50800
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_16
timestamp 1713338890
transform -1 0 7650 0 1 54748
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316528  M2_M1_CDNS_6903358316528_17
timestamp 1713338890
transform 1 0 7414 0 1 54748
box -38 -1496 38 1496
use M2_M1_CDNS_6903358316531  M2_M1_CDNS_6903358316531_0
timestamp 1713338890
transform 1 0 578 0 1 21335
box -146 -146 146 146
use M2_M1_CDNS_6903358316531  M2_M1_CDNS_6903358316531_1
timestamp 1713338890
transform -1 0 14486 0 1 21335
box -146 -146 146 146
use M2_M1_CDNS_6903358316531  M2_M1_CDNS_6903358316531_2
timestamp 1713338890
transform 1 0 578 0 1 56577
box -146 -146 146 146
use M2_M1_CDNS_6903358316531  M2_M1_CDNS_6903358316531_3
timestamp 1713338890
transform -1 0 14486 0 1 56577
box -146 -146 146 146
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_0
timestamp 1713338890
transform 1 0 84 0 1 37197
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_1
timestamp 1713338890
transform 1 0 14980 0 1 37197
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_2
timestamp 1713338890
transform 1 0 14980 0 1 51597
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_3
timestamp 1713338890
transform 1 0 84 0 1 51597
box -38 -686 38 686
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_0
timestamp 1713338890
transform 1 0 6194 0 1 15949
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_1
timestamp 1713338890
transform 1 0 3922 0 1 15949
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_2
timestamp 1713338890
transform 1 0 11142 0 1 15949
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_3
timestamp 1713338890
transform 1 0 8870 0 1 15949
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_4
timestamp 1713338890
transform 1 0 5058 0 1 17324
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_5
timestamp 1713338890
transform 1 0 10006 0 1 17324
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_6
timestamp 1713338890
transform 1 0 5058 0 1 18196
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_7
timestamp 1713338890
transform 1 0 10006 0 1 18196
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_8
timestamp 1713338890
transform 1 0 5058 0 1 19068
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_9
timestamp 1713338890
transform 1 0 10006 0 1 19068
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_10
timestamp 1713338890
transform 1 0 1650 0 1 21335
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_11
timestamp 1713338890
transform 1 0 2786 0 1 21335
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_12
timestamp 1713338890
transform 1 0 5058 0 1 21335
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_13
timestamp 1713338890
transform 1 0 3922 0 1 20443
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_14
timestamp 1713338890
transform 1 0 6194 0 1 20443
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_15
timestamp 1713338890
transform 1 0 8870 0 1 20443
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_16
timestamp 1713338890
transform 1 0 10006 0 1 21335
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_17
timestamp 1713338890
transform 1 0 11142 0 1 20443
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_18
timestamp 1713338890
transform 1 0 12278 0 1 21335
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_19
timestamp 1713338890
transform 1 0 13414 0 1 21335
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_20
timestamp 1713338890
transform 1 0 1650 0 1 56577
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_21
timestamp 1713338890
transform 1 0 2786 0 1 56577
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_22
timestamp 1713338890
transform 1 0 5058 0 1 56577
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_23
timestamp 1713338890
transform 1 0 10006 0 1 56577
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_24
timestamp 1713338890
transform 1 0 12278 0 1 56577
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_25
timestamp 1713338890
transform 1 0 13414 0 1 56577
box -254 -146 254 146
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_0
timestamp 1713338890
transform 1 0 1650 0 1 25138
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_1
timestamp 1713338890
transform 1 0 2786 0 1 25138
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_2
timestamp 1713338890
transform 1 0 5058 0 1 25138
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_3
timestamp 1713338890
transform 1 0 10006 0 1 25138
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_4
timestamp 1713338890
transform 1 0 12278 0 1 25138
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_5
timestamp 1713338890
transform 1 0 13414 0 1 25138
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_6
timestamp 1713338890
transform 1 0 1650 0 1 29086
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_7
timestamp 1713338890
transform 1 0 2786 0 1 29086
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_8
timestamp 1713338890
transform 1 0 5058 0 1 29086
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_9
timestamp 1713338890
transform 1 0 10006 0 1 29086
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_10
timestamp 1713338890
transform 1 0 12278 0 1 29086
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_11
timestamp 1713338890
transform 1 0 13414 0 1 29086
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_12
timestamp 1713338890
transform 1 0 2786 0 1 33034
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_13
timestamp 1713338890
transform 1 0 1650 0 1 33034
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_14
timestamp 1713338890
transform 1 0 5058 0 1 33034
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_15
timestamp 1713338890
transform 1 0 10006 0 1 33034
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_16
timestamp 1713338890
transform 1 0 12278 0 1 33034
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_17
timestamp 1713338890
transform 1 0 13414 0 1 33034
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_18
timestamp 1713338890
transform 1 0 2786 0 1 36982
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_19
timestamp 1713338890
transform 1 0 1650 0 1 36982
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_20
timestamp 1713338890
transform 1 0 5058 0 1 36982
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_21
timestamp 1713338890
transform 1 0 10006 0 1 36982
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_22
timestamp 1713338890
transform 1 0 12278 0 1 36982
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_23
timestamp 1713338890
transform 1 0 2786 0 1 40930
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_24
timestamp 1713338890
transform 1 0 1650 0 1 40930
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_25
timestamp 1713338890
transform 1 0 5058 0 1 40930
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_26
timestamp 1713338890
transform 1 0 10006 0 1 40930
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_27
timestamp 1713338890
transform 1 0 12278 0 1 40930
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_28
timestamp 1713338890
transform 1 0 1650 0 1 44878
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_29
timestamp 1713338890
transform 1 0 2786 0 1 44878
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_30
timestamp 1713338890
transform 1 0 5058 0 1 44878
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_31
timestamp 1713338890
transform 1 0 10006 0 1 44878
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_32
timestamp 1713338890
transform 1 0 12278 0 1 44878
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_33
timestamp 1713338890
transform 1 0 1650 0 1 48826
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_34
timestamp 1713338890
transform 1 0 2786 0 1 48826
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_35
timestamp 1713338890
transform 1 0 5058 0 1 48826
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_36
timestamp 1713338890
transform 1 0 10006 0 1 48826
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_37
timestamp 1713338890
transform 1 0 12278 0 1 48826
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_38
timestamp 1713338890
transform 1 0 1650 0 1 52774
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_39
timestamp 1713338890
transform 1 0 2786 0 1 52774
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_40
timestamp 1713338890
transform 1 0 5058 0 1 52774
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_41
timestamp 1713338890
transform 1 0 10006 0 1 52774
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_42
timestamp 1713338890
transform 1 0 12278 0 1 52774
box -224 -286 224 286
use M2_M1_CDNS_6903358316536  M2_M1_CDNS_6903358316536_43
timestamp 1713338890
transform 1 0 13414 0 1 52774
box -224 -286 224 286
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_0
timestamp 1713338890
transform 1 0 578 0 1 25138
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_1
timestamp 1713338890
transform -1 0 14486 0 1 25138
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_2
timestamp 1713338890
transform 1 0 578 0 1 29086
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_3
timestamp 1713338890
transform -1 0 14486 0 1 29086
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_4
timestamp 1713338890
transform 1 0 578 0 1 33034
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_5
timestamp 1713338890
transform -1 0 14486 0 1 33034
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_6
timestamp 1713338890
transform 1 0 578 0 1 36982
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_7
timestamp 1713338890
transform -1 0 14486 0 1 36982
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_8
timestamp 1713338890
transform 1 0 578 0 1 40930
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_9
timestamp 1713338890
transform -1 0 14486 0 1 40930
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_10
timestamp 1713338890
transform 1 0 578 0 1 44878
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_11
timestamp 1713338890
transform -1 0 14486 0 1 44878
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_12
timestamp 1713338890
transform 1 0 578 0 1 48826
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_13
timestamp 1713338890
transform -1 0 14486 0 1 48826
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_14
timestamp 1713338890
transform 1 0 578 0 1 52774
box -146 -254 146 254
use M2_M1_CDNS_6903358316537  M2_M1_CDNS_6903358316537_15
timestamp 1713338890
transform -1 0 14486 0 1 52774
box -146 -254 146 254
use M2_M1_CDNS_6903358316538  M2_M1_CDNS_6903358316538_0
timestamp 1713338890
transform 1 0 13568 0 1 36982
box -100 -286 100 286
use M2_M1_CDNS_6903358316538  M2_M1_CDNS_6903358316538_1
timestamp 1713338890
transform 1 0 13568 0 1 40930
box -100 -286 100 286
use M2_M1_CDNS_6903358316538  M2_M1_CDNS_6903358316538_2
timestamp 1713338890
transform 1 0 13568 0 1 44878
box -100 -286 100 286
use M2_M1_CDNS_6903358316538  M2_M1_CDNS_6903358316538_3
timestamp 1713338890
transform 1 0 13568 0 1 48826
box -100 -286 100 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_0
timestamp 1713338890
transform 1 0 7289 0 1 25138
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_1
timestamp 1713338890
transform 1 0 7775 0 1 25138
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_2
timestamp 1713338890
transform 1 0 7289 0 1 29086
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_3
timestamp 1713338890
transform 1 0 7775 0 1 29086
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_4
timestamp 1713338890
transform 1 0 7289 0 1 33034
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_5
timestamp 1713338890
transform 1 0 7775 0 1 33034
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_6
timestamp 1713338890
transform 1 0 7289 0 1 36982
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_7
timestamp 1713338890
transform 1 0 7775 0 1 36982
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_8
timestamp 1713338890
transform 1 0 7289 0 1 40930
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_9
timestamp 1713338890
transform 1 0 7775 0 1 40930
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_10
timestamp 1713338890
transform 1 0 7289 0 1 44878
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_11
timestamp 1713338890
transform 1 0 7775 0 1 44878
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_12
timestamp 1713338890
transform 1 0 7289 0 1 48826
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_13
timestamp 1713338890
transform 1 0 7775 0 1 48826
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_14
timestamp 1713338890
transform 1 0 7289 0 1 52774
box -162 -286 162 286
use M2_M1_CDNS_6903358316539  M2_M1_CDNS_6903358316539_15
timestamp 1713338890
transform 1 0 7775 0 1 52774
box -162 -286 162 286
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_0
timestamp 1713338890
transform 1 0 7289 0 1 17324
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_1
timestamp 1713338890
transform 1 0 7775 0 1 17324
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_2
timestamp 1713338890
transform 1 0 7289 0 1 18196
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_3
timestamp 1713338890
transform 1 0 7775 0 1 18196
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_4
timestamp 1713338890
transform 1 0 7289 0 1 19068
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_5
timestamp 1713338890
transform 1 0 7775 0 1 19068
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_6
timestamp 1713338890
transform 1 0 7289 0 1 21335
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_7
timestamp 1713338890
transform 1 0 7775 0 1 21335
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_8
timestamp 1713338890
transform 1 0 7289 0 1 56577
box -200 -146 200 146
use M2_M1_CDNS_6903358316540  M2_M1_CDNS_6903358316540_9
timestamp 1713338890
transform 1 0 7775 0 1 56577
box -200 -146 200 146
use M2_M1_CDNS_6903358316544  M2_M1_CDNS_6903358316544_0
timestamp 1713338890
transform 1 0 1236 0 1 38956
box -100 -1588 100 1588
use M2_M1_CDNS_6903358316544  M2_M1_CDNS_6903358316544_1
timestamp 1713338890
transform 1 0 1236 0 1 42904
box -100 -1588 100 1588
use M2_M1_CDNS_6903358316544  M2_M1_CDNS_6903358316544_2
timestamp 1713338890
transform 1 0 1236 0 1 46852
box -100 -1588 100 1588
use M2_M1_CDNS_6903358316544  M2_M1_CDNS_6903358316544_3
timestamp 1713338890
transform 1 0 1236 0 1 50800
box -100 -1588 100 1588
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_0
timestamp 1713338890
transform 1 0 5058 0 1 16521
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_1
timestamp 1713338890
transform 1 0 10006 0 1 16521
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_2
timestamp 1713338890
transform 1 0 3922 0 1 16888
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_3
timestamp 1713338890
transform 1 0 6194 0 1 16888
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_4
timestamp 1713338890
transform 1 0 11142 0 1 16888
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_5
timestamp 1713338890
transform 1 0 8870 0 1 16888
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_6
timestamp 1713338890
transform 1 0 3922 0 1 17760
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_7
timestamp 1713338890
transform 1 0 6194 0 1 17760
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_8
timestamp 1713338890
transform 1 0 11142 0 1 17760
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_9
timestamp 1713338890
transform 1 0 8870 0 1 17760
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_10
timestamp 1713338890
transform 1 0 3922 0 1 18632
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_11
timestamp 1713338890
transform 1 0 6194 0 1 18632
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_12
timestamp 1713338890
transform 1 0 11142 0 1 18632
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_13
timestamp 1713338890
transform 1 0 8870 0 1 18632
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_14
timestamp 1713338890
transform 1 0 3922 0 1 19504
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_15
timestamp 1713338890
transform 1 0 5058 0 1 19871
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_16
timestamp 1713338890
transform 1 0 6194 0 1 19504
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_17
timestamp 1713338890
transform 1 0 8870 0 1 19504
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_18
timestamp 1713338890
transform 1 0 10006 0 1 19871
box -254 -92 254 92
use M2_M1_CDNS_6903358316546  M2_M1_CDNS_6903358316546_19
timestamp 1713338890
transform 1 0 11142 0 1 19504
box -254 -92 254 92
use M2_M1_CDNS_6903358316547  M2_M1_CDNS_6903358316547_0
timestamp 1713338890
transform 1 0 7289 0 1 16521
box -200 -92 200 92
use M2_M1_CDNS_6903358316547  M2_M1_CDNS_6903358316547_1
timestamp 1713338890
transform 1 0 7775 0 1 16521
box -200 -92 200 92
use M2_M1_CDNS_6903358316547  M2_M1_CDNS_6903358316547_2
timestamp 1713338890
transform 1 0 7289 0 1 19871
box -200 -92 200 92
use M2_M1_CDNS_6903358316547  M2_M1_CDNS_6903358316547_3
timestamp 1713338890
transform 1 0 7775 0 1 19871
box -200 -92 200 92
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_0
timestamp 1713338890
transform 1 0 1082 0 1 11597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_1
timestamp 1713338890
transform 1 0 2218 0 1 11597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_2
timestamp 1713338890
transform 1 0 3922 0 1 11597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_3
timestamp 1713338890
transform 1 0 6194 0 1 11597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_4
timestamp 1713338890
transform -1 0 8870 0 1 11597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_5
timestamp 1713338890
transform -1 0 11142 0 1 11597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_6
timestamp 1713338890
transform -1 0 12846 0 1 11597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_7
timestamp 1713338890
transform -1 0 13982 0 1 11597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_8
timestamp 1713338890
transform 1 0 514 0 1 13197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_9
timestamp 1713338890
transform 1 0 1650 0 1 13197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_10
timestamp 1713338890
transform 1 0 2786 0 1 13197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_11
timestamp 1713338890
transform 1 0 5058 0 1 13197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_12
timestamp 1713338890
transform -1 0 10006 0 1 13197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_13
timestamp 1713338890
transform -1 0 12278 0 1 13197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_14
timestamp 1713338890
transform -1 0 13414 0 1 13197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_15
timestamp 1713338890
transform -1 0 14550 0 1 13197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_16
timestamp 1713338890
transform 1 0 1082 0 1 29197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_17
timestamp 1713338890
transform 1 0 514 0 1 27597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_18
timestamp 1713338890
transform 1 0 1650 0 1 27597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_19
timestamp 1713338890
transform 1 0 2218 0 1 29197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_20
timestamp 1713338890
transform 1 0 2786 0 1 27597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_21
timestamp 1713338890
transform 1 0 3922 0 1 29197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_22
timestamp 1713338890
transform 1 0 6194 0 1 29197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_23
timestamp 1713338890
transform 1 0 5058 0 1 27597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_24
timestamp 1713338890
transform -1 0 8870 0 1 29197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_25
timestamp 1713338890
transform -1 0 11142 0 1 29197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_26
timestamp 1713338890
transform -1 0 10006 0 1 27597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_27
timestamp 1713338890
transform -1 0 12278 0 1 27597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_28
timestamp 1713338890
transform -1 0 12846 0 1 29197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_29
timestamp 1713338890
transform -1 0 13414 0 1 27597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_30
timestamp 1713338890
transform -1 0 13982 0 1 29197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_31
timestamp 1713338890
transform -1 0 14550 0 1 27597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_32
timestamp 1713338890
transform 1 0 2218 0 1 41997
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_33
timestamp 1713338890
transform 1 0 2218 0 1 40397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_34
timestamp 1713338890
transform 1 0 3922 0 1 41997
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_35
timestamp 1713338890
transform 1 0 3922 0 1 40397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_36
timestamp 1713338890
transform 1 0 6194 0 1 40397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_37
timestamp 1713338890
transform 1 0 6194 0 1 41997
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_38
timestamp 1713338890
transform -1 0 11142 0 1 40397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_39
timestamp 1713338890
transform -1 0 11142 0 1 41997
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_40
timestamp 1713338890
transform -1 0 8870 0 1 41997
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_41
timestamp 1713338890
transform -1 0 8870 0 1 40397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_42
timestamp 1713338890
transform -1 0 12846 0 1 40397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_43
timestamp 1713338890
transform -1 0 13982 0 1 41997
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_44
timestamp 1713338890
transform -1 0 12846 0 1 41997
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_45
timestamp 1713338890
transform -1 0 13982 0 1 40397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_46
timestamp 1713338890
transform 1 0 514 0 1 45197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_47
timestamp 1713338890
transform 1 0 1650 0 1 45197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_48
timestamp 1713338890
transform 1 0 2218 0 1 43597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_49
timestamp 1713338890
transform 1 0 2786 0 1 45197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_50
timestamp 1713338890
transform 1 0 6194 0 1 43597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_51
timestamp 1713338890
transform 1 0 3922 0 1 43597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_52
timestamp 1713338890
transform 1 0 5058 0 1 45197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_53
timestamp 1713338890
transform -1 0 11142 0 1 43597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_54
timestamp 1713338890
transform -1 0 8870 0 1 43597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_55
timestamp 1713338890
transform -1 0 10006 0 1 45197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_56
timestamp 1713338890
transform -1 0 12278 0 1 45197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_57
timestamp 1713338890
transform -1 0 12846 0 1 43597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_58
timestamp 1713338890
transform -1 0 13982 0 1 43597
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_59
timestamp 1713338890
transform -1 0 14550 0 1 45197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_60
timestamp 1713338890
transform 1 0 514 0 1 48397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_61
timestamp 1713338890
transform 1 0 1650 0 1 48397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_62
timestamp 1713338890
transform 1 0 2786 0 1 48397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_63
timestamp 1713338890
transform 1 0 2218 0 1 46797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_64
timestamp 1713338890
transform 1 0 3922 0 1 46797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_65
timestamp 1713338890
transform 1 0 6194 0 1 46797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_66
timestamp 1713338890
transform 1 0 5058 0 1 48397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_67
timestamp 1713338890
transform -1 0 11142 0 1 46797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_68
timestamp 1713338890
transform -1 0 10006 0 1 48397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_69
timestamp 1713338890
transform -1 0 8870 0 1 46797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_70
timestamp 1713338890
transform -1 0 12278 0 1 48397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_71
timestamp 1713338890
transform -1 0 12846 0 1 46797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_72
timestamp 1713338890
transform -1 0 13982 0 1 46797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_73
timestamp 1713338890
transform -1 0 14550 0 1 48397
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_74
timestamp 1713338890
transform 1 0 514 0 1 53197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_75
timestamp 1713338890
transform 1 0 1650 0 1 53197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_76
timestamp 1713338890
transform 1 0 2786 0 1 53197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_77
timestamp 1713338890
transform 1 0 5058 0 1 53197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_78
timestamp 1713338890
transform -1 0 10006 0 1 53197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_79
timestamp 1713338890
transform -1 0 12278 0 1 53197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_80
timestamp 1713338890
transform -1 0 13414 0 1 53197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_81
timestamp 1713338890
transform -1 0 14550 0 1 53197
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_82
timestamp 1713338890
transform 1 0 1082 0 1 54797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_83
timestamp 1713338890
transform 1 0 2218 0 1 54797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_84
timestamp 1713338890
transform 1 0 3922 0 1 54797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_85
timestamp 1713338890
transform 1 0 6194 0 1 54797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_86
timestamp 1713338890
transform -1 0 8870 0 1 54797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_87
timestamp 1713338890
transform -1 0 11142 0 1 54797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_88
timestamp 1713338890
transform -1 0 12846 0 1 54797
box -224 -658 224 658
use M3_M2_CDNS_6903358316520  M3_M2_CDNS_6903358316520_89
timestamp 1713338890
transform -1 0 13982 0 1 54797
box -224 -658 224 658
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_0
timestamp 1713338890
transform 1 0 514 0 1 2797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_1
timestamp 1713338890
transform 1 0 2786 0 1 2797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_2
timestamp 1713338890
transform 1 0 1650 0 1 2797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_3
timestamp 1713338890
transform 1 0 5058 0 1 2797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_4
timestamp 1713338890
transform -1 0 10006 0 1 2797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_5
timestamp 1713338890
transform -1 0 12278 0 1 2797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_6
timestamp 1713338890
transform -1 0 13414 0 1 2797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_7
timestamp 1713338890
transform -1 0 14550 0 1 2797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_8
timestamp 1713338890
transform 1 0 514 0 1 5997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_9
timestamp 1713338890
transform 1 0 2786 0 1 5997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_10
timestamp 1713338890
transform 1 0 1650 0 1 5997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_11
timestamp 1713338890
transform 1 0 5058 0 1 5997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_12
timestamp 1713338890
transform -1 0 10006 0 1 5997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_13
timestamp 1713338890
transform -1 0 12278 0 1 5997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_14
timestamp 1713338890
transform -1 0 13414 0 1 5997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_15
timestamp 1713338890
transform -1 0 14550 0 1 5997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_16
timestamp 1713338890
transform 1 0 514 0 1 9197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_17
timestamp 1713338890
transform 1 0 1650 0 1 9197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_18
timestamp 1713338890
transform 1 0 2786 0 1 9197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_19
timestamp 1713338890
transform 1 0 5058 0 1 9197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_20
timestamp 1713338890
transform -1 0 10006 0 1 9197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_21
timestamp 1713338890
transform -1 0 12278 0 1 9197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_22
timestamp 1713338890
transform -1 0 13414 0 1 9197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_23
timestamp 1713338890
transform -1 0 14550 0 1 9197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_24
timestamp 1713338890
transform 1 0 1082 0 1 15597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_25
timestamp 1713338890
transform 1 0 2218 0 1 15597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_26
timestamp 1713338890
transform 1 0 3922 0 1 15597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_27
timestamp 1713338890
transform 1 0 6194 0 1 15597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_28
timestamp 1713338890
transform -1 0 8870 0 1 15597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_29
timestamp 1713338890
transform -1 0 11142 0 1 15597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_30
timestamp 1713338890
transform -1 0 12846 0 1 15597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_31
timestamp 1713338890
transform -1 0 13982 0 1 15597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_32
timestamp 1713338890
transform 1 0 1082 0 1 18797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_33
timestamp 1713338890
transform 1 0 2218 0 1 18797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_34
timestamp 1713338890
transform 1 0 3922 0 1 18797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_35
timestamp 1713338890
transform 1 0 6194 0 1 18797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_36
timestamp 1713338890
transform -1 0 8870 0 1 18797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_37
timestamp 1713338890
transform -1 0 11142 0 1 18797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_38
timestamp 1713338890
transform -1 0 12846 0 1 18797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_39
timestamp 1713338890
transform -1 0 13982 0 1 18797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_40
timestamp 1713338890
transform 1 0 1082 0 1 25197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_41
timestamp 1713338890
transform 1 0 1082 0 1 21997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_42
timestamp 1713338890
transform 1 0 2218 0 1 21997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_43
timestamp 1713338890
transform 1 0 2218 0 1 25197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_44
timestamp 1713338890
transform 1 0 3922 0 1 25197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_45
timestamp 1713338890
transform 1 0 3922 0 1 21997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_46
timestamp 1713338890
transform 1 0 6194 0 1 25197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_47
timestamp 1713338890
transform 1 0 6194 0 1 21997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_48
timestamp 1713338890
transform -1 0 8870 0 1 21997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_49
timestamp 1713338890
transform -1 0 8870 0 1 25197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_50
timestamp 1713338890
transform -1 0 11142 0 1 25197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_51
timestamp 1713338890
transform -1 0 11142 0 1 21997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_52
timestamp 1713338890
transform -1 0 12846 0 1 25197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_53
timestamp 1713338890
transform -1 0 13982 0 1 25197
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_54
timestamp 1713338890
transform -1 0 12846 0 1 21997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_55
timestamp 1713338890
transform -1 0 13982 0 1 21997
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_56
timestamp 1713338890
transform 1 0 1082 0 1 31597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_57
timestamp 1713338890
transform 1 0 2218 0 1 31597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_58
timestamp 1713338890
transform 1 0 3922 0 1 31597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_59
timestamp 1713338890
transform 1 0 6194 0 1 31597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_60
timestamp 1713338890
transform -1 0 11142 0 1 31597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_61
timestamp 1713338890
transform -1 0 8870 0 1 31597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_62
timestamp 1713338890
transform -1 0 12846 0 1 31597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_63
timestamp 1713338890
transform -1 0 13982 0 1 31597
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_64
timestamp 1713338890
transform 1 0 1650 0 1 34797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_65
timestamp 1713338890
transform 1 0 2786 0 1 34797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_66
timestamp 1713338890
transform 1 0 514 0 1 34797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_67
timestamp 1713338890
transform 1 0 5058 0 1 34797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_68
timestamp 1713338890
transform -1 0 10006 0 1 34797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_69
timestamp 1713338890
transform -1 0 14550 0 1 34797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_70
timestamp 1713338890
transform -1 0 13414 0 1 34797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316529  M3_M2_CDNS_6903358316529_71
timestamp 1713338890
transform -1 0 12278 0 1 34797
box -224 -1464 224 1464
use M3_M2_CDNS_6903358316530  M3_M2_CDNS_6903358316530_0
timestamp 1713338890
transform 1 0 2786 0 1 56336
box -224 -596 224 596
use M3_M2_CDNS_6903358316530  M3_M2_CDNS_6903358316530_1
timestamp 1713338890
transform 1 0 1650 0 1 56336
box -224 -596 224 596
use M3_M2_CDNS_6903358316530  M3_M2_CDNS_6903358316530_2
timestamp 1713338890
transform 1 0 514 0 1 56336
box -224 -596 224 596
use M3_M2_CDNS_6903358316530  M3_M2_CDNS_6903358316530_3
timestamp 1713338890
transform 1 0 5058 0 1 56336
box -224 -596 224 596
use M3_M2_CDNS_6903358316530  M3_M2_CDNS_6903358316530_4
timestamp 1713338890
transform -1 0 10006 0 1 56336
box -224 -596 224 596
use M3_M2_CDNS_6903358316530  M3_M2_CDNS_6903358316530_5
timestamp 1713338890
transform -1 0 13414 0 1 56336
box -224 -596 224 596
use M3_M2_CDNS_6903358316530  M3_M2_CDNS_6903358316530_6
timestamp 1713338890
transform -1 0 12278 0 1 56336
box -224 -596 224 596
use M3_M2_CDNS_6903358316530  M3_M2_CDNS_6903358316530_7
timestamp 1713338890
transform -1 0 14550 0 1 56336
box -224 -596 224 596
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_0
timestamp 1713338890
transform 1 0 928 0 1 38797
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_1
timestamp 1713338890
transform -1 0 13260 0 1 37197
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_2
timestamp 1713338890
transform 1 0 1236 0 1 40397
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_3
timestamp 1713338890
transform 1 0 1236 0 1 41997
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_4
timestamp 1713338890
transform 1 0 1236 0 1 43597
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_5
timestamp 1713338890
transform -1 0 13568 0 1 45197
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_6
timestamp 1713338890
transform 1 0 1236 0 1 46797
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_7
timestamp 1713338890
transform -1 0 13568 0 1 48397
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_8
timestamp 1713338890
transform 1 0 928 0 1 49997
box -100 -658 100 658
use M3_M2_CDNS_6903358316532  M3_M2_CDNS_6903358316532_9
timestamp 1713338890
transform -1 0 13260 0 1 51597
box -100 -658 100 658
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_0
timestamp 1713338890
transform 1 0 84 0 1 37197
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_1
timestamp 1713338890
transform 1 0 14980 0 1 37197
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_2
timestamp 1713338890
transform 1 0 14980 0 1 51597
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_3
timestamp 1713338890
transform 1 0 84 0 1 51597
box -38 -686 38 686
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_0
timestamp 1713338890
transform 1 0 7289 0 1 13197
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_1
timestamp 1713338890
transform -1 0 7775 0 1 13197
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_2
timestamp 1713338890
transform 1 0 7289 0 1 27597
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_3
timestamp 1713338890
transform -1 0 7775 0 1 27597
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_4
timestamp 1713338890
transform 1 0 7289 0 1 45197
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_5
timestamp 1713338890
transform -1 0 7775 0 1 45197
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_6
timestamp 1713338890
transform 1 0 7289 0 1 48397
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_7
timestamp 1713338890
transform -1 0 7775 0 1 48397
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_8
timestamp 1713338890
transform 1 0 7289 0 1 53197
box -162 -658 162 658
use M3_M2_CDNS_6903358316541  M3_M2_CDNS_6903358316541_9
timestamp 1713338890
transform -1 0 7775 0 1 53197
box -162 -658 162 658
use M3_M2_CDNS_6903358316542  M3_M2_CDNS_6903358316542_0
timestamp 1713338890
transform -1 0 7775 0 1 56336
box -162 -596 162 596
use M3_M2_CDNS_6903358316542  M3_M2_CDNS_6903358316542_1
timestamp 1713338890
transform 1 0 7289 0 1 56336
box -162 -596 162 596
use M3_M2_CDNS_6903358316543  M3_M2_CDNS_6903358316543_0
timestamp 1713338890
transform 1 0 7289 0 1 2797
box -162 -1464 162 1464
use M3_M2_CDNS_6903358316543  M3_M2_CDNS_6903358316543_1
timestamp 1713338890
transform -1 0 7775 0 1 2797
box -162 -1464 162 1464
use M3_M2_CDNS_6903358316543  M3_M2_CDNS_6903358316543_2
timestamp 1713338890
transform 1 0 7289 0 1 5997
box -162 -1464 162 1464
use M3_M2_CDNS_6903358316543  M3_M2_CDNS_6903358316543_3
timestamp 1713338890
transform -1 0 7775 0 1 5997
box -162 -1464 162 1464
use M3_M2_CDNS_6903358316543  M3_M2_CDNS_6903358316543_4
timestamp 1713338890
transform 1 0 7289 0 1 9197
box -162 -1464 162 1464
use M3_M2_CDNS_6903358316543  M3_M2_CDNS_6903358316543_5
timestamp 1713338890
transform -1 0 7775 0 1 9197
box -162 -1464 162 1464
use M3_M2_CDNS_6903358316543  M3_M2_CDNS_6903358316543_6
timestamp 1713338890
transform 1 0 7289 0 1 34797
box -162 -1464 162 1464
use M3_M2_CDNS_6903358316543  M3_M2_CDNS_6903358316543_7
timestamp 1713338890
transform -1 0 7775 0 1 34797
box -162 -1464 162 1464
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_0
timestamp 1713338890
transform 1 0 878 0 1 21664
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_1
timestamp 1713338890
transform 1 0 4314 0 1 21664
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_2
timestamp 1713338890
transform 1 0 7750 0 1 21664
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_3
timestamp 1713338890
transform 1 0 11186 0 1 21664
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_4
timestamp 1713338890
transform 1 0 878 0 1 25612
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_5
timestamp 1713338890
transform 1 0 4314 0 1 25612
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_6
timestamp 1713338890
transform 1 0 7750 0 1 25612
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_7
timestamp 1713338890
transform 1 0 11186 0 1 25612
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_8
timestamp 1713338890
transform 1 0 878 0 1 29560
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_9
timestamp 1713338890
transform 1 0 4314 0 1 29560
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_10
timestamp 1713338890
transform 1 0 7750 0 1 29560
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_11
timestamp 1713338890
transform 1 0 11186 0 1 29560
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_12
timestamp 1713338890
transform 1 0 878 0 1 33508
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_13
timestamp 1713338890
transform 1 0 4314 0 1 33508
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_14
timestamp 1713338890
transform 1 0 7750 0 1 33508
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_15
timestamp 1713338890
transform 1 0 11186 0 1 33508
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_16
timestamp 1713338890
transform 1 0 878 0 1 37456
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_17
timestamp 1713338890
transform 1 0 4314 0 1 37456
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_18
timestamp 1713338890
transform 1 0 7750 0 1 37456
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_19
timestamp 1713338890
transform 1 0 11186 0 1 37456
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_20
timestamp 1713338890
transform 1 0 878 0 1 41404
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_21
timestamp 1713338890
transform 1 0 4314 0 1 41404
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_22
timestamp 1713338890
transform 1 0 7750 0 1 41404
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_23
timestamp 1713338890
transform 1 0 11186 0 1 41404
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_24
timestamp 1713338890
transform 1 0 878 0 1 45352
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_25
timestamp 1713338890
transform 1 0 4314 0 1 45352
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_26
timestamp 1713338890
transform 1 0 7750 0 1 45352
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_27
timestamp 1713338890
transform 1 0 11186 0 1 45352
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_28
timestamp 1713338890
transform 1 0 878 0 1 49300
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_29
timestamp 1713338890
transform 1 0 4314 0 1 49300
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_30
timestamp 1713338890
transform 1 0 7750 0 1 49300
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_31
timestamp 1713338890
transform 1 0 11186 0 1 49300
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_32
timestamp 1713338890
transform 1 0 878 0 1 53248
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_33
timestamp 1713338890
transform 1 0 4314 0 1 53248
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_34
timestamp 1713338890
transform 1 0 7750 0 1 53248
box -218 -350 3218 3092
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_35
timestamp 1713338890
transform 1 0 11186 0 1 53248
box -218 -350 3218 3092
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_0
timestamp 1713338890
transform 1 0 3532 0 1 16788
box 0 0 8000 200
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_1
timestamp 1713338890
transform 1 0 3532 0 1 17660
box 0 0 8000 200
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_2
timestamp 1713338890
transform 1 0 3532 0 1 18532
box 0 0 8000 200
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_3
timestamp 1713338890
transform 1 0 3532 0 1 19404
box 0 0 8000 200
<< end >>
