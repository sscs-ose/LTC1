* NGSPICE file created from TG_5x_Layout_flat.ext - technology: gf180mcuC

.subckt TG_5x_Layout_flat VIN VOUT VSS VDD CLK
X0 VOUT CLK.t0 VIN.t9 VSS.t8 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 VIN Inverter_Layout_0.OUT.t2 VOUT.t1 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 VOUT Inverter_Layout_0.OUT.t3 VIN.t0 VDD.t6 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 VOUT CLK.t1 VIN.t8 VSS.t7 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 VIN CLK.t3 VOUT.t7 VSS.t3 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 VIN CLK.t4 VOUT.t6 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X6 VOUT CLK.t5 VIN.t7 VSS.t1 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X7 VOUT Inverter_Layout_0.OUT.t4 VIN.t2 VDD.t5 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 VIN Inverter_Layout_0.OUT.t5 VOUT.t10 VDD.t4 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X9 VIN Inverter_Layout_0.OUT.t6 VOUT.t3 VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X10 VIN CLK.t7 VOUT.t4 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 CLK CLK.t7 48.8844
R1 CLK.n4 CLK.t6 34.6755
R2 CLK.n0 CLK.t5 32.4417
R3 CLK.t7 CLK.n3 32.4417
R4 CLK.n1 CLK.n0 23.6425
R5 CLK.n2 CLK.n1 23.6425
R6 CLK.n3 CLK.n2 23.6425
R7 CLK CLK.n4 13.5576
R8 CLK.n4 CLK.t2 13.0362
R9 CLK.n0 CLK.t3 6.51836
R10 CLK.n1 CLK.t0 6.51836
R11 CLK.n2 CLK.t4 6.51836
R12 CLK.n3 CLK.t1 6.51836
R13 VIN.n14 VIN.n0 4.70224
R14 VIN.n7 VIN.n6 3.9605
R15 VIN.n13 VIN.n12 3.50833
R16 VIN.n8 VIN.n2 3.33441
R17 VIN.n7 VIN.n4 3.33441
R18 VIN.n2 VIN.t7 3.2765
R19 VIN.n2 VIN.n1 3.2765
R20 VIN.n6 VIN.t8 3.2765
R21 VIN.n6 VIN.n5 3.2765
R22 VIN.n4 VIN.t9 3.2765
R23 VIN.n4 VIN.n3 3.2765
R24 VIN.n13 VIN.n10 2.88224
R25 VIN.n10 VIN.t0 1.8205
R26 VIN.n10 VIN.n9 1.8205
R27 VIN.n12 VIN.t2 1.8205
R28 VIN.n12 VIN.n11 1.8205
R29 VIN.n8 VIN.n7 0.626587
R30 VIN.n14 VIN.n13 0.626587
R31 VIN.n14 VIN.n8 0.1805
R32 VIN VIN.n14 0.168761
R33 VOUT.n14 VOUT.n0 6.4265
R34 VOUT.n11 VOUT.t4 6.4265
R35 VOUT.n10 VOUT.t1 4.4205
R36 VOUT.n9 VOUT.n8 3.50833
R37 VOUT.n13 VOUT.n2 3.33441
R38 VOUT.n12 VOUT.n4 3.33441
R39 VOUT.n2 VOUT.t7 3.2765
R40 VOUT.n2 VOUT.n1 3.2765
R41 VOUT.n4 VOUT.t6 3.2765
R42 VOUT.n4 VOUT.n3 3.2765
R43 VOUT.n9 VOUT.n6 2.88224
R44 VOUT.n6 VOUT.t3 1.8205
R45 VOUT.n6 VOUT.n5 1.8205
R46 VOUT.n8 VOUT.t10 1.8205
R47 VOUT.n8 VOUT.n7 1.8205
R48 VOUT.n10 VOUT.n9 0.908326
R49 VOUT.n11 VOUT.n10 0.826152
R50 VOUT.n12 VOUT.n11 0.8105
R51 VOUT.n14 VOUT.n13 0.8105
R52 VOUT.n13 VOUT.n12 0.626587
R53 VOUT VOUT.n14 0.303761
R54 VSS.n1 VSS.t0 2254.03
R55 VSS.t3 VSS.t1 1198.16
R56 VSS.t8 VSS.t3 1198.16
R57 VSS.t2 VSS.t8 1198.16
R58 VSS.t7 VSS.t2 1198.16
R59 VSS.t0 VSS.t7 1198.16
R60 VSS.n3 VSS.n0 6.68085
R61 VSS.n3 VSS.n2 2.61175
R62 VSS VSS.n5 2.6005
R63 VSS.n2 VSS.n1 2.6005
R64 VSS.n4 VSS.t4 2.55851
R65 VSS VSS.n3 0.0647857
R66 VSS.n5 VSS.n4 0.0340817
R67 Inverter_Layout_0.OUT Inverter_Layout_0.OUT.t2 51.1321
R68 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.OUT.t5 38.9595
R69 Inverter_Layout_0.OUT.t2 Inverter_Layout_0.OUT.n2 38.9595
R70 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.OUT.n0 23.6425
R71 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.OUT.n1 23.6425
R72 Inverter_Layout_0.OUT.n0 Inverter_Layout_0.OUT.t3 13.0362
R73 Inverter_Layout_0.OUT.n1 Inverter_Layout_0.OUT.t6 13.0362
R74 Inverter_Layout_0.OUT.n2 Inverter_Layout_0.OUT.t4 13.0362
R75 Inverter_Layout_0.OUT Inverter_Layout_0.OUT.t1 6.88041
R76 Inverter_Layout_0.OUT Inverter_Layout_0.OUT.t0 4.70224
R77 VDD.n1 VDD.t7 465.202
R78 VDD.t6 VDD.t4 293.041
R79 VDD.t3 VDD.t6 293.041
R80 VDD.t5 VDD.t3 293.041
R81 VDD.t7 VDD.t5 293.041
R82 VDD.n7 VDD.t0 89.1464
R83 VDD.n3 VDD.n0 4.7942
R84 VDD.n3 VDD.n2 3.19952
R85 VDD.n2 VDD.n1 3.1505
R86 VDD.n6 VDD.n5 3.1505
R87 VDD.n5 VDD.n4 3.1505
R88 VDD VDD.n7 2.46215
R89 VDD VDD.n6 0.0382679
R90 VDD.n6 VDD.n3 0.0270179
C0 VOUT Inverter_Layout_0.OUT 0.165f
C1 VOUT VIN 1.39f
C2 Inverter_Layout_0.OUT VIN 0.0734f
C3 VOUT CLK 0.171f
C4 Inverter_Layout_0.OUT CLK 0.237f
C5 VIN CLK 0.0793f
C6 VIN 0 0.235f
C7 VOUT 0 0.607f
C8 Inverter_Layout_0.OUT 0 0.493f
C9 CLK 0 1.3f
.ends

