** sch_path: /home/shahid/GF180Projects/Top_test3/Top_test/top/xschem/pex_pll_7.sch
**.subckt pex_pll_7
x9 VSS VDD RST_DIV Vdiv net3 pex_CLK_div_110_mag
x11 IPD+ IPD_ net4 net8 LP_op_test VSS VDD_VCO pex_CP_mag
C1 net6 VSS 80.14p m=1
C2 net5 VSS 3.77p m=1
R1 net5 net6 48.84k m=1
x4 net5 VDD LP_op_test S2 VSS net7 pex_a2x1mux_mag
x1 net7 VDD VSS pex_LF_mag
x2 VSS S1 net4 PU_test PU VDD pex_mux_2x1_ibr
x3 VSS S1 net8 PD_test PD VDD pex_mux_2x1_ibr
x5 VSS S1 net2 Vdiv_test Vdiv VDD pex_mux_2x1_ibr
x7 VDD VSS vcntl_test LP_op_test S1 net9 A_MUX_pex
x6 VSS S1 net3 Vo_test VCO_op VDD pex_mux_2x1_ibr
x8 VSS net1 net2 PU PD VDD pex_PFD_layout
x10 VDD_VCO VDD VCO_op VCO_op_bar net9 VSS VCO_PEX
x14 VSS S0 net1 Vref net10 VDD pex_mux_2x1_ibr
x12 VSS VDD RST_DIV Output1 OPA1 OPA0 VCO_op pex_Output_Div_Mag
x13 VSS VDD RST_DIV Output2 OPB1 OPB0 VCO_op pex_Output_Div_Mag
x17 VSS VDD RST_DIV net10 P1 P0 Vref pex_Output_Div_Mag
V12 P1 VSS 0
.save i(v12)
V13 P0 VSS 0
.save i(v13)
VCNTL Vref VSS pulse(3.3 0 0 100p 100p 250n 500n)
.save i(vcntl)
V14 VDD_VCO VSS PWL( 0 0 100n 0 100.001n 3.3)
.save i(v14)
V15 VDD VSS 3.3
.save i(v15)
V16 VSS GND 0
.save i(v16)
V17 RST_DIV VSS PWL( 0 0 10n 0 10.001n 3)
.save i(v17)
V18 F1 VSS 3.3
.save i(v18)
V19 F0 VSS 3.3
.save i(v19)
V20 F2 VSS 3.3
.save i(v20)
V21 OPA0 VSS 3.3
.save i(v21)
V22 OPA1 VSS 3.3
.save i(v22)
V23 OPB0 VSS 3.3
.save i(v23)
V24 OPB1 VSS 0
.save i(v24)
I0 IPD_ VSS 20u
I1 VDD IPD+ 20u
V25 S1 VSS 3.3
.save i(v25)
V26 S0 VSS 3.3
.save i(v26)
V27 S2 VSS 3.3
.save i(v27)
V28 T1 VSS 0
.save i(v28)
V29 T0 VSS 0
.save i(v29)
V30 vcntl_test VSS 1.08
.save i(v30)
V31 Vo_test VSS PWL( 0 0 10n 0 10.001n 3)
.save i(v31)
V32 Vdiv_test VSS pulse(3.3 0 20n 100p 100p 50n 100n)
.save i(v32)
V33 PU_test VSS pulse(3.3 0 50n 100p 100p 75n 100n)
.save i(v33)
V34 PD_test VSS pulse(3.3 0 0 100p 100p 75n 100n)
.save i(v34)
x15 VDD T1 VSS Vco_op Vdiv T0 PU PD test_output pex_mux_4x1_ibr
**** begin user architecture code


.include pex_PFD_layout.spice
.include pex_A_MUX.spice
.include pex_CP_mag.spice
.include pex_a2x1mux_mag.spice
.include pex_LF_mag.spice
.include VCO_PEX.spice
.include pex_CLK_div_110_mag.spice
.include pex_mux_2x1_ibr.spice
.include pex_mux_4x1_ibr.spice
.include pex_Output_Div_Mag.spice
.control
save all
tran 10n 45u
plot v(VCO_op) v(VCO_op_bar)+4
plot v(vcntl)
plot v(Vdiv)
plot v(vref)
**write pll_4.raw
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
* .lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_statistical

**** end user architecture code
**.ends
.GLOBAL GND
.end
