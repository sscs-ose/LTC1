magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1149 -1019 1149 1019
<< metal1 >>
rect -149 13 149 19
rect -149 -13 -143 13
rect 143 -13 149 13
rect -149 -19 149 -13
<< via1 >>
rect -143 -13 143 13
<< metal2 >>
rect -149 13 149 19
rect -149 -13 -143 13
rect 143 -13 149 13
rect -149 -19 149 -13
<< end >>
