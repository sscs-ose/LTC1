magic
tech gf180mcuD
magscale 1 10
timestamp 1713971633
<< checkpaint >>
rect -4075 -2819 7510 3759
<< nwell >>
rect -2001 1624 -917 1632
rect 1083 1624 2885 1631
rect 1990 1043 2885 1624
rect 1083 -739 1128 -159
rect 2199 -177 2400 -151
rect 2199 -642 2352 -177
rect 2107 -715 2444 -642
rect 2199 -739 2352 -715
<< pwell >>
rect -1171 649 -919 1009
rect 1021 647 5127 1016
rect 1136 -87 4626 236
rect 1136 -96 4296 -87
rect 4350 -96 4626 -87
rect 1136 -116 4626 -96
<< psubdiff >>
rect -959 538 -801 556
rect -959 492 -906 538
rect -860 492 -801 538
rect -959 475 -801 492
<< nsubdiff >>
rect 2107 -655 2444 -642
rect 2107 -701 2232 -655
rect 2278 -701 2444 -655
rect 2107 -715 2444 -701
<< psubdiffcont >>
rect -906 492 -860 538
<< nsubdiffcont >>
rect 2232 -701 2278 -655
<< metal1 >>
rect -2075 1660 2321 1706
rect -2075 1035 -2029 1660
rect 1004 1580 2077 1609
rect -1911 1566 -1213 1580
rect -1911 1514 -1902 1566
rect -1850 1514 -1213 1566
rect -1911 1503 -1213 1514
rect -958 1503 -812 1580
rect 1004 1535 1114 1580
rect 2275 1301 2321 1660
rect 4218 1584 5352 1607
rect 4218 1534 5287 1584
rect 5273 1532 5287 1534
rect 5339 1532 5352 1584
rect 5273 1523 5352 1532
rect 2246 1288 2321 1301
rect 2246 1236 2258 1288
rect 2310 1236 2321 1288
rect 2246 1222 2321 1236
rect -1140 1055 -1084 1128
rect -1140 1042 -1050 1055
rect -2075 989 -1738 1035
rect -1140 990 -1117 1042
rect -1065 1035 -1050 1042
rect 1082 1035 1127 1055
rect 1906 1049 1953 1128
rect -1065 990 -706 1035
rect -1140 989 -706 990
rect 1082 989 1364 1035
rect 1906 1002 2219 1049
rect -1140 984 -1050 989
rect 1157 771 1213 989
rect 1145 755 1227 771
rect 1145 703 1160 755
rect 1212 703 1227 755
rect 1145 688 1227 703
rect 78 671 158 684
rect 78 619 92 671
rect 144 666 158 671
rect 144 620 168 666
rect 2172 660 2219 1002
rect 2275 1034 2321 1222
rect 5197 1089 5510 1135
rect 4291 1055 4371 1067
rect 2275 988 2536 1034
rect 4291 1003 4305 1055
rect 4357 1042 4371 1055
rect 4357 1041 4558 1042
rect 4357 1003 4580 1041
rect 4291 996 4580 1003
rect 4291 991 4371 996
rect 3294 673 3416 690
rect 2156 647 2235 660
rect 144 619 158 620
rect 78 607 158 619
rect 2156 595 2169 647
rect 2221 595 2235 647
rect 3294 621 3312 673
rect 3364 666 3416 673
rect 3364 621 3551 666
rect 3294 609 3551 621
rect 3294 603 3416 609
rect 2156 583 2235 595
rect -936 538 -816 556
rect -936 492 -906 538
rect -860 492 -816 538
rect -936 475 -816 492
rect 1033 475 1153 556
rect 2004 542 2081 554
rect 1999 540 2081 542
rect 1999 488 2002 540
rect 2054 488 2081 540
rect 1999 486 2081 488
rect -985 409 -907 424
rect -985 357 -972 409
rect -920 357 -907 409
rect -985 342 -907 357
rect -965 -116 -919 342
rect 1034 337 1163 410
rect 2004 331 2081 486
rect -5 269 85 287
rect -5 217 15 269
rect 67 217 85 269
rect -5 198 85 217
rect 935 72 1011 86
rect 935 20 947 72
rect 999 71 1011 72
rect 999 25 1332 71
rect 999 20 1011 25
rect 935 8 1011 20
rect 855 -90 942 -77
rect -965 -162 -887 -116
rect 855 -142 873 -90
rect 925 -142 942 -90
rect 855 -154 942 -142
rect 1286 -240 1332 25
rect 2172 -104 2219 583
rect 4067 551 4153 553
rect 4051 543 4153 551
rect 2410 532 2468 533
rect 2410 480 2413 532
rect 2465 480 2468 532
rect 2410 479 2468 480
rect 3232 375 3300 531
rect 4051 491 4083 543
rect 4135 491 4153 543
rect 4051 481 4153 491
rect 4051 379 4125 481
rect 2292 263 2381 272
rect 2292 211 2309 263
rect 2361 211 2381 263
rect 2292 210 2381 211
rect 2294 208 2381 210
rect 3194 268 3280 281
rect 4294 278 4343 991
rect 4390 543 4471 559
rect 4390 491 4404 543
rect 4456 491 4471 543
rect 4390 474 4471 491
rect 5235 340 5302 543
rect 3194 216 3211 268
rect 3263 216 3280 268
rect 1888 -150 2219 -104
rect 2302 -163 2369 208
rect 3194 204 3280 216
rect 4266 266 4350 278
rect 4266 214 4282 266
rect 4334 214 4350 266
rect 4266 202 4350 214
rect 4174 82 4256 96
rect 4174 30 4189 82
rect 4241 80 4256 82
rect 4241 34 4506 80
rect 4241 30 4256 34
rect 4174 18 4256 30
rect 4287 -96 4365 -85
rect 4119 -97 4365 -96
rect 4119 -142 4300 -97
rect 4287 -149 4300 -142
rect 4352 -149 4365 -97
rect 4287 -161 4365 -149
rect 4460 -197 4506 34
rect 5464 -105 5510 1089
rect 5195 -107 5510 -105
rect 5127 -151 5510 -107
rect 4460 -243 4574 -197
rect -720 -684 -631 -679
rect -720 -736 -701 -684
rect -649 -736 -631 -684
rect 975 -692 1312 -641
rect 2107 -655 2444 -642
rect 2107 -701 2232 -655
rect 2278 -701 2444 -655
rect 4187 -687 4453 -617
rect 5292 -633 5347 -632
rect 5292 -685 5293 -633
rect 5345 -685 5347 -633
rect 5292 -686 5347 -685
rect 2107 -721 2444 -701
rect -720 -757 -631 -736
<< via1 >>
rect -1902 1514 -1850 1566
rect 5287 1532 5339 1584
rect 2258 1236 2310 1288
rect -1117 990 -1065 1042
rect 1160 703 1212 755
rect 92 619 144 671
rect 4305 1003 4357 1055
rect 2169 595 2221 647
rect 3312 621 3364 673
rect 2002 488 2054 540
rect -972 357 -920 409
rect 15 217 67 269
rect 947 20 999 72
rect 873 -142 925 -90
rect 2413 480 2465 532
rect 4083 491 4135 543
rect 2309 211 2361 263
rect 4404 491 4456 543
rect 3211 216 3263 268
rect 4282 214 4334 266
rect 4189 30 4241 82
rect 4300 -149 4352 -97
rect -701 -736 -649 -684
rect 5293 -685 5345 -633
<< metal2 >>
rect -76 1701 4362 1759
rect -1916 1566 -1833 1580
rect -1916 1514 -1902 1566
rect -1850 1514 -1833 1566
rect -1916 1500 -1833 1514
rect -1908 -756 -1845 1500
rect -1743 -756 -1680 1577
rect -1566 -756 -1503 1582
rect -1400 -756 -1337 1577
rect -1273 -756 -1210 1588
rect -1140 1042 -1050 1055
rect -1140 990 -1117 1042
rect -1065 990 -1050 1042
rect -1140 984 -1050 990
rect -1121 -554 -1062 984
rect -76 684 -18 1701
rect 2246 1296 2320 1301
rect 2194 1293 2320 1296
rect 2114 1288 2320 1293
rect 2114 1236 2258 1288
rect 2310 1236 2320 1288
rect 2114 1228 2320 1236
rect 2114 1004 2179 1228
rect 2246 1222 2320 1228
rect 4304 1067 4362 1701
rect 5273 1584 5357 1607
rect 5273 1532 5287 1584
rect 5339 1532 5357 1584
rect 5273 1523 5357 1532
rect 1792 939 2179 1004
rect 4291 1055 4371 1067
rect 4291 1003 4305 1055
rect 4357 1003 4371 1055
rect 4291 991 4371 1003
rect 1145 755 1227 771
rect 1145 703 1160 755
rect 1212 703 1227 755
rect 1145 688 1227 703
rect -76 671 158 684
rect -76 622 92 671
rect 78 619 92 622
rect 144 619 158 671
rect 1145 635 1209 688
rect 78 607 158 619
rect 1095 577 1209 635
rect -985 418 -907 424
rect 1095 418 1153 577
rect -985 409 1157 418
rect -985 357 -972 409
rect -920 360 1157 409
rect -920 357 -907 360
rect -985 342 -907 357
rect 1792 321 1857 939
rect 3294 673 3416 690
rect 3294 670 3312 673
rect 2200 660 3312 670
rect 2156 647 3312 660
rect 2156 595 2169 647
rect 2221 621 3312 647
rect 3364 670 3416 673
rect 3364 621 3491 670
rect 2221 596 3491 621
rect 2221 595 2235 596
rect 2156 583 2235 595
rect 1987 540 2072 556
rect 4390 553 4471 559
rect 1987 488 2002 540
rect 2054 517 2072 540
rect 4067 543 4471 553
rect 2383 532 2481 539
rect 2383 517 2413 532
rect 2054 488 2413 517
rect 1987 480 2413 488
rect 2465 480 2481 532
rect 4067 491 4083 543
rect 4135 491 4404 543
rect 4456 491 4471 543
rect 4067 483 4471 491
rect 4067 481 4153 483
rect 1987 473 2481 480
rect 4390 474 4471 483
rect 2000 460 2481 473
rect 2000 459 2244 460
rect 2000 445 2058 459
rect -5 271 85 287
rect -17 269 266 271
rect -17 217 15 269
rect 67 217 266 269
rect -17 207 266 217
rect -5 198 85 207
rect 202 79 266 207
rect 1219 256 1857 321
rect 2300 337 4344 404
rect 2300 272 2367 337
rect 3194 274 3280 281
rect 4277 278 4344 337
rect 2292 263 2381 272
rect 935 79 1011 86
rect 202 72 1011 79
rect 202 20 947 72
rect 999 20 1011 72
rect 202 15 1011 20
rect 935 8 1011 15
rect 855 -88 942 -77
rect 1219 -88 1284 256
rect 2292 211 2309 263
rect 2361 211 2381 263
rect 2292 210 2381 211
rect 2294 208 2381 210
rect 3194 268 3580 274
rect 3194 216 3211 268
rect 3263 216 3580 268
rect 3194 211 3580 216
rect 3194 204 3280 211
rect 3517 91 3580 211
rect 4266 266 4350 278
rect 4266 214 4282 266
rect 4334 214 4350 266
rect 4266 202 4350 214
rect 4174 91 4256 96
rect 3517 82 4256 91
rect 3517 30 4189 82
rect 4241 30 4256 82
rect 3517 28 4256 30
rect 4125 26 4256 28
rect 4174 18 4256 26
rect 855 -90 1284 -88
rect 855 -142 873 -90
rect 925 -142 1284 -90
rect 855 -149 1284 -142
rect 4287 -97 4365 -85
rect 4287 -149 4300 -97
rect 4352 -149 4365 -97
rect 855 -154 942 -149
rect 4287 -161 4365 -149
rect 4296 -554 4355 -161
rect -1121 -613 4355 -554
rect 5290 -619 5356 1523
rect 5280 -633 5360 -619
rect -720 -684 -631 -679
rect -720 -736 -701 -684
rect -649 -736 -631 -684
rect 5280 -685 5293 -633
rect 5345 -685 5360 -633
rect 5280 -698 5360 -685
rect -720 -756 -631 -736
rect -1908 -819 -631 -756
use inverter_magic  inverter_magic_2
timestamp 1713185578
transform 1 0 4297 0 1 1051
box 0 -569 1108 580
use inverter_magic  inverter_magic_3
timestamp 1713185578
transform -1 0 5456 0 -1 -159
box 0 -569 1108 580
use inverter_magic  inverter_magic_4
timestamp 1713185578
transform -1 0 2199 0 -1 -159
box 0 -569 1108 580
use inverter_magic  inverter_magic_5
timestamp 1713185578
transform 1 0 -2001 0 1 1044
box 0 -569 1108 580
use inverter_magic  inverter_magic_6
timestamp 1713185578
transform 1 0 1034 0 1 1044
box 0 -569 1108 580
use tg_magic  tg_magic_0
timestamp 1713185578
transform -1 0 1134 0 -1 378
box -2 -52 2031 1117
use tg_magic  tg_magic_1
timestamp 1713185578
transform 1 0 2297 0 1 514
box -2 -52 2031 1117
use tg_magic  tg_magic_2
timestamp 1713185578
transform -1 0 4348 0 -1 378
box -2 -52 2031 1117
use tg_magic  tg_magic_3
timestamp 1713185578
transform 1 0 -917 0 1 515
box -2 -52 2031 1117
<< labels >>
flabel psubdiffcont -883 516 -883 516 0 FreeSans 750 0 0 0 VSS
flabel nsubdiffcont 2255 -678 2255 -678 0 FreeSans 750 0 0 0 VDD
flabel metal1 s -1848 1012 -1848 1012 0 FreeSans 750 0 0 0 CLK
port 1 nsew
flabel metal1 s 5488 450 5488 450 0 FreeSans 750 0 0 0 Q
port 2 nsew
<< end >>
