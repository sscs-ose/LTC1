magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -4162 -2170 4162 2170
<< nwell >>
rect -2162 -170 2162 170
<< pmos >>
rect -1988 -40 -1888 40
rect -1784 -40 -1684 40
rect -1580 -40 -1480 40
rect -1376 -40 -1276 40
rect -1172 -40 -1072 40
rect -968 -40 -868 40
rect -764 -40 -664 40
rect -560 -40 -460 40
rect -356 -40 -256 40
rect -152 -40 -52 40
rect 52 -40 152 40
rect 256 -40 356 40
rect 460 -40 560 40
rect 664 -40 764 40
rect 868 -40 968 40
rect 1072 -40 1172 40
rect 1276 -40 1376 40
rect 1480 -40 1580 40
rect 1684 -40 1784 40
rect 1888 -40 1988 40
<< pdiff >>
rect -2076 23 -1988 40
rect -2076 -23 -2063 23
rect -2017 -23 -1988 23
rect -2076 -40 -1988 -23
rect -1888 23 -1784 40
rect -1888 -23 -1859 23
rect -1813 -23 -1784 23
rect -1888 -40 -1784 -23
rect -1684 23 -1580 40
rect -1684 -23 -1655 23
rect -1609 -23 -1580 23
rect -1684 -40 -1580 -23
rect -1480 23 -1376 40
rect -1480 -23 -1451 23
rect -1405 -23 -1376 23
rect -1480 -40 -1376 -23
rect -1276 23 -1172 40
rect -1276 -23 -1247 23
rect -1201 -23 -1172 23
rect -1276 -40 -1172 -23
rect -1072 23 -968 40
rect -1072 -23 -1043 23
rect -997 -23 -968 23
rect -1072 -40 -968 -23
rect -868 23 -764 40
rect -868 -23 -839 23
rect -793 -23 -764 23
rect -868 -40 -764 -23
rect -664 23 -560 40
rect -664 -23 -635 23
rect -589 -23 -560 23
rect -664 -40 -560 -23
rect -460 23 -356 40
rect -460 -23 -431 23
rect -385 -23 -356 23
rect -460 -40 -356 -23
rect -256 23 -152 40
rect -256 -23 -227 23
rect -181 -23 -152 23
rect -256 -40 -152 -23
rect -52 23 52 40
rect -52 -23 -23 23
rect 23 -23 52 23
rect -52 -40 52 -23
rect 152 23 256 40
rect 152 -23 181 23
rect 227 -23 256 23
rect 152 -40 256 -23
rect 356 23 460 40
rect 356 -23 385 23
rect 431 -23 460 23
rect 356 -40 460 -23
rect 560 23 664 40
rect 560 -23 589 23
rect 635 -23 664 23
rect 560 -40 664 -23
rect 764 23 868 40
rect 764 -23 793 23
rect 839 -23 868 23
rect 764 -40 868 -23
rect 968 23 1072 40
rect 968 -23 997 23
rect 1043 -23 1072 23
rect 968 -40 1072 -23
rect 1172 23 1276 40
rect 1172 -23 1201 23
rect 1247 -23 1276 23
rect 1172 -40 1276 -23
rect 1376 23 1480 40
rect 1376 -23 1405 23
rect 1451 -23 1480 23
rect 1376 -40 1480 -23
rect 1580 23 1684 40
rect 1580 -23 1609 23
rect 1655 -23 1684 23
rect 1580 -40 1684 -23
rect 1784 23 1888 40
rect 1784 -23 1813 23
rect 1859 -23 1888 23
rect 1784 -40 1888 -23
rect 1988 23 2076 40
rect 1988 -23 2017 23
rect 2063 -23 2076 23
rect 1988 -40 2076 -23
<< pdiffc >>
rect -2063 -23 -2017 23
rect -1859 -23 -1813 23
rect -1655 -23 -1609 23
rect -1451 -23 -1405 23
rect -1247 -23 -1201 23
rect -1043 -23 -997 23
rect -839 -23 -793 23
rect -635 -23 -589 23
rect -431 -23 -385 23
rect -227 -23 -181 23
rect -23 -23 23 23
rect 181 -23 227 23
rect 385 -23 431 23
rect 589 -23 635 23
rect 793 -23 839 23
rect 997 -23 1043 23
rect 1201 -23 1247 23
rect 1405 -23 1451 23
rect 1609 -23 1655 23
rect 1813 -23 1859 23
rect 2017 -23 2063 23
<< polysilicon >>
rect -1988 40 -1888 84
rect -1784 40 -1684 84
rect -1580 40 -1480 84
rect -1376 40 -1276 84
rect -1172 40 -1072 84
rect -968 40 -868 84
rect -764 40 -664 84
rect -560 40 -460 84
rect -356 40 -256 84
rect -152 40 -52 84
rect 52 40 152 84
rect 256 40 356 84
rect 460 40 560 84
rect 664 40 764 84
rect 868 40 968 84
rect 1072 40 1172 84
rect 1276 40 1376 84
rect 1480 40 1580 84
rect 1684 40 1784 84
rect 1888 40 1988 84
rect -1988 -84 -1888 -40
rect -1784 -84 -1684 -40
rect -1580 -84 -1480 -40
rect -1376 -84 -1276 -40
rect -1172 -84 -1072 -40
rect -968 -84 -868 -40
rect -764 -84 -664 -40
rect -560 -84 -460 -40
rect -356 -84 -256 -40
rect -152 -84 -52 -40
rect 52 -84 152 -40
rect 256 -84 356 -40
rect 460 -84 560 -40
rect 664 -84 764 -40
rect 868 -84 968 -40
rect 1072 -84 1172 -40
rect 1276 -84 1376 -40
rect 1480 -84 1580 -40
rect 1684 -84 1784 -40
rect 1888 -84 1988 -40
<< metal1 >>
rect -2063 23 -2017 38
rect -2063 -38 -2017 -23
rect -1859 23 -1813 38
rect -1859 -38 -1813 -23
rect -1655 23 -1609 38
rect -1655 -38 -1609 -23
rect -1451 23 -1405 38
rect -1451 -38 -1405 -23
rect -1247 23 -1201 38
rect -1247 -38 -1201 -23
rect -1043 23 -997 38
rect -1043 -38 -997 -23
rect -839 23 -793 38
rect -839 -38 -793 -23
rect -635 23 -589 38
rect -635 -38 -589 -23
rect -431 23 -385 38
rect -431 -38 -385 -23
rect -227 23 -181 38
rect -227 -38 -181 -23
rect -23 23 23 38
rect -23 -38 23 -23
rect 181 23 227 38
rect 181 -38 227 -23
rect 385 23 431 38
rect 385 -38 431 -23
rect 589 23 635 38
rect 589 -38 635 -23
rect 793 23 839 38
rect 793 -38 839 -23
rect 997 23 1043 38
rect 997 -38 1043 -23
rect 1201 23 1247 38
rect 1201 -38 1247 -23
rect 1405 23 1451 38
rect 1405 -38 1451 -23
rect 1609 23 1655 38
rect 1609 -38 1655 -23
rect 1813 23 1859 38
rect 1813 -38 1859 -23
rect 2017 23 2063 38
rect 2017 -38 2063 -23
<< end >>
