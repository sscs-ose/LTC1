magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1019 1045 1019
<< metal1 >>
rect -45 13 45 19
rect -45 -13 -39 13
rect 39 -13 45 13
rect -45 -19 45 -13
<< via1 >>
rect -39 -13 39 13
<< metal2 >>
rect -45 13 45 19
rect -45 -13 -39 13
rect 39 -13 45 13
rect -45 -19 45 -13
<< end >>
