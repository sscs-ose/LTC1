** sch_path: /home/shahid/GF180Projects/CP_PFD_dff_inv_nand_/Xschem/CAP/cap80p_test.sch
**.subckt cap80p_test
V1 IN N pwl 0 0 200n 3.3
.save i(v1)
R2 P IN 100k m=1
x1 N P cap80p
V2 N GND 0
.save i(v2)
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
* .lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_statistical



.control
save all
tran 0.1n 200n
write cap80p_test.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  cap80p.sym # of pins=2
** sym_path: /home/shahid/GF180Projects/CP_PFD_dff_inv_nand_/Xschem/CAP/cap80p.sym
** sch_path: /home/shahid/GF180Projects/CP_PFD_dff_inv_nand_/Xschem/CAP/cap80p.sch
.subckt cap80p N P
*.iopin P
*.iopin N
XC1 P N cap_mim_2f0_m4m5_noshield c_width=25e-6 c_length=25e-6 m=64
.ends

.GLOBAL GND
.end
