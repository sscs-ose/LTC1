* NGSPICE file created from pag_res_magic_flat.ext - technology: gf180mcuC

.subckt pag_res_magic_flat A B G E C H F D VDD
X0 a_2255_5317.t0 a_2535_5015.t0 VDD.t41 ppolyf_u r_width=1u r_length=1u
X1 a_4495_2888.t1 a_3095_1282.t0 VDD.t7 ppolyf_u r_width=1u r_length=1u
X2 a_1695_5015.t0 a_1695_4013.t0 VDD.t19 ppolyf_u r_width=1u r_length=1u
X3 a_3935_5015.t0 a_4775_4363.t0 VDD.t9 ppolyf_u r_width=1u r_length=1u
X4 VDD.t50 VDD.t51 VDD.t2 ppolyf_u r_width=1u r_length=1u
X5 a_7295_4013.t1 a_7015_3711.t0 VDD.t37 ppolyf_u r_width=1u r_length=1u
X6 a_6455_2888.t0 a_5615_2236.t1 VDD.t36 ppolyf_u r_width=1u r_length=1u
X7 a_3375_5015.t1 a_3375_4013.t1 VDD.t6 ppolyf_u r_width=1u r_length=1u
X8 a_8975_2888.t1 a_7575_1282.t1 VDD.t0 ppolyf_u r_width=1u r_length=1u
X9 G.t8 a_1695_5015.t1 VDD.t8 ppolyf_u r_width=1u r_length=1u
X10 a_6175_5015.t1 a_6175_4013.t1 VDD.t10 ppolyf_u r_width=1u r_length=1u
X11 F.t3 a_8975_3711.t1 VDD.t5 ppolyf_u r_width=1u r_length=1u
X12 a_7295_2236.t0 a_8415_2586.t1 VDD.t15 ppolyf_u r_width=1u r_length=1u
X13 a_1135_5317.t0 a_1135_5015.t1 VDD.t25 ppolyf_u r_width=1u r_length=1u
X14 a_3655_5317.t1 a_3095_4665.t0 VDD.t34 ppolyf_u r_width=1u r_length=1u
X15 a_5615_5317.t1 a_5615_5015.t1 VDD.t35 ppolyf_u r_width=1u r_length=1u
X16 a_2815_2888.t0 a_3095_2586.t1 VDD.t27 ppolyf_u r_width=1u r_length=1u
X17 a_3375_4665.t0 a_3375_4363.t0 VDD.t1 ppolyf_u r_width=1u r_length=1u
X18 a_3935_4665.t1 a_5895_4363.t1 VDD.t31 ppolyf_u r_width=1u r_length=1u
X19 a_5055_2888.t0 a_4775_2586.t1 VDD.t13 ppolyf_u r_width=1u r_length=1u
X20 E.t2 E.t3 VDD.t26 ppolyf_u r_width=1u r_length=1u
X21 a_7295_2888.t1 a_7575_2586.t1 VDD.t16 ppolyf_u r_width=1u r_length=1u
X22 a_5335_4665.t0 a_5335_4363.t0 VDD.t21 ppolyf_u r_width=1u r_length=1u
X23 a_7855_4665.t1 a_7855_4363.t1 VDD.t43 ppolyf_u r_width=1u r_length=1u
X24 a_6735_2888.t1 a_7015_2586.t1 VDD.t32 ppolyf_u r_width=1u r_length=1u
X25 G.t0 G.t1 VDD.t20 ppolyf_u r_width=1u r_length=1u
X26 VDD.t46 VDD.t47 VDD.t38 ppolyf_u r_width=1u r_length=1u
X27 a_2255_5317.t1 a_575_3711.t1 VDD.t19 ppolyf_u r_width=1u r_length=1u
X28 a_4495_5317.t1 a_4775_5015.t1 VDD.t9 ppolyf_u r_width=1u r_length=1u
X29 a_1135_5317.t1 a_3375_4665.t1 VDD.t6 ppolyf_u r_width=1u r_length=1u
X30 a_6735_5317.t1 a_5335_4013.t1 VDD.t10 ppolyf_u r_width=1u r_length=1u
X31 a_3655_5317.t0 a_3935_4013.t0 VDD.t7 ppolyf_u r_width=1u r_length=1u
X32 a_5335_2236.t1 a_6175_2586.t1 VDD.t28 ppolyf_u r_width=1u r_length=1u
X33 a_5615_5015.t0 a_5615_4013.t1 VDD.t36 ppolyf_u r_width=1u r_length=1u
X34 a_5615_2888.t1 a_7855_2236.t0 VDD.t24 ppolyf_u r_width=1u r_length=1u
X35 a_8135_5317.t0 a_8415_4013.t0 VDD.t0 ppolyf_u r_width=1u r_length=1u
X36 a_8135_2888.t0 a_7575_2236.t1 VDD.t14 ppolyf_u r_width=1u r_length=1u
X37 B.t1 a_8135_4363.t0 VDD.t15 ppolyf_u r_width=1u r_length=1u
X38 a_1975_5317.t1 a_3375_5015.t0 VDD.t1 ppolyf_u r_width=1u r_length=1u
X39 a_5895_5317.t0 a_5055_4665.t0 VDD.t31 ppolyf_u r_width=1u r_length=1u
X40 a_5055_5317.t1 a_5335_5015.t0 VDD.t21 ppolyf_u r_width=1u r_length=1u
X41 a_6455_5317.t1 a_7855_5015.t1 VDD.t43 ppolyf_u r_width=1u r_length=1u
X42 E.t7 a_855_5015.t1 VDD.t20 ppolyf_u r_width=1u r_length=1u
X43 a_3095_4665.t1 a_3095_4363.t1 VDD.t27 ppolyf_u r_width=1u r_length=1u
X44 a_2815_1584.t0 a_2535_1282.t0 VDD.t42 ppolyf_u r_width=1u r_length=1u
X45 a_5055_4665.t1 a_4775_4363.t1 VDD.t13 ppolyf_u r_width=1u r_length=1u
X46 VDD.t3 VDD.t4 VDD.t2 ppolyf_u r_width=1u r_length=1u
X47 a_7295_2888.t0 a_7015_2586.t0 VDD.t37 ppolyf_u r_width=1u r_length=1u
X48 a_575_4665.t0 A.t1 VDD.t26 ppolyf_u r_width=1u r_length=1u
X49 a_7575_4665.t1 a_7575_4363.t0 VDD.t16 ppolyf_u r_width=1u r_length=1u
X50 a_5895_5317.t1 a_7015_4363.t1 VDD.t32 ppolyf_u r_width=1u r_length=1u
X51 a_8975_2888.t0 D.t1 VDD.t5 ppolyf_u r_width=1u r_length=1u
X52 VDD.t48 VDD.t49 VDD.t38 ppolyf_u r_width=1u r_length=1u
X53 a_4495_5317.t0 a_3095_3711.t0 VDD.t7 ppolyf_u r_width=1u r_length=1u
X54 a_6455_5317.t0 a_5615_4665.t1 VDD.t36 ppolyf_u r_width=1u r_length=1u
X55 a_8975_5317.t1 a_7575_3711.t1 VDD.t0 ppolyf_u r_width=1u r_length=1u
X56 a_1135_1934.t1 C.t2 VDD.t30 ppolyf_u r_width=1u r_length=1u
X57 a_7295_4665.t0 a_8415_5015.t0 VDD.t15 ppolyf_u r_width=1u r_length=1u
X58 a_3935_1584.t1 a_3935_1282.t0 VDD.t29 ppolyf_u r_width=1u r_length=1u
X59 G.t2 G.t3 VDD.t33 ppolyf_u r_width=1u r_length=1u
X60 a_6175_4665.t0 a_5895_4363.t0 VDD.t28 ppolyf_u r_width=1u r_length=1u
X61 a_7855_5015.t0 a_7855_4013.t0 VDD.t24 ppolyf_u r_width=1u r_length=1u
X62 a_6175_4665.t1 a_8135_4363.t1 VDD.t14 ppolyf_u r_width=1u r_length=1u
X63 a_2815_5317.t1 a_3095_5015.t1 VDD.t27 ppolyf_u r_width=1u r_length=1u
X64 a_1415_2888.t3 a_1415_2888.t4 VDD.t42 ppolyf_u r_width=1u r_length=1u
X65 a_5055_5317.t0 a_4775_5015.t0 VDD.t13 ppolyf_u r_width=1u r_length=1u
X66 a_7295_5317.t0 a_7575_5015.t1 VDD.t16 ppolyf_u r_width=1u r_length=1u
X67 E.t4 E.t5 VDD.t26 ppolyf_u r_width=1u r_length=1u
X68 a_6735_5317.t0 a_7015_5015.t0 VDD.t32 ppolyf_u r_width=1u r_length=1u
X69 VDD.t44 VDD.t45 VDD.t38 ppolyf_u r_width=1u r_length=1u
X70 a_2255_1584.t1 a_2535_1282.t1 VDD.t41 ppolyf_u r_width=1u r_length=1u
X71 VDD.t17 VDD.t18 VDD.t2 ppolyf_u r_width=1u r_length=1u
X72 a_7295_4665.t1 a_7015_4363.t0 VDD.t37 ppolyf_u r_width=1u r_length=1u
X73 a_1135_2586.t1 a_1135_1584.t0 VDD.t30 ppolyf_u r_width=1u r_length=1u
X74 a_8415_5015.t1 B.t2 VDD.t5 ppolyf_u r_width=1u r_length=1u
X75 C.t0 a_1415_1934.t1 VDD.t33 ppolyf_u r_width=1u r_length=1u
X76 a_3935_2236.t0 a_3655_1934.t1 VDD.t29 ppolyf_u r_width=1u r_length=1u
X77 a_5335_4665.t1 a_6175_5015.t0 VDD.t28 ppolyf_u r_width=1u r_length=1u
X78 a_1695_1584.t1 a_1695_1282.t1 VDD.t8 ppolyf_u r_width=1u r_length=1u
X79 a_5615_5317.t0 a_7855_4665.t0 VDD.t24 ppolyf_u r_width=1u r_length=1u
X80 a_8135_5317.t1 a_7575_4665.t0 VDD.t14 ppolyf_u r_width=1u r_length=1u
X81 a_2815_4013.t0 a_2535_3711.t1 VDD.t42 ppolyf_u r_width=1u r_length=1u
X82 a_3095_1934.t1 a_1695_1282.t0 VDD.t34 ppolyf_u r_width=1u r_length=1u
X83 a_1135_1584.t1 G.t9 VDD.t25 ppolyf_u r_width=1u r_length=1u
X84 a_5615_1584.t1 a_4215_1282.t1 VDD.t35 ppolyf_u r_width=1u r_length=1u
X85 a_1415_2888.t1 a_1415_2888.t2 VDD.t41 ppolyf_u r_width=1u r_length=1u
X86 a_1135_4363.t1 C.t3 VDD.t30 ppolyf_u r_width=1u r_length=1u
X87 VDD.t22 VDD.t23 VDD.t2 ppolyf_u r_width=1u r_length=1u
X88 a_7295_5317.t1 a_7015_5015.t1 VDD.t37 ppolyf_u r_width=1u r_length=1u
X89 G.t10 G.t11 VDD.t33 ppolyf_u r_width=1u r_length=1u
X90 a_3935_4013.t1 a_3935_3711.t1 VDD.t29 ppolyf_u r_width=1u r_length=1u
X91 a_2255_1584.t0 a_855_2586.t0 VDD.t19 ppolyf_u r_width=1u r_length=1u
X92 a_8975_5317.t0 D.t0 VDD.t5 ppolyf_u r_width=1u r_length=1u
X93 a_4775_1584.t1 a_4495_1282.t1 VDD.t9 ppolyf_u r_width=1u r_length=1u
X94 a_3375_1934.t1 a_4215_1282.t0 VDD.t6 ppolyf_u r_width=1u r_length=1u
X95 a_6735_1584.t0 a_5335_2586.t0 VDD.t10 ppolyf_u r_width=1u r_length=1u
X96 a_1695_2236.t0 a_1415_1934.t0 VDD.t8 ppolyf_u r_width=1u r_length=1u
X97 a_1695_2236.t1 a_3655_1934.t0 VDD.t34 ppolyf_u r_width=1u r_length=1u
X98 a_1135_2236.t0 a_1135_1934.t0 VDD.t25 ppolyf_u r_width=1u r_length=1u
X99 a_5615_2236.t0 a_5615_1934.t0 VDD.t35 ppolyf_u r_width=1u r_length=1u
X100 a_2255_4013.t0 a_2535_3711.t0 VDD.t41 ppolyf_u r_width=1u r_length=1u
X101 a_5335_1934.t1 a_3935_1282.t1 VDD.t31 ppolyf_u r_width=1u r_length=1u
X102 a_3375_1584.t1 a_3375_1282.t0 VDD.t1 ppolyf_u r_width=1u r_length=1u
X103 a_7855_1584.t1 D.t2 VDD.t43 ppolyf_u r_width=1u r_length=1u
X104 a_5335_1584.t1 a_5055_1282.t1 VDD.t21 ppolyf_u r_width=1u r_length=1u
X105 a_575_1282.t1 a_575_1282.t2 VDD.t20 ppolyf_u r_width=1u r_length=1u
X106 a_1695_2586.t0 a_1695_1584.t0 VDD.t19 ppolyf_u r_width=1u r_length=1u
X107 a_3935_2586.t0 a_4775_1934.t0 VDD.t9 ppolyf_u r_width=1u r_length=1u
X108 a_1695_4013.t1 a_1695_3711.t0 VDD.t8 ppolyf_u r_width=1u r_length=1u
X109 a_3375_2586.t0 a_3375_1584.t0 VDD.t6 ppolyf_u r_width=1u r_length=1u
X110 a_1135_4013.t1 G.t7 VDD.t25 ppolyf_u r_width=1u r_length=1u
X111 a_6175_2586.t0 a_6175_1584.t0 VDD.t10 ppolyf_u r_width=1u r_length=1u
X112 a_3095_4363.t0 a_1695_3711.t1 VDD.t34 ppolyf_u r_width=1u r_length=1u
X113 a_3095_2586.t0 a_4495_1282.t0 VDD.t7 ppolyf_u r_width=1u r_length=1u
X114 a_2815_2888.t1 a_2535_2586.t1 VDD.t42 ppolyf_u r_width=1u r_length=1u
X115 a_5615_4013.t0 a_4215_3711.t0 VDD.t35 ppolyf_u r_width=1u r_length=1u
X116 a_5615_1934.t1 a_3375_1282.t1 VDD.t36 ppolyf_u r_width=1u r_length=1u
X117 a_7575_2586.t0 a_8975_1282.t0 VDD.t0 ppolyf_u r_width=1u r_length=1u
X118 a_8415_1584.t0 H.t1 VDD.t15 ppolyf_u r_width=1u r_length=1u
X119 a_3375_2236.t0 a_3375_1934.t0 VDD.t1 ppolyf_u r_width=1u r_length=1u
X120 a_3935_2236.t1 a_5895_1934.t1 VDD.t31 ppolyf_u r_width=1u r_length=1u
X121 a_5335_2236.t0 a_5335_1934.t0 VDD.t21 ppolyf_u r_width=1u r_length=1u
X122 a_1975_2888.t1 a_1135_2236.t1 VDD.t30 ppolyf_u r_width=1u r_length=1u
X123 a_2255_4013.t1 a_855_5015.t0 VDD.t19 ppolyf_u r_width=1u r_length=1u
X124 a_7855_2236.t1 a_7855_1934.t1 VDD.t43 ppolyf_u r_width=1u r_length=1u
X125 G.t4 G.t5 VDD.t20 ppolyf_u r_width=1u r_length=1u
X126 a_4775_4013.t1 a_4495_3711.t0 VDD.t9 ppolyf_u r_width=1u r_length=1u
X127 a_1415_2888.t0 a_575_2236.t1 VDD.t33 ppolyf_u r_width=1u r_length=1u
X128 a_2815_1584.t1 a_3095_1282.t1 VDD.t27 ppolyf_u r_width=1u r_length=1u
X129 a_1415_2888.t5 a_3935_2586.t1 VDD.t29 ppolyf_u r_width=1u r_length=1u
X130 a_3375_4363.t1 a_4215_3711.t1 VDD.t6 ppolyf_u r_width=1u r_length=1u
X131 a_4775_1584.t0 a_5055_1282.t0 VDD.t13 ppolyf_u r_width=1u r_length=1u
X132 a_6735_4013.t0 a_5335_5015.t1 VDD.t10 ppolyf_u r_width=1u r_length=1u
X133 a_7295_1584.t0 a_7575_1282.t0 VDD.t16 ppolyf_u r_width=1u r_length=1u
X134 E.t0 a_575_1282.t0 VDD.t26 ppolyf_u r_width=1u r_length=1u
X135 a_6735_1584.t1 a_7015_1282.t0 VDD.t32 ppolyf_u r_width=1u r_length=1u
X136 VDD.t52 VDD.t53 VDD.t38 ppolyf_u r_width=1u r_length=1u
X137 a_3655_2888.t1 a_3935_1584.t0 VDD.t7 ppolyf_u r_width=1u r_length=1u
X138 a_8135_2888.t1 a_8415_1584.t1 VDD.t0 ppolyf_u r_width=1u r_length=1u
X139 a_5615_2586.t0 a_5615_1584.t0 VDD.t36 ppolyf_u r_width=1u r_length=1u
X140 a_3375_4013.t0 a_3375_3711.t0 VDD.t1 ppolyf_u r_width=1u r_length=1u
X141 a_5335_4363.t1 a_3935_3711.t0 VDD.t31 ppolyf_u r_width=1u r_length=1u
X142 a_2255_2888.t0 a_2535_2586.t0 VDD.t41 ppolyf_u r_width=1u r_length=1u
X143 B.t3 a_8135_1934.t1 VDD.t15 ppolyf_u r_width=1u r_length=1u
X144 a_1415_5317.t2 a_1415_5317.t3 VDD.t42 ppolyf_u r_width=1u r_length=1u
X145 a_5335_4013.t0 a_5055_3711.t1 VDD.t21 ppolyf_u r_width=1u r_length=1u
X146 a_7855_4013.t1 D.t3 VDD.t43 ppolyf_u r_width=1u r_length=1u
X147 a_6175_1584.t1 a_6175_1282.t0 VDD.t28 ppolyf_u r_width=1u r_length=1u
X148 a_575_3711.t2 a_575_3711.t3 VDD.t20 ppolyf_u r_width=1u r_length=1u
X149 a_7855_1934.t0 F.t1 VDD.t24 ppolyf_u r_width=1u r_length=1u
X150 a_7575_1934.t1 a_6175_1282.t1 VDD.t14 ppolyf_u r_width=1u r_length=1u
X151 a_3095_2236.t0 a_3095_1934.t0 VDD.t27 ppolyf_u r_width=1u r_length=1u
X152 G.t6 a_1695_2586.t1 VDD.t8 ppolyf_u r_width=1u r_length=1u
X153 a_7575_2236.t0 a_7575_1934.t0 VDD.t16 ppolyf_u r_width=1u r_length=1u
X154 a_5055_2236.t1 a_4775_1934.t1 VDD.t13 ppolyf_u r_width=1u r_length=1u
X155 a_1135_5015.t0 a_1135_4013.t0 VDD.t30 ppolyf_u r_width=1u r_length=1u
X156 a_3095_5015.t0 a_4495_3711.t1 VDD.t7 ppolyf_u r_width=1u r_length=1u
X157 a_1135_2888.t0 a_1135_2586.t0 VDD.t25 ppolyf_u r_width=1u r_length=1u
X158 a_575_2236.t0 A.t0 VDD.t26 ppolyf_u r_width=1u r_length=1u
X159 VDD.t56 VDD.t57 VDD.t38 ppolyf_u r_width=1u r_length=1u
X160 a_5895_2888.t0 a_7015_1934.t0 VDD.t32 ppolyf_u r_width=1u r_length=1u
X161 a_3655_2888.t0 a_3095_2236.t1 VDD.t34 ppolyf_u r_width=1u r_length=1u
X162 C.t1 a_1415_4363.t0 VDD.t33 ppolyf_u r_width=1u r_length=1u
X163 a_3935_4665.t0 a_3655_4363.t0 VDD.t29 ppolyf_u r_width=1u r_length=1u
X164 a_5615_4363.t1 a_3375_3711.t1 VDD.t36 ppolyf_u r_width=1u r_length=1u
X165 a_7575_5015.t0 a_8975_3711.t0 VDD.t0 ppolyf_u r_width=1u r_length=1u
X166 a_7295_1584.t1 a_7015_1282.t1 VDD.t37 ppolyf_u r_width=1u r_length=1u
X167 VDD.t54 VDD.t55 VDD.t2 ppolyf_u r_width=1u r_length=1u
X168 a_5615_2888.t0 a_5615_2586.t1 VDD.t35 ppolyf_u r_width=1u r_length=1u
X169 a_8415_4013.t1 H.t0 VDD.t15 ppolyf_u r_width=1u r_length=1u
X170 F.t2 a_8975_1282.t1 VDD.t5 ppolyf_u r_width=1u r_length=1u
X171 a_2815_5317.t0 a_2535_5015.t1 VDD.t42 ppolyf_u r_width=1u r_length=1u
X172 a_6175_2236.t1 a_5895_1934.t0 VDD.t28 ppolyf_u r_width=1u r_length=1u
X173 a_2815_4013.t1 a_3095_3711.t1 VDD.t27 ppolyf_u r_width=1u r_length=1u
X174 a_7855_2586.t0 a_7855_1584.t0 VDD.t24 ppolyf_u r_width=1u r_length=1u
X175 a_6175_2236.t0 a_8135_1934.t0 VDD.t14 ppolyf_u r_width=1u r_length=1u
X176 a_2255_2888.t1 a_575_1282.t3 VDD.t19 ppolyf_u r_width=1u r_length=1u
X177 a_1415_5317.t0 a_1415_5317.t1 VDD.t41 ppolyf_u r_width=1u r_length=1u
X178 a_4775_4013.t0 a_5055_3711.t0 VDD.t13 ppolyf_u r_width=1u r_length=1u
X179 a_4495_2888.t0 a_4775_2586.t0 VDD.t9 ppolyf_u r_width=1u r_length=1u
X180 E.t1 a_575_3711.t0 VDD.t26 ppolyf_u r_width=1u r_length=1u
X181 a_7295_4013.t0 a_7575_3711.t0 VDD.t16 ppolyf_u r_width=1u r_length=1u
X182 a_1135_2888.t1 a_3375_2236.t1 VDD.t6 ppolyf_u r_width=1u r_length=1u
X183 a_6735_4013.t1 a_7015_3711.t1 VDD.t32 ppolyf_u r_width=1u r_length=1u
X184 a_6735_2888.t0 a_5335_1584.t0 VDD.t10 ppolyf_u r_width=1u r_length=1u
X185 VDD.t39 VDD.t40 VDD.t38 ppolyf_u r_width=1u r_length=1u
X186 a_1975_5317.t0 a_1135_4665.t1 VDD.t30 ppolyf_u r_width=1u r_length=1u
X187 a_1415_5317.t4 a_575_4665.t1 VDD.t33 ppolyf_u r_width=1u r_length=1u
X188 a_1415_5317.t5 a_3935_5015.t1 VDD.t29 ppolyf_u r_width=1u r_length=1u
X189 a_7295_2236.t1 a_7015_1934.t1 VDD.t37 ppolyf_u r_width=1u r_length=1u
X190 VDD.t11 VDD.t12 VDD.t2 ppolyf_u r_width=1u r_length=1u
X191 a_1695_4665.t1 a_1415_4363.t1 VDD.t8 ppolyf_u r_width=1u r_length=1u
X192 a_1135_4665.t0 a_1135_4363.t0 VDD.t25 ppolyf_u r_width=1u r_length=1u
X193 a_8415_2586.t0 B.t0 VDD.t5 ppolyf_u r_width=1u r_length=1u
X194 a_5895_2888.t1 a_5055_2236.t0 VDD.t31 ppolyf_u r_width=1u r_length=1u
X195 a_1975_2888.t0 a_3375_2586.t1 VDD.t1 ppolyf_u r_width=1u r_length=1u
X196 a_1695_4665.t0 a_3655_4363.t1 VDD.t34 ppolyf_u r_width=1u r_length=1u
X197 a_6175_4013.t0 a_6175_3711.t0 VDD.t28 ppolyf_u r_width=1u r_length=1u
X198 a_7855_4363.t0 F.t0 VDD.t24 ppolyf_u r_width=1u r_length=1u
X199 a_6455_2888.t1 a_7855_2586.t1 VDD.t43 ppolyf_u r_width=1u r_length=1u
X200 a_5055_2888.t1 a_5335_2586.t1 VDD.t21 ppolyf_u r_width=1u r_length=1u
X201 a_5615_4665.t0 a_5615_4363.t0 VDD.t35 ppolyf_u r_width=1u r_length=1u
X202 a_7575_4363.t1 a_6175_3711.t1 VDD.t14 ppolyf_u r_width=1u r_length=1u
X203 E.t6 a_855_2586.t1 VDD.t20 ppolyf_u r_width=1u r_length=1u
R0 a_2255_5317.t0 a_2255_5317.t1 13.3663
R1 a_2535_5015.t0 a_2535_5015.t1 13.3663
R2 VDD.n291 VDD.t5 9.05773
R3 VDD.n375 VDD.t37 9.05773
R4 VDD.n508 VDD.t21 9.05773
R5 VDD.n999 VDD.t1 9.05773
R6 VDD.n901 VDD.t33 9.05773
R7 VDD.n299 VDD.t0 8.23434
R8 VDD.n387 VDD.t32 8.23434
R9 VDD.n522 VDD.t13 8.23434
R10 VDD.n987 VDD.t27 8.23434
R11 VDD.n893 VDD.t25 8.23434
R12 VDD.n617 VDD.t54 7.09079
R13 VDD.n785 VDD.t50 7.09079
R14 VDD.n51 VDD.t52 7.0013
R15 VDD.n194 VDD.t39 7.0013
R16 VDD.n83 VDD.t46 7.00054
R17 VDD.n240 VDD.t44 7.00054
R18 VDD.n74 VDD.t47 7.00019
R19 VDD.n227 VDD.t45 7.00019
R20 VDD.n67 VDD.t56 6.99979
R21 VDD.n217 VDD.t48 6.99979
R22 VDD.n58 VDD.t57 6.99941
R23 VDD.n204 VDD.t49 6.99941
R24 VDD.n44 VDD.t53 6.99677
R25 VDD.n187 VDD.t40 6.99677
R26 VDD.n610 VDD.t55 6.99412
R27 VDD.n778 VDD.t51 6.99412
R28 VDD.n633 VDD.t11 6.92009
R29 VDD.n803 VDD.t17 6.92009
R30 VDD.n626 VDD.t12 6.91844
R31 VDD.n795 VDD.t18 6.91844
R32 VDD.n655 VDD.t4 6.84254
R33 VDD.n561 VDD.t23 6.84254
R34 VDD.n655 VDD.t3 6.4095
R35 VDD.n561 VDD.t22 6.4095
R36 VDD.n280 VDD.t38 6.17588
R37 VDD.n359 VDD.t16 6.17588
R38 VDD.n488 VDD.t35 6.17588
R39 VDD.n1021 VDD.t34 6.17588
R40 VDD.n913 VDD.t8 6.17588
R41 VDD.n311 VDD.t24 5.3525
R42 VDD.n405 VDD.t10 5.3525
R43 VDD.n544 VDD.t9 5.3525
R44 VDD.n969 VDD.t42 5.3525
R45 VDD.n881 VDD.t20 5.3525
R46 VDD.n347 VDD.t43 3.29404
R47 VDD.n467 VDD.t31 3.29404
R48 VDD.n1042 VDD.t29 3.29404
R49 VDD.n925 VDD.t30 3.29404
R50 VDD.n245 VDD.n244 3.1505
R51 VDD.n182 VDD.n181 3.1505
R52 VDD.n184 VDD.n183 3.1505
R53 VDD.n186 VDD.n185 3.1505
R54 VDD.n189 VDD.n188 3.1505
R55 VDD.n191 VDD.n190 3.1505
R56 VDD.n193 VDD.n192 3.1505
R57 VDD.n197 VDD.n196 3.1505
R58 VDD.n200 VDD.n199 3.1505
R59 VDD.n203 VDD.n202 3.1505
R60 VDD.n207 VDD.n206 3.1505
R61 VDD.n210 VDD.n209 3.1505
R62 VDD.n213 VDD.n212 3.1505
R63 VDD.n216 VDD.n215 3.1505
R64 VDD.n220 VDD.n219 3.1505
R65 VDD.n223 VDD.n222 3.1505
R66 VDD.n226 VDD.n225 3.1505
R67 VDD.n230 VDD.n229 3.1505
R68 VDD.n233 VDD.n232 3.1505
R69 VDD.n236 VDD.n235 3.1505
R70 VDD.n239 VDD.n238 3.1505
R71 VDD.n243 VDD.n242 3.1505
R72 VDD.n773 VDD.n562 3.1505
R73 VDD.n824 VDD.n823 3.1505
R74 VDD.n821 VDD.n820 3.1505
R75 VDD.n818 VDD.n817 3.1505
R76 VDD.n816 VDD.n815 3.1505
R77 VDD.n813 VDD.n812 3.1505
R78 VDD.n811 VDD.n810 3.1505
R79 VDD.n808 VDD.n807 3.1505
R80 VDD.n806 VDD.n805 3.1505
R81 VDD.n802 VDD.n801 3.1505
R82 VDD.n800 VDD.n799 3.1505
R83 VDD.n797 VDD.n796 3.1505
R84 VDD.n794 VDD.n793 3.1505
R85 VDD.n791 VDD.n790 3.1505
R86 VDD.n789 VDD.n788 3.1505
R87 VDD.n787 VDD.n786 3.1505
R88 VDD.n784 VDD.n783 3.1505
R89 VDD.n782 VDD.n781 3.1505
R90 VDD.n780 VDD.n779 3.1505
R91 VDD.n777 VDD.n776 3.1505
R92 VDD.n775 VDD.n774 3.1505
R93 VDD.n826 VDD.n825 3.1505
R94 VDD.n178 VDD.n176 3.1505
R95 VDD.n175 VDD.n173 3.1505
R96 VDD.n172 VDD.n170 3.1505
R97 VDD.n169 VDD.n167 3.1505
R98 VDD.n166 VDD.n164 3.1505
R99 VDD.n163 VDD.n161 3.1505
R100 VDD.n160 VDD.n158 3.1505
R101 VDD.n157 VDD.n155 3.1505
R102 VDD.n154 VDD.n152 3.1505
R103 VDD.n151 VDD.n149 3.1505
R104 VDD.n148 VDD.n146 3.1505
R105 VDD.n145 VDD.n143 3.1505
R106 VDD.n142 VDD.n140 3.1505
R107 VDD.n139 VDD.n137 3.1505
R108 VDD.n136 VDD.n134 3.1505
R109 VDD.n133 VDD.n131 3.1505
R110 VDD.n130 VDD.n128 3.1505
R111 VDD.n127 VDD.n125 3.1505
R112 VDD.n124 VDD.n122 3.1505
R113 VDD.n121 VDD.n119 3.1505
R114 VDD.n118 VDD.n116 3.1505
R115 VDD.n115 VDD.n113 3.1505
R116 VDD.n112 VDD.n110 3.1505
R117 VDD.n109 VDD.n107 3.1505
R118 VDD.n106 VDD.n104 3.1505
R119 VDD.n369 VDD.n368 3.1505
R120 VDD.n375 VDD.n374 3.1505
R121 VDD.n381 VDD.n380 3.1505
R122 VDD.n387 VDD.n386 3.1505
R123 VDD.n393 VDD.n392 3.1505
R124 VDD.n399 VDD.n398 3.1505
R125 VDD.n405 VDD.n404 3.1505
R126 VDD.n411 VDD.n410 3.1505
R127 VDD.n417 VDD.n416 3.1505
R128 VDD.n423 VDD.n422 3.1505
R129 VDD.n429 VDD.n428 3.1505
R130 VDD.n435 VDD.n434 3.1505
R131 VDD.n441 VDD.n440 3.1505
R132 VDD.n447 VDD.n446 3.1505
R133 VDD.n453 VDD.n452 3.1505
R134 VDD.n467 VDD.n466 3.1505
R135 VDD.n473 VDD.n472 3.1505
R136 VDD.n479 VDD.n478 3.1505
R137 VDD.n488 VDD.n487 3.1505
R138 VDD.n495 VDD.n494 3.1505
R139 VDD.n502 VDD.n501 3.1505
R140 VDD.n508 VDD.n507 3.1505
R141 VDD.n516 VDD.n515 3.1505
R142 VDD.n522 VDD.n521 3.1505
R143 VDD.n530 VDD.n529 3.1505
R144 VDD.n537 VDD.n536 3.1505
R145 VDD.n544 VDD.n543 3.1505
R146 VDD.n551 VDD.n550 3.1505
R147 VDD.n558 VDD.n557 3.1505
R148 VDD.n1084 VDD.n1083 3.1505
R149 VDD.n1077 VDD.n1076 3.1505
R150 VDD.n1070 VDD.n1069 3.1505
R151 VDD.n1063 VDD.n1062 3.1505
R152 VDD.n1055 VDD.n1054 3.1505
R153 VDD.n1049 VDD.n1048 3.1505
R154 VDD.n1042 VDD.n1041 3.1505
R155 VDD.n1035 VDD.n1034 3.1505
R156 VDD.n1027 VDD.n1026 3.1505
R157 VDD.n1021 VDD.n1020 3.1505
R158 VDD.n1014 VDD.n1013 3.1505
R159 VDD.n1007 VDD.n1006 3.1505
R160 VDD.n999 VDD.n998 3.1505
R161 VDD.n993 VDD.n992 3.1505
R162 VDD.n987 VDD.n986 3.1505
R163 VDD.n981 VDD.n980 3.1505
R164 VDD.n975 VDD.n974 3.1505
R165 VDD.n969 VDD.n968 3.1505
R166 VDD.n963 VDD.n962 3.1505
R167 VDD.n957 VDD.n956 3.1505
R168 VDD.n951 VDD.n950 3.1505
R169 VDD.n694 VDD.n692 3.1505
R170 VDD.n697 VDD.n695 3.1505
R171 VDD.n700 VDD.n698 3.1505
R172 VDD.n703 VDD.n701 3.1505
R173 VDD.n706 VDD.n704 3.1505
R174 VDD.n709 VDD.n707 3.1505
R175 VDD.n712 VDD.n710 3.1505
R176 VDD.n715 VDD.n713 3.1505
R177 VDD.n718 VDD.n716 3.1505
R178 VDD.n721 VDD.n719 3.1505
R179 VDD.n724 VDD.n722 3.1505
R180 VDD.n727 VDD.n725 3.1505
R181 VDD.n730 VDD.n728 3.1505
R182 VDD.n733 VDD.n731 3.1505
R183 VDD.n736 VDD.n734 3.1505
R184 VDD.n739 VDD.n737 3.1505
R185 VDD.n742 VDD.n740 3.1505
R186 VDD.n745 VDD.n743 3.1505
R187 VDD.n748 VDD.n746 3.1505
R188 VDD.n751 VDD.n749 3.1505
R189 VDD.n754 VDD.n752 3.1505
R190 VDD.n757 VDD.n755 3.1505
R191 VDD.n761 VDD.n759 3.1505
R192 VDD.n764 VDD.n762 3.1505
R193 VDD.n767 VDD.n765 3.1505
R194 VDD.n770 VDD.n768 3.1505
R195 VDD.n772 VDD.n563 3.1505
R196 VDD.n180 VDD.n1 3.1505
R197 VDD.n654 VDD.n653 3.1505
R198 VDD.n87 VDD.n86 3.1505
R199 VDD.n649 VDD.n648 3.1505
R200 VDD.n647 VDD.n646 3.1505
R201 VDD.n645 VDD.n644 3.1505
R202 VDD.n643 VDD.n642 3.1505
R203 VDD.n641 VDD.n640 3.1505
R204 VDD.n639 VDD.n638 3.1505
R205 VDD.n637 VDD.n636 3.1505
R206 VDD.n635 VDD.n634 3.1505
R207 VDD.n632 VDD.n631 3.1505
R208 VDD.n630 VDD.n629 3.1505
R209 VDD.n628 VDD.n627 3.1505
R210 VDD.n625 VDD.n624 3.1505
R211 VDD.n623 VDD.n622 3.1505
R212 VDD.n621 VDD.n620 3.1505
R213 VDD.n619 VDD.n618 3.1505
R214 VDD.n616 VDD.n615 3.1505
R215 VDD.n614 VDD.n613 3.1505
R216 VDD.n612 VDD.n611 3.1505
R217 VDD.n609 VDD.n608 3.1505
R218 VDD.n607 VDD.n606 3.1505
R219 VDD.n605 VDD.n604 3.1505
R220 VDD.n651 VDD.n650 3.1505
R221 VDD.n89 VDD.n88 3.1505
R222 VDD.n770 VDD.n769 3.1505
R223 VDD.n767 VDD.n766 3.1505
R224 VDD.n764 VDD.n763 3.1505
R225 VDD.n761 VDD.n760 3.1505
R226 VDD.n757 VDD.n756 3.1505
R227 VDD.n754 VDD.n753 3.1505
R228 VDD.n751 VDD.n750 3.1505
R229 VDD.n748 VDD.n747 3.1505
R230 VDD.n745 VDD.n744 3.1505
R231 VDD.n742 VDD.n741 3.1505
R232 VDD.n739 VDD.n738 3.1505
R233 VDD.n736 VDD.n735 3.1505
R234 VDD.n733 VDD.n732 3.1505
R235 VDD.n730 VDD.n729 3.1505
R236 VDD.n727 VDD.n726 3.1505
R237 VDD.n724 VDD.n723 3.1505
R238 VDD.n721 VDD.n720 3.1505
R239 VDD.n718 VDD.n717 3.1505
R240 VDD.n715 VDD.n714 3.1505
R241 VDD.n712 VDD.n711 3.1505
R242 VDD.n709 VDD.n708 3.1505
R243 VDD.n706 VDD.n705 3.1505
R244 VDD.n703 VDD.n702 3.1505
R245 VDD.n700 VDD.n699 3.1505
R246 VDD.n697 VDD.n696 3.1505
R247 VDD.n694 VDD.n693 3.1505
R248 VDD.n951 VDD.n949 3.1505
R249 VDD.n957 VDD.n955 3.1505
R250 VDD.n963 VDD.n961 3.1505
R251 VDD.n969 VDD.n967 3.1505
R252 VDD.n975 VDD.n973 3.1505
R253 VDD.n981 VDD.n979 3.1505
R254 VDD.n987 VDD.n985 3.1505
R255 VDD.n993 VDD.n991 3.1505
R256 VDD.n999 VDD.n997 3.1505
R257 VDD.n1007 VDD.n1005 3.1505
R258 VDD.n1014 VDD.n1012 3.1505
R259 VDD.n1021 VDD.n1019 3.1505
R260 VDD.n1027 VDD.n1025 3.1505
R261 VDD.n1035 VDD.n1033 3.1505
R262 VDD.n1042 VDD.n1040 3.1505
R263 VDD.n1049 VDD.n1047 3.1505
R264 VDD.n1055 VDD.n1053 3.1505
R265 VDD.n1063 VDD.n1061 3.1505
R266 VDD.n1070 VDD.n1068 3.1505
R267 VDD.n1077 VDD.n1075 3.1505
R268 VDD.n1084 VDD.n1082 3.1505
R269 VDD.n558 VDD.n556 3.1505
R270 VDD.n551 VDD.n549 3.1505
R271 VDD.n544 VDD.n542 3.1505
R272 VDD.n537 VDD.n535 3.1505
R273 VDD.n530 VDD.n528 3.1505
R274 VDD.n522 VDD.n520 3.1505
R275 VDD.n516 VDD.n514 3.1505
R276 VDD.n508 VDD.n506 3.1505
R277 VDD.n502 VDD.n500 3.1505
R278 VDD.n495 VDD.n493 3.1505
R279 VDD.n488 VDD.n486 3.1505
R280 VDD.n479 VDD.n477 3.1505
R281 VDD.n473 VDD.n471 3.1505
R282 VDD.n467 VDD.n465 3.1505
R283 VDD.n453 VDD.n451 3.1505
R284 VDD.n447 VDD.n445 3.1505
R285 VDD.n441 VDD.n439 3.1505
R286 VDD.n435 VDD.n433 3.1505
R287 VDD.n429 VDD.n427 3.1505
R288 VDD.n423 VDD.n421 3.1505
R289 VDD.n417 VDD.n415 3.1505
R290 VDD.n411 VDD.n409 3.1505
R291 VDD.n405 VDD.n403 3.1505
R292 VDD.n399 VDD.n397 3.1505
R293 VDD.n393 VDD.n391 3.1505
R294 VDD.n387 VDD.n385 3.1505
R295 VDD.n381 VDD.n379 3.1505
R296 VDD.n375 VDD.n373 3.1505
R297 VDD.n369 VDD.n367 3.1505
R298 VDD.n106 VDD.n105 3.1505
R299 VDD.n109 VDD.n108 3.1505
R300 VDD.n112 VDD.n111 3.1505
R301 VDD.n115 VDD.n114 3.1505
R302 VDD.n118 VDD.n117 3.1505
R303 VDD.n121 VDD.n120 3.1505
R304 VDD.n124 VDD.n123 3.1505
R305 VDD.n127 VDD.n126 3.1505
R306 VDD.n130 VDD.n129 3.1505
R307 VDD.n133 VDD.n132 3.1505
R308 VDD.n136 VDD.n135 3.1505
R309 VDD.n139 VDD.n138 3.1505
R310 VDD.n142 VDD.n141 3.1505
R311 VDD.n145 VDD.n144 3.1505
R312 VDD.n148 VDD.n147 3.1505
R313 VDD.n151 VDD.n150 3.1505
R314 VDD.n154 VDD.n153 3.1505
R315 VDD.n157 VDD.n156 3.1505
R316 VDD.n160 VDD.n159 3.1505
R317 VDD.n163 VDD.n162 3.1505
R318 VDD.n166 VDD.n165 3.1505
R319 VDD.n169 VDD.n168 3.1505
R320 VDD.n172 VDD.n171 3.1505
R321 VDD.n175 VDD.n174 3.1505
R322 VDD.n178 VDD.n177 3.1505
R323 VDD.n85 VDD.n84 3.1505
R324 VDD.n82 VDD.n81 3.1505
R325 VDD.n80 VDD.n79 3.1505
R326 VDD.n78 VDD.n77 3.1505
R327 VDD.n76 VDD.n75 3.1505
R328 VDD.n73 VDD.n72 3.1505
R329 VDD.n71 VDD.n70 3.1505
R330 VDD.n69 VDD.n68 3.1505
R331 VDD.n66 VDD.n65 3.1505
R332 VDD.n64 VDD.n63 3.1505
R333 VDD.n62 VDD.n61 3.1505
R334 VDD.n60 VDD.n59 3.1505
R335 VDD.n57 VDD.n56 3.1505
R336 VDD.n55 VDD.n54 3.1505
R337 VDD.n53 VDD.n52 3.1505
R338 VDD.n50 VDD.n49 3.1505
R339 VDD.n48 VDD.n47 3.1505
R340 VDD.n46 VDD.n45 3.1505
R341 VDD.n39 VDD.n38 3.1505
R342 VDD.n37 VDD.n36 3.1505
R343 VDD.n35 VDD.n34 3.1505
R344 VDD.n33 VDD.n32 3.1505
R345 VDD.n31 VDD.n30 3.1505
R346 VDD.n287 VDD.n286 3.1505
R347 VDD.n291 VDD.n290 3.1505
R348 VDD.n295 VDD.n294 3.1505
R349 VDD.n299 VDD.n298 3.1505
R350 VDD.n303 VDD.n302 3.1505
R351 VDD.n307 VDD.n306 3.1505
R352 VDD.n311 VDD.n310 3.1505
R353 VDD.n315 VDD.n314 3.1505
R354 VDD.n319 VDD.n318 3.1505
R355 VDD.n323 VDD.n322 3.1505
R356 VDD.n327 VDD.n326 3.1505
R357 VDD.n331 VDD.n330 3.1505
R358 VDD.n335 VDD.n334 3.1505
R359 VDD.n339 VDD.n338 3.1505
R360 VDD.n343 VDD.n342 3.1505
R361 VDD.n347 VDD.n346 3.1505
R362 VDD.n351 VDD.n350 3.1505
R363 VDD.n355 VDD.n354 3.1505
R364 VDD.n359 VDD.n358 3.1505
R365 VDD.n363 VDD.n362 3.1505
R366 VDD.n369 VDD.n366 3.1505
R367 VDD.n375 VDD.n372 3.1505
R368 VDD.n381 VDD.n378 3.1505
R369 VDD.n387 VDD.n384 3.1505
R370 VDD.n393 VDD.n390 3.1505
R371 VDD.n399 VDD.n396 3.1505
R372 VDD.n405 VDD.n402 3.1505
R373 VDD.n411 VDD.n408 3.1505
R374 VDD.n417 VDD.n414 3.1505
R375 VDD.n423 VDD.n420 3.1505
R376 VDD.n429 VDD.n426 3.1505
R377 VDD.n435 VDD.n432 3.1505
R378 VDD.n441 VDD.n438 3.1505
R379 VDD.n447 VDD.n444 3.1505
R380 VDD.n453 VDD.n450 3.1505
R381 VDD.n464 VDD.n463 3.1505
R382 VDD.n467 VDD.n464 3.1505
R383 VDD.n473 VDD.n470 3.1505
R384 VDD.n479 VDD.n476 3.1505
R385 VDD.n485 VDD.n484 3.1505
R386 VDD.n488 VDD.n485 3.1505
R387 VDD.n492 VDD.n491 3.1505
R388 VDD.n495 VDD.n492 3.1505
R389 VDD.n499 VDD.n498 3.1505
R390 VDD.n502 VDD.n499 3.1505
R391 VDD.n508 VDD.n505 3.1505
R392 VDD.n513 VDD.n512 3.1505
R393 VDD.n516 VDD.n513 3.1505
R394 VDD.n522 VDD.n519 3.1505
R395 VDD.n527 VDD.n526 3.1505
R396 VDD.n530 VDD.n527 3.1505
R397 VDD.n534 VDD.n533 3.1505
R398 VDD.n537 VDD.n534 3.1505
R399 VDD.n541 VDD.n540 3.1505
R400 VDD.n544 VDD.n541 3.1505
R401 VDD.n548 VDD.n547 3.1505
R402 VDD.n551 VDD.n548 3.1505
R403 VDD.n555 VDD.n554 3.1505
R404 VDD.n558 VDD.n555 3.1505
R405 VDD.n1081 VDD.n1080 3.1505
R406 VDD.n1084 VDD.n1081 3.1505
R407 VDD.n1074 VDD.n1073 3.1505
R408 VDD.n1077 VDD.n1074 3.1505
R409 VDD.n1067 VDD.n1066 3.1505
R410 VDD.n1070 VDD.n1067 3.1505
R411 VDD.n1060 VDD.n1059 3.1505
R412 VDD.n1063 VDD.n1060 3.1505
R413 VDD.n1055 VDD.n1052 3.1505
R414 VDD.n1046 VDD.n1045 3.1505
R415 VDD.n1049 VDD.n1046 3.1505
R416 VDD.n1039 VDD.n1038 3.1505
R417 VDD.n1042 VDD.n1039 3.1505
R418 VDD.n1032 VDD.n1031 3.1505
R419 VDD.n1035 VDD.n1032 3.1505
R420 VDD.n1027 VDD.n1024 3.1505
R421 VDD.n1018 VDD.n1017 3.1505
R422 VDD.n1021 VDD.n1018 3.1505
R423 VDD.n1011 VDD.n1010 3.1505
R424 VDD.n1014 VDD.n1011 3.1505
R425 VDD.n1004 VDD.n1003 3.1505
R426 VDD.n1007 VDD.n1004 3.1505
R427 VDD.n999 VDD.n996 3.1505
R428 VDD.n993 VDD.n990 3.1505
R429 VDD.n987 VDD.n984 3.1505
R430 VDD.n981 VDD.n978 3.1505
R431 VDD.n975 VDD.n972 3.1505
R432 VDD.n969 VDD.n966 3.1505
R433 VDD.n963 VDD.n960 3.1505
R434 VDD.n957 VDD.n954 3.1505
R435 VDD.n951 VDD.n948 3.1505
R436 VDD.n945 VDD.n944 3.1505
R437 VDD.n941 VDD.n940 3.1505
R438 VDD.n937 VDD.n936 3.1505
R439 VDD.n933 VDD.n932 3.1505
R440 VDD.n929 VDD.n928 3.1505
R441 VDD.n925 VDD.n924 3.1505
R442 VDD.n921 VDD.n920 3.1505
R443 VDD.n917 VDD.n916 3.1505
R444 VDD.n913 VDD.n912 3.1505
R445 VDD.n909 VDD.n908 3.1505
R446 VDD.n905 VDD.n904 3.1505
R447 VDD.n901 VDD.n900 3.1505
R448 VDD.n897 VDD.n896 3.1505
R449 VDD.n893 VDD.n892 3.1505
R450 VDD.n889 VDD.n888 3.1505
R451 VDD.n885 VDD.n884 3.1505
R452 VDD.n881 VDD.n880 3.1505
R453 VDD.n877 VDD.n876 3.1505
R454 VDD.n873 VDD.n872 3.1505
R455 VDD.n869 VDD.n868 3.1505
R456 VDD.n865 VDD.n864 3.1505
R457 VDD.n594 VDD.n593 3.1505
R458 VDD.n596 VDD.n595 3.1505
R459 VDD.n598 VDD.n597 3.1505
R460 VDD.n600 VDD.n599 3.1505
R461 VDD.n602 VDD.n601 3.1505
R462 VDD.n273 VDD.n272 3.1505
R463 VDD.n272 VDD.n271 3.1505
R464 VDD.n850 VDD.n849 3.1505
R465 VDD.n849 VDD.n848 3.1505
R466 VDD.n853 VDD.n852 3.1505
R467 VDD.n852 VDD.n851 3.1505
R468 VDD.n856 VDD.n855 3.1505
R469 VDD.n855 VDD.n854 3.1505
R470 VDD.n859 VDD.n858 3.1505
R471 VDD.n858 VDD.n857 3.1505
R472 VDD.n863 VDD.n862 3.1505
R473 VDD.n862 VDD.n861 3.1505
R474 VDD.n867 VDD.n866 3.1505
R475 VDD.n866 VDD.n865 3.1505
R476 VDD.n871 VDD.n870 3.1505
R477 VDD.n870 VDD.n869 3.1505
R478 VDD.n875 VDD.n874 3.1505
R479 VDD.n874 VDD.n873 3.1505
R480 VDD.n879 VDD.n878 3.1505
R481 VDD.n878 VDD.n877 3.1505
R482 VDD.n883 VDD.n882 3.1505
R483 VDD.n882 VDD.n881 3.1505
R484 VDD.n887 VDD.n886 3.1505
R485 VDD.n886 VDD.n885 3.1505
R486 VDD.n891 VDD.n890 3.1505
R487 VDD.n890 VDD.n889 3.1505
R488 VDD.n895 VDD.n894 3.1505
R489 VDD.n894 VDD.n893 3.1505
R490 VDD.n899 VDD.n898 3.1505
R491 VDD.n898 VDD.n897 3.1505
R492 VDD.n903 VDD.n902 3.1505
R493 VDD.n902 VDD.n901 3.1505
R494 VDD.n907 VDD.n906 3.1505
R495 VDD.n906 VDD.n905 3.1505
R496 VDD.n911 VDD.n910 3.1505
R497 VDD.n910 VDD.n909 3.1505
R498 VDD.n915 VDD.n914 3.1505
R499 VDD.n914 VDD.n913 3.1505
R500 VDD.n919 VDD.n918 3.1505
R501 VDD.n918 VDD.n917 3.1505
R502 VDD.n923 VDD.n922 3.1505
R503 VDD.n922 VDD.n921 3.1505
R504 VDD.n927 VDD.n926 3.1505
R505 VDD.n926 VDD.n925 3.1505
R506 VDD.n931 VDD.n930 3.1505
R507 VDD.n930 VDD.n929 3.1505
R508 VDD.n935 VDD.n934 3.1505
R509 VDD.n934 VDD.n933 3.1505
R510 VDD.n939 VDD.n938 3.1505
R511 VDD.n938 VDD.n937 3.1505
R512 VDD.n943 VDD.n942 3.1505
R513 VDD.n942 VDD.n941 3.1505
R514 VDD.n947 VDD.n946 3.1505
R515 VDD.n946 VDD.n945 3.1505
R516 VDD.n953 VDD.n952 3.1505
R517 VDD.n952 VDD.n951 3.1505
R518 VDD.n959 VDD.n958 3.1505
R519 VDD.n958 VDD.n957 3.1505
R520 VDD.n965 VDD.n964 3.1505
R521 VDD.n964 VDD.n963 3.1505
R522 VDD.n971 VDD.n970 3.1505
R523 VDD.n970 VDD.n969 3.1505
R524 VDD.n977 VDD.n976 3.1505
R525 VDD.n976 VDD.n975 3.1505
R526 VDD.n983 VDD.n982 3.1505
R527 VDD.n982 VDD.n981 3.1505
R528 VDD.n989 VDD.n988 3.1505
R529 VDD.n988 VDD.n987 3.1505
R530 VDD.n995 VDD.n994 3.1505
R531 VDD.n994 VDD.n993 3.1505
R532 VDD.n1001 VDD.n1000 3.1505
R533 VDD.n1000 VDD.n999 3.1505
R534 VDD.n1009 VDD.n1008 3.1505
R535 VDD.n1008 VDD.n1007 3.1505
R536 VDD.n1016 VDD.n1015 3.1505
R537 VDD.n1015 VDD.n1014 3.1505
R538 VDD.n1023 VDD.n1022 3.1505
R539 VDD.n1022 VDD.n1021 3.1505
R540 VDD.n1029 VDD.n1028 3.1505
R541 VDD.n1028 VDD.n1027 3.1505
R542 VDD.n1037 VDD.n1036 3.1505
R543 VDD.n1036 VDD.n1035 3.1505
R544 VDD.n1044 VDD.n1043 3.1505
R545 VDD.n1043 VDD.n1042 3.1505
R546 VDD.n1051 VDD.n1050 3.1505
R547 VDD.n1050 VDD.n1049 3.1505
R548 VDD.n1057 VDD.n1056 3.1505
R549 VDD.n1056 VDD.n1055 3.1505
R550 VDD.n1065 VDD.n1064 3.1505
R551 VDD.n1064 VDD.n1063 3.1505
R552 VDD.n1072 VDD.n1071 3.1505
R553 VDD.n1071 VDD.n1070 3.1505
R554 VDD.n1079 VDD.n1078 3.1505
R555 VDD.n1078 VDD.n1077 3.1505
R556 VDD.n1086 VDD.n1085 3.1505
R557 VDD.n1085 VDD.n1084 3.1505
R558 VDD.n560 VDD.n559 3.1505
R559 VDD.n559 VDD.n558 3.1505
R560 VDD.n553 VDD.n552 3.1505
R561 VDD.n552 VDD.n551 3.1505
R562 VDD.n546 VDD.n545 3.1505
R563 VDD.n545 VDD.n544 3.1505
R564 VDD.n539 VDD.n538 3.1505
R565 VDD.n538 VDD.n537 3.1505
R566 VDD.n532 VDD.n531 3.1505
R567 VDD.n531 VDD.n530 3.1505
R568 VDD.n524 VDD.n523 3.1505
R569 VDD.n523 VDD.n522 3.1505
R570 VDD.n518 VDD.n517 3.1505
R571 VDD.n517 VDD.n516 3.1505
R572 VDD.n510 VDD.n509 3.1505
R573 VDD.n509 VDD.n508 3.1505
R574 VDD.n504 VDD.n503 3.1505
R575 VDD.n503 VDD.n502 3.1505
R576 VDD.n497 VDD.n496 3.1505
R577 VDD.n496 VDD.n495 3.1505
R578 VDD.n490 VDD.n489 3.1505
R579 VDD.n489 VDD.n488 3.1505
R580 VDD.n481 VDD.n480 3.1505
R581 VDD.n480 VDD.n479 3.1505
R582 VDD.n475 VDD.n474 3.1505
R583 VDD.n474 VDD.n473 3.1505
R584 VDD.n469 VDD.n468 3.1505
R585 VDD.n468 VDD.n467 3.1505
R586 VDD.n455 VDD.n454 3.1505
R587 VDD.n454 VDD.n453 3.1505
R588 VDD.n449 VDD.n448 3.1505
R589 VDD.n448 VDD.n447 3.1505
R590 VDD.n443 VDD.n442 3.1505
R591 VDD.n442 VDD.n441 3.1505
R592 VDD.n437 VDD.n436 3.1505
R593 VDD.n436 VDD.n435 3.1505
R594 VDD.n431 VDD.n430 3.1505
R595 VDD.n430 VDD.n429 3.1505
R596 VDD.n425 VDD.n424 3.1505
R597 VDD.n424 VDD.n423 3.1505
R598 VDD.n419 VDD.n418 3.1505
R599 VDD.n418 VDD.n417 3.1505
R600 VDD.n413 VDD.n412 3.1505
R601 VDD.n412 VDD.n411 3.1505
R602 VDD.n407 VDD.n406 3.1505
R603 VDD.n406 VDD.n405 3.1505
R604 VDD.n401 VDD.n400 3.1505
R605 VDD.n400 VDD.n399 3.1505
R606 VDD.n395 VDD.n394 3.1505
R607 VDD.n394 VDD.n393 3.1505
R608 VDD.n389 VDD.n388 3.1505
R609 VDD.n388 VDD.n387 3.1505
R610 VDD.n383 VDD.n382 3.1505
R611 VDD.n382 VDD.n381 3.1505
R612 VDD.n377 VDD.n376 3.1505
R613 VDD.n376 VDD.n375 3.1505
R614 VDD.n371 VDD.n370 3.1505
R615 VDD.n370 VDD.n369 3.1505
R616 VDD.n365 VDD.n364 3.1505
R617 VDD.n364 VDD.n363 3.1505
R618 VDD.n361 VDD.n360 3.1505
R619 VDD.n360 VDD.n359 3.1505
R620 VDD.n357 VDD.n356 3.1505
R621 VDD.n356 VDD.n355 3.1505
R622 VDD.n353 VDD.n352 3.1505
R623 VDD.n352 VDD.n351 3.1505
R624 VDD.n349 VDD.n348 3.1505
R625 VDD.n348 VDD.n347 3.1505
R626 VDD.n345 VDD.n344 3.1505
R627 VDD.n344 VDD.n343 3.1505
R628 VDD.n341 VDD.n340 3.1505
R629 VDD.n340 VDD.n339 3.1505
R630 VDD.n337 VDD.n336 3.1505
R631 VDD.n336 VDD.n335 3.1505
R632 VDD.n333 VDD.n332 3.1505
R633 VDD.n332 VDD.n331 3.1505
R634 VDD.n329 VDD.n328 3.1505
R635 VDD.n328 VDD.n327 3.1505
R636 VDD.n325 VDD.n324 3.1505
R637 VDD.n324 VDD.n323 3.1505
R638 VDD.n321 VDD.n320 3.1505
R639 VDD.n320 VDD.n319 3.1505
R640 VDD.n317 VDD.n316 3.1505
R641 VDD.n316 VDD.n315 3.1505
R642 VDD.n313 VDD.n312 3.1505
R643 VDD.n312 VDD.n311 3.1505
R644 VDD.n309 VDD.n308 3.1505
R645 VDD.n308 VDD.n307 3.1505
R646 VDD.n305 VDD.n304 3.1505
R647 VDD.n304 VDD.n303 3.1505
R648 VDD.n301 VDD.n300 3.1505
R649 VDD.n300 VDD.n299 3.1505
R650 VDD.n297 VDD.n296 3.1505
R651 VDD.n296 VDD.n295 3.1505
R652 VDD.n293 VDD.n292 3.1505
R653 VDD.n292 VDD.n291 3.1505
R654 VDD.n289 VDD.n288 3.1505
R655 VDD.n288 VDD.n287 3.1505
R656 VDD.n285 VDD.n284 3.1505
R657 VDD.n284 VDD.n283 3.1505
R658 VDD.n282 VDD.n281 3.1505
R659 VDD.n281 VDD.n280 3.1505
R660 VDD.n279 VDD.n278 3.1505
R661 VDD.n278 VDD.n277 3.1505
R662 VDD.n276 VDD.n275 3.1505
R663 VDD.n275 VDD.n274 3.1505
R664 VDD.n270 VDD.n269 3.1505
R665 VDD.n847 VDD.n846 3.1505
R666 VDD.n323 VDD.t15 2.47065
R667 VDD.n423 VDD.t36 2.47065
R668 VDD.n1084 VDD.t7 2.47065
R669 VDD.n951 VDD.t41 2.47065
R670 VDD.n869 VDD.t26 2.47065
R671 VDD.n238 VDD.n237 2.39402
R672 VDD.n235 VDD.n234 2.39402
R673 VDD.n232 VDD.n231 2.39402
R674 VDD.n229 VDD.n228 2.39402
R675 VDD.n225 VDD.n224 2.39402
R676 VDD.n222 VDD.n221 2.39402
R677 VDD.n219 VDD.n218 2.39402
R678 VDD.n215 VDD.n214 2.39402
R679 VDD.n212 VDD.n211 2.39402
R680 VDD.n209 VDD.n208 2.39402
R681 VDD.n206 VDD.n205 2.39402
R682 VDD.n202 VDD.n201 2.39402
R683 VDD.n199 VDD.n198 2.39402
R684 VDD.n196 VDD.n195 2.39402
R685 VDD.n267 VDD.n262 1.95449
R686 VDD.n267 VDD.n263 1.95449
R687 VDD.n267 VDD.n264 1.95449
R688 VDD.n267 VDD.n265 1.95449
R689 VDD.n267 VDD.n266 1.95449
R690 VDD.n820 VDD.n819 1.73593
R691 VDD.n815 VDD.n814 1.73593
R692 VDD.n810 VDD.n809 1.73593
R693 VDD.n805 VDD.n804 1.73593
R694 VDD.n799 VDD.n798 1.73593
R695 VDD.n793 VDD.n792 1.73593
R696 VDD.n251 VDD.n249 1.73593
R697 VDD.n251 VDD.n250 1.73541
R698 VDD.n242 VDD.n241 1.41722
R699 VDD.n823 VDD.n822 1.41705
R700 VDD.n844 VDD.n828 1.41673
R701 VDD.n845 VDD.n844 1.38579
R702 VDD.n269 VDD.n268 1.37653
R703 VDD.n248 VDD.n246 1.32556
R704 VDD.n248 VDD.n247 1.3251
R705 VDD.n844 VDD.n839 1.15696
R706 VDD.n844 VDD.n829 1.15696
R707 VDD.n846 VDD.n845 1.07428
R708 VDD.n653 VDD.n652 1.07408
R709 VDD.n1 VDD.n0 1.0274
R710 VDD.n828 VDD.n827 1.0274
R711 VDD.n267 VDD.n248 0.914272
R712 VDD.n267 VDD.n261 0.888554
R713 VDD.n268 VDD.n267 0.888554
R714 VDD.n844 VDD.n843 0.709103
R715 VDD.n844 VDD.n842 0.709103
R716 VDD.n844 VDD.n841 0.709103
R717 VDD.n844 VDD.n840 0.709103
R718 VDD.n844 VDD.n838 0.709103
R719 VDD.n844 VDD.n837 0.709103
R720 VDD.n844 VDD.n836 0.709103
R721 VDD.n844 VDD.n835 0.709103
R722 VDD.n844 VDD.n834 0.709103
R723 VDD.n844 VDD.n833 0.709103
R724 VDD.n844 VDD.n832 0.709103
R725 VDD.n844 VDD.n831 0.709103
R726 VDD.n844 VDD.n830 0.709103
R727 VDD.n267 VDD.n260 0.709103
R728 VDD.n267 VDD.n259 0.709103
R729 VDD.n267 VDD.n258 0.709103
R730 VDD.n267 VDD.n257 0.709103
R731 VDD.n267 VDD.n256 0.709103
R732 VDD.n267 VDD.n255 0.709103
R733 VDD.n267 VDD.n254 0.709103
R734 VDD.n267 VDD.n253 0.709103
R735 VDD.n267 VDD.n252 0.709103
R736 VDD.n267 VDD.n251 0.709103
R737 VDD.n335 VDD.t14 0.412192
R738 VDD.n441 VDD.t28 0.412192
R739 VDD.n1063 VDD.t6 0.412192
R740 VDD.n937 VDD.t19 0.412192
R741 VDD.n857 VDD.t2 0.412192
R742 VDD.n758 VDD.n655 0.329196
R743 VDD.n860 VDD.n561 0.329196
R744 VDD.n40 VDD.n39 0.14675
R745 VDD.n273 VDD.n270 0.14675
R746 VDD.n651 VDD.n649 0.11075
R747 VDD.n649 VDD.n647 0.11075
R748 VDD.n647 VDD.n645 0.11075
R749 VDD.n645 VDD.n643 0.11075
R750 VDD.n643 VDD.n641 0.11075
R751 VDD.n641 VDD.n639 0.11075
R752 VDD.n639 VDD.n637 0.11075
R753 VDD.n637 VDD.n635 0.11075
R754 VDD.n632 VDD.n630 0.11075
R755 VDD.n630 VDD.n628 0.11075
R756 VDD.n625 VDD.n623 0.11075
R757 VDD.n623 VDD.n621 0.11075
R758 VDD.n621 VDD.n619 0.11075
R759 VDD.n616 VDD.n614 0.11075
R760 VDD.n614 VDD.n612 0.11075
R761 VDD.n609 VDD.n607 0.11075
R762 VDD.n607 VDD.n605 0.11075
R763 VDD.n605 VDD.n603 0.11075
R764 VDD.n39 VDD.n37 0.11075
R765 VDD.n37 VDD.n35 0.11075
R766 VDD.n35 VDD.n33 0.11075
R767 VDD.n33 VDD.n31 0.11075
R768 VDD.n31 VDD.n29 0.11075
R769 VDD.n29 VDD.n28 0.11075
R770 VDD.n28 VDD.n27 0.11075
R771 VDD.n27 VDD.n26 0.11075
R772 VDD.n26 VDD.n25 0.11075
R773 VDD.n25 VDD.n24 0.11075
R774 VDD.n24 VDD.n23 0.11075
R775 VDD.n23 VDD.n22 0.11075
R776 VDD.n22 VDD.n21 0.11075
R777 VDD.n21 VDD.n20 0.11075
R778 VDD.n20 VDD.n19 0.11075
R779 VDD.n19 VDD.n18 0.11075
R780 VDD.n18 VDD.n17 0.11075
R781 VDD.n17 VDD.n16 0.11075
R782 VDD.n16 VDD.n15 0.11075
R783 VDD.n15 VDD.n14 0.11075
R784 VDD.n14 VDD.n13 0.11075
R785 VDD.n13 VDD.n12 0.11075
R786 VDD.n12 VDD.n11 0.11075
R787 VDD.n11 VDD.n10 0.11075
R788 VDD.n10 VDD.n9 0.11075
R789 VDD.n9 VDD.n8 0.11075
R790 VDD.n8 VDD.n7 0.11075
R791 VDD.n7 VDD.n6 0.11075
R792 VDD.n6 VDD.n5 0.11075
R793 VDD.n5 VDD.n4 0.11075
R794 VDD.n4 VDD.n3 0.11075
R795 VDD.n3 VDD.n2 0.11075
R796 VDD.n457 VDD.n456 0.11075
R797 VDD.n458 VDD.n457 0.11075
R798 VDD.n459 VDD.n458 0.11075
R799 VDD.n460 VDD.n459 0.11075
R800 VDD.n461 VDD.n460 0.11075
R801 VDD.n462 VDD.n461 0.11075
R802 VDD.n463 VDD.n462 0.11075
R803 VDD.n483 VDD.n482 0.11075
R804 VDD.n484 VDD.n483 0.11075
R805 VDD.n512 VDD.n511 0.11075
R806 VDD.n526 VDD.n525 0.11075
R807 VDD.n1059 VDD.n1058 0.11075
R808 VDD.n1031 VDD.n1030 0.11075
R809 VDD.n1003 VDD.n1002 0.11075
R810 VDD.n565 VDD.n564 0.11075
R811 VDD.n566 VDD.n565 0.11075
R812 VDD.n567 VDD.n566 0.11075
R813 VDD.n568 VDD.n567 0.11075
R814 VDD.n569 VDD.n568 0.11075
R815 VDD.n570 VDD.n569 0.11075
R816 VDD.n571 VDD.n570 0.11075
R817 VDD.n572 VDD.n571 0.11075
R818 VDD.n573 VDD.n572 0.11075
R819 VDD.n574 VDD.n573 0.11075
R820 VDD.n575 VDD.n574 0.11075
R821 VDD.n576 VDD.n575 0.11075
R822 VDD.n577 VDD.n576 0.11075
R823 VDD.n578 VDD.n577 0.11075
R824 VDD.n579 VDD.n578 0.11075
R825 VDD.n580 VDD.n579 0.11075
R826 VDD.n581 VDD.n580 0.11075
R827 VDD.n582 VDD.n581 0.11075
R828 VDD.n583 VDD.n582 0.11075
R829 VDD.n584 VDD.n583 0.11075
R830 VDD.n585 VDD.n584 0.11075
R831 VDD.n586 VDD.n585 0.11075
R832 VDD.n587 VDD.n586 0.11075
R833 VDD.n588 VDD.n587 0.11075
R834 VDD.n589 VDD.n588 0.11075
R835 VDD.n590 VDD.n589 0.11075
R836 VDD.n591 VDD.n590 0.11075
R837 VDD.n592 VDD.n591 0.11075
R838 VDD.n594 VDD.n592 0.11075
R839 VDD.n596 VDD.n594 0.11075
R840 VDD.n598 VDD.n596 0.11075
R841 VDD.n600 VDD.n598 0.11075
R842 VDD.n602 VDD.n600 0.11075
R843 VDD.n87 VDD.n85 0.11075
R844 VDD.n82 VDD.n80 0.11075
R845 VDD.n80 VDD.n78 0.11075
R846 VDD.n78 VDD.n76 0.11075
R847 VDD.n73 VDD.n71 0.11075
R848 VDD.n71 VDD.n69 0.11075
R849 VDD.n66 VDD.n64 0.11075
R850 VDD.n64 VDD.n62 0.11075
R851 VDD.n62 VDD.n60 0.11075
R852 VDD.n57 VDD.n55 0.11075
R853 VDD.n55 VDD.n53 0.11075
R854 VDD.n50 VDD.n48 0.11075
R855 VDD.n48 VDD.n46 0.11075
R856 VDD.n43 VDD.n42 0.11075
R857 VDD.n42 VDD.n41 0.11075
R858 VDD.n826 VDD.n824 0.11075
R859 VDD.n824 VDD.n821 0.11075
R860 VDD.n821 VDD.n818 0.11075
R861 VDD.n818 VDD.n816 0.11075
R862 VDD.n816 VDD.n813 0.11075
R863 VDD.n813 VDD.n811 0.11075
R864 VDD.n811 VDD.n808 0.11075
R865 VDD.n808 VDD.n806 0.11075
R866 VDD.n802 VDD.n800 0.11075
R867 VDD.n800 VDD.n797 0.11075
R868 VDD.n794 VDD.n791 0.11075
R869 VDD.n791 VDD.n789 0.11075
R870 VDD.n789 VDD.n787 0.11075
R871 VDD.n784 VDD.n782 0.11075
R872 VDD.n782 VDD.n780 0.11075
R873 VDD.n777 VDD.n775 0.11075
R874 VDD.n775 VDD.n773 0.11075
R875 VDD.n773 VDD.n772 0.11075
R876 VDD.n245 VDD.n243 0.11075
R877 VDD.n239 VDD.n236 0.11075
R878 VDD.n236 VDD.n233 0.11075
R879 VDD.n233 VDD.n230 0.11075
R880 VDD.n226 VDD.n223 0.11075
R881 VDD.n223 VDD.n220 0.11075
R882 VDD.n216 VDD.n213 0.11075
R883 VDD.n213 VDD.n210 0.11075
R884 VDD.n210 VDD.n207 0.11075
R885 VDD.n203 VDD.n200 0.11075
R886 VDD.n200 VDD.n197 0.11075
R887 VDD.n193 VDD.n191 0.11075
R888 VDD.n191 VDD.n189 0.11075
R889 VDD.n186 VDD.n184 0.11075
R890 VDD.n184 VDD.n182 0.11075
R891 VDD.n276 VDD.n273 0.11075
R892 VDD.n279 VDD.n276 0.11075
R893 VDD.n282 VDD.n279 0.11075
R894 VDD.n285 VDD.n282 0.11075
R895 VDD.n289 VDD.n285 0.11075
R896 VDD.n293 VDD.n289 0.11075
R897 VDD.n297 VDD.n293 0.11075
R898 VDD.n301 VDD.n297 0.11075
R899 VDD.n305 VDD.n301 0.11075
R900 VDD.n309 VDD.n305 0.11075
R901 VDD.n313 VDD.n309 0.11075
R902 VDD.n317 VDD.n313 0.11075
R903 VDD.n321 VDD.n317 0.11075
R904 VDD.n325 VDD.n321 0.11075
R905 VDD.n329 VDD.n325 0.11075
R906 VDD.n333 VDD.n329 0.11075
R907 VDD.n337 VDD.n333 0.11075
R908 VDD.n341 VDD.n337 0.11075
R909 VDD.n345 VDD.n341 0.11075
R910 VDD.n349 VDD.n345 0.11075
R911 VDD.n353 VDD.n349 0.11075
R912 VDD.n357 VDD.n353 0.11075
R913 VDD.n361 VDD.n357 0.11075
R914 VDD.n365 VDD.n361 0.11075
R915 VDD.n371 VDD.n365 0.11075
R916 VDD.n377 VDD.n371 0.11075
R917 VDD.n383 VDD.n377 0.11075
R918 VDD.n389 VDD.n383 0.11075
R919 VDD.n395 VDD.n389 0.11075
R920 VDD.n401 VDD.n395 0.11075
R921 VDD.n407 VDD.n401 0.11075
R922 VDD.n413 VDD.n407 0.11075
R923 VDD.n419 VDD.n413 0.11075
R924 VDD.n425 VDD.n419 0.11075
R925 VDD.n431 VDD.n425 0.11075
R926 VDD.n437 VDD.n431 0.11075
R927 VDD.n443 VDD.n437 0.11075
R928 VDD.n449 VDD.n443 0.11075
R929 VDD.n455 VDD.n449 0.11075
R930 VDD.n469 VDD.n455 0.11075
R931 VDD.n475 VDD.n469 0.11075
R932 VDD.n481 VDD.n475 0.11075
R933 VDD.n490 VDD.n481 0.11075
R934 VDD.n497 VDD.n490 0.11075
R935 VDD.n504 VDD.n497 0.11075
R936 VDD.n510 VDD.n504 0.11075
R937 VDD.n518 VDD.n510 0.11075
R938 VDD.n524 VDD.n518 0.11075
R939 VDD.n532 VDD.n524 0.11075
R940 VDD.n539 VDD.n532 0.11075
R941 VDD.n546 VDD.n539 0.11075
R942 VDD.n553 VDD.n546 0.11075
R943 VDD.n560 VDD.n553 0.11075
R944 VDD.n1086 VDD.n1079 0.11075
R945 VDD.n1079 VDD.n1072 0.11075
R946 VDD.n1072 VDD.n1065 0.11075
R947 VDD.n1065 VDD.n1057 0.11075
R948 VDD.n1057 VDD.n1051 0.11075
R949 VDD.n1051 VDD.n1044 0.11075
R950 VDD.n1044 VDD.n1037 0.11075
R951 VDD.n1037 VDD.n1029 0.11075
R952 VDD.n1029 VDD.n1023 0.11075
R953 VDD.n1023 VDD.n1016 0.11075
R954 VDD.n1016 VDD.n1009 0.11075
R955 VDD.n1009 VDD.n1001 0.11075
R956 VDD.n1001 VDD.n995 0.11075
R957 VDD.n995 VDD.n989 0.11075
R958 VDD.n989 VDD.n983 0.11075
R959 VDD.n983 VDD.n977 0.11075
R960 VDD.n977 VDD.n971 0.11075
R961 VDD.n971 VDD.n965 0.11075
R962 VDD.n965 VDD.n959 0.11075
R963 VDD.n959 VDD.n953 0.11075
R964 VDD.n953 VDD.n947 0.11075
R965 VDD.n947 VDD.n943 0.11075
R966 VDD.n943 VDD.n939 0.11075
R967 VDD.n939 VDD.n935 0.11075
R968 VDD.n935 VDD.n931 0.11075
R969 VDD.n931 VDD.n927 0.11075
R970 VDD.n927 VDD.n923 0.11075
R971 VDD.n923 VDD.n919 0.11075
R972 VDD.n919 VDD.n915 0.11075
R973 VDD.n915 VDD.n911 0.11075
R974 VDD.n911 VDD.n907 0.11075
R975 VDD.n907 VDD.n903 0.11075
R976 VDD.n903 VDD.n899 0.11075
R977 VDD.n899 VDD.n895 0.11075
R978 VDD.n895 VDD.n891 0.11075
R979 VDD.n891 VDD.n887 0.11075
R980 VDD.n887 VDD.n883 0.11075
R981 VDD.n883 VDD.n879 0.11075
R982 VDD.n879 VDD.n875 0.11075
R983 VDD.n875 VDD.n871 0.11075
R984 VDD.n871 VDD.n867 0.11075
R985 VDD.n867 VDD.n863 0.11075
R986 VDD.n859 VDD.n856 0.11075
R987 VDD.n856 VDD.n853 0.11075
R988 VDD.n853 VDD.n850 0.11075
R989 VDD.n850 VDD.n847 0.11075
R990 VDD.n58 VDD.n57 0.109625
R991 VDD.n204 VDD.n203 0.109625
R992 VDD.n85 VDD.n83 0.104
R993 VDD.n243 VDD.n240 0.104
R994 VDD.n863 VDD.n860 0.0995
R995 VDD.n628 VDD.n626 0.096125
R996 VDD.n797 VDD.n795 0.096125
R997 VDD.n179 VDD.n89 0.089375
R998 VDD.n180 VDD.n179 0.089375
R999 VDD.n617 VDD.n616 0.08375
R1000 VDD.n785 VDD.n784 0.08375
R1001 VDD.n51 VDD.n50 0.082625
R1002 VDD.n194 VDD.n193 0.082625
R1003 VDD.n74 VDD.n73 0.0815
R1004 VDD.n227 VDD.n226 0.0815
R1005 VDD.n654 VDD.n651 0.07025
R1006 VDD.n89 VDD.n87 0.07025
R1007 VDD.n847 VDD.n826 0.07025
R1008 VDD.n270 VDD.n245 0.07025
R1009 VDD.n612 VDD.n610 0.069125
R1010 VDD.n46 VDD.n44 0.069125
R1011 VDD.n780 VDD.n778 0.069125
R1012 VDD.n189 VDD.n187 0.069125
R1013 VDD.n635 VDD.n633 0.066875
R1014 VDD.n806 VDD.n803 0.066875
R1015 VDD.n603 VDD.n602 0.06575
R1016 VDD.n41 VDD.n40 0.06575
R1017 VDD.n182 VDD.n180 0.06575
R1018 VDD.n69 VDD.n67 0.062375
R1019 VDD.n220 VDD.n217 0.062375
R1020 VDD.n771 VDD.n654 0.060125
R1021 VDD VDD.n560 0.05675
R1022 VDD VDD.n1086 0.0545
R1023 VDD.n67 VDD.n66 0.048875
R1024 VDD.n217 VDD.n216 0.048875
R1025 VDD.n633 VDD.n632 0.044375
R1026 VDD.n803 VDD.n802 0.044375
R1027 VDD.n610 VDD.n609 0.042125
R1028 VDD.n44 VDD.n43 0.042125
R1029 VDD.n778 VDD.n777 0.042125
R1030 VDD.n187 VDD.n186 0.042125
R1031 VDD.n178 VDD.n175 0.0356394
R1032 VDD.n175 VDD.n172 0.0356394
R1033 VDD.n172 VDD.n169 0.0356394
R1034 VDD.n169 VDD.n166 0.0356394
R1035 VDD.n166 VDD.n163 0.0356394
R1036 VDD.n163 VDD.n160 0.0356394
R1037 VDD.n160 VDD.n157 0.0356394
R1038 VDD.n157 VDD.n154 0.0356394
R1039 VDD.n154 VDD.n151 0.0356394
R1040 VDD.n151 VDD.n148 0.0356394
R1041 VDD.n148 VDD.n145 0.0356394
R1042 VDD.n145 VDD.n142 0.0356394
R1043 VDD.n142 VDD.n139 0.0356394
R1044 VDD.n139 VDD.n136 0.0356394
R1045 VDD.n136 VDD.n133 0.0356394
R1046 VDD.n133 VDD.n130 0.0356394
R1047 VDD.n130 VDD.n127 0.0356394
R1048 VDD.n127 VDD.n124 0.0356394
R1049 VDD.n124 VDD.n121 0.0356394
R1050 VDD.n121 VDD.n118 0.0356394
R1051 VDD.n118 VDD.n115 0.0356394
R1052 VDD.n115 VDD.n112 0.0356394
R1053 VDD.n112 VDD.n109 0.0356394
R1054 VDD.n109 VDD.n106 0.0356394
R1055 VDD.n106 VDD.n103 0.0356394
R1056 VDD.n103 VDD.n102 0.0356394
R1057 VDD.n102 VDD.n101 0.0356394
R1058 VDD.n101 VDD.n100 0.0356394
R1059 VDD.n100 VDD.n99 0.0356394
R1060 VDD.n99 VDD.n98 0.0356394
R1061 VDD.n98 VDD.n97 0.0356394
R1062 VDD.n97 VDD.n96 0.0356394
R1063 VDD.n96 VDD.n95 0.0356394
R1064 VDD.n95 VDD.n94 0.0356394
R1065 VDD.n94 VDD.n93 0.0356394
R1066 VDD.n93 VDD.n92 0.0356394
R1067 VDD.n92 VDD.n91 0.0356394
R1068 VDD.n91 VDD.n90 0.0356394
R1069 VDD.n657 VDD.n656 0.0356394
R1070 VDD.n658 VDD.n657 0.0356394
R1071 VDD.n659 VDD.n658 0.0356394
R1072 VDD.n660 VDD.n659 0.0356394
R1073 VDD.n661 VDD.n660 0.0356394
R1074 VDD.n662 VDD.n661 0.0356394
R1075 VDD.n663 VDD.n662 0.0356394
R1076 VDD.n664 VDD.n663 0.0356394
R1077 VDD.n665 VDD.n664 0.0356394
R1078 VDD.n666 VDD.n665 0.0356394
R1079 VDD.n667 VDD.n666 0.0356394
R1080 VDD.n668 VDD.n667 0.0356394
R1081 VDD.n669 VDD.n668 0.0356394
R1082 VDD.n670 VDD.n669 0.0356394
R1083 VDD.n671 VDD.n670 0.0356394
R1084 VDD.n672 VDD.n671 0.0356394
R1085 VDD.n673 VDD.n672 0.0356394
R1086 VDD.n674 VDD.n673 0.0356394
R1087 VDD.n675 VDD.n674 0.0356394
R1088 VDD.n676 VDD.n675 0.0356394
R1089 VDD.n677 VDD.n676 0.0356394
R1090 VDD.n678 VDD.n677 0.0356394
R1091 VDD.n679 VDD.n678 0.0356394
R1092 VDD.n680 VDD.n679 0.0356394
R1093 VDD.n681 VDD.n680 0.0356394
R1094 VDD.n682 VDD.n681 0.0356394
R1095 VDD.n683 VDD.n682 0.0356394
R1096 VDD.n684 VDD.n683 0.0356394
R1097 VDD.n685 VDD.n684 0.0356394
R1098 VDD.n686 VDD.n685 0.0356394
R1099 VDD.n687 VDD.n686 0.0356394
R1100 VDD.n688 VDD.n687 0.0356394
R1101 VDD.n689 VDD.n688 0.0356394
R1102 VDD.n690 VDD.n689 0.0356394
R1103 VDD.n691 VDD.n690 0.0356394
R1104 VDD.n694 VDD.n691 0.0356394
R1105 VDD.n697 VDD.n694 0.0356394
R1106 VDD.n700 VDD.n697 0.0356394
R1107 VDD.n703 VDD.n700 0.0356394
R1108 VDD.n706 VDD.n703 0.0356394
R1109 VDD.n709 VDD.n706 0.0356394
R1110 VDD.n712 VDD.n709 0.0356394
R1111 VDD.n715 VDD.n712 0.0356394
R1112 VDD.n718 VDD.n715 0.0356394
R1113 VDD.n721 VDD.n718 0.0356394
R1114 VDD.n724 VDD.n721 0.0356394
R1115 VDD.n727 VDD.n724 0.0356394
R1116 VDD.n730 VDD.n727 0.0356394
R1117 VDD.n733 VDD.n730 0.0356394
R1118 VDD.n736 VDD.n733 0.0356394
R1119 VDD.n739 VDD.n736 0.0356394
R1120 VDD.n742 VDD.n739 0.0356394
R1121 VDD.n745 VDD.n742 0.0356394
R1122 VDD.n748 VDD.n745 0.0356394
R1123 VDD.n751 VDD.n748 0.0356394
R1124 VDD.n754 VDD.n751 0.0356394
R1125 VDD.n757 VDD.n754 0.0356394
R1126 VDD.n764 VDD.n761 0.0356394
R1127 VDD.n767 VDD.n764 0.0356394
R1128 VDD.n770 VDD.n767 0.0356394
R1129 VDD.n758 VDD.n757 0.0320538
R1130 VDD.n76 VDD.n74 0.02975
R1131 VDD.n230 VDD.n227 0.02975
R1132 VDD.n53 VDD.n51 0.028625
R1133 VDD.n197 VDD.n194 0.028625
R1134 VDD.n619 VDD.n617 0.0275
R1135 VDD.n787 VDD.n785 0.0275
R1136 VDD.n179 VDD.n178 0.0187869
R1137 VDD.n771 VDD.n770 0.0166355
R1138 VDD.n626 VDD.n625 0.015125
R1139 VDD.n795 VDD.n794 0.015125
R1140 VDD.n772 VDD.n771 0.015125
R1141 VDD.n860 VDD.n859 0.01175
R1142 VDD.n83 VDD.n82 0.00725
R1143 VDD.n240 VDD.n239 0.00725
R1144 VDD.n761 VDD.n758 0.00408566
R1145 VDD.n60 VDD.n58 0.001625
R1146 VDD.n207 VDD.n204 0.001625
R1147 a_4495_2888.t0 a_4495_2888.t1 13.3663
R1148 a_3095_1282.t0 a_3095_1282.t1 12.7459
R1149 a_1695_5015.t0 a_1695_5015.t1 8.90405
R1150 a_1695_4013.t0 a_1695_4013.t1 9.02706
R1151 a_3935_5015.t0 a_3935_5015.t1 15.3118
R1152 a_4775_4363.t0 a_4775_4363.t1 13.5463
R1153 a_7295_4013.t0 a_7295_4013.t1 13.3663
R1154 a_7015_3711.t0 a_7015_3711.t1 13.3663
R1155 a_6455_2888.t0 a_6455_2888.t1 15.6157
R1156 a_5615_2236.t0 a_5615_2236.t1 13.3171
R1157 a_3375_5015.t0 a_3375_5015.t1 13.3172
R1158 a_3375_4013.t0 a_3375_4013.t1 14.6794
R1159 a_8975_2888.t0 a_8975_2888.t1 13.3663
R1160 a_7575_1282.t0 a_7575_1282.t1 12.746
R1161 G G.n13 9.93165
R1162 G.n2 G.t8 8.04282
R1163 G.n9 G.t6 7.0968
R1164 G.n13 G.t9 6.5735
R1165 G.n8 G.t7 6.5735
R1166 G.n10 G.t5 5.27519
R1167 G.n3 G.t1 5.27447
R1168 G.n9 G.t4 5.07521
R1169 G.n2 G.t0 5.07252
R1170 G.n11 G.t2 3.97325
R1171 G G.n8 3.34772
R1172 G.n7 G.t11 3.25137
R1173 G.n12 G.t3 3.21632
R1174 G.n0 G.t10 3.18852
R1175 G.n5 G.n4 2.27388
R1176 G.n11 G.n10 1.9927
R1177 G.n1 G.n0 1.56434
R1178 G.n12 G.n11 1.09431
R1179 G.n7 G.n6 1.08603
R1180 G.n4 G.n3 0.835821
R1181 G.n8 G.n7 0.45775
R1182 G.n13 G.n12 0.457326
R1183 G.n10 G.n9 0.206427
R1184 G.n3 G.n2 0.197719
R1185 G.n6 G.n1 0.0647857
R1186 G.n6 G.n5 0.0647857
R1187 a_6175_5015.t0 a_6175_5015.t1 8.90503
R1188 a_6175_4013.t0 a_6175_4013.t1 9.02698
R1189 F.n0 F.t1 8.86329
R1190 F.n1 F.t0 8.86329
R1191 F.n0 F.t2 8.402
R1192 F.n1 F.t3 8.402
R1193 F F.n0 7.18674
R1194 F F.n1 0.727136
R1195 a_8975_3711.t0 a_8975_3711.t1 13.3663
R1196 a_7295_2236.t0 a_7295_2236.t1 14.6723
R1197 a_8415_2586.t0 a_8415_2586.t1 15.3118
R1198 a_1135_5317.t0 a_1135_5317.t1 18.2801
R1199 a_1135_5015.t0 a_1135_5015.t1 15.1072
R1200 a_3655_5317.t0 a_3655_5317.t1 12.1742
R1201 a_3095_4665.t0 a_3095_4665.t1 8.90515
R1202 a_5615_5317.t0 a_5615_5317.t1 18.2801
R1203 a_5615_5015.t0 a_5615_5015.t1 15.1072
R1204 a_2815_2888.t0 a_2815_2888.t1 13.3663
R1205 a_3095_2586.t0 a_3095_2586.t1 13.8986
R1206 a_3375_4665.t0 a_3375_4665.t1 15.1072
R1207 a_3375_4363.t0 a_3375_4363.t1 15.1112
R1208 a_3935_4665.t0 a_3935_4665.t1 16.7065
R1209 a_5895_4363.t0 a_5895_4363.t1 13.3663
R1210 a_5055_2888.t0 a_5055_2888.t1 13.3663
R1211 a_4775_2586.t0 a_4775_2586.t1 13.5463
R1212 E.n5 E.t0 7.96203
R1213 E.n2 E.t1 7.96203
R1214 E E.n5 7.20855
R1215 E.n3 E.t6 6.95733
R1216 E.n0 E.t7 6.95733
R1217 E.n4 E.t3 6.42124
R1218 E.n1 E.t5 6.42124
R1219 E.n3 E.t2 6.4095
R1220 E.n0 E.t4 6.4095
R1221 E.n5 E.n4 2.55977
R1222 E.n2 E.n1 2.55977
R1223 E E.n2 0.838955
R1224 E.n4 E.n3 0.381128
R1225 E.n1 E.n0 0.381128
R1226 a_7295_2888.t0 a_7295_2888.t1 13.3663
R1227 a_7575_2586.t0 a_7575_2586.t1 13.8986
R1228 a_5335_4665.t0 a_5335_4665.t1 12.1738
R1229 a_5335_4363.t0 a_5335_4363.t1 11.2391
R1230 a_7855_4665.t0 a_7855_4665.t1 15.1072
R1231 a_7855_4363.t0 a_7855_4363.t1 15.1112
R1232 a_6735_2888.t0 a_6735_2888.t1 13.3663
R1233 a_7015_2586.t0 a_7015_2586.t1 13.3663
R1234 a_575_3711.n1 a_575_3711.t1 8.50661
R1235 a_575_3711.n0 a_575_3711.t0 6.84437
R1236 a_575_3711.t2 a_575_3711.n1 5.39199
R1237 a_575_3711.n0 a_575_3711.t3 3.14625
R1238 a_575_3711.n1 a_575_3711.n0 2.04585
R1239 a_4495_5317.t0 a_4495_5317.t1 13.3663
R1240 a_4775_5015.t0 a_4775_5015.t1 13.5463
R1241 a_6735_5317.t0 a_6735_5317.t1 13.3663
R1242 a_5335_4013.t0 a_5335_4013.t1 13.8981
R1243 a_3935_4013.t0 a_3935_4013.t1 11.2396
R1244 a_5335_2236.t0 a_5335_2236.t1 12.1742
R1245 a_6175_2586.t0 a_6175_2586.t1 8.90405
R1246 a_5615_4013.t0 a_5615_4013.t1 15.1112
R1247 a_5615_2888.t0 a_5615_2888.t1 18.2801
R1248 a_7855_2236.t0 a_7855_2236.t1 15.1072
R1249 a_8135_5317.t0 a_8135_5317.t1 12.1742
R1250 a_8415_4013.t0 a_8415_4013.t1 11.2396
R1251 a_8135_2888.t0 a_8135_2888.t1 12.1749
R1252 a_7575_2236.t0 a_7575_2236.t1 8.90503
R1253 B.n0 B.t1 7.9449
R1254 B.n1 B.t3 7.9449
R1255 B.n2 B.n1 7.78834
R1256 B.n0 B.t2 6.789
R1257 B.n1 B.t0 6.789
R1258 B.n2 B.n0 2.25045
R1259 B B.n2 0.1892
R1260 a_8135_4363.t0 a_8135_4363.t1 13.3663
R1261 a_1975_5317.t0 a_1975_5317.t1 15.6157
R1262 a_5895_5317.t0 a_5895_5317.t1 14.6731
R1263 a_5055_4665.t0 a_5055_4665.t1 15.3135
R1264 a_5055_5317.t0 a_5055_5317.t1 13.3663
R1265 a_5335_5015.t0 a_5335_5015.t1 12.7436
R1266 a_6455_5317.t0 a_6455_5317.t1 15.6157
R1267 a_7855_5015.t0 a_7855_5015.t1 13.3181
R1268 a_855_5015.t0 a_855_5015.t1 12.7437
R1269 a_3095_4363.t0 a_3095_4363.t1 9.02696
R1270 a_2815_1584.t0 a_2815_1584.t1 13.3663
R1271 a_2535_1282.t0 a_2535_1282.t1 13.3663
R1272 a_575_4665.t0 a_575_4665.t1 15.3126
R1273 A A.t0 14.9357
R1274 A A.t1 9.04183
R1275 a_7575_4665.t0 a_7575_4665.t1 8.90515
R1276 a_7575_4363.t0 a_7575_4363.t1 9.02687
R1277 a_7015_4363.t0 a_7015_4363.t1 13.3663
R1278 D.n1 D.t0 11.6419
R1279 D.n0 D.t1 11.6419
R1280 D.n0 D.t2 11.1324
R1281 D.n1 D.t3 11.1319
R1282 D D.n0 6.43542
R1283 D D.n1 0.355326
R1284 a_3095_3711.t0 a_3095_3711.t1 12.7459
R1285 a_5615_4665.t0 a_5615_4665.t1 13.3171
R1286 a_8975_5317.t0 a_8975_5317.t1 13.3663
R1287 a_7575_3711.t0 a_7575_3711.t1 12.746
R1288 a_1135_1934.t0 a_1135_1934.t1 14.6793
R1289 C.n1 C.t2 14.2686
R1290 C.n0 C.t3 14.2685
R1291 C.n0 C.t1 10.016
R1292 C.n1 C.t0 10.0155
R1293 C.n2 C.n1 4.97192
R1294 C.n3 C.n2 1.21745
R1295 C.n3 C.n0 0.501554
R1296 C C.n3 0.00595455
R1297 a_7295_4665.t0 a_7295_4665.t1 14.6723
R1298 a_8415_5015.t0 a_8415_5015.t1 15.3132
R1299 a_3935_1584.t0 a_3935_1584.t1 11.2396
R1300 a_3935_1282.t0 a_3935_1282.t1 16.5391
R1301 a_6175_4665.t0 a_6175_4665.t1 16.6921
R1302 a_7855_4013.t0 a_7855_4013.t1 14.6794
R1303 a_2815_5317.t0 a_2815_5317.t1 13.3663
R1304 a_3095_5015.t0 a_3095_5015.t1 13.8986
R1305 a_1415_2888.n2 a_1415_2888.t0 10.5962
R1306 a_1415_2888.n1 a_1415_2888.t5 10.5913
R1307 a_1415_2888.t1 a_1415_2888.n2 4.07589
R1308 a_1415_2888.n1 a_1415_2888.t3 4.07553
R1309 a_1415_2888.n0 a_1415_2888.t2 3.2869
R1310 a_1415_2888.n0 a_1415_2888.t4 3.2859
R1311 a_1415_2888.n2 a_1415_2888.n0 2.26982
R1312 a_1415_2888.n0 a_1415_2888.n1 2.25987
R1313 a_7295_5317.t0 a_7295_5317.t1 13.3663
R1314 a_7575_5015.t0 a_7575_5015.t1 13.8986
R1315 a_7015_5015.t0 a_7015_5015.t1 13.3663
R1316 a_2255_1584.t0 a_2255_1584.t1 13.3663
R1317 a_1135_2586.t0 a_1135_2586.t1 15.1072
R1318 a_1135_1584.t0 a_1135_1584.t1 15.1112
R1319 a_1415_1934.t0 a_1415_1934.t1 13.3663
R1320 a_3935_2236.t0 a_3935_2236.t1 16.7065
R1321 a_3655_1934.t0 a_3655_1934.t1 13.3663
R1322 a_1695_1584.t0 a_1695_1584.t1 9.02706
R1323 a_1695_1282.t0 a_1695_1282.t1 16.5556
R1324 a_2815_4013.t0 a_2815_4013.t1 13.3663
R1325 a_2535_3711.t0 a_2535_3711.t1 13.3663
R1326 a_3095_1934.t0 a_3095_1934.t1 9.02687
R1327 a_5615_1584.t0 a_5615_1584.t1 15.1112
R1328 a_4215_1282.t0 a_4215_1282.t1 15.3136
R1329 a_1135_4363.t0 a_1135_4363.t1 14.6793
R1330 a_3935_3711.t0 a_3935_3711.t1 16.5391
R1331 a_855_2586.t0 a_855_2586.t1 12.7437
R1332 a_4775_1584.t0 a_4775_1584.t1 13.5463
R1333 a_4495_1282.t0 a_4495_1282.t1 13.3663
R1334 a_3375_1934.t0 a_3375_1934.t1 15.1112
R1335 a_6735_1584.t0 a_6735_1584.t1 13.3663
R1336 a_5335_2586.t0 a_5335_2586.t1 12.7437
R1337 a_1695_2236.t0 a_1695_2236.t1 16.6921
R1338 a_1135_2236.t0 a_1135_2236.t1 13.3171
R1339 a_5615_1934.t0 a_5615_1934.t1 14.6793
R1340 a_2255_4013.t0 a_2255_4013.t1 13.3663
R1341 a_5335_1934.t0 a_5335_1934.t1 11.2391
R1342 a_3375_1584.t0 a_3375_1584.t1 14.6794
R1343 a_3375_1282.t0 a_3375_1282.t1 18.9537
R1344 a_7855_1584.t0 a_7855_1584.t1 14.6794
R1345 a_5335_1584.t0 a_5335_1584.t1 13.8984
R1346 a_5055_1282.t0 a_5055_1282.t1 13.3663
R1347 a_575_1282.n1 a_575_1282.t3 8.50661
R1348 a_575_1282.n0 a_575_1282.t0 6.84437
R1349 a_575_1282.t1 a_575_1282.n1 5.39199
R1350 a_575_1282.n0 a_575_1282.t2 3.14625
R1351 a_575_1282.n1 a_575_1282.n0 2.04585
R1352 a_1695_2586.t0 a_1695_2586.t1 8.90405
R1353 a_3935_2586.t0 a_3935_2586.t1 15.3118
R1354 a_4775_1934.t0 a_4775_1934.t1 13.5463
R1355 a_1695_3711.t0 a_1695_3711.t1 16.5556
R1356 a_3375_2586.t0 a_3375_2586.t1 13.3181
R1357 a_1135_4013.t0 a_1135_4013.t1 15.1112
R1358 a_6175_1584.t0 a_6175_1584.t1 9.02706
R1359 a_2535_2586.t0 a_2535_2586.t1 13.3663
R1360 a_4215_3711.t0 a_4215_3711.t1 15.3136
R1361 a_8975_1282.t0 a_8975_1282.t1 13.3663
R1362 a_8415_1584.t0 a_8415_1584.t1 11.2397
R1363 H H.t1 17.0021
R1364 H H.t0 10.2549
R1365 a_3375_2236.t0 a_3375_2236.t1 15.1072
R1366 a_5895_1934.t0 a_5895_1934.t1 13.3663
R1367 a_1975_2888.t0 a_1975_2888.t1 15.6157
R1368 a_7855_1934.t0 a_7855_1934.t1 15.1112
R1369 a_4775_4013.t0 a_4775_4013.t1 13.5463
R1370 a_4495_3711.t0 a_4495_3711.t1 13.3663
R1371 a_575_2236.t0 a_575_2236.t1 15.3126
R1372 a_6735_4013.t0 a_6735_4013.t1 13.3663
R1373 a_7295_1584.t0 a_7295_1584.t1 13.3663
R1374 a_7015_1282.t0 a_7015_1282.t1 13.3663
R1375 a_3655_2888.t0 a_3655_2888.t1 12.1749
R1376 a_5615_2586.t0 a_5615_2586.t1 15.1072
R1377 a_3375_3711.t0 a_3375_3711.t1 18.9537
R1378 a_2255_2888.t0 a_2255_2888.t1 13.3663
R1379 a_8135_1934.t0 a_8135_1934.t1 13.3663
R1380 a_1415_5317.n2 a_1415_5317.t4 10.5962
R1381 a_1415_5317.n1 a_1415_5317.t5 10.5913
R1382 a_1415_5317.t0 a_1415_5317.n2 4.07589
R1383 a_1415_5317.n1 a_1415_5317.t2 4.07553
R1384 a_1415_5317.n0 a_1415_5317.t1 3.2869
R1385 a_1415_5317.n0 a_1415_5317.t3 3.2859
R1386 a_1415_5317.n2 a_1415_5317.n0 2.26982
R1387 a_1415_5317.n0 a_1415_5317.n1 2.25987
R1388 a_5055_3711.t0 a_5055_3711.t1 13.3663
R1389 a_6175_1282.t0 a_6175_1282.t1 16.5556
R1390 a_7575_1934.t0 a_7575_1934.t1 9.02687
R1391 a_3095_2236.t0 a_3095_2236.t1 8.90503
R1392 a_5055_2236.t0 a_5055_2236.t1 15.3135
R1393 a_1135_2888.t0 a_1135_2888.t1 18.2801
R1394 a_5895_2888.t0 a_5895_2888.t1 14.6732
R1395 a_7015_1934.t0 a_7015_1934.t1 13.3663
R1396 a_1415_4363.t0 a_1415_4363.t1 13.3663
R1397 a_3655_4363.t0 a_3655_4363.t1 13.3663
R1398 a_5615_4363.t0 a_5615_4363.t1 14.6793
R1399 a_6175_2236.t0 a_6175_2236.t1 16.6921
R1400 a_7855_2586.t0 a_7855_2586.t1 13.3181
R1401 a_1135_4665.t0 a_1135_4665.t1 13.3171
R1402 a_1695_4665.t0 a_1695_4665.t1 16.6921
R1403 a_6175_3711.t0 a_6175_3711.t1 16.5556
C0 VDD G 4.58f
C1 F D 4.14f
C2 VDD A 1.83f
C3 G A 0.152f
C4 VDD B 3.87f
C5 E C 0.703f
C6 F H 2.98f
C7 D H 0.192f
C8 F VDD 1.95f
C9 VDD E 3.27f
C10 VDD D 3.59f
C11 E G 2.34f
C12 E A 3.29f
C13 VDD C 4.38f
C14 F B 0.195f
C15 G C 1.77f
C16 VDD H 2.57f
C17 A C 2.87f
C18 D B 2.58f
C19 B H 0.0426f
C20 F VSUBS 2.41f
C21 H VSUBS 4.95f
C22 B VSUBS 0.934f
C23 C VSUBS 1.32f
C24 A VSUBS 4.8f
C25 D VSUBS 2.68f
C26 G VSUBS 3.21f
C27 E VSUBS 2.94f
C28 VDD VSUBS 0.154p
C29 a_1415_5317.n0 VSUBS 0.352f
C30 a_1415_5317.t4 VSUBS 0.161f
C31 a_1415_5317.t1 VSUBS 0.0425f
C32 a_1415_5317.t5 VSUBS 0.161f
C33 a_1415_5317.t2 VSUBS 0.0629f
C34 a_1415_5317.n1 VSUBS 0.613f
C35 a_1415_5317.t3 VSUBS 0.0425f
C36 a_1415_5317.n2 VSUBS 0.603f
C37 a_1415_5317.t0 VSUBS 0.0629f
C38 H.t1 VSUBS 1.38f
C39 H.t0 VSUBS 0.444f
C40 a_1415_2888.n0 VSUBS 0.369f
C41 a_1415_2888.t0 VSUBS 0.168f
C42 a_1415_2888.t2 VSUBS 0.0445f
C43 a_1415_2888.t5 VSUBS 0.168f
C44 a_1415_2888.t3 VSUBS 0.0659f
C45 a_1415_2888.n1 VSUBS 0.642f
C46 a_1415_2888.t4 VSUBS 0.0445f
C47 a_1415_2888.n2 VSUBS 0.632f
C48 a_1415_2888.t1 VSUBS 0.0659f
C49 C.t3 VSUBS 0.643f
C50 C.t1 VSUBS 0.276f
C51 C.n0 VSUBS 1.84f
C52 C.t0 VSUBS 0.276f
C53 C.t2 VSUBS 0.643f
C54 C.n1 VSUBS 2.47f
C55 C.n2 VSUBS 0.953f
C56 C.n3 VSUBS 0.18f
C57 D.t1 VSUBS 0.615f
C58 D.t2 VSUBS 0.574f
C59 D.n0 VSUBS 3.88f
C60 D.t3 VSUBS 0.574f
C61 D.t0 VSUBS 0.615f
C62 D.n1 VSUBS 2.6f
C63 A.t1 VSUBS 0.437f
C64 A.t0 VSUBS 1.49f
C65 B.t1 VSUBS 0.247f
C66 B.t2 VSUBS 0.204f
C67 B.n0 VSUBS 1.15f
C68 B.t3 VSUBS 0.247f
C69 B.t0 VSUBS 0.204f
C70 B.n1 VSUBS 2.3f
C71 B.n2 VSUBS 2.08f
C72 E.t1 VSUBS 0.231f
C73 E.t5 VSUBS 0.169f
C74 E.t7 VSUBS 0.183f
C75 E.t4 VSUBS 0.169f
C76 E.n0 VSUBS 0.462f
C77 E.n1 VSUBS 0.644f
C78 E.n2 VSUBS 1.14f
C79 E.t3 VSUBS 0.169f
C80 E.t6 VSUBS 0.183f
C81 E.t2 VSUBS 0.169f
C82 E.n3 VSUBS 0.462f
C83 E.n4 VSUBS 0.644f
C84 E.t0 VSUBS 0.231f
C85 E.n5 VSUBS 2.42f
C86 F.t1 VSUBS 0.319f
C87 F.t2 VSUBS 0.26f
C88 F.n0 VSUBS 2.82f
C89 F.t3 VSUBS 0.26f
C90 F.t0 VSUBS 0.319f
C91 F.n1 VSUBS 1.52f
C92 G.t11 VSUBS 0.0476f
C93 G.t10 VSUBS 0.0454f
C94 G.n0 VSUBS 0.112f
C95 G.n1 VSUBS 0.0288f
C96 G.t8 VSUBS 0.269f
C97 G.t0 VSUBS 0.105f
C98 G.n2 VSUBS 0.695f
C99 G.t1 VSUBS 0.103f
C100 G.n3 VSUBS 0.336f
C101 G.n4 VSUBS 0.191f
C102 G.n5 VSUBS 0.0255f
C103 G.n6 VSUBS 0.162f
C104 G.n7 VSUBS 0.181f
C105 G.t7 VSUBS 0.0693f
C106 G.n8 VSUBS 0.337f
C107 G.t2 VSUBS 0.0676f
C108 G.t6 VSUBS 0.212f
C109 G.t4 VSUBS 0.105f
C110 G.n9 VSUBS 0.754f
C111 G.t5 VSUBS 0.103f
C112 G.n10 VSUBS 0.446f
C113 G.n11 VSUBS 0.39f
C114 G.t3 VSUBS 0.0475f
C115 G.n12 VSUBS 0.186f
C116 G.t9 VSUBS 0.0693f
C117 G.n13 VSUBS 0.825f
C118 VDD.t44 VSUBS 0.00754f
C119 VDD.t45 VSUBS 0.00754f
C120 VDD.t48 VSUBS 0.00754f
C121 VDD.t49 VSUBS 0.00754f
C122 VDD.t39 VSUBS 0.00754f
C123 VDD.t40 VSUBS 0.00754f
C124 VDD.n1 VSUBS 0.00482f
C125 VDD.t46 VSUBS 0.00754f
C126 VDD.t47 VSUBS 0.00754f
C127 VDD.t56 VSUBS 0.00754f
C128 VDD.t57 VSUBS 0.00754f
C129 VDD.t52 VSUBS 0.00754f
C130 VDD.t53 VSUBS 0.00754f
C131 VDD.n2 VSUBS 0.00352f
C132 VDD.n3 VSUBS 0.00352f
C133 VDD.n4 VSUBS 0.00352f
C134 VDD.n5 VSUBS 0.00352f
C135 VDD.n6 VSUBS 0.00352f
C136 VDD.n7 VSUBS 0.00352f
C137 VDD.n8 VSUBS 0.00352f
C138 VDD.n9 VSUBS 0.00352f
C139 VDD.n10 VSUBS 0.00352f
C140 VDD.n11 VSUBS 0.00352f
C141 VDD.n12 VSUBS 0.00352f
C142 VDD.n13 VSUBS 0.00352f
C143 VDD.n14 VSUBS 0.00352f
C144 VDD.n15 VSUBS 0.00352f
C145 VDD.n16 VSUBS 0.00352f
C146 VDD.n17 VSUBS 0.00352f
C147 VDD.n18 VSUBS 0.00352f
C148 VDD.n19 VSUBS 0.00352f
C149 VDD.n20 VSUBS 0.00352f
C150 VDD.n21 VSUBS 0.00352f
C151 VDD.n22 VSUBS 0.00352f
C152 VDD.n23 VSUBS 0.00352f
C153 VDD.n24 VSUBS 0.00352f
C154 VDD.n25 VSUBS 0.00352f
C155 VDD.n26 VSUBS 0.00352f
C156 VDD.n27 VSUBS 0.00352f
C157 VDD.n28 VSUBS 0.00352f
C158 VDD.n29 VSUBS 0.00352f
C159 VDD.n30 VSUBS 0.00352f
C160 VDD.n31 VSUBS 0.00352f
C161 VDD.n32 VSUBS 0.00352f
C162 VDD.n33 VSUBS 0.00352f
C163 VDD.n34 VSUBS 0.00352f
C164 VDD.n35 VSUBS 0.00352f
C165 VDD.n36 VSUBS 0.00352f
C166 VDD.n37 VSUBS 0.00352f
C167 VDD.n38 VSUBS 0.0041f
C168 VDD.n39 VSUBS 0.0041f
C169 VDD.n40 VSUBS 0.00482f
C170 VDD.n41 VSUBS 0.00281f
C171 VDD.n42 VSUBS 0.00352f
C172 VDD.n43 VSUBS 0.00243f
C173 VDD.n44 VSUBS 0.0141f
C174 VDD.n45 VSUBS 0.00352f
C175 VDD.n46 VSUBS 0.00286f
C176 VDD.n47 VSUBS 0.00352f
C177 VDD.n48 VSUBS 0.00352f
C178 VDD.n49 VSUBS 0.00352f
C179 VDD.n50 VSUBS 0.00308f
C180 VDD.n51 VSUBS 0.0141f
C181 VDD.n52 VSUBS 0.00352f
C182 VDD.n53 VSUBS 0.00221f
C183 VDD.n54 VSUBS 0.00352f
C184 VDD.n55 VSUBS 0.00352f
C185 VDD.n56 VSUBS 0.00352f
C186 VDD.n57 VSUBS 0.00351f
C187 VDD.n58 VSUBS 0.0141f
C188 VDD.n59 VSUBS 0.00352f
C189 VDD.n60 VSUBS 0.00178f
C190 VDD.n61 VSUBS 0.00352f
C191 VDD.n62 VSUBS 0.00352f
C192 VDD.n63 VSUBS 0.00352f
C193 VDD.n64 VSUBS 0.00352f
C194 VDD.n65 VSUBS 0.00352f
C195 VDD.n66 VSUBS 0.00254f
C196 VDD.n67 VSUBS 0.0141f
C197 VDD.n68 VSUBS 0.00352f
C198 VDD.n69 VSUBS 0.00275f
C199 VDD.n70 VSUBS 0.00352f
C200 VDD.n71 VSUBS 0.00352f
C201 VDD.n72 VSUBS 0.00352f
C202 VDD.n73 VSUBS 0.00306f
C203 VDD.n74 VSUBS 0.0141f
C204 VDD.n75 VSUBS 0.00352f
C205 VDD.n76 VSUBS 0.00223f
C206 VDD.n77 VSUBS 0.00352f
C207 VDD.n78 VSUBS 0.00352f
C208 VDD.n79 VSUBS 0.00352f
C209 VDD.n80 VSUBS 0.00352f
C210 VDD.n81 VSUBS 0.00352f
C211 VDD.n82 VSUBS 0.00187f
C212 VDD.n83 VSUBS 0.0141f
C213 VDD.n84 VSUBS 0.00352f
C214 VDD.n85 VSUBS 0.00342f
C215 VDD.n86 VSUBS 0.00288f
C216 VDD.n87 VSUBS 0.00288f
C217 VDD.n88 VSUBS 0.00489f
C218 VDD.n89 VSUBS 0.00397f
C219 VDD.n90 VSUBS 0.0111f
C220 VDD.n91 VSUBS 0.0111f
C221 VDD.n92 VSUBS 0.0111f
C222 VDD.n93 VSUBS 0.0111f
C223 VDD.n94 VSUBS 0.0111f
C224 VDD.n95 VSUBS 0.0111f
C225 VDD.n96 VSUBS 0.0111f
C226 VDD.n97 VSUBS 0.0111f
C227 VDD.n98 VSUBS 0.0111f
C228 VDD.n99 VSUBS 0.0111f
C229 VDD.n100 VSUBS 0.0111f
C230 VDD.n101 VSUBS 0.0111f
C231 VDD.n102 VSUBS 0.0111f
C232 VDD.n103 VSUBS 0.0111f
C233 VDD.n104 VSUBS 0.00352f
C234 VDD.n105 VSUBS 0.00352f
C235 VDD.n106 VSUBS 0.0111f
C236 VDD.n107 VSUBS 0.00352f
C237 VDD.n108 VSUBS 0.00352f
C238 VDD.n109 VSUBS 0.0111f
C239 VDD.n110 VSUBS 0.00352f
C240 VDD.n111 VSUBS 0.00352f
C241 VDD.n112 VSUBS 0.0111f
C242 VDD.n113 VSUBS 0.00352f
C243 VDD.n114 VSUBS 0.00352f
C244 VDD.n115 VSUBS 0.0111f
C245 VDD.n116 VSUBS 0.00352f
C246 VDD.n117 VSUBS 0.00352f
C247 VDD.n118 VSUBS 0.0111f
C248 VDD.n119 VSUBS 0.00352f
C249 VDD.n120 VSUBS 0.00352f
C250 VDD.n121 VSUBS 0.0111f
C251 VDD.n122 VSUBS 0.00352f
C252 VDD.n123 VSUBS 0.00352f
C253 VDD.n124 VSUBS 0.0111f
C254 VDD.n125 VSUBS 0.00352f
C255 VDD.n126 VSUBS 0.00352f
C256 VDD.n127 VSUBS 0.0111f
C257 VDD.n128 VSUBS 0.00352f
C258 VDD.n129 VSUBS 0.00352f
C259 VDD.n130 VSUBS 0.0111f
C260 VDD.n131 VSUBS 0.00352f
C261 VDD.n132 VSUBS 0.00352f
C262 VDD.n133 VSUBS 0.0111f
C263 VDD.n134 VSUBS 0.00352f
C264 VDD.n135 VSUBS 0.00352f
C265 VDD.n136 VSUBS 0.0111f
C266 VDD.n137 VSUBS 0.00352f
C267 VDD.n138 VSUBS 0.00352f
C268 VDD.n139 VSUBS 0.0111f
C269 VDD.n140 VSUBS 0.00352f
C270 VDD.n141 VSUBS 0.00352f
C271 VDD.n142 VSUBS 0.0111f
C272 VDD.n143 VSUBS 0.00352f
C273 VDD.n144 VSUBS 0.00352f
C274 VDD.n145 VSUBS 0.0111f
C275 VDD.n146 VSUBS 0.00352f
C276 VDD.n147 VSUBS 0.00352f
C277 VDD.n148 VSUBS 0.0111f
C278 VDD.n149 VSUBS 0.00352f
C279 VDD.n150 VSUBS 0.00352f
C280 VDD.n151 VSUBS 0.0111f
C281 VDD.n152 VSUBS 0.00352f
C282 VDD.n153 VSUBS 0.00352f
C283 VDD.n154 VSUBS 0.0111f
C284 VDD.n155 VSUBS 0.00352f
C285 VDD.n156 VSUBS 0.00352f
C286 VDD.n157 VSUBS 0.0111f
C287 VDD.n158 VSUBS 0.00352f
C288 VDD.n159 VSUBS 0.00352f
C289 VDD.n160 VSUBS 0.0111f
C290 VDD.n161 VSUBS 0.00352f
C291 VDD.n162 VSUBS 0.00352f
C292 VDD.n163 VSUBS 0.0111f
C293 VDD.n164 VSUBS 0.00352f
C294 VDD.n165 VSUBS 0.00352f
C295 VDD.n166 VSUBS 0.0111f
C296 VDD.n167 VSUBS 0.00352f
C297 VDD.n168 VSUBS 0.00352f
C298 VDD.n169 VSUBS 0.0111f
C299 VDD.n170 VSUBS 0.00352f
C300 VDD.n171 VSUBS 0.00352f
C301 VDD.n172 VSUBS 0.0111f
C302 VDD.n173 VSUBS 0.00352f
C303 VDD.n174 VSUBS 0.00352f
C304 VDD.n175 VSUBS 0.0111f
C305 VDD.n176 VSUBS 0.0041f
C306 VDD.n177 VSUBS 0.0041f
C307 VDD.n178 VSUBS 0.00841f
C308 VDD.n179 VSUBS 0.00572f
C309 VDD.n180 VSUBS 0.0039f
C310 VDD.n181 VSUBS 0.00281f
C311 VDD.n182 VSUBS 0.00281f
C312 VDD.n183 VSUBS 0.00352f
C313 VDD.n184 VSUBS 0.00352f
C314 VDD.n185 VSUBS 0.00352f
C315 VDD.n186 VSUBS 0.00243f
C316 VDD.n187 VSUBS 0.0141f
C317 VDD.n188 VSUBS 0.00352f
C318 VDD.n189 VSUBS 0.00286f
C319 VDD.n190 VSUBS 0.00352f
C320 VDD.n191 VSUBS 0.00352f
C321 VDD.n192 VSUBS 0.00352f
C322 VDD.n193 VSUBS 0.00308f
C323 VDD.n194 VSUBS 0.0141f
C324 VDD.n196 VSUBS 0.00352f
C325 VDD.n197 VSUBS 0.00221f
C326 VDD.n199 VSUBS 0.00352f
C327 VDD.n200 VSUBS 0.00352f
C328 VDD.n202 VSUBS 0.00352f
C329 VDD.n203 VSUBS 0.00351f
C330 VDD.n204 VSUBS 0.0141f
C331 VDD.n206 VSUBS 0.00352f
C332 VDD.n207 VSUBS 0.00178f
C333 VDD.n209 VSUBS 0.00352f
C334 VDD.n210 VSUBS 0.00352f
C335 VDD.n212 VSUBS 0.00352f
C336 VDD.n213 VSUBS 0.00352f
C337 VDD.n215 VSUBS 0.00352f
C338 VDD.n216 VSUBS 0.00254f
C339 VDD.n217 VSUBS 0.0141f
C340 VDD.n219 VSUBS 0.00352f
C341 VDD.n220 VSUBS 0.00275f
C342 VDD.n222 VSUBS 0.00352f
C343 VDD.n223 VSUBS 0.00352f
C344 VDD.n225 VSUBS 0.00352f
C345 VDD.n226 VSUBS 0.00306f
C346 VDD.n227 VSUBS 0.0141f
C347 VDD.n229 VSUBS 0.00352f
C348 VDD.n230 VSUBS 0.00223f
C349 VDD.n232 VSUBS 0.00352f
C350 VDD.n233 VSUBS 0.00352f
C351 VDD.n235 VSUBS 0.00352f
C352 VDD.n236 VSUBS 0.00352f
C353 VDD.n238 VSUBS 0.00352f
C354 VDD.n239 VSUBS 0.00187f
C355 VDD.n240 VSUBS 0.0141f
C356 VDD.n242 VSUBS 0.00352f
C357 VDD.n243 VSUBS 0.00342f
C358 VDD.n244 VSUBS 0.00288f
C359 VDD.n245 VSUBS 0.00288f
C360 VDD.n246 VSUBS 0.00281f
C361 VDD.n247 VSUBS 0.00482f
C362 VDD.n249 VSUBS 0.00352f
C363 VDD.n250 VSUBS 0.00352f
C364 VDD.n267 VSUBS 0.339f
C365 VDD.n269 VSUBS 0.00489f
C366 VDD.n270 VSUBS 0.00489f
C367 VDD.n271 VSUBS 0.249f
C368 VDD.n272 VSUBS 0.0041f
C369 VDD.n273 VSUBS 0.0041f
C370 VDD.n274 VSUBS 0.214f
C371 VDD.n275 VSUBS 0.00352f
C372 VDD.n276 VSUBS 0.00352f
C373 VDD.n277 VSUBS 0.181f
C374 VDD.n278 VSUBS 0.00352f
C375 VDD.n279 VSUBS 0.00352f
C376 VDD.t38 VSUBS 0.107f
C377 VDD.n280 VSUBS 0.14f
C378 VDD.n281 VSUBS 0.00352f
C379 VDD.n282 VSUBS 0.00352f
C380 VDD.n283 VSUBS 0.214f
C381 VDD.n284 VSUBS 0.00352f
C382 VDD.n285 VSUBS 0.00352f
C383 VDD.n286 VSUBS 0.00352f
C384 VDD.n287 VSUBS 0.166f
C385 VDD.n288 VSUBS 0.00352f
C386 VDD.n289 VSUBS 0.00352f
C387 VDD.t5 VSUBS 0.107f
C388 VDD.n290 VSUBS 0.00352f
C389 VDD.n291 VSUBS 0.155f
C390 VDD.n292 VSUBS 0.00352f
C391 VDD.n293 VSUBS 0.00352f
C392 VDD.n294 VSUBS 0.00352f
C393 VDD.n295 VSUBS 0.214f
C394 VDD.n296 VSUBS 0.00352f
C395 VDD.n297 VSUBS 0.00352f
C396 VDD.t0 VSUBS 0.107f
C397 VDD.n298 VSUBS 0.00352f
C398 VDD.n299 VSUBS 0.151f
C399 VDD.n300 VSUBS 0.00352f
C400 VDD.n301 VSUBS 0.00352f
C401 VDD.n302 VSUBS 0.00352f
C402 VDD.n303 VSUBS 0.17f
C403 VDD.n304 VSUBS 0.00352f
C404 VDD.n305 VSUBS 0.00352f
C405 VDD.n306 VSUBS 0.00352f
C406 VDD.n307 VSUBS 0.214f
C407 VDD.n308 VSUBS 0.00352f
C408 VDD.n309 VSUBS 0.00352f
C409 VDD.t24 VSUBS 0.107f
C410 VDD.n310 VSUBS 0.00352f
C411 VDD.n311 VSUBS 0.135f
C412 VDD.n312 VSUBS 0.00352f
C413 VDD.n313 VSUBS 0.00352f
C414 VDD.n314 VSUBS 0.00352f
C415 VDD.n315 VSUBS 0.186f
C416 VDD.n316 VSUBS 0.00352f
C417 VDD.n317 VSUBS 0.00352f
C418 VDD.n318 VSUBS 0.00352f
C419 VDD.n319 VSUBS 0.214f
C420 VDD.n320 VSUBS 0.00352f
C421 VDD.n321 VSUBS 0.00352f
C422 VDD.t15 VSUBS 0.107f
C423 VDD.n322 VSUBS 0.00352f
C424 VDD.n323 VSUBS 0.12f
C425 VDD.n324 VSUBS 0.00352f
C426 VDD.n325 VSUBS 0.00352f
C427 VDD.n326 VSUBS 0.00352f
C428 VDD.n327 VSUBS 0.201f
C429 VDD.n328 VSUBS 0.00352f
C430 VDD.n329 VSUBS 0.00352f
C431 VDD.n330 VSUBS 0.00352f
C432 VDD.n331 VSUBS 0.212f
C433 VDD.n332 VSUBS 0.00352f
C434 VDD.n333 VSUBS 0.00352f
C435 VDD.t14 VSUBS 0.107f
C436 VDD.n334 VSUBS 0.00352f
C437 VDD.n335 VSUBS 0.109f
C438 VDD.n336 VSUBS 0.00352f
C439 VDD.n337 VSUBS 0.00352f
C440 VDD.n338 VSUBS 0.00352f
C441 VDD.n339 VSUBS 0.214f
C442 VDD.n340 VSUBS 0.00352f
C443 VDD.n341 VSUBS 0.00352f
C444 VDD.n342 VSUBS 0.00352f
C445 VDD.n343 VSUBS 0.197f
C446 VDD.n344 VSUBS 0.00352f
C447 VDD.n345 VSUBS 0.00352f
C448 VDD.t43 VSUBS 0.107f
C449 VDD.n346 VSUBS 0.00352f
C450 VDD.n347 VSUBS 0.124f
C451 VDD.n348 VSUBS 0.00352f
C452 VDD.n349 VSUBS 0.00352f
C453 VDD.n350 VSUBS 0.00352f
C454 VDD.n351 VSUBS 0.214f
C455 VDD.n352 VSUBS 0.00352f
C456 VDD.n353 VSUBS 0.00352f
C457 VDD.n354 VSUBS 0.00352f
C458 VDD.n355 VSUBS 0.181f
C459 VDD.n356 VSUBS 0.00352f
C460 VDD.n357 VSUBS 0.00352f
C461 VDD.t16 VSUBS 0.107f
C462 VDD.n358 VSUBS 0.00352f
C463 VDD.n359 VSUBS 0.14f
C464 VDD.n360 VSUBS 0.00352f
C465 VDD.n361 VSUBS 0.00352f
C466 VDD.n362 VSUBS 0.00352f
C467 VDD.n363 VSUBS 0.214f
C468 VDD.n364 VSUBS 0.00352f
C469 VDD.n365 VSUBS 0.00352f
C470 VDD.n366 VSUBS 0.00352f
C471 VDD.n367 VSUBS 0.00352f
C472 VDD.n368 VSUBS 0.00352f
C473 VDD.n369 VSUBS 0.166f
C474 VDD.n370 VSUBS 0.00352f
C475 VDD.n371 VSUBS 0.00352f
C476 VDD.t37 VSUBS 0.107f
C477 VDD.n372 VSUBS 0.00352f
C478 VDD.n373 VSUBS 0.00352f
C479 VDD.n374 VSUBS 0.00352f
C480 VDD.n375 VSUBS 0.155f
C481 VDD.n376 VSUBS 0.00352f
C482 VDD.n377 VSUBS 0.00352f
C483 VDD.n378 VSUBS 0.00352f
C484 VDD.n379 VSUBS 0.00352f
C485 VDD.n380 VSUBS 0.00352f
C486 VDD.n381 VSUBS 0.214f
C487 VDD.n382 VSUBS 0.00352f
C488 VDD.n383 VSUBS 0.00352f
C489 VDD.t32 VSUBS 0.107f
C490 VDD.n384 VSUBS 0.00352f
C491 VDD.n385 VSUBS 0.00352f
C492 VDD.n386 VSUBS 0.00352f
C493 VDD.n387 VSUBS 0.151f
C494 VDD.n388 VSUBS 0.00352f
C495 VDD.n389 VSUBS 0.00352f
C496 VDD.n390 VSUBS 0.00352f
C497 VDD.n391 VSUBS 0.00352f
C498 VDD.n392 VSUBS 0.00352f
C499 VDD.n393 VSUBS 0.17f
C500 VDD.n394 VSUBS 0.00352f
C501 VDD.n395 VSUBS 0.00352f
C502 VDD.n396 VSUBS 0.00352f
C503 VDD.n397 VSUBS 0.00352f
C504 VDD.n398 VSUBS 0.00352f
C505 VDD.n399 VSUBS 0.214f
C506 VDD.n400 VSUBS 0.00352f
C507 VDD.n401 VSUBS 0.00352f
C508 VDD.t10 VSUBS 0.107f
C509 VDD.n402 VSUBS 0.00352f
C510 VDD.n403 VSUBS 0.00352f
C511 VDD.n404 VSUBS 0.00352f
C512 VDD.n405 VSUBS 0.135f
C513 VDD.n406 VSUBS 0.00352f
C514 VDD.n407 VSUBS 0.00352f
C515 VDD.n408 VSUBS 0.00352f
C516 VDD.n409 VSUBS 0.00352f
C517 VDD.n410 VSUBS 0.00352f
C518 VDD.n411 VSUBS 0.186f
C519 VDD.n412 VSUBS 0.00352f
C520 VDD.n413 VSUBS 0.00352f
C521 VDD.n414 VSUBS 0.00352f
C522 VDD.n415 VSUBS 0.00352f
C523 VDD.n416 VSUBS 0.00352f
C524 VDD.n417 VSUBS 0.214f
C525 VDD.n418 VSUBS 0.00352f
C526 VDD.n419 VSUBS 0.00352f
C527 VDD.t36 VSUBS 0.107f
C528 VDD.n420 VSUBS 0.00352f
C529 VDD.n421 VSUBS 0.00352f
C530 VDD.n422 VSUBS 0.00352f
C531 VDD.n423 VSUBS 0.12f
C532 VDD.n424 VSUBS 0.00352f
C533 VDD.n425 VSUBS 0.00352f
C534 VDD.n426 VSUBS 0.00352f
C535 VDD.n427 VSUBS 0.00352f
C536 VDD.n428 VSUBS 0.00352f
C537 VDD.n429 VSUBS 0.201f
C538 VDD.n430 VSUBS 0.00352f
C539 VDD.n431 VSUBS 0.00352f
C540 VDD.n432 VSUBS 0.00352f
C541 VDD.n433 VSUBS 0.00352f
C542 VDD.n434 VSUBS 0.00352f
C543 VDD.n435 VSUBS 0.212f
C544 VDD.n436 VSUBS 0.00352f
C545 VDD.n437 VSUBS 0.00352f
C546 VDD.t28 VSUBS 0.107f
C547 VDD.n438 VSUBS 0.00352f
C548 VDD.n439 VSUBS 0.00352f
C549 VDD.n440 VSUBS 0.00352f
C550 VDD.n441 VSUBS 0.109f
C551 VDD.n442 VSUBS 0.00352f
C552 VDD.n443 VSUBS 0.00352f
C553 VDD.n444 VSUBS 0.00352f
C554 VDD.n445 VSUBS 0.00352f
C555 VDD.n446 VSUBS 0.00352f
C556 VDD.n447 VSUBS 0.214f
C557 VDD.n448 VSUBS 0.00352f
C558 VDD.n449 VSUBS 0.00352f
C559 VDD.n450 VSUBS 0.00352f
C560 VDD.n451 VSUBS 0.00352f
C561 VDD.n452 VSUBS 0.00352f
C562 VDD.n453 VSUBS 0.197f
C563 VDD.n454 VSUBS 0.00352f
C564 VDD.n455 VSUBS 0.00352f
C565 VDD.t31 VSUBS 0.107f
C566 VDD.n456 VSUBS 0.00352f
C567 VDD.n457 VSUBS 0.00352f
C568 VDD.n458 VSUBS 0.00352f
C569 VDD.n459 VSUBS 0.00352f
C570 VDD.n460 VSUBS 0.00352f
C571 VDD.n461 VSUBS 0.00352f
C572 VDD.n462 VSUBS 0.00352f
C573 VDD.n463 VSUBS 0.00352f
C574 VDD.n464 VSUBS 0.00352f
C575 VDD.n465 VSUBS 0.00352f
C576 VDD.n466 VSUBS 0.00352f
C577 VDD.n467 VSUBS 0.124f
C578 VDD.n468 VSUBS 0.00352f
C579 VDD.n469 VSUBS 0.00352f
C580 VDD.n470 VSUBS 0.00352f
C581 VDD.n471 VSUBS 0.00352f
C582 VDD.n472 VSUBS 0.00352f
C583 VDD.n473 VSUBS 0.214f
C584 VDD.n474 VSUBS 0.00352f
C585 VDD.n475 VSUBS 0.00352f
C586 VDD.n476 VSUBS 0.00352f
C587 VDD.n477 VSUBS 0.00352f
C588 VDD.n478 VSUBS 0.00352f
C589 VDD.n479 VSUBS 0.181f
C590 VDD.n480 VSUBS 0.00352f
C591 VDD.n481 VSUBS 0.00352f
C592 VDD.t35 VSUBS 0.107f
C593 VDD.n482 VSUBS 0.00352f
C594 VDD.n483 VSUBS 0.00352f
C595 VDD.n484 VSUBS 0.00352f
C596 VDD.n485 VSUBS 0.00352f
C597 VDD.n486 VSUBS 0.00352f
C598 VDD.n487 VSUBS 0.00352f
C599 VDD.n488 VSUBS 0.14f
C600 VDD.n489 VSUBS 0.00352f
C601 VDD.n490 VSUBS 0.00352f
C602 VDD.n491 VSUBS 0.00352f
C603 VDD.n492 VSUBS 0.00352f
C604 VDD.n493 VSUBS 0.00352f
C605 VDD.n494 VSUBS 0.00352f
C606 VDD.n495 VSUBS 0.214f
C607 VDD.n496 VSUBS 0.00352f
C608 VDD.n497 VSUBS 0.00352f
C609 VDD.n498 VSUBS 0.00352f
C610 VDD.n499 VSUBS 0.00352f
C611 VDD.n500 VSUBS 0.00352f
C612 VDD.n501 VSUBS 0.00352f
C613 VDD.n502 VSUBS 0.166f
C614 VDD.n503 VSUBS 0.00352f
C615 VDD.n504 VSUBS 0.00352f
C616 VDD.t21 VSUBS 0.107f
C617 VDD.n505 VSUBS 0.00352f
C618 VDD.n506 VSUBS 0.00352f
C619 VDD.n507 VSUBS 0.00352f
C620 VDD.n508 VSUBS 0.155f
C621 VDD.n509 VSUBS 0.00352f
C622 VDD.n510 VSUBS 0.00352f
C623 VDD.n511 VSUBS 0.00352f
C624 VDD.n512 VSUBS 0.00352f
C625 VDD.n513 VSUBS 0.00352f
C626 VDD.n514 VSUBS 0.00352f
C627 VDD.n515 VSUBS 0.00352f
C628 VDD.n516 VSUBS 0.214f
C629 VDD.n517 VSUBS 0.00352f
C630 VDD.n518 VSUBS 0.00352f
C631 VDD.t13 VSUBS 0.107f
C632 VDD.n519 VSUBS 0.00352f
C633 VDD.n520 VSUBS 0.00352f
C634 VDD.n521 VSUBS 0.00352f
C635 VDD.n522 VSUBS 0.151f
C636 VDD.n523 VSUBS 0.00352f
C637 VDD.n524 VSUBS 0.00352f
C638 VDD.n525 VSUBS 0.00352f
C639 VDD.n526 VSUBS 0.00352f
C640 VDD.n527 VSUBS 0.00352f
C641 VDD.n528 VSUBS 0.00352f
C642 VDD.n529 VSUBS 0.00352f
C643 VDD.n530 VSUBS 0.17f
C644 VDD.n531 VSUBS 0.00352f
C645 VDD.n532 VSUBS 0.00352f
C646 VDD.n533 VSUBS 0.00352f
C647 VDD.n534 VSUBS 0.00352f
C648 VDD.n535 VSUBS 0.00352f
C649 VDD.n536 VSUBS 0.00352f
C650 VDD.n537 VSUBS 0.214f
C651 VDD.n538 VSUBS 0.00352f
C652 VDD.n539 VSUBS 0.00352f
C653 VDD.t9 VSUBS 0.107f
C654 VDD.n540 VSUBS 0.00352f
C655 VDD.n541 VSUBS 0.00352f
C656 VDD.n542 VSUBS 0.00352f
C657 VDD.n543 VSUBS 0.00352f
C658 VDD.n544 VSUBS 0.135f
C659 VDD.n545 VSUBS 0.00352f
C660 VDD.n546 VSUBS 0.00352f
C661 VDD.n547 VSUBS 0.00352f
C662 VDD.n548 VSUBS 0.00352f
C663 VDD.n549 VSUBS 0.00352f
C664 VDD.n550 VSUBS 0.00352f
C665 VDD.n551 VSUBS 0.186f
C666 VDD.n552 VSUBS 0.00352f
C667 VDD.n553 VSUBS 0.00352f
C668 VDD.n554 VSUBS 0.00352f
C669 VDD.n555 VSUBS 0.00352f
C670 VDD.n556 VSUBS 0.00352f
C671 VDD.n557 VSUBS 0.00352f
C672 VDD.n558 VSUBS 0.214f
C673 VDD.n559 VSUBS 0.00352f
C674 VDD.n560 VSUBS 0.00266f
C675 VDD.t22 VSUBS 0.00684f
C676 VDD.t23 VSUBS 0.00719f
C677 VDD.n561 VSUBS 0.014f
C678 VDD.t17 VSUBS 0.0075f
C679 VDD.t18 VSUBS 0.0075f
C680 VDD.t50 VSUBS 0.00761f
C681 VDD.t51 VSUBS 0.00754f
C682 VDD.n562 VSUBS 0.00281f
C683 VDD.n563 VSUBS 0.00424f
C684 VDD.t11 VSUBS 0.0075f
C685 VDD.t12 VSUBS 0.0075f
C686 VDD.t54 VSUBS 0.00761f
C687 VDD.t55 VSUBS 0.00754f
C688 VDD.n564 VSUBS 0.00352f
C689 VDD.n565 VSUBS 0.00352f
C690 VDD.n566 VSUBS 0.00352f
C691 VDD.n567 VSUBS 0.00352f
C692 VDD.n568 VSUBS 0.00352f
C693 VDD.n569 VSUBS 0.00352f
C694 VDD.n570 VSUBS 0.00352f
C695 VDD.n571 VSUBS 0.00352f
C696 VDD.n572 VSUBS 0.00352f
C697 VDD.n573 VSUBS 0.00352f
C698 VDD.n574 VSUBS 0.00352f
C699 VDD.n575 VSUBS 0.00352f
C700 VDD.n576 VSUBS 0.00352f
C701 VDD.n577 VSUBS 0.00352f
C702 VDD.n578 VSUBS 0.00352f
C703 VDD.n579 VSUBS 0.00352f
C704 VDD.n580 VSUBS 0.00352f
C705 VDD.n581 VSUBS 0.00352f
C706 VDD.n582 VSUBS 0.00352f
C707 VDD.n583 VSUBS 0.00352f
C708 VDD.n584 VSUBS 0.00352f
C709 VDD.n585 VSUBS 0.00352f
C710 VDD.n586 VSUBS 0.00352f
C711 VDD.n587 VSUBS 0.00352f
C712 VDD.n588 VSUBS 0.00352f
C713 VDD.n589 VSUBS 0.00352f
C714 VDD.n590 VSUBS 0.00352f
C715 VDD.n591 VSUBS 0.00352f
C716 VDD.n592 VSUBS 0.00352f
C717 VDD.n593 VSUBS 0.00352f
C718 VDD.n594 VSUBS 0.00352f
C719 VDD.n595 VSUBS 0.00352f
C720 VDD.n596 VSUBS 0.00352f
C721 VDD.n597 VSUBS 0.00352f
C722 VDD.n598 VSUBS 0.00352f
C723 VDD.n599 VSUBS 0.00352f
C724 VDD.n600 VSUBS 0.00352f
C725 VDD.n601 VSUBS 0.00352f
C726 VDD.n602 VSUBS 0.00281f
C727 VDD.n603 VSUBS 0.00424f
C728 VDD.n604 VSUBS 0.00281f
C729 VDD.n605 VSUBS 0.00352f
C730 VDD.n606 VSUBS 0.00352f
C731 VDD.n607 VSUBS 0.00352f
C732 VDD.n608 VSUBS 0.00352f
C733 VDD.n609 VSUBS 0.00243f
C734 VDD.n610 VSUBS 0.0142f
C735 VDD.n611 VSUBS 0.00352f
C736 VDD.n612 VSUBS 0.00286f
C737 VDD.n613 VSUBS 0.00352f
C738 VDD.n614 VSUBS 0.00352f
C739 VDD.n615 VSUBS 0.00352f
C740 VDD.n616 VSUBS 0.00309f
C741 VDD.n617 VSUBS 0.0128f
C742 VDD.n618 VSUBS 0.00352f
C743 VDD.n619 VSUBS 0.00219f
C744 VDD.n620 VSUBS 0.00352f
C745 VDD.n621 VSUBS 0.00352f
C746 VDD.n622 VSUBS 0.00352f
C747 VDD.n623 VSUBS 0.00352f
C748 VDD.n624 VSUBS 0.00352f
C749 VDD.n625 VSUBS 0.002f
C750 VDD.n626 VSUBS 0.0156f
C751 VDD.n627 VSUBS 0.00352f
C752 VDD.n628 VSUBS 0.00329f
C753 VDD.n629 VSUBS 0.00352f
C754 VDD.n630 VSUBS 0.00352f
C755 VDD.n631 VSUBS 0.00352f
C756 VDD.n632 VSUBS 0.00246f
C757 VDD.n633 VSUBS 0.0155f
C758 VDD.n634 VSUBS 0.00352f
C759 VDD.n635 VSUBS 0.00282f
C760 VDD.n636 VSUBS 0.00352f
C761 VDD.n637 VSUBS 0.00352f
C762 VDD.n638 VSUBS 0.00352f
C763 VDD.n639 VSUBS 0.00352f
C764 VDD.n640 VSUBS 0.00352f
C765 VDD.n641 VSUBS 0.00352f
C766 VDD.n642 VSUBS 0.00352f
C767 VDD.n643 VSUBS 0.00352f
C768 VDD.n644 VSUBS 0.00352f
C769 VDD.n645 VSUBS 0.00352f
C770 VDD.n646 VSUBS 0.00352f
C771 VDD.n647 VSUBS 0.00352f
C772 VDD.n648 VSUBS 0.00352f
C773 VDD.n649 VSUBS 0.00352f
C774 VDD.n650 VSUBS 0.00288f
C775 VDD.n651 VSUBS 0.00288f
C776 VDD.n653 VSUBS 0.00432f
C777 VDD.n654 VSUBS 0.00351f
C778 VDD.t3 VSUBS 0.00684f
C779 VDD.t4 VSUBS 0.00719f
C780 VDD.n655 VSUBS 0.014f
C781 VDD.n656 VSUBS 0.0111f
C782 VDD.n657 VSUBS 0.0111f
C783 VDD.n658 VSUBS 0.0111f
C784 VDD.n659 VSUBS 0.0111f
C785 VDD.n660 VSUBS 0.0111f
C786 VDD.n661 VSUBS 0.0111f
C787 VDD.n662 VSUBS 0.0111f
C788 VDD.n663 VSUBS 0.0111f
C789 VDD.n664 VSUBS 0.0111f
C790 VDD.n665 VSUBS 0.0111f
C791 VDD.n666 VSUBS 0.0111f
C792 VDD.n667 VSUBS 0.0111f
C793 VDD.n668 VSUBS 0.0111f
C794 VDD.n669 VSUBS 0.0111f
C795 VDD.n670 VSUBS 0.0111f
C796 VDD.n671 VSUBS 0.0111f
C797 VDD.n672 VSUBS 0.0111f
C798 VDD.n673 VSUBS 0.0111f
C799 VDD.n674 VSUBS 0.0111f
C800 VDD.n675 VSUBS 0.0111f
C801 VDD.n676 VSUBS 0.0111f
C802 VDD.n677 VSUBS 0.0111f
C803 VDD.n678 VSUBS 0.0111f
C804 VDD.n679 VSUBS 0.0111f
C805 VDD.n680 VSUBS 0.0111f
C806 VDD.n681 VSUBS 0.0111f
C807 VDD.n682 VSUBS 0.0111f
C808 VDD.n683 VSUBS 0.0111f
C809 VDD.n684 VSUBS 0.0111f
C810 VDD.n685 VSUBS 0.0111f
C811 VDD.n686 VSUBS 0.0111f
C812 VDD.n687 VSUBS 0.0111f
C813 VDD.n688 VSUBS 0.0111f
C814 VDD.n689 VSUBS 0.0111f
C815 VDD.n690 VSUBS 0.0111f
C816 VDD.n691 VSUBS 0.0111f
C817 VDD.n692 VSUBS 0.00352f
C818 VDD.n693 VSUBS 0.00352f
C819 VDD.n694 VSUBS 0.0111f
C820 VDD.n695 VSUBS 0.00352f
C821 VDD.n696 VSUBS 0.00352f
C822 VDD.n697 VSUBS 0.0111f
C823 VDD.n698 VSUBS 0.00352f
C824 VDD.n699 VSUBS 0.00352f
C825 VDD.n700 VSUBS 0.0111f
C826 VDD.n701 VSUBS 0.00352f
C827 VDD.n702 VSUBS 0.00352f
C828 VDD.n703 VSUBS 0.0111f
C829 VDD.n704 VSUBS 0.00352f
C830 VDD.n705 VSUBS 0.00352f
C831 VDD.n706 VSUBS 0.0111f
C832 VDD.n707 VSUBS 0.00352f
C833 VDD.n708 VSUBS 0.00352f
C834 VDD.n709 VSUBS 0.0111f
C835 VDD.n710 VSUBS 0.00352f
C836 VDD.n711 VSUBS 0.00352f
C837 VDD.n712 VSUBS 0.0111f
C838 VDD.n713 VSUBS 0.00352f
C839 VDD.n714 VSUBS 0.00352f
C840 VDD.n715 VSUBS 0.0111f
C841 VDD.n716 VSUBS 0.00352f
C842 VDD.n717 VSUBS 0.00352f
C843 VDD.n718 VSUBS 0.0111f
C844 VDD.n719 VSUBS 0.00352f
C845 VDD.n720 VSUBS 0.00352f
C846 VDD.n721 VSUBS 0.0111f
C847 VDD.n722 VSUBS 0.00352f
C848 VDD.n723 VSUBS 0.00352f
C849 VDD.n724 VSUBS 0.0111f
C850 VDD.n725 VSUBS 0.00352f
C851 VDD.n726 VSUBS 0.00352f
C852 VDD.n727 VSUBS 0.0111f
C853 VDD.n728 VSUBS 0.00352f
C854 VDD.n729 VSUBS 0.00352f
C855 VDD.n730 VSUBS 0.0111f
C856 VDD.n731 VSUBS 0.00352f
C857 VDD.n732 VSUBS 0.00352f
C858 VDD.n733 VSUBS 0.0111f
C859 VDD.n734 VSUBS 0.00352f
C860 VDD.n735 VSUBS 0.00352f
C861 VDD.n736 VSUBS 0.0111f
C862 VDD.n737 VSUBS 0.00352f
C863 VDD.n738 VSUBS 0.00352f
C864 VDD.n739 VSUBS 0.0111f
C865 VDD.n740 VSUBS 0.00352f
C866 VDD.n741 VSUBS 0.00352f
C867 VDD.n742 VSUBS 0.0111f
C868 VDD.n743 VSUBS 0.00352f
C869 VDD.n744 VSUBS 0.00352f
C870 VDD.n745 VSUBS 0.0111f
C871 VDD.n746 VSUBS 0.00352f
C872 VDD.n747 VSUBS 0.00352f
C873 VDD.n748 VSUBS 0.0111f
C874 VDD.n749 VSUBS 0.00352f
C875 VDD.n750 VSUBS 0.00352f
C876 VDD.n751 VSUBS 0.0111f
C877 VDD.n752 VSUBS 0.00352f
C878 VDD.n753 VSUBS 0.00352f
C879 VDD.n754 VSUBS 0.0111f
C880 VDD.n755 VSUBS 0.00352f
C881 VDD.n756 VSUBS 0.00352f
C882 VDD.n757 VSUBS 0.0105f
C883 VDD.n758 VSUBS 0.00944f
C884 VDD.n759 VSUBS 0.00352f
C885 VDD.n760 VSUBS 0.00352f
C886 VDD.n761 VSUBS 0.00609f
C887 VDD.n762 VSUBS 0.00352f
C888 VDD.n763 VSUBS 0.00352f
C889 VDD.n764 VSUBS 0.0111f
C890 VDD.n765 VSUBS 0.00352f
C891 VDD.n766 VSUBS 0.00352f
C892 VDD.n767 VSUBS 0.0111f
C893 VDD.n768 VSUBS 0.00352f
C894 VDD.n769 VSUBS 0.00352f
C895 VDD.n770 VSUBS 0.00807f
C896 VDD.n771 VSUBS 0.00373f
C897 VDD.n772 VSUBS 0.00343f
C898 VDD.n773 VSUBS 0.00352f
C899 VDD.n774 VSUBS 0.00352f
C900 VDD.n775 VSUBS 0.00352f
C901 VDD.n776 VSUBS 0.00352f
C902 VDD.n777 VSUBS 0.00243f
C903 VDD.n778 VSUBS 0.0142f
C904 VDD.n779 VSUBS 0.00352f
C905 VDD.n780 VSUBS 0.00286f
C906 VDD.n781 VSUBS 0.00352f
C907 VDD.n782 VSUBS 0.00352f
C908 VDD.n783 VSUBS 0.00352f
C909 VDD.n784 VSUBS 0.00309f
C910 VDD.n785 VSUBS 0.0128f
C911 VDD.n786 VSUBS 0.00352f
C912 VDD.n787 VSUBS 0.00219f
C913 VDD.n788 VSUBS 0.00352f
C914 VDD.n789 VSUBS 0.00352f
C915 VDD.n790 VSUBS 0.00352f
C916 VDD.n791 VSUBS 0.00352f
C917 VDD.n793 VSUBS 0.00352f
C918 VDD.n794 VSUBS 0.002f
C919 VDD.n795 VSUBS 0.0156f
C920 VDD.n796 VSUBS 0.00352f
C921 VDD.n797 VSUBS 0.00329f
C922 VDD.n799 VSUBS 0.00352f
C923 VDD.n800 VSUBS 0.00352f
C924 VDD.n801 VSUBS 0.00352f
C925 VDD.n802 VSUBS 0.00246f
C926 VDD.n803 VSUBS 0.0155f
C927 VDD.n805 VSUBS 0.00352f
C928 VDD.n806 VSUBS 0.00282f
C929 VDD.n807 VSUBS 0.00352f
C930 VDD.n808 VSUBS 0.00352f
C931 VDD.n810 VSUBS 0.00352f
C932 VDD.n811 VSUBS 0.00352f
C933 VDD.n812 VSUBS 0.00352f
C934 VDD.n813 VSUBS 0.00352f
C935 VDD.n815 VSUBS 0.00352f
C936 VDD.n816 VSUBS 0.00352f
C937 VDD.n817 VSUBS 0.00352f
C938 VDD.n818 VSUBS 0.00352f
C939 VDD.n820 VSUBS 0.00352f
C940 VDD.n821 VSUBS 0.00352f
C941 VDD.n823 VSUBS 0.00352f
C942 VDD.n824 VSUBS 0.00352f
C943 VDD.n825 VSUBS 0.00288f
C944 VDD.n826 VSUBS 0.00288f
C945 VDD.n827 VSUBS 0.00424f
C946 VDD.n844 VSUBS 0.304f
C947 VDD.n846 VSUBS 0.00432f
C948 VDD.n847 VSUBS 0.00432f
C949 VDD.n848 VSUBS 0.214f
C950 VDD.n849 VSUBS 0.00352f
C951 VDD.n850 VSUBS 0.00352f
C952 VDD.n851 VSUBS 0.214f
C953 VDD.n852 VSUBS 0.00352f
C954 VDD.n853 VSUBS 0.00352f
C955 VDD.n854 VSUBS 0.214f
C956 VDD.n855 VSUBS 0.00352f
C957 VDD.n856 VSUBS 0.00352f
C958 VDD.t2 VSUBS 0.107f
C959 VDD.n857 VSUBS 0.109f
C960 VDD.n858 VSUBS 0.00352f
C961 VDD.n859 VSUBS 0.00194f
C962 VDD.n860 VSUBS 0.00567f
C963 VDD.n861 VSUBS 0.212f
C964 VDD.n862 VSUBS 0.00352f
C965 VDD.n863 VSUBS 0.00334f
C966 VDD.n864 VSUBS 0.00352f
C967 VDD.n865 VSUBS 0.201f
C968 VDD.n866 VSUBS 0.00352f
C969 VDD.n867 VSUBS 0.00352f
C970 VDD.t26 VSUBS 0.107f
C971 VDD.n868 VSUBS 0.00352f
C972 VDD.n869 VSUBS 0.12f
C973 VDD.n870 VSUBS 0.00352f
C974 VDD.n871 VSUBS 0.00352f
C975 VDD.n872 VSUBS 0.00352f
C976 VDD.n873 VSUBS 0.214f
C977 VDD.n874 VSUBS 0.00352f
C978 VDD.n875 VSUBS 0.00352f
C979 VDD.n876 VSUBS 0.00352f
C980 VDD.n877 VSUBS 0.186f
C981 VDD.n878 VSUBS 0.00352f
C982 VDD.n879 VSUBS 0.00352f
C983 VDD.t20 VSUBS 0.107f
C984 VDD.n880 VSUBS 0.00352f
C985 VDD.n881 VSUBS 0.135f
C986 VDD.n882 VSUBS 0.00352f
C987 VDD.n883 VSUBS 0.00352f
C988 VDD.n884 VSUBS 0.00352f
C989 VDD.n885 VSUBS 0.214f
C990 VDD.n886 VSUBS 0.00352f
C991 VDD.n887 VSUBS 0.00352f
C992 VDD.n888 VSUBS 0.00352f
C993 VDD.n889 VSUBS 0.17f
C994 VDD.n890 VSUBS 0.00352f
C995 VDD.n891 VSUBS 0.00352f
C996 VDD.t25 VSUBS 0.107f
C997 VDD.n892 VSUBS 0.00352f
C998 VDD.n893 VSUBS 0.151f
C999 VDD.n894 VSUBS 0.00352f
C1000 VDD.n895 VSUBS 0.00352f
C1001 VDD.n896 VSUBS 0.00352f
C1002 VDD.n897 VSUBS 0.214f
C1003 VDD.n898 VSUBS 0.00352f
C1004 VDD.n899 VSUBS 0.00352f
C1005 VDD.t33 VSUBS 0.107f
C1006 VDD.n900 VSUBS 0.00352f
C1007 VDD.n901 VSUBS 0.155f
C1008 VDD.n902 VSUBS 0.00352f
C1009 VDD.n903 VSUBS 0.00352f
C1010 VDD.n904 VSUBS 0.00352f
C1011 VDD.n905 VSUBS 0.166f
C1012 VDD.n906 VSUBS 0.00352f
C1013 VDD.n907 VSUBS 0.00352f
C1014 VDD.n908 VSUBS 0.00352f
C1015 VDD.n909 VSUBS 0.214f
C1016 VDD.n910 VSUBS 0.00352f
C1017 VDD.n911 VSUBS 0.00352f
C1018 VDD.t8 VSUBS 0.107f
C1019 VDD.n912 VSUBS 0.00352f
C1020 VDD.n913 VSUBS 0.14f
C1021 VDD.n914 VSUBS 0.00352f
C1022 VDD.n915 VSUBS 0.00352f
C1023 VDD.n916 VSUBS 0.00352f
C1024 VDD.n917 VSUBS 0.181f
C1025 VDD.n918 VSUBS 0.00352f
C1026 VDD.n919 VSUBS 0.00352f
C1027 VDD.n920 VSUBS 0.00352f
C1028 VDD.n921 VSUBS 0.214f
C1029 VDD.n922 VSUBS 0.00352f
C1030 VDD.n923 VSUBS 0.00352f
C1031 VDD.t30 VSUBS 0.107f
C1032 VDD.n924 VSUBS 0.00352f
C1033 VDD.n925 VSUBS 0.124f
C1034 VDD.n926 VSUBS 0.00352f
C1035 VDD.n927 VSUBS 0.00352f
C1036 VDD.n928 VSUBS 0.00352f
C1037 VDD.n929 VSUBS 0.197f
C1038 VDD.n930 VSUBS 0.00352f
C1039 VDD.n931 VSUBS 0.00352f
C1040 VDD.n932 VSUBS 0.00352f
C1041 VDD.n933 VSUBS 0.214f
C1042 VDD.n934 VSUBS 0.00352f
C1043 VDD.n935 VSUBS 0.00352f
C1044 VDD.t19 VSUBS 0.107f
C1045 VDD.n936 VSUBS 0.00352f
C1046 VDD.n937 VSUBS 0.109f
C1047 VDD.n938 VSUBS 0.00352f
C1048 VDD.n939 VSUBS 0.00352f
C1049 VDD.n940 VSUBS 0.00352f
C1050 VDD.n941 VSUBS 0.212f
C1051 VDD.n942 VSUBS 0.00352f
C1052 VDD.n943 VSUBS 0.00352f
C1053 VDD.n944 VSUBS 0.00352f
C1054 VDD.n945 VSUBS 0.201f
C1055 VDD.n946 VSUBS 0.00352f
C1056 VDD.n947 VSUBS 0.00352f
C1057 VDD.t41 VSUBS 0.107f
C1058 VDD.n948 VSUBS 0.00352f
C1059 VDD.n949 VSUBS 0.00352f
C1060 VDD.n950 VSUBS 0.00352f
C1061 VDD.n951 VSUBS 0.12f
C1062 VDD.n952 VSUBS 0.00352f
C1063 VDD.n953 VSUBS 0.00352f
C1064 VDD.n954 VSUBS 0.00352f
C1065 VDD.n955 VSUBS 0.00352f
C1066 VDD.n956 VSUBS 0.00352f
C1067 VDD.n957 VSUBS 0.214f
C1068 VDD.n958 VSUBS 0.00352f
C1069 VDD.n959 VSUBS 0.00352f
C1070 VDD.n960 VSUBS 0.00352f
C1071 VDD.n961 VSUBS 0.00352f
C1072 VDD.n962 VSUBS 0.00352f
C1073 VDD.n963 VSUBS 0.186f
C1074 VDD.n964 VSUBS 0.00352f
C1075 VDD.n965 VSUBS 0.00352f
C1076 VDD.t42 VSUBS 0.107f
C1077 VDD.n966 VSUBS 0.00352f
C1078 VDD.n967 VSUBS 0.00352f
C1079 VDD.n968 VSUBS 0.00352f
C1080 VDD.n969 VSUBS 0.135f
C1081 VDD.n970 VSUBS 0.00352f
C1082 VDD.n971 VSUBS 0.00352f
C1083 VDD.n972 VSUBS 0.00352f
C1084 VDD.n973 VSUBS 0.00352f
C1085 VDD.n974 VSUBS 0.00352f
C1086 VDD.n975 VSUBS 0.214f
C1087 VDD.n976 VSUBS 0.00352f
C1088 VDD.n977 VSUBS 0.00352f
C1089 VDD.n978 VSUBS 0.00352f
C1090 VDD.n979 VSUBS 0.00352f
C1091 VDD.n980 VSUBS 0.00352f
C1092 VDD.n981 VSUBS 0.17f
C1093 VDD.n982 VSUBS 0.00352f
C1094 VDD.n983 VSUBS 0.00352f
C1095 VDD.t27 VSUBS 0.107f
C1096 VDD.n984 VSUBS 0.00352f
C1097 VDD.n985 VSUBS 0.00352f
C1098 VDD.n986 VSUBS 0.00352f
C1099 VDD.n987 VSUBS 0.151f
C1100 VDD.n988 VSUBS 0.00352f
C1101 VDD.n989 VSUBS 0.00352f
C1102 VDD.n990 VSUBS 0.00352f
C1103 VDD.n991 VSUBS 0.00352f
C1104 VDD.n992 VSUBS 0.00352f
C1105 VDD.n993 VSUBS 0.214f
C1106 VDD.n994 VSUBS 0.00352f
C1107 VDD.n995 VSUBS 0.00352f
C1108 VDD.t1 VSUBS 0.107f
C1109 VDD.n996 VSUBS 0.00352f
C1110 VDD.n997 VSUBS 0.00352f
C1111 VDD.n998 VSUBS 0.00352f
C1112 VDD.n999 VSUBS 0.155f
C1113 VDD.n1000 VSUBS 0.00352f
C1114 VDD.n1001 VSUBS 0.00352f
C1115 VDD.n1002 VSUBS 0.00352f
C1116 VDD.n1003 VSUBS 0.00352f
C1117 VDD.n1004 VSUBS 0.00352f
C1118 VDD.n1005 VSUBS 0.00352f
C1119 VDD.n1006 VSUBS 0.00352f
C1120 VDD.n1007 VSUBS 0.166f
C1121 VDD.n1008 VSUBS 0.00352f
C1122 VDD.n1009 VSUBS 0.00352f
C1123 VDD.n1010 VSUBS 0.00352f
C1124 VDD.n1011 VSUBS 0.00352f
C1125 VDD.n1012 VSUBS 0.00352f
C1126 VDD.n1013 VSUBS 0.00352f
C1127 VDD.n1014 VSUBS 0.214f
C1128 VDD.n1015 VSUBS 0.00352f
C1129 VDD.n1016 VSUBS 0.00352f
C1130 VDD.t34 VSUBS 0.107f
C1131 VDD.n1017 VSUBS 0.00352f
C1132 VDD.n1018 VSUBS 0.00352f
C1133 VDD.n1019 VSUBS 0.00352f
C1134 VDD.n1020 VSUBS 0.00352f
C1135 VDD.n1021 VSUBS 0.14f
C1136 VDD.n1022 VSUBS 0.00352f
C1137 VDD.n1023 VSUBS 0.00352f
C1138 VDD.n1024 VSUBS 0.00352f
C1139 VDD.n1025 VSUBS 0.00352f
C1140 VDD.n1026 VSUBS 0.00352f
C1141 VDD.n1027 VSUBS 0.181f
C1142 VDD.n1028 VSUBS 0.00352f
C1143 VDD.n1029 VSUBS 0.00352f
C1144 VDD.n1030 VSUBS 0.00352f
C1145 VDD.n1031 VSUBS 0.00352f
C1146 VDD.n1032 VSUBS 0.00352f
C1147 VDD.n1033 VSUBS 0.00352f
C1148 VDD.n1034 VSUBS 0.00352f
C1149 VDD.n1035 VSUBS 0.214f
C1150 VDD.n1036 VSUBS 0.00352f
C1151 VDD.n1037 VSUBS 0.00352f
C1152 VDD.t29 VSUBS 0.107f
C1153 VDD.n1038 VSUBS 0.00352f
C1154 VDD.n1039 VSUBS 0.00352f
C1155 VDD.n1040 VSUBS 0.00352f
C1156 VDD.n1041 VSUBS 0.00352f
C1157 VDD.n1042 VSUBS 0.124f
C1158 VDD.n1043 VSUBS 0.00352f
C1159 VDD.n1044 VSUBS 0.00352f
C1160 VDD.n1045 VSUBS 0.00352f
C1161 VDD.n1046 VSUBS 0.00352f
C1162 VDD.n1047 VSUBS 0.00352f
C1163 VDD.n1048 VSUBS 0.00352f
C1164 VDD.n1049 VSUBS 0.197f
C1165 VDD.n1050 VSUBS 0.00352f
C1166 VDD.n1051 VSUBS 0.00352f
C1167 VDD.n1052 VSUBS 0.00352f
C1168 VDD.n1053 VSUBS 0.00352f
C1169 VDD.n1054 VSUBS 0.00352f
C1170 VDD.n1055 VSUBS 0.214f
C1171 VDD.n1056 VSUBS 0.00352f
C1172 VDD.n1057 VSUBS 0.00352f
C1173 VDD.t6 VSUBS 0.107f
C1174 VDD.n1058 VSUBS 0.00352f
C1175 VDD.n1059 VSUBS 0.00352f
C1176 VDD.n1060 VSUBS 0.00352f
C1177 VDD.n1061 VSUBS 0.00352f
C1178 VDD.n1062 VSUBS 0.00352f
C1179 VDD.n1063 VSUBS 0.109f
C1180 VDD.n1064 VSUBS 0.00352f
C1181 VDD.n1065 VSUBS 0.00352f
C1182 VDD.n1066 VSUBS 0.00352f
C1183 VDD.n1067 VSUBS 0.00352f
C1184 VDD.n1068 VSUBS 0.00352f
C1185 VDD.n1069 VSUBS 0.00352f
C1186 VDD.n1070 VSUBS 0.212f
C1187 VDD.n1071 VSUBS 0.00352f
C1188 VDD.n1072 VSUBS 0.00352f
C1189 VDD.n1073 VSUBS 0.00352f
C1190 VDD.n1074 VSUBS 0.00352f
C1191 VDD.n1075 VSUBS 0.00352f
C1192 VDD.n1076 VSUBS 0.00352f
C1193 VDD.n1077 VSUBS 0.201f
C1194 VDD.n1078 VSUBS 0.00352f
C1195 VDD.n1079 VSUBS 0.00352f
C1196 VDD.t7 VSUBS 0.107f
C1197 VDD.n1080 VSUBS 0.00352f
C1198 VDD.n1081 VSUBS 0.00352f
C1199 VDD.n1082 VSUBS 0.00352f
C1200 VDD.n1083 VSUBS 0.00352f
C1201 VDD.n1084 VSUBS 0.12f
C1202 VDD.n1085 VSUBS 0.00352f
C1203 VDD.n1086 VSUBS 0.00263f
.ends

