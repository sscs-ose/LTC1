magic
tech gf180mcuC
magscale 1 10
timestamp 1694074718
<< pwell >>
rect -860 -1104 860 1104
<< nmos >>
rect -748 436 -692 1036
rect -588 436 -532 1036
rect -428 436 -372 1036
rect -268 436 -212 1036
rect -108 436 -52 1036
rect 52 436 108 1036
rect 212 436 268 1036
rect 372 436 428 1036
rect 532 436 588 1036
rect 692 436 748 1036
rect -748 -300 -692 300
rect -588 -300 -532 300
rect -428 -300 -372 300
rect -268 -300 -212 300
rect -108 -300 -52 300
rect 52 -300 108 300
rect 212 -300 268 300
rect 372 -300 428 300
rect 532 -300 588 300
rect 692 -300 748 300
rect -748 -1036 -692 -436
rect -588 -1036 -532 -436
rect -428 -1036 -372 -436
rect -268 -1036 -212 -436
rect -108 -1036 -52 -436
rect 52 -1036 108 -436
rect 212 -1036 268 -436
rect 372 -1036 428 -436
rect 532 -1036 588 -436
rect 692 -1036 748 -436
<< ndiff >>
rect -836 1023 -748 1036
rect -836 449 -823 1023
rect -777 449 -748 1023
rect -836 436 -748 449
rect -692 1023 -588 1036
rect -692 449 -663 1023
rect -617 449 -588 1023
rect -692 436 -588 449
rect -532 1023 -428 1036
rect -532 449 -503 1023
rect -457 449 -428 1023
rect -532 436 -428 449
rect -372 1023 -268 1036
rect -372 449 -343 1023
rect -297 449 -268 1023
rect -372 436 -268 449
rect -212 1023 -108 1036
rect -212 449 -183 1023
rect -137 449 -108 1023
rect -212 436 -108 449
rect -52 1023 52 1036
rect -52 449 -23 1023
rect 23 449 52 1023
rect -52 436 52 449
rect 108 1023 212 1036
rect 108 449 137 1023
rect 183 449 212 1023
rect 108 436 212 449
rect 268 1023 372 1036
rect 268 449 297 1023
rect 343 449 372 1023
rect 268 436 372 449
rect 428 1023 532 1036
rect 428 449 457 1023
rect 503 449 532 1023
rect 428 436 532 449
rect 588 1023 692 1036
rect 588 449 617 1023
rect 663 449 692 1023
rect 588 436 692 449
rect 748 1023 836 1036
rect 748 449 777 1023
rect 823 449 836 1023
rect 748 436 836 449
rect -836 287 -748 300
rect -836 -287 -823 287
rect -777 -287 -748 287
rect -836 -300 -748 -287
rect -692 287 -588 300
rect -692 -287 -663 287
rect -617 -287 -588 287
rect -692 -300 -588 -287
rect -532 287 -428 300
rect -532 -287 -503 287
rect -457 -287 -428 287
rect -532 -300 -428 -287
rect -372 287 -268 300
rect -372 -287 -343 287
rect -297 -287 -268 287
rect -372 -300 -268 -287
rect -212 287 -108 300
rect -212 -287 -183 287
rect -137 -287 -108 287
rect -212 -300 -108 -287
rect -52 287 52 300
rect -52 -287 -23 287
rect 23 -287 52 287
rect -52 -300 52 -287
rect 108 287 212 300
rect 108 -287 137 287
rect 183 -287 212 287
rect 108 -300 212 -287
rect 268 287 372 300
rect 268 -287 297 287
rect 343 -287 372 287
rect 268 -300 372 -287
rect 428 287 532 300
rect 428 -287 457 287
rect 503 -287 532 287
rect 428 -300 532 -287
rect 588 287 692 300
rect 588 -287 617 287
rect 663 -287 692 287
rect 588 -300 692 -287
rect 748 287 836 300
rect 748 -287 777 287
rect 823 -287 836 287
rect 748 -300 836 -287
rect -836 -449 -748 -436
rect -836 -1023 -823 -449
rect -777 -1023 -748 -449
rect -836 -1036 -748 -1023
rect -692 -449 -588 -436
rect -692 -1023 -663 -449
rect -617 -1023 -588 -449
rect -692 -1036 -588 -1023
rect -532 -449 -428 -436
rect -532 -1023 -503 -449
rect -457 -1023 -428 -449
rect -532 -1036 -428 -1023
rect -372 -449 -268 -436
rect -372 -1023 -343 -449
rect -297 -1023 -268 -449
rect -372 -1036 -268 -1023
rect -212 -449 -108 -436
rect -212 -1023 -183 -449
rect -137 -1023 -108 -449
rect -212 -1036 -108 -1023
rect -52 -449 52 -436
rect -52 -1023 -23 -449
rect 23 -1023 52 -449
rect -52 -1036 52 -1023
rect 108 -449 212 -436
rect 108 -1023 137 -449
rect 183 -1023 212 -449
rect 108 -1036 212 -1023
rect 268 -449 372 -436
rect 268 -1023 297 -449
rect 343 -1023 372 -449
rect 268 -1036 372 -1023
rect 428 -449 532 -436
rect 428 -1023 457 -449
rect 503 -1023 532 -449
rect 428 -1036 532 -1023
rect 588 -449 692 -436
rect 588 -1023 617 -449
rect 663 -1023 692 -449
rect 588 -1036 692 -1023
rect 748 -449 836 -436
rect 748 -1023 777 -449
rect 823 -1023 836 -449
rect 748 -1036 836 -1023
<< ndiffc >>
rect -823 449 -777 1023
rect -663 449 -617 1023
rect -503 449 -457 1023
rect -343 449 -297 1023
rect -183 449 -137 1023
rect -23 449 23 1023
rect 137 449 183 1023
rect 297 449 343 1023
rect 457 449 503 1023
rect 617 449 663 1023
rect 777 449 823 1023
rect -823 -287 -777 287
rect -663 -287 -617 287
rect -503 -287 -457 287
rect -343 -287 -297 287
rect -183 -287 -137 287
rect -23 -287 23 287
rect 137 -287 183 287
rect 297 -287 343 287
rect 457 -287 503 287
rect 617 -287 663 287
rect 777 -287 823 287
rect -823 -1023 -777 -449
rect -663 -1023 -617 -449
rect -503 -1023 -457 -449
rect -343 -1023 -297 -449
rect -183 -1023 -137 -449
rect -23 -1023 23 -449
rect 137 -1023 183 -449
rect 297 -1023 343 -449
rect 457 -1023 503 -449
rect 617 -1023 663 -449
rect 777 -1023 823 -449
<< polysilicon >>
rect -748 1036 -692 1080
rect -588 1036 -532 1080
rect -428 1036 -372 1080
rect -268 1036 -212 1080
rect -108 1036 -52 1080
rect 52 1036 108 1080
rect 212 1036 268 1080
rect 372 1036 428 1080
rect 532 1036 588 1080
rect 692 1036 748 1080
rect -748 392 -692 436
rect -588 392 -532 436
rect -428 392 -372 436
rect -268 392 -212 436
rect -108 392 -52 436
rect 52 392 108 436
rect 212 392 268 436
rect 372 392 428 436
rect 532 392 588 436
rect 692 392 748 436
rect -748 300 -692 344
rect -588 300 -532 344
rect -428 300 -372 344
rect -268 300 -212 344
rect -108 300 -52 344
rect 52 300 108 344
rect 212 300 268 344
rect 372 300 428 344
rect 532 300 588 344
rect 692 300 748 344
rect -748 -344 -692 -300
rect -588 -344 -532 -300
rect -428 -344 -372 -300
rect -268 -344 -212 -300
rect -108 -344 -52 -300
rect 52 -344 108 -300
rect 212 -344 268 -300
rect 372 -344 428 -300
rect 532 -344 588 -300
rect 692 -344 748 -300
rect -748 -436 -692 -392
rect -588 -436 -532 -392
rect -428 -436 -372 -392
rect -268 -436 -212 -392
rect -108 -436 -52 -392
rect 52 -436 108 -392
rect 212 -436 268 -392
rect 372 -436 428 -392
rect 532 -436 588 -392
rect 692 -436 748 -392
rect -748 -1080 -692 -1036
rect -588 -1080 -532 -1036
rect -428 -1080 -372 -1036
rect -268 -1080 -212 -1036
rect -108 -1080 -52 -1036
rect 52 -1080 108 -1036
rect 212 -1080 268 -1036
rect 372 -1080 428 -1036
rect 532 -1080 588 -1036
rect 692 -1080 748 -1036
<< metal1 >>
rect -823 1023 -777 1034
rect -823 438 -777 449
rect -663 1023 -617 1034
rect -663 438 -617 449
rect -503 1023 -457 1034
rect -503 438 -457 449
rect -343 1023 -297 1034
rect -343 438 -297 449
rect -183 1023 -137 1034
rect -183 438 -137 449
rect -23 1023 23 1034
rect -23 438 23 449
rect 137 1023 183 1034
rect 137 438 183 449
rect 297 1023 343 1034
rect 297 438 343 449
rect 457 1023 503 1034
rect 457 438 503 449
rect 617 1023 663 1034
rect 617 438 663 449
rect 777 1023 823 1034
rect 777 438 823 449
rect -823 287 -777 298
rect -823 -298 -777 -287
rect -663 287 -617 298
rect -663 -298 -617 -287
rect -503 287 -457 298
rect -503 -298 -457 -287
rect -343 287 -297 298
rect -343 -298 -297 -287
rect -183 287 -137 298
rect -183 -298 -137 -287
rect -23 287 23 298
rect -23 -298 23 -287
rect 137 287 183 298
rect 137 -298 183 -287
rect 297 287 343 298
rect 297 -298 343 -287
rect 457 287 503 298
rect 457 -298 503 -287
rect 617 287 663 298
rect 617 -298 663 -287
rect 777 287 823 298
rect 777 -298 823 -287
rect -823 -449 -777 -438
rect -823 -1034 -777 -1023
rect -663 -449 -617 -438
rect -663 -1034 -617 -1023
rect -503 -449 -457 -438
rect -503 -1034 -457 -1023
rect -343 -449 -297 -438
rect -343 -1034 -297 -1023
rect -183 -449 -137 -438
rect -183 -1034 -137 -1023
rect -23 -449 23 -438
rect -23 -1034 23 -1023
rect 137 -449 183 -438
rect 137 -1034 183 -1023
rect 297 -449 343 -438
rect 297 -1034 343 -1023
rect 457 -449 503 -438
rect 457 -1034 503 -1023
rect 617 -449 663 -438
rect 617 -1034 663 -1023
rect 777 -449 823 -438
rect 777 -1034 823 -1023
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 3 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
