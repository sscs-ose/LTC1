* NGSPICE file created from ppolyf_u_WRMTN3_flat.ext - technology: gf180mcuC

.subckt ppolyf_u_WRMTN3_flat VDD VSS VINP VINN OUT VC VD VX VA VB VBS2 VBS3 VBIASN
+ IBIAS2 VBIASN2 IBIAS3 IBIAS OUTo VP c_mid
X0 VDD IBIAS3.t78 OUTo.t78 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1 VSS.t128 VSS.t127 VSS.t128 VSS.t90 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X2 VDD.t419 VDD.t418 VDD.t419 VDD.t353 pfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X3 OUTo IBIAS3.t79 VDD.t262 VDD.t29 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X4 VDD IBIAS3.t34 IBIAS3.t35 VDD.t12 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X5 VSS OUT.t30 OUTo.t154 VSS.t49 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X6 VDD IBIAS.t6 VBS3.t7 VDD.t311 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X7 VA VBS2.t4 VX.t17 VDD.t436 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X8 VSS VX.t20 VC.t15 VSS.t52 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X9 VSS VX.t21 VC.t14 VSS.t57 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X10 VDD IBIAS3.t80 OUTo.t77 VDD.t18 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X11 OUTo IBIAS3.t81 VDD.t257 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X12 VD VBS3.t8 OUT.t20 VSS.t153 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X13 VDD.t417 VDD.t416 VDD.t417 VDD.t333 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X14 VC VX.t22 VSS.t161 VSS.t55 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X15 OUTo IBIAS3.t82 VDD.t256 VDD.t82 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X16 VX.t7 VX.t6 VX.t7 VSS.t39 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X17 VSS.t126 VSS.t125 VSS.t126 VSS.t84 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X18 VP VINP.t0 VD.t0 VDD.t7 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X19 IBIAS3 VBIASN2.t20 VSS.t208 VSS.t174 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X20 VX VBS3.t9 VC.t23 VSS.t12 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X21 VSS OUT.t31 OUTo.t155 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X22 VD.t64 VD.t63 VD.t64 VSS.t3 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X23 OUTo OUT.t32 VSS.t241 VSS.t26 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X24 OUTo IBIAS3.t83 VDD.t255 VDD.t34 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X25 VSS VD.t47 VD.t48 VSS.t0 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X26 OUTo IBIAS3.t84 VDD.t254 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X27 VDD IBIAS3.t85 OUTo.t76 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X28 VDD IBIAS3.t86 OUTo.t75 VDD.t147 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X29 VDD.t415 VDD.t414 VDD.t415 VDD.t339 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X30 VSS VX.t23 VD.t16 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X31 VC VINN.t0 VP.t51 VDD.t434 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X32 c_mid.t4 OUT.t0 cap_mim_2f0_m4m5_noshield c_width=24u c_length=15.5u
X33 OUTo OUT.t33 VSS.t242 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X34 OUT.t18 OUT.t17 OUT.t18 VSS.t39 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X35 OUTo IBIAS3.t87 VDD.t249 VDD.t76 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X36 VDD IBIAS3.t88 OUTo.t74 VDD.t65 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X37 VD VD.t45 VSS.t20 VSS.t19 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X38 VP IBIAS.t7 VDD.t315 VDD.t314 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X39 VBS2 VBIASN.t4 VSS.t269 VSS.t268 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.56u
X40 VC.t39 VC.t38 VC.t39 VDD.t301 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X41 VC.t37 VC.t36 VC.t37 VDD.t301 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X42 VDD.t413 VDD.t412 VDD.t413 VDD.t366 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X43 VDD IBIAS3.t32 IBIAS3.t33 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X44 VSS VX.t24 VC.t12 VSS.t57 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X45 VD VINP.t1 VP.t30 VDD.t437 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X46 VDD IBIAS3.t89 OUTo.t73 VDD.t108 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X47 OUTo OUT.t34 VSS.t230 VSS.t31 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X48 VDD IBIAS3.t90 OUTo.t72 VDD.t147 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X49 VSS OUT.t35 OUTo.t150 VSS.t35 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X50 VB.t15 VB.t14 VB.t15 VDD.t282 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X51 VDD VBS2.t1 VBS2.t2 VDD.t308 pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.56u
X52 VDD IBIAS3.t91 OUTo.t71 VDD.t65 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X53 OUTo IBIAS3.t92 VDD.t239 VDD.t82 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X54 OUTo OUT.t36 VSS.t233 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X55 VSS VBIASN2.t21 IBIAS3.t74 VSS.t176 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X56 VSS.t124 VSS.t122 VSS.t124 VSS.t123 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=0.56u
X57 IBIAS3 VBIASN2.t22 VSS.t203 VSS.t174 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X58 VDD IBIAS3.t30 IBIAS3.t31 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X59 VDD IBIAS3.t93 OUTo.t70 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X60 IBIAS IBIAS.t4 VDD.t302 VDD.t286 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X61 VP VINP.t2 VD.t31 VDD.t438 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X62 IBIAS3 IBIAS3.t36 VDD.t234 VDD.t89 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X63 VDD IBIAS3.t95 OUTo.t69 VDD.t108 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X64 VDD.t411 VDD.t410 VDD.t411 VDD.t366 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X65 VBIASN VBIASN.t2 VSS.t267 VSS.t266 nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.56u
X66 VSS OUT.t37 OUTo.t152 VSS.t41 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X67 VDD.t409 VDD.t408 VDD.t409 VDD.t363 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X68 VA VBS2.t5 VX.t16 VDD.t436 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X69 OUTo IBIAS3.t96 VDD.t230 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X70 OUTo OUT.t38 VSS.t236 VSS.t26 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X71 VX VBS3.t10 VC.t22 VSS.t11 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X72 OUTo IBIAS3.t97 VDD.t229 VDD.t34 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X73 VDD.t407 VDD.t406 VDD.t407 VDD.t350 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X74 VDD.t405 VDD.t404 VDD.t405 VDD.t339 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X75 VSS OUT.t39 OUTo.t158 VSS.t44 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X76 VBIASN2 IBIAS2.t5 VDD.t285 VDD.t284 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X77 VDD.t403 VDD.t402 VDD.t403 VDD.t333 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X78 VSS VBIASN2.t23 IBIAS3.t76 VSS.t192 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X79 VDD IBIAS3.t98 OUTo.t68 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X80 VDD IBIAS.t9 VP.t14 VDD.t290 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X81 VP VINN.t1 VC.t56 VDD.t428 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X82 c_mid.t1 OUTo.t141 VDD.t307 ppolyf_u r_width=0.8u r_length=6.46u
X83 VP IBIAS.t10 VDD.t455 VDD.t314 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X84 VBS3 IBIAS.t11 VDD.t457 VDD.t456 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X85 VDD IBIAS3.t99 OUTo.t67 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X86 VSS VX.t25 VC.t11 VSS.t6 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X87 VA.t15 VA.t14 VA.t15 VDD.t282 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X88 VSS VBIASN2.t24 IBIAS3.t71 VSS.t176 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X89 VP IBIAS.t12 VDD.t458 VDD.t326 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X90 VDD IBIAS3.t100 OUTo.t66 VDD.t50 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X91 OUTo OUT.t40 VSS.t245 VSS.t47 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X92 OUTo IBIAS3.t101 VDD.t222 VDD.t34 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X93 VDD.t401 VDD.t400 VDD.t401 VDD.t363 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X94 VDD.t399 VDD.t398 VDD.t399 VDD.t358 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X95 VDD IBIAS3.t102 OUTo.t65 VDD.t55 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X96 VSS.t121 VSS.t120 VSS.t121 VSS.t84 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X97 VSS OUT.t41 OUTo.t160 VSS.t49 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X98 VC VX.t26 VSS.t139 VSS.t4 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X99 VP IBIAS.t13 VDD.t462 VDD.t326 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X100 IBIAS3 VBIASN2.t25 VSS.t198 VSS.t190 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X101 VDD.t460 VDD.t461 VDD.t459 ppolyf_u r_width=0.8u r_length=6.46u
X102 OUTo OUT.t42 VSS.t248 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X103 VDD IBIAS3.t103 OUTo.t64 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X104 VSS.t119 VSS.t118 VSS.t119 VSS.t106 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X105 VD VX.t27 VSS.t166 VSS.t9 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X106 VSS VC.t50 VC.t51 VSS.t156 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X107 OUT.t16 OUT.t15 OUT.t16 VSS.t39 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X108 VC VX.t28 VSS.t167 VSS.t142 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X109 VDD IBIAS3.t104 OUTo.t63 VDD.t55 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X110 IBIAS2 IBIAS2.t3 VDD.t9 VDD.t8 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X111 VSS OUT.t43 OUTo.t162 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X112 VDD IBIAS3.t28 IBIAS3.t29 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X113 VC VINN.t2 VP.t48 VDD.t429 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X114 OUTo IBIAS3.t105 VDD.t213 VDD.t45 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X115 VC VINN.t3 VP.t49 VDD.t429 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X116 OUTo OUT.t44 VSS.t221 VSS.t31 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X117 VDD IBIAS3.t106 OUTo.t62 VDD.t15 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X118 VSS OUT.t45 OUTo.t145 VSS.t41 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X119 VDD.t397 VDD.t396 VDD.t397 VDD.t363 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X120 VC VBS3.t11 VX.t11 VSS.t165 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X121 VDD.t395 VDD.t394 VDD.t395 VDD.t358 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X122 VDD IBIAS.t14 VA.t7 VDD.t293 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X123 IBIAS3 IBIAS3.t42 VDD.t210 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X124 VDD IBIAS.t15 VP.t10 VDD.t272 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X125 VP.t47 VP.t46 VP.t47 VDD.t435 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X126 VB VBS2.t6 OUT.t28 VDD.t439 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X127 c_mid.t2 OUTo.t142 VDD.t321 ppolyf_u r_width=0.8u r_length=6.46u
X128 OUTo IBIAS3.t108 VDD.t209 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X129 VBIASN2 VBIASN2.t17 VSS.t207 VSS.t172 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X130 VDD.t393 VDD.t391 VDD.t393 VDD.t392 pfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=0.56u
X131 VBIASN2 IBIAS2.t7 VDD.t276 VDD.t275 pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X132 OUTo IBIAS3.t109 VDD.t208 VDD.t29 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X133 VDD IBIAS.t16 VP.t9 VDD.t272 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X134 OUTo IBIAS3.t110 VDD.t207 VDD.t68 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X135 VC VX.t29 VSS.t168 VSS.t4 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X136 VDD IBIAS3.t111 OUTo.t61 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X137 VDD.t390 VDD.t389 VDD.t390 VDD.t333 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X138 VD VX.t30 VSS.t143 VSS.t142 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X139 VDD.t388 VDD.t387 VDD.t388 VDD.t333 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X140 OUTo IBIAS3.t112 VDD.t204 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X141 VSS OUT.t46 OUTo.t146 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X142 VSS.t117 VSS.t116 VSS.t117 VSS.t90 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X143 VDD.t386 VDD.t385 VDD.t386 VDD.t363 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X144 VC VBS3.t12 VX.t10 VSS.t153 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X145 VDD.t384 VDD.t383 VDD.t384 VDD.t358 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X146 VSS VD.t43 VD.t44 VSS.t16 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X147 VC VC.t48 VSS.t152 VSS.t151 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X148 IBIAS3 IBIAS3.t38 VDD.t203 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X149 VP.t45 VP.t44 VP.t45 VDD.t435 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X150 VDD.t382 VDD.t381 VDD.t382 VDD.t339 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X151 VD VBS3.t13 OUT.t21 VSS.t165 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X152 VSS VBIASN2.t27 IBIAS3.t73 VSS.t192 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X153 VD.t62 VD.t61 VD.t62 VSS.t164 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X154 VD.t60 VD.t59 VD.t60 VDD.t301 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X155 VP VINP.t3 VD.t34 VDD.t7 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X156 VDD.t380 VDD.t379 VDD.t380 VDD.t366 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X157 VSS VBS3.t2 VBS3.t3 VSS.t213 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X158 VSS OUT.t47 OUTo.t147 VSS.t49 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X159 VP.t43 VP.t42 VP.t43 VDD.t435 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X160 VDD IBIAS3.t114 OUTo.t60 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X161 VSS.t115 VSS.t114 VSS.t115 VSS.t84 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X162 OUTo IBIAS3.t115 VDD.t200 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X163 VC VX.t31 VSS.t144 VSS.t142 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X164 VDD.t378 VDD.t377 VDD.t378 VDD.t350 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X165 OUTo IBIAS3.t116 VDD.t199 VDD.t76 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X166 VDD.t376 VDD.t375 VDD.t376 VDD.t336 pfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=1u
X167 VDD IBIAS3.t117 OUTo.t59 VDD.t18 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X168 c_mid.t0 OUTo.t120 VDD.t265 ppolyf_u r_width=0.8u r_length=6.46u
X169 VDD IBIAS3.t118 OUTo.t58 VDD.t15 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X170 VC VINN.t4 VP.t50 VDD.t434 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X171 IBIAS3 VBIASN2.t28 VSS.t191 VSS.t190 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X172 VA.t13 VA.t12 VA.t13 VDD.t282 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X173 VSS OUT.t48 OUTo.t148 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X174 VDD IBIAS3.t119 OUTo.t57 VDD.t65 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X175 OUTo OUT.t49 VSS.t281 VSS.t31 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X176 VSS.t113 VSS.t112 VSS.t113 VSS.t106 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X177 OUTo OUT.t50 VSS.t282 VSS.t26 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X178 VDD IBIAS3.t120 OUTo.t56 VDD.t10 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X179 VDD IBIAS3.t121 OUTo.t55 VDD.t147 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X180 VD VINP.t4 VP.t27 VDD.t298 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X181 c_mid.t3 OUTo.t163 VDD.t447 ppolyf_u r_width=0.8u r_length=6.46u
X182 VDD.t374 VDD.t373 VDD.t374 VDD.t350 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X183 OUT VBS2.t7 VB.t18 VDD.t420 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X184 IBIAS3 IBIAS3.t52 VDD.t188 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X185 VD VINP.t5 VP.t26 VDD.t298 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X186 OUTo IBIAS3.t123 VDD.t187 VDD.t87 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X187 OUTo IBIAS3.t124 VDD.t186 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X188 VD VD.t41 VSS.t63 VSS.t62 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X189 OUTo OUT.t51 VSS.t283 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X190 OUTo IBIAS3.t125 VDD.t185 VDD.t87 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X191 VDD IBIAS3.t126 OUTo.t54 VDD.t18 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X192 VX.t5 VX.t4 VX.t5 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X193 VDD.t372 VDD.t370 VDD.t372 VDD.t371 pfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=0.56u
X194 VSS VBIASN2.t29 IBIAS3.t69 VSS.t192 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X195 VDD IBIAS.t17 VB.t7 VDD.t293 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X196 OUTo IBIAS3.t127 VDD.t182 VDD.t39 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X197 VBIASN2 VBIASN2.t15 VSS.t206 VSS.t172 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X198 VSS.t111 VSS.t110 VSS.t111 VSS.t90 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X199 VP IBIAS.t18 VDD.t454 VDD.t326 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X200 VSS.t109 VSS.t108 VSS.t109 VSS.t90 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X201 VDD.t369 VDD.t368 VDD.t369 VDD.t366 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X202 VP VINP.t6 VD.t35 VDD.t442 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X203 VDD IBIAS.t19 VP.t7 VDD.t272 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X204 VP VINP.t7 VD.t36 VDD.t442 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X205 c_mid.t5 OUT.t29 cap_mim_2f0_m4m5_noshield c_width=24u c_length=15.5u
X206 VD.t58 VD.t57 VD.t58 VSS.t164 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X207 VB VBS2.t8 OUT.t24 VDD.t439 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X208 VDD IBIAS3.t128 OUTo.t53 VDD.t147 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X209 VSS OUT.t52 OUTo.t182 VSS.t35 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X210 VDD IBIAS3.t129 OUTo.t52 VDD.t59 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X211 IBIAS3 IBIAS3.t48 VDD.t176 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X212 VDD IBIAS3.t131 OUTo.t51 VDD.t108 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X213 VDD.t445 VDD.t446 VDD.t444 ppolyf_u r_width=0.8u r_length=6.46u
X214 VB IBIAS.t20 VDD.t330 VDD.t1 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X215 IBIAS3 VBIASN2.t31 VSS.t195 VSS.t190 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X216 VDD.t367 VDD.t365 VDD.t367 VDD.t366 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X217 OUT VBS3.t14 VD.t22 VSS.t12 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X218 OUT.t14 OUT.t13 OUT.t14 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X219 VSS.t107 VSS.t105 VSS.t107 VSS.t106 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X220 VSS VX.t32 VD.t13 VSS.t52 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X221 VDD IBIAS2.t8 VBIASN2.t4 VDD.t318 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X222 VC.t35 VC.t34 VC.t35 VDD.t300 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X223 VDD IBIAS3.t132 OUTo.t50 VDD.t50 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X224 VSS OUT.t53 OUTo.t183 VSS.t44 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X225 VC.t33 VC.t32 VC.t33 VDD.t300 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X226 IBIAS3 VBIASN2.t32 VSS.t186 VSS.t182 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X227 VD VINP.t8 VP.t23 VDD.t429 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X228 VDD IBIAS3.t133 OUTo.t49 VDD.t108 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X229 VSS VX.t33 VD.t12 VSS.t52 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X230 OUTo OUT.t54 VSS.t76 VSS.t26 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X231 OUTo IBIAS3.t134 VDD.t170 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X232 VDD IBIAS3.t135 OUTo.t48 VDD.t10 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X233 VA IBIAS.t21 VDD.t331 VDD.t322 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X234 VC.t31 VC.t30 VC.t31 VSS.t3 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X235 OUTo OUT.t55 VSS.t77 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X236 VD VX.t34 VSS.t56 VSS.t55 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X237 VBIASN2 VBIASN2.t13 VSS.t173 VSS.t172 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X238 VB.t13 VB.t12 VB.t13 VDD.t282 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X239 VA IBIAS.t22 VDD.t2 VDD.t1 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X240 OUTo IBIAS3.t136 VDD.t167 VDD.t29 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X241 VC VC.t46 VSS.t150 VSS.t149 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X242 VBS3 IBIAS.t23 VDD.t4 VDD.t3 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X243 VDD IBIAS3.t137 OUTo.t47 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X244 OUTo OUT.t56 VSS.t78 VSS.t47 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X245 IBIAS3 IBIAS3.t50 VDD.t161 VDD.t89 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X246 VD VBS3.t15 OUT.t23 VSS.t153 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X247 OUTo IBIAS3.t139 VDD.t164 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X248 VSS VBIASN2.t34 IBIAS3.t66 VSS.t179 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X249 VC VBS3.t16 VX.t9 VSS.t165 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X250 VDD IBIAS3.t140 OUTo.t46 VDD.t50 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X251 OUTo IBIAS3.t141 VDD.t160 VDD.t87 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X252 VSS VX.t35 VD.t10 VSS.t57 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X253 VD VD.t39 VSS.t61 VSS.t60 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X254 VDD IBIAS3.t142 OUTo.t45 VDD.t10 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X255 VSS.t104 VSS.t103 VSS.t104 VSS.t87 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X256 VBIASN IBIAS.t24 VDD.t6 VDD.t5 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.56u
X257 VDD.t364 VDD.t362 VDD.t364 VDD.t363 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X258 IBIAS2 VBIASN.t6 VSS.t22 VSS.t21 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.56u
X259 OUT VBS2.t9 VB.t16 VDD.t420 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X260 VDD.t361 VDD.t360 VDD.t361 VDD.t358 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X261 VSS.t102 VSS.t101 VSS.t102 VSS.t84 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X262 IBIAS3 IBIAS3.t44 VDD.t157 VDD.t89 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X263 OUTo OUT.t57 VSS.t80 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X264 VDD.t359 VDD.t357 VDD.t359 VDD.t358 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X265 IBIAS3 IBIAS3.t46 VDD.t152 VDD.t89 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X266 VDD IBIAS3.t145 OUTo.t44 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X267 VSS VX.t36 VD.t9 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X268 VC.t29 VC.t28 VC.t29 VSS.t3 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X269 VB IBIAS.t25 VDD.t323 VDD.t322 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X270 VSS VD.t37 VD.t38 VSS.t13 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X271 VDD IBIAS3.t146 OUTo.t43 VDD.t15 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X272 OUTo IBIAS3.t147 VDD.t151 VDD.t87 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X273 VSS OUT.t58 OUTo.t140 VSS.t35 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X274 VBIASN2 IBIAS2.t9 VDD.t467 VDD.t284 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X275 VDD IBIAS.t26 VB.t4 VDD.t266 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X276 OUTo IBIAS3.t148 VDD.t150 VDD.t68 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X277 OUTo OUT.t59 VSS.t40 VSS.t31 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X278 VSS VX.t37 VC.t6 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X279 VDD IBIAS2.t10 VBIASN2.t1 VDD.t277 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X280 VDD IBIAS3.t149 OUTo.t42 VDD.t147 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X281 VSS OUT.t60 OUTo.t127 VSS.t41 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X282 IBIAS3 IBIAS3.t4 VDD.t135 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X283 VSS OUT.t61 OUTo.t128 VSS.t44 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X284 VD VX.t38 VSS.t134 VSS.t55 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X285 VDD IBIAS3.t151 OUTo.t41 VDD.t59 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X286 VDD IBIAS3.t152 OUTo.t40 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X287 VP IBIAS.t27 VDD.t327 VDD.t326 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X288 VP IBIAS.t28 VDD.t468 VDD.t314 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X289 VDD IBIAS3.t153 OUTo.t39 VDD.t55 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X290 VX VBS3.t17 VC.t18 VSS.t11 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X291 VD.t56 VD.t55 VD.t56 VDD.t301 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X292 IBIAS3 VBIASN2.t35 VSS.t189 VSS.t182 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X293 VC VINN.t5 VP.t53 VDD.t298 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X294 OUTo IBIAS3.t154 VDD.t140 VDD.t68 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X295 OUTo IBIAS3.t155 VDD.t139 VDD.t68 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X296 OUTo OUT.t62 VSS.t48 VSS.t47 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X297 OUTo IBIAS3.t156 VDD.t138 VDD.t45 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X298 VP IBIAS.t29 VDD.t469 VDD.t314 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X299 VSS.t100 VSS.t99 VSS.t100 VSS.t90 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X300 VSS VX.t39 VD.t7 VSS.t57 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X301 VSS OUT.t63 OUTo.t130 VSS.t49 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X302 VB IBIAS.t30 VDD.t470 VDD.t1 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X303 VDD IBIAS3.t157 OUTo.t38 VDD.t59 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X304 VX.t3 VX.t2 VX.t3 VSS.t39 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X305 VC VINN.t6 VP.t54 VDD.t437 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X306 OUTo IBIAS3.t158 VDD.t134 VDD.t45 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X307 VC VINN.t7 VP.t55 VDD.t437 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X308 VP VINN.t8 VC.t65 VDD.t442 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X309 VSS VBIASN2.t36 IBIAS3.t62 VSS.t179 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X310 VDD IBIAS3.t159 OUTo.t37 VDD.t55 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X311 OUTo IBIAS3.t160 VDD.t131 VDD.t39 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X312 VSS.t98 VSS.t97 VSS.t98 VSS.t84 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X313 VDD.t356 VDD.t355 VDD.t356 VDD.t350 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X314 VDD.t354 VDD.t352 VDD.t354 VDD.t353 pfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X315 VBIASN2 IBIAS2.t11 VDD.t449 VDD.t275 pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X316 VDD IBIAS3.t161 OUTo.t36 VDD.t18 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X317 VSS.t96 VSS.t95 VSS.t96 VSS.t87 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X318 VP VINN.t9 VC.t66 VDD.t438 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X319 VP VINN.t10 VC.t67 VDD.t438 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X320 OUTo OUT.t64 VSS.t27 VSS.t26 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X321 VSS VX.t40 VC.t5 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X322 OUT VBS3.t18 VD.t20 VSS.t11 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X323 IBIAS3 IBIAS3.t40 VDD.t128 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X324 VSS OUT.t65 OUTo.t122 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X325 OUTo IBIAS3.t163 VDD.t127 VDD.t45 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X326 OUTo OUT.t66 VSS.t32 VSS.t31 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X327 VC VC.t44 VSS.t148 VSS.t147 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X328 VDD IBIAS.t2 IBIAS.t3 VDD.t5 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X329 OUTo IBIAS3.t164 VDD.t126 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X330 OUTo OUT.t67 VSS.t34 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X331 IBIAS3 VBIASN2.t37 VSS.t183 VSS.t182 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X332 VA IBIAS.t31 VDD.t421 VDD.t322 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X333 VSS.t94 VSS.t92 VSS.t94 VSS.t93 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=0.56u
X334 OUTo IBIAS3.t165 VDD.t125 VDD.t39 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X335 VD.t54 VD.t53 VD.t54 VDD.t300 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X336 VDD IBIAS3.t26 IBIAS3.t27 VDD.t12 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X337 VP.t41 VP.t40 VP.t41 VDD.t435 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.56u
X338 OUT.t12 OUT.t11 OUT.t12 VDD.t299 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X339 IBIAS3 IBIAS3.t58 VDD.t122 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X340 OUTo IBIAS3.t167 VDD.t121 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X341 VSS VX.t41 VD.t6 VSS.t6 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X342 VSS VBIASN2.t11 VBIASN2.t12 VSS.t169 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X343 VBIASN IBIAS.t32 VDD.t423 VDD.t422 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.56u
X344 VDD IBIAS3.t24 IBIAS3.t25 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X345 VP VINP.t9 VD.t67 VDD.t428 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X346 VP VINP.t10 VD.t27 VDD.t428 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X347 VSS OUT.t68 OUTo.t125 VSS.t35 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X348 VDD IBIAS.t33 VB.t2 VDD.t266 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X349 VSS VBIASN2.t38 IBIAS3.t64 VSS.t179 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X350 OUTo IBIAS3.t168 VDD.t118 VDD.t76 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X351 OUTo IBIAS3.t169 VDD.t117 VDD.t29 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X352 VSS.t91 VSS.t89 VSS.t91 VSS.t90 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X353 OUTo IBIAS3.t170 VDD.t116 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X354 IBIAS3 IBIAS3.t0 VDD.t115 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X355 VDD IBIAS3.t22 IBIAS3.t23 VDD.t12 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X356 VSS OUT.t69 OUTo.t169 VSS.t49 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X357 VP.t39 VP.t38 VP.t39 VDD.t0 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.56u
X358 VC VX.t42 VSS.t294 VSS.t9 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X359 VSS VX.t43 VC.t3 VSS.t6 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X360 OUTo IBIAS3.t172 VDD.t112 VDD.t39 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X361 OUTo IBIAS3.t173 VDD.t111 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X362 VDD IBIAS3.t174 OUTo.t35 VDD.t108 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X363 VSS.t88 VSS.t86 VSS.t88 VSS.t87 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X364 OUTo IBIAS3.t175 VDD.t107 VDD.t82 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X365 VB IBIAS.t34 VDD.t430 VDD.t322 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X366 VSS VC.t42 VC.t43 VSS.t216 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X367 VD VINP.t11 VP.t20 VDD.t429 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X368 VSS VBIASN.t7 VBS2.t0 VSS.t23 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.56u
X369 VDD.t351 VDD.t349 VDD.t351 VDD.t350 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X370 VDD IBIAS.t35 VA.t3 VDD.t266 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X371 VD VX.t44 VSS.t297 VSS.t142 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X372 VB.t11 VB.t10 VB.t11 VDD.t283 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.56u
X373 VDD IBIAS3.t20 IBIAS3.t21 VDD.t12 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X374 VDD IBIAS3.t176 OUTo.t34 VDD.t59 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X375 VDD IBIAS3.t177 OUTo.t33 VDD.t50 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X376 VSS OUT.t70 OUTo.t170 VSS.t44 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X377 VDD IBIAS3.t178 OUTo.t32 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X378 VA IBIAS.t36 VDD.t433 VDD.t1 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X379 VD VX.t45 VSS.t5 VSS.t4 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X380 OUTo OUT.t71 VSS.t262 VSS.t26 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X381 VDD IBIAS3.t179 OUTo.t31 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X382 VDD IBIAS3.t180 OUTo.t30 VDD.t10 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X383 OUTo IBIAS3.t181 VDD.t94 VDD.t82 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X384 OUTo OUT.t72 VSS.t263 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X385 OUT VBS3.t19 VD.t19 VSS.t11 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X386 VSS VX.t46 VD.t3 VSS.t6 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X387 OUTo IBIAS3.t182 VDD.t93 VDD.t76 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X388 VD VX.t47 VSS.t10 VSS.t9 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X389 IBIAS3 IBIAS3.t54 VDD.t92 VDD.t91 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X390 VC.t27 VC.t26 VC.t27 VSS.t164 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X391 VA.t11 VA.t10 VA.t11 VDD.t283 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.56u
X392 VBS3 VBS3.t0 VSS.t155 VSS.t154 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X393 VSS OUT.t73 OUTo.t173 VSS.t44 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X394 OUTo OUT.t74 VSS.t251 VSS.t47 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X395 IBIAS3 IBIAS3.t2 VDD.t90 VDD.t89 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X396 VDD IBIAS.t37 VP.t3 VDD.t290 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X397 OUTo IBIAS3.t185 VDD.t88 VDD.t87 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X398 VX VBS2.t10 VA.t17 VDD.t443 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X399 VDD IBIAS3.t186 OUTo.t29 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X400 VX.t1 VX.t0 VX.t1 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X401 VSS OUT.t75 OUTo.t165 VSS.t35 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X402 VC VX.t48 VSS.t64 VSS.t9 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X403 OUTo IBIAS3.t187 VDD.t83 VDD.t82 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X404 OUTo OUT.t76 VSS.t254 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X405 VDD IBIAS3.t188 OUTo.t28 VDD.t65 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X406 VDD IBIAS.t38 VB.t0 VDD.t293 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X407 VSS VBIASN2.t9 VBIASN2.t10 VSS.t169 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X408 VDD.t348 VDD.t346 VDD.t348 VDD.t347 pfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=0.56u
X409 VDD IBIAS3.t18 IBIAS3.t19 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X410 VP.t37 VP.t36 VP.t37 VDD.t0 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.56u
X411 VDD IBIAS2.t12 VBIASN2.t5 VDD.t318 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X412 OUT.t10 OUT.t9 OUT.t10 VDD.t299 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X413 VX VBS3.t21 VC.t17 VSS.t12 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X414 OUT.t8 OUT.t7 OUT.t8 VDD.t289 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X415 VP VINN.t11 VC.t62 VDD.t7 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X416 OUTo IBIAS3.t189 VDD.t77 VDD.t76 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X417 VDD IBIAS3.t16 IBIAS3.t17 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X418 VDD IBIAS.t39 VA.t1 VDD.t293 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X419 VP VINN.t12 VC.t63 VDD.t7 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X420 VC.t25 VC.t24 VC.t25 VSS.t164 nfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X421 VD VINP.t12 VP.t19 VDD.t437 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X422 VDD IBIAS.t40 VA.t0 VDD.t266 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X423 VP.t35 VP.t34 VP.t35 VDD.t0 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.56u
X424 OUTo IBIAS3.t190 VDD.t73 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X425 VDD IBIAS3.t191 OUTo.t27 VDD.t70 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X426 VSS OUT.t77 OUTo.t167 VSS.t41 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X427 OUTo IBIAS3.t192 VDD.t69 VDD.t68 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X428 OUT VBS3.t22 VD.t18 VSS.t12 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X429 VD VINP.t13 VP.t18 VDD.t434 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X430 VDD IBIAS3.t193 OUTo.t26 VDD.t65 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X431 OUTo IBIAS3.t194 VDD.t64 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X432 VD VINP.t14 VP.t17 VDD.t434 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X433 VDD IBIAS.t41 VBS3.t4 VDD.t269 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.56u
X434 OUTo OUT.t78 VSS.t257 VSS.t47 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X435 VD VX.t49 VSS.t65 VSS.t4 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X436 VP VINP.t15 VD.t33 VDD.t438 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X437 VC VINN.t13 VP.t60 VDD.t298 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X438 VDD.t345 VDD.t344 VDD.t345 VDD.t339 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X439 VSS OUT.t79 OUTo.t174 VSS.t44 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X440 VDD IBIAS3.t14 IBIAS3.t15 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X441 IBIAS2 IBIAS2.t1 VDD.t448 VDD.t8 pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X442 VDD IBIAS.t42 VP.t2 VDD.t272 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X443 VDD IBIAS3.t195 OUTo.t25 VDD.t59 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X444 VC VBS3.t23 VX.t8 VSS.t153 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X445 VDD IBIAS.t43 VP.t1 VDD.t290 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X446 VD VBS3.t24 OUT.t26 VSS.t165 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X447 VDD IBIAS3.t12 IBIAS3.t13 VDD.t52 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X448 VDD IBIAS3.t196 OUTo.t24 VDD.t55 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X449 VDD IBIAS3.t197 OUTo.t23 VDD.t50 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X450 VDD.t343 VDD.t341 VDD.t343 VDD.t342 pfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=0.56u
X451 VSS VBIASN2.t7 VBIASN2.t8 VSS.t169 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X452 VP VINN.t14 VC.t60 VDD.t442 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X453 VDD IBIAS.t44 VP.t0 VDD.t290 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X454 OUTo OUT.t80 VSS.t272 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X455 OUTo OUT.t81 VSS.t273 VSS.t47 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X456 OUTo IBIAS3.t198 VDD.t49 VDD.t48 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X457 OUTo IBIAS3.t199 VDD.t47 VDD.t34 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X458 VSS OUT.t82 OUTo.t177 VSS.t49 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X459 VP VINN.t15 VC.t61 VDD.t428 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X460 VDD.t340 VDD.t338 VDD.t340 VDD.t339 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X461 IBIAS3 VBIASN2.t39 VSS.t175 VSS.t174 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X462 VB.t9 VB.t8 VB.t9 VDD.t283 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.56u
X463 OUTo OUT.t83 VSS.t276 VSS.t79 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X464 OUTo IBIAS3.t200 VDD.t46 VDD.t45 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X465 VSS VX.t50 VC.t1 VSS.t52 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X466 VDD IBIAS2.t14 VBIASN2.t2 VDD.t277 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X467 OUTo IBIAS3.t201 VDD.t44 VDD.t43 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X468 IBIAS3 IBIAS3.t56 VDD.t42 VDD.t41 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X469 OUTo IBIAS3.t203 VDD.t40 VDD.t39 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X470 VSS.t85 VSS.t83 VSS.t85 VSS.t84 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X471 OUTo IBIAS3.t204 VDD.t38 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X472 VSS OUT.t84 OUTo.t131 VSS.t28 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X473 VDD IBIAS3.t10 IBIAS3.t11 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X474 VD.t52 VD.t51 VD.t52 VDD.t300 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X475 OUTo IBIAS3.t205 VDD.t35 VDD.t34 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X476 VDD IBIAS3.t8 IBIAS3.t9 VDD.t12 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X477 VDD IBIAS3.t206 OUTo.t22 VDD.t15 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X478 VSS OUT.t85 OUTo.t132 VSS.t41 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X479 VX VBS2.t11 VA.t16 VDD.t443 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X480 VD.t50 VD.t49 VD.t50 VSS.t3 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X481 OUTo OUT.t86 VSS.t72 VSS.t31 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X482 VSS OUT.t87 OUTo.t134 VSS.t41 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X483 OUT.t6 OUT.t5 OUT.t6 VDD.t289 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X484 OUTo IBIAS3.t207 VDD.t30 VDD.t29 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X485 OUTo IBIAS3.t208 VDD.t27 VDD.t26 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X486 OUTo OUT.t88 VSS.t75 VSS.t33 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X487 VDD.t337 VDD.t335 VDD.t337 VDD.t336 pfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=1u
X488 VP.t33 VP.t32 VP.t33 VDD.t0 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.56u
X489 VSS VC.t40 VC.t41 VSS.t278 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X490 VDD IBIAS3.t6 IBIAS3.t7 VDD.t23 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X491 OUTo IBIAS3.t209 VDD.t22 VDD.t21 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X492 VDD.t334 VDD.t332 VDD.t334 VDD.t333 pfet_03v3 ad=0.78p pd=3.52u as=0 ps=0 w=3u l=0.28u
X493 VC VX.t51 VSS.t277 VSS.t55 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X494 VDD IBIAS.t0 IBIAS.t1 VDD.t286 pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.56u
X495 VDD IBIAS3.t210 OUTo.t21 VDD.t18 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X496 VSS VBIASN2.t40 IBIAS3.t61 VSS.t176 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X497 VDD IBIAS3.t211 OUTo.t20 VDD.t15 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X498 OUT.t4 OUT.t3 OUT.t4 VSS.t38 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X499 VDD IBIAS3.t212 OUTo.t19 VDD.t10 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X500 VA.t9 VA.t8 VA.t9 VDD.t283 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.56u
X501 VSS OUT.t89 OUTo.t143 VSS.t35 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
R0 IBIAS3.n119 IBIAS3.t191 57.4713
R1 IBIAS3.n123 IBIAS3.t208 57.4713
R2 IBIAS3.n341 IBIAS3.t85 57.4713
R3 IBIAS3.n345 IBIAS3.t87 57.4713
R4 IBIAS3.n229 IBIAS3.t174 57.4713
R5 IBIAS3.n233 IBIAS3.t192 57.4713
R6 IBIAS3.n80 IBIAS3.t152 42.888
R7 IBIAS3.n81 IBIAS3.t198 42.888
R8 IBIAS3.n82 IBIAS3.t90 42.888
R9 IBIAS3.n83 IBIAS3.t163 42.888
R10 IBIAS3.n84 IBIAS3.t14 42.888
R11 IBIAS3.n89 IBIAS3.t48 42.888
R12 IBIAS3.n88 IBIAS3.t159 42.888
R13 IBIAS3.n87 IBIAS3.t205 42.888
R14 IBIAS3.n86 IBIAS3.t140 42.888
R15 IBIAS3.n59 IBIAS3.t114 42.888
R16 IBIAS3.n60 IBIAS3.t108 42.888
R17 IBIAS3.n61 IBIAS3.t149 42.888
R18 IBIAS3.n62 IBIAS3.t156 42.888
R19 IBIAS3.n63 IBIAS3.t12 42.888
R20 IBIAS3.n68 IBIAS3.t56 42.888
R21 IBIAS3.n67 IBIAS3.t102 42.888
R22 IBIAS3.n66 IBIAS3.t97 42.888
R23 IBIAS3.n64 IBIAS3.t139 42.888
R24 IBIAS3.n44 IBIAS3.t197 42.888
R25 IBIAS3.n45 IBIAS3.t83 42.888
R26 IBIAS3.n46 IBIAS3.t104 42.888
R27 IBIAS3.n47 IBIAS3.t40 42.888
R28 IBIAS3.n42 IBIAS3.t18 42.888
R29 IBIAS3.n41 IBIAS3.t105 42.888
R30 IBIAS3.n40 IBIAS3.t128 42.888
R31 IBIAS3.n39 IBIAS3.t190 42.888
R32 IBIAS3.n38 IBIAS3.t78 42.888
R33 IBIAS3.n43 IBIAS3.t134 42.888
R34 IBIAS3.n65 IBIAS3.t100 42.888
R35 IBIAS3.n85 IBIAS3.t170 42.888
R36 IBIAS3.n302 IBIAS3.t186 42.888
R37 IBIAS3.n303 IBIAS3.t79 42.888
R38 IBIAS3.n304 IBIAS3.t103 42.888
R39 IBIAS3.n305 IBIAS3.t181 42.888
R40 IBIAS3.n306 IBIAS3.t6 42.888
R41 IBIAS3.n311 IBIAS3.t46 42.888
R42 IBIAS3.n310 IBIAS3.t193 42.888
R43 IBIAS3.n309 IBIAS3.t84 42.888
R44 IBIAS3.n308 IBIAS3.t157 42.888
R45 IBIAS3.n281 IBIAS3.t99 42.888
R46 IBIAS3.n282 IBIAS3.t136 42.888
R47 IBIAS3.n283 IBIAS3.t179 42.888
R48 IBIAS3.n284 IBIAS3.t187 42.888
R49 IBIAS3.n285 IBIAS3.t32 42.888
R50 IBIAS3.n290 IBIAS3.t36 42.888
R51 IBIAS3.n289 IBIAS3.t88 42.888
R52 IBIAS3.n288 IBIAS3.t124 42.888
R53 IBIAS3.n286 IBIAS3.t168 42.888
R54 IBIAS3.n266 IBIAS3.t176 42.888
R55 IBIAS3.n267 IBIAS3.t201 42.888
R56 IBIAS3.n268 IBIAS3.t119 42.888
R57 IBIAS3.n269 IBIAS3.t44 42.888
R58 IBIAS3.n264 IBIAS3.t24 42.888
R59 IBIAS3.n263 IBIAS3.t92 42.888
R60 IBIAS3.n262 IBIAS3.t111 42.888
R61 IBIAS3.n261 IBIAS3.t169 42.888
R62 IBIAS3.n260 IBIAS3.t93 42.888
R63 IBIAS3.n265 IBIAS3.t116 42.888
R64 IBIAS3.n287 IBIAS3.t129 42.888
R65 IBIAS3.n307 IBIAS3.t189 42.888
R66 IBIAS3.n190 IBIAS3.t133 42.888
R67 IBIAS3.n191 IBIAS3.t165 42.888
R68 IBIAS3.n192 IBIAS3.t211 42.888
R69 IBIAS3.n193 IBIAS3.t147 42.888
R70 IBIAS3.n194 IBIAS3.t20 42.888
R71 IBIAS3.n199 IBIAS3.t38 42.888
R72 IBIAS3.n198 IBIAS3.t142 42.888
R73 IBIAS3.n197 IBIAS3.t173 42.888
R74 IBIAS3.n196 IBIAS3.t126 42.888
R75 IBIAS3.n169 IBIAS3.t89 42.888
R76 IBIAS3.n170 IBIAS3.t127 42.888
R77 IBIAS3.n171 IBIAS3.t118 42.888
R78 IBIAS3.n172 IBIAS3.t125 42.888
R79 IBIAS3.n173 IBIAS3.t26 42.888
R80 IBIAS3.n178 IBIAS3.t0 42.888
R81 IBIAS3.n177 IBIAS3.t212 42.888
R82 IBIAS3.n176 IBIAS3.t112 42.888
R83 IBIAS3.n174 IBIAS3.t110 42.888
R84 IBIAS3.n154 IBIAS3.t80 42.888
R85 IBIAS3.n155 IBIAS3.t204 42.888
R86 IBIAS3.n156 IBIAS3.t120 42.888
R87 IBIAS3.n157 IBIAS3.t54 42.888
R88 IBIAS3.n152 IBIAS3.t8 42.888
R89 IBIAS3.n151 IBIAS3.t123 42.888
R90 IBIAS3.n150 IBIAS3.t146 42.888
R91 IBIAS3.n149 IBIAS3.t172 42.888
R92 IBIAS3.n148 IBIAS3.t95 42.888
R93 IBIAS3.n153 IBIAS3.t155 42.888
R94 IBIAS3.n175 IBIAS3.t210 42.888
R95 IBIAS3.n195 IBIAS3.t154 42.888
R96 IBIAS3.n101 IBIAS3.t145 42.6273
R97 IBIAS3.n102 IBIAS3.t194 42.6273
R98 IBIAS3.n103 IBIAS3.t86 42.6273
R99 IBIAS3.n104 IBIAS3.t158 42.6273
R100 IBIAS3.n105 IBIAS3.t16 42.6273
R101 IBIAS3.n110 IBIAS3.t52 42.6273
R102 IBIAS3.n109 IBIAS3.t153 42.6273
R103 IBIAS3.n108 IBIAS3.t199 42.6273
R104 IBIAS3.n106 IBIAS3.t164 42.6273
R105 IBIAS3.n107 IBIAS3.t132 42.6273
R106 IBIAS3.n323 IBIAS3.t178 42.6273
R107 IBIAS3.n324 IBIAS3.t207 42.6273
R108 IBIAS3.n325 IBIAS3.t98 42.6273
R109 IBIAS3.n326 IBIAS3.t175 42.6273
R110 IBIAS3.n327 IBIAS3.t10 42.6273
R111 IBIAS3.n332 IBIAS3.t50 42.6273
R112 IBIAS3.n331 IBIAS3.t188 42.6273
R113 IBIAS3.n330 IBIAS3.t81 42.6273
R114 IBIAS3.n328 IBIAS3.t182 42.6273
R115 IBIAS3.n329 IBIAS3.t151 42.6273
R116 IBIAS3.n211 IBIAS3.t131 42.6273
R117 IBIAS3.n212 IBIAS3.t160 42.6273
R118 IBIAS3.n213 IBIAS3.t206 42.6273
R119 IBIAS3.n214 IBIAS3.t141 42.6273
R120 IBIAS3.n215 IBIAS3.t22 42.6273
R121 IBIAS3.n220 IBIAS3.t42 42.6273
R122 IBIAS3.n219 IBIAS3.t135 42.6273
R123 IBIAS3.n218 IBIAS3.t167 42.6273
R124 IBIAS3.n216 IBIAS3.t148 42.6273
R125 IBIAS3.n217 IBIAS3.t117 42.6273
R126 IBIAS3.n119 IBIAS3.t96 42.4969
R127 IBIAS3.n120 IBIAS3.t121 42.4969
R128 IBIAS3.n121 IBIAS3.t200 42.4969
R129 IBIAS3.n122 IBIAS3.t30 42.4969
R130 IBIAS3.n126 IBIAS3.t58 42.4969
R131 IBIAS3.n125 IBIAS3.t196 42.4969
R132 IBIAS3.n124 IBIAS3.t101 42.4969
R133 IBIAS3.n123 IBIAS3.t177 42.4969
R134 IBIAS3.n341 IBIAS3.t109 42.4969
R135 IBIAS3.n342 IBIAS3.t137 42.4969
R136 IBIAS3.n343 IBIAS3.t82 42.4969
R137 IBIAS3.n344 IBIAS3.t28 42.4969
R138 IBIAS3.n348 IBIAS3.t2 42.4969
R139 IBIAS3.n347 IBIAS3.t91 42.4969
R140 IBIAS3.n346 IBIAS3.t115 42.4969
R141 IBIAS3.n345 IBIAS3.t195 42.4969
R142 IBIAS3.n229 IBIAS3.t203 42.4969
R143 IBIAS3.n230 IBIAS3.t106 42.4969
R144 IBIAS3.n231 IBIAS3.t185 42.4969
R145 IBIAS3.n232 IBIAS3.t34 42.4969
R146 IBIAS3.n236 IBIAS3.t4 42.4969
R147 IBIAS3.n235 IBIAS3.t180 42.4969
R148 IBIAS3.n234 IBIAS3.t209 42.4969
R149 IBIAS3.n233 IBIAS3.t161 42.4969
R150 IBIAS3.n22 IBIAS3.n21 14.9749
R151 IBIAS3.n23 IBIAS3.n22 14.9749
R152 IBIAS3.n24 IBIAS3.n23 14.9749
R153 IBIAS3.n28 IBIAS3.n27 14.9749
R154 IBIAS3.n27 IBIAS3.n26 14.9749
R155 IBIAS3.n26 IBIAS3.n25 14.9749
R156 IBIAS3.n39 IBIAS3.n38 14.9749
R157 IBIAS3.n40 IBIAS3.n39 14.9749
R158 IBIAS3.n41 IBIAS3.n40 14.9749
R159 IBIAS3.n42 IBIAS3.n41 14.9749
R160 IBIAS3.n47 IBIAS3.n46 14.9749
R161 IBIAS3.n46 IBIAS3.n45 14.9749
R162 IBIAS3.n45 IBIAS3.n44 14.9749
R163 IBIAS3.n44 IBIAS3.n43 14.9749
R164 IBIAS3.n60 IBIAS3.n59 14.9749
R165 IBIAS3.n61 IBIAS3.n60 14.9749
R166 IBIAS3.n62 IBIAS3.n61 14.9749
R167 IBIAS3.n63 IBIAS3.n62 14.9749
R168 IBIAS3.n68 IBIAS3.n67 14.9749
R169 IBIAS3.n67 IBIAS3.n66 14.9749
R170 IBIAS3.n66 IBIAS3.n65 14.9749
R171 IBIAS3.n65 IBIAS3.n64 14.9749
R172 IBIAS3.n81 IBIAS3.n80 14.9749
R173 IBIAS3.n82 IBIAS3.n81 14.9749
R174 IBIAS3.n83 IBIAS3.n82 14.9749
R175 IBIAS3.n84 IBIAS3.n83 14.9749
R176 IBIAS3.n89 IBIAS3.n88 14.9749
R177 IBIAS3.n88 IBIAS3.n87 14.9749
R178 IBIAS3.n87 IBIAS3.n86 14.9749
R179 IBIAS3.n86 IBIAS3.n85 14.9749
R180 IBIAS3.n102 IBIAS3.n101 14.9749
R181 IBIAS3.n103 IBIAS3.n102 14.9749
R182 IBIAS3.n104 IBIAS3.n103 14.9749
R183 IBIAS3.n105 IBIAS3.n104 14.9749
R184 IBIAS3.n110 IBIAS3.n109 14.9749
R185 IBIAS3.n109 IBIAS3.n108 14.9749
R186 IBIAS3.n108 IBIAS3.n107 14.9749
R187 IBIAS3.n107 IBIAS3.n106 14.9749
R188 IBIAS3.n120 IBIAS3.n119 14.9749
R189 IBIAS3.n121 IBIAS3.n120 14.9749
R190 IBIAS3.n122 IBIAS3.n121 14.9749
R191 IBIAS3.n126 IBIAS3.n125 14.9749
R192 IBIAS3.n125 IBIAS3.n124 14.9749
R193 IBIAS3.n124 IBIAS3.n123 14.9749
R194 IBIAS3.n244 IBIAS3.n243 14.9749
R195 IBIAS3.n245 IBIAS3.n244 14.9749
R196 IBIAS3.n246 IBIAS3.n245 14.9749
R197 IBIAS3.n250 IBIAS3.n249 14.9749
R198 IBIAS3.n249 IBIAS3.n248 14.9749
R199 IBIAS3.n248 IBIAS3.n247 14.9749
R200 IBIAS3.n261 IBIAS3.n260 14.9749
R201 IBIAS3.n262 IBIAS3.n261 14.9749
R202 IBIAS3.n263 IBIAS3.n262 14.9749
R203 IBIAS3.n264 IBIAS3.n263 14.9749
R204 IBIAS3.n269 IBIAS3.n268 14.9749
R205 IBIAS3.n268 IBIAS3.n267 14.9749
R206 IBIAS3.n267 IBIAS3.n266 14.9749
R207 IBIAS3.n266 IBIAS3.n265 14.9749
R208 IBIAS3.n282 IBIAS3.n281 14.9749
R209 IBIAS3.n283 IBIAS3.n282 14.9749
R210 IBIAS3.n284 IBIAS3.n283 14.9749
R211 IBIAS3.n285 IBIAS3.n284 14.9749
R212 IBIAS3.n290 IBIAS3.n289 14.9749
R213 IBIAS3.n289 IBIAS3.n288 14.9749
R214 IBIAS3.n288 IBIAS3.n287 14.9749
R215 IBIAS3.n287 IBIAS3.n286 14.9749
R216 IBIAS3.n303 IBIAS3.n302 14.9749
R217 IBIAS3.n304 IBIAS3.n303 14.9749
R218 IBIAS3.n305 IBIAS3.n304 14.9749
R219 IBIAS3.n306 IBIAS3.n305 14.9749
R220 IBIAS3.n311 IBIAS3.n310 14.9749
R221 IBIAS3.n310 IBIAS3.n309 14.9749
R222 IBIAS3.n309 IBIAS3.n308 14.9749
R223 IBIAS3.n308 IBIAS3.n307 14.9749
R224 IBIAS3.n324 IBIAS3.n323 14.9749
R225 IBIAS3.n325 IBIAS3.n324 14.9749
R226 IBIAS3.n326 IBIAS3.n325 14.9749
R227 IBIAS3.n327 IBIAS3.n326 14.9749
R228 IBIAS3.n332 IBIAS3.n331 14.9749
R229 IBIAS3.n331 IBIAS3.n330 14.9749
R230 IBIAS3.n330 IBIAS3.n329 14.9749
R231 IBIAS3.n329 IBIAS3.n328 14.9749
R232 IBIAS3.n342 IBIAS3.n341 14.9749
R233 IBIAS3.n343 IBIAS3.n342 14.9749
R234 IBIAS3.n344 IBIAS3.n343 14.9749
R235 IBIAS3.n348 IBIAS3.n347 14.9749
R236 IBIAS3.n347 IBIAS3.n346 14.9749
R237 IBIAS3.n346 IBIAS3.n345 14.9749
R238 IBIAS3.n132 IBIAS3.n131 14.9749
R239 IBIAS3.n133 IBIAS3.n132 14.9749
R240 IBIAS3.n134 IBIAS3.n133 14.9749
R241 IBIAS3.n138 IBIAS3.n137 14.9749
R242 IBIAS3.n137 IBIAS3.n136 14.9749
R243 IBIAS3.n136 IBIAS3.n135 14.9749
R244 IBIAS3.n149 IBIAS3.n148 14.9749
R245 IBIAS3.n150 IBIAS3.n149 14.9749
R246 IBIAS3.n151 IBIAS3.n150 14.9749
R247 IBIAS3.n152 IBIAS3.n151 14.9749
R248 IBIAS3.n157 IBIAS3.n156 14.9749
R249 IBIAS3.n156 IBIAS3.n155 14.9749
R250 IBIAS3.n155 IBIAS3.n154 14.9749
R251 IBIAS3.n154 IBIAS3.n153 14.9749
R252 IBIAS3.n170 IBIAS3.n169 14.9749
R253 IBIAS3.n171 IBIAS3.n170 14.9749
R254 IBIAS3.n172 IBIAS3.n171 14.9749
R255 IBIAS3.n173 IBIAS3.n172 14.9749
R256 IBIAS3.n178 IBIAS3.n177 14.9749
R257 IBIAS3.n177 IBIAS3.n176 14.9749
R258 IBIAS3.n176 IBIAS3.n175 14.9749
R259 IBIAS3.n175 IBIAS3.n174 14.9749
R260 IBIAS3.n191 IBIAS3.n190 14.9749
R261 IBIAS3.n192 IBIAS3.n191 14.9749
R262 IBIAS3.n193 IBIAS3.n192 14.9749
R263 IBIAS3.n194 IBIAS3.n193 14.9749
R264 IBIAS3.n199 IBIAS3.n198 14.9749
R265 IBIAS3.n198 IBIAS3.n197 14.9749
R266 IBIAS3.n197 IBIAS3.n196 14.9749
R267 IBIAS3.n196 IBIAS3.n195 14.9749
R268 IBIAS3.n212 IBIAS3.n211 14.9749
R269 IBIAS3.n213 IBIAS3.n212 14.9749
R270 IBIAS3.n214 IBIAS3.n213 14.9749
R271 IBIAS3.n215 IBIAS3.n214 14.9749
R272 IBIAS3.n220 IBIAS3.n219 14.9749
R273 IBIAS3.n219 IBIAS3.n218 14.9749
R274 IBIAS3.n218 IBIAS3.n217 14.9749
R275 IBIAS3.n217 IBIAS3.n216 14.9749
R276 IBIAS3.n230 IBIAS3.n229 14.9749
R277 IBIAS3.n231 IBIAS3.n230 14.9749
R278 IBIAS3.n232 IBIAS3.n231 14.9749
R279 IBIAS3.n236 IBIAS3.n235 14.9749
R280 IBIAS3.n235 IBIAS3.n234 14.9749
R281 IBIAS3.n234 IBIAS3.n233 14.9749
R282 IBIAS3.n127 IBIAS3.n122 7.86204
R283 IBIAS3.n349 IBIAS3.n344 7.86204
R284 IBIAS3.n237 IBIAS3.n232 7.86204
R285 IBIAS3.n69 IBIAS3.n63 7.76845
R286 IBIAS3.n90 IBIAS3.n84 7.76845
R287 IBIAS3.n291 IBIAS3.n285 7.76845
R288 IBIAS3.n312 IBIAS3.n306 7.76845
R289 IBIAS3.n179 IBIAS3.n173 7.76845
R290 IBIAS3.n200 IBIAS3.n194 7.76845
R291 IBIAS3.n29 IBIAS3.n24 7.67486
R292 IBIAS3.n111 IBIAS3.n105 7.67486
R293 IBIAS3.n251 IBIAS3.n246 7.67486
R294 IBIAS3.n333 IBIAS3.n327 7.67486
R295 IBIAS3.n139 IBIAS3.n134 7.67486
R296 IBIAS3.n221 IBIAS3.n215 7.67486
R297 IBIAS3.n48 IBIAS3.n42 7.58127
R298 IBIAS3.n270 IBIAS3.n264 7.58127
R299 IBIAS3.n158 IBIAS3.n152 7.58127
R300 IBIAS3.n48 IBIAS3.n47 7.39409
R301 IBIAS3.n270 IBIAS3.n269 7.39409
R302 IBIAS3.n158 IBIAS3.n157 7.39409
R303 IBIAS3.n29 IBIAS3.n28 7.3005
R304 IBIAS3.n111 IBIAS3.n110 7.3005
R305 IBIAS3.n251 IBIAS3.n250 7.3005
R306 IBIAS3.n333 IBIAS3.n332 7.3005
R307 IBIAS3.n139 IBIAS3.n138 7.3005
R308 IBIAS3.n221 IBIAS3.n220 7.3005
R309 IBIAS3.n69 IBIAS3.n68 7.20691
R310 IBIAS3.n90 IBIAS3.n89 7.20691
R311 IBIAS3.n291 IBIAS3.n290 7.20691
R312 IBIAS3.n312 IBIAS3.n311 7.20691
R313 IBIAS3.n179 IBIAS3.n178 7.20691
R314 IBIAS3.n200 IBIAS3.n199 7.20691
R315 IBIAS3.n127 IBIAS3.n126 7.11332
R316 IBIAS3.n349 IBIAS3.n348 7.11332
R317 IBIAS3.n237 IBIAS3.n236 7.11332
R318 IBIAS3.n30 IBIAS3.n29 4.30071
R319 IBIAS3.n252 IBIAS3.n251 4.30071
R320 IBIAS3.n128 IBIAS3.n127 4.23696
R321 IBIAS3.n350 IBIAS3.n349 4.23696
R322 IBIAS3.n238 IBIAS3.n237 4.23696
R323 IBIAS3.n140 IBIAS3.n139 4.2258
R324 IBIAS3.n49 IBIAS3.n48 4.0005
R325 IBIAS3.n70 IBIAS3.n69 4.0005
R326 IBIAS3.n91 IBIAS3.n90 4.0005
R327 IBIAS3.n112 IBIAS3.n111 4.0005
R328 IBIAS3.n271 IBIAS3.n270 4.0005
R329 IBIAS3.n292 IBIAS3.n291 4.0005
R330 IBIAS3.n313 IBIAS3.n312 4.0005
R331 IBIAS3.n334 IBIAS3.n333 4.0005
R332 IBIAS3.n222 IBIAS3.n221 4.0005
R333 IBIAS3.n201 IBIAS3.n200 4.0005
R334 IBIAS3.n180 IBIAS3.n179 4.0005
R335 IBIAS3.n159 IBIAS3.n158 4.0005
R336 IBIAS3.n372 IBIAS3.n371 2.61298
R337 IBIAS3.n412 IBIAS3.n411 2.61298
R338 IBIAS3.n241 IBIAS3.n240 1.89565
R339 IBIAS3.n395 IBIAS3.n394 1.82618
R340 IBIAS3.n11 IBIAS3.n10 1.82586
R341 IBIAS3.n406 IBIAS3.t76 1.73227
R342 IBIAS3.n365 IBIAS3.n364 1.73042
R343 IBIAS3.n34 IBIAS3.n33 1.63706
R344 IBIAS3.n256 IBIAS3.n255 1.63706
R345 IBIAS3.n76 IBIAS3.n75 1.6369
R346 IBIAS3.n298 IBIAS3.n297 1.6369
R347 IBIAS3.n186 IBIAS3.n185 1.6369
R348 IBIAS3.n55 IBIAS3.n54 1.63685
R349 IBIAS3.n277 IBIAS3.n276 1.63685
R350 IBIAS3.n165 IBIAS3.n164 1.63685
R351 IBIAS3.n97 IBIAS3.n96 1.63682
R352 IBIAS3.n319 IBIAS3.n318 1.63682
R353 IBIAS3.n207 IBIAS3.n206 1.63682
R354 IBIAS3.n228 IBIAS3.n227 1.63483
R355 IBIAS3.n353 IBIAS3.n352 1.44752
R356 IBIAS3.n363 IBIAS3.n362 1.4267
R357 IBIAS3.n405 IBIAS3.n404 1.4257
R358 IBIAS3.n37 IBIAS3.n31 1.20341
R359 IBIAS3.n259 IBIAS3.n253 1.20341
R360 IBIAS3.n147 IBIAS3.n141 1.20341
R361 IBIAS3.n118 IBIAS3.n117 1.18592
R362 IBIAS3.n340 IBIAS3.n339 1.18592
R363 IBIAS3.n144 IBIAS3.n143 1.18481
R364 IBIAS3.n402 IBIAS3.n386 1.16943
R365 IBIAS3.n18 IBIAS3.n2 1.16928
R366 IBIAS3.n418 IBIAS3.n405 1.14806
R367 IBIAS3.n378 IBIAS3.n363 1.14599
R368 IBIAS3.n17 IBIAS3.n16 1.1255
R369 IBIAS3.n14 IBIAS3.n13 1.1255
R370 IBIAS3.n8 IBIAS3.n7 1.1255
R371 IBIAS3.n401 IBIAS3.n400 1.1255
R372 IBIAS3.n398 IBIAS3.n397 1.1255
R373 IBIAS3.n392 IBIAS3.n391 1.1255
R374 IBIAS3.n130 IBIAS3.n129 1.1255
R375 IBIAS3.n52 IBIAS3.n51 1.1255
R376 IBIAS3.n58 IBIAS3.n57 1.1255
R377 IBIAS3.n73 IBIAS3.n72 1.1255
R378 IBIAS3.n79 IBIAS3.n78 1.1255
R379 IBIAS3.n94 IBIAS3.n93 1.1255
R380 IBIAS3.n100 IBIAS3.n99 1.1255
R381 IBIAS3.n115 IBIAS3.n114 1.1255
R382 IBIAS3.n37 IBIAS3.n36 1.1255
R383 IBIAS3.n352 IBIAS3.n351 1.1255
R384 IBIAS3.n274 IBIAS3.n273 1.1255
R385 IBIAS3.n280 IBIAS3.n279 1.1255
R386 IBIAS3.n295 IBIAS3.n294 1.1255
R387 IBIAS3.n301 IBIAS3.n300 1.1255
R388 IBIAS3.n316 IBIAS3.n315 1.1255
R389 IBIAS3.n322 IBIAS3.n321 1.1255
R390 IBIAS3.n337 IBIAS3.n336 1.1255
R391 IBIAS3.n259 IBIAS3.n258 1.1255
R392 IBIAS3.n210 IBIAS3.n209 1.1255
R393 IBIAS3.n204 IBIAS3.n203 1.1255
R394 IBIAS3.n189 IBIAS3.n188 1.1255
R395 IBIAS3.n183 IBIAS3.n182 1.1255
R396 IBIAS3.n168 IBIAS3.n167 1.1255
R397 IBIAS3.n162 IBIAS3.n161 1.1255
R398 IBIAS3.n147 IBIAS3.n146 1.1255
R399 IBIAS3.n240 IBIAS3.n239 1.1255
R400 IBIAS3.n225 IBIAS3.n224 1.1255
R401 IBIAS3.n377 IBIAS3.n376 1.1255
R402 IBIAS3.n374 IBIAS3.n373 1.1255
R403 IBIAS3.n368 IBIAS3.n367 1.1255
R404 IBIAS3.n417 IBIAS3.n416 1.1255
R405 IBIAS3.n414 IBIAS3.n413 1.1255
R406 IBIAS3.n409 IBIAS3.n408 1.1255
R407 IBIAS3.n383 IBIAS3.n18 1.12215
R408 IBIAS3.n358 IBIAS3.n357 1.1167
R409 IBIAS3.n403 IBIAS3.n402 1.0896
R410 IBIAS3.n386 IBIAS3.n385 1.06753
R411 IBIAS3.n2 IBIAS3.n1 1.06753
R412 IBIAS3 IBIAS3.n403 1.02107
R413 IBIAS3.n241 IBIAS3.n130 1.01814
R414 IBIAS3.n368 IBIAS3.n365 0.925791
R415 IBIAS3.n8 IBIAS3.n5 0.92452
R416 IBIAS3.n392 IBIAS3.n389 0.92446
R417 IBIAS3.n409 IBIAS3.n406 0.924202
R418 IBIAS3.n389 IBIAS3.n388 0.912989
R419 IBIAS3.n5 IBIAS3.n4 0.912902
R420 IBIAS3.n380 IBIAS3.n379 0.895909
R421 IBIAS3.n404 IBIAS3.t69 0.8195
R422 IBIAS3.n411 IBIAS3.t73 0.8195
R423 IBIAS3.n1 IBIAS3.t64 0.8195
R424 IBIAS3.n1 IBIAS3.n0 0.8195
R425 IBIAS3.n10 IBIAS3.t62 0.8195
R426 IBIAS3.n10 IBIAS3.n9 0.8195
R427 IBIAS3.n4 IBIAS3.t66 0.8195
R428 IBIAS3.n4 IBIAS3.n3 0.8195
R429 IBIAS3.n385 IBIAS3.t71 0.8195
R430 IBIAS3.n385 IBIAS3.n384 0.8195
R431 IBIAS3.n394 IBIAS3.t74 0.8195
R432 IBIAS3.n394 IBIAS3.n393 0.8195
R433 IBIAS3.n388 IBIAS3.t61 0.8195
R434 IBIAS3.n388 IBIAS3.n387 0.8195
R435 IBIAS3.n362 IBIAS3.n361 0.8195
R436 IBIAS3.n371 IBIAS3.n370 0.8195
R437 IBIAS3.n359 IBIAS3.n358 0.7655
R438 IBIAS3.n33 IBIAS3.t19 0.607167
R439 IBIAS3.n33 IBIAS3.n32 0.607167
R440 IBIAS3.n54 IBIAS3.t13 0.607167
R441 IBIAS3.n54 IBIAS3.n53 0.607167
R442 IBIAS3.n75 IBIAS3.t15 0.607167
R443 IBIAS3.n75 IBIAS3.n74 0.607167
R444 IBIAS3.n96 IBIAS3.t17 0.607167
R445 IBIAS3.n96 IBIAS3.n95 0.607167
R446 IBIAS3.n117 IBIAS3.t31 0.607167
R447 IBIAS3.n117 IBIAS3.n116 0.607167
R448 IBIAS3.n255 IBIAS3.t25 0.607167
R449 IBIAS3.n255 IBIAS3.n254 0.607167
R450 IBIAS3.n276 IBIAS3.t33 0.607167
R451 IBIAS3.n276 IBIAS3.n275 0.607167
R452 IBIAS3.n297 IBIAS3.t7 0.607167
R453 IBIAS3.n297 IBIAS3.n296 0.607167
R454 IBIAS3.n318 IBIAS3.t11 0.607167
R455 IBIAS3.n318 IBIAS3.n317 0.607167
R456 IBIAS3.n339 IBIAS3.t29 0.607167
R457 IBIAS3.n339 IBIAS3.n338 0.607167
R458 IBIAS3.n164 IBIAS3.t27 0.607167
R459 IBIAS3.n164 IBIAS3.n163 0.607167
R460 IBIAS3.n185 IBIAS3.t21 0.607167
R461 IBIAS3.n185 IBIAS3.n184 0.607167
R462 IBIAS3.n206 IBIAS3.t23 0.607167
R463 IBIAS3.n206 IBIAS3.n205 0.607167
R464 IBIAS3.n227 IBIAS3.t35 0.607167
R465 IBIAS3.n227 IBIAS3.n226 0.607167
R466 IBIAS3.n143 IBIAS3.t9 0.607167
R467 IBIAS3.n143 IBIAS3.n142 0.607167
R468 IBIAS3.n379 IBIAS3.n378 0.547622
R469 IBIAS3.n115 IBIAS3.n100 0.433037
R470 IBIAS3.n337 IBIAS3.n322 0.433037
R471 IBIAS3.n225 IBIAS3.n210 0.433037
R472 IBIAS3.n52 IBIAS3.n37 0.426993
R473 IBIAS3.n274 IBIAS3.n259 0.426993
R474 IBIAS3.n162 IBIAS3.n147 0.426993
R475 IBIAS3.n94 IBIAS3.n79 0.420948
R476 IBIAS3.n316 IBIAS3.n301 0.420948
R477 IBIAS3.n204 IBIAS3.n189 0.420948
R478 IBIAS3.n73 IBIAS3.n58 0.414231
R479 IBIAS3.n295 IBIAS3.n280 0.414231
R480 IBIAS3.n183 IBIAS3.n168 0.414231
R481 IBIAS3.n17 IBIAS3.n14 0.372342
R482 IBIAS3.n401 IBIAS3.n398 0.372342
R483 IBIAS3.n377 IBIAS3.n374 0.372342
R484 IBIAS3.n417 IBIAS3.n414 0.372342
R485 IBIAS3.n223 IBIAS3.n222 0.350735
R486 IBIAS3.n242 IBIAS3.n241 0.335978
R487 IBIAS3.n92 IBIAS3.n91 0.320899
R488 IBIAS3.n314 IBIAS3.n313 0.320899
R489 IBIAS3.n202 IBIAS3.n201 0.320899
R490 IBIAS3.n50 IBIAS3.n49 0.318657
R491 IBIAS3.n272 IBIAS3.n271 0.318657
R492 IBIAS3.n160 IBIAS3.n159 0.318657
R493 IBIAS3.n71 IBIAS3.n70 0.314173
R494 IBIAS3.n293 IBIAS3.n292 0.314173
R495 IBIAS3.n181 IBIAS3.n180 0.314173
R496 IBIAS3.n403 IBIAS3.n383 0.264793
R497 IBIAS3.n113 IBIAS3.n112 0.259738
R498 IBIAS3.n335 IBIAS3.n334 0.259738
R499 IBIAS3 IBIAS3.n418 0.197079
R500 IBIAS3.n36 IBIAS3.n35 0.192197
R501 IBIAS3.n258 IBIAS3.n257 0.192197
R502 IBIAS3.n146 IBIAS3.n145 0.192197
R503 IBIAS3.n78 IBIAS3.n77 0.183344
R504 IBIAS3.n300 IBIAS3.n299 0.183344
R505 IBIAS3.n188 IBIAS3.n187 0.183344
R506 IBIAS3.n57 IBIAS3.n56 0.180394
R507 IBIAS3.n279 IBIAS3.n278 0.180394
R508 IBIAS3.n167 IBIAS3.n166 0.180394
R509 IBIAS3.n99 IBIAS3.n98 0.178918
R510 IBIAS3.n321 IBIAS3.n320 0.178918
R511 IBIAS3.n209 IBIAS3.n208 0.178918
R512 IBIAS3.n114 IBIAS3.n113 0.172302
R513 IBIAS3.n336 IBIAS3.n335 0.172302
R514 IBIAS3.n129 IBIAS3.n128 0.161213
R515 IBIAS3.n351 IBIAS3.n350 0.161213
R516 IBIAS3.n239 IBIAS3.n238 0.161213
R517 IBIAS3.n141 IBIAS3.n140 0.141318
R518 IBIAS3.n383 IBIAS3.n382 0.117852
R519 IBIAS3.n18 IBIAS3.n17 0.0920789
R520 IBIAS3.n14 IBIAS3.n8 0.0920789
R521 IBIAS3.n402 IBIAS3.n401 0.0920789
R522 IBIAS3.n398 IBIAS3.n392 0.0920789
R523 IBIAS3.n378 IBIAS3.n377 0.0920789
R524 IBIAS3.n374 IBIAS3.n368 0.0920789
R525 IBIAS3.n418 IBIAS3.n417 0.0920789
R526 IBIAS3.n414 IBIAS3.n409 0.0920789
R527 IBIAS3.n13 IBIAS3.n12 0.0860505
R528 IBIAS3.n397 IBIAS3.n396 0.0860505
R529 IBIAS3.n16 IBIAS3.n15 0.0806418
R530 IBIAS3.n400 IBIAS3.n399 0.0806418
R531 IBIAS3.n224 IBIAS3.n223 0.0793147
R532 IBIAS3.n373 IBIAS3.n369 0.0785711
R533 IBIAS3.n58 IBIAS3.n52 0.0784104
R534 IBIAS3.n79 IBIAS3.n73 0.0784104
R535 IBIAS3.n100 IBIAS3.n94 0.0784104
R536 IBIAS3.n130 IBIAS3.n115 0.0784104
R537 IBIAS3.n280 IBIAS3.n274 0.0784104
R538 IBIAS3.n301 IBIAS3.n295 0.0784104
R539 IBIAS3.n322 IBIAS3.n316 0.0784104
R540 IBIAS3.n352 IBIAS3.n337 0.0784104
R541 IBIAS3.n168 IBIAS3.n162 0.0784104
R542 IBIAS3.n189 IBIAS3.n183 0.0784104
R543 IBIAS3.n210 IBIAS3.n204 0.0784104
R544 IBIAS3.n240 IBIAS3.n225 0.0784104
R545 IBIAS3.n93 IBIAS3.n92 0.0713702
R546 IBIAS3.n315 IBIAS3.n314 0.0713702
R547 IBIAS3.n203 IBIAS3.n202 0.0713702
R548 IBIAS3.n51 IBIAS3.n50 0.0707069
R549 IBIAS3.n273 IBIAS3.n272 0.0707069
R550 IBIAS3.n161 IBIAS3.n160 0.0707069
R551 IBIAS3.n413 IBIAS3.n410 0.0703936
R552 IBIAS3.n72 IBIAS3.n71 0.0693796
R553 IBIAS3.n294 IBIAS3.n293 0.0693796
R554 IBIAS3.n182 IBIAS3.n181 0.0693796
R555 IBIAS3.n31 IBIAS3.n30 0.0653931
R556 IBIAS3.n253 IBIAS3.n252 0.0653931
R557 IBIAS3.n129 IBIAS3.n118 0.0570651
R558 IBIAS3.n351 IBIAS3.n340 0.0570651
R559 IBIAS3.n146 IBIAS3.n144 0.0483228
R560 IBIAS3.n391 IBIAS3.n390 0.0459639
R561 IBIAS3.n7 IBIAS3.n6 0.0450361
R562 IBIAS3.n13 IBIAS3.n11 0.0432191
R563 IBIAS3.n397 IBIAS3.n395 0.0425445
R564 IBIAS3.n239 IBIAS3.n228 0.0381228
R565 IBIAS3.n356 IBIAS3.n355 0.038
R566 IBIAS3.n416 IBIAS3.n415 0.0347237
R567 IBIAS3.n376 IBIAS3.n375 0.0318359
R568 IBIAS3.n99 IBIAS3.n97 0.0311692
R569 IBIAS3.n321 IBIAS3.n319 0.0311692
R570 IBIAS3.n209 IBIAS3.n207 0.0311692
R571 IBIAS3.n57 IBIAS3.n55 0.0305887
R572 IBIAS3.n279 IBIAS3.n277 0.0305887
R573 IBIAS3.n167 IBIAS3.n165 0.0305887
R574 IBIAS3.n78 IBIAS3.n76 0.0294265
R575 IBIAS3.n300 IBIAS3.n298 0.0294265
R576 IBIAS3.n188 IBIAS3.n186 0.0294265
R577 IBIAS3.n381 IBIAS3.n380 0.0274649
R578 IBIAS3.n382 IBIAS3.n381 0.0262757
R579 IBIAS3.n36 IBIAS3.n34 0.0262212
R580 IBIAS3.n258 IBIAS3.n256 0.0262212
R581 IBIAS3.n355 IBIAS3.n354 0.0258619
R582 IBIAS3.n413 IBIAS3.n412 0.0233115
R583 IBIAS3.n373 IBIAS3.n372 0.0233115
R584 IBIAS3.n379 IBIAS3.n360 0.0201693
R585 IBIAS3.n20 IBIAS3.n19 0.0201693
R586 IBIAS3.n408 IBIAS3.n407 0.0198639
R587 IBIAS3.n357 IBIAS3.n242 0.019595
R588 IBIAS3.n357 IBIAS3.n356 0.019595
R589 IBIAS3.n367 IBIAS3.n366 0.0179463
R590 IBIAS3.n354 IBIAS3.n353 0.0134309
R591 IBIAS3.n358 IBIAS3.n20 0.0105847
R592 IBIAS3.n360 IBIAS3.n359 0.0105847
R593 OUTo.n1 OUTo.t163 5.17489
R594 OUTo.n23 OUTo.t142 5.15289
R595 OUTo.n18 OUTo.t120 4.43476
R596 OUTo.n8 OUTo.t141 3.01175
R597 OUTo.n9 OUTo.n8 2.8714
R598 OUTo.n283 OUTo.n282 2.58542
R599 OUTo.n430 OUTo.n429 2.58542
R600 OUTo.n28 OUTo.n24 2.28927
R601 OUTo.n12 OUTo.n3 2.28927
R602 OUTo.n267 OUTo.n266 2.25086
R603 OUTo.n279 OUTo.n245 2.25086
R604 OUTo.n237 OUTo.n236 2.25086
R605 OUTo.n274 OUTo.n273 2.25086
R606 OUTo.n318 OUTo.n317 2.25086
R607 OUTo.n329 OUTo.n328 2.25086
R608 OUTo.n414 OUTo.n413 2.25086
R609 OUTo.n426 OUTo.n392 2.25086
R610 OUTo.n384 OUTo.n383 2.25086
R611 OUTo.n421 OUTo.n420 2.25086
R612 OUTo.n465 OUTo.n464 2.25086
R613 OUTo.n476 OUTo.n475 2.25086
R614 OUTo.n12 OUTo.n11 2.2505
R615 OUTo.n16 OUTo.n15 2.2505
R616 OUTo.n28 OUTo.n27 2.2505
R617 OUTo.n285 OUTo.n284 2.2473
R618 OUTo.n224 OUTo.n188 2.2473
R619 OUTo.n275 OUTo.n250 2.2473
R620 OUTo.n332 OUTo.n331 2.2473
R621 OUTo.n432 OUTo.n431 2.2473
R622 OUTo.n371 OUTo.n335 2.2473
R623 OUTo.n422 OUTo.n397 2.2473
R624 OUTo.n479 OUTo.n478 2.2473
R625 OUTo.n262 OUTo.n261 2.2473
R626 OUTo.n242 OUTo.n241 2.2473
R627 OUTo.n231 OUTo.n230 2.2473
R628 OUTo.n321 OUTo.n320 2.2473
R629 OUTo.n409 OUTo.n408 2.2473
R630 OUTo.n389 OUTo.n388 2.2473
R631 OUTo.n378 OUTo.n377 2.2473
R632 OUTo.n468 OUTo.n467 2.2473
R633 OUTo.n249 OUTo.n248 1.8413
R634 OUTo.n396 OUTo.n395 1.8413
R635 OUTo.n167 OUTo.n166 1.63699
R636 OUTo.n660 OUTo.n659 1.63699
R637 OUTo.n176 OUTo.n175 1.63689
R638 OUTo.n669 OUTo.n668 1.63689
R639 OUTo.n765 OUTo.n764 1.63687
R640 OUTo.n78 OUTo.n77 1.63687
R641 OUTo.n613 OUTo.n612 1.63687
R642 OUTo.n774 OUTo.n773 1.63672
R643 OUTo.n87 OUTo.n86 1.63672
R644 OUTo.n622 OUTo.n621 1.63672
R645 OUTo.n727 OUTo.n726 1.63667
R646 OUTo.n736 OUTo.n735 1.63667
R647 OUTo.n575 OUTo.n574 1.63667
R648 OUTo.n584 OUTo.n583 1.63667
R649 OUTo.n41 OUTo.n40 1.63667
R650 OUTo.n50 OUTo.n49 1.63667
R651 OUTo.n537 OUTo.n536 1.63664
R652 OUTo.n121 OUTo.n120 1.63664
R653 OUTo.n689 OUTo.n688 1.63664
R654 OUTo.n158 OUTo.n157 1.63649
R655 OUTo.n651 OUTo.n650 1.63649
R656 OUTo.n500 OUTo.n499 1.63649
R657 OUTo.n555 OUTo.n554 1.63642
R658 OUTo.n139 OUTo.n138 1.63642
R659 OUTo.n707 OUTo.n706 1.63642
R660 OUTo.n783 OUTo.n782 1.63582
R661 OUTo.n96 OUTo.n95 1.63582
R662 OUTo.n631 OUTo.n630 1.63582
R663 OUTo.n546 OUTo.n545 1.63562
R664 OUTo.n130 OUTo.n129 1.63562
R665 OUTo.n698 OUTo.n697 1.63562
R666 OUTo.n745 OUTo.n744 1.63523
R667 OUTo.n593 OUTo.n592 1.63523
R668 OUTo.n59 OUTo.n58 1.63523
R669 OUTo.n518 OUTo.n517 1.63265
R670 OUTo.n509 OUTo.n508 1.63126
R671 OUTo.n213 OUTo.n212 1.49783
R672 OUTo.n201 OUTo.n200 1.49783
R673 OUTo.n295 OUTo.n294 1.49783
R674 OUTo.n305 OUTo.n304 1.49783
R675 OUTo.n360 OUTo.n359 1.49783
R676 OUTo.n348 OUTo.n347 1.49783
R677 OUTo.n442 OUTo.n441 1.49783
R678 OUTo.n452 OUTo.n451 1.49783
R679 OUTo.n206 OUTo.n205 1.49759
R680 OUTo.n221 OUTo.n220 1.49759
R681 OUTo.n310 OUTo.n309 1.49759
R682 OUTo.n299 OUTo.n298 1.49759
R683 OUTo.n353 OUTo.n352 1.49759
R684 OUTo.n368 OUTo.n367 1.49759
R685 OUTo.n457 OUTo.n456 1.49759
R686 OUTo.n446 OUTo.n445 1.49759
R687 OUTo.n204 OUTo.n203 1.42962
R688 OUTo.n351 OUTo.n350 1.42962
R689 OUTo.n211 OUTo.n210 1.42935
R690 OUTo.n229 OUTo.n228 1.42935
R691 OUTo.n358 OUTo.n357 1.42935
R692 OUTo.n376 OUTo.n375 1.42935
R693 OUTo.n308 OUTo.n307 1.42817
R694 OUTo.n327 OUTo.n326 1.42817
R695 OUTo.n455 OUTo.n454 1.42817
R696 OUTo.n474 OUTo.n473 1.42817
R697 OUTo.n293 OUTo.n292 1.42798
R698 OUTo.n440 OUTo.n439 1.42798
R699 OUTo.n566 OUTo.n528 1.34531
R700 OUTo.n196 OUTo.n195 1.29129
R701 OUTo.n216 OUTo.n215 1.29129
R702 OUTo.n253 OUTo.n252 1.29129
R703 OUTo.n343 OUTo.n342 1.29129
R704 OUTo.n363 OUTo.n362 1.29129
R705 OUTo.n400 OUTo.n399 1.29129
R706 OUTo.n680 OUTo.n679 1.2545
R707 OUTo.n718 OUTo.n717 1.25382
R708 OUTo.n566 OUTo.n565 1.25338
R709 OUTo.n756 OUTo.n755 1.2527
R710 OUTo.n604 OUTo.n603 1.2527
R711 OUTo.n794 OUTo.n793 1.25047
R712 OUTo.n642 OUTo.n641 1.25047
R713 OUTo.n527 OUTo.n526 1.24873
R714 OUTo.n793 OUTo.n792 1.17148
R715 OUTo.n106 OUTo.n105 1.17148
R716 OUTo.n641 OUTo.n640 1.17148
R717 OUTo.n755 OUTo.n754 1.17097
R718 OUTo.n603 OUTo.n602 1.17097
R719 OUTo.n69 OUTo.n68 1.17097
R720 OUTo.n565 OUTo.n564 1.17063
R721 OUTo.n149 OUTo.n148 1.17063
R722 OUTo.n717 OUTo.n716 1.17063
R723 OUTo.n186 OUTo.n185 1.17046
R724 OUTo.n679 OUTo.n678 1.17046
R725 OUTo.n528 OUTo.n527 1.15251
R726 OUTo.n257 OUTo.n254 1.12719
R727 OUTo.n404 OUTo.n401 1.12719
R728 OUTo.n257 OUTo.n256 1.12669
R729 OUTo.n404 OUTo.n403 1.12669
R730 OUTo.n730 OUTo.n729 1.1255
R731 OUTo.n724 OUTo.n723 1.1255
R732 OUTo.n739 OUTo.n738 1.1255
R733 OUTo.n733 OUTo.n732 1.1255
R734 OUTo.n748 OUTo.n747 1.1255
R735 OUTo.n742 OUTo.n741 1.1255
R736 OUTo.n751 OUTo.n750 1.1255
R737 OUTo.n578 OUTo.n577 1.1255
R738 OUTo.n572 OUTo.n571 1.1255
R739 OUTo.n587 OUTo.n586 1.1255
R740 OUTo.n581 OUTo.n580 1.1255
R741 OUTo.n596 OUTo.n595 1.1255
R742 OUTo.n590 OUTo.n589 1.1255
R743 OUTo.n599 OUTo.n598 1.1255
R744 OUTo.n540 OUTo.n539 1.1255
R745 OUTo.n534 OUTo.n533 1.1255
R746 OUTo.n549 OUTo.n548 1.1255
R747 OUTo.n543 OUTo.n542 1.1255
R748 OUTo.n558 OUTo.n557 1.1255
R749 OUTo.n552 OUTo.n551 1.1255
R750 OUTo.n561 OUTo.n560 1.1255
R751 OUTo.n768 OUTo.n767 1.1255
R752 OUTo.n762 OUTo.n761 1.1255
R753 OUTo.n777 OUTo.n776 1.1255
R754 OUTo.n771 OUTo.n770 1.1255
R755 OUTo.n786 OUTo.n785 1.1255
R756 OUTo.n780 OUTo.n779 1.1255
R757 OUTo.n789 OUTo.n788 1.1255
R758 OUTo.n81 OUTo.n80 1.1255
R759 OUTo.n75 OUTo.n74 1.1255
R760 OUTo.n90 OUTo.n89 1.1255
R761 OUTo.n84 OUTo.n83 1.1255
R762 OUTo.n99 OUTo.n98 1.1255
R763 OUTo.n93 OUTo.n92 1.1255
R764 OUTo.n102 OUTo.n101 1.1255
R765 OUTo.n44 OUTo.n43 1.1255
R766 OUTo.n38 OUTo.n37 1.1255
R767 OUTo.n53 OUTo.n52 1.1255
R768 OUTo.n47 OUTo.n46 1.1255
R769 OUTo.n62 OUTo.n61 1.1255
R770 OUTo.n56 OUTo.n55 1.1255
R771 OUTo.n65 OUTo.n64 1.1255
R772 OUTo.n124 OUTo.n123 1.1255
R773 OUTo.n118 OUTo.n117 1.1255
R774 OUTo.n133 OUTo.n132 1.1255
R775 OUTo.n127 OUTo.n126 1.1255
R776 OUTo.n142 OUTo.n141 1.1255
R777 OUTo.n136 OUTo.n135 1.1255
R778 OUTo.n145 OUTo.n144 1.1255
R779 OUTo.n161 OUTo.n160 1.1255
R780 OUTo.n155 OUTo.n154 1.1255
R781 OUTo.n170 OUTo.n169 1.1255
R782 OUTo.n164 OUTo.n163 1.1255
R783 OUTo.n179 OUTo.n178 1.1255
R784 OUTo.n173 OUTo.n172 1.1255
R785 OUTo.n182 OUTo.n181 1.1255
R786 OUTo.n616 OUTo.n615 1.1255
R787 OUTo.n610 OUTo.n609 1.1255
R788 OUTo.n625 OUTo.n624 1.1255
R789 OUTo.n619 OUTo.n618 1.1255
R790 OUTo.n634 OUTo.n633 1.1255
R791 OUTo.n628 OUTo.n627 1.1255
R792 OUTo.n637 OUTo.n636 1.1255
R793 OUTo.n654 OUTo.n653 1.1255
R794 OUTo.n648 OUTo.n647 1.1255
R795 OUTo.n663 OUTo.n662 1.1255
R796 OUTo.n657 OUTo.n656 1.1255
R797 OUTo.n672 OUTo.n671 1.1255
R798 OUTo.n666 OUTo.n665 1.1255
R799 OUTo.n675 OUTo.n674 1.1255
R800 OUTo.n692 OUTo.n691 1.1255
R801 OUTo.n686 OUTo.n685 1.1255
R802 OUTo.n701 OUTo.n700 1.1255
R803 OUTo.n695 OUTo.n694 1.1255
R804 OUTo.n710 OUTo.n709 1.1255
R805 OUTo.n704 OUTo.n703 1.1255
R806 OUTo.n713 OUTo.n712 1.1255
R807 OUTo.n497 OUTo.n496 1.1255
R808 OUTo.n503 OUTo.n502 1.1255
R809 OUTo.n506 OUTo.n505 1.1255
R810 OUTo.n512 OUTo.n511 1.1255
R811 OUTo.n515 OUTo.n514 1.1255
R812 OUTo.n521 OUTo.n520 1.1255
R813 OUTo.n524 OUTo.n523 1.1255
R814 OUTo.n11 OUTo.n10 1.1255
R815 OUTo.n798 OUTo.n491 1.1255
R816 OUTo.n112 OUTo.n111 1.1255
R817 OUTo.n24 OUTo.n23 1.12469
R818 OUTo.n3 OUTo.n1 1.12241
R819 OUTo.n240 OUTo.n239 1.06972
R820 OUTo.n387 OUTo.n386 1.06972
R821 OUTo.n316 OUTo.n315 1.06956
R822 OUTo.n463 OUTo.n462 1.06956
R823 OUTo.n762 OUTo.n759 1.05314
R824 OUTo.n75 OUTo.n72 1.05314
R825 OUTo.n610 OUTo.n607 1.05314
R826 OUTo.n724 OUTo.n721 1.04551
R827 OUTo.n572 OUTo.n569 1.04551
R828 OUTo.n38 OUTo.n35 1.04551
R829 OUTo.n155 OUTo.n152 1.03013
R830 OUTo.n648 OUTo.n645 1.03013
R831 OUTo.n497 OUTo.n494 1.02996
R832 OUTo.n534 OUTo.n531 1.02977
R833 OUTo.n118 OUTo.n115 1.02977
R834 OUTo.n686 OUTo.n683 1.02977
R835 OUTo.n185 OUTo.n184 0.964358
R836 OUTo.n678 OUTo.n677 0.964358
R837 OUTo.n564 OUTo.n563 0.96424
R838 OUTo.n148 OUTo.n147 0.96424
R839 OUTo.n716 OUTo.n715 0.96424
R840 OUTo.n754 OUTo.n753 0.964059
R841 OUTo.n602 OUTo.n601 0.964059
R842 OUTo.n68 OUTo.n67 0.964059
R843 OUTo.n792 OUTo.n791 0.963815
R844 OUTo.n105 OUTo.n104 0.963815
R845 OUTo.n640 OUTo.n639 0.963815
R846 OUTo.n192 OUTo.n191 0.915267
R847 OUTo.n339 OUTo.n338 0.915267
R848 OUTo.n289 OUTo.n288 0.91305
R849 OUTo.n436 OUTo.n435 0.91305
R850 OUTo.n494 OUTo.n493 0.809647
R851 OUTo.n531 OUTo.n530 0.80933
R852 OUTo.n115 OUTo.n114 0.80933
R853 OUTo.n683 OUTo.n682 0.80933
R854 OUTo.n152 OUTo.n151 0.808908
R855 OUTo.n645 OUTo.n644 0.808908
R856 OUTo.n759 OUTo.n758 0.806374
R857 OUTo.n72 OUTo.n71 0.806374
R858 OUTo.n607 OUTo.n606 0.806374
R859 OUTo.n721 OUTo.n720 0.80586
R860 OUTo.n569 OUTo.n568 0.80586
R861 OUTo.n35 OUTo.n34 0.80586
R862 OUTo.n290 OUTo.n289 0.745852
R863 OUTo.n437 OUTo.n436 0.745852
R864 OUTo.n193 OUTo.n192 0.743777
R865 OUTo.n340 OUTo.n339 0.743777
R866 OUTo.n192 OUTo.n189 0.680835
R867 OUTo.n339 OUTo.n336 0.680835
R868 OUTo.n487 OUTo.n186 0.665425
R869 OUTo.n490 OUTo.n149 0.664754
R870 OUTo.n110 OUTo.n69 0.66341
R871 OUTo.n107 OUTo.n106 0.661396
R872 OUTo.n297 OUTo.n296 0.621961
R873 OUTo.n444 OUTo.n443 0.621961
R874 OUTo.n303 OUTo.n302 0.619651
R875 OUTo.n450 OUTo.n449 0.619651
R876 OUTo.n219 OUTo.n218 0.615708
R877 OUTo.n366 OUTo.n365 0.615708
R878 OUTo.n199 OUTo.n198 0.61192
R879 OUTo.n346 OUTo.n345 0.61192
R880 OUTo.n744 OUTo.t75 0.607167
R881 OUTo.n744 OUTo.n743 0.607167
R882 OUTo.n735 OUTo.t72 0.607167
R883 OUTo.n735 OUTo.n734 0.607167
R884 OUTo.n726 OUTo.t42 0.607167
R885 OUTo.n726 OUTo.n725 0.607167
R886 OUTo.n720 OUTo.t53 0.607167
R887 OUTo.n720 OUTo.n719 0.607167
R888 OUTo.n753 OUTo.t55 0.607167
R889 OUTo.n753 OUTo.n752 0.607167
R890 OUTo.n592 OUTo.t22 0.607167
R891 OUTo.n592 OUTo.n591 0.607167
R892 OUTo.n583 OUTo.t20 0.607167
R893 OUTo.n583 OUTo.n582 0.607167
R894 OUTo.n574 OUTo.t58 0.607167
R895 OUTo.n574 OUTo.n573 0.607167
R896 OUTo.n568 OUTo.t43 0.607167
R897 OUTo.n568 OUTo.n567 0.607167
R898 OUTo.n601 OUTo.t62 0.607167
R899 OUTo.n601 OUTo.n600 0.607167
R900 OUTo.n554 OUTo.t48 0.607167
R901 OUTo.n554 OUTo.n553 0.607167
R902 OUTo.n545 OUTo.t45 0.607167
R903 OUTo.n545 OUTo.n544 0.607167
R904 OUTo.n536 OUTo.t19 0.607167
R905 OUTo.n536 OUTo.n535 0.607167
R906 OUTo.n530 OUTo.t56 0.607167
R907 OUTo.n530 OUTo.n529 0.607167
R908 OUTo.n563 OUTo.t30 0.607167
R909 OUTo.n563 OUTo.n562 0.607167
R910 OUTo.n782 OUTo.t44 0.607167
R911 OUTo.n782 OUTo.n781 0.607167
R912 OUTo.n773 OUTo.t40 0.607167
R913 OUTo.n773 OUTo.n772 0.607167
R914 OUTo.n764 OUTo.t60 0.607167
R915 OUTo.n764 OUTo.n763 0.607167
R916 OUTo.n758 OUTo.t78 0.607167
R917 OUTo.n758 OUTo.n757 0.607167
R918 OUTo.n791 OUTo.t27 0.607167
R919 OUTo.n791 OUTo.n790 0.607167
R920 OUTo.n95 OUTo.t32 0.607167
R921 OUTo.n95 OUTo.n94 0.607167
R922 OUTo.n86 OUTo.t29 0.607167
R923 OUTo.n86 OUTo.n85 0.607167
R924 OUTo.n77 OUTo.t67 0.607167
R925 OUTo.n77 OUTo.n76 0.607167
R926 OUTo.n71 OUTo.t70 0.607167
R927 OUTo.n71 OUTo.n70 0.607167
R928 OUTo.n104 OUTo.t76 0.607167
R929 OUTo.n104 OUTo.n103 0.607167
R930 OUTo.n58 OUTo.t68 0.607167
R931 OUTo.n58 OUTo.n57 0.607167
R932 OUTo.n49 OUTo.t64 0.607167
R933 OUTo.n49 OUTo.n48 0.607167
R934 OUTo.n40 OUTo.t31 0.607167
R935 OUTo.n40 OUTo.n39 0.607167
R936 OUTo.n34 OUTo.t61 0.607167
R937 OUTo.n34 OUTo.n33 0.607167
R938 OUTo.n67 OUTo.t47 0.607167
R939 OUTo.n67 OUTo.n66 0.607167
R940 OUTo.n138 OUTo.t28 0.607167
R941 OUTo.n138 OUTo.n137 0.607167
R942 OUTo.n129 OUTo.t26 0.607167
R943 OUTo.n129 OUTo.n128 0.607167
R944 OUTo.n120 OUTo.t74 0.607167
R945 OUTo.n120 OUTo.n119 0.607167
R946 OUTo.n114 OUTo.t57 0.607167
R947 OUTo.n114 OUTo.n113 0.607167
R948 OUTo.n147 OUTo.t71 0.607167
R949 OUTo.n147 OUTo.n146 0.607167
R950 OUTo.n175 OUTo.t41 0.607167
R951 OUTo.n175 OUTo.n174 0.607167
R952 OUTo.n166 OUTo.t38 0.607167
R953 OUTo.n166 OUTo.n165 0.607167
R954 OUTo.n157 OUTo.t52 0.607167
R955 OUTo.n157 OUTo.n156 0.607167
R956 OUTo.n151 OUTo.t34 0.607167
R957 OUTo.n151 OUTo.n150 0.607167
R958 OUTo.n184 OUTo.t25 0.607167
R959 OUTo.n184 OUTo.n183 0.607167
R960 OUTo.n630 OUTo.t51 0.607167
R961 OUTo.n630 OUTo.n629 0.607167
R962 OUTo.n621 OUTo.t49 0.607167
R963 OUTo.n621 OUTo.n620 0.607167
R964 OUTo.n612 OUTo.t73 0.607167
R965 OUTo.n612 OUTo.n611 0.607167
R966 OUTo.n606 OUTo.t69 0.607167
R967 OUTo.n606 OUTo.n605 0.607167
R968 OUTo.n639 OUTo.t35 0.607167
R969 OUTo.n639 OUTo.n638 0.607167
R970 OUTo.n668 OUTo.t50 0.607167
R971 OUTo.n668 OUTo.n667 0.607167
R972 OUTo.n659 OUTo.t46 0.607167
R973 OUTo.n659 OUTo.n658 0.607167
R974 OUTo.n650 OUTo.t66 0.607167
R975 OUTo.n650 OUTo.n649 0.607167
R976 OUTo.n644 OUTo.t23 0.607167
R977 OUTo.n644 OUTo.n643 0.607167
R978 OUTo.n677 OUTo.t33 0.607167
R979 OUTo.n677 OUTo.n676 0.607167
R980 OUTo.n706 OUTo.t39 0.607167
R981 OUTo.n706 OUTo.n705 0.607167
R982 OUTo.n697 OUTo.t37 0.607167
R983 OUTo.n697 OUTo.n696 0.607167
R984 OUTo.n688 OUTo.t65 0.607167
R985 OUTo.n688 OUTo.n687 0.607167
R986 OUTo.n682 OUTo.t63 0.607167
R987 OUTo.n682 OUTo.n681 0.607167
R988 OUTo.n715 OUTo.t24 0.607167
R989 OUTo.n715 OUTo.n714 0.607167
R990 OUTo.n493 OUTo.t77 0.607167
R991 OUTo.n493 OUTo.n492 0.607167
R992 OUTo.n499 OUTo.t21 0.607167
R993 OUTo.n499 OUTo.n498 0.607167
R994 OUTo.n508 OUTo.t54 0.607167
R995 OUTo.n508 OUTo.n507 0.607167
R996 OUTo.n517 OUTo.t59 0.607167
R997 OUTo.n517 OUTo.n516 0.607167
R998 OUTo.n526 OUTo.t36 0.607167
R999 OUTo.n526 OUTo.n525 0.607167
R1000 OUTo.n481 OUTo.n480 0.596332
R1001 OUTo.n30 OUTo.n29 0.553515
R1002 OUTo.n248 OUTo.t150 0.5465
R1003 OUTo.n248 OUTo.n247 0.5465
R1004 OUTo.n239 OUTo.t128 0.5465
R1005 OUTo.n239 OUTo.n238 0.5465
R1006 OUTo.n210 OUTo.t155 0.5465
R1007 OUTo.n210 OUTo.n209 0.5465
R1008 OUTo.n215 OUTo.t148 0.5465
R1009 OUTo.n215 OUTo.n214 0.5465
R1010 OUTo.n307 OUTo.t122 0.5465
R1011 OUTo.n307 OUTo.n306 0.5465
R1012 OUTo.n191 OUTo.t132 0.5465
R1013 OUTo.n191 OUTo.n190 0.5465
R1014 OUTo.n252 OUTo.t145 0.5465
R1015 OUTo.n252 OUTo.n251 0.5465
R1016 OUTo.n288 OUTo.t127 0.5465
R1017 OUTo.n288 OUTo.n287 0.5465
R1018 OUTo.n203 OUTo.t169 0.5465
R1019 OUTo.n203 OUTo.n202 0.5465
R1020 OUTo.n195 OUTo.t154 0.5465
R1021 OUTo.n195 OUTo.n194 0.5465
R1022 OUTo.n292 OUTo.t147 0.5465
R1023 OUTo.n292 OUTo.n291 0.5465
R1024 OUTo.n282 OUTo.t174 0.5465
R1025 OUTo.n282 OUTo.n281 0.5465
R1026 OUTo.n326 OUTo.t158 0.5465
R1027 OUTo.n326 OUTo.n325 0.5465
R1028 OUTo.n228 OUTo.t165 0.5465
R1029 OUTo.n228 OUTo.n227 0.5465
R1030 OUTo.n315 OUTo.t182 0.5465
R1031 OUTo.n315 OUTo.n314 0.5465
R1032 OUTo.n395 OUTo.t143 0.5465
R1033 OUTo.n395 OUTo.n394 0.5465
R1034 OUTo.n386 OUTo.t183 0.5465
R1035 OUTo.n386 OUTo.n385 0.5465
R1036 OUTo.n357 OUTo.t131 0.5465
R1037 OUTo.n357 OUTo.n356 0.5465
R1038 OUTo.n362 OUTo.t162 0.5465
R1039 OUTo.n362 OUTo.n361 0.5465
R1040 OUTo.n454 OUTo.t146 0.5465
R1041 OUTo.n454 OUTo.n453 0.5465
R1042 OUTo.n338 OUTo.t167 0.5465
R1043 OUTo.n338 OUTo.n337 0.5465
R1044 OUTo.n399 OUTo.t152 0.5465
R1045 OUTo.n399 OUTo.n398 0.5465
R1046 OUTo.n435 OUTo.t134 0.5465
R1047 OUTo.n435 OUTo.n434 0.5465
R1048 OUTo.n350 OUTo.t130 0.5465
R1049 OUTo.n350 OUTo.n349 0.5465
R1050 OUTo.n342 OUTo.t177 0.5465
R1051 OUTo.n342 OUTo.n341 0.5465
R1052 OUTo.n439 OUTo.t160 0.5465
R1053 OUTo.n439 OUTo.n438 0.5465
R1054 OUTo.n429 OUTo.t170 0.5465
R1055 OUTo.n429 OUTo.n428 0.5465
R1056 OUTo.n473 OUTo.t173 0.5465
R1057 OUTo.n473 OUTo.n472 0.5465
R1058 OUTo.n375 OUTo.t125 0.5465
R1059 OUTo.n375 OUTo.n374 0.5465
R1060 OUTo.n462 OUTo.t140 0.5465
R1061 OUTo.n462 OUTo.n461 0.5465
R1062 OUTo.n486 OUTo.n485 0.449699
R1063 OUTo.n164 OUTo.n161 0.435052
R1064 OUTo.n657 OUTo.n654 0.435052
R1065 OUTo.n506 OUTo.n503 0.435052
R1066 OUTo.n751 OUTo.n748 0.424978
R1067 OUTo.n599 OUTo.n596 0.424978
R1068 OUTo.n789 OUTo.n786 0.424978
R1069 OUTo.n102 OUTo.n99 0.424978
R1070 OUTo.n65 OUTo.n62 0.424978
R1071 OUTo.n637 OUTo.n634 0.424978
R1072 OUTo.n680 OUTo.n642 0.421386
R1073 OUTo.n552 OUTo.n549 0.419604
R1074 OUTo.n561 OUTo.n558 0.419604
R1075 OUTo.n136 OUTo.n133 0.419604
R1076 OUTo.n145 OUTo.n142 0.419604
R1077 OUTo.n704 OUTo.n701 0.419604
R1078 OUTo.n713 OUTo.n710 0.419604
R1079 OUTo.n733 OUTo.n730 0.416918
R1080 OUTo.n581 OUTo.n578 0.416918
R1081 OUTo.n47 OUTo.n44 0.416918
R1082 OUTo.n543 OUTo.n540 0.412216
R1083 OUTo.n127 OUTo.n124 0.412216
R1084 OUTo.n173 OUTo.n170 0.412216
R1085 OUTo.n666 OUTo.n663 0.412216
R1086 OUTo.n695 OUTo.n692 0.412216
R1087 OUTo.n515 OUTo.n512 0.412216
R1088 OUTo.n483 OUTo.n482 0.411509
R1089 OUTo.n742 OUTo.n739 0.40953
R1090 OUTo.n590 OUTo.n587 0.40953
R1091 OUTo.n771 OUTo.n768 0.40953
R1092 OUTo.n84 OUTo.n81 0.40953
R1093 OUTo.n56 OUTo.n53 0.40953
R1094 OUTo.n619 OUTo.n616 0.40953
R1095 OUTo.n780 OUTo.n777 0.408858
R1096 OUTo.n93 OUTo.n90 0.408858
R1097 OUTo.n628 OUTo.n625 0.408858
R1098 OUTo.n182 OUTo.n179 0.404828
R1099 OUTo.n675 OUTo.n672 0.404828
R1100 OUTo.n524 OUTo.n521 0.404828
R1101 OUTo.n795 OUTo.n794 0.404501
R1102 OUTo.n484 OUTo.n286 0.401659
R1103 OUTo.n481 OUTo.n433 0.401659
R1104 OUTo.n485 OUTo.n243 0.40111
R1105 OUTo.n483 OUTo.n333 0.40111
R1106 OUTo.n482 OUTo.n390 0.40111
R1107 OUTo.n163 OUTo.n162 0.197963
R1108 OUTo.n656 OUTo.n655 0.197963
R1109 OUTo.n484 OUTo.n483 0.195723
R1110 OUTo.n485 OUTo.n484 0.195455
R1111 OUTo.n482 OUTo.n481 0.195455
R1112 OUTo.n761 OUTo.n760 0.191535
R1113 OUTo.n74 OUTo.n73 0.191535
R1114 OUTo.n172 OUTo.n171 0.191535
R1115 OUTo.n609 OUTo.n608 0.191535
R1116 OUTo.n665 OUTo.n664 0.191535
R1117 OUTo.n770 OUTo.n769 0.181892
R1118 OUTo.n788 OUTo.n787 0.181892
R1119 OUTo.n83 OUTo.n82 0.181892
R1120 OUTo.n101 OUTo.n100 0.181892
R1121 OUTo.n618 OUTo.n617 0.181892
R1122 OUTo.n636 OUTo.n635 0.181892
R1123 OUTo.n750 OUTo.n749 0.180285
R1124 OUTo.n598 OUTo.n597 0.180285
R1125 OUTo.n64 OUTo.n63 0.180285
R1126 OUTo.n502 OUTo.n501 0.179788
R1127 OUTo.n723 OUTo.n722 0.178677
R1128 OUTo.n732 OUTo.n731 0.178677
R1129 OUTo.n571 OUTo.n570 0.178677
R1130 OUTo.n580 OUTo.n579 0.178677
R1131 OUTo.n560 OUTo.n559 0.178677
R1132 OUTo.n37 OUTo.n36 0.178677
R1133 OUTo.n46 OUTo.n45 0.178677
R1134 OUTo.n144 OUTo.n143 0.178677
R1135 OUTo.n712 OUTo.n711 0.178677
R1136 OUTo.n533 OUTo.n532 0.17707
R1137 OUTo.n117 OUTo.n116 0.17707
R1138 OUTo.n181 OUTo.n180 0.17707
R1139 OUTo.n674 OUTo.n673 0.17707
R1140 OUTo.n685 OUTo.n684 0.17707
R1141 OUTo.n551 OUTo.n550 0.175463
R1142 OUTo.n135 OUTo.n134 0.175463
R1143 OUTo.n154 OUTo.n153 0.175463
R1144 OUTo.n647 OUTo.n646 0.175463
R1145 OUTo.n703 OUTo.n702 0.175463
R1146 OUTo.n604 OUTo.n566 0.174925
R1147 OUTo.n756 OUTo.n718 0.174904
R1148 OUTo.n218 OUTo.n217 0.173016
R1149 OUTo.n198 OUTo.n197 0.173016
R1150 OUTo.n365 OUTo.n364 0.173016
R1151 OUTo.n345 OUTo.n344 0.173016
R1152 OUTo.n542 OUTo.n541 0.172249
R1153 OUTo.n779 OUTo.n778 0.172249
R1154 OUTo.n92 OUTo.n91 0.172249
R1155 OUTo.n126 OUTo.n125 0.172249
R1156 OUTo.n627 OUTo.n626 0.172249
R1157 OUTo.n694 OUTo.n693 0.172249
R1158 OUTo.n250 OUTo.n246 0.171541
R1159 OUTo.n397 OUTo.n393 0.171541
R1160 OUTo.n741 OUTo.n740 0.170642
R1161 OUTo.n589 OUTo.n588 0.170642
R1162 OUTo.n55 OUTo.n54 0.170642
R1163 OUTo.n320 OUTo.n319 0.165639
R1164 OUTo.n467 OUTo.n466 0.165639
R1165 OUTo.n520 OUTo.n519 0.163716
R1166 OUTo.n256 OUTo.n255 0.160498
R1167 OUTo.n403 OUTo.n402 0.160498
R1168 OUTo.n511 OUTo.n510 0.157288
R1169 OUTo.n236 OUTo.n235 0.156072
R1170 OUTo.n383 OUTo.n382 0.156072
R1171 OUTo.n258 OUTo.n257 0.156069
R1172 OUTo.n405 OUTo.n404 0.156069
R1173 OUTo.n323 OUTo.n322 0.146476
R1174 OUTo.n470 OUTo.n469 0.146476
R1175 OUTo.n264 OUTo.n263 0.145927
R1176 OUTo.n270 OUTo.n269 0.145927
R1177 OUTo.n277 OUTo.n276 0.145927
R1178 OUTo.n208 OUTo.n207 0.145927
R1179 OUTo.n223 OUTo.n222 0.145927
R1180 OUTo.n233 OUTo.n232 0.145927
R1181 OUTo.n301 OUTo.n300 0.145927
R1182 OUTo.n411 OUTo.n410 0.145927
R1183 OUTo.n417 OUTo.n416 0.145927
R1184 OUTo.n424 OUTo.n423 0.145927
R1185 OUTo.n355 OUTo.n354 0.145927
R1186 OUTo.n370 OUTo.n369 0.145927
R1187 OUTo.n380 OUTo.n379 0.145927
R1188 OUTo.n448 OUTo.n447 0.145927
R1189 OUTo.n312 OUTo.n311 0.145378
R1190 OUTo.n459 OUTo.n458 0.145378
R1191 OUTo.n9 OUTo.n7 0.0943502
R1192 OUTo.n718 OUTo.n680 0.0918478
R1193 OUTo.n642 OUTo.n604 0.0913143
R1194 OUTo.n794 OUTo.n756 0.0913143
R1195 OUTo.n505 OUTo.n504 0.090779
R1196 OUTo.n514 OUTo.n513 0.0879126
R1197 OUTo.n747 OUTo.n746 0.0848204
R1198 OUTo.n595 OUTo.n594 0.0848204
R1199 OUTo.n61 OUTo.n60 0.0848204
R1200 OUTo.n548 OUTo.n547 0.0841023
R1201 OUTo.n785 OUTo.n784 0.0841023
R1202 OUTo.n98 OUTo.n97 0.0841023
R1203 OUTo.n132 OUTo.n131 0.0841023
R1204 OUTo.n633 OUTo.n632 0.0841023
R1205 OUTo.n700 OUTo.n699 0.0841023
R1206 OUTo.n557 OUTo.n556 0.0826652
R1207 OUTo.n141 OUTo.n140 0.0826652
R1208 OUTo.n160 OUTo.n159 0.0826652
R1209 OUTo.n653 OUTo.n652 0.0826652
R1210 OUTo.n709 OUTo.n708 0.0826652
R1211 OUTo.n169 OUTo.n167 0.082645
R1212 OUTo.n662 OUTo.n660 0.082645
R1213 OUTo.n539 OUTo.n538 0.0819463
R1214 OUTo.n123 OUTo.n122 0.0819463
R1215 OUTo.n691 OUTo.n690 0.0819463
R1216 OUTo.n523 OUTo.n522 0.0814496
R1217 OUTo.n729 OUTo.n728 0.0812272
R1218 OUTo.n738 OUTo.n737 0.0812272
R1219 OUTo.n577 OUTo.n576 0.0812272
R1220 OUTo.n586 OUTo.n585 0.0812272
R1221 OUTo.n43 OUTo.n42 0.0812272
R1222 OUTo.n52 OUTo.n51 0.0812272
R1223 OUTo.n496 OUTo.n495 0.0807304
R1224 OUTo.n178 OUTo.n176 0.0805961
R1225 OUTo.n671 OUTo.n669 0.0805961
R1226 OUTo.n767 OUTo.n765 0.080303
R1227 OUTo.n80 OUTo.n78 0.080303
R1228 OUTo.n615 OUTo.n613 0.080303
R1229 OUTo.n776 OUTo.n775 0.0797883
R1230 OUTo.n89 OUTo.n88 0.0797883
R1231 OUTo.n624 OUTo.n623 0.0797883
R1232 OUTo.n730 OUTo.n724 0.0784104
R1233 OUTo.n739 OUTo.n733 0.0784104
R1234 OUTo.n748 OUTo.n742 0.0784104
R1235 OUTo.n755 OUTo.n751 0.0784104
R1236 OUTo.n578 OUTo.n572 0.0784104
R1237 OUTo.n587 OUTo.n581 0.0784104
R1238 OUTo.n596 OUTo.n590 0.0784104
R1239 OUTo.n603 OUTo.n599 0.0784104
R1240 OUTo.n540 OUTo.n534 0.0784104
R1241 OUTo.n549 OUTo.n543 0.0784104
R1242 OUTo.n558 OUTo.n552 0.0784104
R1243 OUTo.n565 OUTo.n561 0.0784104
R1244 OUTo.n768 OUTo.n762 0.0784104
R1245 OUTo.n777 OUTo.n771 0.0784104
R1246 OUTo.n786 OUTo.n780 0.0784104
R1247 OUTo.n793 OUTo.n789 0.0784104
R1248 OUTo.n81 OUTo.n75 0.0784104
R1249 OUTo.n90 OUTo.n84 0.0784104
R1250 OUTo.n99 OUTo.n93 0.0784104
R1251 OUTo.n106 OUTo.n102 0.0784104
R1252 OUTo.n44 OUTo.n38 0.0784104
R1253 OUTo.n53 OUTo.n47 0.0784104
R1254 OUTo.n62 OUTo.n56 0.0784104
R1255 OUTo.n69 OUTo.n65 0.0784104
R1256 OUTo.n124 OUTo.n118 0.0784104
R1257 OUTo.n133 OUTo.n127 0.0784104
R1258 OUTo.n142 OUTo.n136 0.0784104
R1259 OUTo.n149 OUTo.n145 0.0784104
R1260 OUTo.n161 OUTo.n155 0.0784104
R1261 OUTo.n170 OUTo.n164 0.0784104
R1262 OUTo.n179 OUTo.n173 0.0784104
R1263 OUTo.n186 OUTo.n182 0.0784104
R1264 OUTo.n616 OUTo.n610 0.0784104
R1265 OUTo.n625 OUTo.n619 0.0784104
R1266 OUTo.n634 OUTo.n628 0.0784104
R1267 OUTo.n641 OUTo.n637 0.0784104
R1268 OUTo.n654 OUTo.n648 0.0784104
R1269 OUTo.n663 OUTo.n657 0.0784104
R1270 OUTo.n672 OUTo.n666 0.0784104
R1271 OUTo.n679 OUTo.n675 0.0784104
R1272 OUTo.n692 OUTo.n686 0.0784104
R1273 OUTo.n701 OUTo.n695 0.0784104
R1274 OUTo.n710 OUTo.n704 0.0784104
R1275 OUTo.n717 OUTo.n713 0.0784104
R1276 OUTo.n503 OUTo.n497 0.0784104
R1277 OUTo.n512 OUTo.n506 0.0784104
R1278 OUTo.n521 OUTo.n515 0.0784104
R1279 OUTo.n528 OUTo.n524 0.0784104
R1280 OUTo.n776 OUTo.n774 0.0770706
R1281 OUTo.n89 OUTo.n87 0.0770706
R1282 OUTo.n624 OUTo.n622 0.0770706
R1283 OUTo.n729 OUTo.n727 0.0758918
R1284 OUTo.n738 OUTo.n736 0.0758918
R1285 OUTo.n577 OUTo.n575 0.0758918
R1286 OUTo.n586 OUTo.n584 0.0758918
R1287 OUTo.n43 OUTo.n41 0.0758918
R1288 OUTo.n52 OUTo.n50 0.0758918
R1289 OUTo.n767 OUTo.n766 0.0754658
R1290 OUTo.n80 OUTo.n79 0.0754658
R1291 OUTo.n178 OUTo.n177 0.0754658
R1292 OUTo.n615 OUTo.n614 0.0754658
R1293 OUTo.n671 OUTo.n670 0.0754658
R1294 OUTo.n539 OUTo.n537 0.0753017
R1295 OUTo.n123 OUTo.n121 0.0753017
R1296 OUTo.n691 OUTo.n689 0.0753017
R1297 OUTo.n557 OUTo.n555 0.0744132
R1298 OUTo.n141 OUTo.n139 0.0744132
R1299 OUTo.n709 OUTo.n707 0.0744132
R1300 OUTo.n160 OUTo.n158 0.0743729
R1301 OUTo.n653 OUTo.n651 0.0743729
R1302 OUTo.n785 OUTo.n783 0.0735187
R1303 OUTo.n98 OUTo.n96 0.0735187
R1304 OUTo.n633 OUTo.n631 0.0735187
R1305 OUTo.n548 OUTo.n546 0.0732202
R1306 OUTo.n132 OUTo.n130 0.0732202
R1307 OUTo.n700 OUTo.n698 0.0732202
R1308 OUTo OUTo.n112 0.0730539
R1309 OUTo.n747 OUTo.n745 0.0726227
R1310 OUTo.n595 OUTo.n593 0.0726227
R1311 OUTo.n61 OUTo.n59 0.0726227
R1312 OUTo.n169 OUTo.n168 0.0725795
R1313 OUTo.n662 OUTo.n661 0.0725795
R1314 OUTo.n284 OUTo.n283 0.0705602
R1315 OUTo.n431 OUTo.n430 0.0705602
R1316 OUTo.n298 OUTo.n297 0.0693681
R1317 OUTo.n445 OUTo.n444 0.0693681
R1318 OUTo.n304 OUTo.n303 0.0687718
R1319 OUTo.n331 OUTo.n330 0.0687718
R1320 OUTo.n451 OUTo.n450 0.0687718
R1321 OUTo.n478 OUTo.n477 0.0687718
R1322 OUTo OUTo.n798 0.0686231
R1323 OUTo.n245 OUTo.n244 0.0678863
R1324 OUTo.n392 OUTo.n391 0.0678863
R1325 OUTo.n273 OUTo.n272 0.0672896
R1326 OUTo.n420 OUTo.n419 0.0672896
R1327 OUTo.n22 OUTo.n21 0.0671964
R1328 OUTo.n220 OUTo.n219 0.0649012
R1329 OUTo.n188 OUTo.n187 0.0649012
R1330 OUTo.n367 OUTo.n366 0.0649012
R1331 OUTo.n335 OUTo.n334 0.0649012
R1332 OUTo.n200 OUTo.n199 0.0643037
R1333 OUTo.n347 OUTo.n346 0.0643037
R1334 OUTo.n797 OUTo.n796 0.0581
R1335 OUTo.n32 OUTo.n31 0.0575462
R1336 OUTo.n489 OUTo.n488 0.056049
R1337 OUTo.n109 OUTo.n108 0.0555148
R1338 OUTo.n217 OUTo.n216 0.0538329
R1339 OUTo.n254 OUTo.n253 0.0538329
R1340 OUTo.n197 OUTo.n196 0.0538329
R1341 OUTo.n364 OUTo.n363 0.0538329
R1342 OUTo.n401 OUTo.n400 0.0538329
R1343 OUTo.n344 OUTo.n343 0.0538329
R1344 OUTo.n284 OUTo.n280 0.0534224
R1345 OUTo.n431 OUTo.n427 0.0534224
R1346 OUTo.n317 OUTo.n316 0.045622
R1347 OUTo.n464 OUTo.n463 0.045622
R1348 OUTo.n241 OUTo.n240 0.0445215
R1349 OUTo.n388 OUTo.n387 0.0445215
R1350 OUTo.n511 OUTo.n509 0.043333
R1351 OUTo.n520 OUTo.n518 0.0413095
R1352 OUTo.n19 OUTo.n18 0.0406142
R1353 OUTo.n16 OUTo.n12 0.0392692
R1354 OUTo.n502 OUTo.n500 0.0348512
R1355 OUTo.n31 OUTo.n30 0.0337308
R1356 OUTo.n112 OUTo.n32 0.0337308
R1357 OUTo.n798 OUTo.n797 0.0337308
R1358 OUTo.n796 OUTo.n795 0.0337308
R1359 OUTo.n250 OUTo.n249 0.0317394
R1360 OUTo.n397 OUTo.n396 0.0317394
R1361 OUTo.n6 OUTo.n5 0.028625
R1362 OUTo.n15 OUTo.n14 0.028625
R1363 OUTo.n29 OUTo.n16 0.0268077
R1364 OUTo.n21 OUTo.n20 0.0262143
R1365 OUTo.n27 OUTo.n26 0.0262143
R1366 OUTo.n294 OUTo.n293 0.0253785
R1367 OUTo.n441 OUTo.n440 0.0253785
R1368 OUTo.n309 OUTo.n308 0.0251875
R1369 OUTo.n328 OUTo.n327 0.0251875
R1370 OUTo.n456 OUTo.n455 0.0251875
R1371 OUTo.n475 OUTo.n474 0.0251875
R1372 OUTo.n23 OUTo.n22 0.0247138
R1373 OUTo.n10 OUTo.n4 0.0242491
R1374 OUTo.n212 OUTo.n211 0.0229088
R1375 OUTo.n230 OUTo.n229 0.0229088
R1376 OUTo.n359 OUTo.n358 0.0229088
R1377 OUTo.n377 OUTo.n376 0.0229088
R1378 OUTo.n205 OUTo.n204 0.0222846
R1379 OUTo.n352 OUTo.n351 0.0222846
R1380 OUTo.n24 OUTo.n17 0.0205893
R1381 OUTo.n111 OUTo.n110 0.0181261
R1382 OUTo.n491 OUTo.n490 0.017592
R1383 OUTo.n487 OUTo.n486 0.0173249
R1384 OUTo.n108 OUTo.n107 0.0167908
R1385 OUTo.n10 OUTo.n9 0.0159927
R1386 OUTo.n488 OUTo.n487 0.0157226
R1387 OUTo.n490 OUTo.n489 0.0154555
R1388 OUTo.n110 OUTo.n109 0.0149214
R1389 OUTo.n29 OUTo.n28 0.0129615
R1390 OUTo.n221 OUTo.n213 0.0118709
R1391 OUTo.n206 OUTo.n201 0.0118709
R1392 OUTo.n310 OUTo.n305 0.0118709
R1393 OUTo.n299 OUTo.n295 0.0118709
R1394 OUTo.n368 OUTo.n360 0.0118709
R1395 OUTo.n353 OUTo.n348 0.0118709
R1396 OUTo.n457 OUTo.n452 0.0118709
R1397 OUTo.n446 OUTo.n442 0.0118709
R1398 OUTo.n213 OUTo.n208 0.0115229
R1399 OUTo.n201 OUTo.n193 0.0115229
R1400 OUTo.n295 OUTo.n290 0.0115229
R1401 OUTo.n305 OUTo.n301 0.0115229
R1402 OUTo.n360 OUTo.n355 0.0115229
R1403 OUTo.n348 OUTo.n340 0.0115229
R1404 OUTo.n442 OUTo.n437 0.0115229
R1405 OUTo.n452 OUTo.n448 0.0115229
R1406 OUTo.n222 OUTo.n221 0.0112206
R1407 OUTo.n207 OUTo.n206 0.0112206
R1408 OUTo.n300 OUTo.n299 0.0112206
R1409 OUTo.n311 OUTo.n310 0.0112206
R1410 OUTo.n369 OUTo.n368 0.0112206
R1411 OUTo.n354 OUTo.n353 0.0112206
R1412 OUTo.n447 OUTo.n446 0.0112206
R1413 OUTo.n458 OUTo.n457 0.0112206
R1414 OUTo.n1 OUTo.n0 0.0107848
R1415 OUTo.n274 OUTo.n271 0.00917073
R1416 OUTo.n279 OUTo.n278 0.00917073
R1417 OUTo.n285 OUTo.n279 0.00917073
R1418 OUTo.n275 OUTo.n274 0.00917073
R1419 OUTo.n329 OUTo.n324 0.00917073
R1420 OUTo.n332 OUTo.n329 0.00917073
R1421 OUTo.n421 OUTo.n418 0.00917073
R1422 OUTo.n426 OUTo.n425 0.00917073
R1423 OUTo.n432 OUTo.n426 0.00917073
R1424 OUTo.n422 OUTo.n421 0.00917073
R1425 OUTo.n476 OUTo.n471 0.00917073
R1426 OUTo.n479 OUTo.n476 0.00917073
R1427 OUTo.n262 OUTo.n260 0.00917073
R1428 OUTo.n267 OUTo.n265 0.00917073
R1429 OUTo.n268 OUTo.n267 0.00917073
R1430 OUTo.n260 OUTo.n259 0.00917073
R1431 OUTo.n237 OUTo.n234 0.00917073
R1432 OUTo.n242 OUTo.n237 0.00917073
R1433 OUTo.n318 OUTo.n313 0.00917073
R1434 OUTo.n321 OUTo.n318 0.00917073
R1435 OUTo.n409 OUTo.n407 0.00917073
R1436 OUTo.n414 OUTo.n412 0.00917073
R1437 OUTo.n415 OUTo.n414 0.00917073
R1438 OUTo.n407 OUTo.n406 0.00917073
R1439 OUTo.n384 OUTo.n381 0.00917073
R1440 OUTo.n389 OUTo.n384 0.00917073
R1441 OUTo.n465 OUTo.n460 0.00917073
R1442 OUTo.n468 OUTo.n465 0.00917073
R1443 OUTo.n286 OUTo.n285 0.00839636
R1444 OUTo.n278 OUTo.n277 0.00839636
R1445 OUTo.n225 OUTo.n224 0.00839636
R1446 OUTo.n224 OUTo.n223 0.00839636
R1447 OUTo.n271 OUTo.n270 0.00839636
R1448 OUTo.n276 OUTo.n275 0.00839636
R1449 OUTo.n333 OUTo.n332 0.00839636
R1450 OUTo.n324 OUTo.n323 0.00839636
R1451 OUTo.n433 OUTo.n432 0.00839636
R1452 OUTo.n425 OUTo.n424 0.00839636
R1453 OUTo.n372 OUTo.n371 0.00839636
R1454 OUTo.n371 OUTo.n370 0.00839636
R1455 OUTo.n418 OUTo.n417 0.00839636
R1456 OUTo.n423 OUTo.n422 0.00839636
R1457 OUTo.n480 OUTo.n479 0.00839636
R1458 OUTo.n471 OUTo.n470 0.00839636
R1459 OUTo.n259 OUTo.n258 0.00839636
R1460 OUTo.n269 OUTo.n268 0.00839636
R1461 OUTo.n263 OUTo.n262 0.00839636
R1462 OUTo.n265 OUTo.n264 0.00839636
R1463 OUTo.n232 OUTo.n231 0.00839636
R1464 OUTo.n234 OUTo.n233 0.00839636
R1465 OUTo.n243 OUTo.n242 0.00839636
R1466 OUTo.n231 OUTo.n226 0.00839636
R1467 OUTo.n322 OUTo.n321 0.00839636
R1468 OUTo.n313 OUTo.n312 0.00839636
R1469 OUTo.n406 OUTo.n405 0.00839636
R1470 OUTo.n416 OUTo.n415 0.00839636
R1471 OUTo.n410 OUTo.n409 0.00839636
R1472 OUTo.n412 OUTo.n411 0.00839636
R1473 OUTo.n379 OUTo.n378 0.00839636
R1474 OUTo.n381 OUTo.n380 0.00839636
R1475 OUTo.n390 OUTo.n389 0.00839636
R1476 OUTo.n378 OUTo.n373 0.00839636
R1477 OUTo.n469 OUTo.n468 0.00839636
R1478 OUTo.n460 OUTo.n459 0.00839636
R1479 OUTo.n20 OUTo.n19 0.00692857
R1480 OUTo.n27 OUTo.n25 0.00692857
R1481 OUTo.n7 OUTo.n6 0.00451786
R1482 OUTo.n15 OUTo.n13 0.00451786
R1483 OUTo.n3 OUTo.n2 0.00210714
R1484 OUTo.n226 OUTo.n225 0.00104878
R1485 OUTo.n373 OUTo.n372 0.00104878
R1486 VDD.t307 VDD.t447 128.756
R1487 VDD.t265 VDD.t321 128.756
R1488 VDD.n532 VDD.t459 112.593
R1489 VDD.n467 VDD.t444 112.593
R1490 VDD.n418 VDD.t307 64.3782
R1491 VDD.n418 VDD.t265 64.3782
R1492 VDD.n638 VDD.t377 45.7877
R1493 VDD.n725 VDD.t332 45.7877
R1494 VDD.n1137 VDD.t398 45.7877
R1495 VDD.n1932 VDD.t412 45.7877
R1496 VDD.n1217 VDD.t344 45.7877
R1497 VDD.n375 VDD.t396 45.7559
R1498 VDD.n388 VDD.t408 45.7559
R1499 VDD.n311 VDD.t373 45.7559
R1500 VDD.n319 VDD.t349 45.7559
R1501 VDD.n251 VDD.t416 45.7559
R1502 VDD.n261 VDD.t389 45.7559
R1503 VDD.n187 VDD.t394 45.7559
R1504 VDD.n195 VDD.t357 45.7559
R1505 VDD.n62 VDD.t410 45.7559
R1506 VDD.n70 VDD.t379 45.7559
R1507 VDD.n126 VDD.t338 45.7559
R1508 VDD.n136 VDD.t414 45.7559
R1509 VDD.n388 VDD.t385 45.6574
R1510 VDD.n319 VDD.t406 45.6574
R1511 VDD.n261 VDD.t402 45.6574
R1512 VDD.n195 VDD.t383 45.6574
R1513 VDD.n70 VDD.t365 45.6574
R1514 VDD.n136 VDD.t381 45.6574
R1515 VDD.n429 VDD.t362 45.6255
R1516 VDD.n382 VDD.t400 45.6255
R1517 VDD.n638 VDD.t355 45.6255
R1518 VDD.n725 VDD.t387 45.6255
R1519 VDD.n1137 VDD.t360 45.6255
R1520 VDD.n1932 VDD.t368 45.6255
R1521 VDD.n1217 VDD.t404 45.6255
R1522 VDD.n1317 VDD.t353 25.8626
R1523 VDD.n1613 VDD.t346 23.622
R1524 VDD.n1844 VDD.t370 23.622
R1525 VDD.n1853 VDD.t341 23.0774
R1526 VDD.n1702 VDD.t391 23.0774
R1527 VDD.n1796 VDD.t311 22.3774
R1528 VDD.n1043 VDD.t336 21.2649
R1529 VDD.n1683 VDD.t289 19.3637
R1530 VDD.n1825 VDD.t456 17.4048
R1531 VDD.n1837 VDD.t269 15.4157
R1532 VDD.n964 VDD.t284 13.2189
R1533 VDD.n2329 VDD.t272 12.698
R1534 VDD.n990 VDD.t8 12.0695
R1535 VDD.n2690 VDD.t443 11.6184
R1536 VDD.n2484 VDD.t7 11.4588
R1537 VDD.n1830 VDD.t308 11.4376
R1538 VDD.n1586 VDD.t366 11.2284
R1539 VDD.n610 VDD.t350 11.2284
R1540 VDD.n954 VDD.t358 11.2284
R1541 VDD.n2310 VDD.t0 11.005
R1542 VDD.n1527 VDD.t108 10.7506
R1543 VDD.n551 VDD.t84 10.7506
R1544 VDD.n895 VDD.t70 10.7506
R1545 VDD.n1815 VDD.t286 10.4431
R1546 VDD.n2455 VDD.t429 10.4172
R1547 VDD.n1039 VDD.t375 9.9285
R1548 VDD.n2711 VDD.t299 9.89723
R1549 VDD.n1325 VDD.t418 9.8555
R1550 VDD.n1325 VDD.t352 9.7095
R1551 VDD.n1039 VDD.t335 9.6365
R1552 VDD.n3121 VDD.t293 9.61159
R1553 VDD.n1792 VDD.t392 9.44854
R1554 VDD.n1546 VDD.t87 9.31727
R1555 VDD.n570 VDD.t82 9.31727
R1556 VDD.n914 VDD.t45 9.31727
R1557 VDD.n2177 VDD.t282 9.16456
R1558 VDD.n1680 VDD.t420 9.03664
R1559 VDD.n2498 VDD.t434 8.85467
R1560 VDD.n1566 VDD.t21 8.83949
R1561 VDD.n590 VDD.t43 8.83949
R1562 VDD.n934 VDD.t34 8.83949
R1563 VDD.n1053 VDD.t277 8.62119
R1564 VDD.n1802 VDD.t3 8.45401
R1565 VDD.n2493 VDD.t438 8.33383
R1566 VDD.n2186 VDD.t1 7.15294
R1567 VDD.n421 VDD.t445 7.11063
R1568 VDD.n534 VDD.t460 7.09044
R1569 VDD.n531 VDD.t461 7.01175
R1570 VDD.n424 VDD.t446 7.01175
R1571 VDD.n1563 VDD.t10 6.92836
R1572 VDD.n587 VDD.t65 6.92836
R1573 VDD.n931 VDD.t55 6.92836
R1574 VDD.n2463 VDD.t300 6.77133
R1575 VDD.n2210 VDD.t283 6.70591
R1576 VDD.n1550 VDD.t12 6.45057
R1577 VDD.n574 VDD.t23 6.45057
R1578 VDD.n918 VDD.t52 6.45057
R1579 VDD.n2345 VDD.t314 5.92601
R1580 VDD.n2486 VDD.t437 5.72967
R1581 VDD.n1790 VDD.t347 5.47042
R1582 VDD.n1523 VDD.t339 5.01722
R1583 VDD.n547 VDD.t363 5.01722
R1584 VDD.n891 VDD.t333 5.01722
R1585 VDD.n2323 VDD.t326 4.79734
R1586 VDD.n1579 VDD.t68 4.53944
R1587 VDD.n603 VDD.t76 4.53944
R1588 VDD.n947 VDD.t26 4.53944
R1589 VDD.n1799 VDD.t422 4.47589
R1590 VDD.n2469 VDD.t298 4.16717
R1591 VDD.n1533 VDD.t39 4.06166
R1592 VDD.n557 VDD.t29 4.06166
R1593 VDD.n901 VDD.t48 4.06166
R1594 VDD.n1022 VDD.t275 4.02349
R1595 VDD.n389 VDD.n388 4.0005
R1596 VDD.n376 VDD.n375 4.0005
R1597 VDD.n383 VDD.n382 4.0005
R1598 VDD.n430 VDD.n429 4.0005
R1599 VDD.n320 VDD.n319 4.0005
R1600 VDD.n312 VDD.n311 4.0005
R1601 VDD.n314 VDD.n313 4.0005
R1602 VDD.n639 VDD.n638 4.0005
R1603 VDD.n262 VDD.n261 4.0005
R1604 VDD.n252 VDD.n251 4.0005
R1605 VDD.n256 VDD.n255 4.0005
R1606 VDD.n726 VDD.n725 4.0005
R1607 VDD.n196 VDD.n195 4.0005
R1608 VDD.n188 VDD.n187 4.0005
R1609 VDD.n190 VDD.n189 4.0005
R1610 VDD.n1138 VDD.n1137 4.0005
R1611 VDD.n71 VDD.n70 4.0005
R1612 VDD.n63 VDD.n62 4.0005
R1613 VDD.n65 VDD.n64 4.0005
R1614 VDD.n1933 VDD.n1932 4.0005
R1615 VDD.n137 VDD.n136 4.0005
R1616 VDD.n127 VDD.n126 4.0005
R1617 VDD.n131 VDD.n130 4.0005
R1618 VDD.n1218 VDD.n1217 4.0005
R1619 VDD.n1853 VDD.t343 3.92171
R1620 VDD.n1702 VDD.t393 3.92171
R1621 VDD.n2449 VDD.n2448 3.54139
R1622 VDD.n981 VDD.t276 3.5105
R1623 VDD.n982 VDD.t449 3.5105
R1624 VDD.n526 VDD.n524 3.48636
R1625 VDD.n1387 VDD.n1385 3.48636
R1626 VDD.n1461 VDD.n1459 3.48636
R1627 VDD.n2754 VDD.n2753 3.48583
R1628 VDD.n2754 VDD.n2751 3.48583
R1629 VDD.n2908 VDD.n2906 3.48583
R1630 VDD.n850 VDD.n849 3.48583
R1631 VDD.n809 VDD.n807 3.48583
R1632 VDD.n809 VDD.n808 3.48583
R1633 VDD.n792 VDD.n791 3.48583
R1634 VDD.n771 VDD.n769 3.48583
R1635 VDD.n792 VDD.n790 3.48583
R1636 VDD.n828 VDD.n826 3.48583
R1637 VDD.n850 VDD.n848 3.48583
R1638 VDD.n471 VDD.n469 3.48583
R1639 VDD.n459 VDD.n457 3.48583
R1640 VDD.n459 VDD.n458 3.48583
R1641 VDD.n510 VDD.n508 3.48583
R1642 VDD.n510 VDD.n509 3.48583
R1643 VDD.n526 VDD.n525 3.48583
R1644 VDD.n292 VDD.n290 3.48583
R1645 VDD.n1387 VDD.n1386 3.48583
R1646 VDD.n1404 VDD.n1403 3.48583
R1647 VDD.n1404 VDD.n1402 3.48583
R1648 VDD.n1425 VDD.n1424 3.48583
R1649 VDD.n1425 VDD.n1423 3.48583
R1650 VDD.n1442 VDD.n1441 3.48583
R1651 VDD.n1461 VDD.n1460 3.48583
R1652 VDD.n1479 VDD.n1478 3.48583
R1653 VDD.n1479 VDD.n1477 3.48583
R1654 VDD.n1499 VDD.n1498 3.48583
R1655 VDD.n1499 VDD.n1497 3.48583
R1656 VDD.n154 VDD.n153 3.48583
R1657 VDD.n1284 VDD.n1282 3.48569
R1658 VDD.n1294 VDD.n1290 3.48569
R1659 VDD.n1294 VDD.n1293 3.48569
R1660 VDD.n2771 VDD.n2770 3.48569
R1661 VDD.n2792 VDD.n2791 3.48569
R1662 VDD.n1673 VDD.n1672 3.48569
R1663 VDD.n1759 VDD.n1758 3.48569
R1664 VDD.n1751 VDD.n1750 3.48569
R1665 VDD.n1743 VDD.n1741 3.48569
R1666 VDD.n1884 VDD.n1881 3.48569
R1667 VDD.n1434 VDD.n1432 3.48569
R1668 VDD.n1415 VDD.n1413 3.48569
R1669 VDD.n1396 VDD.n1394 3.48569
R1670 VDD.n1379 VDD.n1377 3.48569
R1671 VDD.n279 VDD.n278 3.48569
R1672 VDD.n866 VDD.n865 3.48569
R1673 VDD.n626 VDD.n624 3.48569
R1674 VDD.n762 VDD.n760 3.48569
R1675 VDD.n782 VDD.n780 3.48569
R1676 VDD.n801 VDD.n799 3.48569
R1677 VDD.n306 VDD.n301 3.48569
R1678 VDD.n182 VDD.n181 3.48569
R1679 VDD.n168 VDD.n167 3.48569
R1680 VDD.n2062 VDD.n2060 3.48569
R1681 VDD.n2042 VDD.n2040 3.48569
R1682 VDD.n2164 VDD.n2162 3.48569
R1683 VDD.n1602 VDD.n1600 3.48569
R1684 VDD.n479 VDD.n478 3.4853
R1685 VDD.n2792 VDD.n2790 3.48517
R1686 VDD.n2771 VDD.n2769 3.48517
R1687 VDD.n2908 VDD.n2907 3.48517
R1688 VDD.n1623 VDD.n1621 3.48517
R1689 VDD.n1759 VDD.n1757 3.48517
R1690 VDD.n1751 VDD.n1749 3.48517
R1691 VDD.n1743 VDD.n1742 3.48517
R1692 VDD.n1884 VDD.n1883 3.48517
R1693 VDD.n1434 VDD.n1433 3.48517
R1694 VDD.n1415 VDD.n1414 3.48517
R1695 VDD.n1396 VDD.n1395 3.48517
R1696 VDD.n1379 VDD.n1378 3.48517
R1697 VDD.n279 VDD.n277 3.48517
R1698 VDD.n866 VDD.n864 3.48517
R1699 VDD.n306 VDD.n305 3.48517
R1700 VDD.n801 VDD.n800 3.48517
R1701 VDD.n782 VDD.n781 3.48517
R1702 VDD.n762 VDD.n761 3.48517
R1703 VDD.n626 VDD.n625 3.48517
R1704 VDD.n428 VDD.n426 3.48517
R1705 VDD.n182 VDD.n180 3.48517
R1706 VDD.n168 VDD.n166 3.48517
R1707 VDD.n57 VDD.n56 3.48517
R1708 VDD.n2164 VDD.n2163 3.48517
R1709 VDD.n2062 VDD.n2061 3.48517
R1710 VDD.n2042 VDD.n2041 3.48517
R1711 VDD.n1602 VDD.n1601 3.48517
R1712 VDD.n2449 VDD.n2447 3.48517
R1713 VDD.n1616 VDD.n1615 3.48503
R1714 VDD.n1616 VDD.n1614 3.48503
R1715 VDD.n1620 VDD.n1619 3.48503
R1716 VDD.n1620 VDD.n1618 3.48503
R1717 VDD.n1623 VDD.n1622 3.48503
R1718 VDD.n1769 VDD.n1768 3.48503
R1719 VDD.n1769 VDD.n1765 3.48503
R1720 VDD.n1852 VDD.n1850 3.48503
R1721 VDD.n1852 VDD.n1851 3.48503
R1722 VDD.n1506 VDD.n1505 3.48503
R1723 VDD.n1506 VDD.n1504 3.48503
R1724 VDD.n1489 VDD.n1488 3.48503
R1725 VDD.n57 VDD.n55 3.48503
R1726 VDD.n2079 VDD.n2077 3.48503
R1727 VDD.n2079 VDD.n2078 3.48503
R1728 VDD.n1809 VDD.t5 3.48136
R1729 VDD.n1805 VDD.n1795 3.46514
R1730 VDD.n1836 VDD.n1829 3.46514
R1731 VDD.n1921 VDD.n1843 3.46514
R1732 VDD.n1822 VDD.n1821 3.46514
R1733 VDD.n1860 VDD.n1855 3.42447
R1734 VDD.n1714 VDD.n1705 3.42447
R1735 VDD.n1727 VDD.n1703 3.42447
R1736 VDD.n3128 VDD.t322 3.3532
R1737 VDD.n432 VDD.t364 3.20717
R1738 VDD.n641 VDD.t356 3.20717
R1739 VDD.n637 VDD.t378 3.20717
R1740 VDD.n316 VDD.t374 3.20717
R1741 VDD.n318 VDD.t351 3.20717
R1742 VDD.n322 VDD.t407 3.20717
R1743 VDD.n1140 VDD.t361 3.20717
R1744 VDD.n728 VDD.t388 3.20717
R1745 VDD.n724 VDD.t334 3.20717
R1746 VDD.n1136 VDD.t399 3.20717
R1747 VDD.n192 VDD.t395 3.20717
R1748 VDD.n194 VDD.t359 3.20717
R1749 VDD.n198 VDD.t384 3.20717
R1750 VDD.n1935 VDD.t369 3.20717
R1751 VDD.n1931 VDD.t413 3.20717
R1752 VDD.n67 VDD.t411 3.20717
R1753 VDD.n69 VDD.t380 3.20717
R1754 VDD.n73 VDD.t367 3.20717
R1755 VDD.n1220 VDD.t405 3.20717
R1756 VDD.n1216 VDD.t345 3.20717
R1757 VDD.n828 VDD.n827 3.16765
R1758 VDD.n771 VDD.n770 3.16765
R1759 VDD.n471 VDD.n470 3.16765
R1760 VDD.n292 VDD.n291 3.16765
R1761 VDD.n635 VDD.n634 3.16712
R1762 VDD.n507 VDD.n506 3.16696
R1763 VDD.n528 VDD.n527 3.16696
R1764 VDD.n1284 VDD.n1283 3.16682
R1765 VDD.n2900 VDD.n2899 3.16022
R1766 VDD.n533 VDD.n532 3.1505
R1767 VDD.n423 VDD.n422 3.1505
R1768 VDD.n468 VDD.n467 3.1505
R1769 VDD.n1126 VDD.n1125 3.1505
R1770 VDD.n969 VDD.n968 3.1505
R1771 VDD.n1301 VDD.n1300 3.1505
R1772 VDD.n1226 VDD.n1225 3.1505
R1773 VDD.n1225 VDD.n1224 3.1505
R1774 VDD.n1313 VDD.n1312 3.1505
R1775 VDD.n1312 VDD.n1311 3.1505
R1776 VDD.n1316 VDD.n1315 3.1505
R1777 VDD.n1315 VDD.n1314 3.1505
R1778 VDD.n1318 VDD.n1317 3.1505
R1779 VDD.n1320 VDD.n1319 3.1505
R1780 VDD.n1306 VDD.n1305 3.1505
R1781 VDD.n1305 VDD.n1304 3.1505
R1782 VDD.n966 VDD.n965 3.1505
R1783 VDD.n965 VDD.n964 3.1505
R1784 VDD.n968 VDD.n967 3.1505
R1785 VDD.n1010 VDD.n1009 3.1505
R1786 VDD.n1012 VDD.n1011 3.1505
R1787 VDD.n1008 VDD.n1007 3.1505
R1788 VDD.n1007 VDD.n1006 3.1505
R1789 VDD.n998 VDD.n997 3.1505
R1790 VDD.n997 VDD.n996 3.1505
R1791 VDD.n991 VDD.n990 3.1505
R1792 VDD.n993 VDD.n992 3.1505
R1793 VDD.n989 VDD.n988 3.1505
R1794 VDD.n988 VDD.n987 3.1505
R1795 VDD.n986 VDD.n985 3.1505
R1796 VDD.n985 VDD.n984 3.1505
R1797 VDD.n1027 VDD.n1026 3.1505
R1798 VDD.n1026 VDD.n1025 3.1505
R1799 VDD.n1024 VDD.n1023 3.1505
R1800 VDD.n1023 VDD.n1022 3.1505
R1801 VDD.n1021 VDD.n1020 3.1505
R1802 VDD.n1020 VDD.n1019 3.1505
R1803 VDD.n1018 VDD.n1017 3.1505
R1804 VDD.n1017 VDD.n1016 3.1505
R1805 VDD.n1055 VDD.n1054 3.1505
R1806 VDD.n1054 VDD.n1053 3.1505
R1807 VDD.n1052 VDD.n1051 3.1505
R1808 VDD.n1051 VDD.n1050 3.1505
R1809 VDD.n1048 VDD.n1047 3.1505
R1810 VDD.n1047 VDD.n1046 3.1505
R1811 VDD.n1045 VDD.n1044 3.1505
R1812 VDD.n1044 VDD.n1043 3.1505
R1813 VDD.n1067 VDD.n1066 3.1505
R1814 VDD.n1066 VDD.n1065 3.1505
R1815 VDD.n1061 VDD.n1060 3.1505
R1816 VDD.n1063 VDD.n1062 3.1505
R1817 VDD.n1124 VDD.n1123 3.1505
R1818 VDD.n1119 VDD.n1118 3.1505
R1819 VDD.n1117 VDD.n1116 3.1505
R1820 VDD.n1114 VDD.n1113 3.1505
R1821 VDD.n1112 VDD.n1111 3.1505
R1822 VDD.n1109 VDD.n1108 3.1505
R1823 VDD.n1107 VDD.n1106 3.1505
R1824 VDD.n1104 VDD.n1103 3.1505
R1825 VDD.n1102 VDD.n1101 3.1505
R1826 VDD.n1099 VDD.n1098 3.1505
R1827 VDD.n1097 VDD.n1096 3.1505
R1828 VDD.n1094 VDD.n1093 3.1505
R1829 VDD.n1092 VDD.n1091 3.1505
R1830 VDD.n1089 VDD.n1088 3.1505
R1831 VDD.n1087 VDD.n1086 3.1505
R1832 VDD.n1084 VDD.n1083 3.1505
R1833 VDD.n1082 VDD.n1081 3.1505
R1834 VDD.n1080 VDD.n1079 3.1505
R1835 VDD.n1078 VDD.n1077 3.1505
R1836 VDD.n1076 VDD.n1075 3.1505
R1837 VDD.n1074 VDD.n1073 3.1505
R1838 VDD.n1072 VDD.n1071 3.1505
R1839 VDD.n1036 VDD.n1035 3.1505
R1840 VDD.n1034 VDD.n1033 3.1505
R1841 VDD.n971 VDD.n970 3.1505
R1842 VDD.n973 VDD.n972 3.1505
R1843 VDD.n975 VDD.n974 3.1505
R1844 VDD.n977 VDD.n976 3.1505
R1845 VDD.n979 VDD.n978 3.1505
R1846 VDD.n1231 VDD.n1230 3.1505
R1847 VDD.n1233 VDD.n1232 3.1505
R1848 VDD.n1235 VDD.n1234 3.1505
R1849 VDD.n1237 VDD.n1236 3.1505
R1850 VDD.n1240 VDD.n1239 3.1505
R1851 VDD.n1242 VDD.n1241 3.1505
R1852 VDD.n1244 VDD.n1243 3.1505
R1853 VDD.n1246 VDD.n1245 3.1505
R1854 VDD.n1248 VDD.n1247 3.1505
R1855 VDD.n1250 VDD.n1249 3.1505
R1856 VDD.n1253 VDD.n1252 3.1505
R1857 VDD.n1255 VDD.n1254 3.1505
R1858 VDD.n1257 VDD.n1256 3.1505
R1859 VDD.n1259 VDD.n1258 3.1505
R1860 VDD.n1262 VDD.n1261 3.1505
R1861 VDD.n1299 VDD.n1298 3.1505
R1862 VDD.n1297 VDD.n1296 3.1505
R1863 VDD.n1289 VDD.n1288 3.1505
R1864 VDD.n1287 VDD.n1286 3.1505
R1865 VDD.n1281 VDD.n1280 3.1505
R1866 VDD.n1279 VDD.n1278 3.1505
R1867 VDD.n1276 VDD.n1229 3.1505
R1868 VDD.n1276 VDD.n1227 3.1505
R1869 VDD.n1267 VDD.n1266 3.1505
R1870 VDD.n1270 VDD.n1269 3.1505
R1871 VDD.n1275 VDD.n1274 3.1505
R1872 VDD.n1272 VDD.n1271 3.1505
R1873 VDD.n1264 VDD.n1263 3.1505
R1874 VDD.n1694 VDD.n1693 3.1505
R1875 VDD.n1693 VDD.n1692 3.1505
R1876 VDD.n2719 VDD.n2718 3.1505
R1877 VDD.n2718 VDD.n2717 3.1505
R1878 VDD.n2716 VDD.n2715 3.1505
R1879 VDD.n2715 VDD.n2714 3.1505
R1880 VDD.n2713 VDD.n2712 3.1505
R1881 VDD.n2712 VDD.n2711 3.1505
R1882 VDD.n2710 VDD.n2709 3.1505
R1883 VDD.n2709 VDD.n2708 3.1505
R1884 VDD.n2707 VDD.n2706 3.1505
R1885 VDD.n2706 VDD.n2705 3.1505
R1886 VDD.n2704 VDD.n2703 3.1505
R1887 VDD.n2703 VDD.n2702 3.1505
R1888 VDD.n2701 VDD.n2700 3.1505
R1889 VDD.n2700 VDD.n2699 3.1505
R1890 VDD.n2698 VDD.n2697 3.1505
R1891 VDD.n2697 VDD.n2696 3.1505
R1892 VDD.n2695 VDD.n2694 3.1505
R1893 VDD.n2694 VDD.n2693 3.1505
R1894 VDD.n2692 VDD.n2691 3.1505
R1895 VDD.n2691 VDD.n2690 3.1505
R1896 VDD.n1676 VDD.n1675 3.1505
R1897 VDD.n1675 VDD.n1674 3.1505
R1898 VDD.n1679 VDD.n1678 3.1505
R1899 VDD.n1678 VDD.n1677 3.1505
R1900 VDD.n1682 VDD.n1681 3.1505
R1901 VDD.n1681 VDD.n1680 3.1505
R1902 VDD.n1685 VDD.n1684 3.1505
R1903 VDD.n1684 VDD.n1683 3.1505
R1904 VDD.n1688 VDD.n1687 3.1505
R1905 VDD.n1687 VDD.n1686 3.1505
R1906 VDD.n1691 VDD.n1690 3.1505
R1907 VDD.n1690 VDD.n1689 3.1505
R1908 VDD.n1696 VDD.n1695 3.1505
R1909 VDD.n2794 VDD.n2793 3.1505
R1910 VDD.n2750 VDD.n2749 3.1505
R1911 VDD.n2748 VDD.n2747 3.1505
R1912 VDD.n2775 VDD.n2774 3.1505
R1913 VDD.n2773 VDD.n2772 3.1505
R1914 VDD.n2796 VDD.n2795 3.1505
R1915 VDD.n2729 VDD.n2728 3.1505
R1916 VDD.n2726 VDD.n2725 3.1505
R1917 VDD.n2756 VDD.n2755 3.1505
R1918 VDD.n2724 VDD.n2723 3.1505
R1919 VDD.n2722 VDD.n2721 3.1505
R1920 VDD.n2853 VDD.n2852 3.1505
R1921 VDD.n2589 VDD.n2588 3.1505
R1922 VDD.n2587 VDD.n2586 3.1505
R1923 VDD.n2584 VDD.n2583 3.1505
R1924 VDD.n2582 VDD.n2581 3.1505
R1925 VDD.n2579 VDD.n2578 3.1505
R1926 VDD.n2577 VDD.n2576 3.1505
R1927 VDD.n2574 VDD.n2573 3.1505
R1928 VDD.n2572 VDD.n2571 3.1505
R1929 VDD.n2569 VDD.n2568 3.1505
R1930 VDD.n2567 VDD.n2566 3.1505
R1931 VDD.n2564 VDD.n2563 3.1505
R1932 VDD.n2562 VDD.n2561 3.1505
R1933 VDD.n2559 VDD.n2558 3.1505
R1934 VDD.n2557 VDD.n2556 3.1505
R1935 VDD.n2554 VDD.n2553 3.1505
R1936 VDD.n2552 VDD.n2551 3.1505
R1937 VDD.n2550 VDD.n2549 3.1505
R1938 VDD.n2548 VDD.n2547 3.1505
R1939 VDD.n2546 VDD.n2545 3.1505
R1940 VDD.n2544 VDD.n2543 3.1505
R1941 VDD.n2542 VDD.n2541 3.1505
R1942 VDD.n2540 VDD.n2539 3.1505
R1943 VDD.n2538 VDD.n2537 3.1505
R1944 VDD.n2536 VDD.n2535 3.1505
R1945 VDD.n2534 VDD.n2533 3.1505
R1946 VDD.n2532 VDD.n2531 3.1505
R1947 VDD.n2530 VDD.n2529 3.1505
R1948 VDD.n2528 VDD.n2527 3.1505
R1949 VDD.n2526 VDD.n2525 3.1505
R1950 VDD.n2524 VDD.n2523 3.1505
R1951 VDD.n2522 VDD.n2521 3.1505
R1952 VDD.n2520 VDD.n2519 3.1505
R1953 VDD.n2518 VDD.n2517 3.1505
R1954 VDD.n2845 VDD.n2844 3.1505
R1955 VDD.n2847 VDD.n2846 3.1505
R1956 VDD.n2849 VDD.n2848 3.1505
R1957 VDD.n2851 VDD.n2850 3.1505
R1958 VDD.n2895 VDD.n2894 3.1505
R1959 VDD.n2893 VDD.n2892 3.1505
R1960 VDD.n2891 VDD.n2890 3.1505
R1961 VDD.n2889 VDD.n2888 3.1505
R1962 VDD.n2887 VDD.n2886 3.1505
R1963 VDD.n2885 VDD.n2884 3.1505
R1964 VDD.n2883 VDD.n2882 3.1505
R1965 VDD.n2881 VDD.n2880 3.1505
R1966 VDD.n2879 VDD.n2878 3.1505
R1967 VDD.n2877 VDD.n2876 3.1505
R1968 VDD.n2875 VDD.n2874 3.1505
R1969 VDD.n2873 VDD.n2872 3.1505
R1970 VDD.n2871 VDD.n2870 3.1505
R1971 VDD.n2869 VDD.n2868 3.1505
R1972 VDD.n2867 VDD.n2866 3.1505
R1973 VDD.n2865 VDD.n2864 3.1505
R1974 VDD.n2863 VDD.n2862 3.1505
R1975 VDD.n2861 VDD.n2860 3.1505
R1976 VDD.n2859 VDD.n2858 3.1505
R1977 VDD.n2857 VDD.n2856 3.1505
R1978 VDD.n2855 VDD.n2854 3.1505
R1979 VDD.n2897 VDD.n2896 3.1505
R1980 VDD.n2668 VDD.n2667 3.1505
R1981 VDD.n2621 VDD.n2620 3.1505
R1982 VDD.n2624 VDD.n2623 3.1505
R1983 VDD.n2627 VDD.n2626 3.1505
R1984 VDD.n2619 VDD.n2618 3.1505
R1985 VDD.n2688 VDD.n2687 3.1505
R1986 VDD.n2732 VDD.n2731 3.1505
R1987 VDD.n2671 VDD.n2670 3.1505
R1988 VDD.n2673 VDD.n2672 3.1505
R1989 VDD.n2676 VDD.n2675 3.1505
R1990 VDD.n2678 VDD.n2677 3.1505
R1991 VDD.n2681 VDD.n2680 3.1505
R1992 VDD.n2683 VDD.n2682 3.1505
R1993 VDD.n2686 VDD.n2685 3.1505
R1994 VDD.n2734 VDD.n2733 3.1505
R1995 VDD.n2737 VDD.n2736 3.1505
R1996 VDD.n2745 VDD.n2744 3.1505
R1997 VDD.n2759 VDD.n2758 3.1505
R1998 VDD.n2740 VDD.n2739 3.1505
R1999 VDD.n2742 VDD.n2741 3.1505
R2000 VDD.n2767 VDD.n2766 3.1505
R2001 VDD.n2764 VDD.n2763 3.1505
R2002 VDD.n2778 VDD.n2777 3.1505
R2003 VDD.n2762 VDD.n2761 3.1505
R2004 VDD.n2781 VDD.n2780 3.1505
R2005 VDD.n2788 VDD.n2787 3.1505
R2006 VDD.n2783 VDD.n2782 3.1505
R2007 VDD.n2786 VDD.n2785 3.1505
R2008 VDD.n2800 VDD.n2799 3.1505
R2009 VDD.n2807 VDD.n2806 3.1505
R2010 VDD.n2810 VDD.n2809 3.1505
R2011 VDD.n2802 VDD.n2801 3.1505
R2012 VDD.n2805 VDD.n2804 3.1505
R2013 VDD.n2818 VDD.n2817 3.1505
R2014 VDD.n2812 VDD.n2811 3.1505
R2015 VDD.n2815 VDD.n2814 3.1505
R2016 VDD.n2902 VDD.n2901 3.1505
R2017 VDD.n2590 VDD.n2516 3.1505
R2018 VDD.n2614 VDD.n2613 3.1505
R2019 VDD.n2465 VDD.n2464 3.1505
R2020 VDD.n2492 VDD.n2491 3.1505
R2021 VDD.n2491 VDD.n2490 3.1505
R2022 VDD.n2495 VDD.n2494 3.1505
R2023 VDD.n2494 VDD.n2493 3.1505
R2024 VDD.n2499 VDD.n2498 3.1505
R2025 VDD.n2497 VDD.n2496 3.1505
R2026 VDD.n2480 VDD.n2479 3.1505
R2027 VDD.n2479 VDD.n2478 3.1505
R2028 VDD.n2483 VDD.n2482 3.1505
R2029 VDD.n2482 VDD.n2481 3.1505
R2030 VDD.n2487 VDD.n2486 3.1505
R2031 VDD.n2485 VDD.n2484 3.1505
R2032 VDD.n2468 VDD.n2467 3.1505
R2033 VDD.n2467 VDD.n2466 3.1505
R2034 VDD.n2471 VDD.n2470 3.1505
R2035 VDD.n2470 VDD.n2469 3.1505
R2036 VDD.n2475 VDD.n2474 3.1505
R2037 VDD.n2473 VDD.n2472 3.1505
R2038 VDD.n2454 VDD.n2453 3.1505
R2039 VDD.n2453 VDD.n2452 3.1505
R2040 VDD.n2457 VDD.n2456 3.1505
R2041 VDD.n2456 VDD.n2455 3.1505
R2042 VDD.n2464 VDD.n2463 3.1505
R2043 VDD.n2461 VDD.n2460 3.1505
R2044 VDD.n2459 VDD.n2458 3.1505
R2045 VDD.n2371 VDD.n2370 3.1505
R2046 VDD.n3059 VDD.n3058 3.1505
R2047 VDD.n3089 VDD.n3088 3.1505
R2048 VDD.n3092 VDD.n3091 3.1505
R2049 VDD.n3067 VDD.n3066 3.1505
R2050 VDD.n3046 VDD.n3045 3.1505
R2051 VDD.n3061 VDD.n3060 3.1505
R2052 VDD.n3064 VDD.n3063 3.1505
R2053 VDD.n3049 VDD.n3048 3.1505
R2054 VDD.n3056 VDD.n3055 3.1505
R2055 VDD.n3051 VDD.n3050 3.1505
R2056 VDD.n3053 VDD.n3052 3.1505
R2057 VDD.n3036 VDD.n3035 3.1505
R2058 VDD.n3043 VDD.n3042 3.1505
R2059 VDD.n3038 VDD.n3037 3.1505
R2060 VDD.n3040 VDD.n3039 3.1505
R2061 VDD.n3024 VDD.n3023 3.1505
R2062 VDD.n3032 VDD.n3031 3.1505
R2063 VDD.n3012 VDD.n3011 3.1505
R2064 VDD.n3027 VDD.n3026 3.1505
R2065 VDD.n3029 VDD.n3028 3.1505
R2066 VDD.n3020 VDD.n3019 3.1505
R2067 VDD.n3017 VDD.n3016 3.1505
R2068 VDD.n2924 VDD.n2923 3.1505
R2069 VDD.n3015 VDD.n3014 3.1505
R2070 VDD.n2927 VDD.n2926 3.1505
R2071 VDD.n3009 VDD.n3008 3.1505
R2072 VDD.n3007 VDD.n3006 3.1505
R2073 VDD.n3004 VDD.n3003 3.1505
R2074 VDD.n3097 VDD.n3096 3.1505
R2075 VDD.n3087 VDD.n3086 3.1505
R2076 VDD.n3085 VDD.n3084 3.1505
R2077 VDD.n3082 VDD.n3081 3.1505
R2078 VDD.n3080 VDD.n3079 3.1505
R2079 VDD.n2369 VDD.n2368 3.1505
R2080 VDD.n2300 VDD.n2299 3.1505
R2081 VDD.n2299 VDD.n2298 3.1505
R2082 VDD.n2303 VDD.n2302 3.1505
R2083 VDD.n2302 VDD.n2301 3.1505
R2084 VDD.n2306 VDD.n2305 3.1505
R2085 VDD.n2305 VDD.n2304 3.1505
R2086 VDD.n2309 VDD.n2308 3.1505
R2087 VDD.n2308 VDD.n2307 3.1505
R2088 VDD.n2312 VDD.n2311 3.1505
R2089 VDD.n2311 VDD.n2310 3.1505
R2090 VDD.n2315 VDD.n2314 3.1505
R2091 VDD.n2314 VDD.n2313 3.1505
R2092 VDD.n2318 VDD.n2317 3.1505
R2093 VDD.n2317 VDD.n2316 3.1505
R2094 VDD.n2321 VDD.n2320 3.1505
R2095 VDD.n2320 VDD.n2319 3.1505
R2096 VDD.n2325 VDD.n2324 3.1505
R2097 VDD.n2324 VDD.n2323 3.1505
R2098 VDD.n2328 VDD.n2327 3.1505
R2099 VDD.n2327 VDD.n2326 3.1505
R2100 VDD.n2331 VDD.n2330 3.1505
R2101 VDD.n2330 VDD.n2329 3.1505
R2102 VDD.n2334 VDD.n2333 3.1505
R2103 VDD.n2333 VDD.n2332 3.1505
R2104 VDD.n2344 VDD.n2343 3.1505
R2105 VDD.n2343 VDD.n2342 3.1505
R2106 VDD.n2347 VDD.n2346 3.1505
R2107 VDD.n2346 VDD.n2345 3.1505
R2108 VDD.n2350 VDD.n2349 3.1505
R2109 VDD.n2349 VDD.n2348 3.1505
R2110 VDD.n2353 VDD.n2352 3.1505
R2111 VDD.n2352 VDD.n2351 3.1505
R2112 VDD.n2356 VDD.n2355 3.1505
R2113 VDD.n2355 VDD.n2354 3.1505
R2114 VDD.n2359 VDD.n2358 3.1505
R2115 VDD.n2358 VDD.n2357 3.1505
R2116 VDD.n2362 VDD.n2361 3.1505
R2117 VDD.n2361 VDD.n2360 3.1505
R2118 VDD.n2365 VDD.n2364 3.1505
R2119 VDD.n2364 VDD.n2363 3.1505
R2120 VDD.n2367 VDD.n2366 3.1505
R2121 VDD.n2296 VDD.n2295 3.1505
R2122 VDD.n2278 VDD.n2277 3.1505
R2123 VDD.n2275 VDD.n2274 3.1505
R2124 VDD.n2273 VDD.n2272 3.1505
R2125 VDD.n2270 VDD.n2269 3.1505
R2126 VDD.n2268 VDD.n2267 3.1505
R2127 VDD.n2265 VDD.n2264 3.1505
R2128 VDD.n2263 VDD.n2262 3.1505
R2129 VDD.n2260 VDD.n2259 3.1505
R2130 VDD.n2258 VDD.n2257 3.1505
R2131 VDD.n2255 VDD.n2254 3.1505
R2132 VDD.n2253 VDD.n2252 3.1505
R2133 VDD.n2250 VDD.n2249 3.1505
R2134 VDD.n2248 VDD.n2247 3.1505
R2135 VDD.n2246 VDD.n2245 3.1505
R2136 VDD.n2244 VDD.n2243 3.1505
R2137 VDD.n2242 VDD.n2241 3.1505
R2138 VDD.n2240 VDD.n2239 3.1505
R2139 VDD.n2238 VDD.n2237 3.1505
R2140 VDD.n2236 VDD.n2235 3.1505
R2141 VDD.n2234 VDD.n2233 3.1505
R2142 VDD.n2232 VDD.n2231 3.1505
R2143 VDD.n2230 VDD.n2229 3.1505
R2144 VDD.n2228 VDD.n2227 3.1505
R2145 VDD.n2226 VDD.n2225 3.1505
R2146 VDD.n2938 VDD.n2937 3.1505
R2147 VDD.n2940 VDD.n2939 3.1505
R2148 VDD.n2942 VDD.n2941 3.1505
R2149 VDD.n2944 VDD.n2943 3.1505
R2150 VDD.n2946 VDD.n2945 3.1505
R2151 VDD.n2948 VDD.n2947 3.1505
R2152 VDD.n2950 VDD.n2949 3.1505
R2153 VDD.n2952 VDD.n2951 3.1505
R2154 VDD.n2954 VDD.n2953 3.1505
R2155 VDD.n2956 VDD.n2955 3.1505
R2156 VDD.n2280 VDD.n2279 3.1505
R2157 VDD.n2992 VDD.n2991 3.1505
R2158 VDD.n2958 VDD.n2957 3.1505
R2159 VDD.n2961 VDD.n2960 3.1505
R2160 VDD.n2967 VDD.n2966 3.1505
R2161 VDD.n2969 VDD.n2968 3.1505
R2162 VDD.n2975 VDD.n2974 3.1505
R2163 VDD.n2981 VDD.n2980 3.1505
R2164 VDD.n2984 VDD.n2983 3.1505
R2165 VDD.n2987 VDD.n2986 3.1505
R2166 VDD.n2994 VDD.n2993 3.1505
R2167 VDD.n2996 VDD.n2995 3.1505
R2168 VDD.n3002 VDD.n3001 3.1505
R2169 VDD.n2597 VDD.n2596 3.1505
R2170 VDD.n2595 VDD.n2594 3.1505
R2171 VDD.n2592 VDD.n2591 3.1505
R2172 VDD.n2914 VDD.n2905 3.1505
R2173 VDD.n2913 VDD.n2912 3.1505
R2174 VDD.n2910 VDD.n2909 3.1505
R2175 VDD.n2822 VDD.n2821 3.1505
R2176 VDD.n2842 VDD.n2841 3.1505
R2177 VDD.n1641 VDD.n1640 3.1505
R2178 VDD.n1639 VDD.n1638 3.1505
R2179 VDD.n1637 VDD.n1636 3.1505
R2180 VDD.n1635 VDD.n1634 3.1505
R2181 VDD.n1633 VDD.n1632 3.1505
R2182 VDD.n1631 VDD.n1630 3.1505
R2183 VDD.n1629 VDD.n1628 3.1505
R2184 VDD.n1627 VDD.n1626 3.1505
R2185 VDD.n1625 VDD.n1624 3.1505
R2186 VDD.n2824 VDD.n2823 3.1505
R2187 VDD.n2826 VDD.n2825 3.1505
R2188 VDD.n2828 VDD.n2827 3.1505
R2189 VDD.n2830 VDD.n2829 3.1505
R2190 VDD.n2832 VDD.n2831 3.1505
R2191 VDD.n2834 VDD.n2833 3.1505
R2192 VDD.n2836 VDD.n2835 3.1505
R2193 VDD.n2838 VDD.n2837 3.1505
R2194 VDD.n2840 VDD.n2839 3.1505
R2195 VDD.n1654 VDD.n1617 3.1505
R2196 VDD.n1643 VDD.n1642 3.1505
R2197 VDD.n1700 VDD.n1699 3.1505
R2198 VDD.n1698 VDD.n1697 3.1505
R2199 VDD.n1665 VDD.n1664 3.1505
R2200 VDD.n1668 VDD.n1667 3.1505
R2201 VDD.n1656 VDD.n1655 3.1505
R2202 VDD.n1659 VDD.n1658 3.1505
R2203 VDD.n1651 VDD.n1650 3.1505
R2204 VDD.n1653 VDD.n1652 3.1505
R2205 VDD.n1646 VDD.n1645 3.1505
R2206 VDD.n1648 VDD.n1647 3.1505
R2207 VDD.n1663 VDD.n1661 3.1505
R2208 VDD.n1663 VDD.n1662 3.1505
R2209 VDD.n1779 VDD.n1778 3.1505
R2210 VDD.n1756 VDD.n1755 3.1505
R2211 VDD.n1748 VDD.n1747 3.1505
R2212 VDD.n1746 VDD.n1745 3.1505
R2213 VDD.n1754 VDD.n1753 3.1505
R2214 VDD.n1762 VDD.n1761 3.1505
R2215 VDD.n1764 VDD.n1763 3.1505
R2216 VDD.n1772 VDD.n1771 3.1505
R2217 VDD.n1774 VDD.n1773 3.1505
R2218 VDD.n1777 VDD.n1776 3.1505
R2219 VDD.n1740 VDD.n1739 3.1505
R2220 VDD.n1871 VDD.n1870 3.1505
R2221 VDD.n1869 VDD.n1868 3.1505
R2222 VDD.n1866 VDD.n1865 3.1505
R2223 VDD.n1864 VDD.n1863 3.1505
R2224 VDD.n1862 VDD.n1861 3.1505
R2225 VDD.n1859 VDD.n1858 3.1505
R2226 VDD.n1857 VDD.n1856 3.1505
R2227 VDD.n1707 VDD.n1706 3.1505
R2228 VDD.n1709 VDD.n1708 3.1505
R2229 VDD.n1711 VDD.n1710 3.1505
R2230 VDD.n1713 VDD.n1712 3.1505
R2231 VDD.n1716 VDD.n1715 3.1505
R2232 VDD.n1718 VDD.n1717 3.1505
R2233 VDD.n1720 VDD.n1719 3.1505
R2234 VDD.n1722 VDD.n1721 3.1505
R2235 VDD.n1724 VDD.n1723 3.1505
R2236 VDD.n1726 VDD.n1725 3.1505
R2237 VDD.n1729 VDD.n1728 3.1505
R2238 VDD.n1731 VDD.n1730 3.1505
R2239 VDD.n1734 VDD.n1733 3.1505
R2240 VDD.n1736 VDD.n1735 3.1505
R2241 VDD.n1738 VDD.n1737 3.1505
R2242 VDD.n1873 VDD.n1872 3.1505
R2243 VDD.n1888 VDD.n1887 3.1505
R2244 VDD.n1897 VDD.n1896 3.1505
R2245 VDD.n1907 VDD.n1906 3.1505
R2246 VDD.n1912 VDD.n1911 3.1505
R2247 VDD.n1909 VDD.n1908 3.1505
R2248 VDD.n1904 VDD.n1902 3.1505
R2249 VDD.n1904 VDD.n1903 3.1505
R2250 VDD.n1900 VDD.n1899 3.1505
R2251 VDD.n1895 VDD.n1893 3.1505
R2252 VDD.n1895 VDD.n1894 3.1505
R2253 VDD.n1891 VDD.n1890 3.1505
R2254 VDD.n1886 VDD.n1885 3.1505
R2255 VDD.n1880 VDD.n1879 3.1505
R2256 VDD.n1878 VDD.n1877 3.1505
R2257 VDD.n1875 VDD.n1874 3.1505
R2258 VDD.n1917 VDD.n1916 3.1505
R2259 VDD.n1808 VDD.n1807 3.1505
R2260 VDD.n1846 VDD.n1845 3.1505
R2261 VDD.n1848 VDD.n1847 3.1505
R2262 VDD.n1916 VDD.n1915 3.1505
R2263 VDD.n1920 VDD.n1919 3.1505
R2264 VDD.n1919 VDD.n1918 3.1505
R2265 VDD.n1840 VDD.n1839 3.1505
R2266 VDD.n1838 VDD.n1837 3.1505
R2267 VDD.n1832 VDD.n1831 3.1505
R2268 VDD.n1831 VDD.n1830 3.1505
R2269 VDD.n1835 VDD.n1834 3.1505
R2270 VDD.n1834 VDD.n1833 3.1505
R2271 VDD.n1826 VDD.n1825 3.1505
R2272 VDD.n1824 VDD.n1823 3.1505
R2273 VDD.n1811 VDD.n1810 3.1505
R2274 VDD.n1810 VDD.n1809 3.1505
R2275 VDD.n1814 VDD.n1813 3.1505
R2276 VDD.n1813 VDD.n1812 3.1505
R2277 VDD.n1807 VDD.n1806 3.1505
R2278 VDD.n1798 VDD.n1797 3.1505
R2279 VDD.n1797 VDD.n1796 3.1505
R2280 VDD.n1801 VDD.n1800 3.1505
R2281 VDD.n1800 VDD.n1799 3.1505
R2282 VDD.n1804 VDD.n1803 3.1505
R2283 VDD.n1803 VDD.n1802 3.1505
R2284 VDD.n1793 VDD.n1792 3.1505
R2285 VDD.n1791 VDD.n1790 3.1505
R2286 VDD.n1789 VDD.n1788 3.1505
R2287 VDD.n1788 VDD.n1787 3.1505
R2288 VDD.n1785 VDD.n1784 3.1505
R2289 VDD.n1784 VDD.n1783 3.1505
R2290 VDD.n1782 VDD.n1781 3.1505
R2291 VDD.n1816 VDD.n1815 3.1505
R2292 VDD.n1818 VDD.n1817 3.1505
R2293 VDD.n175 VDD.n174 3.1505
R2294 VDD.n1468 VDD.n1467 3.1505
R2295 VDD.n1449 VDD.n1448 3.1505
R2296 VDD.n1429 VDD.n1428 3.1505
R2297 VDD.n1410 VDD.n1409 3.1505
R2298 VDD.n1393 VDD.n1392 3.1505
R2299 VDD.n1376 VDD.n1375 3.1505
R2300 VDD.n1215 VDD.n1213 3.1505
R2301 VDD.n173 VDD.n172 3.1505
R2302 VDD.n1508 VDD.n1507 3.1505
R2303 VDD.n1503 VDD.n1502 3.1505
R2304 VDD.n1491 VDD.n1490 3.1505
R2305 VDD.n1486 VDD.n1485 3.1505
R2306 VDD.n1483 VDD.n1482 3.1505
R2307 VDD.n1472 VDD.n1469 3.1505
R2308 VDD.n1472 VDD.n1471 3.1505
R2309 VDD.n1465 VDD.n1464 3.1505
R2310 VDD.n1453 VDD.n1450 3.1505
R2311 VDD.n1453 VDD.n1452 3.1505
R2312 VDD.n1446 VDD.n1445 3.1505
R2313 VDD.n1431 VDD.n1430 3.1505
R2314 VDD.n1412 VDD.n1411 3.1505
R2315 VDD.n1408 VDD.n1407 3.1505
R2316 VDD.n1391 VDD.n1390 3.1505
R2317 VDD.n1374 VDD.n1373 3.1505
R2318 VDD.n1135 VDD.n1134 3.1505
R2319 VDD.n1215 VDD.n1214 3.1505
R2320 VDD.n185 VDD.n184 3.1505
R2321 VDD.n747 VDD.n746 3.1505
R2322 VDD.n744 VDD.n743 3.1505
R2323 VDD.n742 VDD.n741 3.1505
R2324 VDD.n739 VDD.n738 3.1505
R2325 VDD.n737 VDD.n736 3.1505
R2326 VDD.n1154 VDD.n1153 3.1505
R2327 VDD.n1156 VDD.n1155 3.1505
R2328 VDD.n1159 VDD.n1158 3.1505
R2329 VDD.n1161 VDD.n1160 3.1505
R2330 VDD.n1173 VDD.n1172 3.1505
R2331 VDD.n1175 VDD.n1174 3.1505
R2332 VDD.n1187 VDD.n1186 3.1505
R2333 VDD.n1189 VDD.n1188 3.1505
R2334 VDD.n1196 VDD.n1195 3.1505
R2335 VDD.n1204 VDD.n1203 3.1505
R2336 VDD.n1206 VDD.n1205 3.1505
R2337 VDD.n1210 VDD.n1209 3.1505
R2338 VDD.n1212 VDD.n1211 3.1505
R2339 VDD.n749 VDD.n748 3.1505
R2340 VDD.n287 VDD.n286 3.1505
R2341 VDD.n825 VDD.n824 3.1505
R2342 VDD.n632 VDD.n631 3.1505
R2343 VDD.n723 VDD.n722 3.1505
R2344 VDD.n629 VDD.n628 3.1505
R2345 VDD.n766 VDD.n765 3.1505
R2346 VDD.n768 VDD.n767 3.1505
R2347 VDD.n787 VDD.n786 3.1505
R2348 VDD.n789 VDD.n788 3.1505
R2349 VDD.n785 VDD.n784 3.1505
R2350 VDD.n804 VDD.n803 3.1505
R2351 VDD.n806 VDD.n805 3.1505
R2352 VDD.n823 VDD.n822 3.1505
R2353 VDD.n843 VDD.n842 3.1505
R2354 VDD.n845 VDD.n844 3.1505
R2355 VDD.n847 VDD.n846 3.1505
R2356 VDD.n863 VDD.n862 3.1505
R2357 VDD.n274 VDD.n273 3.1505
R2358 VDD.n276 VDD.n275 3.1505
R2359 VDD.n282 VDD.n281 3.1505
R2360 VDD.n285 VDD.n284 3.1505
R2361 VDD.n757 VDD.n756 3.1505
R2362 VDD.n777 VDD.n776 3.1505
R2363 VDD.n775 VDD.n774 3.1505
R2364 VDD.n796 VDD.n795 3.1505
R2365 VDD.n834 VDD.n833 3.1505
R2366 VDD.n832 VDD.n831 3.1505
R2367 VDD.n854 VDD.n853 3.1505
R2368 VDD.n870 VDD.n869 3.1505
R2369 VDD.n309 VDD.n308 3.1505
R2370 VDD.n300 VDD.n299 3.1505
R2371 VDD.n298 VDD.n297 3.1505
R2372 VDD.n877 VDD.n874 3.1505
R2373 VDD.n877 VDD.n876 3.1505
R2374 VDD.n873 VDD.n872 3.1505
R2375 VDD.n861 VDD.n859 3.1505
R2376 VDD.n861 VDD.n860 3.1505
R2377 VDD.n857 VDD.n856 3.1505
R2378 VDD.n841 VDD.n839 3.1505
R2379 VDD.n841 VDD.n840 3.1505
R2380 VDD.n837 VDD.n836 3.1505
R2381 VDD.n820 VDD.n818 3.1505
R2382 VDD.n820 VDD.n819 3.1505
R2383 VDD.n816 VDD.n815 3.1505
R2384 VDD.n813 VDD.n812 3.1505
R2385 VDD.n798 VDD.n797 3.1505
R2386 VDD.n779 VDD.n778 3.1505
R2387 VDD.n759 VDD.n758 3.1505
R2388 VDD.n623 VDD.n622 3.1505
R2389 VDD.n621 VDD.n620 3.1505
R2390 VDD.n716 VDD.n715 3.1505
R2391 VDD.n448 VDD.n447 3.1505
R2392 VDD.n445 VDD.n444 3.1505
R2393 VDD.n443 VDD.n442 3.1505
R2394 VDD.n440 VDD.n439 3.1505
R2395 VDD.n438 VDD.n437 3.1505
R2396 VDD.n672 VDD.n671 3.1505
R2397 VDD.n674 VDD.n673 3.1505
R2398 VDD.n677 VDD.n676 3.1505
R2399 VDD.n679 VDD.n678 3.1505
R2400 VDD.n681 VDD.n680 3.1505
R2401 VDD.n684 VDD.n683 3.1505
R2402 VDD.n686 VDD.n685 3.1505
R2403 VDD.n688 VDD.n687 3.1505
R2404 VDD.n691 VDD.n690 3.1505
R2405 VDD.n693 VDD.n692 3.1505
R2406 VDD.n695 VDD.n694 3.1505
R2407 VDD.n697 VDD.n696 3.1505
R2408 VDD.n700 VDD.n699 3.1505
R2409 VDD.n702 VDD.n701 3.1505
R2410 VDD.n704 VDD.n703 3.1505
R2411 VDD.n707 VDD.n706 3.1505
R2412 VDD.n709 VDD.n708 3.1505
R2413 VDD.n712 VDD.n711 3.1505
R2414 VDD.n714 VDD.n713 3.1505
R2415 VDD.n450 VDD.n449 3.1505
R2416 VDD.n519 VDD.n518 3.1505
R2417 VDD.n517 VDD.n516 3.1505
R2418 VDD.n505 VDD.n504 3.1505
R2419 VDD.n503 VDD.n502 3.1505
R2420 VDD.n476 VDD.n475 3.1505
R2421 VDD.n466 VDD.n465 3.1505
R2422 VDD.n455 VDD.n454 3.1505
R2423 VDD.n453 VDD.n452 3.1505
R2424 VDD.n464 VDD.n463 3.1505
R2425 VDD.n461 VDD.n460 3.1505
R2426 VDD.n474 VDD.n473 3.1505
R2427 VDD.n483 VDD.n482 3.1505
R2428 VDD.n485 VDD.n484 3.1505
R2429 VDD.n488 VDD.n487 3.1505
R2430 VDD.n491 VDD.n490 3.1505
R2431 VDD.n494 VDD.n493 3.1505
R2432 VDD.n497 VDD.n496 3.1505
R2433 VDD.n500 VDD.n499 3.1505
R2434 VDD.n420 VDD.n419 3.1505
R2435 VDD.n419 VDD.n418 3.1505
R2436 VDD.n513 VDD.n512 3.1505
R2437 VDD.n529 VDD.n521 3.1505
R2438 VDD.n405 VDD.n404 3.1505
R2439 VDD.n407 VDD.n406 3.1505
R2440 VDD.n410 VDD.n409 3.1505
R2441 VDD.n413 VDD.n412 3.1505
R2442 VDD.n416 VDD.n415 3.1505
R2443 VDD.n402 VDD.n401 3.1505
R2444 VDD.n539 VDD.n538 3.1505
R2445 VDD.n542 VDD.n541 3.1505
R2446 VDD.n541 VDD.n540 3.1505
R2447 VDD.n546 VDD.n545 3.1505
R2448 VDD.n545 VDD.n544 3.1505
R2449 VDD.n549 VDD.n548 3.1505
R2450 VDD.n548 VDD.n547 3.1505
R2451 VDD.n553 VDD.n552 3.1505
R2452 VDD.n552 VDD.n551 3.1505
R2453 VDD.n556 VDD.n555 3.1505
R2454 VDD.n555 VDD.n554 3.1505
R2455 VDD.n559 VDD.n558 3.1505
R2456 VDD.n558 VDD.n557 3.1505
R2457 VDD.n562 VDD.n561 3.1505
R2458 VDD.n561 VDD.n560 3.1505
R2459 VDD.n566 VDD.n565 3.1505
R2460 VDD.n565 VDD.n564 3.1505
R2461 VDD.n569 VDD.n568 3.1505
R2462 VDD.n568 VDD.n567 3.1505
R2463 VDD.n572 VDD.n571 3.1505
R2464 VDD.n571 VDD.n570 3.1505
R2465 VDD.n576 VDD.n575 3.1505
R2466 VDD.n575 VDD.n574 3.1505
R2467 VDD.n579 VDD.n578 3.1505
R2468 VDD.n578 VDD.n577 3.1505
R2469 VDD.n582 VDD.n581 3.1505
R2470 VDD.n581 VDD.n580 3.1505
R2471 VDD.n586 VDD.n585 3.1505
R2472 VDD.n585 VDD.n584 3.1505
R2473 VDD.n589 VDD.n588 3.1505
R2474 VDD.n588 VDD.n587 3.1505
R2475 VDD.n592 VDD.n591 3.1505
R2476 VDD.n591 VDD.n590 3.1505
R2477 VDD.n595 VDD.n594 3.1505
R2478 VDD.n594 VDD.n593 3.1505
R2479 VDD.n599 VDD.n598 3.1505
R2480 VDD.n598 VDD.n597 3.1505
R2481 VDD.n602 VDD.n601 3.1505
R2482 VDD.n601 VDD.n600 3.1505
R2483 VDD.n605 VDD.n604 3.1505
R2484 VDD.n604 VDD.n603 3.1505
R2485 VDD.n609 VDD.n608 3.1505
R2486 VDD.n608 VDD.n607 3.1505
R2487 VDD.n612 VDD.n611 3.1505
R2488 VDD.n611 VDD.n610 3.1505
R2489 VDD.n616 VDD.n615 3.1505
R2490 VDD.n615 VDD.n614 3.1505
R2491 VDD.n618 VDD.n617 3.1505
R2492 VDD.n295 VDD.n294 3.1505
R2493 VDD.n883 VDD.n882 3.1505
R2494 VDD.n886 VDD.n885 3.1505
R2495 VDD.n885 VDD.n884 3.1505
R2496 VDD.n890 VDD.n889 3.1505
R2497 VDD.n889 VDD.n888 3.1505
R2498 VDD.n893 VDD.n892 3.1505
R2499 VDD.n892 VDD.n891 3.1505
R2500 VDD.n897 VDD.n896 3.1505
R2501 VDD.n896 VDD.n895 3.1505
R2502 VDD.n900 VDD.n899 3.1505
R2503 VDD.n899 VDD.n898 3.1505
R2504 VDD.n903 VDD.n902 3.1505
R2505 VDD.n902 VDD.n901 3.1505
R2506 VDD.n906 VDD.n905 3.1505
R2507 VDD.n905 VDD.n904 3.1505
R2508 VDD.n910 VDD.n909 3.1505
R2509 VDD.n909 VDD.n908 3.1505
R2510 VDD.n913 VDD.n912 3.1505
R2511 VDD.n912 VDD.n911 3.1505
R2512 VDD.n916 VDD.n915 3.1505
R2513 VDD.n915 VDD.n914 3.1505
R2514 VDD.n920 VDD.n919 3.1505
R2515 VDD.n919 VDD.n918 3.1505
R2516 VDD.n923 VDD.n922 3.1505
R2517 VDD.n922 VDD.n921 3.1505
R2518 VDD.n926 VDD.n925 3.1505
R2519 VDD.n925 VDD.n924 3.1505
R2520 VDD.n930 VDD.n929 3.1505
R2521 VDD.n929 VDD.n928 3.1505
R2522 VDD.n933 VDD.n932 3.1505
R2523 VDD.n932 VDD.n931 3.1505
R2524 VDD.n936 VDD.n935 3.1505
R2525 VDD.n935 VDD.n934 3.1505
R2526 VDD.n939 VDD.n938 3.1505
R2527 VDD.n938 VDD.n937 3.1505
R2528 VDD.n943 VDD.n942 3.1505
R2529 VDD.n942 VDD.n941 3.1505
R2530 VDD.n946 VDD.n945 3.1505
R2531 VDD.n945 VDD.n944 3.1505
R2532 VDD.n949 VDD.n948 3.1505
R2533 VDD.n948 VDD.n947 3.1505
R2534 VDD.n953 VDD.n952 3.1505
R2535 VDD.n952 VDD.n951 3.1505
R2536 VDD.n956 VDD.n955 3.1505
R2537 VDD.n955 VDD.n954 3.1505
R2538 VDD.n960 VDD.n959 3.1505
R2539 VDD.n959 VDD.n958 3.1505
R2540 VDD.n962 VDD.n961 3.1505
R2541 VDD.n1515 VDD.n1514 3.1505
R2542 VDD.n1518 VDD.n1517 3.1505
R2543 VDD.n1517 VDD.n1516 3.1505
R2544 VDD.n1522 VDD.n1521 3.1505
R2545 VDD.n1521 VDD.n1520 3.1505
R2546 VDD.n1525 VDD.n1524 3.1505
R2547 VDD.n1524 VDD.n1523 3.1505
R2548 VDD.n1529 VDD.n1528 3.1505
R2549 VDD.n1528 VDD.n1527 3.1505
R2550 VDD.n1532 VDD.n1531 3.1505
R2551 VDD.n1531 VDD.n1530 3.1505
R2552 VDD.n1535 VDD.n1534 3.1505
R2553 VDD.n1534 VDD.n1533 3.1505
R2554 VDD.n1538 VDD.n1537 3.1505
R2555 VDD.n1537 VDD.n1536 3.1505
R2556 VDD.n1542 VDD.n1541 3.1505
R2557 VDD.n1541 VDD.n1540 3.1505
R2558 VDD.n1545 VDD.n1544 3.1505
R2559 VDD.n1544 VDD.n1543 3.1505
R2560 VDD.n1548 VDD.n1547 3.1505
R2561 VDD.n1547 VDD.n1546 3.1505
R2562 VDD.n1552 VDD.n1551 3.1505
R2563 VDD.n1551 VDD.n1550 3.1505
R2564 VDD.n1555 VDD.n1554 3.1505
R2565 VDD.n1554 VDD.n1553 3.1505
R2566 VDD.n1558 VDD.n1557 3.1505
R2567 VDD.n1557 VDD.n1556 3.1505
R2568 VDD.n1562 VDD.n1561 3.1505
R2569 VDD.n1561 VDD.n1560 3.1505
R2570 VDD.n1565 VDD.n1564 3.1505
R2571 VDD.n1564 VDD.n1563 3.1505
R2572 VDD.n1568 VDD.n1567 3.1505
R2573 VDD.n1567 VDD.n1566 3.1505
R2574 VDD.n1571 VDD.n1570 3.1505
R2575 VDD.n1570 VDD.n1569 3.1505
R2576 VDD.n1575 VDD.n1574 3.1505
R2577 VDD.n1574 VDD.n1573 3.1505
R2578 VDD.n1578 VDD.n1577 3.1505
R2579 VDD.n1577 VDD.n1576 3.1505
R2580 VDD.n1581 VDD.n1580 3.1505
R2581 VDD.n1580 VDD.n1579 3.1505
R2582 VDD.n1585 VDD.n1584 3.1505
R2583 VDD.n1584 VDD.n1583 3.1505
R2584 VDD.n1588 VDD.n1587 3.1505
R2585 VDD.n1587 VDD.n1586 3.1505
R2586 VDD.n1592 VDD.n1591 3.1505
R2587 VDD.n1591 VDD.n1590 3.1505
R2588 VDD.n1594 VDD.n1593 3.1505
R2589 VDD.n1367 VDD.n1366 3.1505
R2590 VDD.n1399 VDD.n1398 3.1505
R2591 VDD.n1420 VDD.n1419 3.1505
R2592 VDD.n1418 VDD.n1417 3.1505
R2593 VDD.n1437 VDD.n1436 3.1505
R2594 VDD.n1474 VDD.n1473 3.1505
R2595 VDD.n1494 VDD.n1493 3.1505
R2596 VDD.n149 VDD.n148 3.1505
R2597 VDD.n162 VDD.n161 3.1505
R2598 VDD.n157 VDD.n156 3.1505
R2599 VDD.n160 VDD.n159 3.1505
R2600 VDD.n151 VDD.n150 3.1505
R2601 VDD.n1496 VDD.n1495 3.1505
R2602 VDD.n1476 VDD.n1475 3.1505
R2603 VDD.n1458 VDD.n1457 3.1505
R2604 VDD.n1456 VDD.n1455 3.1505
R2605 VDD.n1439 VDD.n1438 3.1505
R2606 VDD.n1422 VDD.n1421 3.1505
R2607 VDD.n1401 VDD.n1400 3.1505
R2608 VDD.n1384 VDD.n1383 3.1505
R2609 VDD.n1382 VDD.n1381 3.1505
R2610 VDD.n171 VDD.n170 3.1505
R2611 VDD.n1362 VDD.n1361 3.1505
R2612 VDD.n1359 VDD.n1358 3.1505
R2613 VDD.n1357 VDD.n1356 3.1505
R2614 VDD.n1354 VDD.n1353 3.1505
R2615 VDD.n1352 VDD.n1351 3.1505
R2616 VDD.n1349 VDD.n1348 3.1505
R2617 VDD.n1347 VDD.n1346 3.1505
R2618 VDD.n1954 VDD.n1953 3.1505
R2619 VDD.n1956 VDD.n1955 3.1505
R2620 VDD.n1968 VDD.n1967 3.1505
R2621 VDD.n1970 VDD.n1969 3.1505
R2622 VDD.n1977 VDD.n1976 3.1505
R2623 VDD.n1985 VDD.n1984 3.1505
R2624 VDD.n1987 VDD.n1986 3.1505
R2625 VDD.n1991 VDD.n1990 3.1505
R2626 VDD.n1993 VDD.n1992 3.1505
R2627 VDD.n1365 VDD.n1364 3.1505
R2628 VDD.n2161 VDD.n2160 3.1505
R2629 VDD.n2141 VDD.n2140 3.1505
R2630 VDD.n2120 VDD.n2119 3.1505
R2631 VDD.n2098 VDD.n2097 3.1505
R2632 VDD.n2076 VDD.n2075 3.1505
R2633 VDD.n2057 VDD.n2056 3.1505
R2634 VDD.n2037 VDD.n2036 3.1505
R2635 VDD.n1599 VDD.n1598 3.1505
R2636 VDD.n60 VDD.n59 3.1505
R2637 VDD.n50 VDD.n49 3.1505
R2638 VDD.n48 VDD.n47 3.1505
R2639 VDD.n2166 VDD.n2165 3.1505
R2640 VDD.n2143 VDD.n2142 3.1505
R2641 VDD.n2147 VDD.n2145 3.1505
R2642 VDD.n2147 VDD.n2146 3.1505
R2643 VDD.n2122 VDD.n2121 3.1505
R2644 VDD.n2126 VDD.n2124 3.1505
R2645 VDD.n2126 VDD.n2125 3.1505
R2646 VDD.n2117 VDD.n2116 3.1505
R2647 VDD.n2102 VDD.n2100 3.1505
R2648 VDD.n2102 VDD.n2101 3.1505
R2649 VDD.n2095 VDD.n2094 3.1505
R2650 VDD.n2081 VDD.n2080 3.1505
R2651 VDD.n2059 VDD.n2058 3.1505
R2652 VDD.n2039 VDD.n2038 3.1505
R2653 VDD.n2035 VDD.n2034 3.1505
R2654 VDD.n1597 VDD.n1596 3.1505
R2655 VDD.n1930 VDD.n1929 3.1505
R2656 VDD.n1996 VDD.n1994 3.1505
R2657 VDD.n1996 VDD.n1995 3.1505
R2658 VDD.n2028 VDD.n1999 3.1505
R2659 VDD.n30 VDD.n29 3.1505
R2660 VDD.n27 VDD.n26 3.1505
R2661 VDD.n22 VDD.n21 3.1505
R2662 VDD.n24 VDD.n23 3.1505
R2663 VDD.n19 VDD.n18 3.1505
R2664 VDD.n16 VDD.n15 3.1505
R2665 VDD.n11 VDD.n10 3.1505
R2666 VDD.n13 VDD.n12 3.1505
R2667 VDD.n2149 VDD.n2148 3.1505
R2668 VDD.n2156 VDD.n2155 3.1505
R2669 VDD.n2151 VDD.n2150 3.1505
R2670 VDD.n2153 VDD.n2152 3.1505
R2671 VDD.n2129 VDD.n2128 3.1505
R2672 VDD.n2136 VDD.n2135 3.1505
R2673 VDD.n2133 VDD.n2132 3.1505
R2674 VDD.n2105 VDD.n2104 3.1505
R2675 VDD.n2131 VDD.n2130 3.1505
R2676 VDD.n2113 VDD.n2112 3.1505
R2677 VDD.n2110 VDD.n2109 3.1505
R2678 VDD.n2083 VDD.n2082 3.1505
R2679 VDD.n2108 VDD.n2107 3.1505
R2680 VDD.n2086 VDD.n2085 3.1505
R2681 VDD.n2065 VDD.n2064 3.1505
R2682 VDD.n2089 VDD.n2088 3.1505
R2683 VDD.n2091 VDD.n2090 3.1505
R2684 VDD.n2068 VDD.n2067 3.1505
R2685 VDD.n2072 VDD.n2071 3.1505
R2686 VDD.n2045 VDD.n2044 3.1505
R2687 VDD.n2070 VDD.n2069 3.1505
R2688 VDD.n2047 VDD.n2046 3.1505
R2689 VDD.n2053 VDD.n2052 3.1505
R2690 VDD.n1605 VDD.n1604 3.1505
R2691 VDD.n2049 VDD.n2048 3.1505
R2692 VDD.n2051 VDD.n2050 3.1505
R2693 VDD.n1611 VDD.n1610 3.1505
R2694 VDD.n1607 VDD.n1606 3.1505
R2695 VDD.n1609 VDD.n1608 3.1505
R2696 VDD.n1998 VDD.n1997 3.1505
R2697 VDD.n2023 VDD.n2022 3.1505
R2698 VDD.n2025 VDD.n2024 3.1505
R2699 VDD.n2027 VDD.n2026 3.1505
R2700 VDD.n2021 VDD.n2020 3.1505
R2701 VDD.n2030 VDD.n2029 3.1505
R2702 VDD.n43 VDD.n42 3.1505
R2703 VDD.n46 VDD.n45 3.1505
R2704 VDD.n45 VDD.n44 3.1505
R2705 VDD.n2209 VDD.n2208 3.1505
R2706 VDD.n2211 VDD.n2210 3.1505
R2707 VDD.n2215 VDD.n2214 3.1505
R2708 VDD.n2214 VDD.n2213 3.1505
R2709 VDD.n3115 VDD.n3114 3.1505
R2710 VDD.n3114 VDD.n3113 3.1505
R2711 VDD.n3112 VDD.n3111 3.1505
R2712 VDD.n3111 VDD.n3110 3.1505
R2713 VDD.n3108 VDD.n3107 3.1505
R2714 VDD.n2665 VDD.n2664 3.1505
R2715 VDD.n2630 VDD.n2629 3.1505
R2716 VDD.n2612 VDD.n2611 3.1505
R2717 VDD.n2606 VDD.n2605 3.1505
R2718 VDD.n2451 VDD.n2450 3.1505
R2719 VDD.n3074 VDD.n3073 3.1505
R2720 VDD.n3071 VDD.n3070 3.1505
R2721 VDD.n2375 VDD.n2374 3.1505
R2722 VDD.n2378 VDD.n2377 3.1505
R2723 VDD.n2385 VDD.n2384 3.1505
R2724 VDD.n2383 VDD.n2382 3.1505
R2725 VDD.n2380 VDD.n2379 3.1505
R2726 VDD.n2388 VDD.n2387 3.1505
R2727 VDD.n2395 VDD.n2394 3.1505
R2728 VDD.n2393 VDD.n2392 3.1505
R2729 VDD.n2390 VDD.n2389 3.1505
R2730 VDD.n2398 VDD.n2397 3.1505
R2731 VDD.n2405 VDD.n2404 3.1505
R2732 VDD.n2403 VDD.n2402 3.1505
R2733 VDD.n2400 VDD.n2399 3.1505
R2734 VDD.n2407 VDD.n2406 3.1505
R2735 VDD.n2415 VDD.n2414 3.1505
R2736 VDD.n2412 VDD.n2411 3.1505
R2737 VDD.n2409 VDD.n2408 3.1505
R2738 VDD.n2417 VDD.n2416 3.1505
R2739 VDD.n2425 VDD.n2424 3.1505
R2740 VDD.n2422 VDD.n2421 3.1505
R2741 VDD.n2419 VDD.n2418 3.1505
R2742 VDD.n2427 VDD.n2426 3.1505
R2743 VDD.n2442 VDD.n2441 3.1505
R2744 VDD.n2439 VDD.n2438 3.1505
R2745 VDD.n2436 VDD.n2435 3.1505
R2746 VDD.n2434 VDD.n2433 3.1505
R2747 VDD.n2431 VDD.n2430 3.1505
R2748 VDD.n2429 VDD.n2428 3.1505
R2749 VDD.n3077 VDD.n3076 3.1505
R2750 VDD.n2446 VDD.n2445 3.1505
R2751 VDD.n2444 VDD.n2443 3.1505
R2752 VDD.n2608 VDD.n2607 3.1505
R2753 VDD.n2610 VDD.n2609 3.1505
R2754 VDD.n2632 VDD.n2631 3.1505
R2755 VDD.n3100 VDD.n3099 3.1505
R2756 VDD.n2662 VDD.n2661 3.1505
R2757 VDD.n2017 VDD.n2016 3.1505
R2758 VDD.n2015 VDD.n2014 3.1505
R2759 VDD.n2013 VDD.n2012 3.1505
R2760 VDD.n2011 VDD.n2010 3.1505
R2761 VDD.n2009 VDD.n2008 3.1505
R2762 VDD.n2007 VDD.n2006 3.1505
R2763 VDD.n2005 VDD.n2004 3.1505
R2764 VDD.n2637 VDD.n2636 3.1505
R2765 VDD.n2639 VDD.n2638 3.1505
R2766 VDD.n2641 VDD.n2640 3.1505
R2767 VDD.n2643 VDD.n2642 3.1505
R2768 VDD.n2645 VDD.n2644 3.1505
R2769 VDD.n2648 VDD.n2647 3.1505
R2770 VDD.n2650 VDD.n2649 3.1505
R2771 VDD.n2652 VDD.n2651 3.1505
R2772 VDD.n2654 VDD.n2653 3.1505
R2773 VDD.n2656 VDD.n2655 3.1505
R2774 VDD.n2658 VDD.n2657 3.1505
R2775 VDD.n2660 VDD.n2659 3.1505
R2776 VDD.n2019 VDD.n2018 3.1505
R2777 VDD.n2173 VDD.n2172 3.1505
R2778 VDD.n2172 VDD.n2171 3.1505
R2779 VDD.n2176 VDD.n2175 3.1505
R2780 VDD.n2175 VDD.n2174 3.1505
R2781 VDD.n2179 VDD.n2178 3.1505
R2782 VDD.n2178 VDD.n2177 3.1505
R2783 VDD.n2182 VDD.n2181 3.1505
R2784 VDD.n2181 VDD.n2180 3.1505
R2785 VDD.n2185 VDD.n2184 3.1505
R2786 VDD.n2184 VDD.n2183 3.1505
R2787 VDD.n2188 VDD.n2187 3.1505
R2788 VDD.n2187 VDD.n2186 3.1505
R2789 VDD.n2192 VDD.n2191 3.1505
R2790 VDD.n2191 VDD.n2190 3.1505
R2791 VDD.n2195 VDD.n2194 3.1505
R2792 VDD.n2194 VDD.n2193 3.1505
R2793 VDD.n2198 VDD.n2197 3.1505
R2794 VDD.n2197 VDD.n2196 3.1505
R2795 VDD.n3130 VDD.n3129 3.1505
R2796 VDD.n3129 VDD.n3128 3.1505
R2797 VDD.n3127 VDD.n3126 3.1505
R2798 VDD.n3126 VDD.n3125 3.1505
R2799 VDD.n3123 VDD.n3122 3.1505
R2800 VDD.n3122 VDD.n3121 3.1505
R2801 VDD.n3120 VDD.n3119 3.1505
R2802 VDD.n3119 VDD.n3118 3.1505
R2803 VDD.n2472 VDD.t428 3.1255
R2804 VDD.n2316 VDD.t290 3.10434
R2805 VDD.n2598 VDD.n2595 2.84812
R2806 VDD.n1540 VDD.t15 2.62831
R2807 VDD.n564 VDD.t97 2.62831
R2808 VDD.n908 VDD.t147 2.62831
R2809 VDD.n391 VDD.n372 2.6005
R2810 VDD.n387 VDD.n374 2.6005
R2811 VDD.n385 VDD.n378 2.6005
R2812 VDD.n381 VDD.n380 2.6005
R2813 VDD.n436 VDD.n435 2.6005
R2814 VDD.n369 VDD.n362 2.6005
R2815 VDD.n368 VDD.n364 2.6005
R2816 VDD.n367 VDD.n366 2.6005
R2817 VDD.n667 VDD.n666 2.6005
R2818 VDD.n670 VDD.n669 2.6005
R2819 VDD.n360 VDD.n353 2.6005
R2820 VDD.n359 VDD.n355 2.6005
R2821 VDD.n358 VDD.n357 2.6005
R2822 VDD.n661 VDD.n660 2.6005
R2823 VDD.n664 VDD.n663 2.6005
R2824 VDD.n351 VDD.n344 2.6005
R2825 VDD.n350 VDD.n346 2.6005
R2826 VDD.n349 VDD.n348 2.6005
R2827 VDD.n655 VDD.n654 2.6005
R2828 VDD.n658 VDD.n657 2.6005
R2829 VDD.n342 VDD.n335 2.6005
R2830 VDD.n341 VDD.n337 2.6005
R2831 VDD.n340 VDD.n339 2.6005
R2832 VDD.n649 VDD.n648 2.6005
R2833 VDD.n652 VDD.n651 2.6005
R2834 VDD.n332 VDD.n324 2.6005
R2835 VDD.n330 VDD.n325 2.6005
R2836 VDD.n328 VDD.n326 2.6005
R2837 VDD.n643 VDD.n642 2.6005
R2838 VDD.n646 VDD.n645 2.6005
R2839 VDD.n264 VDD.n248 2.6005
R2840 VDD.n260 VDD.n250 2.6005
R2841 VDD.n258 VDD.n254 2.6005
R2842 VDD.n731 VDD.n730 2.6005
R2843 VDD.n735 VDD.n734 2.6005
R2844 VDD.n245 VDD.n238 2.6005
R2845 VDD.n244 VDD.n240 2.6005
R2846 VDD.n243 VDD.n242 2.6005
R2847 VDD.n1149 VDD.n1148 2.6005
R2848 VDD.n1152 VDD.n1151 2.6005
R2849 VDD.n236 VDD.n229 2.6005
R2850 VDD.n235 VDD.n231 2.6005
R2851 VDD.n234 VDD.n233 2.6005
R2852 VDD.n1164 VDD.n1163 2.6005
R2853 VDD.n1167 VDD.n1166 2.6005
R2854 VDD.n227 VDD.n220 2.6005
R2855 VDD.n226 VDD.n222 2.6005
R2856 VDD.n225 VDD.n224 2.6005
R2857 VDD.n1178 VDD.n1177 2.6005
R2858 VDD.n1181 VDD.n1180 2.6005
R2859 VDD.n218 VDD.n211 2.6005
R2860 VDD.n217 VDD.n213 2.6005
R2861 VDD.n216 VDD.n215 2.6005
R2862 VDD.n1143 VDD.n1142 2.6005
R2863 VDD.n1146 VDD.n1145 2.6005
R2864 VDD.n208 VDD.n200 2.6005
R2865 VDD.n206 VDD.n201 2.6005
R2866 VDD.n204 VDD.n202 2.6005
R2867 VDD.n1198 VDD.n1197 2.6005
R2868 VDD.n1201 VDD.n1200 2.6005
R2869 VDD.n111 VDD.n104 2.6005
R2870 VDD.n110 VDD.n106 2.6005
R2871 VDD.n109 VDD.n108 2.6005
R2872 VDD.n1944 VDD.n1943 2.6005
R2873 VDD.n1947 VDD.n1946 2.6005
R2874 VDD.n1004 VDD.n1000 2.6005
R2875 VDD.n1003 VDD.n1002 2.6005
R2876 VDD.n1038 VDD.n1032 2.6005
R2877 VDD.n1042 VDD.n1030 2.6005
R2878 VDD.n1328 VDD.n1322 2.6005
R2879 VDD.n1324 VDD.n1323 2.6005
R2880 VDD.n2978 VDD.n2977 2.6005
R2881 VDD.n2222 VDD.n2221 2.6005
R2882 VDD.n2223 VDD.n2219 2.6005
R2883 VDD.n2224 VDD.n2217 2.6005
R2884 VDD.n2933 VDD.n2932 2.6005
R2885 VDD.n2930 VDD.n2929 2.6005
R2886 VDD.n2339 VDD.n2338 2.6005
R2887 VDD.n2340 VDD.n2336 2.6005
R2888 VDD.n102 VDD.n95 2.6005
R2889 VDD.n101 VDD.n97 2.6005
R2890 VDD.n100 VDD.n99 2.6005
R2891 VDD.n1959 VDD.n1958 2.6005
R2892 VDD.n1962 VDD.n1961 2.6005
R2893 VDD.n93 VDD.n86 2.6005
R2894 VDD.n92 VDD.n88 2.6005
R2895 VDD.n91 VDD.n90 2.6005
R2896 VDD.n1938 VDD.n1937 2.6005
R2897 VDD.n1941 VDD.n1940 2.6005
R2898 VDD.n83 VDD.n75 2.6005
R2899 VDD.n81 VDD.n76 2.6005
R2900 VDD.n79 VDD.n77 2.6005
R2901 VDD.n1979 VDD.n1978 2.6005
R2902 VDD.n1982 VDD.n1981 2.6005
R2903 VDD.n139 VDD.n123 2.6005
R2904 VDD.n135 VDD.n125 2.6005
R2905 VDD.n133 VDD.n129 2.6005
R2906 VDD.n1335 VDD.n1334 2.6005
R2907 VDD.n1339 VDD.n1338 2.6005
R2908 VDD.n120 VDD.n113 2.6005
R2909 VDD.n119 VDD.n115 2.6005
R2910 VDD.n118 VDD.n117 2.6005
R2911 VDD.n1342 VDD.n1341 2.6005
R2912 VDD.n1345 VDD.n1344 2.6005
R2913 VDD.n2635 VDD.n2634 2.6005
R2914 VDD.n2205 VDD.n2204 2.6005
R2915 VDD.n2206 VDD.n2202 2.6005
R2916 VDD.n2207 VDD.n2200 2.6005
R2917 VDD.n2002 VDD.n2001 2.6005
R2918 VDD.n6 VDD.n5 2.6005
R2919 VDD.n7 VDD.n3 2.6005
R2920 VDD.n8 VDD.n1 2.6005
R2921 VDD.n1839 VDD.t342 2.48683
R2922 VDD.n2626 VDD.n2625 2.40832
R2923 VDD.n2623 VDD.n2622 2.40832
R2924 VDD.n631 VDD.n630 2.40832
R2925 VDD.n502 VDD.n501 2.40832
R2926 VDD.n499 VDD.n498 2.40832
R2927 VDD.n496 VDD.n495 2.40832
R2928 VDD.n493 VDD.n492 2.40832
R2929 VDD.n490 VDD.n489 2.40832
R2930 VDD.n487 VDD.n486 2.40832
R2931 VDD.n512 VDD.n511 2.40832
R2932 VDD.n521 VDD.n520 2.40832
R2933 VDD.n412 VDD.n411 2.40832
R2934 VDD.n409 VDD.n408 2.40832
R2935 VDD.n2705 VDD.t439 2.15196
R2936 VDD.n1573 VDD.t18 2.15052
R2937 VDD.n597 VDD.t59 2.15052
R2938 VDD.n941 VDD.t50 2.15052
R2939 VDD.n2206 VDD.n2205 2.03528
R2940 VDD.n7 VDD.n6 2.03528
R2941 VDD.n2207 VDD.n2206 2.03137
R2942 VDD.n8 VDD.n7 2.03137
R2943 VDD.n2351 VDD.t435 1.97567
R2944 VDD.n1040 VDD.n1039 1.96766
R2945 VDD.n1326 VDD.n1325 1.96766
R2946 VDD.n533 VDD.n531 1.93067
R2947 VDD.n2085 VDD.n2084 1.79846
R2948 VDD.n2067 VDD.n2066 1.79846
R2949 VDD.n2441 VDD.n2440 1.79846
R2950 VDD.n2433 VDD.n2432 1.79846
R2951 VDD.n2107 VDD.n2106 1.75914
R2952 VDD.n2438 VDD.n2437 1.75914
R2953 VDD.n3076 VDD.n3075 1.75914
R2954 VDD.n1064 VDD.n1061 1.74343
R2955 VDD.n994 VDD.n991 1.74343
R2956 VDD.n1013 VDD.n1010 1.74343
R2957 VDD.n1321 VDD.n1318 1.74343
R2958 VDD.n1123 VDD.n1122 1.74343
R2959 VDD.n2964 VDD.n2962 1.74343
R2960 VDD.n1849 VDD.n1846 1.74343
R2961 VDD.n1819 VDD.n1816 1.74343
R2962 VDD.n635 VDD.n633 1.74343
R2963 VDD.n752 VDD.n750 1.74343
R2964 VDD.n479 VDD.n477 1.74343
R2965 VDD.n1442 VDD.n1440 1.74343
R2966 VDD.n154 VDD.n152 1.74343
R2967 VDD.n1370 VDD.n1368 1.74343
R2968 VDD.n1950 VDD.n1948 1.74343
R2969 VDD.n1223 VDD.n1221 1.74343
R2970 VDD.n2212 VDD.n2209 1.74343
R2971 VDD.n1321 VDD.n1320 1.7429
R2972 VDD.n1013 VDD.n1012 1.7429
R2973 VDD.n994 VDD.n993 1.7429
R2974 VDD.n1064 VDD.n1063 1.7429
R2975 VDD.n2964 VDD.n2963 1.7429
R2976 VDD.n1849 VDD.n1848 1.7429
R2977 VDD.n1819 VDD.n1818 1.7429
R2978 VDD.n752 VDD.n751 1.7429
R2979 VDD.n1455 VDD.n1454 1.7429
R2980 VDD.n159 VDD.n158 1.7429
R2981 VDD.n1370 VDD.n1369 1.7429
R2982 VDD.n1223 VDD.n1222 1.7429
R2983 VDD.n1950 VDD.n1949 1.7429
R2984 VDD.n2212 VDD.n2211 1.7429
R2985 VDD.n26 VDD.n25 1.74276
R2986 VDD.n21 VDD.n20 1.74276
R2987 VDD.n15 VDD.n14 1.74276
R2988 VDD.n10 VDD.n9 1.74276
R2989 VDD.n2155 VDD.n2154 1.74276
R2990 VDD.n2135 VDD.n2134 1.74276
R2991 VDD.n2112 VDD.n2111 1.74276
R2992 VDD.n2088 VDD.n2087 1.74276
R2993 VDD.n1116 VDD.n1115 1.74276
R2994 VDD.n1111 VDD.n1110 1.74276
R2995 VDD.n1106 VDD.n1105 1.74276
R2996 VDD.n1101 VDD.n1100 1.74276
R2997 VDD.n1096 VDD.n1095 1.74276
R2998 VDD.n1091 VDD.n1090 1.74276
R2999 VDD.n1086 VDD.n1085 1.74276
R3000 VDD.n1229 VDD.n1228 1.74276
R3001 VDD.n1269 VDD.n1268 1.74276
R3002 VDD.n1274 VDD.n1273 1.74276
R3003 VDD.n2586 VDD.n2585 1.74276
R3004 VDD.n2581 VDD.n2580 1.74276
R3005 VDD.n2576 VDD.n2575 1.74276
R3006 VDD.n2571 VDD.n2570 1.74276
R3007 VDD.n2566 VDD.n2565 1.74276
R3008 VDD.n2561 VDD.n2560 1.74276
R3009 VDD.n2556 VDD.n2555 1.74276
R3010 VDD.n2736 VDD.n2735 1.74276
R3011 VDD.n2817 VDD.n2816 1.74276
R3012 VDD.n2899 VDD.n2898 1.74276
R3013 VDD.n2670 VDD.n2669 1.74276
R3014 VDD.n2675 VDD.n2674 1.74276
R3015 VDD.n2680 VDD.n2679 1.74276
R3016 VDD.n2685 VDD.n2684 1.74276
R3017 VDD.n2744 VDD.n2743 1.74276
R3018 VDD.n2739 VDD.n2738 1.74276
R3019 VDD.n2766 VDD.n2765 1.74276
R3020 VDD.n2761 VDD.n2760 1.74276
R3021 VDD.n2780 VDD.n2779 1.74276
R3022 VDD.n2785 VDD.n2784 1.74276
R3023 VDD.n2799 VDD.n2798 1.74276
R3024 VDD.n2804 VDD.n2803 1.74276
R3025 VDD.n2814 VDD.n2813 1.74276
R3026 VDD.n2462 VDD.n2459 1.74276
R3027 VDD.n2476 VDD.n2473 1.74276
R3028 VDD.n2488 VDD.n2485 1.74276
R3029 VDD.n2500 VDD.n2497 1.74276
R3030 VDD.n2500 VDD.n2499 1.74276
R3031 VDD.n2488 VDD.n2487 1.74276
R3032 VDD.n2476 VDD.n2475 1.74276
R3033 VDD.n2462 VDD.n2461 1.74276
R3034 VDD.n3079 VDD.n3078 1.74276
R3035 VDD.n3084 VDD.n3083 1.74276
R3036 VDD.n3096 VDD.n3095 1.74276
R3037 VDD.n3066 VDD.n3065 1.74276
R3038 VDD.n3048 VDD.n3047 1.74276
R3039 VDD.n3035 VDD.n3034 1.74276
R3040 VDD.n3023 VDD.n3022 1.74276
R3041 VDD.n3006 VDD.n3005 1.74276
R3042 VDD.n2926 VDD.n2925 1.74276
R3043 VDD.n3014 VDD.n3013 1.74276
R3044 VDD.n3019 VDD.n3018 1.74276
R3045 VDD.n3026 VDD.n3025 1.74276
R3046 VDD.n3031 VDD.n3030 1.74276
R3047 VDD.n3042 VDD.n3041 1.74276
R3048 VDD.n3055 VDD.n3054 1.74276
R3049 VDD.n3063 VDD.n3062 1.74276
R3050 VDD.n3091 VDD.n3090 1.74276
R3051 VDD.n2277 VDD.n2276 1.74276
R3052 VDD.n2272 VDD.n2271 1.74276
R3053 VDD.n2267 VDD.n2266 1.74276
R3054 VDD.n2262 VDD.n2261 1.74276
R3055 VDD.n2257 VDD.n2256 1.74276
R3056 VDD.n2252 VDD.n2251 1.74276
R3057 VDD.n2999 VDD.n2997 1.74276
R3058 VDD.n2990 VDD.n2988 1.74276
R3059 VDD.n2936 VDD.n2934 1.74276
R3060 VDD.n2972 VDD.n2970 1.74276
R3061 VDD.n2999 VDD.n2998 1.74276
R3062 VDD.n2990 VDD.n2989 1.74276
R3063 VDD.n2936 VDD.n2935 1.74276
R3064 VDD.n2972 VDD.n2971 1.74276
R3065 VDD.n2912 VDD.n2911 1.74276
R3066 VDD.n1673 VDD.n1669 1.74276
R3067 VDD.n1667 VDD.n1666 1.74276
R3068 VDD.n1658 VDD.n1657 1.74276
R3069 VDD.n1661 VDD.n1660 1.74276
R3070 VDD.n1776 VDD.n1775 1.74276
R3071 VDD.n1902 VDD.n1901 1.74276
R3072 VDD.n1899 VDD.n1898 1.74276
R3073 VDD.n1893 VDD.n1892 1.74276
R3074 VDD.n1890 VDD.n1889 1.74276
R3075 VDD.n1841 VDD.n1838 1.74276
R3076 VDD.n1827 VDD.n1824 1.74276
R3077 VDD.n1794 VDD.n1791 1.74276
R3078 VDD.n1841 VDD.n1840 1.74276
R3079 VDD.n1827 VDD.n1826 1.74276
R3080 VDD.n1794 VDD.n1793 1.74276
R3081 VDD.n1489 VDD.n1487 1.74276
R3082 VDD.n1471 VDD.n1470 1.74276
R3083 VDD.n1452 VDD.n1451 1.74276
R3084 VDD.n1485 VDD.n1484 1.74276
R3085 VDD.n1467 VDD.n1466 1.74276
R3086 VDD.n1448 VDD.n1447 1.74276
R3087 VDD.n1170 VDD.n1168 1.74276
R3088 VDD.n1184 VDD.n1182 1.74276
R3089 VDD.n1193 VDD.n1191 1.74276
R3090 VDD.n1193 VDD.n1192 1.74276
R3091 VDD.n1184 VDD.n1183 1.74276
R3092 VDD.n1170 VDD.n1169 1.74276
R3093 VDD.n297 VDD.n296 1.74276
R3094 VDD.n872 VDD.n871 1.74276
R3095 VDD.n859 VDD.n858 1.74276
R3096 VDD.n856 VDD.n855 1.74276
R3097 VDD.n839 VDD.n838 1.74276
R3098 VDD.n836 VDD.n835 1.74276
R3099 VDD.n818 VDD.n817 1.74276
R3100 VDD.n815 VDD.n814 1.74276
R3101 VDD.n719 VDD.n717 1.74276
R3102 VDD.n719 VDD.n718 1.74276
R3103 VDD.n876 VDD.n875 1.74276
R3104 VDD.n428 VDD.n427 1.74276
R3105 VDD.n1965 VDD.n1963 1.74276
R3106 VDD.n1974 VDD.n1972 1.74276
R3107 VDD.n1974 VDD.n1973 1.74276
R3108 VDD.n1965 VDD.n1964 1.74276
R3109 VDD.n2160 VDD.n2159 1.74276
R3110 VDD.n2145 VDD.n2144 1.74276
R3111 VDD.n2140 VDD.n2139 1.74276
R3112 VDD.n2124 VDD.n2123 1.74276
R3113 VDD.n2119 VDD.n2118 1.74276
R3114 VDD.n2100 VDD.n2099 1.74276
R3115 VDD.n2097 VDD.n2096 1.74276
R3116 VDD.n2104 VDD.n2103 1.74276
R3117 VDD.n2128 VDD.n2127 1.74276
R3118 VDD.n2414 VDD.n2413 1.74276
R3119 VDD.n2424 VDD.n2423 1.74276
R3120 VDD.n3070 VDD.n3069 1.74276
R3121 VDD.n2377 VDD.n2376 1.74276
R3122 VDD.n2382 VDD.n2381 1.74276
R3123 VDD.n2387 VDD.n2386 1.74276
R3124 VDD.n2392 VDD.n2391 1.74276
R3125 VDD.n2397 VDD.n2396 1.74276
R3126 VDD.n2402 VDD.n2401 1.74276
R3127 VDD.n2411 VDD.n2410 1.74276
R3128 VDD.n2421 VDD.n2420 1.74276
R3129 VDD.n534 VDD.n533 1.7105
R3130 VDD.n2478 VDD.t442 1.563
R3131 VDD.n1918 VDD.t371 1.4923
R3132 VDD.n2728 VDD.n2727 1.441
R3133 VDD.n2618 VDD.n2617 1.42472
R3134 VDD.n2593 VDD.n2592 1.42472
R3135 VDD.n415 VDD.n414 1.42472
R3136 VDD.n1278 VDD.n1277 1.42456
R3137 VDD.n2667 VDD.n2666 1.42456
R3138 VDD.n2598 VDD.n2597 1.42456
R3139 VDD.n1911 VDD.n1910 1.42456
R3140 VDD.n1906 VDD.n1905 1.42456
R3141 VDD.n284 VDD.n283 1.42456
R3142 VDD.n822 VDD.n821 1.42456
R3143 VDD.n765 VDD.n764 1.42456
R3144 VDD.n722 VDD.n721 1.42456
R3145 VDD.n404 VDD.n403 1.42456
R3146 VDD.n516 VDD.n515 1.42456
R3147 VDD.n482 VDD.n481 1.42456
R3148 VDD.n463 VDD.n462 1.42456
R3149 VDD.n42 VDD.n41 1.36443
R3150 VDD.n3107 VDD.n3106 1.36443
R3151 VDD.n2664 VDD.n2663 1.36443
R3152 VDD.n2516 VDD.n2515 1.351
R3153 VDD.n2295 VDD.n2294 1.351
R3154 VDD.n2821 VDD.n2820 1.351
R3155 VDD.n2193 VDD.t266 1.34158
R3156 VDD.n2224 VDD.n2223 1.27435
R3157 VDD.n2223 VDD.n2222 1.27435
R3158 VDD.n2340 VDD.n2339 1.27435
R3159 VDD.n2933 VDD.n2930 1.27435
R3160 VDD.n2617 VDD.n2616 1.15215
R3161 VDD.n2599 VDD.n2593 1.15215
R3162 VDD.n2599 VDD.n2598 1.15196
R3163 VDD.n2646 VDD.n2635 1.1255
R3164 VDD.n2003 VDD.n2002 1.1255
R3165 VDD.n369 VDD.n368 1.0864
R3166 VDD.n368 VDD.n367 1.0864
R3167 VDD.n670 VDD.n667 1.0864
R3168 VDD.n360 VDD.n359 1.0864
R3169 VDD.n359 VDD.n358 1.0864
R3170 VDD.n664 VDD.n661 1.0864
R3171 VDD.n351 VDD.n350 1.0864
R3172 VDD.n350 VDD.n349 1.0864
R3173 VDD.n658 VDD.n655 1.0864
R3174 VDD.n342 VDD.n341 1.0864
R3175 VDD.n341 VDD.n340 1.0864
R3176 VDD.n652 VDD.n649 1.0864
R3177 VDD.n245 VDD.n244 1.0864
R3178 VDD.n244 VDD.n243 1.0864
R3179 VDD.n1152 VDD.n1149 1.0864
R3180 VDD.n236 VDD.n235 1.0864
R3181 VDD.n235 VDD.n234 1.0864
R3182 VDD.n1167 VDD.n1164 1.0864
R3183 VDD.n227 VDD.n226 1.0864
R3184 VDD.n226 VDD.n225 1.0864
R3185 VDD.n1181 VDD.n1178 1.0864
R3186 VDD.n218 VDD.n217 1.0864
R3187 VDD.n217 VDD.n216 1.0864
R3188 VDD.n1146 VDD.n1143 1.0864
R3189 VDD.n111 VDD.n110 1.0864
R3190 VDD.n110 VDD.n109 1.0864
R3191 VDD.n1947 VDD.n1944 1.0864
R3192 VDD.n102 VDD.n101 1.0864
R3193 VDD.n101 VDD.n100 1.0864
R3194 VDD.n1962 VDD.n1959 1.0864
R3195 VDD.n93 VDD.n92 1.0864
R3196 VDD.n92 VDD.n91 1.0864
R3197 VDD.n1941 VDD.n1938 1.0864
R3198 VDD.n120 VDD.n119 1.0864
R3199 VDD.n119 VDD.n118 1.0864
R3200 VDD.n1345 VDD.n1342 1.0864
R3201 VDD.n2721 VDD.n2720 1.07528
R3202 VDD.n424 VDD.n423 1.04661
R3203 VDD.n2591 VDD.t301 1.04217
R3204 VDD.n3124 VDD.n2207 1.03159
R3205 VDD.n2189 VDD.n8 1.03159
R3206 VDD.n2979 VDD.n2978 0.968
R3207 VDD.n2985 VDD.n2933 0.968
R3208 VDD.n1795 VDD.t4 0.9105
R3209 VDD.n1795 VDD.t348 0.9105
R3210 VDD.n1829 VDD.t457 0.9105
R3211 VDD.n1829 VDD.n1828 0.9105
R3212 VDD.n1843 VDD.t372 0.9105
R3213 VDD.n1843 VDD.n1842 0.9105
R3214 VDD.n1002 VDD.t448 0.9105
R3215 VDD.n1002 VDD.n1001 0.9105
R3216 VDD.n1000 VDD.t9 0.9105
R3217 VDD.n1000 VDD.n999 0.9105
R3218 VDD.n1323 VDD.t285 0.9105
R3219 VDD.n1323 VDD.t354 0.9105
R3220 VDD.n1322 VDD.t467 0.9105
R3221 VDD.n1322 VDD.t419 0.9105
R3222 VDD.n1030 VDD.t376 0.9105
R3223 VDD.n1030 VDD.n1029 0.9105
R3224 VDD.n1032 VDD.t337 0.9105
R3225 VDD.n1032 VDD.n1031 0.9105
R3226 VDD.n1855 VDD.n1854 0.9105
R3227 VDD.n1705 VDD.t6 0.9105
R3228 VDD.n1705 VDD.n1704 0.9105
R3229 VDD.n1703 VDD.t423 0.9105
R3230 VDD.n1821 VDD.t302 0.9105
R3231 VDD.n1821 VDD.n1820 0.9105
R3232 VDD.n2515 VDD.n2514 0.901
R3233 VDD.n2294 VDD.n2293 0.901
R3234 VDD.n2322 VDD.n2224 0.9005
R3235 VDD.n2341 VDD.n2340 0.9005
R3236 VDD.n41 VDD.n40 0.894284
R3237 VDD.n3106 VDD.n3105 0.894284
R3238 VDD.n40 VDD.n37 0.894284
R3239 VDD.n1786 VDD.n1613 0.843086
R3240 VDD.n1914 VDD.n1844 0.843086
R3241 VDD.n421 VDD.n417 0.794848
R3242 VDD.n563 VDD.n369 0.788369
R3243 VDD.n573 VDD.n360 0.788369
R3244 VDD.n583 VDD.n351 0.788369
R3245 VDD.n596 VDD.n342 0.788369
R3246 VDD.n907 VDD.n245 0.788369
R3247 VDD.n917 VDD.n236 0.788369
R3248 VDD.n927 VDD.n227 0.788369
R3249 VDD.n940 VDD.n218 0.788369
R3250 VDD.n1549 VDD.n111 0.788369
R3251 VDD.n1559 VDD.n102 0.788369
R3252 VDD.n1572 VDD.n93 0.788369
R3253 VDD.n1539 VDD.n120 0.788369
R3254 VDD.n1004 VDD.n1003 0.75425
R3255 VDD.n982 VDD.n981 0.75425
R3256 VDD.n1952 VDD.n1947 0.715603
R3257 VDD.n1171 VDD.n1167 0.710091
R3258 VDD.n1185 VDD.n1181 0.710091
R3259 VDD.n1966 VDD.n1962 0.710091
R3260 VDD.n1363 VDD.n1220 0.710091
R3261 VDD.n1329 VDD.n1321 0.705355
R3262 VDD.n1014 VDD.n1013 0.705355
R3263 VDD.n995 VDD.n994 0.705355
R3264 VDD.n1127 VDD.n1064 0.705355
R3265 VDD.n1122 VDD.n1121 0.705355
R3266 VDD.n1293 VDD.n1292 0.705355
R3267 VDD.n2757 VDD.n2754 0.705355
R3268 VDD.n2753 VDD.n2752 0.705355
R3269 VDD.n2965 VDD.n2964 0.705355
R3270 VDD.n2914 VDD.n2908 0.705355
R3271 VDD.n1672 VDD.n1671 0.705355
R3272 VDD.n1744 VDD.n1743 0.705355
R3273 VDD.n1752 VDD.n1751 0.705355
R3274 VDD.n1760 VDD.n1759 0.705355
R3275 VDD.n1886 VDD.n1884 0.705355
R3276 VDD.n1913 VDD.n1849 0.705355
R3277 VDD.n1822 VDD.n1819 0.705355
R3278 VDD.n1435 VDD.n1434 0.705355
R3279 VDD.n1416 VDD.n1415 0.705355
R3280 VDD.n1397 VDD.n1396 0.705355
R3281 VDD.n1380 VDD.n1379 0.705355
R3282 VDD.n772 VDD.n771 0.705355
R3283 VDD.n793 VDD.n792 0.705355
R3284 VDD.n810 VDD.n809 0.705355
R3285 VDD.n829 VDD.n828 0.705355
R3286 VDD.n851 VDD.n850 0.705355
R3287 VDD.n636 VDD.n635 0.705355
R3288 VDD.n753 VDD.n752 0.705355
R3289 VDD.n802 VDD.n801 0.705355
R3290 VDD.n783 VDD.n782 0.705355
R3291 VDD.n763 VDD.n762 0.705355
R3292 VDD.n627 VDD.n626 0.705355
R3293 VDD.n461 VDD.n459 0.705355
R3294 VDD.n472 VDD.n471 0.705355
R3295 VDD.n480 VDD.n479 0.705355
R3296 VDD.n513 VDD.n510 0.705355
R3297 VDD.n513 VDD.n507 0.705355
R3298 VDD.n524 VDD.n523 0.705355
R3299 VDD.n529 VDD.n526 0.705355
R3300 VDD.n529 VDD.n528 0.705355
R3301 VDD.n307 VDD.n306 0.705355
R3302 VDD.n293 VDD.n292 0.705355
R3303 VDD.n290 VDD.n289 0.705355
R3304 VDD.n183 VDD.n182 0.705355
R3305 VDD.n155 VDD.n154 0.705355
R3306 VDD.n1500 VDD.n1499 0.705355
R3307 VDD.n1480 VDD.n1479 0.705355
R3308 VDD.n1462 VDD.n1461 0.705355
R3309 VDD.n1443 VDD.n1442 0.705355
R3310 VDD.n1426 VDD.n1425 0.705355
R3311 VDD.n1405 VDD.n1404 0.705355
R3312 VDD.n1388 VDD.n1387 0.705355
R3313 VDD.n165 VDD.n164 0.705355
R3314 VDD.n1371 VDD.n1370 0.705355
R3315 VDD.n166 VDD.n165 0.705355
R3316 VDD.n1363 VDD.n1223 0.705355
R3317 VDD.n1952 VDD.n1950 0.705355
R3318 VDD.n2166 VDD.n2164 0.705355
R3319 VDD.n2063 VDD.n2062 0.705355
R3320 VDD.n2043 VDD.n2042 0.705355
R3321 VDD.n1603 VDD.n1602 0.705355
R3322 VDD.n2215 VDD.n2212 0.705355
R3323 VDD.n2451 VDD.n2449 0.705355
R3324 VDD.n1285 VDD.n1284 0.705118
R3325 VDD.n1295 VDD.n1294 0.705118
R3326 VDD.n2797 VDD.n2792 0.705118
R3327 VDD.n2776 VDD.n2771 0.705118
R3328 VDD.n2514 VDD.n2513 0.705118
R3329 VDD.n2514 VDD.n2512 0.705118
R3330 VDD.n2514 VDD.n2511 0.705118
R3331 VDD.n2514 VDD.n2510 0.705118
R3332 VDD.n2514 VDD.n2509 0.705118
R3333 VDD.n2514 VDD.n2508 0.705118
R3334 VDD.n2514 VDD.n2507 0.705118
R3335 VDD.n2514 VDD.n2506 0.705118
R3336 VDD.n2514 VDD.n2505 0.705118
R3337 VDD.n2514 VDD.n2504 0.705118
R3338 VDD.n2514 VDD.n2503 0.705118
R3339 VDD.n2501 VDD.n2500 0.705118
R3340 VDD.n2489 VDD.n2488 0.705118
R3341 VDD.n2477 VDD.n2476 0.705118
R3342 VDD.n2465 VDD.n2462 0.705118
R3343 VDD.n3095 VDD.n3094 0.705118
R3344 VDD.n2293 VDD.n2292 0.705118
R3345 VDD.n2293 VDD.n2291 0.705118
R3346 VDD.n2293 VDD.n2290 0.705118
R3347 VDD.n2293 VDD.n2289 0.705118
R3348 VDD.n2293 VDD.n2288 0.705118
R3349 VDD.n2293 VDD.n2287 0.705118
R3350 VDD.n2293 VDD.n2286 0.705118
R3351 VDD.n2293 VDD.n2285 0.705118
R3352 VDD.n2293 VDD.n2284 0.705118
R3353 VDD.n2293 VDD.n2283 0.705118
R3354 VDD.n2293 VDD.n2282 0.705118
R3355 VDD.n3000 VDD.n2999 0.705118
R3356 VDD.n2992 VDD.n2990 0.705118
R3357 VDD.n2982 VDD.n2936 0.705118
R3358 VDD.n2973 VDD.n2972 0.705118
R3359 VDD.n1701 VDD.n1673 0.705118
R3360 VDD.n1654 VDD.n1616 0.705118
R3361 VDD.n1649 VDD.n1620 0.705118
R3362 VDD.n1644 VDD.n1623 0.705118
R3363 VDD.n1768 VDD.n1767 0.705118
R3364 VDD.n1770 VDD.n1769 0.705118
R3365 VDD.n1876 VDD.n1852 0.705118
R3366 VDD.n1883 VDD.n1882 0.705118
R3367 VDD.n1921 VDD.n1841 0.705118
R3368 VDD.n1836 VDD.n1827 0.705118
R3369 VDD.n1805 VDD.n1794 0.705118
R3370 VDD.n1509 VDD.n1506 0.705118
R3371 VDD.n1492 VDD.n1489 0.705118
R3372 VDD.n179 VDD.n178 0.705118
R3373 VDD.n179 VDD.n177 0.705118
R3374 VDD.n180 VDD.n179 0.705118
R3375 VDD.n1194 VDD.n1193 0.705118
R3376 VDD.n1185 VDD.n1184 0.705118
R3377 VDD.n1171 VDD.n1170 0.705118
R3378 VDD.n280 VDD.n279 0.705118
R3379 VDD.n867 VDD.n866 0.705118
R3380 VDD.n720 VDD.n719 0.705118
R3381 VDD.n304 VDD.n303 0.705118
R3382 VDD.n451 VDD.n428 0.705118
R3383 VDD.n305 VDD.n304 0.705118
R3384 VDD.n169 VDD.n168 0.705118
R3385 VDD.n1975 VDD.n1974 0.705118
R3386 VDD.n1966 VDD.n1965 0.705118
R3387 VDD.n58 VDD.n57 0.705118
R3388 VDD.n2081 VDD.n2079 0.705118
R3389 VDD.n55 VDD.n54 0.705118
R3390 VDD.n54 VDD.n53 0.705118
R3391 VDD.n54 VDD.n52 0.705118
R3392 VDD.n40 VDD.n33 0.705118
R3393 VDD.n40 VDD.n39 0.705118
R3394 VDD.n40 VDD.n38 0.705118
R3395 VDD.n3105 VDD.n3102 0.705118
R3396 VDD.n40 VDD.n35 0.69693
R3397 VDD.n40 VDD.n31 0.69693
R3398 VDD.n3105 VDD.n3104 0.69693
R3399 VDD.n1038 VDD.n1037 0.690969
R3400 VDD.n981 VDD.n980 0.690969
R3401 VDD.n446 VDD.n432 0.688041
R3402 VDD.n441 VDD.n436 0.688041
R3403 VDD.n675 VDD.n670 0.688041
R3404 VDD.n682 VDD.n664 0.688041
R3405 VDD.n689 VDD.n658 0.688041
R3406 VDD.n698 VDD.n652 0.688041
R3407 VDD.n705 VDD.n646 0.688041
R3408 VDD.n710 VDD.n641 0.688041
R3409 VDD.n745 VDD.n728 0.688041
R3410 VDD.n740 VDD.n735 0.688041
R3411 VDD.n1157 VDD.n1152 0.688041
R3412 VDD.n1190 VDD.n1146 0.688041
R3413 VDD.n1202 VDD.n1201 0.688041
R3414 VDD.n1207 VDD.n1140 0.688041
R3415 VDD.n1971 VDD.n1941 0.688041
R3416 VDD.n1983 VDD.n1982 0.688041
R3417 VDD.n1988 VDD.n1935 0.688041
R3418 VDD.n1360 VDD.n1339 0.688041
R3419 VDD.n1350 VDD.n1345 0.688041
R3420 VDD.n1127 VDD.n1070 0.687706
R3421 VDD.n1329 VDD.n1328 0.687706
R3422 VDD.n40 VDD.n36 0.677271
R3423 VDD.n40 VDD.n34 0.677271
R3424 VDD.n40 VDD.n32 0.677271
R3425 VDD.n3105 VDD.n3103 0.677271
R3426 VDD.n3105 VDD.n3101 0.677271
R3427 VDD.n1005 VDD.n1004 0.665656
R3428 VDD.n1049 VDD.n1042 0.665656
R3429 VDD.n983 VDD.n982 0.665656
R3430 VDD.n1310 VDD.n1309 0.665656
R3431 VDD.n1 VDD.t433 0.607167
R3432 VDD.n1 VDD.n0 0.607167
R3433 VDD.n3 VDD.t330 0.607167
R3434 VDD.n3 VDD.n2 0.607167
R3435 VDD.n5 VDD.t470 0.607167
R3436 VDD.n5 VDD.n4 0.607167
R3437 VDD.n2001 VDD.t2 0.607167
R3438 VDD.n2001 VDD.n2000 0.607167
R3439 VDD.n435 VDD.n434 0.607167
R3440 VDD.n380 VDD.t401 0.607167
R3441 VDD.n380 VDD.n379 0.607167
R3442 VDD.n378 VDD.t397 0.607167
R3443 VDD.n378 VDD.n377 0.607167
R3444 VDD.n374 VDD.t409 0.607167
R3445 VDD.n374 VDD.n373 0.607167
R3446 VDD.n372 VDD.t386 0.607167
R3447 VDD.n372 VDD.n371 0.607167
R3448 VDD.n669 VDD.t208 0.607167
R3449 VDD.n669 VDD.n668 0.607167
R3450 VDD.n666 VDD.t30 0.607167
R3451 VDD.n666 VDD.n665 0.607167
R3452 VDD.n366 VDD.t262 0.607167
R3453 VDD.n366 VDD.n365 0.607167
R3454 VDD.n364 VDD.t167 0.607167
R3455 VDD.n364 VDD.n363 0.607167
R3456 VDD.n362 VDD.t117 0.607167
R3457 VDD.n362 VDD.n361 0.607167
R3458 VDD.n663 VDD.t256 0.607167
R3459 VDD.n663 VDD.n662 0.607167
R3460 VDD.n660 VDD.t107 0.607167
R3461 VDD.n660 VDD.n659 0.607167
R3462 VDD.n357 VDD.t94 0.607167
R3463 VDD.n357 VDD.n356 0.607167
R3464 VDD.n355 VDD.t83 0.607167
R3465 VDD.n355 VDD.n354 0.607167
R3466 VDD.n353 VDD.t239 0.607167
R3467 VDD.n353 VDD.n352 0.607167
R3468 VDD.n657 VDD.t90 0.607167
R3469 VDD.n657 VDD.n656 0.607167
R3470 VDD.n654 VDD.t161 0.607167
R3471 VDD.n654 VDD.n653 0.607167
R3472 VDD.n348 VDD.t152 0.607167
R3473 VDD.n348 VDD.n347 0.607167
R3474 VDD.n346 VDD.t234 0.607167
R3475 VDD.n346 VDD.n345 0.607167
R3476 VDD.n344 VDD.t157 0.607167
R3477 VDD.n344 VDD.n343 0.607167
R3478 VDD.n651 VDD.t200 0.607167
R3479 VDD.n651 VDD.n650 0.607167
R3480 VDD.n648 VDD.t257 0.607167
R3481 VDD.n648 VDD.n647 0.607167
R3482 VDD.n339 VDD.t254 0.607167
R3483 VDD.n339 VDD.n338 0.607167
R3484 VDD.n337 VDD.t186 0.607167
R3485 VDD.n337 VDD.n336 0.607167
R3486 VDD.n335 VDD.t44 0.607167
R3487 VDD.n335 VDD.n334 0.607167
R3488 VDD.n645 VDD.t249 0.607167
R3489 VDD.n642 VDD.t93 0.607167
R3490 VDD.n326 VDD.t77 0.607167
R3491 VDD.n325 VDD.t118 0.607167
R3492 VDD.n324 VDD.t199 0.607167
R3493 VDD.n1200 VDD.t27 0.607167
R3494 VDD.n734 VDD.n733 0.607167
R3495 VDD.n730 VDD.n729 0.607167
R3496 VDD.n254 VDD.t417 0.607167
R3497 VDD.n254 VDD.n253 0.607167
R3498 VDD.n250 VDD.t390 0.607167
R3499 VDD.n250 VDD.n249 0.607167
R3500 VDD.n248 VDD.t403 0.607167
R3501 VDD.n248 VDD.n247 0.607167
R3502 VDD.n1151 VDD.t230 0.607167
R3503 VDD.n1151 VDD.n1150 0.607167
R3504 VDD.n1148 VDD.t64 0.607167
R3505 VDD.n1148 VDD.n1147 0.607167
R3506 VDD.n242 VDD.t49 0.607167
R3507 VDD.n242 VDD.n241 0.607167
R3508 VDD.n240 VDD.t209 0.607167
R3509 VDD.n240 VDD.n239 0.607167
R3510 VDD.n238 VDD.t73 0.607167
R3511 VDD.n238 VDD.n237 0.607167
R3512 VDD.n1166 VDD.t46 0.607167
R3513 VDD.n1166 VDD.n1165 0.607167
R3514 VDD.n1163 VDD.t134 0.607167
R3515 VDD.n1163 VDD.n1162 0.607167
R3516 VDD.n233 VDD.t127 0.607167
R3517 VDD.n233 VDD.n232 0.607167
R3518 VDD.n231 VDD.t138 0.607167
R3519 VDD.n231 VDD.n230 0.607167
R3520 VDD.n229 VDD.t213 0.607167
R3521 VDD.n229 VDD.n228 0.607167
R3522 VDD.n1180 VDD.t122 0.607167
R3523 VDD.n1180 VDD.n1179 0.607167
R3524 VDD.n1177 VDD.t188 0.607167
R3525 VDD.n1177 VDD.n1176 0.607167
R3526 VDD.n224 VDD.t176 0.607167
R3527 VDD.n224 VDD.n223 0.607167
R3528 VDD.n222 VDD.t42 0.607167
R3529 VDD.n222 VDD.n221 0.607167
R3530 VDD.n220 VDD.t128 0.607167
R3531 VDD.n220 VDD.n219 0.607167
R3532 VDD.n1145 VDD.t222 0.607167
R3533 VDD.n1145 VDD.n1144 0.607167
R3534 VDD.n1142 VDD.t47 0.607167
R3535 VDD.n1142 VDD.n1141 0.607167
R3536 VDD.n215 VDD.t35 0.607167
R3537 VDD.n215 VDD.n214 0.607167
R3538 VDD.n213 VDD.t229 0.607167
R3539 VDD.n213 VDD.n212 0.607167
R3540 VDD.n211 VDD.t255 0.607167
R3541 VDD.n211 VDD.n210 0.607167
R3542 VDD.n1197 VDD.t126 0.607167
R3543 VDD.n202 VDD.t116 0.607167
R3544 VDD.n201 VDD.t164 0.607167
R3545 VDD.n200 VDD.t170 0.607167
R3546 VDD.n1946 VDD.t88 0.607167
R3547 VDD.n1946 VDD.n1945 0.607167
R3548 VDD.n1943 VDD.t160 0.607167
R3549 VDD.n1943 VDD.n1942 0.607167
R3550 VDD.n108 VDD.t151 0.607167
R3551 VDD.n108 VDD.n107 0.607167
R3552 VDD.n106 VDD.t185 0.607167
R3553 VDD.n106 VDD.n105 0.607167
R3554 VDD.n104 VDD.t187 0.607167
R3555 VDD.n104 VDD.n103 0.607167
R3556 VDD.n2336 VDD.t455 0.607167
R3557 VDD.n2336 VDD.n2335 0.607167
R3558 VDD.n2338 VDD.t468 0.607167
R3559 VDD.n2338 VDD.n2337 0.607167
R3560 VDD.n2929 VDD.t469 0.607167
R3561 VDD.n2929 VDD.n2928 0.607167
R3562 VDD.n2932 VDD.t315 0.607167
R3563 VDD.n2932 VDD.n2931 0.607167
R3564 VDD.n2217 VDD.t327 0.607167
R3565 VDD.n2217 VDD.n2216 0.607167
R3566 VDD.n2219 VDD.t458 0.607167
R3567 VDD.n2219 VDD.n2218 0.607167
R3568 VDD.n2221 VDD.t462 0.607167
R3569 VDD.n2221 VDD.n2220 0.607167
R3570 VDD.n2977 VDD.t454 0.607167
R3571 VDD.n2977 VDD.n2976 0.607167
R3572 VDD.n1981 VDD.t69 0.607167
R3573 VDD.n1961 VDD.t135 0.607167
R3574 VDD.n1961 VDD.n1960 0.607167
R3575 VDD.n1958 VDD.t210 0.607167
R3576 VDD.n1958 VDD.n1957 0.607167
R3577 VDD.n99 VDD.t203 0.607167
R3578 VDD.n99 VDD.n98 0.607167
R3579 VDD.n97 VDD.t115 0.607167
R3580 VDD.n97 VDD.n96 0.607167
R3581 VDD.n95 VDD.t92 0.607167
R3582 VDD.n95 VDD.n94 0.607167
R3583 VDD.n1940 VDD.t22 0.607167
R3584 VDD.n1940 VDD.n1939 0.607167
R3585 VDD.n1937 VDD.t121 0.607167
R3586 VDD.n1937 VDD.n1936 0.607167
R3587 VDD.n90 VDD.t111 0.607167
R3588 VDD.n90 VDD.n89 0.607167
R3589 VDD.n88 VDD.t204 0.607167
R3590 VDD.n88 VDD.n87 0.607167
R3591 VDD.n86 VDD.t38 0.607167
R3592 VDD.n86 VDD.n85 0.607167
R3593 VDD.n1978 VDD.t150 0.607167
R3594 VDD.n77 VDD.t140 0.607167
R3595 VDD.n76 VDD.t207 0.607167
R3596 VDD.n75 VDD.t139 0.607167
R3597 VDD.n1338 VDD.n1337 0.607167
R3598 VDD.n1334 VDD.n1333 0.607167
R3599 VDD.n129 VDD.t340 0.607167
R3600 VDD.n129 VDD.n128 0.607167
R3601 VDD.n125 VDD.t415 0.607167
R3602 VDD.n125 VDD.n124 0.607167
R3603 VDD.n123 VDD.t382 0.607167
R3604 VDD.n123 VDD.n122 0.607167
R3605 VDD.n1344 VDD.t40 0.607167
R3606 VDD.n1344 VDD.n1343 0.607167
R3607 VDD.n1341 VDD.t131 0.607167
R3608 VDD.n1341 VDD.n1340 0.607167
R3609 VDD.n117 VDD.t125 0.607167
R3610 VDD.n117 VDD.n116 0.607167
R3611 VDD.n115 VDD.t182 0.607167
R3612 VDD.n115 VDD.n114 0.607167
R3613 VDD.n113 VDD.t112 0.607167
R3614 VDD.n113 VDD.n112 0.607167
R3615 VDD.n2200 VDD.t430 0.607167
R3616 VDD.n2200 VDD.n2199 0.607167
R3617 VDD.n2202 VDD.t331 0.607167
R3618 VDD.n2202 VDD.n2201 0.607167
R3619 VDD.n2204 VDD.t421 0.607167
R3620 VDD.n2204 VDD.n2203 0.607167
R3621 VDD.n2634 VDD.t323 0.607167
R3622 VDD.n2634 VDD.n2633 0.607167
R3623 VDD.n1121 VDD.n1120 0.575213
R3624 VDD.n1011 VDD.t318 0.575213
R3625 VDD.n1292 VDD.n1291 0.575213
R3626 VDD.n400 VDD.n399 0.502139
R3627 VDD.n392 VDD.n391 0.502139
R3628 VDD.n333 VDD.n332 0.502139
R3629 VDD.n323 VDD.n322 0.502139
R3630 VDD.n272 VDD.n271 0.502139
R3631 VDD.n265 VDD.n264 0.502139
R3632 VDD.n209 VDD.n208 0.502139
R3633 VDD.n199 VDD.n198 0.502139
R3634 VDD.n84 VDD.n83 0.502139
R3635 VDD.n74 VDD.n73 0.502139
R3636 VDD.n147 VDD.n146 0.502139
R3637 VDD.n140 VDD.n139 0.502139
R3638 VDD.n1767 VDD.n1766 0.497765
R3639 VDD.n395 VDD.n394 0.490336
R3640 VDD.n385 VDD.n384 0.490336
R3641 VDD.n328 VDD.n327 0.490336
R3642 VDD.n316 VDD.n315 0.490336
R3643 VDD.n640 VDD.n637 0.490336
R3644 VDD.n644 VDD.n643 0.490336
R3645 VDD.n267 VDD.n266 0.490336
R3646 VDD.n258 VDD.n257 0.490336
R3647 VDD.n732 VDD.n731 0.490336
R3648 VDD.n727 VDD.n724 0.490336
R3649 VDD.n204 VDD.n203 0.490336
R3650 VDD.n192 VDD.n191 0.490336
R3651 VDD.n1139 VDD.n1136 0.490336
R3652 VDD.n1199 VDD.n1198 0.490336
R3653 VDD.n79 VDD.n78 0.490336
R3654 VDD.n67 VDD.n66 0.490336
R3655 VDD.n1934 VDD.n1931 0.490336
R3656 VDD.n1980 VDD.n1979 0.490336
R3657 VDD.n142 VDD.n141 0.490336
R3658 VDD.n133 VDD.n132 0.490336
R3659 VDD.n1336 VDD.n1335 0.490336
R3660 VDD.n1219 VDD.n1216 0.490336
R3661 VDD.n399 VDD.n398 0.488861
R3662 VDD.n391 VDD.n390 0.488861
R3663 VDD.n390 VDD.n387 0.488861
R3664 VDD.n387 VDD.n386 0.488861
R3665 VDD.n398 VDD.n397 0.488861
R3666 VDD.n397 VDD.n396 0.488861
R3667 VDD.n396 VDD.n395 0.488861
R3668 VDD.n386 VDD.n385 0.488861
R3669 VDD.n332 VDD.n331 0.488861
R3670 VDD.n322 VDD.n321 0.488861
R3671 VDD.n321 VDD.n318 0.488861
R3672 VDD.n318 VDD.n317 0.488861
R3673 VDD.n331 VDD.n330 0.488861
R3674 VDD.n330 VDD.n329 0.488861
R3675 VDD.n329 VDD.n328 0.488861
R3676 VDD.n317 VDD.n316 0.488861
R3677 VDD.n271 VDD.n270 0.488861
R3678 VDD.n264 VDD.n263 0.488861
R3679 VDD.n263 VDD.n260 0.488861
R3680 VDD.n260 VDD.n259 0.488861
R3681 VDD.n270 VDD.n269 0.488861
R3682 VDD.n269 VDD.n268 0.488861
R3683 VDD.n268 VDD.n267 0.488861
R3684 VDD.n259 VDD.n258 0.488861
R3685 VDD.n208 VDD.n207 0.488861
R3686 VDD.n198 VDD.n197 0.488861
R3687 VDD.n197 VDD.n194 0.488861
R3688 VDD.n194 VDD.n193 0.488861
R3689 VDD.n207 VDD.n206 0.488861
R3690 VDD.n206 VDD.n205 0.488861
R3691 VDD.n205 VDD.n204 0.488861
R3692 VDD.n193 VDD.n192 0.488861
R3693 VDD.n83 VDD.n82 0.488861
R3694 VDD.n73 VDD.n72 0.488861
R3695 VDD.n72 VDD.n69 0.488861
R3696 VDD.n69 VDD.n68 0.488861
R3697 VDD.n82 VDD.n81 0.488861
R3698 VDD.n81 VDD.n80 0.488861
R3699 VDD.n80 VDD.n79 0.488861
R3700 VDD.n68 VDD.n67 0.488861
R3701 VDD.n146 VDD.n145 0.488861
R3702 VDD.n139 VDD.n138 0.488861
R3703 VDD.n138 VDD.n135 0.488861
R3704 VDD.n135 VDD.n134 0.488861
R3705 VDD.n145 VDD.n144 0.488861
R3706 VDD.n144 VDD.n143 0.488861
R3707 VDD.n143 VDD.n142 0.488861
R3708 VDD.n134 VDD.n133 0.488861
R3709 VDD.n384 VDD.n381 0.487385
R3710 VDD.n394 VDD.n393 0.487385
R3711 VDD.n432 VDD.n431 0.487385
R3712 VDD.n436 VDD.n433 0.487385
R3713 VDD.n646 VDD.n644 0.487385
R3714 VDD.n641 VDD.n640 0.487385
R3715 VDD.n728 VDD.n727 0.487385
R3716 VDD.n735 VDD.n732 0.487385
R3717 VDD.n1201 VDD.n1199 0.487385
R3718 VDD.n1140 VDD.n1139 0.487385
R3719 VDD.n1982 VDD.n1980 0.487385
R3720 VDD.n1935 VDD.n1934 0.487385
R3721 VDD.n1220 VDD.n1219 0.487385
R3722 VDD.n1339 VDD.n1336 0.487385
R3723 VDD.n1671 VDD.n1670 0.430793
R3724 VDD.n2696 VDD.t436 0.430793
R3725 VDD.n2920 VDD.n2919 0.3518
R3726 VDD.n1070 VDD.n1069 0.329562
R3727 VDD.n1042 VDD.n1041 0.329562
R3728 VDD.n1309 VDD.n1308 0.32675
R3729 VDD.n1328 VDD.n1327 0.32675
R3730 VDD.n1327 VDD.n1324 0.322531
R3731 VDD.n1308 VDD.n1307 0.322531
R3732 VDD.n2055 VDD.n2054 0.3218
R3733 VDD.n2074 VDD.n2073 0.3218
R3734 VDD.n2093 VDD.n2092 0.3218
R3735 VDD.n2115 VDD.n2114 0.3218
R3736 VDD.n2138 VDD.n2137 0.3218
R3737 VDD.n2158 VDD.n2157 0.3218
R3738 VDD.n2033 VDD.n1612 0.3218
R3739 VDD.n2032 VDD.n2031 0.3218
R3740 VDD.n1041 VDD.n1038 0.319719
R3741 VDD.n1069 VDD.n1068 0.319719
R3742 VDD.n1928 VDD.n1805 0.2993
R3743 VDD.n1926 VDD.n1836 0.2993
R3744 VDD.n1925 VDD.n1921 0.2993
R3745 VDD.n1927 VDD.n1822 0.2993
R3746 VDD.n425 VDD.n424 0.297674
R3747 VDD.n1372 VDD.n1133 0.294837
R3748 VDD.n421 VDD.n420 0.293978
R3749 VDD.n2032 VDD.n1928 0.2921
R3750 VDD.n1867 VDD.n1853 0.286017
R3751 VDD.n1732 VDD.n1702 0.286017
R3752 VDD.n3094 VDD.n3093 0.282667
R3753 VDD.n2293 VDD.n2281 0.282667
R3754 VDD.n2616 VDD.n2615 0.260917
R3755 VDD.n2514 VDD.n2502 0.260917
R3756 VDD.n1363 VDD.n1332 0.2561
R3757 VDD.n1928 VDD.n1927 0.24575
R3758 VDD.n165 VDD.n163 0.239392
R3759 VDD.n1556 VDD.t91 0.239392
R3760 VDD.n54 VDD.n51 0.239392
R3761 VDD.n523 VDD.n522 0.239392
R3762 VDD.n580 VDD.t89 0.239392
R3763 VDD.n304 VDD.n302 0.239392
R3764 VDD.n289 VDD.n288 0.239392
R3765 VDD.n924 VDD.t41 0.239392
R3766 VDD.n179 VDD.n176 0.239392
R3767 VDD.n537 VDD.n536 0.239186
R3768 VDD.n3010 VDD.n2922 0.21425
R3769 VDD.n2055 VDD.n2043 0.19895
R3770 VDD.n2074 VDD.n2063 0.19895
R3771 VDD.n2093 VDD.n2081 0.19895
R3772 VDD.n2115 VDD.n2102 0.19895
R3773 VDD.n2138 VDD.n2126 0.19895
R3774 VDD.n2158 VDD.n2147 0.19895
R3775 VDD.n2167 VDD.n2166 0.19895
R3776 VDD.n2033 VDD.n1603 0.19895
R3777 VDD.n2032 VDD.n1996 0.19895
R3778 VDD.n2170 VDD.n2169 0.197926
R3779 VDD.n1041 VDD.n1040 0.18407
R3780 VDD.n1058 VDD.n1057 0.1805
R3781 VDD.n1059 VDD.n1058 0.1805
R3782 VDD.n1330 VDD.n1303 0.1805
R3783 VDD.n1926 VDD.n1925 0.1805
R3784 VDD.n1927 VDD.n1926 0.1805
R3785 VDD.n1130 VDD.n1129 0.1805
R3786 VDD.n1131 VDD.n1130 0.1805
R3787 VDD.n1132 VDD.n1131 0.1805
R3788 VDD.n1332 VDD.n1331 0.1805
R3789 VDD.n1327 VDD.n1326 0.18047
R3790 VDD.n550 VDD.n392 0.177549
R3791 VDD.n543 VDD.n400 0.177549
R3792 VDD.n613 VDD.n323 0.177549
R3793 VDD.n606 VDD.n333 0.177549
R3794 VDD.n894 VDD.n265 0.177549
R3795 VDD.n887 VDD.n272 0.177549
R3796 VDD.n957 VDD.n199 0.177549
R3797 VDD.n950 VDD.n209 0.177549
R3798 VDD.n1589 VDD.n74 0.177549
R3799 VDD.n1582 VDD.n84 0.177549
R3800 VDD.n1526 VDD.n140 0.177549
R3801 VDD.n1519 VDD.n147 0.177549
R3802 VDD.n536 VDD.n535 0.176669
R3803 VDD.n514 VDD.n513 0.173106
R3804 VDD.n530 VDD.n529 0.173106
R3805 VDD.n1925 VDD.n1924 0.1715
R3806 VDD.n1133 VDD.n1132 0.17105
R3807 VDD.n472 VDD.n468 0.1697
R3808 VDD.n461 VDD.n456 0.1697
R3809 VDD.n451 VDD.n425 0.1697
R3810 VDD.n2922 VDD.n2604 0.167375
R3811 VDD.n1780 VDD.n1701 0.1535
R3812 VDD.n3068 VDD.n3057 0.1505
R3813 VDD.n3057 VDD.n3044 0.1505
R3814 VDD.n3044 VDD.n3033 0.1505
R3815 VDD.n3033 VDD.n3021 0.1505
R3816 VDD.n3021 VDD.n3010 0.1505
R3817 VDD.n2604 VDD.n2603 0.1505
R3818 VDD.n2603 VDD.n2602 0.1505
R3819 VDD.n2602 VDD.n2601 0.1505
R3820 VDD.n2601 VDD.n2600 0.1505
R3821 VDD.n2921 VDD.n2920 0.1505
R3822 VDD.n2919 VDD.n2918 0.1505
R3823 VDD.n2918 VDD.n2917 0.1505
R3824 VDD.n2917 VDD.n2916 0.1505
R3825 VDD.n2916 VDD.n2915 0.1505
R3826 VDD.n2915 VDD.n2904 0.1505
R3827 VDD.n1952 VDD.n1951 0.14675
R3828 VDD.n1133 VDD.n1015 0.134122
R3829 VDD.n1332 VDD.n1330 0.13145
R3830 VDD.n1129 VDD.n1128 0.13145
R3831 VDD.n1132 VDD.n1059 0.13145
R3832 VDD.n2922 VDD.n2921 0.12875
R3833 VDD.n1015 VDD.n1014 0.127235
R3834 VDD.n773 VDD.n763 0.12695
R3835 VDD.n794 VDD.n783 0.12695
R3836 VDD.n811 VDD.n802 0.12695
R3837 VDD.n830 VDD.n820 0.12695
R3838 VDD.n852 VDD.n841 0.12695
R3839 VDD.n868 VDD.n861 0.12695
R3840 VDD.n878 VDD.n877 0.12695
R3841 VDD.n755 VDD.n627 0.12695
R3842 VDD.n754 VDD.n720 0.12695
R3843 VDD.n2917 VDD.n2776 0.12515
R3844 VDD.n2916 VDD.n2797 0.12515
R3845 VDD.n2918 VDD.n2757 0.12515
R3846 VDD.n2915 VDD.n2914 0.12515
R3847 VDD.n1128 VDD.n1127 0.1247
R3848 VDD.n1330 VDD.n1329 0.1247
R3849 VDD.n1372 VDD.n1215 0.12425
R3850 VDD.n1389 VDD.n1380 0.12425
R3851 VDD.n1406 VDD.n1397 0.12425
R3852 VDD.n1427 VDD.n1416 0.12425
R3853 VDD.n1444 VDD.n1435 0.12425
R3854 VDD.n1463 VDD.n1453 0.12425
R3855 VDD.n1481 VDD.n1472 0.12425
R3856 VDD.n1501 VDD.n1492 0.12425
R3857 VDD.n1510 VDD.n1509 0.12425
R3858 VDD.n1372 VDD.n1371 0.12065
R3859 VDD.n1389 VDD.n1388 0.12065
R3860 VDD.n1406 VDD.n1405 0.12065
R3861 VDD.n1427 VDD.n1426 0.12065
R3862 VDD.n1444 VDD.n1443 0.12065
R3863 VDD.n1463 VDD.n1462 0.12065
R3864 VDD.n1481 VDD.n1480 0.12065
R3865 VDD.n1501 VDD.n1500 0.12065
R3866 VDD.n2919 VDD.n2746 0.11885
R3867 VDD.n2918 VDD.n2768 0.11885
R3868 VDD.n2917 VDD.n2789 0.11885
R3869 VDD.n2916 VDD.n2808 0.11885
R3870 VDD.n2915 VDD.n2819 0.11885
R3871 VDD.n2904 VDD.n2903 0.11885
R3872 VDD.n773 VDD.n772 0.11795
R3873 VDD.n794 VDD.n793 0.11795
R3874 VDD.n811 VDD.n810 0.11795
R3875 VDD.n830 VDD.n829 0.11795
R3876 VDD.n852 VDD.n851 0.11795
R3877 VDD.n868 VDD.n867 0.11795
R3878 VDD.n755 VDD.n636 0.11795
R3879 VDD.n754 VDD.n753 0.11795
R3880 VDD.n3109 VDD.n2373 0.117525
R3881 VDD.n3072 VDD.n3068 0.113
R3882 VDD.n2922 VDD.n2451 0.10925
R3883 VDD.n2904 VDD.n2843 0.1031
R3884 VDD.n2919 VDD.n2730 0.1031
R3885 VDD.n1057 VDD.n1056 0.10265
R3886 VDD.n1058 VDD.n1028 0.10265
R3887 VDD.n1303 VDD.n1302 0.10265
R3888 VDD.n392 VDD.n370 0.0990135
R3889 VDD.n390 VDD.n389 0.0990135
R3890 VDD.n386 VDD.n376 0.0990135
R3891 VDD.n384 VDD.n383 0.0990135
R3892 VDD.n323 VDD.n310 0.0990135
R3893 VDD.n321 VDD.n320 0.0990135
R3894 VDD.n317 VDD.n312 0.0990135
R3895 VDD.n315 VDD.n314 0.0990135
R3896 VDD.n640 VDD.n639 0.0990135
R3897 VDD.n265 VDD.n246 0.0990135
R3898 VDD.n263 VDD.n262 0.0990135
R3899 VDD.n259 VDD.n252 0.0990135
R3900 VDD.n257 VDD.n256 0.0990135
R3901 VDD.n199 VDD.n186 0.0990135
R3902 VDD.n197 VDD.n196 0.0990135
R3903 VDD.n193 VDD.n188 0.0990135
R3904 VDD.n191 VDD.n190 0.0990135
R3905 VDD.n1139 VDD.n1138 0.0990135
R3906 VDD.n74 VDD.n61 0.0990135
R3907 VDD.n72 VDD.n71 0.0990135
R3908 VDD.n68 VDD.n63 0.0990135
R3909 VDD.n66 VDD.n65 0.0990135
R3910 VDD.n1934 VDD.n1933 0.0990135
R3911 VDD.n140 VDD.n121 0.0990135
R3912 VDD.n138 VDD.n137 0.0990135
R3913 VDD.n134 VDD.n127 0.0990135
R3914 VDD.n132 VDD.n131 0.0990135
R3915 VDD.n1512 VDD.n1511 0.0969286
R3916 VDD.n2169 VDD.n1595 0.095826
R3917 VDD.n880 VDD.n879 0.095551
R3918 VDD.n431 VDD.n430 0.0953649
R3919 VDD.n727 VDD.n726 0.0953649
R3920 VDD.n1219 VDD.n1218 0.0953649
R3921 VDD.n2601 VDD.n2501 0.0941
R3922 VDD.n2602 VDD.n2489 0.0941
R3923 VDD.n2603 VDD.n2477 0.0941
R3924 VDD.n2604 VDD.n2465 0.0941
R3925 VDD.n2600 VDD.n2599 0.0941
R3926 VDD.n514 VDD.n421 0.0938803
R3927 VDD.n535 VDD.n534 0.0938803
R3928 VDD.n2434 VDD.n2431 0.0932551
R3929 VDD.n2015 VDD.n2013 0.0932551
R3930 VDD.n2007 VDD.n2005 0.0932551
R3931 VDD.n2643 VDD.n2641 0.0932551
R3932 VDD.n2652 VDD.n2650 0.0932551
R3933 VDD.n2660 VDD.n2658 0.0932551
R3934 VDD.n773 VDD.n755 0.0923367
R3935 VDD.n794 VDD.n773 0.0923367
R3936 VDD.n811 VDD.n794 0.0923367
R3937 VDD.n830 VDD.n811 0.0923367
R3938 VDD.n852 VDD.n830 0.0923367
R3939 VDD.n878 VDD.n868 0.0923367
R3940 VDD.n868 VDD.n852 0.0923367
R3941 VDD.n1389 VDD.n1372 0.0923367
R3942 VDD.n1406 VDD.n1389 0.0923367
R3943 VDD.n1427 VDD.n1406 0.0923367
R3944 VDD.n1444 VDD.n1427 0.0923367
R3945 VDD.n1463 VDD.n1444 0.0923367
R3946 VDD.n1481 VDD.n1463 0.0923367
R3947 VDD.n1510 VDD.n1501 0.0923367
R3948 VDD.n1501 VDD.n1481 0.0923367
R3949 VDD.n755 VDD.n754 0.0923367
R3950 VDD.n879 VDD.n878 0.0923367
R3951 VDD.n1511 VDD.n1510 0.0923367
R3952 VDD.n2169 VDD.n2168 0.09185
R3953 VDD.n2055 VDD.n2033 0.0905
R3954 VDD.n2074 VDD.n2055 0.0905
R3955 VDD.n2093 VDD.n2074 0.0905
R3956 VDD.n2115 VDD.n2093 0.0905
R3957 VDD.n2138 VDD.n2115 0.0905
R3958 VDD.n2158 VDD.n2138 0.0905
R3959 VDD.n2167 VDD.n2158 0.0905
R3960 VDD.n2168 VDD.n2167 0.0905
R3961 VDD.n2033 VDD.n2032 0.0905
R3962 VDD.n1700 VDD.n1698 0.0886633
R3963 VDD.n2724 VDD.n2722 0.0886633
R3964 VDD.n2446 VDD.n2444 0.0886633
R3965 VDD.n43 VDD.n30 0.0886633
R3966 VDD.n13 VDD.n11 0.0886633
R3967 VDD.n2133 VDD.n2131 0.0886633
R3968 VDD.n1609 VDD.n1607 0.0886633
R3969 VDD.n2027 VDD.n2025 0.0886633
R3970 VDD.n2639 VDD.n2637 0.0886633
R3971 VDD.n2656 VDD.n2654 0.0886633
R3972 VDD.n2296 VDD.n2280 0.088625
R3973 VDD.n2280 VDD.n2278 0.088625
R3974 VDD.n2278 VDD.n2275 0.088625
R3975 VDD.n2275 VDD.n2273 0.088625
R3976 VDD.n2273 VDD.n2270 0.088625
R3977 VDD.n2270 VDD.n2268 0.088625
R3978 VDD.n2268 VDD.n2265 0.088625
R3979 VDD.n2265 VDD.n2263 0.088625
R3980 VDD.n2263 VDD.n2260 0.088625
R3981 VDD.n2260 VDD.n2258 0.088625
R3982 VDD.n2258 VDD.n2255 0.088625
R3983 VDD.n2255 VDD.n2253 0.088625
R3984 VDD.n2253 VDD.n2250 0.088625
R3985 VDD.n2250 VDD.n2248 0.088625
R3986 VDD.n2248 VDD.n2246 0.088625
R3987 VDD.n2246 VDD.n2244 0.088625
R3988 VDD.n2244 VDD.n2242 0.088625
R3989 VDD.n2242 VDD.n2240 0.088625
R3990 VDD.n2240 VDD.n2238 0.088625
R3991 VDD.n2238 VDD.n2236 0.088625
R3992 VDD.n2236 VDD.n2234 0.088625
R3993 VDD.n2234 VDD.n2232 0.088625
R3994 VDD.n2232 VDD.n2230 0.088625
R3995 VDD.n2230 VDD.n2228 0.088625
R3996 VDD.n2228 VDD.n2226 0.088625
R3997 VDD.n2940 VDD.n2938 0.088625
R3998 VDD.n2942 VDD.n2940 0.088625
R3999 VDD.n2944 VDD.n2942 0.088625
R4000 VDD.n2946 VDD.n2944 0.088625
R4001 VDD.n2948 VDD.n2946 0.088625
R4002 VDD.n2950 VDD.n2948 0.088625
R4003 VDD.n2952 VDD.n2950 0.088625
R4004 VDD.n2954 VDD.n2952 0.088625
R4005 VDD.n2956 VDD.n2954 0.088625
R4006 VDD.n2958 VDD.n2956 0.088625
R4007 VDD.n2730 VDD.n2729 0.0877449
R4008 VDD.n2373 VDD.n2372 0.0872537
R4009 VDD.n1599 VDD.n1597 0.0868265
R4010 VDD.n2037 VDD.n2035 0.0868265
R4011 VDD.n2098 VDD.n2095 0.0868265
R4012 VDD.n2120 VDD.n2117 0.0868265
R4013 VDD.n151 VDD.n149 0.0868265
R4014 VDD.n1496 VDD.n1494 0.0868265
R4015 VDD.n1476 VDD.n1474 0.0868265
R4016 VDD.n1458 VDD.n1456 0.0868265
R4017 VDD.n1422 VDD.n1420 0.0868265
R4018 VDD.n1401 VDD.n1399 0.0868265
R4019 VDD.n1384 VDD.n1382 0.0868265
R4020 VDD.n50 VDD.n48 0.0868265
R4021 VDD.n162 VDD.n160 0.0868265
R4022 VDD.n160 VDD.n157 0.0868265
R4023 VDD.n466 VDD.n464 0.0868265
R4024 VDD.n476 VDD.n474 0.0868265
R4025 VDD.n503 VDD.n500 0.0868265
R4026 VDD.n500 VDD.n497 0.0868265
R4027 VDD.n497 VDD.n494 0.0868265
R4028 VDD.n494 VDD.n491 0.0868265
R4029 VDD.n491 VDD.n488 0.0868265
R4030 VDD.n488 VDD.n485 0.0868265
R4031 VDD.n485 VDD.n483 0.0868265
R4032 VDD.n519 VDD.n517 0.0868265
R4033 VDD.n300 VDD.n298 0.0868265
R4034 VDD.n837 VDD.n834 0.0868265
R4035 VDD.n816 VDD.n813 0.0868265
R4036 VDD.n779 VDD.n777 0.0868265
R4037 VDD.n759 VDD.n757 0.0868265
R4038 VDD.n455 VDD.n453 0.0868265
R4039 VDD.n450 VDD.n448 0.0868265
R4040 VDD.n445 VDD.n443 0.0868265
R4041 VDD.n440 VDD.n438 0.0868265
R4042 VDD.n674 VDD.n672 0.0868265
R4043 VDD.n679 VDD.n677 0.0868265
R4044 VDD.n681 VDD.n679 0.0868265
R4045 VDD.n686 VDD.n684 0.0868265
R4046 VDD.n688 VDD.n686 0.0868265
R4047 VDD.n693 VDD.n691 0.0868265
R4048 VDD.n695 VDD.n693 0.0868265
R4049 VDD.n697 VDD.n695 0.0868265
R4050 VDD.n702 VDD.n700 0.0868265
R4051 VDD.n704 VDD.n702 0.0868265
R4052 VDD.n709 VDD.n707 0.0868265
R4053 VDD.n714 VDD.n712 0.0868265
R4054 VDD.n623 VDD.n621 0.0868265
R4055 VDD.n845 VDD.n843 0.0868265
R4056 VDD.n789 VDD.n787 0.0868265
R4057 VDD.n768 VDD.n766 0.0868265
R4058 VDD.n632 VDD.n629 0.0868265
R4059 VDD.n825 VDD.n823 0.0868265
R4060 VDD.n276 VDD.n274 0.0868265
R4061 VDD.n287 VDD.n285 0.0868265
R4062 VDD.n285 VDD.n282 0.0868265
R4063 VDD.n1376 VDD.n1374 0.0868265
R4064 VDD.n1393 VDD.n1391 0.0868265
R4065 VDD.n1410 VDD.n1408 0.0868265
R4066 VDD.n1449 VDD.n1446 0.0868265
R4067 VDD.n1468 VDD.n1465 0.0868265
R4068 VDD.n1486 VDD.n1483 0.0868265
R4069 VDD.n749 VDD.n747 0.0868265
R4070 VDD.n744 VDD.n742 0.0868265
R4071 VDD.n739 VDD.n737 0.0868265
R4072 VDD.n1156 VDD.n1154 0.0868265
R4073 VDD.n1161 VDD.n1159 0.0868265
R4074 VDD.n1175 VDD.n1173 0.0868265
R4075 VDD.n1189 VDD.n1187 0.0868265
R4076 VDD.n1206 VDD.n1204 0.0868265
R4077 VDD.n1212 VDD.n1210 0.0868265
R4078 VDD.n1801 VDD.n1798 0.0868265
R4079 VDD.n1804 VDD.n1801 0.0868265
R4080 VDD.n1814 VDD.n1811 0.0868265
R4081 VDD.n1835 VDD.n1832 0.0868265
R4082 VDD.n1920 VDD.n1917 0.0868265
R4083 VDD.n1912 VDD.n1909 0.0868265
R4084 VDD.n1909 VDD.n1907 0.0868265
R4085 VDD.n1900 VDD.n1897 0.0868265
R4086 VDD.n1891 VDD.n1888 0.0868265
R4087 VDD.n1880 VDD.n1878 0.0868265
R4088 VDD.n969 VDD.n966 0.0868265
R4089 VDD.n1048 VDD.n1045 0.0868265
R4090 VDD.n1021 VDD.n1018 0.0868265
R4091 VDD.n1024 VDD.n1021 0.0868265
R4092 VDD.n989 VDD.n986 0.0868265
R4093 VDD.n1281 VDD.n1279 0.0868265
R4094 VDD.n1289 VDD.n1287 0.0868265
R4095 VDD.n1299 VDD.n1297 0.0868265
R4096 VDD.n1316 VDD.n1313 0.0868265
R4097 VDD.n1082 VDD.n1080 0.0868265
R4098 VDD.n1080 VDD.n1078 0.0868265
R4099 VDD.n1078 VDD.n1076 0.0868265
R4100 VDD.n1076 VDD.n1074 0.0868265
R4101 VDD.n1074 VDD.n1072 0.0868265
R4102 VDD.n1036 VDD.n1034 0.0868265
R4103 VDD.n973 VDD.n971 0.0868265
R4104 VDD.n975 VDD.n973 0.0868265
R4105 VDD.n977 VDD.n975 0.0868265
R4106 VDD.n1233 VDD.n1231 0.0868265
R4107 VDD.n1235 VDD.n1233 0.0868265
R4108 VDD.n1237 VDD.n1235 0.0868265
R4109 VDD.n1242 VDD.n1240 0.0868265
R4110 VDD.n1244 VDD.n1242 0.0868265
R4111 VDD.n1246 VDD.n1244 0.0868265
R4112 VDD.n1248 VDD.n1246 0.0868265
R4113 VDD.n1250 VDD.n1248 0.0868265
R4114 VDD.n1255 VDD.n1253 0.0868265
R4115 VDD.n1257 VDD.n1255 0.0868265
R4116 VDD.n1259 VDD.n1257 0.0868265
R4117 VDD.n1124 VDD.n1119 0.0868265
R4118 VDD.n1119 VDD.n1117 0.0868265
R4119 VDD.n1117 VDD.n1114 0.0868265
R4120 VDD.n1114 VDD.n1112 0.0868265
R4121 VDD.n1112 VDD.n1109 0.0868265
R4122 VDD.n1109 VDD.n1107 0.0868265
R4123 VDD.n1107 VDD.n1104 0.0868265
R4124 VDD.n1104 VDD.n1102 0.0868265
R4125 VDD.n1102 VDD.n1099 0.0868265
R4126 VDD.n1099 VDD.n1097 0.0868265
R4127 VDD.n1097 VDD.n1094 0.0868265
R4128 VDD.n1094 VDD.n1092 0.0868265
R4129 VDD.n1092 VDD.n1089 0.0868265
R4130 VDD.n1089 VDD.n1087 0.0868265
R4131 VDD.n1087 VDD.n1084 0.0868265
R4132 VDD.n1275 VDD.n1272 0.0868265
R4133 VDD.n1272 VDD.n1270 0.0868265
R4134 VDD.n1270 VDD.n1267 0.0868265
R4135 VDD.n1873 VDD.n1871 0.0868265
R4136 VDD.n1871 VDD.n1869 0.0868265
R4137 VDD.n1866 VDD.n1864 0.0868265
R4138 VDD.n1864 VDD.n1862 0.0868265
R4139 VDD.n1859 VDD.n1857 0.0868265
R4140 VDD.n1709 VDD.n1707 0.0868265
R4141 VDD.n1711 VDD.n1709 0.0868265
R4142 VDD.n1713 VDD.n1711 0.0868265
R4143 VDD.n1718 VDD.n1716 0.0868265
R4144 VDD.n1720 VDD.n1718 0.0868265
R4145 VDD.n1722 VDD.n1720 0.0868265
R4146 VDD.n1724 VDD.n1722 0.0868265
R4147 VDD.n1726 VDD.n1724 0.0868265
R4148 VDD.n1731 VDD.n1729 0.0868265
R4149 VDD.n1736 VDD.n1734 0.0868265
R4150 VDD.n1738 VDD.n1736 0.0868265
R4151 VDD.n1748 VDD.n1746 0.0868265
R4152 VDD.n1756 VDD.n1754 0.0868265
R4153 VDD.n1764 VDD.n1762 0.0868265
R4154 VDD.n1659 VDD.n1656 0.0868265
R4155 VDD.n1653 VDD.n1651 0.0868265
R4156 VDD.n1648 VDD.n1646 0.0868265
R4157 VDD.n1641 VDD.n1639 0.0868265
R4158 VDD.n1639 VDD.n1637 0.0868265
R4159 VDD.n1637 VDD.n1635 0.0868265
R4160 VDD.n1635 VDD.n1633 0.0868265
R4161 VDD.n1633 VDD.n1631 0.0868265
R4162 VDD.n1631 VDD.n1629 0.0868265
R4163 VDD.n1629 VDD.n1627 0.0868265
R4164 VDD.n1627 VDD.n1625 0.0868265
R4165 VDD.n2826 VDD.n2824 0.0868265
R4166 VDD.n2828 VDD.n2826 0.0868265
R4167 VDD.n2830 VDD.n2828 0.0868265
R4168 VDD.n2832 VDD.n2830 0.0868265
R4169 VDD.n2834 VDD.n2832 0.0868265
R4170 VDD.n2836 VDD.n2834 0.0868265
R4171 VDD.n2838 VDD.n2836 0.0868265
R4172 VDD.n2840 VDD.n2838 0.0868265
R4173 VDD.n2750 VDD.n2748 0.0868265
R4174 VDD.n2775 VDD.n2773 0.0868265
R4175 VDD.n2796 VDD.n2794 0.0868265
R4176 VDD.n1668 VDD.n1665 0.0868265
R4177 VDD.n1696 VDD.n1694 0.0868265
R4178 VDD.n1694 VDD.n1691 0.0868265
R4179 VDD.n1691 VDD.n1688 0.0868265
R4180 VDD.n1688 VDD.n1685 0.0868265
R4181 VDD.n1685 VDD.n1682 0.0868265
R4182 VDD.n1682 VDD.n1679 0.0868265
R4183 VDD.n1679 VDD.n1676 0.0868265
R4184 VDD.n2695 VDD.n2692 0.0868265
R4185 VDD.n2698 VDD.n2695 0.0868265
R4186 VDD.n2701 VDD.n2698 0.0868265
R4187 VDD.n2704 VDD.n2701 0.0868265
R4188 VDD.n2707 VDD.n2704 0.0868265
R4189 VDD.n2710 VDD.n2707 0.0868265
R4190 VDD.n2713 VDD.n2710 0.0868265
R4191 VDD.n2716 VDD.n2713 0.0868265
R4192 VDD.n2719 VDD.n2716 0.0868265
R4193 VDD.n2729 VDD.n2726 0.0868265
R4194 VDD.n2495 VDD.n2492 0.0868265
R4195 VDD.n2483 VDD.n2480 0.0868265
R4196 VDD.n2471 VDD.n2468 0.0868265
R4197 VDD.n2457 VDD.n2454 0.0868265
R4198 VDD.n2619 VDD.n2614 0.0868265
R4199 VDD.n2627 VDD.n2624 0.0868265
R4200 VDD.n2624 VDD.n2621 0.0868265
R4201 VDD.n2688 VDD.n2686 0.0868265
R4202 VDD.n2686 VDD.n2683 0.0868265
R4203 VDD.n2683 VDD.n2681 0.0868265
R4204 VDD.n2681 VDD.n2678 0.0868265
R4205 VDD.n2678 VDD.n2676 0.0868265
R4206 VDD.n2676 VDD.n2673 0.0868265
R4207 VDD.n2673 VDD.n2671 0.0868265
R4208 VDD.n2734 VDD.n2732 0.0868265
R4209 VDD.n2737 VDD.n2734 0.0868265
R4210 VDD.n2745 VDD.n2742 0.0868265
R4211 VDD.n2742 VDD.n2740 0.0868265
R4212 VDD.n2767 VDD.n2764 0.0868265
R4213 VDD.n2764 VDD.n2762 0.0868265
R4214 VDD.n2781 VDD.n2778 0.0868265
R4215 VDD.n2788 VDD.n2786 0.0868265
R4216 VDD.n2786 VDD.n2783 0.0868265
R4217 VDD.n2807 VDD.n2805 0.0868265
R4218 VDD.n2805 VDD.n2802 0.0868265
R4219 VDD.n2818 VDD.n2815 0.0868265
R4220 VDD.n2815 VDD.n2812 0.0868265
R4221 VDD.n2897 VDD.n2895 0.0868265
R4222 VDD.n2895 VDD.n2893 0.0868265
R4223 VDD.n2893 VDD.n2891 0.0868265
R4224 VDD.n2891 VDD.n2889 0.0868265
R4225 VDD.n2889 VDD.n2887 0.0868265
R4226 VDD.n2887 VDD.n2885 0.0868265
R4227 VDD.n2885 VDD.n2883 0.0868265
R4228 VDD.n2883 VDD.n2881 0.0868265
R4229 VDD.n2881 VDD.n2879 0.0868265
R4230 VDD.n2879 VDD.n2877 0.0868265
R4231 VDD.n2877 VDD.n2875 0.0868265
R4232 VDD.n2875 VDD.n2873 0.0868265
R4233 VDD.n2873 VDD.n2871 0.0868265
R4234 VDD.n2871 VDD.n2869 0.0868265
R4235 VDD.n2869 VDD.n2867 0.0868265
R4236 VDD.n2867 VDD.n2865 0.0868265
R4237 VDD.n2865 VDD.n2863 0.0868265
R4238 VDD.n2863 VDD.n2861 0.0868265
R4239 VDD.n2861 VDD.n2859 0.0868265
R4240 VDD.n2859 VDD.n2857 0.0868265
R4241 VDD.n2857 VDD.n2855 0.0868265
R4242 VDD.n2589 VDD.n2587 0.0868265
R4243 VDD.n2587 VDD.n2584 0.0868265
R4244 VDD.n2584 VDD.n2582 0.0868265
R4245 VDD.n2582 VDD.n2579 0.0868265
R4246 VDD.n2579 VDD.n2577 0.0868265
R4247 VDD.n2577 VDD.n2574 0.0868265
R4248 VDD.n2574 VDD.n2572 0.0868265
R4249 VDD.n2572 VDD.n2569 0.0868265
R4250 VDD.n2569 VDD.n2567 0.0868265
R4251 VDD.n2567 VDD.n2564 0.0868265
R4252 VDD.n2564 VDD.n2562 0.0868265
R4253 VDD.n2562 VDD.n2559 0.0868265
R4254 VDD.n2559 VDD.n2557 0.0868265
R4255 VDD.n2557 VDD.n2554 0.0868265
R4256 VDD.n2554 VDD.n2552 0.0868265
R4257 VDD.n2552 VDD.n2550 0.0868265
R4258 VDD.n2550 VDD.n2548 0.0868265
R4259 VDD.n2548 VDD.n2546 0.0868265
R4260 VDD.n2546 VDD.n2544 0.0868265
R4261 VDD.n2544 VDD.n2542 0.0868265
R4262 VDD.n2542 VDD.n2540 0.0868265
R4263 VDD.n2540 VDD.n2538 0.0868265
R4264 VDD.n2538 VDD.n2536 0.0868265
R4265 VDD.n2536 VDD.n2534 0.0868265
R4266 VDD.n2534 VDD.n2532 0.0868265
R4267 VDD.n2532 VDD.n2530 0.0868265
R4268 VDD.n2530 VDD.n2528 0.0868265
R4269 VDD.n2528 VDD.n2526 0.0868265
R4270 VDD.n2526 VDD.n2524 0.0868265
R4271 VDD.n2524 VDD.n2522 0.0868265
R4272 VDD.n2522 VDD.n2520 0.0868265
R4273 VDD.n2520 VDD.n2518 0.0868265
R4274 VDD.n2847 VDD.n2845 0.0868265
R4275 VDD.n2849 VDD.n2847 0.0868265
R4276 VDD.n2851 VDD.n2849 0.0868265
R4277 VDD.n2853 VDD.n2851 0.0868265
R4278 VDD.n2436 VDD.n2434 0.0868265
R4279 VDD.n2431 VDD.n2429 0.0868265
R4280 VDD.n2422 VDD.n2419 0.0868265
R4281 VDD.n2412 VDD.n2409 0.0868265
R4282 VDD.n2403 VDD.n2400 0.0868265
R4283 VDD.n2393 VDD.n2390 0.0868265
R4284 VDD.n2383 VDD.n2380 0.0868265
R4285 VDD.n2969 VDD.n2967 0.0868265
R4286 VDD.n2996 VDD.n2994 0.0868265
R4287 VDD.n3007 VDD.n3004 0.0868265
R4288 VDD.n3017 VDD.n3015 0.0868265
R4289 VDD.n3029 VDD.n3027 0.0868265
R4290 VDD.n3040 VDD.n3038 0.0868265
R4291 VDD.n3053 VDD.n3051 0.0868265
R4292 VDD.n3064 VDD.n3061 0.0868265
R4293 VDD.n3092 VDD.n3089 0.0868265
R4294 VDD.n2371 VDD.n2369 0.0868265
R4295 VDD.n3082 VDD.n3080 0.0868265
R4296 VDD.n3085 VDD.n3082 0.0868265
R4297 VDD.n2913 VDD.n2910 0.0868265
R4298 VDD.n1779 VDD.n1777 0.0868265
R4299 VDD.n1777 VDD.n1774 0.0868265
R4300 VDD.n1774 VDD.n1772 0.0868265
R4301 VDD.n1956 VDD.n1954 0.0868265
R4302 VDD.n1970 VDD.n1968 0.0868265
R4303 VDD.n1987 VDD.n1985 0.0868265
R4304 VDD.n1993 VDD.n1991 0.0868265
R4305 VDD.n1359 VDD.n1357 0.0868265
R4306 VDD.n1354 VDD.n1352 0.0868265
R4307 VDD.n1349 VDD.n1347 0.0868265
R4308 VDD.n175 VDD.n173 0.0868265
R4309 VDD.n416 VDD.n413 0.0868265
R4310 VDD.n413 VDD.n410 0.0868265
R4311 VDD.n410 VDD.n407 0.0868265
R4312 VDD.n407 VDD.n405 0.0868265
R4313 VDD.n405 VDD.n402 0.0868265
R4314 VDD.n27 VDD.n24 0.0868265
R4315 VDD.n24 VDD.n22 0.0868265
R4316 VDD.n22 VDD.n19 0.0868265
R4317 VDD.n16 VDD.n13 0.0868265
R4318 VDD.n2156 VDD.n2153 0.0868265
R4319 VDD.n2153 VDD.n2151 0.0868265
R4320 VDD.n2136 VDD.n2133 0.0868265
R4321 VDD.n2113 VDD.n2110 0.0868265
R4322 VDD.n2110 VDD.n2108 0.0868265
R4323 VDD.n2086 VDD.n2083 0.0868265
R4324 VDD.n2091 VDD.n2089 0.0868265
R4325 VDD.n2068 VDD.n2065 0.0868265
R4326 VDD.n2072 VDD.n2070 0.0868265
R4327 VDD.n2047 VDD.n2045 0.0868265
R4328 VDD.n2053 VDD.n2051 0.0868265
R4329 VDD.n2051 VDD.n2049 0.0868265
R4330 VDD.n1611 VDD.n1609 0.0868265
R4331 VDD.n2030 VDD.n2028 0.0868265
R4332 VDD.n2028 VDD.n2027 0.0868265
R4333 VDD.n2025 VDD.n2023 0.0868265
R4334 VDD.n2023 VDD.n2021 0.0868265
R4335 VDD.n2019 VDD.n2017 0.0868265
R4336 VDD.n2017 VDD.n2015 0.0868265
R4337 VDD.n2013 VDD.n2011 0.0868265
R4338 VDD.n2011 VDD.n2009 0.0868265
R4339 VDD.n2009 VDD.n2007 0.0868265
R4340 VDD.n2641 VDD.n2639 0.0868265
R4341 VDD.n2645 VDD.n2643 0.0868265
R4342 VDD.n2650 VDD.n2648 0.0868265
R4343 VDD.n2654 VDD.n2652 0.0868265
R4344 VDD.n2658 VDD.n2656 0.0868265
R4345 VDD.n2662 VDD.n2660 0.0868265
R4346 VDD.n2439 VDD.n2436 0.0866336
R4347 VDD.n2610 VDD.n2608 0.0853043
R4348 VDD.n1654 VDD.n1653 0.0849898
R4349 VDD.n2768 VDD.n2759 0.0849898
R4350 VDD.n3072 VDD.n3071 0.0849898
R4351 VDD.n2092 VDD.n2091 0.0849898
R4352 VDD.n677 VDD.n675 0.0840714
R4353 VDD.n1159 VDD.n1157 0.0840714
R4354 VDD.n2981 VDD.n2979 0.0840714
R4355 VDD.n1350 VDD.n1349 0.0840714
R4356 VDD.n464 VDD.n461 0.0831531
R4357 VDD.n529 VDD.n519 0.0831531
R4358 VDD.n513 VDD.n505 0.0822347
R4359 VDD.n448 VDD.n446 0.0822347
R4360 VDD.n747 VDD.n745 0.0822347
R4361 VDD.n1888 VDD.n1886 0.0822347
R4362 VDD.n1729 VDD.n1727 0.0822347
R4363 VDD.n2992 VDD.n2987 0.0822347
R4364 VDD.n3056 VDD.n3053 0.0814388
R4365 VDD.n2114 VDD.n2105 0.0813163
R4366 VDD.n3009 VDD.n3007 0.0804592
R4367 VDD.n1886 VDD.n1880 0.080398
R4368 VDD.n1716 VDD.n1714 0.080398
R4369 VDD.n2994 VDD.n2992 0.080398
R4370 VDD.n2914 VDD.n2913 0.080398
R4371 VDD.n461 VDD.n455 0.0794796
R4372 VDD.n2465 VDD.n2457 0.0794796
R4373 VDD.n2385 VDD.n2383 0.0790225
R4374 VDD.n1262 VDD.n1260 0.0785612
R4375 VDD.n1860 VDD.n1859 0.0785612
R4376 VDD.n2599 VDD.n2590 0.0785612
R4377 VDD.n530 VDD.n514 0.0780352
R4378 VDD.n2166 VDD.n2161 0.0776429
R4379 VDD.n1656 VDD.n1654 0.0776429
R4380 VDD.n1357 VDD.n1355 0.0767245
R4381 VDD.n2081 VDD.n2076 0.0758061
R4382 VDD.n1251 VDD.n1250 0.0758061
R4383 VDD.n1127 VDD.n1126 0.0748878
R4384 VDD.n877 VDD.n873 0.0739694
R4385 VDD.n689 VDD.n688 0.0739694
R4386 VDD.n280 VDD.n276 0.0739694
R4387 VDD.n1279 VDD.n1276 0.0739694
R4388 VDD.n1770 VDD.n1764 0.0739694
R4389 VDD.n802 VDD.n798 0.0721327
R4390 VDD.n810 VDD.n804 0.0721327
R4391 VDD.n1265 VDD.n1264 0.0721327
R4392 VDD.n1782 VDD.n1780 0.0721327
R4393 VDD.n155 VDD.n151 0.0712143
R4394 VDD.n1056 VDD.n1055 0.0712143
R4395 VDD.n1509 VDD.n1503 0.0712143
R4396 VDD.n28 VDD.n27 0.0712143
R4397 VDD.n1822 VDD.n1814 0.0702959
R4398 VDD.n2005 VDD.n2003 0.0702959
R4399 VDD.n3043 VDD.n3040 0.0696837
R4400 VDD.n2395 VDD.n2393 0.0695746
R4401 VDD.n1913 VDD.n1912 0.069389
R4402 VDD.n1443 VDD.n1439 0.0693775
R4403 VDD.n185 VDD.n183 0.0693775
R4404 VDD.n1435 VDD.n1429 0.0693775
R4405 VDD.n1173 VDD.n1171 0.0693775
R4406 VDD.n1869 VDD.n1867 0.0693775
R4407 VDD.n1954 VDD.n1952 0.0693775
R4408 VDD.n171 VDD.n169 0.0693775
R4409 VDD.n2073 VDD.n2072 0.0693775
R4410 VDD.n1746 VDD.n1744 0.0684592
R4411 VDD.n2137 VDD.n2129 0.0675408
R4412 VDD.n2031 VDD.n1998 0.0675408
R4413 VDD.n309 VDD.n307 0.0666224
R4414 VDD.n1052 VDD.n1049 0.0666224
R4415 VDD.n1037 VDD.n1036 0.0666224
R4416 VDD.n2789 VDD.n2788 0.0666224
R4417 VDD.n295 VDD.n293 0.0666224
R4418 VDD.n700 VDD.n698 0.0647857
R4419 VDD.n2819 VDD.n2810 0.0647857
R4420 VDD.n2843 VDD.n2842 0.0647857
R4421 VDD.n1786 VDD.n1785 0.0638673
R4422 VDD.n1329 VDD.n1316 0.0638673
R4423 VDD.n60 VDD.n58 0.062949
R4424 VDD.n1649 VDD.n1648 0.062949
R4425 VDD.n2746 VDD.n2737 0.062949
R4426 VDD.n3087 VDD.n3085 0.0628265
R4427 VDD.n2405 VDD.n2403 0.0627854
R4428 VDD.n1914 VDD.n1913 0.0620306
R4429 VDD.n2903 VDD.n2902 0.0620306
R4430 VDD.n474 VDD.n472 0.0611122
R4431 VDD.n880 VDD.n619 0.0605319
R4432 VDD.n1897 VDD.n1895 0.0601939
R4433 VDD.n2757 VDD.n2750 0.0601939
R4434 VDD.n2967 VDD.n2965 0.0601939
R4435 VDD.n2982 VDD.n2981 0.0601939
R4436 VDD.n2648 VDD.n2646 0.0601939
R4437 VDD.n1014 VDD.n1008 0.0592755
R4438 VDD.n1512 VDD.n963 0.0592084
R4439 VDD.n3097 VDD.n3092 0.0589082
R4440 VDD.n980 VDD.n977 0.0583571
R4441 VDD.n1876 VDD.n1875 0.0583571
R4442 VDD.n2689 VDD.n2668 0.0583571
R4443 VDD.n3002 VDD.n3000 0.0583571
R4444 VDD.n3117 VDD.n3116 0.0582241
R4445 VDD.n3032 VDD.n3029 0.0579286
R4446 VDD.n1513 VDD.n1512 0.0574437
R4447 VDD.n705 VDD.n704 0.0574388
R4448 VDD.n1202 VDD.n1196 0.0574388
R4449 VDD.n2477 VDD.n2471 0.0574388
R4450 VDD.n1983 VDD.n1977 0.0574388
R4451 VDD.n1734 VDD.n1732 0.0565204
R4452 VDD.n881 VDD.n880 0.0561201
R4453 VDD.n2147 VDD.n2141 0.055602
R4454 VDD.n443 VDD.n441 0.055602
R4455 VDD.n712 VDD.n710 0.055602
R4456 VDD.n742 VDD.n740 0.055602
R4457 VDD.n1665 VDD.n1663 0.055602
R4458 VDD.n1362 VDD.n1360 0.055602
R4459 VDD.n17 VDD.n16 0.055602
R4460 VDD.n2054 VDD.n2053 0.055602
R4461 VDD.n995 VDD.n989 0.0546837
R4462 VDD.n2985 VDD.n2984 0.0546837
R4463 VDD.n2063 VDD.n2057 0.0537653
R4464 VDD.n1612 VDD.n1605 0.0537653
R4465 VDD.n2415 VDD.n2412 0.0533376
R4466 VDD.n1805 VDD.n1804 0.0528469
R4467 VDD.n1008 VDD.n1005 0.0528469
R4468 VDD.n1240 VDD.n1238 0.0528469
R4469 VDD.n861 VDD.n857 0.0519286
R4470 VDD.n867 VDD.n863 0.0519286
R4471 VDD.n1287 VDD.n1285 0.0519286
R4472 VDD.n1760 VDD.n1756 0.0519286
R4473 VDD.n2157 VDD.n2149 0.0519286
R4474 VDD.n2628 VDD.n2627 0.0510102
R4475 VDD.n783 VDD.n779 0.0500918
R4476 VDD.n793 VDD.n789 0.0500918
R4477 VDD.n2451 VDD.n2446 0.0500918
R4478 VDD.n2632 VDD.n2630 0.049618
R4479 VDD.n1365 VDD.n1363 0.0491735
R4480 VDD.n1500 VDD.n1496 0.0491735
R4481 VDD.n684 VDD.n682 0.0491735
R4482 VDD.n1492 VDD.n1486 0.0491735
R4483 VDD.n1028 VDD.n1027 0.0491735
R4484 VDD.n2378 VDD.n2375 0.0491106
R4485 VDD.n1836 VDD.n1835 0.0482551
R4486 VDD.n1426 VDD.n1422 0.0473367
R4487 VDD.n1416 VDD.n1410 0.0473367
R4488 VDD.n1187 VDD.n1185 0.0473367
R4489 VDD.n1208 VDD.n1207 0.0473367
R4490 VDD.n1302 VDD.n1301 0.0473367
R4491 VDD.n1968 VDD.n1966 0.0473367
R4492 VDD.n1989 VDD.n1988 0.0473367
R4493 VDD.n3067 VDD.n3064 0.0471531
R4494 VDD.n2425 VDD.n2422 0.0465484
R4495 VDD.n841 VDD.n832 0.0464184
R4496 VDD.n851 VDD.n847 0.0464184
R4497 VDD.n1295 VDD.n1289 0.0464184
R4498 VDD.n1754 VDD.n1752 0.0464184
R4499 VDD.n3020 VDD.n3017 0.0461735
R4500 VDD.n513 VDD.n503 0.0455
R4501 VDD.n1698 VDD.n1696 0.0455
R4502 VDD.n2043 VDD.n2039 0.0445816
R4503 VDD.n2808 VDD.n2807 0.0445816
R4504 VDD.n1643 VDD.n1641 0.0436633
R4505 VDD.n2722 VDD.n2719 0.0436633
R4506 VDD.n2961 VDD.n2959 0.0436633
R4507 VDD.n2021 VDD.n2019 0.0436633
R4508 VDD.n2126 VDD.n2122 0.0427449
R4509 VDD.n1785 VDD.n1782 0.0427449
R4510 VDD.n1264 VDD.n1262 0.0427449
R4511 VDD.n2842 VDD.n2840 0.0427449
R4512 VDD.n1701 VDD.n1668 0.0427449
R4513 VDD.n2808 VDD.n2800 0.0427449
R4514 VDD.n2590 VDD.n2589 0.0427449
R4515 VDD.n2372 VDD.n2371 0.0427449
R4516 VDD.n1301 VDD.n1299 0.0427449
R4517 VDD.n1084 VDD.n1082 0.0427449
R4518 VDD.n1126 VDD.n1124 0.0427449
R4519 VDD.n1875 VDD.n1873 0.0427449
R4520 VDD.n1740 VDD.n1738 0.0427449
R4521 VDD.n2855 VDD.n2853 0.0427449
R4522 VDD.n3004 VDD.n3002 0.0427449
R4523 VDD.n46 VDD.n43 0.0418265
R4524 VDD.n1595 VDD.n60 0.0418265
R4525 VDD.n619 VDD.n309 0.0418265
R4526 VDD.n963 VDD.n185 0.0418265
R4527 VDD.n537 VDD.n416 0.0418265
R4528 VDD.n881 VDD.n295 0.0418265
R4529 VDD.n1513 VDD.n171 0.0418265
R4530 VDD.n2157 VDD.n2156 0.0418265
R4531 VDD.n2927 VDD.n2924 0.0412755
R4532 VDD.n3010 VDD.n2427 0.0411849
R4533 VDD.n1644 VDD.n1643 0.0409082
R4534 VDD.n536 VDD.n530 0.0408433
R4535 VDD.n3049 VDD.n3046 0.0407857
R4536 VDD.n2921 VDD.n2606 0.040774
R4537 VDD.n2309 VDD.n2306 0.0404057
R4538 VDD.n2306 VDD.n2303 0.0404057
R4539 VDD.n2303 VDD.n2300 0.0404057
R4540 VDD.n1302 VDD.n1226 0.0399898
R4541 VDD.n1612 VDD.n1611 0.0399898
R4542 VDD.n2612 VDD.n2610 0.0391301
R4543 VDD.n2442 VDD.n2439 0.0391301
R4544 VDD.n483 VDD.n480 0.0390714
R4545 VDD.n2921 VDD.n2628 0.03875
R4546 VDD.n2920 VDD.n2689 0.03875
R4547 VDD.n3057 VDD.n3056 0.0386429
R4548 VDD.n682 VDD.n681 0.0381531
R4549 VDD.n1907 VDD.n1904 0.0381531
R4550 VDD.n1904 VDD.n1900 0.0381531
R4551 VDD.n1028 VDD.n1024 0.0381531
R4552 VDD.n2776 VDD.n2775 0.0381531
R4553 VDD.n2973 VDD.n2969 0.0381531
R4554 VDD.n2975 VDD.n2973 0.0381531
R4555 VDD.n19 VDD.n17 0.0381531
R4556 VDD.n2054 VDD.n2047 0.0381531
R4557 VDD.n3010 VDD.n3009 0.0377857
R4558 VDD.n480 VDD.n476 0.0372347
R4559 VDD.n2312 VDD.n2309 0.0365357
R4560 VDD.n2628 VDD.n2619 0.0363163
R4561 VDD.n2170 VDD.n46 0.035398
R4562 VDD.n1646 VDD.n1644 0.035398
R4563 VDD.n2489 VDD.n2483 0.035398
R4564 VDD.n1923 VDD.n1922 0.0352439
R4565 VDD.n1005 VDD.n998 0.0344796
R4566 VDD.n1238 VDD.n1237 0.0344796
R4567 VDD.n3115 VDD.n3112 0.0344179
R4568 VDD.n3068 VDD.n2385 0.0337877
R4569 VDD.n2126 VDD.n2120 0.0335612
R4570 VDD.n1701 VDD.n1700 0.0335612
R4571 VDD.n2665 VDD.n2662 0.0335151
R4572 VDD.n3021 VDD.n3012 0.0335
R4573 VDD.n2920 VDD.n2665 0.0333767
R4574 VDD.n2987 VDD.n2985 0.0326429
R4575 VDD.n3068 VDD.n3059 0.0326429
R4576 VDD.n3021 VDD.n2417 0.0321438
R4577 VDD.n2043 VDD.n2037 0.0317245
R4578 VDD.n441 VDD.n440 0.0317245
R4579 VDD.n710 VDD.n709 0.0317245
R4580 VDD.n740 VDD.n739 0.0317245
R4581 VDD.n1207 VDD.n1206 0.0317245
R4582 VDD.n1988 VDD.n1987 0.0317245
R4583 VDD.n1360 VDD.n1359 0.0317245
R4584 VDD.n1732 VDD.n1731 0.0308061
R4585 VDD.n841 VDD.n837 0.0298878
R4586 VDD.n707 VDD.n705 0.0298878
R4587 VDD.n851 VDD.n845 0.0298878
R4588 VDD.n1204 VDD.n1202 0.0298878
R4589 VDD.n1297 VDD.n1295 0.0298878
R4590 VDD.n1752 VDD.n1748 0.0298878
R4591 VDD.n1985 VDD.n1983 0.0298878
R4592 VDD.n1996 VDD.n1993 0.0298878
R4593 VDD.n1426 VDD.n1418 0.0289694
R4594 VDD.n1416 VDD.n1412 0.0289694
R4595 VDD.n1185 VDD.n1175 0.0289694
R4596 VDD.n1194 VDD.n1190 0.0289694
R4597 VDD.n986 VDD.n983 0.0289694
R4598 VDD.n980 VDD.n979 0.0289694
R4599 VDD.n2689 VDD.n2688 0.0289694
R4600 VDD.n1966 VDD.n1956 0.0289694
R4601 VDD.n1975 VDD.n1971 0.0289694
R4602 VDD.n3044 VDD.n3043 0.0283571
R4603 VDD.n763 VDD.n759 0.028051
R4604 VDD.n772 VDD.n768 0.028051
R4605 VDD.n3057 VDD.n2395 0.0276233
R4606 VDD.n1480 VDD.n1476 0.0271327
R4607 VDD.n1472 VDD.n1468 0.0271327
R4608 VDD.n1363 VDD.n1362 0.0271327
R4609 VDD.n1492 VDD.n1491 0.0271327
R4610 VDD.n2646 VDD.n2645 0.0271327
R4611 VDD.n3116 VDD.n2215 0.0268793
R4612 VDD.n783 VDD.n775 0.0262143
R4613 VDD.n720 VDD.n714 0.0262143
R4614 VDD.n793 VDD.n785 0.0262143
R4615 VDD.n753 VDD.n749 0.0262143
R4616 VDD.n1921 VDD.n1920 0.0262143
R4617 VDD.n2137 VDD.n2136 0.0262143
R4618 VDD.n2031 VDD.n2030 0.0262143
R4619 VDD.n1405 VDD.n1401 0.0252959
R4620 VDD.n1397 VDD.n1393 0.0252959
R4621 VDD.n1196 VDD.n1194 0.0252959
R4622 VDD.n1977 VDD.n1975 0.0252959
R4623 VDD.n3033 VDD.n2407 0.0251575
R4624 VDD.n861 VDD.n854 0.0243775
R4625 VDD.n1285 VDD.n1281 0.0243775
R4626 VDD.n1762 VDD.n1760 0.0243775
R4627 VDD.n2746 VDD.n2745 0.0243775
R4628 VDD.n2073 VDD.n2068 0.0243775
R4629 VDD.n2367 VDD.n2365 0.0238702
R4630 VDD.n2365 VDD.n2362 0.0238702
R4631 VDD.n2362 VDD.n2359 0.0238702
R4632 VDD.n2359 VDD.n2356 0.0238702
R4633 VDD.n2356 VDD.n2353 0.0238702
R4634 VDD.n2353 VDD.n2350 0.0238702
R4635 VDD.n2350 VDD.n2347 0.0238702
R4636 VDD.n2347 VDD.n2344 0.0238702
R4637 VDD.n2334 VDD.n2331 0.0238702
R4638 VDD.n2331 VDD.n2328 0.0238702
R4639 VDD.n2328 VDD.n2325 0.0238702
R4640 VDD.n2321 VDD.n2318 0.0238702
R4641 VDD.n2318 VDD.n2315 0.0238702
R4642 VDD.n2315 VDD.n2312 0.0238702
R4643 VDD.n1371 VDD.n1365 0.0234592
R4644 VDD.n1215 VDD.n1212 0.0234592
R4645 VDD.n1805 VDD.n1789 0.0234592
R4646 VDD.n1789 VDD.n1786 0.0234592
R4647 VDD.n2843 VDD.n2822 0.0234592
R4648 VDD.n3033 VDD.n3024 0.0232143
R4649 VDD.n2325 VDD.n2322 0.0231243
R4650 VDD.n2063 VDD.n2059 0.0225408
R4651 VDD.n698 VDD.n697 0.0225408
R4652 VDD.n1190 VDD.n1189 0.0225408
R4653 VDD.n2819 VDD.n2818 0.0225408
R4654 VDD.n1971 VDD.n1970 0.0225408
R4655 VDD.n30 VDD.n28 0.0225408
R4656 VDD.n3098 VDD.n3087 0.0223571
R4657 VDD.n998 VDD.n995 0.0216225
R4658 VDD.n2147 VDD.n2143 0.0207041
R4659 VDD.n1014 VDD.n969 0.0207041
R4660 VDD.n1049 VDD.n1048 0.0207041
R4661 VDD.n1663 VDD.n1659 0.0207041
R4662 VDD.n2789 VDD.n2781 0.0207041
R4663 VDD.n3044 VDD.n2405 0.020637
R4664 VDD.n2300 VDD.n2297 0.0204528
R4665 VDD.n3108 VDD.n3100 0.0193235
R4666 VDD.n3077 VDD.n3074 0.0193235
R4667 VDD.n3044 VDD.n2398 0.0189932
R4668 VDD.n3098 VDD.n3097 0.0189286
R4669 VDD.n453 VDD.n451 0.0188673
R4670 VDD.n2900 VDD.n2897 0.0186539
R4671 VDD.n3100 VDD.n3098 0.0185392
R4672 VDD.n3033 VDD.n3032 0.0180714
R4673 VDD.n1878 VDD.n1876 0.017949
R4674 VDD.n1867 VDD.n1866 0.017949
R4675 VDD.n3000 VDD.n2996 0.017949
R4676 VDD.n542 VDD.n539 0.017488
R4677 VDD.n549 VDD.n546 0.017488
R4678 VDD.n556 VDD.n553 0.017488
R4679 VDD.n559 VDD.n556 0.017488
R4680 VDD.n562 VDD.n559 0.017488
R4681 VDD.n569 VDD.n566 0.017488
R4682 VDD.n572 VDD.n569 0.017488
R4683 VDD.n579 VDD.n576 0.017488
R4684 VDD.n582 VDD.n579 0.017488
R4685 VDD.n589 VDD.n586 0.017488
R4686 VDD.n592 VDD.n589 0.017488
R4687 VDD.n595 VDD.n592 0.017488
R4688 VDD.n602 VDD.n599 0.017488
R4689 VDD.n605 VDD.n602 0.017488
R4690 VDD.n612 VDD.n609 0.017488
R4691 VDD.n618 VDD.n616 0.017488
R4692 VDD.n886 VDD.n883 0.017488
R4693 VDD.n893 VDD.n890 0.017488
R4694 VDD.n900 VDD.n897 0.017488
R4695 VDD.n903 VDD.n900 0.017488
R4696 VDD.n906 VDD.n903 0.017488
R4697 VDD.n913 VDD.n910 0.017488
R4698 VDD.n916 VDD.n913 0.017488
R4699 VDD.n923 VDD.n920 0.017488
R4700 VDD.n926 VDD.n923 0.017488
R4701 VDD.n933 VDD.n930 0.017488
R4702 VDD.n936 VDD.n933 0.017488
R4703 VDD.n939 VDD.n936 0.017488
R4704 VDD.n946 VDD.n943 0.017488
R4705 VDD.n949 VDD.n946 0.017488
R4706 VDD.n956 VDD.n953 0.017488
R4707 VDD.n962 VDD.n960 0.017488
R4708 VDD.n1518 VDD.n1515 0.017488
R4709 VDD.n1525 VDD.n1522 0.017488
R4710 VDD.n1532 VDD.n1529 0.017488
R4711 VDD.n1535 VDD.n1532 0.017488
R4712 VDD.n1538 VDD.n1535 0.017488
R4713 VDD.n1545 VDD.n1542 0.017488
R4714 VDD.n1548 VDD.n1545 0.017488
R4715 VDD.n1555 VDD.n1552 0.017488
R4716 VDD.n1558 VDD.n1555 0.017488
R4717 VDD.n1565 VDD.n1562 0.017488
R4718 VDD.n1568 VDD.n1565 0.017488
R4719 VDD.n1571 VDD.n1568 0.017488
R4720 VDD.n1578 VDD.n1575 0.017488
R4721 VDD.n1581 VDD.n1578 0.017488
R4722 VDD.n1588 VDD.n1585 0.017488
R4723 VDD.n1594 VDD.n1592 0.017488
R4724 VDD.n3109 VDD.n3108 0.0171667
R4725 VDD.n566 VDD.n563 0.0169458
R4726 VDD.n910 VDD.n907 0.0169458
R4727 VDD.n1542 VDD.n1539 0.0169458
R4728 VDD.n543 VDD.n542 0.0165843
R4729 VDD.n887 VDD.n886 0.0165843
R4730 VDD.n1519 VDD.n1518 0.0165843
R4731 VDD.n1895 VDD.n1891 0.0161122
R4732 VDD.n1056 VDD.n1052 0.0161122
R4733 VDD.n2797 VDD.n2796 0.0161122
R4734 VDD.n2757 VDD.n2756 0.0161122
R4735 VDD.n2965 VDD.n2961 0.0161122
R4736 VDD.n2984 VDD.n2982 0.0161122
R4737 VDD.n3112 VDD.n3109 0.0156119
R4738 VDD.n3116 VDD.n3115 0.0152761
R4739 VDD.n472 VDD.n466 0.0151939
R4740 VDD.n1267 VDD.n1265 0.0151939
R4741 VDD.n1780 VDD.n1779 0.0151939
R4742 VDD.n2341 VDD.n2334 0.0151685
R4743 VDD.n583 VDD.n582 0.0149578
R4744 VDD.n927 VDD.n926 0.0149578
R4745 VDD.n1559 VDD.n1558 0.0149578
R4746 VDD.n2176 VDD.n2173 0.0147031
R4747 VDD.n2188 VDD.n2185 0.0147031
R4748 VDD.n3033 VDD.n2415 0.0144726
R4749 VDD.n2195 VDD.n2192 0.014
R4750 VDD.n2179 VDD.n2176 0.0137188
R4751 VDD.n2182 VDD.n2179 0.0137188
R4752 VDD.n2185 VDD.n2182 0.0137188
R4753 VDD.n2198 VDD.n2195 0.0137188
R4754 VDD.n3130 VDD.n3127 0.0137188
R4755 VDD.n3123 VDD.n3120 0.0137188
R4756 VDD.n58 VDD.n50 0.0133571
R4757 VDD.n451 VDD.n450 0.0133571
R4758 VDD.n691 VDD.n689 0.0133571
R4759 VDD.n1651 VDD.n1649 0.0133571
R4760 VDD.n2501 VDD.n2495 0.0133571
R4761 VDD.n599 VDD.n596 0.0131506
R4762 VDD.n943 VDD.n940 0.0131506
R4763 VDD.n1575 VDD.n1572 0.0131506
R4764 VDD.n3044 VDD.n3036 0.0129286
R4765 VDD.n1329 VDD.n1306 0.0124388
R4766 VDD.n2114 VDD.n2113 0.0124388
R4767 VDD VDD.n3130 0.0121719
R4768 VDD.n3057 VDD.n2388 0.0120068
R4769 VDD.n606 VDD.n605 0.0117048
R4770 VDD.n950 VDD.n949 0.0117048
R4771 VDD.n1582 VDD.n1581 0.0117048
R4772 VDD.n2102 VDD.n2098 0.0115204
R4773 VDD.n1253 VDD.n1251 0.0115204
R4774 VDD.n550 VDD.n549 0.0113434
R4775 VDD.n616 VDD.n613 0.0113434
R4776 VDD.n894 VDD.n893 0.0113434
R4777 VDD.n960 VDD.n957 0.0113434
R4778 VDD.n1526 VDD.n1525 0.0113434
R4779 VDD.n1592 VDD.n1589 0.0113434
R4780 VDD.n2189 VDD.n2188 0.0111875
R4781 VDD.n2903 VDD.n2900 0.0110413
R4782 VDD.n1917 VDD.n1914 0.010602
R4783 VDD.n1355 VDD.n1354 0.010602
R4784 VDD.n576 VDD.n573 0.0100783
R4785 VDD.n920 VDD.n917 0.0100783
R4786 VDD.n1552 VDD.n1549 0.0100783
R4787 VDD.n1603 VDD.n1599 0.00968367
R4788 VDD.n307 VDD.n300 0.00968367
R4789 VDD.n293 VDD.n287 0.00968367
R4790 VDD.n3124 VDD.n3123 0.00964062
R4791 VDD.n1924 VDD.n1923 0.00956098
R4792 VDD.n2344 VDD.n2341 0.00920166
R4793 VDD.n1371 VDD.n1367 0.00876531
R4794 VDD.n1215 VDD.n1135 0.00876531
R4795 VDD.n1210 VDD.n1208 0.00876531
R4796 VDD.n1313 VDD.n1310 0.00876531
R4797 VDD.n1260 VDD.n1259 0.00876531
R4798 VDD.n1862 VDD.n1860 0.00876531
R4799 VDD.n1991 VDD.n1989 0.00876531
R4800 VDD.n2092 VDD.n2086 0.00876531
R4801 VDD.n3068 VDD.n3067 0.00864286
R4802 VDD.n2173 VDD.n2170 0.008375
R4803 VDD.n573 VDD.n572 0.00790964
R4804 VDD.n917 VDD.n916 0.00790964
R4805 VDD.n1549 VDD.n1548 0.00790964
R4806 VDD.n820 VDD.n816 0.00784694
R4807 VDD.n829 VDD.n825 0.00784694
R4808 VDD.n1744 VDD.n1740 0.00784694
R4809 VDD.n3021 VDD.n3020 0.00778571
R4810 VDD.n3120 VDD.n3117 0.00767187
R4811 VDD.n3021 VDD.n2425 0.0074863
R4812 VDD.n1443 VDD.n1437 0.00692857
R4813 VDD.n169 VDD.n162 0.00692857
R4814 VDD.n1435 VDD.n1431 0.00692857
R4815 VDD.n1171 VDD.n1161 0.00692857
R4816 VDD.n1714 VDD.n1713 0.00692857
R4817 VDD.n183 VDD.n175 0.00692857
R4818 VDD.n553 VDD.n550 0.00664458
R4819 VDD.n613 VDD.n612 0.00664458
R4820 VDD.n897 VDD.n894 0.00664458
R4821 VDD.n957 VDD.n956 0.00664458
R4822 VDD.n1529 VDD.n1526 0.00664458
R4823 VDD.n1589 VDD.n1588 0.00664458
R4824 VDD.n609 VDD.n606 0.00628313
R4825 VDD.n953 VDD.n950 0.00628313
R4826 VDD.n1585 VDD.n1582 0.00628313
R4827 VDD.n2920 VDD.n2632 0.00625342
R4828 VDD.n627 VDD.n623 0.0060102
R4829 VDD.n720 VDD.n716 0.0060102
R4830 VDD.n636 VDD.n632 0.0060102
R4831 VDD.n753 VDD.n723 0.0060102
R4832 VDD.n1822 VDD.n1808 0.0060102
R4833 VDD.n3068 VDD.n2378 0.00584247
R4834 VDD.n1462 VDD.n1458 0.00509184
R4835 VDD.n157 VDD.n155 0.00509184
R4836 VDD.n446 VDD.n445 0.00509184
R4837 VDD.n1453 VDD.n1449 0.00509184
R4838 VDD.n745 VDD.n744 0.00509184
R4839 VDD.n1727 VDD.n1726 0.00509184
R4840 VDD.n1509 VDD.n1508 0.00509184
R4841 VDD.n596 VDD.n595 0.00483735
R4842 VDD.n940 VDD.n939 0.00483735
R4843 VDD.n1572 VDD.n1571 0.00483735
R4844 VDD.n3127 VDD.n3124 0.00457813
R4845 VDD.n802 VDD.n796 0.00417347
R4846 VDD.n810 VDD.n806 0.00417347
R4847 VDD.n3010 VDD.n2927 0.0035
R4848 VDD.n1388 VDD.n1384 0.0032551
R4849 VDD.n675 VDD.n674 0.0032551
R4850 VDD.n1380 VDD.n1376 0.0032551
R4851 VDD.n1157 VDD.n1156 0.0032551
R4852 VDD.n2979 VDD.n2975 0.0032551
R4853 VDD.n1352 VDD.n1350 0.0032551
R4854 VDD.n2192 VDD.n2189 0.00303125
R4855 VDD VDD.n2198 0.00303125
R4856 VDD.n586 VDD.n583 0.00303012
R4857 VDD.n930 VDD.n927 0.00303012
R4858 VDD.n1562 VDD.n1559 0.00303012
R4859 VDD.n3057 VDD.n3049 0.00264286
R4860 VDD.n1996 VDD.n1930 0.00233673
R4861 VDD.n877 VDD.n870 0.00233673
R4862 VDD.n282 VDD.n280 0.00233673
R4863 VDD.n1276 VDD.n1275 0.00233673
R4864 VDD.n2768 VDD.n2767 0.00233673
R4865 VDD.n1772 VDD.n1770 0.00233673
R4866 VDD.n2297 VDD.n2296 0.00186203
R4867 VDD.n2921 VDD.n2612 0.00173288
R4868 VDD.n1127 VDD.n1067 0.00141837
R4869 VDD.n2730 VDD.n2724 0.00141837
R4870 VDD.n2959 VDD.n2958 0.00141837
R4871 VDD.n546 VDD.n543 0.00140361
R4872 VDD.n890 VDD.n887 0.00140361
R4873 VDD.n1522 VDD.n1519 0.00140361
R4874 VDD.n3010 VDD.n2442 0.00132192
R4875 VDD.n2322 VDD.n2321 0.00124586
R4876 VDD.n563 VDD.n562 0.00104217
R4877 VDD.n907 VDD.n906 0.00104217
R4878 VDD.n1539 VDD.n1538 0.00104217
R4879 VDD.n3098 VDD.n3077 0.000892157
R4880 VDD.n3074 VDD.n3072 0.000892157
R4881 VDD.n2372 VDD.n2367 0.000748619
R4882 VDD.n539 VDD.n537 0.000680723
R4883 VDD.n619 VDD.n618 0.000680723
R4884 VDD.n883 VDD.n881 0.000680723
R4885 VDD.n963 VDD.n962 0.000680723
R4886 VDD.n1515 VDD.n1513 0.000680723
R4887 VDD.n1595 VDD.n1594 0.000680723
R4888 VSS.n841 VSS.n840 33926.4
R4889 VSS.n880 VSS.n874 33926.4
R4890 VSS.n1937 VSS.n1936 13208.8
R4891 VSS.n1938 VSS.n1937 12616
R4892 VSS.n878 VSS.n875 7574.75
R4893 VSS.n879 VSS.n878 5135.34
R4894 VSS.n881 VSS.n880 4288.97
R4895 VSS.n880 VSS.n879 2442.17
R4896 VSS.n878 VSS.n877 936.442
R4897 VSS.n877 VSS.n876 328.005
R4898 VSS.n1942 VSS.n1938 216.931
R4899 VSS.n1308 VSS.n1307 121.826
R4900 VSS.n970 VSS.t116 46.7987
R4901 VSS.n976 VSS.t99 46.7987
R4902 VSS.n937 VSS.t101 46.7987
R4903 VSS.n774 VSS.t97 46.7987
R4904 VSS.n720 VSS.t108 46.7987
R4905 VSS.n718 VSS.t89 46.7987
R4906 VSS.n785 VSS.t120 46.6684
R4907 VSS.n461 VSS.t114 46.6684
R4908 VSS.n976 VSS.t110 46.0557
R4909 VSS.n937 VSS.t125 46.0557
R4910 VSS.n774 VSS.t83 46.0557
R4911 VSS.n718 VSS.t127 46.0557
R4912 VSS.n1765 VSS.t6 31.935
R4913 VSS.n1987 VSS.t39 28.4397
R4914 VSS.n1423 VSS.t21 28.1645
R4915 VSS.n1910 VSS.t9 26.6126
R4916 VSS.n1518 VSS.t4 25.282
R4917 VSS.n1268 VSS.t122 23.9247
R4918 VSS.n1190 VSS.t16 23.5797
R4919 VSS.n208 VSS.t192 23.4
R4920 VSS.n114 VSS.t92 23.2729
R4921 VSS.n1931 VSS.t165 22.4873
R4922 VSS.n1897 VSS.t3 21.2902
R4923 VSS.n2145 VSS.t278 20.3048
R4924 VSS.n2129 VSS.t123 20.3048
R4925 VSS.n1172 VSS.t266 18.9949
R4926 VSS.n1146 VSS.t84 18.8616
R4927 VSS.n1089 VSS.t90 18.0757
R4928 VSS.n198 VSS.t182 17.0758
R4929 VSS.n1223 VSS.t62 17.0299
R4930 VSS.n1958 VSS.t153 16.5349
R4931 VSS.n1103 VSS.t49 16.5039
R4932 VSS.n1514 VSS.t129 15.9677
R4933 VSS.n1132 VSS.t31 15.7181
R4934 VSS.n1395 VSS.t23 15.065
R4935 VSS.n1231 VSS.t154 15.065
R4936 VSS.n1913 VSS.t52 14.6371
R4937 VSS.n858 VSS.t174 12.9675
R4938 VSS.n1119 VSS.t47 12.5746
R4939 VSS.n1116 VSS.t28 11.7887
R4940 VSS.n256 VSS.t176 10.7516
R4941 VSS.n174 VSS.t112 9.892
R4942 VSS.n302 VSS.t103 9.8555
R4943 VSS.n170 VSS.t105 9.7825
R4944 VSS.n304 VSS.t86 9.7825
R4945 VSS.n302 VSS.t95 9.7095
R4946 VSS.n174 VSS.t118 9.673
R4947 VSS.n1768 VSS.t55 9.31473
R4948 VSS.n868 VSS.t179 9.0381
R4949 VSS.n1136 VSS.t44 8.64516
R4950 VSS.n885 VSS.t190 8.22194
R4951 VSS.n1508 VSS.t142 7.98412
R4952 VSS.n1099 VSS.t26 7.85928
R4953 VSS.n842 VSS.t87 7.46634
R4954 VSS.n1952 VSS.t38 7.27563
R4955 VSS.n224 VSS.t106 6.95711
R4956 VSS.n1197 VSS.t13 6.55028
R4957 VSS.n1093 VSS.t41 6.28753
R4958 VSS.n1142 VSS.t33 5.50165
R4959 VSS.n117 VSS.n116 5.05985
R4960 VSS.n1406 VSS.t267 4.72519
R4961 VSS.n1922 VSS.t11 4.63013
R4962 VSS.t13 VSS.t216 4.58534
R4963 VSS.t60 VSS.t147 4.58534
R4964 VSS.t156 VSS.t0 4.58534
R4965 VSS.t62 VSS.t149 4.58534
R4966 VSS.n285 VSS.t172 4.42743
R4967 VSS.n1167 VSS.n1164 4.27059
R4968 VSS.n1240 VSS.t63 4.27059
R4969 VSS.n2162 VSS.n1461 4.25968
R4970 VSS.n2128 VSS.t150 4.25968
R4971 VSS.n971 VSS.n970 4.0005
R4972 VSS.n977 VSS.n976 4.0005
R4973 VSS.n719 VSS.n718 4.0005
R4974 VSS.n721 VSS.n720 4.0005
R4975 VSS.n462 VSS.n461 4.0005
R4976 VSS.n775 VSS.n774 4.0005
R4977 VSS.n786 VSS.n785 4.0005
R4978 VSS.n938 VSS.n937 4.0005
R4979 VSS.n113 VSS.t94 3.9695
R4980 VSS.n1267 VSS.t124 3.9695
R4981 VSS.n177 VSS.t119 3.9695
R4982 VSS.n173 VSS.t113 3.9695
R4983 VSS.n169 VSS.t107 3.9695
R4984 VSS.n326 VSS.t88 3.9695
R4985 VSS.n307 VSS.t96 3.9695
R4986 VSS.n309 VSS.t104 3.9695
R4987 VSS.n882 VSS.n881 3.92989
R4988 VSS.n1247 VSS.n1239 3.74619
R4989 VSS.n1214 VSS.n1209 3.72459
R4990 VSS.n2152 VSS.n1463 3.71368
R4991 VSS.n2138 VSS.n1974 3.71368
R4992 VSS.n940 VSS.t126 3.6965
R4993 VSS.n936 VSS.t102 3.6965
R4994 VSS.n788 VSS.t121 3.6965
R4995 VSS.n777 VSS.t85 3.6965
R4996 VSS.n773 VSS.t98 3.6965
R4997 VSS.n464 VSS.t115 3.6965
R4998 VSS.n474 VSS.n472 3.30215
R4999 VSS.n324 VSS.n323 3.30215
R5000 VSS.n86 VSS.n84 3.30215
R5001 VSS.n549 VSS.n547 3.30158
R5002 VSS.n474 VSS.n473 3.30158
R5003 VSS.n485 VSS.n484 3.30158
R5004 VSS.n493 VSS.n492 3.30158
R5005 VSS.n502 VSS.n501 3.30158
R5006 VSS.n502 VSS.n500 3.30158
R5007 VSS.n917 VSS.n916 3.30158
R5008 VSS.n106 VSS.n103 3.30158
R5009 VSS.n86 VSS.n85 3.30158
R5010 VSS.n1604 VSS.n1602 3.30147
R5011 VSS.n1622 VSS.n1620 3.30147
R5012 VSS.n1587 VSS.n1584 3.30147
R5013 VSS.n1647 VSS.n1645 3.30147
R5014 VSS.n1651 VSS.n1650 3.30147
R5015 VSS.n95 VSS.n93 3.30147
R5016 VSS.n2101 VSS.n2099 3.30147
R5017 VSS.n2093 VSS.n2091 3.30147
R5018 VSS.n2023 VSS.n2021 3.30147
R5019 VSS.n2109 VSS.n2108 3.30147
R5020 VSS.n1683 VSS.n1682 3.30147
R5021 VSS.n1310 VSS.n1306 3.30147
R5022 VSS.n1433 VSS.n1431 3.30147
R5023 VSS.n1447 VSS.n1446 3.30147
R5024 VSS.n2174 VSS.n2171 3.30147
R5025 VSS.n1299 VSS.n1297 3.30101
R5026 VSS.n1447 VSS.n1445 3.30091
R5027 VSS.n1754 VSS.n1753 3.30091
R5028 VSS.n1647 VSS.n1646 3.30091
R5029 VSS.n1622 VSS.n1621 3.30091
R5030 VSS.n1604 VSS.n1603 3.30091
R5031 VSS.n1587 VSS.n1586 3.30091
R5032 VSS.n1651 VSS.n1649 3.30091
R5033 VSS.n31 VSS.n30 3.30091
R5034 VSS.n95 VSS.n94 3.30091
R5035 VSS.n2109 VSS.n2107 3.30091
R5036 VSS.n2023 VSS.n2022 3.30091
R5037 VSS.n2093 VSS.n2092 3.30091
R5038 VSS.n2101 VSS.n2100 3.30091
R5039 VSS.n1683 VSS.n1681 3.30091
R5040 VSS.n1433 VSS.n1432 3.30091
R5041 VSS.n2174 VSS.n2173 3.30091
R5042 VSS.n2153 VSS.t151 3.27539
R5043 VSS.n2135 VSS.t156 3.27539
R5044 VSS.n1186 VSS.n1185 3.1505
R5045 VSS.n1219 VSS.n1218 3.1505
R5046 VSS.n1694 VSS.n1693 3.1505
R5047 VSS.n1773 VSS.n1772 3.1505
R5048 VSS.n1776 VSS.n1775 3.1505
R5049 VSS.n1779 VSS.n1778 3.1505
R5050 VSS.n1691 VSS.n1690 3.1505
R5051 VSS.n1497 VSS.n1496 3.1505
R5052 VSS.n1500 VSS.n1499 3.1505
R5053 VSS.n1503 VSS.n1502 3.1505
R5054 VSS.n1688 VSS.n1687 3.1505
R5055 VSS.n1488 VSS.n1487 3.1505
R5056 VSS.n1491 VSS.n1490 3.1505
R5057 VSS.n1494 VSS.n1493 3.1505
R5058 VSS.n1715 VSS.n1714 3.1505
R5059 VSS.n1782 VSS.n1781 3.1505
R5060 VSS.n1785 VSS.n1784 3.1505
R5061 VSS.n1788 VSS.n1787 3.1505
R5062 VSS.n635 VSS.n634 3.1505
R5063 VSS.n975 VSS.n974 3.1505
R5064 VSS.n981 VSS.n980 3.1505
R5065 VSS.n969 VSS.n968 3.1505
R5066 VSS.n966 VSS.n965 3.1505
R5067 VSS.n645 VSS.n644 3.1505
R5068 VSS.n249 VSS.n248 3.1505
R5069 VSS.n252 VSS.n251 3.1505
R5070 VSS.n255 VSS.n254 3.1505
R5071 VSS.n185 VSS.n184 3.1505
R5072 VSS.n188 VSS.n187 3.1505
R5073 VSS.n191 VSS.n190 3.1505
R5074 VSS.n268 VSS.n267 3.1505
R5075 VSS.n271 VSS.n270 3.1505
R5076 VSS.n274 VSS.n273 3.1505
R5077 VSS.n295 VSS.n294 3.1505
R5078 VSS.n298 VSS.n297 3.1505
R5079 VSS.n301 VSS.n300 3.1505
R5080 VSS.n381 VSS.n379 3.1505
R5081 VSS.n681 VSS.n680 3.1505
R5082 VSS.n678 VSS.n677 3.1505
R5083 VSS.n384 VSS.n383 3.1505
R5084 VSS.n555 VSS.n553 3.1505
R5085 VSS.n951 VSS.n950 3.1505
R5086 VSS.n948 VSS.n947 3.1505
R5087 VSS.n558 VSS.n557 3.1505
R5088 VSS.n687 VSS.n686 3.1505
R5089 VSS.n684 VSS.n683 3.1505
R5090 VSS.n387 VSS.n386 3.1505
R5091 VSS.n957 VSS.n956 3.1505
R5092 VSS.n954 VSS.n953 3.1505
R5093 VSS.n667 VSS.n666 3.1505
R5094 VSS.n696 VSS.n695 3.1505
R5095 VSS.n693 VSS.n692 3.1505
R5096 VSS.n390 VSS.n389 3.1505
R5097 VSS.n963 VSS.n962 3.1505
R5098 VSS.n960 VSS.n959 3.1505
R5099 VSS.n656 VSS.n655 3.1505
R5100 VSS.n705 VSS.n704 3.1505
R5101 VSS.n702 VSS.n701 3.1505
R5102 VSS.n393 VSS.n392 3.1505
R5103 VSS.n729 VSS.n728 3.1505
R5104 VSS.n396 VSS.n395 3.1505
R5105 VSS.n725 VSS.n724 3.1505
R5106 VSS.n766 VSS.n765 3.1505
R5107 VSS.n769 VSS.n768 3.1505
R5108 VSS.n942 VSS.n941 3.1505
R5109 VSS.n945 VSS.n944 3.1505
R5110 VSS.n1422 VSS.n1421 3.1505
R5111 VSS.t87 VSS.n841 3.14401
R5112 VSS.n31 VSS.n29 3.04657
R5113 VSS.n1299 VSS.n1298 3.04657
R5114 VSS.n549 VSS.n548 2.99152
R5115 VSS.n106 VSS.n105 2.99146
R5116 VSS.n1754 VSS.n1752 2.99137
R5117 VSS.n1310 VSS.n1309 2.9908
R5118 VSS.n279 VSS.n276 2.79116
R5119 VSS.n552 VSS.n551 2.79049
R5120 VSS.n287 VSS.n284 2.79049
R5121 VSS.n1903 VSS.t57 2.66171
R5122 VSS.n1288 VSS.n1271 2.60143
R5123 VSS.n1533 VSS.n1485 2.60143
R5124 VSS.n369 VSS.n368 2.60143
R5125 VSS.n1341 VSS.n1340 2.60143
R5126 VSS.n1750 VSS.n1685 2.60142
R5127 VSS.n1888 VSS.n1887 2.6005
R5128 VSS.n1863 VSS.n1862 2.6005
R5129 VSS.n1860 VSS.n1859 2.6005
R5130 VSS.n1857 VSS.n1856 2.6005
R5131 VSS.n1854 VSS.n1853 2.6005
R5132 VSS.n1851 VSS.n1850 2.6005
R5133 VSS.n1848 VSS.n1847 2.6005
R5134 VSS.n1845 VSS.n1844 2.6005
R5135 VSS.n1842 VSS.n1841 2.6005
R5136 VSS.n1839 VSS.n1838 2.6005
R5137 VSS.n1836 VSS.n1835 2.6005
R5138 VSS.n1833 VSS.n1832 2.6005
R5139 VSS.n1830 VSS.n1829 2.6005
R5140 VSS.n1827 VSS.n1826 2.6005
R5141 VSS.n1824 VSS.n1823 2.6005
R5142 VSS.n1822 VSS.n1821 2.6005
R5143 VSS.n1820 VSS.n1819 2.6005
R5144 VSS.n1818 VSS.n1817 2.6005
R5145 VSS.n1816 VSS.n1815 2.6005
R5146 VSS.n1814 VSS.n1813 2.6005
R5147 VSS.n1812 VSS.n1811 2.6005
R5148 VSS.n1810 VSS.n1809 2.6005
R5149 VSS.n1808 VSS.n1807 2.6005
R5150 VSS.n1806 VSS.n1805 2.6005
R5151 VSS.n1804 VSS.n1803 2.6005
R5152 VSS.n1802 VSS.n1801 2.6005
R5153 VSS.n1800 VSS.n1799 2.6005
R5154 VSS.n1798 VSS.n1797 2.6005
R5155 VSS.n1796 VSS.n1795 2.6005
R5156 VSS.n1794 VSS.n1793 2.6005
R5157 VSS.n1792 VSS.n1791 2.6005
R5158 VSS.n1790 VSS.n1789 2.6005
R5159 VSS.n1696 VSS.n1695 2.6005
R5160 VSS.n1698 VSS.n1697 2.6005
R5161 VSS.n1700 VSS.n1699 2.6005
R5162 VSS.n1532 VSS.n1531 2.6005
R5163 VSS.n1531 VSS.n1530 2.6005
R5164 VSS.n1626 VSS.n1625 2.6005
R5165 VSS.n1628 VSS.n1627 2.6005
R5166 VSS.n1606 VSS.n1605 2.6005
R5167 VSS.n1608 VSS.n1607 2.6005
R5168 VSS.n1589 VSS.n1588 2.6005
R5169 VSS.n1592 VSS.n1591 2.6005
R5170 VSS.n1568 VSS.n1567 2.6005
R5171 VSS.n1571 VSS.n1570 2.6005
R5172 VSS.n1574 VSS.n1566 2.6005
R5173 VSS.n1574 VSS.n1573 2.6005
R5174 VSS.n1549 VSS.n1548 2.6005
R5175 VSS.n1552 VSS.n1551 2.6005
R5176 VSS.n1555 VSS.n1547 2.6005
R5177 VSS.n1555 VSS.n1554 2.6005
R5178 VSS.n1481 VSS.n1480 2.6005
R5179 VSS.n1484 VSS.n1483 2.6005
R5180 VSS.n1536 VSS.n1479 2.6005
R5181 VSS.n1536 VSS.n1535 2.6005
R5182 VSS.n1624 VSS.n1623 2.6005
R5183 VSS.n1653 VSS.n1652 2.6005
R5184 VSS.n1655 VSS.n1654 2.6005
R5185 VSS.n1641 VSS.n1640 2.6005
R5186 VSS.n1643 VSS.n1642 2.6005
R5187 VSS.n1702 VSS.n1701 2.6005
R5188 VSS.n1749 VSS.n1748 2.6005
R5189 VSS.n1747 VSS.n1746 2.6005
R5190 VSS.n1745 VSS.n1744 2.6005
R5191 VSS.n1743 VSS.n1742 2.6005
R5192 VSS.n1741 VSS.n1740 2.6005
R5193 VSS.n1738 VSS.n1737 2.6005
R5194 VSS.n1736 VSS.n1735 2.6005
R5195 VSS.n1734 VSS.n1733 2.6005
R5196 VSS.n1731 VSS.n1730 2.6005
R5197 VSS.n1729 VSS.n1728 2.6005
R5198 VSS.n1727 VSS.n1726 2.6005
R5199 VSS.n1724 VSS.n1723 2.6005
R5200 VSS.n1722 VSS.n1721 2.6005
R5201 VSS.n1720 VSS.n1719 2.6005
R5202 VSS.n1718 VSS.n1717 2.6005
R5203 VSS.n1712 VSS.n1711 2.6005
R5204 VSS.n1710 VSS.n1709 2.6005
R5205 VSS.n1708 VSS.n1707 2.6005
R5206 VSS.n1706 VSS.n1705 2.6005
R5207 VSS.n1704 VSS.n1703 2.6005
R5208 VSS.n1890 VSS.n1889 2.6005
R5209 VSS.n1893 VSS.n1892 2.6005
R5210 VSS.n1892 VSS.n1891 2.6005
R5211 VSS.n1896 VSS.n1895 2.6005
R5212 VSS.n1895 VSS.n1894 2.6005
R5213 VSS.n1899 VSS.n1898 2.6005
R5214 VSS.n1898 VSS.n1897 2.6005
R5215 VSS.n1902 VSS.n1901 2.6005
R5216 VSS.n1901 VSS.n1900 2.6005
R5217 VSS.n1905 VSS.n1904 2.6005
R5218 VSS.n1904 VSS.n1903 2.6005
R5219 VSS.n1909 VSS.n1908 2.6005
R5220 VSS.n1908 VSS.n1907 2.6005
R5221 VSS.n1912 VSS.n1911 2.6005
R5222 VSS.n1911 VSS.n1910 2.6005
R5223 VSS.n1915 VSS.n1914 2.6005
R5224 VSS.n1914 VSS.n1913 2.6005
R5225 VSS.n1918 VSS.n1917 2.6005
R5226 VSS.n1917 VSS.n1916 2.6005
R5227 VSS.n1770 VSS.n1769 2.6005
R5228 VSS.n1769 VSS.n1768 2.6005
R5229 VSS.n1767 VSS.n1766 2.6005
R5230 VSS.n1766 VSS.n1765 2.6005
R5231 VSS.n1506 VSS.n1505 2.6005
R5232 VSS.n1505 VSS.n1504 2.6005
R5233 VSS.n1510 VSS.n1509 2.6005
R5234 VSS.n1509 VSS.n1508 2.6005
R5235 VSS.n1513 VSS.n1512 2.6005
R5236 VSS.n1512 VSS.n1511 2.6005
R5237 VSS.n1516 VSS.n1515 2.6005
R5238 VSS.n1515 VSS.n1514 2.6005
R5239 VSS.n1520 VSS.n1519 2.6005
R5240 VSS.n1519 VSS.n1518 2.6005
R5241 VSS.n1523 VSS.n1522 2.6005
R5242 VSS.n1522 VSS.n1521 2.6005
R5243 VSS.n1526 VSS.n1525 2.6005
R5244 VSS.n1525 VSS.n1524 2.6005
R5245 VSS.n1529 VSS.n1528 2.6005
R5246 VSS.n1528 VSS.n1527 2.6005
R5247 VSS.n410 VSS.n409 2.6005
R5248 VSS.n538 VSS.n535 2.6005
R5249 VSS.n623 VSS.n580 2.6005
R5250 VSS.n661 VSS.n660 2.6005
R5251 VSS.n573 VSS.n560 2.6005
R5252 VSS.n1080 VSS.n1079 2.6005
R5253 VSS.n1034 VSS.n1033 2.6005
R5254 VSS.n1031 VSS.n1030 2.6005
R5255 VSS.n1028 VSS.n1027 2.6005
R5256 VSS.n1025 VSS.n1024 2.6005
R5257 VSS.n1022 VSS.n1021 2.6005
R5258 VSS.n1019 VSS.n1018 2.6005
R5259 VSS.n1016 VSS.n1015 2.6005
R5260 VSS.n1013 VSS.n1012 2.6005
R5261 VSS.n1010 VSS.n1009 2.6005
R5262 VSS.n1007 VSS.n1006 2.6005
R5263 VSS.n1005 VSS.n1004 2.6005
R5264 VSS.n1003 VSS.n1002 2.6005
R5265 VSS.n1001 VSS.n1000 2.6005
R5266 VSS.n999 VSS.n998 2.6005
R5267 VSS.n997 VSS.n996 2.6005
R5268 VSS.n995 VSS.n994 2.6005
R5269 VSS.n993 VSS.n992 2.6005
R5270 VSS.n991 VSS.n990 2.6005
R5271 VSS.n989 VSS.n988 2.6005
R5272 VSS.n562 VSS.n561 2.6005
R5273 VSS.n564 VSS.n563 2.6005
R5274 VSS.n566 VSS.n565 2.6005
R5275 VSS.n568 VSS.n567 2.6005
R5276 VSS.n570 VSS.n569 2.6005
R5277 VSS.n572 VSS.n571 2.6005
R5278 VSS.n575 VSS.n574 2.6005
R5279 VSS.n578 VSS.n577 2.6005
R5280 VSS.n630 VSS.n629 2.6005
R5281 VSS.n632 VSS.n631 2.6005
R5282 VSS.n638 VSS.n637 2.6005
R5283 VSS.n648 VSS.n647 2.6005
R5284 VSS.n650 VSS.n649 2.6005
R5285 VSS.n659 VSS.n658 2.6005
R5286 VSS.n670 VSS.n669 2.6005
R5287 VSS.n672 VSS.n671 2.6005
R5288 VSS.n675 VSS.n674 2.6005
R5289 VSS.n755 VSS.n754 2.6005
R5290 VSS.n757 VSS.n756 2.6005
R5291 VSS.n760 VSS.n759 2.6005
R5292 VSS.n790 VSS.n550 2.6005
R5293 VSS.n315 VSS.n314 2.6005
R5294 VSS.n900 VSS.n899 2.6005
R5295 VSS.n902 VSS.n901 2.6005
R5296 VSS.n906 VSS.n905 2.6005
R5297 VSS.n897 VSS.n896 2.6005
R5298 VSS.n927 VSS.n926 2.6005
R5299 VSS.n924 VSS.n923 2.6005
R5300 VSS.n525 VSS.n524 2.6005
R5301 VSS.n504 VSS.n503 2.6005
R5302 VSS.n490 VSS.n489 2.6005
R5303 VSS.n480 VSS.n479 2.6005
R5304 VSS.n476 VSS.n475 2.6005
R5305 VSS.n478 VSS.n477 2.6005
R5306 VSS.n487 VSS.n486 2.6005
R5307 VSS.n482 VSS.n481 2.6005
R5308 VSS.n495 VSS.n494 2.6005
R5309 VSS.n499 VSS.n498 2.6005
R5310 VSS.n506 VSS.n505 2.6005
R5311 VSS.n509 VSS.n508 2.6005
R5312 VSS.n511 VSS.n510 2.6005
R5313 VSS.n367 VSS.n366 2.6005
R5314 VSS.n364 VSS.n363 2.6005
R5315 VSS.n362 VSS.n361 2.6005
R5316 VSS.n360 VSS.n359 2.6005
R5317 VSS.n357 VSS.n356 2.6005
R5318 VSS.n355 VSS.n354 2.6005
R5319 VSS.n353 VSS.n352 2.6005
R5320 VSS.n351 VSS.n350 2.6005
R5321 VSS.n349 VSS.n348 2.6005
R5322 VSS.n346 VSS.n345 2.6005
R5323 VSS.n344 VSS.n343 2.6005
R5324 VSS.n342 VSS.n341 2.6005
R5325 VSS.n340 VSS.n339 2.6005
R5326 VSS.n372 VSS.n371 2.6005
R5327 VSS.n519 VSS.n518 2.6005
R5328 VSS.n377 VSS.n376 2.6005
R5329 VSS.n516 VSS.n515 2.6005
R5330 VSS.n513 VSS.n512 2.6005
R5331 VSS.n522 VSS.n521 2.6005
R5332 VSS.n531 VSS.n530 2.6005
R5333 VSS.n375 VSS.n374 2.6005
R5334 VSS.n534 VSS.n533 2.6005
R5335 VSS.n471 VSS.n470 2.6005
R5336 VSS.n622 VSS.n621 2.6005
R5337 VSS.n620 VSS.n619 2.6005
R5338 VSS.n618 VSS.n617 2.6005
R5339 VSS.n616 VSS.n615 2.6005
R5340 VSS.n614 VSS.n613 2.6005
R5341 VSS.n612 VSS.n611 2.6005
R5342 VSS.n610 VSS.n609 2.6005
R5343 VSS.n608 VSS.n607 2.6005
R5344 VSS.n606 VSS.n605 2.6005
R5345 VSS.n604 VSS.n603 2.6005
R5346 VSS.n602 VSS.n601 2.6005
R5347 VSS.n600 VSS.n599 2.6005
R5348 VSS.n598 VSS.n597 2.6005
R5349 VSS.n596 VSS.n595 2.6005
R5350 VSS.n594 VSS.n593 2.6005
R5351 VSS.n592 VSS.n591 2.6005
R5352 VSS.n590 VSS.n589 2.6005
R5353 VSS.n588 VSS.n587 2.6005
R5354 VSS.n586 VSS.n585 2.6005
R5355 VSS.n584 VSS.n583 2.6005
R5356 VSS.n582 VSS.n581 2.6005
R5357 VSS.n400 VSS.n399 2.6005
R5358 VSS.n402 VSS.n401 2.6005
R5359 VSS.n404 VSS.n403 2.6005
R5360 VSS.n406 VSS.n405 2.6005
R5361 VSS.n408 VSS.n407 2.6005
R5362 VSS.n782 VSS.n781 2.6005
R5363 VSS.n772 VSS.n771 2.6005
R5364 VSS.n764 VSS.n763 2.6005
R5365 VSS.n762 VSS.n761 2.6005
R5366 VSS.n751 VSS.n750 2.6005
R5367 VSS.n748 VSS.n747 2.6005
R5368 VSS.n746 VSS.n745 2.6005
R5369 VSS.n743 VSS.n742 2.6005
R5370 VSS.n741 VSS.n740 2.6005
R5371 VSS.n738 VSS.n737 2.6005
R5372 VSS.n736 VSS.n735 2.6005
R5373 VSS.n732 VSS.n731 2.6005
R5374 VSS.n717 VSS.n716 2.6005
R5375 VSS.n715 VSS.n714 2.6005
R5376 VSS.n625 VSS.n624 2.6005
R5377 VSS.n528 VSS.n527 2.6005
R5378 VSS.n541 VSS.n540 2.6005
R5379 VSS.n818 VSS.n817 2.6005
R5380 VSS.n815 VSS.n814 2.6005
R5381 VSS.n813 VSS.n812 2.6005
R5382 VSS.n803 VSS.n802 2.6005
R5383 VSS.n805 VSS.n804 2.6005
R5384 VSS.n801 VSS.n800 2.6005
R5385 VSS.n798 VSS.n797 2.6005
R5386 VSS.n795 VSS.n794 2.6005
R5387 VSS.n793 VSS.n792 2.6005
R5388 VSS.n537 VSS.n536 2.6005
R5389 VSS.n546 VSS.n545 2.6005
R5390 VSS.n317 VSS.n316 2.6005
R5391 VSS.n319 VSS.n318 2.6005
R5392 VSS.n325 VSS.n321 2.6005
R5393 VSS.n821 VSS.n820 2.6005
R5394 VSS.n824 VSS.n823 2.6005
R5395 VSS.n826 VSS.n825 2.6005
R5396 VSS.n884 VSS.n883 2.6005
R5397 VSS.n883 VSS.n882 2.6005
R5398 VSS.n873 VSS.n872 2.6005
R5399 VSS.n872 VSS.n871 2.6005
R5400 VSS.n870 VSS.n869 2.6005
R5401 VSS.n869 VSS.n868 2.6005
R5402 VSS.n867 VSS.n866 2.6005
R5403 VSS.n866 VSS.n865 2.6005
R5404 VSS.n863 VSS.n862 2.6005
R5405 VSS.n862 VSS.n861 2.6005
R5406 VSS.n860 VSS.n859 2.6005
R5407 VSS.n859 VSS.n858 2.6005
R5408 VSS.n857 VSS.n856 2.6005
R5409 VSS.n856 VSS.n855 2.6005
R5410 VSS.n854 VSS.n853 2.6005
R5411 VSS.n853 VSS.n852 2.6005
R5412 VSS.n851 VSS.n850 2.6005
R5413 VSS.n850 VSS.n849 2.6005
R5414 VSS.n847 VSS.n846 2.6005
R5415 VSS.n846 VSS.n845 2.6005
R5416 VSS.n844 VSS.n843 2.6005
R5417 VSS.n843 VSS.n842 2.6005
R5418 VSS.n839 VSS.n838 2.6005
R5419 VSS.n838 VSS.n837 2.6005
R5420 VSS.n835 VSS.n834 2.6005
R5421 VSS.n834 VSS.n833 2.6005
R5422 VSS.n832 VSS.n810 2.6005
R5423 VSS.n831 VSS.n830 2.6005
R5424 VSS.n908 VSS.n907 2.6005
R5425 VSS.n911 VSS.n910 2.6005
R5426 VSS.n919 VSS.n918 2.6005
R5427 VSS.n922 VSS.n921 2.6005
R5428 VSS.n930 VSS.n929 2.6005
R5429 VSS.n892 VSS.n891 2.6005
R5430 VSS.n895 VSS.n894 2.6005
R5431 VSS.n935 VSS.n934 2.6005
R5432 VSS.n1155 VSS.n1154 2.6005
R5433 VSS.n1154 VSS.n1153 2.6005
R5434 VSS.n1151 VSS.n1150 2.6005
R5435 VSS.n1150 VSS.n1149 2.6005
R5436 VSS.n1148 VSS.n1147 2.6005
R5437 VSS.n1147 VSS.n1146 2.6005
R5438 VSS.n1144 VSS.n1143 2.6005
R5439 VSS.n1143 VSS.n1142 2.6005
R5440 VSS.n1141 VSS.n1140 2.6005
R5441 VSS.n1140 VSS.n1139 2.6005
R5442 VSS.n1138 VSS.n1137 2.6005
R5443 VSS.n1137 VSS.n1136 2.6005
R5444 VSS.n1134 VSS.n1133 2.6005
R5445 VSS.n1133 VSS.n1132 2.6005
R5446 VSS.n1131 VSS.n1130 2.6005
R5447 VSS.n1130 VSS.n1129 2.6005
R5448 VSS.n1128 VSS.n1127 2.6005
R5449 VSS.n1127 VSS.n1126 2.6005
R5450 VSS.n1124 VSS.n1123 2.6005
R5451 VSS.n1123 VSS.n1122 2.6005
R5452 VSS.n1121 VSS.n1120 2.6005
R5453 VSS.n1120 VSS.n1119 2.6005
R5454 VSS.n1118 VSS.n1117 2.6005
R5455 VSS.n1117 VSS.n1116 2.6005
R5456 VSS.n1115 VSS.n1114 2.6005
R5457 VSS.n1114 VSS.n1113 2.6005
R5458 VSS.n1111 VSS.n1110 2.6005
R5459 VSS.n1110 VSS.n1109 2.6005
R5460 VSS.n1108 VSS.n1107 2.6005
R5461 VSS.n1107 VSS.n1106 2.6005
R5462 VSS.n1105 VSS.n1104 2.6005
R5463 VSS.n1104 VSS.n1103 2.6005
R5464 VSS.n1101 VSS.n1100 2.6005
R5465 VSS.n1100 VSS.n1099 2.6005
R5466 VSS.n1098 VSS.n1097 2.6005
R5467 VSS.n1097 VSS.n1096 2.6005
R5468 VSS.n1095 VSS.n1094 2.6005
R5469 VSS.n1094 VSS.n1093 2.6005
R5470 VSS.n1091 VSS.n1090 2.6005
R5471 VSS.n1090 VSS.n1089 2.6005
R5472 VSS.n1088 VSS.n1087 2.6005
R5473 VSS.n1087 VSS.n1086 2.6005
R5474 VSS.n1084 VSS.n1083 2.6005
R5475 VSS.n1083 VSS.n1082 2.6005
R5476 VSS.n987 VSS.n986 2.6005
R5477 VSS.n411 VSS.n398 2.6005
R5478 VSS.n413 VSS.n412 2.6005
R5479 VSS.n416 VSS.n415 2.6005
R5480 VSS.n418 VSS.n417 2.6005
R5481 VSS.n421 VSS.n420 2.6005
R5482 VSS.n423 VSS.n422 2.6005
R5483 VSS.n425 VSS.n424 2.6005
R5484 VSS.n428 VSS.n427 2.6005
R5485 VSS.n430 VSS.n429 2.6005
R5486 VSS.n432 VSS.n431 2.6005
R5487 VSS.n435 VSS.n434 2.6005
R5488 VSS.n437 VSS.n436 2.6005
R5489 VSS.n439 VSS.n438 2.6005
R5490 VSS.n441 VSS.n440 2.6005
R5491 VSS.n444 VSS.n443 2.6005
R5492 VSS.n446 VSS.n445 2.6005
R5493 VSS.n448 VSS.n447 2.6005
R5494 VSS.n451 VSS.n450 2.6005
R5495 VSS.n453 VSS.n452 2.6005
R5496 VSS.n455 VSS.n454 2.6005
R5497 VSS.n458 VSS.n457 2.6005
R5498 VSS.n460 VSS.n459 2.6005
R5499 VSS.n467 VSS.n466 2.6005
R5500 VSS.n469 VSS.n468 2.6005
R5501 VSS.n234 VSS.n233 2.6005
R5502 VSS.n76 VSS.n75 2.6005
R5503 VSS.n338 VSS.n337 2.6005
R5504 VSS.n336 VSS.n335 2.6005
R5505 VSS.n333 VSS.n332 2.6005
R5506 VSS.n331 VSS.n330 2.6005
R5507 VSS.n329 VSS.n328 2.6005
R5508 VSS.n34 VSS.n33 2.6005
R5509 VSS.n36 VSS.n35 2.6005
R5510 VSS.n38 VSS.n37 2.6005
R5511 VSS.n41 VSS.n40 2.6005
R5512 VSS.n43 VSS.n42 2.6005
R5513 VSS.n45 VSS.n44 2.6005
R5514 VSS.n47 VSS.n46 2.6005
R5515 VSS.n49 VSS.n48 2.6005
R5516 VSS.n51 VSS.n50 2.6005
R5517 VSS.n54 VSS.n53 2.6005
R5518 VSS.n56 VSS.n55 2.6005
R5519 VSS.n58 VSS.n57 2.6005
R5520 VSS.n60 VSS.n59 2.6005
R5521 VSS.n62 VSS.n61 2.6005
R5522 VSS.n65 VSS.n64 2.6005
R5523 VSS.n67 VSS.n66 2.6005
R5524 VSS.n69 VSS.n68 2.6005
R5525 VSS.n72 VSS.n71 2.6005
R5526 VSS.n79 VSS.n78 2.6005
R5527 VSS.n82 VSS.n81 2.6005
R5528 VSS.n98 VSS.n97 2.6005
R5529 VSS.n101 VSS.n100 2.6005
R5530 VSS.n129 VSS.n128 2.6005
R5531 VSS.n132 VSS.n131 2.6005
R5532 VSS.n135 VSS.n134 2.6005
R5533 VSS.n150 VSS.n149 2.6005
R5534 VSS.n154 VSS.n153 2.6005
R5535 VSS.n148 VSS.n147 2.6005
R5536 VSS.n20 VSS.n19 2.6005
R5537 VSS.n89 VSS.n88 2.6005
R5538 VSS.n91 VSS.n90 2.6005
R5539 VSS.n22 VSS.n21 2.6005
R5540 VSS.n25 VSS.n24 2.6005
R5541 VSS.n27 VSS.n26 2.6005
R5542 VSS.n144 VSS.n143 2.6005
R5543 VSS.n158 VSS.n157 2.6005
R5544 VSS.n161 VSS.n160 2.6005
R5545 VSS.n164 VSS.n163 2.6005
R5546 VSS.n238 VSS.n237 2.6005
R5547 VSS.n237 VSS.n236 2.6005
R5548 VSS.n242 VSS.n241 2.6005
R5549 VSS.n241 VSS.n240 2.6005
R5550 VSS.n229 VSS.n228 2.6005
R5551 VSS.n228 VSS.n227 2.6005
R5552 VSS.n226 VSS.n225 2.6005
R5553 VSS.n225 VSS.n224 2.6005
R5554 VSS.n223 VSS.n222 2.6005
R5555 VSS.n222 VSS.n221 2.6005
R5556 VSS.n219 VSS.n218 2.6005
R5557 VSS.n218 VSS.n217 2.6005
R5558 VSS.n216 VSS.n215 2.6005
R5559 VSS.n215 VSS.n214 2.6005
R5560 VSS.n213 VSS.n212 2.6005
R5561 VSS.n212 VSS.n211 2.6005
R5562 VSS.n210 VSS.n209 2.6005
R5563 VSS.n209 VSS.n208 2.6005
R5564 VSS.n207 VSS.n206 2.6005
R5565 VSS.n206 VSS.n205 2.6005
R5566 VSS.n203 VSS.n202 2.6005
R5567 VSS.n202 VSS.n201 2.6005
R5568 VSS.n200 VSS.n199 2.6005
R5569 VSS.n199 VSS.n198 2.6005
R5570 VSS.n197 VSS.n196 2.6005
R5571 VSS.n196 VSS.n195 2.6005
R5572 VSS.n194 VSS.n193 2.6005
R5573 VSS.n193 VSS.n192 2.6005
R5574 VSS.n258 VSS.n257 2.6005
R5575 VSS.n257 VSS.n256 2.6005
R5576 VSS.n261 VSS.n260 2.6005
R5577 VSS.n260 VSS.n259 2.6005
R5578 VSS.n265 VSS.n264 2.6005
R5579 VSS.n264 VSS.n263 2.6005
R5580 VSS.n286 VSS.n285 2.6005
R5581 VSS.n284 VSS.n283 2.6005
R5582 VSS.n281 VSS.n280 2.6005
R5583 VSS.n290 VSS.n289 2.6005
R5584 VSS.n276 VSS.n275 2.6005
R5585 VSS.n278 VSS.n277 2.6005
R5586 VSS.n887 VSS.n886 2.6005
R5587 VSS.n886 VSS.n885 2.6005
R5588 VSS.n2124 VSS.n2123 2.6005
R5589 VSS.n2098 VSS.n2097 2.6005
R5590 VSS.n2090 VSS.n2089 2.6005
R5591 VSS.n2020 VSS.n2019 2.6005
R5592 VSS.n2015 VSS.n2014 2.6005
R5593 VSS.n1169 VSS.n1168 2.6005
R5594 VSS.n1166 VSS.n1165 2.6005
R5595 VSS.n1207 VSS.n1206 2.6005
R5596 VSS.n1216 VSS.n1215 2.6005
R5597 VSS.n1213 VSS.n1212 2.6005
R5598 VSS.n1211 VSS.n1210 2.6005
R5599 VSS.n1246 VSS.n1245 2.6005
R5600 VSS.n1244 VSS.n1243 2.6005
R5601 VSS.n1242 VSS.n1241 2.6005
R5602 VSS.n1249 VSS.n1248 2.6005
R5603 VSS.n2018 VSS.n2017 2.6005
R5604 VSS.n2088 VSS.n2087 2.6005
R5605 VSS.n2096 VSS.n2095 2.6005
R5606 VSS.n2104 VSS.n2103 2.6005
R5607 VSS.n2106 VSS.n2105 2.6005
R5608 VSS.n2112 VSS.n2111 2.6005
R5609 VSS.n2114 VSS.n2113 2.6005
R5610 VSS.n2117 VSS.n2116 2.6005
R5611 VSS.n1294 VSS.n1293 2.6005
R5612 VSS.n1296 VSS.n1295 2.6005
R5613 VSS.n1291 VSS.n1290 2.6005
R5614 VSS.n1305 VSS.n1304 2.6005
R5615 VSS.n1302 VSS.n1301 2.6005
R5616 VSS.n2120 VSS.n2119 2.6005
R5617 VSS.n2127 VSS.n2126 2.6005
R5618 VSS.n2126 VSS.n2125 2.6005
R5619 VSS.n2131 VSS.n2130 2.6005
R5620 VSS.n2130 VSS.n2129 2.6005
R5621 VSS.n2134 VSS.n2133 2.6005
R5622 VSS.n2133 VSS.n2132 2.6005
R5623 VSS.n2137 VSS.n2136 2.6005
R5624 VSS.n2136 VSS.n2135 2.6005
R5625 VSS.n2141 VSS.n2140 2.6005
R5626 VSS.n2140 VSS.n2139 2.6005
R5627 VSS.n2144 VSS.n2143 2.6005
R5628 VSS.n2143 VSS.n2142 2.6005
R5629 VSS.n2147 VSS.n2146 2.6005
R5630 VSS.n2146 VSS.n2145 2.6005
R5631 VSS.n2151 VSS.n2150 2.6005
R5632 VSS.n2150 VSS.n2149 2.6005
R5633 VSS.n2155 VSS.n2154 2.6005
R5634 VSS.n2154 VSS.n2153 2.6005
R5635 VSS.n2158 VSS.n2157 2.6005
R5636 VSS.n2157 VSS.n2156 2.6005
R5637 VSS.n2161 VSS.n2160 2.6005
R5638 VSS.n2160 VSS.n2159 2.6005
R5639 VSS.n2165 VSS.n2164 2.6005
R5640 VSS.n2164 VSS.n2163 2.6005
R5641 VSS.n2185 VSS.n2184 2.6005
R5642 VSS.n1338 VSS.n1337 2.6005
R5643 VSS.n1336 VSS.n1335 2.6005
R5644 VSS.n1334 VSS.n1333 2.6005
R5645 VSS.n1332 VSS.n1331 2.6005
R5646 VSS.n1330 VSS.n1329 2.6005
R5647 VSS.n1328 VSS.n1327 2.6005
R5648 VSS.n1326 VSS.n1325 2.6005
R5649 VSS.n1324 VSS.n1323 2.6005
R5650 VSS.n1322 VSS.n1321 2.6005
R5651 VSS.n1320 VSS.n1319 2.6005
R5652 VSS.n1318 VSS.n1317 2.6005
R5653 VSS.n1316 VSS.n1315 2.6005
R5654 VSS.n1314 VSS.n1313 2.6005
R5655 VSS.n1312 VSS.n1311 2.6005
R5656 VSS.n1668 VSS.n1667 2.6005
R5657 VSS.n1670 VSS.n1669 2.6005
R5658 VSS.n1672 VSS.n1671 2.6005
R5659 VSS.n1674 VSS.n1673 2.6005
R5660 VSS.n1666 VSS.n1665 2.6005
R5661 VSS.n1632 VSS.n1631 2.6005
R5662 VSS.n1612 VSS.n1611 2.6005
R5663 VSS.n1594 VSS.n1593 2.6005
R5664 VSS.n1576 VSS.n1575 2.6005
R5665 VSS.n1557 VSS.n1556 2.6005
R5666 VSS.n1538 VSS.n1537 2.6005
R5667 VSS.n1470 VSS.n1469 2.6005
R5668 VSS.n1468 VSS.n1467 2.6005
R5669 VSS.n1678 VSS.n1677 2.6005
R5670 VSS.n1676 VSS.n1675 2.6005
R5671 VSS.n1680 VSS.n1679 2.6005
R5672 VSS.n1935 VSS.n1934 2.6005
R5673 VSS.n1465 VSS.n1464 2.6005
R5674 VSS.n1639 VSS.n1636 2.6005
R5675 VSS.n1664 VSS.n1662 2.6005
R5676 VSS.n1659 VSS.n1658 2.6005
R5677 VSS.n1661 VSS.n1660 2.6005
R5678 VSS.n1664 VSS.n1663 2.6005
R5679 VSS.n1635 VSS.n1634 2.6005
R5680 VSS.n1639 VSS.n1638 2.6005
R5681 VSS.n1615 VSS.n1614 2.6005
R5682 VSS.n1619 VSS.n1616 2.6005
R5683 VSS.n1597 VSS.n1596 2.6005
R5684 VSS.n1619 VSS.n1618 2.6005
R5685 VSS.n1601 VSS.n1598 2.6005
R5686 VSS.n1579 VSS.n1578 2.6005
R5687 VSS.n1601 VSS.n1600 2.6005
R5688 VSS.n1583 VSS.n1580 2.6005
R5689 VSS.n1560 VSS.n1559 2.6005
R5690 VSS.n1583 VSS.n1582 2.6005
R5691 VSS.n1564 VSS.n1562 2.6005
R5692 VSS.n1541 VSS.n1540 2.6005
R5693 VSS.n1564 VSS.n1563 2.6005
R5694 VSS.n1545 VSS.n1542 2.6005
R5695 VSS.n1473 VSS.n1472 2.6005
R5696 VSS.n1545 VSS.n1544 2.6005
R5697 VSS.n1477 VSS.n1474 2.6005
R5698 VSS.n1477 VSS.n1476 2.6005
R5699 VSS.n1945 VSS.n1944 2.6005
R5700 VSS.n1994 VSS.n1993 2.6005
R5701 VSS.n1948 VSS.n1947 2.6005
R5702 VSS.n1947 VSS.n1946 2.6005
R5703 VSS.n1951 VSS.n1950 2.6005
R5704 VSS.n1950 VSS.n1949 2.6005
R5705 VSS.n1954 VSS.n1953 2.6005
R5706 VSS.n1953 VSS.n1952 2.6005
R5707 VSS.n1957 VSS.n1956 2.6005
R5708 VSS.n1956 VSS.n1955 2.6005
R5709 VSS.n1960 VSS.n1959 2.6005
R5710 VSS.n1959 VSS.n1958 2.6005
R5711 VSS.n1963 VSS.n1962 2.6005
R5712 VSS.n1962 VSS.n1961 2.6005
R5713 VSS.n1966 VSS.n1965 2.6005
R5714 VSS.n1965 VSS.n1964 2.6005
R5715 VSS.n1969 VSS.n1968 2.6005
R5716 VSS.n1968 VSS.n1967 2.6005
R5717 VSS.n1972 VSS.n1971 2.6005
R5718 VSS.n1971 VSS.n1970 2.6005
R5719 VSS.n1933 VSS.n1932 2.6005
R5720 VSS.n1932 VSS.n1931 2.6005
R5721 VSS.n1930 VSS.n1929 2.6005
R5722 VSS.n1929 VSS.n1928 2.6005
R5723 VSS.n1927 VSS.n1926 2.6005
R5724 VSS.n1926 VSS.n1925 2.6005
R5725 VSS.n1924 VSS.n1923 2.6005
R5726 VSS.n1923 VSS.n1922 2.6005
R5727 VSS.n1986 VSS.n1985 2.6005
R5728 VSS.n1985 VSS.n1984 2.6005
R5729 VSS.n1989 VSS.n1988 2.6005
R5730 VSS.n1988 VSS.n1987 2.6005
R5731 VSS.n1992 VSS.n1991 2.6005
R5732 VSS.n1991 VSS.n1990 2.6005
R5733 VSS.n1995 VSS.n1994 2.6005
R5734 VSS.n1996 VSS.n1983 2.6005
R5735 VSS.n1982 VSS.n1981 2.6005
R5736 VSS.n1979 VSS.n1978 2.6005
R5737 VSS.n1976 VSS.n1975 2.6005
R5738 VSS.n2083 VSS.n2082 2.6005
R5739 VSS.n2079 VSS.n2078 2.6005
R5740 VSS.n2076 VSS.n2075 2.6005
R5741 VSS.n2073 VSS.n2072 2.6005
R5742 VSS.n2069 VSS.n2068 2.6005
R5743 VSS.n2065 VSS.n2064 2.6005
R5744 VSS.n2062 VSS.n2061 2.6005
R5745 VSS.n2059 VSS.n2058 2.6005
R5746 VSS.n2055 VSS.n2054 2.6005
R5747 VSS.n2051 VSS.n2050 2.6005
R5748 VSS.n2048 VSS.n2047 2.6005
R5749 VSS.n2045 VSS.n2044 2.6005
R5750 VSS.n2041 VSS.n2040 2.6005
R5751 VSS.n2038 VSS.n2037 2.6005
R5752 VSS.n2029 VSS.n2028 2.6005
R5753 VSS.n2032 VSS.n2031 2.6005
R5754 VSS.n2034 VSS.n2033 2.6005
R5755 VSS.n2026 VSS.n2025 2.6005
R5756 VSS.n1264 VSS.n1263 2.6005
R5757 VSS.n1261 VSS.n1260 2.6005
R5758 VSS.n1257 VSS.n1256 2.6005
R5759 VSS.n1368 VSS.n1367 2.6005
R5760 VSS.n1364 VSS.n1363 2.6005
R5761 VSS.n1362 VSS.n1361 2.6005
R5762 VSS.n1360 VSS.n1359 2.6005
R5763 VSS.n1343 VSS.n1342 2.6005
R5764 VSS.n1346 VSS.n1345 2.6005
R5765 VSS.n1352 VSS.n1351 2.6005
R5766 VSS.n1350 VSS.n1349 2.6005
R5767 VSS.n1354 VSS.n1353 2.6005
R5768 VSS.n1356 VSS.n1355 2.6005
R5769 VSS.n1366 VSS.n1365 2.6005
R5770 VSS.n1252 VSS.n1251 2.6005
R5771 VSS.n1255 VSS.n1254 2.6005
R5772 VSS.n2010 VSS.n2009 2.6005
R5773 VSS.n2001 VSS.n2000 2.6005
R5774 VSS.n1999 VSS.n1998 2.6005
R5775 VSS.n2012 VSS.n2011 2.6005
R5776 VSS.n1372 VSS.n1371 2.6005
R5777 VSS.n1374 VSS.n1373 2.6005
R5778 VSS.n1189 VSS.n1188 2.6005
R5779 VSS.n1394 VSS.n1393 2.6005
R5780 VSS.n1397 VSS.n1396 2.6005
R5781 VSS.n1396 VSS.n1395 2.6005
R5782 VSS.n1393 VSS.n1392 2.6005
R5783 VSS.n1171 VSS.n1170 2.6005
R5784 VSS.n1173 VSS.n1172 2.6005
R5785 VSS.n1196 VSS.n1195 2.6005
R5786 VSS.n1195 VSS.n1194 2.6005
R5787 VSS.n1199 VSS.n1198 2.6005
R5788 VSS.n1198 VSS.n1197 2.6005
R5789 VSS.n1201 VSS.n1200 2.6005
R5790 VSS.n1203 VSS.n1202 2.6005
R5791 VSS.n1192 VSS.n1191 2.6005
R5792 VSS.n1191 VSS.n1190 2.6005
R5793 VSS.n1188 VSS.n1187 2.6005
R5794 VSS.n1230 VSS.t60 2.6005
R5795 VSS.n1232 VSS.n1231 2.6005
R5796 VSS.n1229 VSS.n1228 2.6005
R5797 VSS.n1228 VSS.n1227 2.6005
R5798 VSS.n1225 VSS.n1224 2.6005
R5799 VSS.n1224 VSS.n1223 2.6005
R5800 VSS.n1222 VSS.n1221 2.6005
R5801 VSS.n1221 VSS.n1220 2.6005
R5802 VSS.n1377 VSS.n1376 2.6005
R5803 VSS.n1376 VSS.n1375 2.6005
R5804 VSS.n1403 VSS.n1402 2.6005
R5805 VSS.n1402 VSS.n1401 2.6005
R5806 VSS.n121 VSS.n120 2.6005
R5807 VSS.n120 VSS.t93 2.6005
R5808 VSS.n126 VSS.n125 2.6005
R5809 VSS.n125 VSS.n124 2.6005
R5810 VSS.n1400 VSS.n1399 2.6005
R5811 VSS.n1399 VSS.n1398 2.6005
R5812 VSS.n112 VSS.n111 2.6005
R5813 VSS.n111 VSS.n110 2.6005
R5814 VSS.n119 VSS.n118 2.6005
R5815 VSS.n118 VSS.n117 2.6005
R5816 VSS.n109 VSS.n108 2.6005
R5817 VSS.n17 VSS.n0 2.6005
R5818 VSS.n16 VSS.n15 2.6005
R5819 VSS.n13 VSS.n12 2.6005
R5820 VSS.n11 VSS.n10 2.6005
R5821 VSS.n9 VSS.n8 2.6005
R5822 VSS.n6 VSS.n5 2.6005
R5823 VSS.n4 VSS.n3 2.6005
R5824 VSS.n2 VSS.n1 2.6005
R5825 VSS.n1418 VSS.n1417 2.6005
R5826 VSS.n1416 VSS.n1415 2.6005
R5827 VSS.n1414 VSS.n1413 2.6005
R5828 VSS.n1412 VSS.n1411 2.6005
R5829 VSS.n1410 VSS.n1409 2.6005
R5830 VSS.n1408 VSS.n1407 2.6005
R5831 VSS.n1405 VSS.n1404 2.6005
R5832 VSS.n1178 VSS.n1177 2.6005
R5833 VSS.n1180 VSS.n1179 2.6005
R5834 VSS.n1182 VSS.n1181 2.6005
R5835 VSS.n1273 VSS.n1272 2.6005
R5836 VSS.n1275 VSS.n1274 2.6005
R5837 VSS.n1277 VSS.n1276 2.6005
R5838 VSS.n1279 VSS.n1278 2.6005
R5839 VSS.n1282 VSS.n1281 2.6005
R5840 VSS.n1284 VSS.n1283 2.6005
R5841 VSS.n1287 VSS.n1286 2.6005
R5842 VSS.n1424 VSS.n1423 2.6005
R5843 VSS.n1426 VSS.n1425 2.6005
R5844 VSS.n140 VSS.n138 2.6005
R5845 VSS.n140 VSS.n139 2.6005
R5846 VSS.n1388 VSS.n1387 2.6005
R5847 VSS.n1390 VSS.n1389 2.6005
R5848 VSS.n1435 VSS.n1434 2.6005
R5849 VSS.n1454 VSS.n1453 2.6005
R5850 VSS.n1452 VSS.n1451 2.6005
R5851 VSS.n1449 VSS.n1448 2.6005
R5852 VSS.n1437 VSS.n1436 2.6005
R5853 VSS.n1440 VSS.n1439 2.6005
R5854 VSS.n1443 VSS.n1442 2.6005
R5855 VSS.n2170 VSS.n2169 2.6005
R5856 VSS.n1456 VSS.n1455 2.6005
R5857 VSS.n2167 VSS.n2166 2.6005
R5858 VSS.n2179 VSS.n2178 2.6005
R5859 VSS.n2181 VSS.n2180 2.6005
R5860 VSS.n2176 VSS.n2175 2.6005
R5861 VSS.n1159 VSS.n1157 2.6005
R5862 VSS.n1159 VSS.n1158 2.6005
R5863 VSS.n1260 VSS.n1258 2.41715
R5864 VSS.n2037 VSS.n2035 2.41715
R5865 VSS.n2047 VSS.n2046 2.41715
R5866 VSS.n2050 VSS.n2049 2.41715
R5867 VSS.n2054 VSS.n2052 2.41715
R5868 VSS.n2061 VSS.n2060 2.41715
R5869 VSS.n2064 VSS.n2063 2.41715
R5870 VSS.n2068 VSS.n2066 2.41715
R5871 VSS.n2075 VSS.n2074 2.41715
R5872 VSS.n2078 VSS.n2077 2.41715
R5873 VSS.n2082 VSS.n2080 2.41715
R5874 VSS.n1978 VSS.n1977 2.41715
R5875 VSS.n1826 VSS.n1825 2.41715
R5876 VSS.n1829 VSS.n1828 2.41715
R5877 VSS.n1832 VSS.n1831 2.41715
R5878 VSS.n1835 VSS.n1834 2.41715
R5879 VSS.n1838 VSS.n1837 2.41715
R5880 VSS.n1841 VSS.n1840 2.41715
R5881 VSS.n1844 VSS.n1843 2.41715
R5882 VSS.n1847 VSS.n1846 2.41715
R5883 VSS.n1850 VSS.n1849 2.41715
R5884 VSS.n1853 VSS.n1852 2.41715
R5885 VSS.n1856 VSS.n1855 2.41715
R5886 VSS.n1859 VSS.n1858 2.41715
R5887 VSS.n1862 VSS.n1861 2.41715
R5888 VSS.n1009 VSS.n1008 2.41715
R5889 VSS.n1012 VSS.n1011 2.41715
R5890 VSS.n1015 VSS.n1014 2.41715
R5891 VSS.n1018 VSS.n1017 2.41715
R5892 VSS.n1021 VSS.n1020 2.41715
R5893 VSS.n1024 VSS.n1023 2.41715
R5894 VSS.n1027 VSS.n1026 2.41715
R5895 VSS.n1030 VSS.n1029 2.41715
R5896 VSS.n1033 VSS.n1032 2.41715
R5897 VSS.n905 VSS.n903 2.41715
R5898 VSS.n291 VSS.n290 2.41715
R5899 VSS.n282 VSS.n281 2.41715
R5900 VSS.n905 VSS.n904 2.41715
R5901 VSS.n1260 VSS.n1259 2.41715
R5902 VSS.n1263 VSS.n1262 2.41715
R5903 VSS.n2037 VSS.n2036 2.41715
R5904 VSS.n2040 VSS.n2039 2.41715
R5905 VSS.n2054 VSS.n2053 2.41715
R5906 VSS.n2068 VSS.n2067 2.41715
R5907 VSS.n2082 VSS.n2081 2.41715
R5908 VSS.n1109 VSS.t79 2.35814
R5909 VSS.n175 VSS.n174 1.96785
R5910 VSS.n305 VSS.n304 1.96785
R5911 VSS.n171 VSS.n170 1.96766
R5912 VSS.n303 VSS.n302 1.96766
R5913 VSS.n1187 VSS.t213 1.96543
R5914 VSS.n289 VSS.t169 1.89776
R5915 VSS.n664 VSS.n662 1.65132
R5916 VSS.n653 VSS.n651 1.65132
R5917 VSS.n641 VSS.n639 1.65132
R5918 VSS.n524 VSS.n523 1.65132
R5919 VSS.n485 VSS.n483 1.65132
R5920 VSS.n493 VSS.n491 1.65132
R5921 VSS.n515 VSS.n514 1.65132
R5922 VSS.n690 VSS.n689 1.65132
R5923 VSS.n699 VSS.n698 1.65132
R5924 VSS.n708 VSS.n707 1.65132
R5925 VSS.n545 VSS.n544 1.65132
R5926 VSS.n917 VSS.n912 1.65132
R5927 VSS.n929 VSS.n928 1.65132
R5928 VSS.n233 VSS.n232 1.65132
R5929 VSS.n1233 VSS.n1230 1.65132
R5930 VSS.n1204 VSS.n1201 1.65132
R5931 VSS.n1174 VSS.n1171 1.65132
R5932 VSS.n1427 VSS.n1424 1.65132
R5933 VSS.n690 VSS.n688 1.65076
R5934 VSS.n699 VSS.n697 1.65076
R5935 VSS.n708 VSS.n706 1.65076
R5936 VSS.n641 VSS.n640 1.65076
R5937 VSS.n653 VSS.n652 1.65076
R5938 VSS.n664 VSS.n663 1.65076
R5939 VSS.n321 VSS.n320 1.65076
R5940 VSS.n910 VSS.n909 1.65076
R5941 VSS.n518 VSS.n517 1.65076
R5942 VSS.n508 VSS.n507 1.65076
R5943 VSS.n540 VSS.n539 1.65076
R5944 VSS.n324 VSS.n322 1.65076
R5945 VSS.n24 VSS.n23 1.65076
R5946 VSS.n1174 VSS.n1173 1.65076
R5947 VSS.n1204 VSS.n1203 1.65076
R5948 VSS.n1233 VSS.n1232 1.65076
R5949 VSS.n1427 VSS.n1426 1.65076
R5950 VSS.n1451 VSS.n1450 1.65065
R5951 VSS.n2169 VSS.n2168 1.65065
R5952 VSS.n1237 VSS.n1235 1.65065
R5953 VSS.n2116 VSS.n2115 1.65065
R5954 VSS.n1566 VSS.n1565 1.65065
R5955 VSS.n1547 VSS.n1546 1.65065
R5956 VSS.n1479 VSS.n1478 1.65065
R5957 VSS.n1483 VSS.n1482 1.65065
R5958 VSS.n1551 VSS.n1550 1.65065
R5959 VSS.n1570 VSS.n1569 1.65065
R5960 VSS.n134 VSS.n133 1.65065
R5961 VSS.n153 VSS.n152 1.65065
R5962 VSS.n160 VSS.n159 1.65065
R5963 VSS.n533 VSS.n532 1.65065
R5964 VSS.n792 VSS.n791 1.65065
R5965 VSS.n797 VSS.n796 1.65065
R5966 VSS.n812 VSS.n811 1.65065
R5967 VSS.n817 VSS.n816 1.65065
R5968 VSS.n823 VSS.n822 1.65065
R5969 VSS.n830 VSS.n829 1.65065
R5970 VSS.n780 VSS.n778 1.65065
R5971 VSS.n780 VSS.n779 1.65065
R5972 VSS.n800 VSS.n799 1.65065
R5973 VSS.n147 VSS.n146 1.65065
R5974 VSS.n1237 VSS.n1236 1.65065
R5975 VSS.n1634 VSS.n1633 1.65065
R5976 VSS.n1614 VSS.n1613 1.65065
R5977 VSS.n1618 VSS.n1617 1.65065
R5978 VSS.n1596 VSS.n1595 1.65065
R5979 VSS.n1600 VSS.n1599 1.65065
R5980 VSS.n1578 VSS.n1577 1.65065
R5981 VSS.n1582 VSS.n1581 1.65065
R5982 VSS.n1559 VSS.n1558 1.65065
R5983 VSS.n1540 VSS.n1539 1.65065
R5984 VSS.n1544 VSS.n1543 1.65065
R5985 VSS.n1472 VSS.n1471 1.65065
R5986 VSS.n1476 VSS.n1475 1.65065
R5987 VSS.n1467 VSS.n1466 1.65065
R5988 VSS.n1638 VSS.n1637 1.65065
R5989 VSS.n1562 VSS.n1561 1.65065
R5990 VSS.n2009 VSS.n2008 1.65065
R5991 VSS.n138 VSS.n137 1.65065
R5992 VSS.n1439 VSS.n1438 1.65065
R5993 VSS.n1126 VSS.t35 1.57226
R5994 VSS.n1779 VSS.n1776 1.4405
R5995 VSS.n1503 VSS.n1500 1.4405
R5996 VSS.n1494 VSS.n1491 1.4405
R5997 VSS.n1788 VSS.n1785 1.4405
R5998 VSS.n1776 VSS.n1773 1.4369
R5999 VSS.n1500 VSS.n1497 1.4369
R6000 VSS.n1491 VSS.n1488 1.4369
R6001 VSS.n1785 VSS.n1782 1.4369
R6002 VSS.n279 VSS.n278 1.39588
R6003 VSS.n1254 VSS.n1253 1.39588
R6004 VSS.n921 VSS.n920 1.39588
R6005 VSS.n894 VSS.n893 1.39588
R6006 VSS.n1345 VSS.n1344 1.39574
R6007 VSS.n2028 VSS.n2027 1.39574
R6008 VSS.n2031 VSS.n2030 1.39574
R6009 VSS.n1981 VSS.n1980 1.39574
R6010 VSS.n1304 VSS.n1303 1.39574
R6011 VSS.n1887 VSS.n1886 1.39574
R6012 VSS.n1079 VSS.n1078 1.39574
R6013 VSS.n926 VSS.n925 1.39574
R6014 VSS.n899 VSS.n898 1.39574
R6015 VSS.n934 VSS.n933 1.39574
R6016 VSS.n784 VSS.n783 1.39574
R6017 VSS.n78 VSS.n77 1.39574
R6018 VSS.n287 VSS.n286 1.39574
R6019 VSS.n371 VSS.n370 1.39574
R6020 VSS.n374 VSS.n373 1.39574
R6021 VSS.n1885 VSS.n1865 1.39293
R6022 VSS.n1885 VSS.n1866 1.39293
R6023 VSS.n1885 VSS.n1867 1.39293
R6024 VSS.n1885 VSS.n1868 1.39293
R6025 VSS.n1885 VSS.n1869 1.39293
R6026 VSS.n1885 VSS.n1870 1.39293
R6027 VSS.n1885 VSS.n1871 1.39293
R6028 VSS.n1885 VSS.n1872 1.39293
R6029 VSS.n1885 VSS.n1873 1.39293
R6030 VSS.n1885 VSS.n1874 1.39293
R6031 VSS.n1885 VSS.n1875 1.39293
R6032 VSS.n1885 VSS.n1876 1.39293
R6033 VSS.n1885 VSS.n1877 1.39293
R6034 VSS.n1885 VSS.n1878 1.39293
R6035 VSS.n1885 VSS.n1879 1.39293
R6036 VSS.n1885 VSS.n1880 1.39293
R6037 VSS.n1885 VSS.n1881 1.39293
R6038 VSS.n1885 VSS.n1882 1.39293
R6039 VSS.n1885 VSS.n1883 1.39293
R6040 VSS.n1885 VSS.n1884 1.39293
R6041 VSS.n1077 VSS.n1035 1.39293
R6042 VSS.n1077 VSS.n1036 1.39293
R6043 VSS.n1077 VSS.n1037 1.39293
R6044 VSS.n1077 VSS.n1038 1.39293
R6045 VSS.n1077 VSS.n1039 1.39293
R6046 VSS.n1077 VSS.n1040 1.39293
R6047 VSS.n1077 VSS.n1041 1.39293
R6048 VSS.n1077 VSS.n1042 1.39293
R6049 VSS.n1077 VSS.n1043 1.39293
R6050 VSS.n1077 VSS.n1044 1.39293
R6051 VSS.n1077 VSS.n1045 1.39293
R6052 VSS.n1077 VSS.n1046 1.39293
R6053 VSS.n1077 VSS.n1047 1.39293
R6054 VSS.n1077 VSS.n1048 1.39293
R6055 VSS.n1077 VSS.n1051 1.39293
R6056 VSS.n1077 VSS.n1052 1.39293
R6057 VSS.n1077 VSS.n1053 1.39293
R6058 VSS.n1077 VSS.n1054 1.39293
R6059 VSS.n1077 VSS.n1055 1.39293
R6060 VSS.n1077 VSS.n1056 1.39293
R6061 VSS.n1077 VSS.n1057 1.39293
R6062 VSS.n1077 VSS.n1058 1.39293
R6063 VSS.n1077 VSS.n1059 1.39293
R6064 VSS.n1077 VSS.n1060 1.39293
R6065 VSS.n1077 VSS.n1061 1.39293
R6066 VSS.n1077 VSS.n1062 1.39293
R6067 VSS.n1077 VSS.n1063 1.39293
R6068 VSS.n1077 VSS.n1064 1.39293
R6069 VSS.n1077 VSS.n1065 1.39293
R6070 VSS.n1077 VSS.n1066 1.39293
R6071 VSS.n1077 VSS.n1067 1.39293
R6072 VSS.n1077 VSS.n1068 1.39293
R6073 VSS.n1077 VSS.n1069 1.39293
R6074 VSS.n1077 VSS.n1070 1.39293
R6075 VSS.n1077 VSS.n1071 1.39293
R6076 VSS.n1077 VSS.n1072 1.39293
R6077 VSS.n1077 VSS.n1073 1.39293
R6078 VSS.n1077 VSS.n1074 1.39293
R6079 VSS.n292 VSS.n288 1.39293
R6080 VSS.n292 VSS.n282 1.39293
R6081 VSS.n292 VSS.n291 1.39293
R6082 VSS.n1293 VSS.n1292 1.3824
R6083 VSS.n2123 VSS.n2122 1.34121
R6084 VSS.n2184 VSS.n2183 1.34121
R6085 VSS.n19 VSS.n18 1.3407
R6086 VSS.n527 VSS.n526 1.3407
R6087 VSS.n1998 VSS.n1997 1.3407
R6088 VSS.n1944 VSS.n1943 1.34055
R6089 VSS.n1524 VSS.t164 1.3311
R6090 VSS.n1387 VSS.n1386 1.33029
R6091 VSS.n2017 VSS.n2016 1.32978
R6092 VSS.n1967 VSS.t12 1.32325
R6093 VSS.n2153 VSS.t19 1.31046
R6094 VSS.t151 VSS.t268 1.31046
R6095 VSS.n969 VSS.n966 1.0864
R6096 VSS.n681 VSS.n678 1.0864
R6097 VSS.n951 VSS.n948 1.0864
R6098 VSS.n687 VSS.n684 1.0864
R6099 VSS.n957 VSS.n954 1.0864
R6100 VSS.n696 VSS.n693 1.0864
R6101 VSS.n963 VSS.n960 1.0864
R6102 VSS.n705 VSS.n702 1.0864
R6103 VSS.n1271 VSS.n1270 1.07937
R6104 VSS.n1340 VSS.n1339 1.0792
R6105 VSS.n580 VSS.n579 1.0792
R6106 VSS.n1157 VSS.n1156 1.0792
R6107 VSS.n1885 VSS.n1864 1.01553
R6108 VSS.n1725 VSS.n1694 0.9455
R6109 VSS.n1732 VSS.n1691 0.9455
R6110 VSS.n1739 VSS.n1688 0.9455
R6111 VSS.n1716 VSS.n1715 0.9455
R6112 VSS.n789 VSS.n788 0.915105
R6113 VSS.n668 VSS.n667 0.913698
R6114 VSS.n657 VSS.n656 0.913698
R6115 VSS.n1919 VSS.n1779 0.9131
R6116 VSS.n1507 VSS.n1503 0.9131
R6117 VSS.n1517 VSS.n1494 0.9131
R6118 VSS.n1906 VSS.n1788 0.9131
R6119 VSS.n628 VSS.n559 0.891647
R6120 VSS.n636 VSS.n635 0.891647
R6121 VSS.n646 VSS.n645 0.891647
R6122 VSS.n456 VSS.n381 0.891647
R6123 VSS.n449 VSS.n384 0.891647
R6124 VSS.n758 VSS.n555 0.891647
R6125 VSS.n673 VSS.n558 0.891647
R6126 VSS.n442 VSS.n387 0.891647
R6127 VSS.n433 VSS.n390 0.891647
R6128 VSS.n426 VSS.n393 0.891647
R6129 VSS.n419 VSS.n396 0.891647
R6130 VSS.n414 VSS.n397 0.891647
R6131 VSS.n465 VSS.n464 0.891647
R6132 VSS.n782 VSS.n777 0.864941
R6133 VSS.n744 VSS.n687 0.863534
R6134 VSS.n739 VSS.n696 0.863534
R6135 VSS.n1085 VSS.n985 0.841484
R6136 VSS.n1092 VSS.n981 0.841484
R6137 VSS.n1102 VSS.n969 0.841484
R6138 VSS.n749 VSS.n681 0.841484
R6139 VSS.n1135 VSS.n951 0.841484
R6140 VSS.n1125 VSS.n957 0.841484
R6141 VSS.n1112 VSS.n963 0.841484
R6142 VSS.n734 VSS.n705 0.841484
R6143 VSS.n730 VSS.n729 0.841484
R6144 VSS.n713 VSS.n712 0.841484
R6145 VSS.n770 VSS.n769 0.841484
R6146 VSS.n1145 VSS.n945 0.841484
R6147 VSS.n1152 VSS.n940 0.841484
R6148 VSS.n1421 VSS.t22 0.8195
R6149 VSS.n1421 VSS.n1420 0.8195
R6150 VSS.n1185 VSS.t269 0.8195
R6151 VSS.n1185 VSS.n1184 0.8195
R6152 VSS.n1218 VSS.t155 0.8195
R6153 VSS.n300 VSS.t175 0.8195
R6154 VSS.n300 VSS.n299 0.8195
R6155 VSS.n297 VSS.t208 0.8195
R6156 VSS.n297 VSS.n296 0.8195
R6157 VSS.n294 VSS.t203 0.8195
R6158 VSS.n294 VSS.n293 0.8195
R6159 VSS.n273 VSS.t198 0.8195
R6160 VSS.n273 VSS.n272 0.8195
R6161 VSS.n270 VSS.t191 0.8195
R6162 VSS.n270 VSS.n269 0.8195
R6163 VSS.n267 VSS.t195 0.8195
R6164 VSS.n267 VSS.n266 0.8195
R6165 VSS.n254 VSS.t207 0.8195
R6166 VSS.n254 VSS.n253 0.8195
R6167 VSS.n251 VSS.t206 0.8195
R6168 VSS.n251 VSS.n250 0.8195
R6169 VSS.n248 VSS.t173 0.8195
R6170 VSS.n248 VSS.n247 0.8195
R6171 VSS.n190 VSS.t186 0.8195
R6172 VSS.n190 VSS.n189 0.8195
R6173 VSS.n187 VSS.t189 0.8195
R6174 VSS.n187 VSS.n186 0.8195
R6175 VSS.n184 VSS.t183 0.8195
R6176 VSS.n184 VSS.n183 0.8195
R6177 VSS.n292 VSS.n279 0.804703
R6178 VSS.n1077 VSS.n1049 0.804703
R6179 VSS.n1077 VSS.n1075 0.804703
R6180 VSS.n1886 VSS.n1885 0.804503
R6181 VSS.n789 VSS.n552 0.804503
R6182 VSS.n1078 VSS.n1077 0.804503
R6183 VSS.n789 VSS.n784 0.804503
R6184 VSS.n292 VSS.n287 0.804503
R6185 VSS.n1428 VSS.n1422 0.784447
R6186 VSS.n1193 VSS.n1186 0.762397
R6187 VSS.n1226 VSS.n1219 0.762397
R6188 VSS.n123 VSS.n122 0.762397
R6189 VSS.n1186 VSS.n1183 0.75619
R6190 VSS.n1422 VSS.n1419 0.75619
R6191 VSS.n252 VSS.n249 0.75425
R6192 VSS.n255 VSS.n252 0.75425
R6193 VSS.n188 VSS.n185 0.75425
R6194 VSS.n191 VSS.n188 0.75425
R6195 VSS.n271 VSS.n268 0.75425
R6196 VSS.n274 VSS.n271 0.75425
R6197 VSS.n298 VSS.n295 0.75425
R6198 VSS.n301 VSS.n298 0.75425
R6199 VSS.n2148 VSS.n1972 0.733671
R6200 VSS.n292 VSS.n274 0.731479
R6201 VSS.n262 VSS.n255 0.723312
R6202 VSS.n204 VSS.n191 0.723312
R6203 VSS.n220 VSS.n182 0.723312
R6204 VSS.n230 VSS.n177 0.723312
R6205 VSS.n848 VSS.n309 0.723312
R6206 VSS.n836 VSS.n313 0.723312
R6207 VSS.n864 VSS.n301 0.723312
R6208 VSS.n358 VSS.n327 0.665656
R6209 VSS.n365 VSS.n326 0.665656
R6210 VSS.n1077 VSS.n1050 0.631461
R6211 VSS.n1077 VSS.n1076 0.631461
R6212 VSS.n105 VSS.n104 0.631461
R6213 VSS.n2122 VSS.n2121 0.631461
R6214 VSS.n1943 VSS.n1942 0.631226
R6215 VSS.n1309 VSS.n1308 0.631226
R6216 VSS.n1209 VSS.t20 0.5465
R6217 VSS.n1209 VSS.n1208 0.5465
R6218 VSS.n1239 VSS.t61 0.5465
R6219 VSS.n1239 VSS.n1238 0.5465
R6220 VSS.n1463 VSS.t152 0.5465
R6221 VSS.n1463 VSS.n1462 0.5465
R6222 VSS.n1974 VSS.t148 0.5465
R6223 VSS.n1974 VSS.n1973 0.5465
R6224 VSS.n1787 VSS.t10 0.5465
R6225 VSS.n1787 VSS.n1786 0.5465
R6226 VSS.n1784 VSS.t294 0.5465
R6227 VSS.n1784 VSS.n1783 0.5465
R6228 VSS.n1781 VSS.t64 0.5465
R6229 VSS.n1781 VSS.n1780 0.5465
R6230 VSS.n1714 VSS.t166 0.5465
R6231 VSS.n1714 VSS.n1713 0.5465
R6232 VSS.n1778 VSS.t161 0.5465
R6233 VSS.n1778 VSS.n1777 0.5465
R6234 VSS.n1775 VSS.t56 0.5465
R6235 VSS.n1775 VSS.n1774 0.5465
R6236 VSS.n1772 VSS.t134 0.5465
R6237 VSS.n1772 VSS.n1771 0.5465
R6238 VSS.n1693 VSS.t277 0.5465
R6239 VSS.n1693 VSS.n1692 0.5465
R6240 VSS.n1502 VSS.t143 0.5465
R6241 VSS.n1502 VSS.n1501 0.5465
R6242 VSS.n1499 VSS.t167 0.5465
R6243 VSS.n1499 VSS.n1498 0.5465
R6244 VSS.n1496 VSS.t144 0.5465
R6245 VSS.n1496 VSS.n1495 0.5465
R6246 VSS.n1690 VSS.t297 0.5465
R6247 VSS.n1690 VSS.n1689 0.5465
R6248 VSS.n1493 VSS.t139 0.5465
R6249 VSS.n1493 VSS.n1492 0.5465
R6250 VSS.n1490 VSS.t5 0.5465
R6251 VSS.n1490 VSS.n1489 0.5465
R6252 VSS.n1487 VSS.t65 0.5465
R6253 VSS.n1487 VSS.n1486 0.5465
R6254 VSS.n1687 VSS.t168 0.5465
R6255 VSS.n1687 VSS.n1686 0.5465
R6256 VSS.n980 VSS.t111 0.5465
R6257 VSS.n980 VSS.n979 0.5465
R6258 VSS.n974 VSS.t100 0.5465
R6259 VSS.n974 VSS.n973 0.5465
R6260 VSS.n634 VSS.t117 0.5465
R6261 VSS.n634 VSS.n633 0.5465
R6262 VSS.n644 VSS.t241 0.5465
R6263 VSS.n644 VSS.n643 0.5465
R6264 VSS.n965 VSS.t282 0.5465
R6265 VSS.n965 VSS.n964 0.5465
R6266 VSS.n968 VSS.t27 0.5465
R6267 VSS.n968 VSS.n967 0.5465
R6268 VSS.n944 VSS.t77 0.5465
R6269 VSS.n941 VSS.t75 0.5465
R6270 VSS.n768 VSS.t283 0.5465
R6271 VSS.n765 VSS.t242 0.5465
R6272 VSS.n379 VSS.t263 0.5465
R6273 VSS.n724 VSS.t91 0.5465
R6274 VSS.n724 VSS.n723 0.5465
R6275 VSS.n728 VSS.t128 0.5465
R6276 VSS.n728 VSS.n727 0.5465
R6277 VSS.n383 VSS.t281 0.5465
R6278 VSS.n383 VSS.n382 0.5465
R6279 VSS.n677 VSS.t32 0.5465
R6280 VSS.n677 VSS.n676 0.5465
R6281 VSS.n680 VSS.t72 0.5465
R6282 VSS.n680 VSS.n679 0.5465
R6283 VSS.n553 VSS.t34 0.5465
R6284 VSS.n557 VSS.t221 0.5465
R6285 VSS.n557 VSS.n556 0.5465
R6286 VSS.n947 VSS.t40 0.5465
R6287 VSS.n947 VSS.n946 0.5465
R6288 VSS.n950 VSS.t230 0.5465
R6289 VSS.n950 VSS.n949 0.5465
R6290 VSS.n386 VSS.t48 0.5465
R6291 VSS.n386 VSS.n385 0.5465
R6292 VSS.n683 VSS.t273 0.5465
R6293 VSS.n683 VSS.n682 0.5465
R6294 VSS.n686 VSS.t245 0.5465
R6295 VSS.n686 VSS.n685 0.5465
R6296 VSS.n666 VSS.t78 0.5465
R6297 VSS.n666 VSS.n665 0.5465
R6298 VSS.n953 VSS.t251 0.5465
R6299 VSS.n953 VSS.n952 0.5465
R6300 VSS.n956 VSS.t257 0.5465
R6301 VSS.n956 VSS.n955 0.5465
R6302 VSS.n389 VSS.t276 0.5465
R6303 VSS.n389 VSS.n388 0.5465
R6304 VSS.n692 VSS.t248 0.5465
R6305 VSS.n692 VSS.n691 0.5465
R6306 VSS.n695 VSS.t80 0.5465
R6307 VSS.n695 VSS.n694 0.5465
R6308 VSS.n655 VSS.t254 0.5465
R6309 VSS.n655 VSS.n654 0.5465
R6310 VSS.n959 VSS.t233 0.5465
R6311 VSS.n959 VSS.n958 0.5465
R6312 VSS.n962 VSS.t272 0.5465
R6313 VSS.n962 VSS.n961 0.5465
R6314 VSS.n392 VSS.t236 0.5465
R6315 VSS.n392 VSS.n391 0.5465
R6316 VSS.n701 VSS.t76 0.5465
R6317 VSS.n701 VSS.n700 0.5465
R6318 VSS.n704 VSS.t262 0.5465
R6319 VSS.n704 VSS.n703 0.5465
R6320 VSS.n395 VSS.t109 0.5465
R6321 VSS.n395 VSS.n394 0.5465
R6322 VSS.n1921 VSS.n1920 0.524768
R6323 VSS.n978 VSS.n975 0.491811
R6324 VSS.n984 VSS.n983 0.491811
R6325 VSS.n711 VSS.n710 0.491811
R6326 VSS.n726 VSS.n725 0.491811
R6327 VSS.n776 VSS.n773 0.491811
R6328 VSS.n767 VSS.n766 0.491811
R6329 VSS.n939 VSS.n936 0.491811
R6330 VSS.n943 VSS.n942 0.491811
R6331 VSS.n381 VSS.n380 0.490336
R6332 VSS.n555 VSS.n554 0.490336
R6333 VSS.n464 VSS.n463 0.490336
R6334 VSS.n788 VSS.n787 0.490336
R6335 VSS.n975 VSS.n972 0.484434
R6336 VSS.n983 VSS.n982 0.484434
R6337 VSS.n985 VSS.n984 0.484434
R6338 VSS.n981 VSS.n978 0.484434
R6339 VSS.n729 VSS.n726 0.484434
R6340 VSS.n710 VSS.n709 0.484434
R6341 VSS.n712 VSS.n711 0.484434
R6342 VSS.n725 VSS.n722 0.484434
R6343 VSS.n769 VSS.n767 0.484434
R6344 VSS.n777 VSS.n776 0.484434
R6345 VSS.n945 VSS.n943 0.484434
R6346 VSS.n940 VSS.n939 0.484434
R6347 VSS.n1630 VSS.n1622 0.476417
R6348 VSS.n1610 VSS.n1604 0.476417
R6349 VSS.n1592 VSS.n1587 0.476417
R6350 VSS.n1648 VSS.n1647 0.476417
R6351 VSS.n1657 VSS.n1651 0.476417
R6352 VSS.n1755 VSS.n1754 0.476417
R6353 VSS.n642 VSS.n641 0.476417
R6354 VSS.n657 VSS.n653 0.476417
R6355 VSS.n668 VSS.n664 0.476417
R6356 VSS.n476 VSS.n474 0.476417
R6357 VSS.n915 VSS.n914 0.476417
R6358 VSS.n487 VSS.n485 0.476417
R6359 VSS.n915 VSS.n913 0.476417
R6360 VSS.n495 VSS.n493 0.476417
R6361 VSS.n504 VSS.n502 0.476417
R6362 VSS.n744 VSS.n690 0.476417
R6363 VSS.n739 VSS.n699 0.476417
R6364 VSS.n733 VSS.n708 0.476417
R6365 VSS.n325 VSS.n324 0.476417
R6366 VSS.n790 VSS.n549 0.476417
R6367 VSS.n919 VSS.n917 0.476417
R6368 VSS.n916 VSS.n915 0.476417
R6369 VSS.n232 VSS.n231 0.476417
R6370 VSS.n87 VSS.n86 0.476417
R6371 VSS.n32 VSS.n31 0.476417
R6372 VSS.n96 VSS.n95 0.476417
R6373 VSS.n107 VSS.n106 0.476417
R6374 VSS.n2024 VSS.n2023 0.476417
R6375 VSS.n2094 VSS.n2093 0.476417
R6376 VSS.n2102 VSS.n2101 0.476417
R6377 VSS.n2110 VSS.n2109 0.476417
R6378 VSS.n1300 VSS.n1299 0.476417
R6379 VSS.n1684 VSS.n1683 0.476417
R6380 VSS.n1372 VSS.n1310 0.476417
R6381 VSS.n1175 VSS.n1174 0.476417
R6382 VSS.n1205 VSS.n1204 0.476417
R6383 VSS.n1234 VSS.n1233 0.476417
R6384 VSS.n1428 VSS.n1427 0.476417
R6385 VSS.n1443 VSS.n1433 0.476417
R6386 VSS.n1458 VSS.n1447 0.476417
R6387 VSS.n2176 VSS.n2174 0.476417
R6388 VSS.n1586 VSS.n1585 0.476176
R6389 VSS.n782 VSS.n780 0.476176
R6390 VSS.n829 VSS.n828 0.476176
R6391 VSS.n1247 VSS.n1237 0.476176
R6392 VSS.n1942 VSS.n1941 0.476176
R6393 VSS.n1942 VSS.n1939 0.476176
R6394 VSS.n1942 VSS.n1940 0.476176
R6395 VSS.n2007 VSS.n2003 0.476176
R6396 VSS.n2007 VSS.n2004 0.476176
R6397 VSS.n2007 VSS.n2006 0.476176
R6398 VSS.n2007 VSS.n2005 0.476176
R6399 VSS.n2007 VSS.n2002 0.476176
R6400 VSS.n2008 VSS.n2007 0.476176
R6401 VSS.n2173 VSS.n2172 0.476176
R6402 VSS.n1972 VSS.n1921 0.455622
R6403 VSS.n1268 VSS.n1267 0.431879
R6404 VSS.n114 VSS.n113 0.416362
R6405 VSS.n828 VSS.n827 0.393439
R6406 VSS.n1161 VSS.n1160 0.347167
R6407 VSS.n176 VSS.n173 0.328156
R6408 VSS.n181 VSS.n180 0.328156
R6409 VSS.n309 VSS.n308 0.328156
R6410 VSS.n313 VSS.n312 0.328156
R6411 VSS.n173 VSS.n172 0.325344
R6412 VSS.n180 VSS.n179 0.325344
R6413 VSS.n311 VSS.n310 0.325344
R6414 VSS.n307 VSS.n306 0.325344
R6415 VSS.n179 VSS.n178 0.323938
R6416 VSS.n172 VSS.n169 0.323938
R6417 VSS.n182 VSS.n181 0.321125
R6418 VSS.n177 VSS.n176 0.321125
R6419 VSS.n312 VSS.n311 0.321125
R6420 VSS.n308 VSS.n307 0.321125
R6421 VSS.n1385 VSS.n1169 0.307168
R6422 VSS.n156 VSS.n155 0.298318
R6423 VSS.n1162 VSS.n1161 0.297833
R6424 VSS.n142 VSS.n141 0.2912
R6425 VSS.n488 VSS.n476 0.224477
R6426 VSS.n115 VSS.n114 0.219293
R6427 VSS.n1269 VSS.n1268 0.203776
R6428 VSS.n166 VSS.n165 0.190706
R6429 VSS.n167 VSS.n166 0.18545
R6430 VSS.n1459 VSS.n1444 0.18545
R6431 VSS.n176 VSS.n175 0.181095
R6432 VSS.n1381 VSS.n1380 0.1805
R6433 VSS.n1380 VSS.n1379 0.1805
R6434 VSS.n172 VSS.n171 0.18047
R6435 VSS.n306 VSS.n305 0.179637
R6436 VSS.n308 VSS.n303 0.17927
R6437 VSS.n1921 VSS.n1764 0.173915
R6438 VSS.n932 VSS.n931 0.162432
R6439 VSS.n1358 VSS.n1348 0.157022
R6440 VSS.n1370 VSS.n1358 0.157022
R6441 VSS.n2057 VSS.n2043 0.157022
R6442 VSS.n2071 VSS.n2057 0.157022
R6443 VSS.n2085 VSS.n2071 0.157022
R6444 VSS.n2086 VSS.n2085 0.157022
R6445 VSS.n1459 VSS.n1458 0.148531
R6446 VSS.n1757 VSS.n1756 0.146841
R6447 VSS.n1758 VSS.n1757 0.146841
R6448 VSS.n1759 VSS.n1758 0.146841
R6449 VSS.n1760 VSS.n1759 0.146841
R6450 VSS.n1761 VSS.n1760 0.146841
R6451 VSS.n1762 VSS.n1761 0.146841
R6452 VSS.n1763 VSS.n1762 0.146841
R6453 VSS.n1764 VSS.n1763 0.146841
R6454 VSS.n1379 VSS.n1266 0.14495
R6455 VSS.n107 VSS.n102 0.1445
R6456 VSS.n87 VSS.n83 0.1445
R6457 VSS.n1382 VSS.n1381 0.1409
R6458 VSS.n161 VSS.n158 0.1405
R6459 VSS.n238 VSS.n234 0.1405
R6460 VSS.n135 VSS.n132 0.1405
R6461 VSS.n168 VSS.n167 0.14045
R6462 VSS.n1460 VSS.n1459 0.14045
R6463 VSS.n79 VSS.n76 0.139071
R6464 VSS.n1163 VSS.n1162 0.135
R6465 VSS.n1160 VSS.n932 0.133795
R6466 VSS.n1444 VSS.n1443 0.132253
R6467 VSS.n488 VSS.n487 0.129705
R6468 VSS.n496 VSS.n495 0.129705
R6469 VSS.n573 VSS.n572 0.1265
R6470 VSS.n572 VSS.n570 0.1265
R6471 VSS.n570 VSS.n568 0.1265
R6472 VSS.n568 VSS.n566 0.1265
R6473 VSS.n566 VSS.n564 0.1265
R6474 VSS.n564 VSS.n562 0.1265
R6475 VSS.n991 VSS.n989 0.1265
R6476 VSS.n993 VSS.n991 0.1265
R6477 VSS.n995 VSS.n993 0.1265
R6478 VSS.n997 VSS.n995 0.1265
R6479 VSS.n999 VSS.n997 0.1265
R6480 VSS.n1001 VSS.n999 0.1265
R6481 VSS.n1003 VSS.n1001 0.1265
R6482 VSS.n1005 VSS.n1003 0.1265
R6483 VSS.n1007 VSS.n1005 0.1265
R6484 VSS.n1010 VSS.n1007 0.1265
R6485 VSS.n1013 VSS.n1010 0.1265
R6486 VSS.n1016 VSS.n1013 0.1265
R6487 VSS.n1019 VSS.n1016 0.1265
R6488 VSS.n1022 VSS.n1019 0.1265
R6489 VSS.n1025 VSS.n1022 0.1265
R6490 VSS.n1028 VSS.n1025 0.1265
R6491 VSS.n1031 VSS.n1028 0.1265
R6492 VSS.n1034 VSS.n1031 0.1265
R6493 VSS.n1080 VSS.n1034 0.1265
R6494 VSS.n101 VSS.n99 0.124786
R6495 VSS.n808 VSS.n325 0.122321
R6496 VSS.n807 VSS.n790 0.122321
R6497 VSS.n832 VSS.n809 0.121759
R6498 VSS.n246 VSS.n245 0.120384
R6499 VSS.n1163 VSS.n168 0.1184
R6500 VSS.n2187 VSS.n1460 0.1184
R6501 VSS.n164 VSS.n162 0.117643
R6502 VSS.n130 VSS.n129 0.116214
R6503 VSS.n166 VSS.n156 0.11435
R6504 VSS.n1444 VSS.n1430 0.11435
R6505 VSS.n1381 VSS.n1205 0.1139
R6506 VSS.n1380 VSS.n1234 0.1139
R6507 VSS.n1429 VSS.n1428 0.1139
R6508 VSS.n520 VSS.n497 0.112659
R6509 VSS.n789 VSS.n782 0.112306
R6510 VSS.n807 VSS.n543 0.111977
R6511 VSS.n1430 VSS.n1391 0.109591
R6512 VSS.n156 VSS.n142 0.10895
R6513 VSS.n1430 VSS.n1429 0.10895
R6514 VSS.n1756 VSS.n1684 0.10805
R6515 VSS.n1764 VSS.n1477 0.10805
R6516 VSS.n1763 VSS.n1545 0.10805
R6517 VSS.n1762 VSS.n1564 0.10805
R6518 VSS.n1761 VSS.n1583 0.10805
R6519 VSS.n1760 VSS.n1601 0.10805
R6520 VSS.n1759 VSS.n1619 0.10805
R6521 VSS.n1758 VSS.n1639 0.10805
R6522 VSS.n1757 VSS.n1664 0.10805
R6523 VSS.n543 VSS.n542 0.107536
R6524 VSS.n807 VSS.n806 0.107536
R6525 VSS.n543 VSS.n529 0.106571
R6526 VSS.n543 VSS.n520 0.105841
R6527 VSS.n808 VSS.n807 0.103795
R6528 VSS.n82 VSS.n80 0.101929
R6529 VSS.n2043 VSS.n2024 0.09995
R6530 VSS.n1996 VSS.n1995 0.0963696
R6531 VSS.n1995 VSS.n1992 0.0963696
R6532 VSS.n1992 VSS.n1989 0.0963696
R6533 VSS.n1989 VSS.n1986 0.0963696
R6534 VSS.n1927 VSS.n1924 0.0963696
R6535 VSS.n1930 VSS.n1927 0.0963696
R6536 VSS.n1933 VSS.n1930 0.0963696
R6537 VSS.n1972 VSS.n1933 0.0963696
R6538 VSS.n1972 VSS.n1969 0.0963696
R6539 VSS.n1969 VSS.n1966 0.0963696
R6540 VSS.n1966 VSS.n1963 0.0963696
R6541 VSS.n1963 VSS.n1960 0.0963696
R6542 VSS.n1960 VSS.n1957 0.0963696
R6543 VSS.n1957 VSS.n1954 0.0963696
R6544 VSS.n1954 VSS.n1951 0.0963696
R6545 VSS.n1951 VSS.n1948 0.0963696
R6546 VSS.n1948 VSS.n1945 0.0963696
R6547 VSS.n809 VSS.n808 0.0956136
R6548 VSS.n972 VSS.n971 0.0953
R6549 VSS.n978 VSS.n977 0.0953
R6550 VSS.n726 VSS.n719 0.0953
R6551 VSS.n722 VSS.n721 0.0953
R6552 VSS.n463 VSS.n462 0.0953
R6553 VSS.n776 VSS.n775 0.0953
R6554 VSS.n787 VSS.n786 0.0953
R6555 VSS.n939 VSS.n938 0.0953
R6556 VSS.n154 VSS.n151 0.0947857
R6557 VSS.n1380 VSS.n1247 0.09365
R6558 VSS.n75 VSS.n74 0.0926053
R6559 VSS.n237 VSS.n235 0.0926053
R6560 VSS.n1379 VSS.n1378 0.0923
R6561 VSS.n142 VSS.n127 0.0923
R6562 VSS.n1758 VSS.n1648 0.09185
R6563 VSS.n1759 VSS.n1630 0.09185
R6564 VSS.n1760 VSS.n1610 0.09185
R6565 VSS.n1761 VSS.n1592 0.09185
R6566 VSS.n1762 VSS.n1574 0.09185
R6567 VSS.n1763 VSS.n1555 0.09185
R6568 VSS.n1764 VSS.n1536 0.09185
R6569 VSS.n1757 VSS.n1657 0.09185
R6570 VSS.n1756 VSS.n1755 0.09185
R6571 VSS.n1162 VSS.n246 0.0915425
R6572 VSS.n1225 VSS.n1222 0.0914278
R6573 VSS.n121 VSS.n119 0.0914278
R6574 VSS.n1397 VSS.n1394 0.0914278
R6575 VSS.n1192 VSS.n1189 0.0914278
R6576 VSS.n1199 VSS.n1196 0.0914278
R6577 VSS.n1468 VSS.n1465 0.0914278
R6578 VSS.n1473 VSS.n1470 0.0914278
R6579 VSS.n1541 VSS.n1538 0.0914278
R6580 VSS.n1560 VSS.n1557 0.0914278
R6581 VSS.n1579 VSS.n1576 0.0914278
R6582 VSS.n1597 VSS.n1594 0.0914278
R6583 VSS.n1615 VSS.n1612 0.0914278
R6584 VSS.n1635 VSS.n1632 0.0914278
R6585 VSS.n1661 VSS.n1659 0.0914278
R6586 VSS.n1678 VSS.n1676 0.0914278
R6587 VSS.n1680 VSS.n1678 0.0914278
R6588 VSS.n1305 VSS.n1302 0.0914278
R6589 VSS.n1296 VSS.n1294 0.0914278
R6590 VSS.n1213 VSS.n1211 0.0914278
R6591 VSS.n1246 VSS.n1244 0.0914278
R6592 VSS.n1244 VSS.n1242 0.0914278
R6593 VSS.n2020 VSS.n2018 0.0914278
R6594 VSS.n2090 VSS.n2088 0.0914278
R6595 VSS.n2098 VSS.n2096 0.0914278
R6596 VSS.n1626 VSS.n1624 0.0914278
R6597 VSS.n1571 VSS.n1568 0.0914278
R6598 VSS.n1552 VSS.n1549 0.0914278
R6599 VSS.n1484 VSS.n1481 0.0914278
R6600 VSS.n1655 VSS.n1653 0.0914278
R6601 VSS.n1643 VSS.n1641 0.0914278
R6602 VSS.n2106 VSS.n2104 0.0914278
R6603 VSS.n2114 VSS.n2112 0.0914278
R6604 VSS.n2117 VSS.n2114 0.0914278
R6605 VSS.n2124 VSS.n2120 0.0914278
R6606 VSS.n91 VSS.n89 0.0914278
R6607 VSS.n25 VSS.n22 0.0914278
R6608 VSS.n27 VSS.n25 0.0914278
R6609 VSS.n364 VSS.n362 0.0914278
R6610 VSS.n362 VSS.n360 0.0914278
R6611 VSS.n357 VSS.n355 0.0914278
R6612 VSS.n355 VSS.n353 0.0914278
R6613 VSS.n353 VSS.n351 0.0914278
R6614 VSS.n351 VSS.n349 0.0914278
R6615 VSS.n346 VSS.n344 0.0914278
R6616 VSS.n344 VSS.n342 0.0914278
R6617 VSS.n342 VSS.n340 0.0914278
R6618 VSS.n340 VSS.n338 0.0914278
R6619 VSS.n338 VSS.n336 0.0914278
R6620 VSS.n333 VSS.n331 0.0914278
R6621 VSS.n331 VSS.n329 0.0914278
R6622 VSS.n36 VSS.n34 0.0914278
R6623 VSS.n38 VSS.n36 0.0914278
R6624 VSS.n43 VSS.n41 0.0914278
R6625 VSS.n45 VSS.n43 0.0914278
R6626 VSS.n47 VSS.n45 0.0914278
R6627 VSS.n49 VSS.n47 0.0914278
R6628 VSS.n51 VSS.n49 0.0914278
R6629 VSS.n56 VSS.n54 0.0914278
R6630 VSS.n58 VSS.n56 0.0914278
R6631 VSS.n60 VSS.n58 0.0914278
R6632 VSS.n62 VSS.n60 0.0914278
R6633 VSS.n67 VSS.n65 0.0914278
R6634 VSS.n69 VSS.n67 0.0914278
R6635 VSS.n372 VSS.n369 0.0914278
R6636 VSS.n377 VSS.n375 0.0914278
R6637 VSS.n534 VSS.n531 0.0914278
R6638 VSS.n541 VSS.n538 0.0914278
R6639 VSS.n538 VSS.n537 0.0914278
R6640 VSS.n795 VSS.n793 0.0914278
R6641 VSS.n798 VSS.n795 0.0914278
R6642 VSS.n801 VSS.n798 0.0914278
R6643 VSS.n805 VSS.n803 0.0914278
R6644 VSS.n815 VSS.n813 0.0914278
R6645 VSS.n818 VSS.n815 0.0914278
R6646 VSS.n824 VSS.n821 0.0914278
R6647 VSS.n826 VSS.n824 0.0914278
R6648 VSS.n831 VSS.n826 0.0914278
R6649 VSS.n1338 VSS.n1336 0.0914278
R6650 VSS.n1336 VSS.n1334 0.0914278
R6651 VSS.n1334 VSS.n1332 0.0914278
R6652 VSS.n1332 VSS.n1330 0.0914278
R6653 VSS.n1330 VSS.n1328 0.0914278
R6654 VSS.n1328 VSS.n1326 0.0914278
R6655 VSS.n1326 VSS.n1324 0.0914278
R6656 VSS.n1324 VSS.n1322 0.0914278
R6657 VSS.n1322 VSS.n1320 0.0914278
R6658 VSS.n1320 VSS.n1318 0.0914278
R6659 VSS.n1318 VSS.n1316 0.0914278
R6660 VSS.n1316 VSS.n1314 0.0914278
R6661 VSS.n1314 VSS.n1312 0.0914278
R6662 VSS.n1670 VSS.n1668 0.0914278
R6663 VSS.n1672 VSS.n1670 0.0914278
R6664 VSS.n1674 VSS.n1672 0.0914278
R6665 VSS.n1352 VSS.n1350 0.0914278
R6666 VSS.n1354 VSS.n1352 0.0914278
R6667 VSS.n1362 VSS.n1360 0.0914278
R6668 VSS.n1364 VSS.n1362 0.0914278
R6669 VSS.n1368 VSS.n1366 0.0914278
R6670 VSS.n1255 VSS.n1252 0.0914278
R6671 VSS.n1257 VSS.n1255 0.0914278
R6672 VSS.n1261 VSS.n1257 0.0914278
R6673 VSS.n2029 VSS.n2026 0.0914278
R6674 VSS.n2032 VSS.n2029 0.0914278
R6675 VSS.n2034 VSS.n2032 0.0914278
R6676 VSS.n2038 VSS.n2034 0.0914278
R6677 VSS.n2048 VSS.n2045 0.0914278
R6678 VSS.n2051 VSS.n2048 0.0914278
R6679 VSS.n2062 VSS.n2059 0.0914278
R6680 VSS.n2065 VSS.n2062 0.0914278
R6681 VSS.n2076 VSS.n2073 0.0914278
R6682 VSS.n2079 VSS.n2076 0.0914278
R6683 VSS.n1979 VSS.n1976 0.0914278
R6684 VSS.n1982 VSS.n1979 0.0914278
R6685 VSS.n2012 VSS.n2010 0.0914278
R6686 VSS.n2010 VSS.n2001 0.0914278
R6687 VSS.n2001 VSS.n1999 0.0914278
R6688 VSS.n1377 VSS.n1374 0.0914278
R6689 VSS.n1403 VSS.n1400 0.0914278
R6690 VSS.n112 VSS.n109 0.0914278
R6691 VSS.n17 VSS.n16 0.0914278
R6692 VSS.n13 VSS.n11 0.0914278
R6693 VSS.n11 VSS.n9 0.0914278
R6694 VSS.n6 VSS.n4 0.0914278
R6695 VSS.n4 VSS.n2 0.0914278
R6696 VSS.n1418 VSS.n1416 0.0914278
R6697 VSS.n1416 VSS.n1414 0.0914278
R6698 VSS.n1414 VSS.n1412 0.0914278
R6699 VSS.n1412 VSS.n1410 0.0914278
R6700 VSS.n1410 VSS.n1408 0.0914278
R6701 VSS.n1180 VSS.n1178 0.0914278
R6702 VSS.n1275 VSS.n1273 0.0914278
R6703 VSS.n1277 VSS.n1275 0.0914278
R6704 VSS.n1279 VSS.n1277 0.0914278
R6705 VSS.n1284 VSS.n1282 0.0914278
R6706 VSS.n1440 VSS.n1437 0.0914278
R6707 VSS.n1452 VSS.n1449 0.0914278
R6708 VSS.n1454 VSS.n1452 0.0914278
R6709 VSS.n2170 VSS.n2167 0.0914278
R6710 VSS.n2181 VSS.n2179 0.0914278
R6711 VSS.n1372 VSS.n1305 0.0905
R6712 VSS.n1700 VSS.n1698 0.0905
R6713 VSS.n1698 VSS.n1696 0.0905
R6714 VSS.n1792 VSS.n1790 0.0905
R6715 VSS.n1794 VSS.n1792 0.0905
R6716 VSS.n1796 VSS.n1794 0.0905
R6717 VSS.n1798 VSS.n1796 0.0905
R6718 VSS.n1800 VSS.n1798 0.0905
R6719 VSS.n1802 VSS.n1800 0.0905
R6720 VSS.n1804 VSS.n1802 0.0905
R6721 VSS.n1806 VSS.n1804 0.0905
R6722 VSS.n1808 VSS.n1806 0.0905
R6723 VSS.n1810 VSS.n1808 0.0905
R6724 VSS.n1812 VSS.n1810 0.0905
R6725 VSS.n1814 VSS.n1812 0.0905
R6726 VSS.n1816 VSS.n1814 0.0905
R6727 VSS.n1818 VSS.n1816 0.0905
R6728 VSS.n1820 VSS.n1818 0.0905
R6729 VSS.n1822 VSS.n1820 0.0905
R6730 VSS.n1824 VSS.n1822 0.0905
R6731 VSS.n1827 VSS.n1824 0.0905
R6732 VSS.n1830 VSS.n1827 0.0905
R6733 VSS.n1833 VSS.n1830 0.0905
R6734 VSS.n1836 VSS.n1833 0.0905
R6735 VSS.n1839 VSS.n1836 0.0905
R6736 VSS.n1842 VSS.n1839 0.0905
R6737 VSS.n1845 VSS.n1842 0.0905
R6738 VSS.n1848 VSS.n1845 0.0905
R6739 VSS.n1851 VSS.n1848 0.0905
R6740 VSS.n1854 VSS.n1851 0.0905
R6741 VSS.n1857 VSS.n1854 0.0905
R6742 VSS.n1860 VSS.n1857 0.0905
R6743 VSS.n1863 VSS.n1860 0.0905
R6744 VSS.n1888 VSS.n1863 0.0905
R6745 VSS.n1533 VSS.n1532 0.0905
R6746 VSS.n1749 VSS.n1747 0.0905
R6747 VSS.n1747 VSS.n1745 0.0905
R6748 VSS.n1745 VSS.n1743 0.0905
R6749 VSS.n1743 VSS.n1741 0.0905
R6750 VSS.n1738 VSS.n1736 0.0905
R6751 VSS.n1736 VSS.n1734 0.0905
R6752 VSS.n1731 VSS.n1729 0.0905
R6753 VSS.n1729 VSS.n1727 0.0905
R6754 VSS.n1724 VSS.n1722 0.0905
R6755 VSS.n1722 VSS.n1720 0.0905
R6756 VSS.n1720 VSS.n1718 0.0905
R6757 VSS.n1712 VSS.n1710 0.0905
R6758 VSS.n1710 VSS.n1708 0.0905
R6759 VSS.n1708 VSS.n1706 0.0905
R6760 VSS.n1706 VSS.n1704 0.0905
R6761 VSS.n1704 VSS.n1702 0.0905
R6762 VSS.n480 VSS.n478 0.0905
R6763 VSS.n911 VSS.n908 0.0905
R6764 VSS.n661 VSS.n659 0.0905
R6765 VSS.n632 VSS.n630 0.0905
R6766 VSS.n650 VSS.n648 0.0905
R6767 VSS.n319 VSS.n317 0.0905
R6768 VSS.n895 VSS.n892 0.0905
R6769 VSS.n806 VSS.n805 0.0905
R6770 VSS.n509 VSS.n506 0.0905
R6771 VSS.n525 VSS.n522 0.0905
R6772 VSS.n764 VSS.n762 0.0905
R6773 VSS.n757 VSS.n755 0.0905
R6774 VSS.n672 VSS.n670 0.0905
R6775 VSS.n748 VSS.n746 0.0905
R6776 VSS.n743 VSS.n741 0.0905
R6777 VSS.n738 VSS.n736 0.0905
R6778 VSS.n717 VSS.n715 0.0905
R6779 VSS.n413 VSS.n411 0.0905
R6780 VSS.n418 VSS.n416 0.0905
R6781 VSS.n423 VSS.n421 0.0905
R6782 VSS.n425 VSS.n423 0.0905
R6783 VSS.n430 VSS.n428 0.0905
R6784 VSS.n432 VSS.n430 0.0905
R6785 VSS.n437 VSS.n435 0.0905
R6786 VSS.n439 VSS.n437 0.0905
R6787 VSS.n441 VSS.n439 0.0905
R6788 VSS.n446 VSS.n444 0.0905
R6789 VSS.n448 VSS.n446 0.0905
R6790 VSS.n453 VSS.n451 0.0905
R6791 VSS.n455 VSS.n453 0.0905
R6792 VSS.n460 VSS.n458 0.0905
R6793 VSS.n469 VSS.n467 0.0905
R6794 VSS.n625 VSS.n623 0.0905
R6795 VSS.n410 VSS.n408 0.0905
R6796 VSS.n408 VSS.n406 0.0905
R6797 VSS.n406 VSS.n404 0.0905
R6798 VSS.n404 VSS.n402 0.0905
R6799 VSS.n402 VSS.n400 0.0905
R6800 VSS.n584 VSS.n582 0.0905
R6801 VSS.n586 VSS.n584 0.0905
R6802 VSS.n588 VSS.n586 0.0905
R6803 VSS.n590 VSS.n588 0.0905
R6804 VSS.n592 VSS.n590 0.0905
R6805 VSS.n594 VSS.n592 0.0905
R6806 VSS.n596 VSS.n594 0.0905
R6807 VSS.n598 VSS.n596 0.0905
R6808 VSS.n600 VSS.n598 0.0905
R6809 VSS.n602 VSS.n600 0.0905
R6810 VSS.n604 VSS.n602 0.0905
R6811 VSS.n606 VSS.n604 0.0905
R6812 VSS.n608 VSS.n606 0.0905
R6813 VSS.n610 VSS.n608 0.0905
R6814 VSS.n612 VSS.n610 0.0905
R6815 VSS.n614 VSS.n612 0.0905
R6816 VSS.n616 VSS.n614 0.0905
R6817 VSS.n618 VSS.n616 0.0905
R6818 VSS.n620 VSS.n618 0.0905
R6819 VSS.n622 VSS.n620 0.0905
R6820 VSS.n1343 VSS.n1341 0.0905
R6821 VSS.n1750 VSS.n1749 0.0895816
R6822 VSS.n1294 VSS.n1291 0.0895722
R6823 VSS.n22 VSS.n20 0.0895722
R6824 VSS.n1372 VSS.n1370 0.08915
R6825 VSS.n1590 VSS.n1589 0.0886443
R6826 VSS.n1159 VSS.n935 0.0877449
R6827 VSS.n819 VSS.n818 0.0877165
R6828 VSS.n1727 VSS.n1725 0.0868265
R6829 VSS.n1441 VSS.n1435 0.0858608
R6830 VSS.n1684 VSS.n1680 0.084933
R6831 VSS.n1183 VSS.n1180 0.084933
R6832 VSS.n1265 VSS.n1264 0.0840052
R6833 VSS.n2177 VSS.n2170 0.0840052
R6834 VSS.n504 VSS.n499 0.0831531
R6835 VSS.n1300 VSS.n1296 0.0830773
R6836 VSS.n7 VSS.n6 0.0830773
R6837 VSS.n115 VSS.n112 0.0821495
R6838 VSS.n16 VSS.n14 0.0821495
R6839 VSS.n1609 VSS.n1606 0.0812216
R6840 VSS.n433 VSS.n432 0.080398
R6841 VSS.n890 VSS.n889 0.0796667
R6842 VSS.n487 VSS.n480 0.0794796
R6843 VSS.n924 VSS.n922 0.0788281
R6844 VSS.n2118 VSS.n2086 0.07835
R6845 VSS.n889 VSS.n888 0.0778333
R6846 VSS.n444 VSS.n442 0.0776429
R6847 VSS.n578 VSS.n576 0.0776429
R6848 VSS.n52 VSS.n51 0.0756546
R6849 VSS.n922 VSS.n919 0.0748878
R6850 VSS.n1289 VSS.n1288 0.0747268
R6851 VSS.n1217 VSS.n1207 0.0747268
R6852 VSS.n89 VSS.n87 0.0747268
R6853 VSS.n542 VSS.n534 0.0747268
R6854 VSS.n1629 VSS.n1626 0.073799
R6855 VSS.n516 VSS.n513 0.0732992
R6856 VSS.n1216 VSS.n1214 0.0728711
R6857 VSS.n902 VSS.n900 0.0726849
R6858 VSS.n347 VSS.n346 0.0719433
R6859 VSS.n1381 VSS.n1217 0.0716
R6860 VSS.n1379 VSS.n1250 0.0716
R6861 VSS.n753 VSS.n752 0.0716
R6862 VSS.n627 VSS.n626 0.0716
R6863 VSS.n2013 VSS.n1982 0.0710155
R6864 VSS.n520 VSS.n378 0.0703456
R6865 VSS.n1716 VSS.n1712 0.0702959
R6866 VSS.n378 VSS.n377 0.0700876
R6867 VSS.n897 VSS.n895 0.0696134
R6868 VSS.n511 VSS.n509 0.068999
R6869 VSS.n1348 VSS.n1347 0.06845
R6870 VSS.n1358 VSS.n1357 0.06845
R6871 VSS.n2086 VSS.n2013 0.06845
R6872 VSS.n2043 VSS.n2042 0.06845
R6873 VSS.n2057 VSS.n2056 0.06845
R6874 VSS.n2071 VSS.n2070 0.06845
R6875 VSS.n2085 VSS.n2084 0.06845
R6876 VSS.n1370 VSS.n1369 0.06845
R6877 VSS.n1266 VSS.n1265 0.06845
R6878 VSS.n244 VSS.n243 0.0682606
R6879 VSS.n141 VSS.n135 0.0676429
R6880 VSS.n496 VSS.n488 0.0666364
R6881 VSS.n1644 VSS.n1643 0.0663763
R6882 VSS.n1385 VSS.n1384 0.0663286
R6883 VSS.n414 VSS.n413 0.0657041
R6884 VSS.n1161 VSS.n890 0.0656667
R6885 VSS.n360 VSS.n358 0.0654485
R6886 VSS VSS.n1163 0.0651667
R6887 VSS.n1383 VSS.n1176 0.0639126
R6888 VSS.n790 VSS.n789 0.0638673
R6889 VSS.n1160 VSS.n1159 0.0636667
R6890 VSS.n2084 VSS.n2079 0.0635928
R6891 VSS.n576 VSS.n573 0.0635
R6892 VSS.n1081 VSS.n1080 0.0635
R6893 VSS.n2187 VSS.n2186 0.0635
R6894 VSS.n1734 VSS.n1732 0.062949
R6895 VSS.n467 VSS.n465 0.062949
R6896 VSS.n770 VSS.n764 0.0620306
R6897 VSS.n758 VSS.n757 0.0620306
R6898 VSS.n456 VSS.n455 0.0620306
R6899 VSS.n73 VSS.n72 0.0617371
R6900 VSS.n127 VSS.n126 0.0617371
R6901 VSS.n1226 VSS.n1225 0.0608093
R6902 VSS.n1347 VSS.n1346 0.0608093
R6903 VSS.n1282 VSS.n1280 0.0608093
R6904 VSS.n2096 VSS.n2094 0.0598814
R6905 VSS.n325 VSS.n319 0.0592755
R6906 VSS.n1656 VSS.n1655 0.0589536
R6907 VSS.n367 VSS.n365 0.0589536
R6908 VSS.n638 VSS.n636 0.0583571
R6909 VSS.n732 VSS.n730 0.0583571
R6910 VSS.n421 VSS.n419 0.0583571
R6911 VSS.n65 VSS.n63 0.0580258
R6912 VSS.n39 VSS.n38 0.0570979
R6913 VSS.n659 VSS.n657 0.0565204
R6914 VSS.n741 VSS.n739 0.0565204
R6915 VSS.n426 VSS.n425 0.0565204
R6916 VSS.n497 VSS.n496 0.0564091
R6917 VSS.n2070 VSS.n2065 0.0561701
R6918 VSS.n1406 VSS.n1405 0.0552423
R6919 VSS.n1477 VSS.n1473 0.0533866
R6920 VSS.n334 VSS.n333 0.0533866
R6921 VSS.n72 VSS.n70 0.0533866
R6922 VSS.n1357 VSS.n1356 0.0533866
R6923 VSS.n1176 VSS.n1175 0.0529571
R6924 VSS.n782 VSS.n772 0.0528469
R6925 VSS.n789 VSS.n760 0.0528469
R6926 VSS.n675 VSS.n673 0.0528469
R6927 VSS.n751 VSS.n749 0.0528469
R6928 VSS.n451 VSS.n449 0.0528469
R6929 VSS.n1428 VSS.n1397 0.0524588
R6930 VSS.n2104 VSS.n2102 0.0524588
R6931 VSS.n2118 VSS.n2117 0.0524588
R6932 VSS.n1739 VSS.n1738 0.0519286
R6933 VSS.n1205 VSS.n1199 0.0506031
R6934 VSS.n2042 VSS.n2041 0.0506031
R6935 VSS.n495 VSS.n490 0.0500918
R6936 VSS.n529 VSS.n525 0.0500918
R6937 VSS.n1169 VSS.n1167 0.0496753
R6938 VSS.n1285 VSS.n1284 0.0496753
R6939 VSS.n670 VSS.n668 0.0491735
R6940 VSS.n746 VSS.n744 0.0491735
R6941 VSS.n2056 VSS.n2051 0.0487474
R6942 VSS.n628 VSS.n627 0.0482551
R6943 VSS.n753 VSS.n675 0.0473367
R6944 VSS.n752 VSS.n751 0.0473367
R6945 VSS.n369 VSS.n367 0.0468918
R6946 VSS.n1341 VSS.n1338 0.0468918
R6947 VSS.n151 VSS.n150 0.0462143
R6948 VSS.n1945 VSS.n1935 0.0459639
R6949 VSS.n1545 VSS.n1541 0.0459639
R6950 VSS.n1676 VSS.n1674 0.0459639
R6951 VSS.n2018 VSS.n2015 0.0459639
R6952 VSS.n20 VSS.n17 0.0459639
R6953 VSS.n832 VSS.n831 0.0459639
R6954 VSS.n1369 VSS.n1364 0.0459639
R6955 VSS.n1369 VSS.n1368 0.0459639
R6956 VSS.n1999 VSS.n1996 0.0459639
R6957 VSS.n1288 VSS.n1287 0.0459639
R6958 VSS.n2182 VSS.n2181 0.0459639
R6959 VSS.n1702 VSS.n1700 0.0455
R6960 VSS.n1890 VSS.n1888 0.0455
R6961 VSS.n471 VSS.n469 0.0455
R6962 VSS.n411 VSS.n410 0.0455
R6963 VSS.n623 VSS.n622 0.0455
R6964 VSS.n2112 VSS.n2110 0.0450361
R6965 VSS.n325 VSS.n315 0.0445816
R6966 VSS.n755 VSS.n753 0.0436633
R6967 VSS.n1374 VSS.n1372 0.0431804
R6968 VSS.n2110 VSS.n2106 0.0431804
R6969 VSS.n2056 VSS.n2055 0.0431804
R6970 VSS.n1167 VSS.n1166 0.0422526
R6971 VSS.n1287 VSS.n1285 0.0422526
R6972 VSS.n2042 VSS.n2038 0.0413247
R6973 VSS.n529 VSS.n528 0.0409082
R6974 VSS.n1388 VSS.n1385 0.0406143
R6975 VSS.n2179 VSS.n2177 0.0403969
R6976 VSS.n790 VSS.n546 0.0399898
R6977 VSS.n2120 VSS.n2118 0.0394691
R6978 VSS.n1741 VSS.n1739 0.0390714
R6979 VSS.n487 VSS.n482 0.0390714
R6980 VSS.n80 VSS.n79 0.0390714
R6981 VSS.n1564 VSS.n1560 0.0385412
R6982 VSS.n336 VSS.n334 0.0385412
R6983 VSS.n70 VSS.n69 0.0385412
R6984 VSS.n1357 VSS.n1354 0.0385412
R6985 VSS.n668 VSS.n661 0.0381531
R6986 VSS.n673 VSS.n672 0.0381531
R6987 VSS.n749 VSS.n748 0.0381531
R6988 VSS.n744 VSS.n743 0.0381531
R6989 VSS.n449 VSS.n448 0.0381531
R6990 VSS.n1383 VSS.n1382 0.037699
R6991 VSS.n1408 VSS.n1406 0.0366856
R6992 VSS.n2102 VSS.n2098 0.0357577
R6993 VSS.n2070 VSS.n2069 0.0357577
R6994 VSS.n1428 VSS.n1403 0.0357577
R6995 VSS.n506 VSS.n504 0.035398
R6996 VSS.n1477 VSS.n1468 0.0348299
R6997 VSS.n41 VSS.n39 0.0348299
R6998 VSS.n648 VSS.n646 0.0344796
R6999 VSS.n736 VSS.n734 0.0344796
R7000 VSS.n428 VSS.n426 0.0344796
R7001 VSS.n63 VSS.n62 0.0339021
R7002 VSS.n2127 VSS.n2124 0.0336891
R7003 VSS.n245 VSS.n244 0.0335116
R7004 VSS.n365 VSS.n364 0.0329742
R7005 VSS.n1391 VSS.n1390 0.0329
R7006 VSS.n919 VSS.n911 0.0326429
R7007 VSS.n636 VSS.n632 0.0326429
R7008 VSS.n730 VSS.n717 0.0326429
R7009 VSS.n419 VSS.n418 0.0326429
R7010 VSS.n1532 VSS.n1529 0.0317362
R7011 VSS.n476 VSS.n471 0.0317245
R7012 VSS.n1205 VSS.n1193 0.0311186
R7013 VSS.n1229 VSS.n1226 0.0311186
R7014 VSS.n1583 VSS.n1579 0.0311186
R7015 VSS.n1347 VSS.n1343 0.0311186
R7016 VSS.n1419 VSS.n1418 0.0311186
R7017 VSS.n1280 VSS.n1279 0.0311186
R7018 VSS.n657 VSS.n650 0.0308061
R7019 VSS.n739 VSS.n738 0.0308061
R7020 VSS.n927 VSS.n924 0.0302973
R7021 VSS.n906 VSS.n902 0.0302973
R7022 VSS.n519 VSS.n516 0.0302973
R7023 VSS.n1234 VSS.n1229 0.0301907
R7024 VSS.n1242 VSS.n1240 0.0301907
R7025 VSS.n127 VSS.n121 0.0301907
R7026 VSS.n646 VSS.n642 0.0298878
R7027 VSS.n734 VSS.n733 0.0298878
R7028 VSS.n932 VSS.n897 0.0296892
R7029 VSS.n520 VSS.n511 0.0293851
R7030 VSS.n772 VSS.n770 0.0289694
R7031 VSS.n760 VSS.n758 0.0289694
R7032 VSS.n458 VSS.n456 0.0289694
R7033 VSS.n2094 VSS.n2090 0.0283351
R7034 VSS.n2084 VSS.n2083 0.0283351
R7035 VSS.n1732 VSS.n1731 0.028051
R7036 VSS.n465 VSS.n460 0.028051
R7037 VSS.n358 VSS.n357 0.0264794
R7038 VSS.n931 VSS.n930 0.0263446
R7039 VSS.n155 VSS.n144 0.0262143
R7040 VSS.n261 VSS.n258 0.0258448
R7041 VSS.n197 VSS.n194 0.0258448
R7042 VSS.n200 VSS.n197 0.0258448
R7043 VSS.n203 VSS.n200 0.0258448
R7044 VSS.n210 VSS.n207 0.0258448
R7045 VSS.n213 VSS.n210 0.0258448
R7046 VSS.n216 VSS.n213 0.0258448
R7047 VSS.n219 VSS.n216 0.0258448
R7048 VSS.n226 VSS.n223 0.0258448
R7049 VSS.n229 VSS.n226 0.0258448
R7050 VSS.n835 VSS.n832 0.0258448
R7051 VSS.n844 VSS.n839 0.0258448
R7052 VSS.n847 VSS.n844 0.0258448
R7053 VSS.n854 VSS.n851 0.0258448
R7054 VSS.n857 VSS.n854 0.0258448
R7055 VSS.n860 VSS.n857 0.0258448
R7056 VSS.n863 VSS.n860 0.0258448
R7057 VSS.n870 VSS.n867 0.0258448
R7058 VSS.n873 VSS.n870 0.0258448
R7059 VSS.n884 VSS.n873 0.0258448
R7060 VSS.n887 VSS.n884 0.0258448
R7061 VSS.n1529 VSS.n1526 0.0257
R7062 VSS.n1526 VSS.n1523 0.0257
R7063 VSS.n1523 VSS.n1520 0.0257
R7064 VSS.n1516 VSS.n1513 0.0257
R7065 VSS.n1513 VSS.n1510 0.0257
R7066 VSS.n1770 VSS.n1767 0.0257
R7067 VSS.n1918 VSS.n1915 0.0257
R7068 VSS.n1915 VSS.n1912 0.0257
R7069 VSS.n1912 VSS.n1909 0.0257
R7070 VSS.n1905 VSS.n1902 0.0257
R7071 VSS.n1902 VSS.n1899 0.0257
R7072 VSS.n1899 VSS.n1896 0.0257
R7073 VSS.n1896 VSS.n1893 0.0257
R7074 VSS.n1893 VSS.n1890 0.0257
R7075 VSS.n416 VSS.n414 0.0252959
R7076 VSS.n630 VSS.n628 0.0252959
R7077 VSS.n715 VSS.n713 0.0252959
R7078 VSS.n132 VSS.n130 0.0247857
R7079 VSS.n1378 VSS.n1377 0.0246237
R7080 VSS.n2161 VSS.n2158 0.0245984
R7081 VSS.n2158 VSS.n2155 0.0245984
R7082 VSS.n2147 VSS.n2144 0.0245984
R7083 VSS.n2144 VSS.n2141 0.0245984
R7084 VSS.n2137 VSS.n2134 0.0245984
R7085 VSS.n2134 VSS.n2131 0.0245984
R7086 VSS.n2182 VSS.n2165 0.0243525
R7087 VSS.n888 VSS.n265 0.0237759
R7088 VSS.n1601 VSS.n1597 0.0236959
R7089 VSS.n1457 VSS.n1456 0.0236959
R7090 VSS.n642 VSS.n638 0.0234592
R7091 VSS.n733 VSS.n732 0.0234592
R7092 VSS.n162 VSS.n161 0.0233571
R7093 VSS.n1534 VSS.n1533 0.022768
R7094 VSS.n109 VSS.n107 0.0218402
R7095 VSS.n378 VSS.n372 0.0218402
R7096 VSS.n204 VSS.n203 0.0214483
R7097 VSS.n2155 VSS.n2152 0.0214016
R7098 VSS.n2138 VSS.n2137 0.0214016
R7099 VSS.n888 VSS.n292 0.0213333
R7100 VSS.n2024 VSS.n2020 0.0209124
R7101 VSS.n107 VSS.n91 0.0209124
R7102 VSS.n2013 VSS.n2012 0.0209124
R7103 VSS.n2151 VSS.n2148 0.0209098
R7104 VSS.n1718 VSS.n1716 0.0207041
R7105 VSS.n867 VSS.n864 0.0204138
R7106 VSS.n1906 VSS.n1905 0.0200429
R7107 VSS.n1534 VSS.n1484 0.0199845
R7108 VSS.n349 VSS.n347 0.0199845
R7109 VSS.n155 VSS.n154 0.0190714
R7110 VSS.n102 VSS.n101 0.0190714
R7111 VSS.n1214 VSS.n1213 0.0190567
R7112 VSS.n848 VSS.n847 0.0186034
R7113 VSS.n1091 VSS.n1088 0.0185738
R7114 VSS.n1098 VSS.n1095 0.0185738
R7115 VSS.n1101 VSS.n1098 0.0185738
R7116 VSS.n1108 VSS.n1105 0.0185738
R7117 VSS.n1111 VSS.n1108 0.0185738
R7118 VSS.n1118 VSS.n1115 0.0185738
R7119 VSS.n1121 VSS.n1118 0.0185738
R7120 VSS.n1124 VSS.n1121 0.0185738
R7121 VSS.n1131 VSS.n1128 0.0185738
R7122 VSS.n1134 VSS.n1131 0.0185738
R7123 VSS.n1141 VSS.n1138 0.0185738
R7124 VSS.n1144 VSS.n1141 0.0185738
R7125 VSS.n1151 VSS.n1148 0.0185738
R7126 VSS.n1391 VSS.n1388 0.0185
R7127 VSS.n1378 VSS.n1269 0.0181289
R7128 VSS.n1510 VSS.n1507 0.0179857
R7129 VSS.n627 VSS.n578 0.017949
R7130 VSS.n626 VSS.n625 0.017949
R7131 VSS.n1159 VSS.n1155 0.0177036
R7132 VSS.n242 VSS.n239 0.017569
R7133 VSS.n1920 VSS.n1919 0.0172143
R7134 VSS.n1217 VSS.n1216 0.017201
R7135 VSS.n542 VSS.n541 0.017201
R7136 VSS.n836 VSS.n835 0.0167931
R7137 VSS.n1112 VSS.n1111 0.0165451
R7138 VSS.n223 VSS.n220 0.0165345
R7139 VSS.n265 VSS.n262 0.0162759
R7140 VSS.n1619 VSS.n1615 0.0162732
R7141 VSS.n1291 VSS.n1289 0.0162732
R7142 VSS.n54 VSS.n52 0.0162732
R7143 VSS.n76 VSS.n73 0.0162732
R7144 VSS.n99 VSS.n98 0.0162143
R7145 VSS.n1084 VSS.n1081 0.0159918
R7146 VSS.n1128 VSS.n1125 0.0159918
R7147 VSS.n2165 VSS.n2162 0.0152541
R7148 VSS.n2128 VSS.n2127 0.0150082
R7149 VSS.n888 VSS.n887 0.0149828
R7150 VSS.n1517 VSS.n1516 0.0149
R7151 VSS.n1629 VSS.n1628 0.0144175
R7152 VSS.n1085 VSS.n1084 0.0135943
R7153 VSS.n87 VSS.n27 0.0134897
R7154 VSS.n442 VSS.n441 0.0133571
R7155 VSS.n576 VSS.n575 0.0133571
R7156 VSS.n1155 VSS.n1152 0.013041
R7157 VSS.n1145 VSS.n1144 0.0128566
R7158 VSS.n1553 VSS.n1552 0.0125619
R7159 VSS.n243 VSS.n242 0.0123966
R7160 VSS.n2186 VSS.n2185 0.0123033
R7161 VSS.n1095 VSS.n1092 0.0121189
R7162 VSS.n1102 VSS.n1101 0.01175
R7163 VSS.n1520 VSS.n1517 0.0113
R7164 VSS.n230 VSS.n229 0.0111034
R7165 VSS.n1138 VSS.n1135 0.0110123
R7166 VSS.n435 VSS.n433 0.010602
R7167 VSS.n155 VSS.n148 0.0103182
R7168 VSS.n2131 VSS.n2128 0.0100902
R7169 VSS.n262 VSS.n261 0.010069
R7170 VSS.n2162 VSS.n2161 0.00984426
R7171 VSS.n220 VSS.n219 0.00981034
R7172 VSS.n119 VSS.n115 0.00977835
R7173 VSS.n14 VSS.n13 0.00977835
R7174 VSS.n1457 VSS.n1454 0.00977835
R7175 VSS.n839 VSS.n836 0.00955172
R7176 VSS.n1639 VSS.n1635 0.00885052
R7177 VSS.n126 VSS.n123 0.00885052
R7178 VSS.n9 VSS.n7 0.00885052
R7179 VSS.n1441 VSS.n1440 0.00885052
R7180 VSS.n102 VSS.n96 0.0086
R7181 VSS.n83 VSS.n32 0.0086
R7182 VSS.n141 VSS.n140 0.0086
R7183 VSS.n1507 VSS.n1506 0.00821429
R7184 VSS.n148 VSS.n145 0.00813636
R7185 VSS.n1135 VSS.n1134 0.00806148
R7186 VSS.n1920 VSS.n1770 0.00795714
R7187 VSS.n1247 VSS.n1246 0.00792268
R7188 VSS.n1265 VSS.n1261 0.00792268
R7189 VSS.n851 VSS.n848 0.00774138
R7190 VSS.n165 VSS.n164 0.00764286
R7191 VSS.n83 VSS.n82 0.00764286
R7192 VSS.n1105 VSS.n1102 0.00732377
R7193 VSS.n1193 VSS.n1192 0.00699485
R7194 VSS.n1609 VSS.n1608 0.00699485
R7195 VSS.n1183 VSS.n1182 0.00699485
R7196 VSS.n1092 VSS.n1091 0.00695492
R7197 VSS.n96 VSS.n92 0.0068
R7198 VSS.n32 VSS.n28 0.0068
R7199 VSS.n140 VSS.n136 0.0068
R7200 VSS.n239 VSS.n238 0.00632512
R7201 VSS.n1384 VSS.n1383 0.00624272
R7202 VSS.n1148 VSS.n1145 0.00621721
R7203 VSS.n1909 VSS.n1906 0.00615714
R7204 VSS.n1751 VSS.n1750 0.00606701
R7205 VSS.n1152 VSS.n1151 0.00603279
R7206 VSS.n864 VSS.n863 0.00593103
R7207 VSS.n1088 VSS.n1085 0.00547951
R7208 VSS.n1302 VSS.n1300 0.00513918
R7209 VSS.n1572 VSS.n1571 0.00513918
R7210 VSS.n207 VSS.n204 0.00489655
R7211 VSS.n931 VSS.n927 0.0044527
R7212 VSS.n821 VSS.n819 0.00421134
R7213 VSS.n2148 VSS.n2147 0.00418852
R7214 VSS.n1725 VSS.n1724 0.00417347
R7215 VSS.n2152 VSS.n2151 0.00369672
R7216 VSS.n2141 VSS.n2138 0.00369672
R7217 VSS.n243 VSS.n230 0.00334483
R7218 VSS.n1684 VSS.n1666 0.00328351
R7219 VSS.n1081 VSS.n987 0.00308197
R7220 VSS.n1125 VSS.n1124 0.00308197
R7221 VSS.n1115 VSS.n1112 0.00252869
R7222 VSS VSS.n2187 0.0025
R7223 VSS.n1250 VSS.n1249 0.00235567
R7224 VSS.n1919 VSS.n1918 0.00152857
R7225 VSS.n1664 VSS.n1661 0.00142783
R7226 VSS.n806 VSS.n801 0.00142783
R7227 VSS.n520 VSS.n519 0.00141216
R7228 VSS.n932 VSS.n906 0.00110811
R7229 VSS.n1648 VSS.n1644 0.00095
R7230 VSS.n1630 VSS.n1629 0.00095
R7231 VSS.n1610 VSS.n1609 0.00095
R7232 VSS.n1592 VSS.n1590 0.00095
R7233 VSS.n1574 VSS.n1572 0.00095
R7234 VSS.n1555 VSS.n1553 0.00095
R7235 VSS.n1536 VSS.n1534 0.00095
R7236 VSS.n1657 VSS.n1656 0.00095
R7237 VSS.n1755 VSS.n1751 0.00095
R7238 VSS.n1458 VSS.n1457 0.00084749
R7239 VSS.n2177 VSS.n2176 0.00084749
R7240 VSS.n1443 VSS.n1441 0.000809278
R7241 VSS.n2185 VSS.n2182 0.000745902
R7242 OUT.n30 OUT.t17 55.2511
R7243 OUT.n17 OUT.t3 53.6484
R7244 OUT.n32 OUT.t13 52.4934
R7245 OUT.n15 OUT.t15 51.4031
R7246 OUT.n76 OUT.t60 50.0802
R7247 OUT.n179 OUT.t87 50.0802
R7248 OUT.n195 OUT.t9 50.0561
R7249 OUT.n1 OUT.t5 49.577
R7250 OUT.n1 OUT.t7 48.7525
R7251 OUT.n195 OUT.t11 48.2735
R7252 OUT.n60 OUT.t85 47.8988
R7253 OUT.n128 OUT.t77 47.8988
R7254 OUT.n85 OUT.t51 47.7394
R7255 OUT.n157 OUT.t55 47.7394
R7256 OUT.n38 OUT.t72 47.5312
R7257 OUT.n106 OUT.t67 47.5312
R7258 OUT.n75 OUT.t71 43.8005
R7259 OUT.n94 OUT.t47 43.8005
R7260 OUT.n96 OUT.t57 43.8005
R7261 OUT.n78 OUT.t65 43.8005
R7262 OUT.n80 OUT.t40 43.8005
R7263 OUT.n87 OUT.t52 43.8005
R7264 OUT.n89 OUT.t86 43.8005
R7265 OUT.n83 OUT.t39 43.8005
R7266 OUT.n178 OUT.t64 43.8005
R7267 OUT.n171 OUT.t41 43.8005
R7268 OUT.n173 OUT.t80 43.8005
R7269 OUT.n165 OUT.t46 43.8005
R7270 OUT.n167 OUT.t78 43.8005
R7271 OUT.n159 OUT.t58 43.8005
R7272 OUT.n161 OUT.t34 43.8005
R7273 OUT.n155 OUT.t73 43.8005
R7274 OUT.n36 OUT.t61 43.5398
R7275 OUT.n42 OUT.t49 43.5398
R7276 OUT.n40 OUT.t75 43.5398
R7277 OUT.n48 OUT.t62 43.5398
R7278 OUT.n46 OUT.t31 43.5398
R7279 OUT.n54 OUT.t83 43.5398
R7280 OUT.n52 OUT.t69 43.5398
R7281 OUT.n59 OUT.t38 43.5398
R7282 OUT.n104 OUT.t53 43.5398
R7283 OUT.n110 OUT.t44 43.5398
R7284 OUT.n108 OUT.t68 43.5398
R7285 OUT.n116 OUT.t56 43.5398
R7286 OUT.n114 OUT.t84 43.5398
R7287 OUT.n122 OUT.t76 43.5398
R7288 OUT.n120 OUT.t63 43.5398
R7289 OUT.n127 OUT.t32 43.5398
R7290 OUT.t60 OUT.n73 43.4094
R7291 OUT.t71 OUT.n74 43.4094
R7292 OUT.t47 OUT.n93 43.4094
R7293 OUT.t57 OUT.n95 43.4094
R7294 OUT.t65 OUT.n77 43.4094
R7295 OUT.t40 OUT.n79 43.4094
R7296 OUT.t52 OUT.n86 43.4094
R7297 OUT.t86 OUT.n88 43.4094
R7298 OUT.t39 OUT.n82 43.4094
R7299 OUT.t61 OUT.n35 43.4094
R7300 OUT.t49 OUT.n41 43.4094
R7301 OUT.t75 OUT.n39 43.4094
R7302 OUT.t62 OUT.n47 43.4094
R7303 OUT.t31 OUT.n45 43.4094
R7304 OUT.t83 OUT.n53 43.4094
R7305 OUT.t69 OUT.n51 43.4094
R7306 OUT.t38 OUT.n58 43.4094
R7307 OUT.t85 OUT.n57 43.4094
R7308 OUT.t72 OUT.n37 43.4094
R7309 OUT.t51 OUT.n84 43.4094
R7310 OUT.t87 OUT.n176 43.4094
R7311 OUT.t64 OUT.n177 43.4094
R7312 OUT.t41 OUT.n170 43.4094
R7313 OUT.t80 OUT.n172 43.4094
R7314 OUT.t46 OUT.n164 43.4094
R7315 OUT.t78 OUT.n166 43.4094
R7316 OUT.t58 OUT.n158 43.4094
R7317 OUT.t34 OUT.n160 43.4094
R7318 OUT.t73 OUT.n154 43.4094
R7319 OUT.t53 OUT.n103 43.4094
R7320 OUT.t44 OUT.n109 43.4094
R7321 OUT.t68 OUT.n107 43.4094
R7322 OUT.t56 OUT.n115 43.4094
R7323 OUT.t84 OUT.n113 43.4094
R7324 OUT.t76 OUT.n121 43.4094
R7325 OUT.t63 OUT.n119 43.4094
R7326 OUT.t32 OUT.n126 43.4094
R7327 OUT.t77 OUT.n125 43.4094
R7328 OUT.t67 OUT.n105 43.4094
R7329 OUT.t55 OUT.n156 43.4094
R7330 OUT.n57 OUT.t45 43.2791
R7331 OUT.n74 OUT.t54 43.2791
R7332 OUT.n51 OUT.t30 43.2791
R7333 OUT.n53 OUT.t42 43.2791
R7334 OUT.n77 OUT.t48 43.2791
R7335 OUT.n47 OUT.t81 43.2791
R7336 OUT.n86 OUT.t35 43.2791
R7337 OUT.n41 OUT.t66 43.2791
R7338 OUT.n37 OUT.t33 43.2791
R7339 OUT.n35 OUT.t79 43.2791
R7340 OUT.n125 OUT.t37 43.2791
R7341 OUT.n177 OUT.t50 43.2791
R7342 OUT.n170 OUT.t82 43.2791
R7343 OUT.n172 OUT.t36 43.2791
R7344 OUT.n164 OUT.t43 43.2791
R7345 OUT.n166 OUT.t74 43.2791
R7346 OUT.n158 OUT.t89 43.2791
R7347 OUT.n109 OUT.t59 43.2791
R7348 OUT.n156 OUT.t88 43.2791
R7349 OUT.n154 OUT.t70 43.2791
R7350 OUT.n49 OUT.n46 4.88467
R7351 OUT.n117 OUT.n114 4.88467
R7352 OUT.n43 OUT.n40 4.72712
R7353 OUT.n111 OUT.n108 4.72712
R7354 OUT.n81 OUT.n78 4.56957
R7355 OUT.n168 OUT.n165 4.56957
R7356 OUT.n85 OUT.n83 4.46453
R7357 OUT.n157 OUT.n155 4.46453
R7358 OUT.n38 OUT.n36 4.41201
R7359 OUT.n106 OUT.n104 4.41201
R7360 OUT.n90 OUT.n89 4.35949
R7361 OUT.n162 OUT.n161 4.35949
R7362 OUT.n55 OUT.n52 4.30697
R7363 OUT.n123 OUT.n120 4.30697
R7364 OUT.n185 OUT.n184 4.283
R7365 OUT.n97 OUT.n94 4.25446
R7366 OUT.n174 OUT.n171 4.25446
R7367 OUT.n97 OUT.n96 4.14942
R7368 OUT.n174 OUT.n173 4.14942
R7369 OUT.n55 OUT.n54 4.0969
R7370 OUT.n123 OUT.n122 4.0969
R7371 OUT.n60 OUT.n59 4.04439
R7372 OUT.n90 OUT.n87 4.04439
R7373 OUT.n128 OUT.n127 4.04439
R7374 OUT.n162 OUT.n159 4.04439
R7375 OUT.n197 OUT.n195 4.0005
R7376 OUT.n2 OUT.n1 4.0005
R7377 OUT.n76 OUT.n75 3.88683
R7378 OUT.n179 OUT.n178 3.88683
R7379 OUT.n91 OUT.n85 3.86999
R7380 OUT.n163 OUT.n157 3.86999
R7381 OUT.n31 OUT.n29 3.86659
R7382 OUT.n112 OUT.n106 3.86201
R7383 OUT.n44 OUT.n38 3.85966
R7384 OUT.n16 OUT.n14 3.83724
R7385 OUT.n81 OUT.n80 3.83431
R7386 OUT.n168 OUT.n167 3.83431
R7387 OUT.n43 OUT.n42 3.67676
R7388 OUT.n111 OUT.n110 3.67676
R7389 OUT.n61 OUT.n60 3.62694
R7390 OUT.n56 OUT.n55 3.62694
R7391 OUT.n44 OUT.n43 3.62694
R7392 OUT.n91 OUT.n90 3.62694
R7393 OUT.n98 OUT.n97 3.62694
R7394 OUT.n118 OUT.n117 3.62694
R7395 OUT.n163 OUT.n162 3.62694
R7396 OUT.n92 OUT.n81 3.62672
R7397 OUT.n99 OUT.n76 3.62672
R7398 OUT.n129 OUT.n128 3.62672
R7399 OUT.n180 OUT.n179 3.62672
R7400 OUT.n175 OUT.n174 3.62672
R7401 OUT.n169 OUT.n168 3.62672
R7402 OUT.n50 OUT.n49 3.62642
R7403 OUT.n112 OUT.n111 3.62642
R7404 OUT.n124 OUT.n123 3.62642
R7405 OUT.n49 OUT.n48 3.51921
R7406 OUT.n117 OUT.n116 3.51921
R7407 OUT.n186 OUT.n26 3.45519
R7408 OUT.n189 OUT.n22 3.37867
R7409 OUT.n187 OUT.n24 3.23061
R7410 OUT.n199 OUT.n198 3.02196
R7411 OUT.n201 OUT.n200 2.6005
R7412 OUT.n18 OUT.n16 2.32876
R7413 OUT.n33 OUT.n31 2.31115
R7414 OUT.n137 OUT.t0 2.28772
R7415 OUT.n136 OUT.t29 2.27583
R7416 OUT.n190 OUT.n189 1.83428
R7417 OUT.n185 OUT.n34 1.71595
R7418 OUT.n11 OUT.n10 1.63529
R7419 OUT.n142 OUT.n141 1.14106
R7420 OUT.n64 OUT.n63 1.1255
R7421 OUT.n69 OUT.n68 1.1255
R7422 OUT.n72 OUT.n71 1.1255
R7423 OUT.n102 OUT.n101 1.1255
R7424 OUT.n132 OUT.n131 1.1255
R7425 OUT.n143 OUT.n142 1.1255
R7426 OUT.n145 OUT.n144 1.1255
R7427 OUT.n148 OUT.n147 1.1255
R7428 OUT.n151 OUT.n150 1.1255
R7429 OUT.n193 OUT.n192 1.1255
R7430 OUT.n192 OUT.n191 1.11366
R7431 OUT.n184 OUT.n183 1.11352
R7432 OUT.n21 OUT.n20 1.04336
R7433 OUT.n64 OUT.n62 0.972114
R7434 OUT.n34 OUT.n27 0.933803
R7435 OUT.n5 OUT.n4 0.837772
R7436 OUT OUT.n203 0.768041
R7437 OUT.n187 OUT.n186 0.712763
R7438 OUT.n181 OUT.n180 0.677331
R7439 OUT.n10 OUT.t6 0.607167
R7440 OUT.n10 OUT.n9 0.607167
R7441 OUT.n4 OUT.t8 0.607167
R7442 OUT.n4 OUT.n3 0.607167
R7443 OUT.n200 OUT.t24 0.607167
R7444 OUT.n200 OUT.t10 0.607167
R7445 OUT.n198 OUT.t28 0.607167
R7446 OUT.n198 OUT.t12 0.607167
R7447 OUT.n26 OUT.t26 0.5465
R7448 OUT.n26 OUT.n25 0.5465
R7449 OUT.n24 OUT.t21 0.5465
R7450 OUT.n24 OUT.n23 0.5465
R7451 OUT.n14 OUT.t16 0.5465
R7452 OUT.n14 OUT.n13 0.5465
R7453 OUT.n20 OUT.t23 0.5465
R7454 OUT.n20 OUT.t4 0.5465
R7455 OUT.n27 OUT.t20 0.5465
R7456 OUT.n27 OUT.t14 0.5465
R7457 OUT.n29 OUT.t18 0.5465
R7458 OUT.n29 OUT.n28 0.5465
R7459 OUT OUT.n194 0.545119
R7460 OUT.n188 OUT.n187 0.54055
R7461 OUT.n62 OUT.n61 0.536124
R7462 OUT.n186 OUT.n185 0.535757
R7463 OUT.n100 OUT.n99 0.522126
R7464 OUT.n130 OUT.n129 0.519913
R7465 OUT.n202 OUT.n201 0.507573
R7466 OUT.n201 OUT.n199 0.435134
R7467 OUT.n143 OUT.n132 0.423314
R7468 OUT.n137 OUT.n136 0.421821
R7469 OUT.n102 OUT.n72 0.36188
R7470 OUT.n34 OUT.n33 0.332105
R7471 OUT.n31 OUT.n30 0.277411
R7472 OUT.n7 OUT.n6 0.254037
R7473 OUT.n124 OUT.n118 0.248269
R7474 OUT.n56 OUT.n50 0.247603
R7475 OUT.n175 OUT.n169 0.24375
R7476 OUT.n98 OUT.n92 0.243505
R7477 OUT.n129 OUT.n124 0.238996
R7478 OUT.n50 OUT.n44 0.237941
R7479 OUT.n61 OUT.n56 0.237592
R7480 OUT.n118 OUT.n112 0.237275
R7481 OUT.n180 OUT.n175 0.235635
R7482 OUT.n99 OUT.n98 0.234886
R7483 OUT.n92 OUT.n91 0.231198
R7484 OUT.n169 OUT.n163 0.231198
R7485 OUT.n19 OUT.n18 0.21963
R7486 OUT.n6 OUT.n5 0.216907
R7487 OUT.n153 OUT.n151 0.192005
R7488 OUT.n8 OUT.n7 0.173915
R7489 OUT.n22 OUT.n21 0.169406
R7490 OUT.n101 OUT.n100 0.164572
R7491 OUT.n131 OUT.n130 0.163731
R7492 OUT.n33 OUT.n32 0.160935
R7493 OUT.n18 OUT.n17 0.158978
R7494 OUT.n16 OUT.n15 0.157022
R7495 OUT.n189 OUT.n188 0.130578
R7496 OUT.n197 OUT.n196 0.122534
R7497 OUT.n2 OUT.n0 0.121008
R7498 OUT.n193 OUT.n11 0.107094
R7499 OUT.n192 OUT.n12 0.10705
R7500 OUT.n203 OUT.n202 0.101492
R7501 OUT.n22 OUT.n19 0.0813159
R7502 OUT.n6 OUT.n2 0.0615169
R7503 OUT.n199 OUT.n197 0.0554153
R7504 OUT.n194 OUT.n193 0.0528411
R7505 OUT.n65 OUT.n64 0.0468918
R7506 OUT.n72 OUT.n69 0.0468918
R7507 OUT.n145 OUT.n143 0.0468918
R7508 OUT.n151 OUT.n148 0.0468918
R7509 OUT.n132 OUT.n102 0.0455
R7510 OUT.n68 OUT.n67 0.0453454
R7511 OUT.n69 OUT.n65 0.0453454
R7512 OUT.n148 OUT.n145 0.0453454
R7513 OUT.n138 OUT.n137 0.0374422
R7514 OUT.n136 OUT.n135 0.0369463
R7515 OUT.n191 OUT.n190 0.0329324
R7516 OUT.n147 OUT.n146 0.0306981
R7517 OUT.n184 OUT.n153 0.0275
R7518 OUT.n183 OUT.n181 0.0259538
R7519 OUT.n183 OUT.n182 0.0259538
R7520 OUT.n67 OUT.n66 0.024329
R7521 OUT.n71 OUT.n70 0.0239592
R7522 OUT.n11 OUT.n8 0.0227109
R7523 OUT.n153 OUT.n152 0.0185
R7524 OUT.n150 OUT.n149 0.0163584
R7525 OUT.n134 OUT.n133 0.0125661
R7526 OUT.n141 OUT.n139 0.00711157
R7527 OUT.n141 OUT.n140 0.00595455
R7528 OUT.n139 OUT.n138 0.000830579
R7529 OUT.n135 OUT.n134 0.000830579
R7530 IBIAS.n33 IBIAS.t20 30.6996
R7531 IBIAS.n34 IBIAS.t35 30.6996
R7532 IBIAS.n47 IBIAS.t38 29.7219
R7533 IBIAS.n54 IBIAS.t30 29.5264
R7534 IBIAS.n55 IBIAS.t40 29.5264
R7535 IBIAS.n57 IBIAS.t25 28.6139
R7536 IBIAS.n54 IBIAS.t22 28.6139
R7537 IBIAS.n55 IBIAS.t33 28.6139
R7538 IBIAS.n56 IBIAS.t14 28.6139
R7539 IBIAS.n47 IBIAS.t17 28.5487
R7540 IBIAS.n11 IBIAS.t41 28.2228
R7541 IBIAS.n42 IBIAS.t21 27.8317
R7542 IBIAS.n33 IBIAS.t36 27.4407
R7543 IBIAS.n34 IBIAS.t26 27.4407
R7544 IBIAS.n36 IBIAS.t34 27.4407
R7545 IBIAS.n37 IBIAS.t39 27.4407
R7546 IBIAS.n52 IBIAS.t31 27.1148
R7547 IBIAS.n22 IBIAS.t23 24.3089
R7548 IBIAS.n72 IBIAS.t37 24.0514
R7549 IBIAS.n0 IBIAS.t10 24.0514
R7550 IBIAS.n65 IBIAS.t9 23.921
R7551 IBIAS.n68 IBIAS.t44 23.921
R7552 IBIAS.n72 IBIAS.t43 23.921
R7553 IBIAS.n2 IBIAS.t7 23.921
R7554 IBIAS.n5 IBIAS.t29 23.921
R7555 IBIAS.n0 IBIAS.t28 23.921
R7556 IBIAS.n73 IBIAS.t12 23.921
R7557 IBIAS.n69 IBIAS.t13 23.921
R7558 IBIAS.n6 IBIAS.t16 23.921
R7559 IBIAS.n1 IBIAS.t15 23.921
R7560 IBIAS.n67 IBIAS.t18 23.7907
R7561 IBIAS.n4 IBIAS.t42 23.7907
R7562 IBIAS.n80 IBIAS.t19 19.5541
R7563 IBIAS.n63 IBIAS.t27 19.5541
R7564 IBIAS.n23 IBIAS.t6 19.163
R7565 IBIAS.n22 IBIAS.t32 19.0326
R7566 IBIAS.n20 IBIAS.t24 19.0326
R7567 IBIAS.n11 IBIAS.t11 15.9041
R7568 IBIAS.n12 IBIAS.t2 15.9041
R7569 IBIAS.n29 IBIAS.t4 15.9041
R7570 IBIAS.n21 IBIAS.t0 15.513
R7571 IBIAS.n20 IBIAS.n19 12.9251
R7572 IBIAS.n12 IBIAS.n11 12.3193
R7573 IBIAS.n29 IBIAS.n28 12.3193
R7574 IBIAS.n21 IBIAS.n20 11.897
R7575 IBIAS.n55 IBIAS.n54 10.8005
R7576 IBIAS.n57 IBIAS.n56 10.8005
R7577 IBIAS.n45 IBIAS.n44 10.8005
R7578 IBIAS.n46 IBIAS.n45 10.8005
R7579 IBIAS.n34 IBIAS.n33 10.8005
R7580 IBIAS.n48 IBIAS.n47 10.7505
R7581 IBIAS.n38 IBIAS.n37 10.7505
R7582 IBIAS.n73 IBIAS.n72 10.4005
R7583 IBIAS.n69 IBIAS.n68 10.4005
R7584 IBIAS.n66 IBIAS.n65 10.4005
R7585 IBIAS.n1 IBIAS.n0 10.4005
R7586 IBIAS.n6 IBIAS.n5 10.4005
R7587 IBIAS.n3 IBIAS.n2 10.4005
R7588 IBIAS.n58 IBIAS.n55 9.3005
R7589 IBIAS.n23 IBIAS.n22 7.77919
R7590 IBIAS.n24 IBIAS.n23 6.40568
R7591 IBIAS.n35 IBIAS.n34 5.4005
R7592 IBIAS.n71 IBIAS.n67 5.27954
R7593 IBIAS.n7 IBIAS.n4 5.27781
R7594 IBIAS.n16 IBIAS.n15 4.5005
R7595 IBIAS.n84 IBIAS.n83 4.5005
R7596 IBIAS.n39 IBIAS.n35 4.11457
R7597 IBIAS.n59 IBIAS.n58 4.0077
R7598 IBIAS.n39 IBIAS.n38 4.0005
R7599 IBIAS.n51 IBIAS.n50 4.0005
R7600 IBIAS.n49 IBIAS.n48 4.0005
R7601 IBIAS.n43 IBIAS.n42 4.0005
R7602 IBIAS.n41 IBIAS.n40 4.0005
R7603 IBIAS.n53 IBIAS.n52 4.0005
R7604 IBIAS.n25 IBIAS.n24 4.0005
R7605 IBIAS.n75 IBIAS.n74 4.0005
R7606 IBIAS.n71 IBIAS.n70 4.0005
R7607 IBIAS.n8 IBIAS.n1 4.0005
R7608 IBIAS.n7 IBIAS.n6 4.0005
R7609 IBIAS.n25 IBIAS.t1 3.91084
R7610 IBIAS.n24 IBIAS.n21 3.85789
R7611 IBIAS.n31 IBIAS.n30 2.8805
R7612 IBIAS.n77 IBIAS.n64 2.8805
R7613 IBIAS.n30 IBIAS.n29 2.79503
R7614 IBIAS.n62 IBIAS.n60 2.70728
R7615 IBIAS.n26 IBIAS.n18 2.6005
R7616 IBIAS.n81 IBIAS.n80 2.35719
R7617 IBIAS.n60 IBIAS.n59 2.29351
R7618 IBIAS.n60 IBIAS.n32 1.98864
R7619 IBIAS.n15 IBIAS.n12 1.93956
R7620 IBIAS.n14 IBIAS.n13 1.54034
R7621 IBIAS.n58 IBIAS.n57 1.5005
R7622 IBIAS.n43 IBIAS.n41 1.47165
R7623 IBIAS.n53 IBIAS.n51 1.43012
R7624 IBIAS.n83 IBIAS.n82 1.3855
R7625 IBIAS.n75 IBIAS.n71 1.27954
R7626 IBIAS.n8 IBIAS.n7 1.27435
R7627 IBIAS.n76 IBIAS.n75 1.25103
R7628 IBIAS.n87 IBIAS.n8 1.24838
R7629 IBIAS.n64 IBIAS.n63 0.977665
R7630 IBIAS.n79 IBIAS.n62 0.945657
R7631 IBIAS.n26 IBIAS.n25 0.942312
R7632 IBIAS.n18 IBIAS.t3 0.9105
R7633 IBIAS.n18 IBIAS.n17 0.9105
R7634 IBIAS.n32 IBIAS.n16 0.782929
R7635 IBIAS.n32 IBIAS.n31 0.779848
R7636 IBIAS.n27 IBIAS.n26 0.421045
R7637 IBIAS.n74 IBIAS.n73 0.261214
R7638 IBIAS.n49 IBIAS.n43 0.185692
R7639 IBIAS.n82 IBIAS.n81 0.172941
R7640 IBIAS.n15 IBIAS.n14 0.171594
R7641 IBIAS.n51 IBIAS.n49 0.166654
R7642 IBIAS.n59 IBIAS.n53 0.161415
R7643 IBIAS.n41 IBIAS.n39 0.137231
R7644 IBIAS.n67 IBIAS.n66 0.130857
R7645 IBIAS.n4 IBIAS.n3 0.130857
R7646 IBIAS.n79 IBIAS.n78 0.0851369
R7647 IBIAS.n70 IBIAS.n69 0.0656786
R7648 IBIAS.n48 IBIAS.n46 0.0505
R7649 IBIAS.n38 IBIAS.n36 0.0505
R7650 IBIAS.n87 IBIAS.n86 0.046625
R7651 IBIAS.n31 IBIAS.n27 0.0246667
R7652 IBIAS.n84 IBIAS.n79 0.023695
R7653 IBIAS.n85 IBIAS.n84 0.023
R7654 IBIAS.n62 IBIAS.n61 0.0189615
R7655 IBIAS.n78 IBIAS.n77 0.0186513
R7656 IBIAS.n10 IBIAS.n9 0.01175
R7657 IBIAS IBIAS.n87 0.00725
R7658 IBIAS.n86 IBIAS.n85 0.003875
R7659 IBIAS.n77 IBIAS.n76 0.00325363
R7660 IBIAS.n16 IBIAS.n10 0.00175
R7661 VBS3.n42 VBS3.t17 56.0541
R7662 VBS3.n42 VBS3.t10 55.5326
R7663 VBS3.n43 VBS3.t18 47.3201
R7664 VBS3.n44 VBS3.t11 47.3201
R7665 VBS3.n46 VBS3.t21 47.3201
R7666 VBS3.n45 VBS3.t8 47.3201
R7667 VBS3.n44 VBS3.t24 47.3201
R7668 VBS3.n46 VBS3.t14 47.3201
R7669 VBS3.n52 VBS3.t9 47.3201
R7670 VBS3.n49 VBS3.t19 47.3201
R7671 VBS3.n50 VBS3.t13 47.3201
R7672 VBS3.n50 VBS3.t16 47.3201
R7673 VBS3.n51 VBS3.t12 47.3201
R7674 VBS3.n51 VBS3.t15 47.3201
R7675 VBS3.n52 VBS3.t22 47.3201
R7676 VBS3.n45 VBS3.t23 47.3201
R7677 VBS3.n50 VBS3.n49 18.8981
R7678 VBS3.n52 VBS3.n51 18.8981
R7679 VBS3.n42 VBS3.n41 18.8981
R7680 VBS3.n40 VBS3.n39 18.8981
R7681 VBS3.n44 VBS3.n43 18.8981
R7682 VBS3.n46 VBS3.n45 18.8981
R7683 VBS3.n27 VBS3.t0 17.8034
R7684 VBS3.n48 VBS3.n42 17.4226
R7685 VBS3.n23 VBS3.t2 17.2468
R7686 VBS3.n41 VBS3.n40 9.41985
R7687 VBS3.n48 VBS3.n47 6.66569
R7688 VBS3.n54 VBS3.n53 6.13751
R7689 VBS3.n47 VBS3.n44 5.12227
R7690 VBS3.n53 VBS3.n52 4.82792
R7691 VBS3.n53 VBS3.n50 4.59244
R7692 VBS3.n12 VBS3.n11 4.50092
R7693 VBS3.n38 VBS3.n34 4.5005
R7694 VBS3.n38 VBS3.n37 4.5005
R7695 VBS3.n20 VBS3.n19 4.5005
R7696 VBS3.n18 VBS3.n17 4.5005
R7697 VBS3.n15 VBS3.n14 4.5005
R7698 VBS3.n47 VBS3.n46 4.29808
R7699 VBS3.n31 VBS3.n26 3.56947
R7700 VBS3.n34 VBS3.n33 2.2505
R7701 VBS3.n2 VBS3.n1 2.08733
R7702 VBS3.n11 VBS3.n10 1.50499
R7703 VBS3.n4 VBS3.n3 1.49676
R7704 VBS3.n9 VBS3.n8 1.4966
R7705 VBS3.n28 VBS3.n27 1.43031
R7706 VBS3.n24 VBS3.n23 1.42468
R7707 VBS3.n6 VBS3.t7 0.9105
R7708 VBS3.n6 VBS3.n5 0.9105
R7709 VBS3.n1 VBS3.t4 0.9105
R7710 VBS3.n1 VBS3.n0 0.9105
R7711 VBS3 VBS3.n54 0.824379
R7712 VBS3.n26 VBS3.t3 0.8195
R7713 VBS3.n26 VBS3.n25 0.8195
R7714 VBS3.n7 VBS3.n6 0.805572
R7715 VBS3.n54 VBS3.n48 0.4185
R7716 VBS3.n8 VBS3.n7 0.0613454
R7717 VBS3.n32 VBS3.n31 0.0365
R7718 VBS3.n31 VBS3.n30 0.0275
R7719 VBS3 VBS3.n38 0.0269953
R7720 VBS3.n30 VBS3.n29 0.0212
R7721 VBS3.n33 VBS3.n32 0.0194
R7722 VBS3.n9 VBS3.n4 0.0144547
R7723 VBS3.n10 VBS3.n9 0.0141896
R7724 VBS3.n4 VBS3.n2 0.0137198
R7725 VBS3.n22 VBS3.n21 0.00900394
R7726 VBS3.n33 VBS3.n24 0.0086
R7727 VBS3.n13 VBS3.n12 0.00849065
R7728 VBS3.n29 VBS3.n28 0.0068
R7729 VBS3.n34 VBS3.n22 0.00655042
R7730 VBS3.n17 VBS3.n16 0.00503782
R7731 VBS3.n15 VBS3.n13 0.00428505
R7732 VBS3.n37 VBS3.n36 0.00262598
R7733 VBS3.n20 VBS3.n18 0.00218224
R7734 VBS3.n18 VBS3.n15 0.00134112
R7735 VBS3.n36 VBS3.n35 0.00120866
R7736 VBS3.n38 VBS3.n20 0.000920561
R7737 VBS2.n6 VBS2.t7 70.1735
R7738 VBS2.n12 VBS2.t6 45.8988
R7739 VBS2.n8 VBS2.t9 44.8434
R7740 VBS2.n9 VBS2.t11 44.8434
R7741 VBS2.n6 VBS2.t10 44.8434
R7742 VBS2.n10 VBS2.t5 44.8434
R7743 VBS2.n7 VBS2.t4 44.8434
R7744 VBS2.n11 VBS2.t8 44.8434
R7745 VBS2.t6 VBS2.n11 44.8434
R7746 VBS2.n12 VBS2.n7 24.2752
R7747 VBS2.n9 VBS2.n8 22.8527
R7748 VBS2.n11 VBS2.n10 22.8527
R7749 VBS2.n18 VBS2.t1 20.237
R7750 VBS2.n15 VBS2.n12 16.3334
R7751 VBS2.n7 VBS2.n6 14.0728
R7752 VBS2.n10 VBS2.n9 12.6962
R7753 VBS2.n20 VBS2.n19 5.11604
R7754 VBS2.n16 VBS2.n15 4.5005
R7755 VBS2.n20 VBS2.t0 4.44846
R7756 VBS2.n18 VBS2.t2 3.90373
R7757 VBS2.n22 VBS2.n21 3.5729
R7758 VBS2.n23 VBS2.n17 2.24666
R7759 VBS2.n14 VBS2.n13 2.22224
R7760 VBS2.n21 VBS2.n18 1.78171
R7761 VBS2.n21 VBS2.n20 1.27289
R7762 VBS2.n15 VBS2.n14 0.317891
R7763 VBS2.n4 VBS2.n3 0.0548396
R7764 VBS2.n5 VBS2.n4 0.0242736
R7765 VBS2.n27 VBS2.n0 0.0167
R7766 VBS2.n2 VBS2.n1 0.014934
R7767 VBS2.n3 VBS2.n2 0.0132358
R7768 VBS2 VBS2.n28 0.0106887
R7769 VBS2.n23 VBS2.n22 0.0102832
R7770 VBS2.n28 VBS2.n27 0.00983962
R7771 VBS2.n24 VBS2.n23 0.00968321
R7772 VBS2.n17 VBS2.n16 0.00474528
R7773 VBS2.n16 VBS2.n5 0.00389623
R7774 VBS2.n27 VBS2.n26 0.0011
R7775 VBS2.n26 VBS2.n25 0.0011
R7776 VBS2.n25 VBS2.n24 0.0011
R7777 VX.n35 VX.t0 52.4934
R7778 VX.n51 VX.t2 52.1689
R7779 VX.n38 VX.t4 51.5691
R7780 VX.n45 VX.t6 50.3958
R7781 VX.n5 VX.t49 45.8862
R7782 VX.n6 VX.t40 45.8862
R7783 VX.n7 VX.t31 45.8862
R7784 VX.n8 VX.t46 45.8862
R7785 VX.n12 VX.t38 45.8862
R7786 VX.n11 VX.t20 45.8862
R7787 VX.n10 VX.t48 45.8862
R7788 VX.n9 VX.t39 45.8862
R7789 VX.n5 VX.t29 45.6255
R7790 VX.n6 VX.t23 45.6255
R7791 VX.n7 VX.t44 45.6255
R7792 VX.n8 VX.t25 45.6255
R7793 VX.n12 VX.t51 45.6255
R7794 VX.n11 VX.t32 45.6255
R7795 VX.n10 VX.t27 45.6255
R7796 VX.n19 VX.t47 45.6255
R7797 VX.n14 VX.t26 45.6255
R7798 VX.n23 VX.t45 45.6255
R7799 VX.n15 VX.t36 45.6255
R7800 VX.n24 VX.t37 45.6255
R7801 VX.n16 VX.t30 45.6255
R7802 VX.n25 VX.t28 45.6255
R7803 VX.n17 VX.t43 45.6255
R7804 VX.n26 VX.t41 45.6255
R7805 VX.n21 VX.t22 45.6255
R7806 VX.n30 VX.t34 45.6255
R7807 VX.n20 VX.t33 45.6255
R7808 VX.n29 VX.t50 45.6255
R7809 VX.n18 VX.t24 45.6255
R7810 VX.n27 VX.t35 45.6255
R7811 VX.n28 VX.t42 45.6255
R7812 VX.n9 VX.t21 45.6255
R7813 VX.n15 VX.n14 11.9189
R7814 VX.n16 VX.n15 11.9189
R7815 VX.n17 VX.n16 11.9189
R7816 VX.n21 VX.n20 11.9189
R7817 VX.n20 VX.n19 11.9189
R7818 VX.n19 VX.n18 11.9189
R7819 VX.n24 VX.n23 11.9189
R7820 VX.n25 VX.n24 11.9189
R7821 VX.n26 VX.n25 11.9189
R7822 VX.n30 VX.n29 11.9189
R7823 VX.n29 VX.n28 11.9189
R7824 VX.n28 VX.n27 11.9189
R7825 VX.n6 VX.n5 11.9189
R7826 VX.n7 VX.n6 11.9189
R7827 VX.n8 VX.n7 11.9189
R7828 VX.n12 VX.n11 11.9189
R7829 VX.n11 VX.n10 11.9189
R7830 VX.n10 VX.n9 11.9189
R7831 VX.n32 VX.n22 6.32873
R7832 VX.n22 VX.n17 6.10866
R7833 VX.n31 VX.n26 6.03417
R7834 VX.n13 VX.n8 6.03417
R7835 VX.n31 VX.n30 5.88519
R7836 VX.n13 VX.n12 5.88519
R7837 VX.n32 VX.n31 5.88439
R7838 VX.n33 VX.n13 5.88428
R7839 VX.n22 VX.n21 5.8107
R7840 VX.n59 VX.n58 5.66239
R7841 VX.n61 VX.n60 5.59128
R7842 VX.n34 VX.n33 5.43287
R7843 VX.n2 VX.n0 4.61117
R7844 VX.n62 VX.t17 4.61117
R7845 VX.n34 VX.n4 4.2863
R7846 VX.n2 VX.n1 3.20717
R7847 VX.n62 VX.t16 3.20717
R7848 VX.n39 VX.n37 3.1505
R7849 VX.n52 VX.n50 3.1505
R7850 VX.n41 VX.n40 2.60725
R7851 VX.n59 VX.n56 2.50615
R7852 VX.n60 VX.n34 2.2505
R7853 VX.n46 VX.n44 1.78546
R7854 VX.n41 VX.n39 1.45274
R7855 VX.n53 VX.n52 1.40137
R7856 VX.n55 VX.n47 1.27585
R7857 VX.n56 VX.n55 1.15061
R7858 VX.n60 VX.n59 1.13035
R7859 VX.n55 VX.n54 1.12656
R7860 VX.n56 VX.n42 1.1178
R7861 VX.n61 VX.n2 0.921572
R7862 VX.n52 VX.n51 0.863826
R7863 VX.n39 VX.n38 0.851587
R7864 VX.n36 VX.n35 0.800639
R7865 VX.n46 VX.n45 0.775265
R7866 VX VX.n62 0.7619
R7867 VX.n58 VX.t11 0.5465
R7868 VX.n58 VX.n57 0.5465
R7869 VX.n40 VX.t10 0.5465
R7870 VX.n40 VX.t1 0.5465
R7871 VX.n37 VX.t8 0.5465
R7872 VX.n37 VX.t5 0.5465
R7873 VX.n44 VX.t7 0.5465
R7874 VX.n44 VX.n43 0.5465
R7875 VX.n50 VX.t3 0.5465
R7876 VX.n50 VX.n49 0.5465
R7877 VX.n4 VX.t9 0.5465
R7878 VX.n4 VX.n3 0.5465
R7879 VX.n33 VX.n32 0.4455
R7880 VX.n42 VX.n36 0.405068
R7881 VX VX.n61 0.154524
R7882 VX.n47 VX.n46 0.115871
R7883 VX.n54 VX.n53 0.0721087
R7884 VX.n42 VX.n41 0.0331417
R7885 VX.n54 VX.n48 0.032107
R7886 VA.n27 VA.t10 33.7219
R7887 VA.n22 VA.t12 33.5264
R7888 VA.n5 VA.t14 30.5282
R7889 VA.n1 VA.t8 30.3978
R7890 VA.n13 VA.n12 7.3045
R7891 VA VA.n29 5.2068
R7892 VA.n14 VA.n13 4.87764
R7893 VA.n19 VA.n18 3.60336
R7894 VA.n25 VA.n19 3.4268
R7895 VA.n12 VA.n9 3.26712
R7896 VA.n12 VA.n11 3.25833
R7897 VA.n23 VA.n21 3.16819
R7898 VA.n29 VA.n28 3.16468
R7899 VA.n24 VA.n23 2.80761
R7900 VA.n19 VA.n16 2.6005
R7901 VA.n26 VA.n25 2.34348
R7902 VA.n7 VA.n2 1.92616
R7903 VA.n13 VA.n7 1.72443
R7904 VA.n7 VA.n6 1.22918
R7905 VA.n2 VA.n0 1.19523
R7906 VA.n6 VA.n4 1.19326
R7907 VA.n6 VA.n5 0.683691
R7908 VA.n2 VA.n1 0.660465
R7909 VA.n28 VA.t7 0.607167
R7910 VA.n28 VA.t11 0.607167
R7911 VA.n21 VA.t13 0.607167
R7912 VA.n21 VA.n20 0.607167
R7913 VA.n18 VA.t16 0.607167
R7914 VA.n18 VA.n17 0.607167
R7915 VA.n16 VA.t17 0.607167
R7916 VA.n16 VA.n15 0.607167
R7917 VA.n9 VA.t3 0.607167
R7918 VA.n9 VA.n8 0.607167
R7919 VA.n11 VA.t0 0.607167
R7920 VA.n11 VA.n10 0.607167
R7921 VA.n4 VA.t15 0.607167
R7922 VA.n4 VA.n3 0.607167
R7923 VA.n0 VA.t1 0.607167
R7924 VA.n0 VA.t9 0.607167
R7925 VA VA.n26 0.431462
R7926 VA.n26 VA.n14 0.125115
R7927 VA.n23 VA.n22 0.0534007
R7928 VA.n29 VA.n27 0.0444286
R7929 VA.n25 VA.n24 0.0146322
R7930 VC.n34 VC.t38 56.2889
R7931 VC.n10 VC.t32 55.9277
R7932 VC.n31 VC.t34 55.8956
R7933 VC.n13 VC.t36 55.4158
R7934 VC.n76 VC.t26 55.0018
R7935 VC.n79 VC.t28 54.9998
R7936 VC.n43 VC.t24 54.9964
R7937 VC.n46 VC.t30 54.9896
R7938 VC.n95 VC.t42 47.1352
R7939 VC.n83 VC.t46 47.1036
R7940 VC.n86 VC.t50 44.8434
R7941 VC.n106 VC.t44 44.8434
R7942 VC.n100 VC.t40 44.8434
R7943 VC.n97 VC.t48 44.8434
R7944 VC.n58 VC.t23 5.58454
R7945 VC.n60 VC.t17 5.58454
R7946 VC.n53 VC.n52 5.58454
R7947 VC.n55 VC.n54 5.58454
R7948 VC.n115 VC.n114 4.35225
R7949 VC.n96 VC.n95 4.03836
R7950 VC.n109 VC.n108 4.0005
R7951 VC.n88 VC.n87 4.0005
R7952 VC.n102 VC.n101 4.0005
R7953 VC.n99 VC.n98 4.0005
R7954 VC.n58 VC.n57 3.6965
R7955 VC.n60 VC.n59 3.6965
R7956 VC.n53 VC.t18 3.6965
R7957 VC.n55 VC.t22 3.6965
R7958 VC.n89 VC.n85 3.62641
R7959 VC.n103 VC.n92 3.62641
R7960 VC.n96 VC.n94 3.62641
R7961 VC.n71 VC.n68 3.4441
R7962 VC.n62 VC.n56 3.09912
R7963 VC.n5 VC.n4 3.0681
R7964 VC.n2 VC.n1 3.06142
R7965 VC.n63 VC.n62 3.03192
R7966 VC.n48 VC.n47 2.62105
R7967 VC.n45 VC.n40 2.62099
R7968 VC.n44 VC.n42 2.62076
R7969 VC.n81 VC.n80 2.61951
R7970 VC.n78 VC.n73 2.61951
R7971 VC.n77 VC.n75 2.61862
R7972 VC.n71 VC.n70 2.61099
R7973 VC.n66 VC.n65 2.61045
R7974 VC.n63 VC.n51 2.6061
R7975 VC.n24 VC.n23 2.52173
R7976 VC.n19 VC.n18 2.52114
R7977 VC.n36 VC.n35 2.44199
R7978 VC.n33 VC.n28 2.44109
R7979 VC.n32 VC.n30 2.44021
R7980 VC.n11 VC.n9 2.43525
R7981 VC.n15 VC.n14 2.43469
R7982 VC.n12 VC.n7 2.43462
R7983 VC.n101 VC.n100 2.37724
R7984 VC.n98 VC.n97 2.29236
R7985 VC.n116 VC.n71 2.25886
R7986 VC.n117 VC.n66 2.25826
R7987 VC.n26 VC.n2 2.25371
R7988 VC.n21 VC.n5 2.25371
R7989 VC.n62 VC.n61 2.2505
R7990 VC.n20 VC.n19 2.2505
R7991 VC.n25 VC.n24 2.2505
R7992 VC.n115 VC.n82 2.2505
R7993 VC.n118 VC.n49 2.2505
R7994 VC.n87 VC.n86 2.20748
R7995 VC.n108 VC.n105 2.03771
R7996 VC.n107 VC.n106 2.03771
R7997 VC.n20 VC.n16 1.47548
R7998 VC.n90 VC.n83 1.33644
R7999 VC.n11 VC.n10 1.33543
R8000 VC.n32 VC.n31 1.332
R8001 VC.n15 VC.n13 1.32509
R8002 VC.n36 VC.n34 1.32446
R8003 VC.n48 VC.n46 1.31314
R8004 VC.n44 VC.n43 1.31277
R8005 VC.n81 VC.n79 1.31213
R8006 VC.n77 VC.n76 1.30769
R8007 VC.n113 VC.n90 1.16492
R8008 VC.n113 VC.n112 1.14768
R8009 VC.n38 VC.n37 1.09748
R8010 VC.n61 VC.n58 1.06058
R8011 VC.n56 VC.n53 1.06058
R8012 VC.n12 VC.n11 0.89438
R8013 VC.n33 VC.n32 0.893512
R8014 VC.n78 VC.n77 0.847423
R8015 VC.n45 VC.n44 0.844344
R8016 VC.n66 VC.n63 0.836178
R8017 VC.n38 VC.n26 0.809115
R8018 VC.n61 VC.n60 0.768847
R8019 VC.n56 VC.n55 0.768847
R8020 VC.n118 VC.n117 0.6713
R8021 VC.n35 VC.t66 0.607167
R8022 VC.n35 VC.t39 0.607167
R8023 VC.n28 VC.t62 0.607167
R8024 VC.n28 VC.n27 0.607167
R8025 VC.n30 VC.t35 0.607167
R8026 VC.n30 VC.n29 0.607167
R8027 VC.n14 VC.t67 0.607167
R8028 VC.n14 VC.t37 0.607167
R8029 VC.n7 VC.t63 0.607167
R8030 VC.n7 VC.n6 0.607167
R8031 VC.n9 VC.t33 0.607167
R8032 VC.n9 VC.n8 0.607167
R8033 VC.n23 VC.t65 0.607167
R8034 VC.n23 VC.n22 0.607167
R8035 VC.n1 VC.t61 0.607167
R8036 VC.n1 VC.n0 0.607167
R8037 VC.n18 VC.t60 0.607167
R8038 VC.n18 VC.n17 0.607167
R8039 VC.n4 VC.t56 0.607167
R8040 VC.n4 VC.n3 0.607167
R8041 VC.n25 VC.n21 0.595192
R8042 VC.n37 VC.n36 0.587054
R8043 VC.n16 VC.n15 0.583766
R8044 VC.n70 VC.t1 0.5465
R8045 VC.n70 VC.n69 0.5465
R8046 VC.n68 VC.t6 0.5465
R8047 VC.n68 VC.n67 0.5465
R8048 VC.n65 VC.t15 0.5465
R8049 VC.n65 VC.n64 0.5465
R8050 VC.n51 VC.t5 0.5465
R8051 VC.n51 VC.n50 0.5465
R8052 VC.n47 VC.t14 0.5465
R8053 VC.n47 VC.t31 0.5465
R8054 VC.n40 VC.t11 0.5465
R8055 VC.n40 VC.n39 0.5465
R8056 VC.n42 VC.t25 0.5465
R8057 VC.n42 VC.n41 0.5465
R8058 VC.n80 VC.t12 0.5465
R8059 VC.n80 VC.t29 0.5465
R8060 VC.n73 VC.t3 0.5465
R8061 VC.n73 VC.n72 0.5465
R8062 VC.n75 VC.t27 0.5465
R8063 VC.n75 VC.n74 0.5465
R8064 VC.n85 VC.t51 0.5465
R8065 VC.n85 VC.n84 0.5465
R8066 VC.n92 VC.t41 0.5465
R8067 VC.n92 VC.n91 0.5465
R8068 VC.n94 VC.t43 0.5465
R8069 VC.n94 VC.n93 0.5465
R8070 VC.n117 VC.n116 0.4811
R8071 VC VC.n38 0.466021
R8072 VC.n82 VC.n78 0.389361
R8073 VC VC.n118 0.3845
R8074 VC.n82 VC.n81 0.383642
R8075 VC.n49 VC.n45 0.376674
R8076 VC.n49 VC.n48 0.368178
R8077 VC.n116 VC.n115 0.2891
R8078 VC.n16 VC.n12 0.235408
R8079 VC.n37 VC.n33 0.226622
R8080 VC.n108 VC.n107 0.170267
R8081 VC.n102 VC.n99 0.154071
R8082 VC.n112 VC.n111 0.0943913
R8083 VC.n89 VC.n88 0.0390714
R8084 VC.n99 VC.n96 0.0383571
R8085 VC.n103 VC.n102 0.0383571
R8086 VC.n104 VC.n103 0.0212143
R8087 VC.n90 VC.n89 0.0184638
R8088 VC.n109 VC.n104 0.0176429
R8089 VC.n112 VC.n110 0.0109665
R8090 VC.n114 VC.n113 0.0078125
R8091 VC.n110 VC.n109 0.00192857
R8092 VC.n21 VC.n20 0.00119231
R8093 VC.n26 VC.n25 0.00119231
R8094 VD.n24 VD.t59 56.2443
R8095 VD.n7 VD.t51 55.924
R8096 VD.n15 VD.t55 55.5592
R8097 VD.n2 VD.t53 55.5578
R8098 VD.n73 VD.t49 55.0033
R8099 VD.n62 VD.t63 54.9998
R8100 VD.n71 VD.t61 54.9984
R8101 VD.n60 VD.t57 54.9949
R8102 VD.n92 VD.t37 47.1352
R8103 VD.n85 VD.t41 47.1036
R8104 VD.n94 VD.t45 44.8434
R8105 VD.n97 VD.t43 44.8434
R8106 VD.n103 VD.t39 44.8434
R8107 VD.n111 VD.t47 44.8434
R8108 VD.n46 VD.t19 5.39224
R8109 VD.n42 VD.n41 5.38071
R8110 VD.n43 VD.n42 5.11785
R8111 VD.n47 VD.n46 5.06689
R8112 VD.n42 VD.t20 4.77202
R8113 VD.n48 VD.t22 4.77006
R8114 VD.n46 VD.n45 4.76049
R8115 VD.n44 VD.n39 4.44941
R8116 VD.n120 VD.n119 4.09427
R8117 VD.n93 VD.n92 4.03836
R8118 VD.n113 VD.n112 4.0005
R8119 VD.n106 VD.n105 4.0005
R8120 VD.n96 VD.n95 4.0005
R8121 VD.n99 VD.n98 4.0005
R8122 VD.n93 VD.n91 3.62641
R8123 VD.n100 VD.n89 3.62641
R8124 VD.n114 VD.n87 3.62641
R8125 VD.n84 VD.n81 3.44138
R8126 VD.n50 VD.n49 3.28338
R8127 VD.n14 VD.n13 3.12963
R8128 VD.n37 VD.n36 3.12513
R8129 VD.n56 VD.n52 3.07277
R8130 VD.n49 VD.n44 2.6551
R8131 VD.n61 VD.n59 2.61997
R8132 VD.n67 VD.n66 2.61988
R8133 VD.n78 VD.n77 2.61927
R8134 VD.n72 VD.n70 2.61922
R8135 VD.n75 VD.n74 2.61864
R8136 VD.n64 VD.n63 2.61837
R8137 VD.n84 VD.n83 2.61079
R8138 VD.n14 VD.n11 2.57348
R8139 VD.n37 VD.n34 2.5726
R8140 VD.n3 VD.n1 2.43744
R8141 VD.n20 VD.n19 2.43742
R8142 VD.n29 VD.n28 2.43722
R8143 VD.n17 VD.n16 2.43707
R8144 VD.n26 VD.n25 2.43662
R8145 VD.n8 VD.n6 2.43646
R8146 VD.n98 VD.n97 2.37724
R8147 VD.n95 VD.n94 2.29236
R8148 VD.n32 VD.n4 2.27729
R8149 VD.n23 VD.n9 2.27621
R8150 VD.n120 VD.n84 2.25741
R8151 VD.n22 VD.n21 2.2505
R8152 VD.n31 VD.n30 2.2505
R8153 VD.n49 VD.n48 2.2505
R8154 VD.n123 VD.n57 2.2505
R8155 VD.n122 VD.n68 2.2505
R8156 VD.n121 VD.n79 2.2505
R8157 VD.n56 VD.n55 2.24525
R8158 VD.n112 VD.n111 2.20748
R8159 VD.n105 VD.n102 2.03771
R8160 VD.n104 VD.n103 2.03771
R8161 VD.n22 VD.n14 1.90471
R8162 VD.n43 VD.n40 1.89811
R8163 VD.n47 VD.t18 1.88742
R8164 VD.n55 VD.n54 1.48765
R8165 VD.n115 VD.n85 1.33719
R8166 VD.n8 VD.n7 1.33324
R8167 VD.n26 VD.n24 1.32423
R8168 VD.n17 VD.n15 1.32296
R8169 VD.n3 VD.n2 1.32289
R8170 VD.n61 VD.n60 1.31297
R8171 VD.n72 VD.n71 1.31199
R8172 VD.n75 VD.n73 1.31004
R8173 VD.n64 VD.n62 1.30945
R8174 VD.n116 VD.n115 1.20065
R8175 VD.n44 VD.n43 1.16362
R8176 VD.n38 VD.n37 1.09748
R8177 VD.n20 VD.n17 0.902773
R8178 VD.n29 VD.n26 0.899324
R8179 VD.n48 VD.n47 0.881391
R8180 VD.n78 VD.n75 0.850388
R8181 VD.n67 VD.n64 0.850347
R8182 VD VD.n38 0.76296
R8183 VD VD.n123 0.755218
R8184 VD.n121 VD.n120 0.731668
R8185 VD.n36 VD.t35 0.607167
R8186 VD.n36 VD.n35 0.607167
R8187 VD.n34 VD.t67 0.607167
R8188 VD.n34 VD.n33 0.607167
R8189 VD.n13 VD.t36 0.607167
R8190 VD.n13 VD.n12 0.607167
R8191 VD.n11 VD.t27 0.607167
R8192 VD.n11 VD.n10 0.607167
R8193 VD.n19 VD.t34 0.607167
R8194 VD.n19 VD.n18 0.607167
R8195 VD.n16 VD.t31 0.607167
R8196 VD.n16 VD.t56 0.607167
R8197 VD.n6 VD.t52 0.607167
R8198 VD.n6 VD.n5 0.607167
R8199 VD.n28 VD.t0 0.607167
R8200 VD.n28 VD.n27 0.607167
R8201 VD.n25 VD.t33 0.607167
R8202 VD.n25 VD.t60 0.607167
R8203 VD.n1 VD.t54 0.607167
R8204 VD.n1 VD.n0 0.607167
R8205 VD.n31 VD.n23 0.593808
R8206 VD.n83 VD.t9 0.5465
R8207 VD.n83 VD.n82 0.5465
R8208 VD.n81 VD.t12 0.5465
R8209 VD.n81 VD.n80 0.5465
R8210 VD.n77 VD.t6 0.5465
R8211 VD.n77 VD.n76 0.5465
R8212 VD.n74 VD.t10 0.5465
R8213 VD.n74 VD.t50 0.5465
R8214 VD.n70 VD.t62 0.5465
R8215 VD.n70 VD.n69 0.5465
R8216 VD.n66 VD.t3 0.5465
R8217 VD.n66 VD.n65 0.5465
R8218 VD.n63 VD.t7 0.5465
R8219 VD.n63 VD.t64 0.5465
R8220 VD.n59 VD.t58 0.5465
R8221 VD.n59 VD.n58 0.5465
R8222 VD.n54 VD.t16 0.5465
R8223 VD.n54 VD.n53 0.5465
R8224 VD.n52 VD.t13 0.5465
R8225 VD.n52 VD.n51 0.5465
R8226 VD.n91 VD.t38 0.5465
R8227 VD.n91 VD.n90 0.5465
R8228 VD.n89 VD.t44 0.5465
R8229 VD.n89 VD.n88 0.5465
R8230 VD.n87 VD.t48 0.5465
R8231 VD.n87 VD.n86 0.5465
R8232 VD.n122 VD.n121 0.528018
R8233 VD.n4 VD.n3 0.500303
R8234 VD.n9 VD.n8 0.493909
R8235 VD.n68 VD.n61 0.392883
R8236 VD.n79 VD.n72 0.392063
R8237 VD.n79 VD.n78 0.38736
R8238 VD.n38 VD.n32 0.381269
R8239 VD.n68 VD.n67 0.380664
R8240 VD.n123 VD.n122 0.319113
R8241 VD.n30 VD.n29 0.203821
R8242 VD.n21 VD.n20 0.202321
R8243 VD.n105 VD.n104 0.170267
R8244 VD.n99 VD.n96 0.154071
R8245 VD.n110 VD.n109 0.0790714
R8246 VD.n117 VD.n116 0.062375
R8247 VD.n113 VD.n110 0.0490714
R8248 VD.n114 VD.n113 0.0390714
R8249 VD.n96 VD.n93 0.0383571
R8250 VD.n100 VD.n99 0.0383571
R8251 VD.n101 VD.n100 0.0212143
R8252 VD.n115 VD.n114 0.0187151
R8253 VD.n106 VD.n101 0.0176429
R8254 VD.n109 VD.n108 0.0176429
R8255 VD.n118 VD.n117 0.014
R8256 VD.n57 VD.n50 0.0139871
R8257 VD.n57 VD.n56 0.0124995
R8258 VD.n108 VD.n107 0.00621429
R8259 VD.n119 VD.n118 0.005
R8260 VD.n107 VD.n106 0.00192857
R8261 VD.n23 VD.n22 0.00119231
R8262 VD.n32 VD.n31 0.00119231
R8263 VINP.n5 VINP.t14 56.8887
R8264 VINP.n3 VINP.t1 56.8887
R8265 VINP.n2 VINP.t3 56.8887
R8266 VINP.n0 VINP.t10 56.8887
R8267 VINP.n12 VINP.t13 56.8887
R8268 VINP.n10 VINP.t12 56.8887
R8269 VINP.n9 VINP.t0 56.8887
R8270 VINP.n7 VINP.t9 56.8887
R8271 VINP.n0 VINP.t11 56.8325
R8272 VINP.n7 VINP.t8 56.8325
R8273 VINP.n4 VINP.t7 56.7951
R8274 VINP.n1 VINP.t5 56.7951
R8275 VINP.n11 VINP.t6 56.7951
R8276 VINP.n8 VINP.t4 56.7951
R8277 VINP.n13 VINP.t15 55.496
R8278 VINP.n6 VINP.t2 55.495
R8279 VINP.n14 VINP.n13 4.1806
R8280 VINP.n14 VINP.n6 2.99939
R8281 VINP.n16 VINP.n14 1.23127
R8282 VINP.n16 VINP.n15 1.13036
R8283 VINP.n2 VINP.n1 0.223893
R8284 VINP.n4 VINP.n3 0.223893
R8285 VINP.n9 VINP.n8 0.223893
R8286 VINP.n11 VINP.n10 0.223893
R8287 VINP.n1 VINP.n0 0.223455
R8288 VINP.n5 VINP.n4 0.223455
R8289 VINP.n8 VINP.n7 0.223455
R8290 VINP.n12 VINP.n11 0.223455
R8291 VINP.n3 VINP.n2 0.222578
R8292 VINP.n10 VINP.n9 0.222578
R8293 VINP.n6 VINP.n5 0.196877
R8294 VINP.n13 VINP.n12 0.182267
R8295 VINP VINP.n16 0.0468226
R8296 VP.n34 VP.t46 23.9862
R8297 VP.n51 VP.t40 23.9862
R8298 VP.n51 VP.t42 23.9862
R8299 VP.n40 VP.t44 23.9862
R8300 VP.n1 VP.t32 23.9862
R8301 VP.n16 VP.t38 23.9862
R8302 VP.n16 VP.t34 23.9862
R8303 VP.n6 VP.t36 23.9862
R8304 VP.n35 VP.n34 4.0005
R8305 VP.n41 VP.n40 4.0005
R8306 VP.n52 VP.n51 4.0005
R8307 VP.n2 VP.n1 4.0005
R8308 VP.n7 VP.n6 4.0005
R8309 VP.n17 VP.n16 4.0005
R8310 VP.n25 VP.n22 3.87435
R8311 VP.n57 VP.n56 3.53247
R8312 VP.n58 VP.n20 3.34268
R8313 VP.n57 VP.n31 3.34139
R8314 VP.n36 VP.n33 3.19242
R8315 VP.n3 VP.n0 3.19069
R8316 VP.n100 VP.n99 2.82155
R8317 VP.n78 VP.n77 2.81436
R8318 VP.n67 VP.n66 2.80891
R8319 VP.n89 VP.n88 2.80587
R8320 VP.n39 VP.n38 2.6005
R8321 VP.n45 VP.n44 2.6005
R8322 VP.n56 VP.n55 2.6005
R8323 VP.n31 VP.n30 2.6005
R8324 VP.n28 VP.n27 2.6005
R8325 VP.n25 VP.n24 2.6005
R8326 VP.n5 VP.n4 2.6005
R8327 VP.n10 VP.n9 2.6005
R8328 VP.n20 VP.n19 2.6005
R8329 VP.n68 VP.n62 2.40247
R8330 VP.n69 VP.n60 2.40119
R8331 VP.n67 VP.n64 2.40107
R8332 VP.n80 VP.n71 2.40102
R8333 VP.n78 VP.n75 2.40095
R8334 VP.n89 VP.n86 2.40032
R8335 VP.n79 VP.n73 2.40025
R8336 VP.n91 VP.n82 2.39998
R8337 VP.n100 VP.n97 2.39924
R8338 VP.n90 VP.n84 2.39922
R8339 VP.n101 VP.n95 2.39889
R8340 VP.n102 VP.n93 2.39852
R8341 VP.n28 VP.n25 1.27435
R8342 VP.n31 VP.n28 1.27435
R8343 VP.n103 VP.n102 1.1476
R8344 VP.n104 VP.n80 0.775433
R8345 VP.n105 VP.n69 0.772829
R8346 VP.n103 VP.n91 0.772356
R8347 VP.n55 VP.t41 0.607167
R8348 VP.n55 VP.n54 0.607167
R8349 VP.n44 VP.t43 0.607167
R8350 VP.n44 VP.n43 0.607167
R8351 VP.n38 VP.t45 0.607167
R8352 VP.n38 VP.n37 0.607167
R8353 VP.n33 VP.t47 0.607167
R8354 VP.n33 VP.n32 0.607167
R8355 VP.n22 VP.t7 0.607167
R8356 VP.n22 VP.n21 0.607167
R8357 VP.n24 VP.t10 0.607167
R8358 VP.n24 VP.n23 0.607167
R8359 VP.n27 VP.t9 0.607167
R8360 VP.n27 VP.n26 0.607167
R8361 VP.n30 VP.t2 0.607167
R8362 VP.n30 VP.n29 0.607167
R8363 VP.n19 VP.t14 0.607167
R8364 VP.n19 VP.t39 0.607167
R8365 VP.n9 VP.t0 0.607167
R8366 VP.n9 VP.t35 0.607167
R8367 VP.n4 VP.t1 0.607167
R8368 VP.n4 VP.t37 0.607167
R8369 VP.n0 VP.t3 0.607167
R8370 VP.n0 VP.t33 0.607167
R8371 VP.n60 VP.t17 0.607167
R8372 VP.n60 VP.n59 0.607167
R8373 VP.n62 VP.t55 0.607167
R8374 VP.n62 VP.n61 0.607167
R8375 VP.n64 VP.t26 0.607167
R8376 VP.n64 VP.n63 0.607167
R8377 VP.n66 VP.t49 0.607167
R8378 VP.n66 VP.n65 0.607167
R8379 VP.n71 VP.t50 0.607167
R8380 VP.n71 VP.n70 0.607167
R8381 VP.n73 VP.t30 0.607167
R8382 VP.n73 VP.n72 0.607167
R8383 VP.n75 VP.t60 0.607167
R8384 VP.n75 VP.n74 0.607167
R8385 VP.n77 VP.t20 0.607167
R8386 VP.n77 VP.n76 0.607167
R8387 VP.n82 VP.t51 0.607167
R8388 VP.n82 VP.n81 0.607167
R8389 VP.n84 VP.t19 0.607167
R8390 VP.n84 VP.n83 0.607167
R8391 VP.n86 VP.t53 0.607167
R8392 VP.n86 VP.n85 0.607167
R8393 VP.n88 VP.t23 0.607167
R8394 VP.n88 VP.n87 0.607167
R8395 VP.n93 VP.t18 0.607167
R8396 VP.n93 VP.n92 0.607167
R8397 VP.n95 VP.t54 0.607167
R8398 VP.n95 VP.n94 0.607167
R8399 VP.n97 VP.t27 0.607167
R8400 VP.n97 VP.n96 0.607167
R8401 VP.n99 VP.t48 0.607167
R8402 VP.n99 VP.n98 0.607167
R8403 VP.n48 VP.n47 0.590692
R8404 VP.n42 VP.n39 0.590692
R8405 VP.n45 VP.n42 0.590692
R8406 VP.n53 VP.n45 0.590692
R8407 VP.n49 VP.n48 0.590692
R8408 VP.n50 VP.n49 0.590692
R8409 VP.n56 VP.n53 0.590692
R8410 VP.n12 VP.n11 0.590692
R8411 VP.n13 VP.n12 0.590692
R8412 VP.n5 VP.n3 0.590692
R8413 VP.n8 VP.n5 0.590692
R8414 VP.n10 VP.n8 0.590692
R8415 VP.n18 VP.n10 0.590692
R8416 VP.n14 VP.n13 0.590692
R8417 VP.n15 VP.n14 0.590692
R8418 VP.n20 VP.n18 0.590692
R8419 VP.n47 VP.n46 0.588962
R8420 VP.n39 VP.n36 0.588962
R8421 VP.n90 VP.n89 0.420294
R8422 VP.n102 VP.n101 0.415949
R8423 VP.n68 VP.n67 0.414607
R8424 VP.n79 VP.n78 0.41384
R8425 VP.n69 VP.n68 0.412846
R8426 VP.n91 VP.n90 0.41173
R8427 VP.n80 VP.n79 0.410757
R8428 VP.n101 VP.n100 0.408775
R8429 VP.n104 VP.n103 0.383554
R8430 VP.n105 VP.n104 0.380451
R8431 VP.n106 VP.n105 0.374046
R8432 VP.n106 VP.n58 0.221732
R8433 VP.n58 VP.n57 0.192027
R8434 VP.n3 VP.n2 0.183833
R8435 VP.n8 VP.n7 0.183833
R8436 VP.n42 VP.n41 0.182167
R8437 VP.n53 VP.n52 0.182167
R8438 VP.n18 VP.n17 0.182167
R8439 VP.n36 VP.n35 0.1805
R8440 VP.n52 VP.n50 0.178833
R8441 VP.n17 VP.n15 0.178833
R8442 VP VP.n106 0.0105385
R8443 VBIASN2.n5 VBIASN2.n4 20.2258
R8444 VBIASN2.n34 VBIASN2.n33 20.2258
R8445 VBIASN2.n36 VBIASN2.n35 20.2258
R8446 VBIASN2.n3 VBIASN2.n2 20.2258
R8447 VBIASN2.n9 VBIASN2.t22 19.8861
R8448 VBIASN2.n14 VBIASN2.t29 19.8861
R8449 VBIASN2.n81 VBIASN2.t23 19.8861
R8450 VBIASN2.n75 VBIASN2.t39 19.8861
R8451 VBIASN2.n80 VBIASN2.n79 14.8581
R8452 VBIASN2.n13 VBIASN2.n12 14.8581
R8453 VBIASN2.n74 VBIASN2.n73 14.8581
R8454 VBIASN2.n8 VBIASN2.n7 14.8581
R8455 VBIASN2.n83 VBIASN2.n82 11.2888
R8456 VBIASN2.n82 VBIASN2.n81 11.2888
R8457 VBIASN2.n15 VBIASN2.n14 11.2888
R8458 VBIASN2.n16 VBIASN2.n15 11.2888
R8459 VBIASN2.n11 VBIASN2.n10 11.2888
R8460 VBIASN2.n77 VBIASN2.n76 11.2888
R8461 VBIASN2.n76 VBIASN2.n75 11.2888
R8462 VBIASN2.n10 VBIASN2.n9 11.2888
R8463 VBIASN2.n79 VBIASN2.t27 9.7825
R8464 VBIASN2.n73 VBIASN2.t20 9.7825
R8465 VBIASN2.n37 VBIASN2.n36 7.44744
R8466 VBIASN2.n6 VBIASN2.n5 7.39445
R8467 VBIASN2.n6 VBIASN2.n3 7.34145
R8468 VBIASN2.n80 VBIASN2.t35 7.3005
R8469 VBIASN2.t32 VBIASN2.n80 7.3005
R8470 VBIASN2.n81 VBIASN2.t32 7.3005
R8471 VBIASN2.n14 VBIASN2.t37 7.3005
R8472 VBIASN2.t37 VBIASN2.n13 7.3005
R8473 VBIASN2.n15 VBIASN2.t24 7.3005
R8474 VBIASN2.n11 VBIASN2.t7 7.3005
R8475 VBIASN2.n16 VBIASN2.t13 7.3005
R8476 VBIASN2.n34 VBIASN2.t15 7.3005
R8477 VBIASN2.n33 VBIASN2.t21 7.3005
R8478 VBIASN2.n82 VBIASN2.t40 7.3005
R8479 VBIASN2.n83 VBIASN2.t17 7.3005
R8480 VBIASN2.n76 VBIASN2.t25 7.3005
R8481 VBIASN2.n74 VBIASN2.t36 7.3005
R8482 VBIASN2.t34 VBIASN2.n74 7.3005
R8483 VBIASN2.n75 VBIASN2.t34 7.3005
R8484 VBIASN2.n9 VBIASN2.t38 7.3005
R8485 VBIASN2.t38 VBIASN2.n8 7.3005
R8486 VBIASN2.n10 VBIASN2.t31 7.3005
R8487 VBIASN2.n35 VBIASN2.t28 7.3005
R8488 VBIASN2.n36 VBIASN2.t9 7.3005
R8489 VBIASN2.n77 VBIASN2.t11 7.3005
R8490 VBIASN2.n37 VBIASN2.n34 7.28845
R8491 VBIASN2.n17 VBIASN2.n16 4.62994
R8492 VBIASN2.n17 VBIASN2.n11 4.36021
R8493 VBIASN2 VBIASN2.n78 4.06727
R8494 VBIASN2.n85 VBIASN2.n84 4.06631
R8495 VBIASN2.n84 VBIASN2.n83 2.86592
R8496 VBIASN2.n78 VBIASN2.n77 2.7977
R8497 VBIASN2.n32 VBIASN2.n31 2.61477
R8498 VBIASN2.n24 VBIASN2.n23 2.60633
R8499 VBIASN2.n41 VBIASN2.n1 1.84256
R8500 VBIASN2.n18 VBIASN2.n17 1.466
R8501 VBIASN2.n64 VBIASN2.n63 1.23809
R8502 VBIASN2.n71 VBIASN2.n70 1.19902
R8503 VBIASN2.n66 VBIASN2.n65 1.19015
R8504 VBIASN2.n65 VBIASN2.n64 1.15853
R8505 VBIASN2.n61 VBIASN2.n60 1.1255
R8506 VBIASN2.n46 VBIASN2.n43 0.993901
R8507 VBIASN2.n51 VBIASN2.n48 0.97786
R8508 VBIASN2.n25 VBIASN2.n6 0.915407
R8509 VBIASN2.n38 VBIASN2.n37 0.915407
R8510 VBIASN2.n55 VBIASN2.n51 0.915349
R8511 VBIASN2.n43 VBIASN2.t2 0.9105
R8512 VBIASN2.n43 VBIASN2.n42 0.9105
R8513 VBIASN2.n63 VBIASN2.t1 0.9105
R8514 VBIASN2.n63 VBIASN2.n62 0.9105
R8515 VBIASN2.n48 VBIASN2.t5 0.9105
R8516 VBIASN2.n48 VBIASN2.n47 0.9105
R8517 VBIASN2.n53 VBIASN2.t4 0.9105
R8518 VBIASN2.n53 VBIASN2.n52 0.9105
R8519 VBIASN2.n55 VBIASN2.n54 0.868849
R8520 VBIASN2.n1 VBIASN2.t12 0.8195
R8521 VBIASN2.n1 VBIASN2.n0 0.8195
R8522 VBIASN2.n23 VBIASN2.t8 0.8195
R8523 VBIASN2.n23 VBIASN2.n22 0.8195
R8524 VBIASN2.n31 VBIASN2.t10 0.8195
R8525 VBIASN2.n31 VBIASN2.n30 0.8195
R8526 VBIASN2.n54 VBIASN2.n53 0.812856
R8527 VBIASN2.n58 VBIASN2.n46 0.640451
R8528 VBIASN2.n57 VBIASN2.n56 0.54098
R8529 VBIASN2.n68 VBIASN2.n67 0.299021
R8530 VBIASN2.n70 VBIASN2.n69 0.255923
R8531 VBIASN2.n26 VBIASN2.n25 0.241301
R8532 VBIASN2.n85 VBIASN2.n72 0.211633
R8533 VBIASN2.n61 VBIASN2.n58 0.210289
R8534 VBIASN2.n25 VBIASN2.n24 0.170557
R8535 VBIASN2.n39 VBIASN2.n38 0.163625
R8536 VBIASN2.n40 VBIASN2.n39 0.123337
R8537 VBIASN2.n38 VBIASN2.n32 0.113727
R8538 VBIASN2.n71 VBIASN2.n41 0.0894192
R8539 VBIASN2.n29 VBIASN2.n28 0.0860505
R8540 VBIASN2.n65 VBIASN2.n61 0.0740211
R8541 VBIASN2.n67 VBIASN2.n66 0.0740211
R8542 VBIASN2.n69 VBIASN2.n68 0.0740211
R8543 VBIASN2.n27 VBIASN2.n26 0.0692314
R8544 VBIASN2.n21 VBIASN2.n20 0.0599134
R8545 VBIASN2.n45 VBIASN2.n44 0.0586492
R8546 VBIASN2.n51 VBIASN2.n50 0.0584622
R8547 VBIASN2.n50 VBIASN2.n49 0.0572429
R8548 VBIASN2.n60 VBIASN2.n59 0.0513104
R8549 VBIASN2.n20 VBIASN2.n19 0.0497072
R8550 VBIASN2.n19 VBIASN2.n18 0.0418468
R8551 VBIASN2.n46 VBIASN2.n45 0.040877
R8552 VBIASN2.n24 VBIASN2.n21 0.0347237
R8553 VBIASN2.n72 VBIASN2.n71 0.0248899
R8554 VBIASN2.n28 VBIASN2.n27 0.0233115
R8555 VBIASN2.n41 VBIASN2.n40 0.0209255
R8556 VBIASN2.n32 VBIASN2.n29 0.0202472
R8557 VBIASN2.n58 VBIASN2.n57 0.0143462
R8558 VBIASN2.n56 VBIASN2.n55 0.00631525
R8559 VBIASN2.n85 VBIASN2 0.00146774
R8560 VINN.n0 VINN.t10 54.2657
R8561 VINN.n10 VINN.t9 54.2657
R8562 VINN.n4 VINN.t13 53.6747
R8563 VINN.n4 VINN.t5 53.6747
R8564 VINN.n5 VINN.t14 53.6747
R8565 VINN.n5 VINN.t8 53.6747
R8566 VINN.n3 VINN.t1 53.6282
R8567 VINN.n3 VINN.t15 53.6282
R8568 VINN.n6 VINN.t4 53.6282
R8569 VINN.n6 VINN.t0 53.6282
R8570 VINN.n0 VINN.t7 53.5872
R8571 VINN.n1 VINN.t12 53.5872
R8572 VINN.n11 VINN.t11 53.5872
R8573 VINN.n10 VINN.t6 53.5872
R8574 VINN.n2 VINN.t3 52.426
R8575 VINN.n12 VINN.t2 52.3838
R8576 VINN.n13 VINN.n9 4.69366
R8577 VINN.n7 VINN.n6 4.25764
R8578 VINN.n13 VINN.n12 4.17098
R8579 VINN.n7 VINN.n5 4.0005
R8580 VINN.n8 VINN.n4 4.0005
R8581 VINN.n9 VINN.n3 4.0005
R8582 VINN.n14 VINN.n2 2.99912
R8583 VINN VINN.n14 1.56656
R8584 VINN VINN.n15 1.19503
R8585 VINN.n14 VINN.n13 1.16283
R8586 VINN.n8 VINN.n7 0.768714
R8587 VINN.n12 VINN.n11 0.72402
R8588 VINN.n2 VINN.n1 0.713688
R8589 VINN.n1 VINN.n0 0.257643
R8590 VINN.n11 VINN.n10 0.257643
R8591 VINN.n9 VINN.n8 0.257643
R8592 c_mid.n6 c_mid.t3 7.12295
R8593 c_mid.n35 c_mid.t2 5.14938
R8594 c_mid.n30 c_mid.t0 4.4346
R8595 c_mid.n5 c_mid.t1 3.01175
R8596 c_mid.n0 c_mid.t4 2.37396
R8597 c_mid c_mid.n38 2.26149
R8598 c_mid.n2 c_mid.n1 2.2505
R8599 c_mid.n3 c_mid.n2 2.2505
R8600 c_mid.n14 c_mid.n13 2.2505
R8601 c_mid.n20 c_mid.n19 2.2505
R8602 c_mid.n26 c_mid.n25 2.2505
R8603 c_mid.n37 c_mid.n36 2.2505
R8604 c_mid.n0 c_mid.t5 2.2505
R8605 c_mid.n4 c_mid.n3 2.2505
R8606 c_mid.n15 c_mid.n14 2.2505
R8607 c_mid.n16 c_mid.n15 2.2505
R8608 c_mid.n22 c_mid.n21 2.2505
R8609 c_mid.n21 c_mid.n20 2.2505
R8610 c_mid.n27 c_mid.n26 2.2505
R8611 c_mid.n28 c_mid.n27 2.2505
R8612 c_mid.n38 c_mid.n37 2.2505
R8613 c_mid.n7 c_mid.n5 2.10922
R8614 c_mid.n13 c_mid.n12 1.1255
R8615 c_mid.n36 c_mid.n35 1.12478
R8616 c_mid.n4 c_mid.n0 0.862121
R8617 c_mid.n7 c_mid.n6 0.101266
R8618 c_mid.n11 c_mid.n10 0.0684091
R8619 c_mid.n34 c_mid.n33 0.0684091
R8620 c_mid.n31 c_mid.n30 0.0413161
R8621 c_mid.n12 c_mid.n11 0.0405909
R8622 c_mid.n9 c_mid.n8 0.0266818
R8623 c_mid.n19 c_mid.n18 0.0266818
R8624 c_mid.n35 c_mid.n34 0.0263556
R8625 c_mid.n33 c_mid.n32 0.0242273
R8626 c_mid.n25 c_mid.n24 0.0242273
R8627 c_mid.n36 c_mid.n29 0.0234091
R8628 c_mid.n16 c_mid.n4 0.0210128
R8629 c_mid.n22 c_mid.n16 0.0210128
R8630 c_mid.n28 c_mid.n22 0.0210128
R8631 c_mid.n12 c_mid.n7 0.0160874
R8632 c_mid c_mid.n28 0.0100238
R8633 c_mid.n32 c_mid.n31 0.0095
R8634 c_mid.n25 c_mid.n23 0.0095
R8635 c_mid.n10 c_mid.n9 0.00704545
R8636 c_mid.n19 c_mid.n17 0.00704545
R8637 VBIASN.n22 VBIASN.t4 33.7891
R8638 VBIASN.n0 VBIASN.t6 27.1669
R8639 VBIASN.n23 VBIASN.t2 15.9041
R8640 VBIASN.n0 VBIASN.t7 15.9041
R8641 VBIASN.n1 VBIASN.n0 9.49741
R8642 VBIASN.n13 VBIASN.n12 5.04476
R8643 VBIASN.n29 VBIASN.n20 4.39933
R8644 VBIASN.n25 VBIASN.n24 4.0005
R8645 VBIASN.n5 VBIASN.n4 2.54282
R8646 VBIASN.n10 VBIASN.n9 2.42521
R8647 VBIASN.n18 VBIASN.n17 2.24796
R8648 VBIASN.n11 VBIASN.n5 1.51386
R8649 VBIASN.n11 VBIASN.n10 1.49826
R8650 VBIASN.n2 VBIASN.n1 1.43944
R8651 VBIASN.n24 VBIASN.n23 1.14764
R8652 VBIASN.n7 VBIASN.n6 0.893
R8653 VBIASN.n14 VBIASN.n13 0.834626
R8654 VBIASN.n13 VBIASN.n11 0.754852
R8655 VBIASN.n24 VBIASN.n21 0.209071
R8656 VBIASN.n23 VBIASN.n22 0.156929
R8657 VBIASN.n29 VBIASN.n28 0.0433939
R8658 VBIASN.n5 VBIASN.n3 0.0408598
R8659 VBIASN.n28 VBIASN.n27 0.0205
R8660 VBIASN.n19 VBIASN.n18 0.0193182
R8661 VBIASN VBIASN.n19 0.0111364
R8662 VBIASN.n9 VBIASN.n8 0.0104275
R8663 VBIASN.n9 VBIASN.n7 0.00904126
R8664 VBIASN.n16 VBIASN.n15 0.0086203
R8665 VBIASN.n17 VBIASN.n16 0.00708199
R8666 VBIASN.n17 VBIASN.n14 0.00708199
R8667 VBIASN.n18 VBIASN.n2 0.00622727
R8668 VBIASN.n27 VBIASN.n26 0.0055
R8669 VBIASN.n26 VBIASN.n25 0.00383333
R8670 VBIASN VBIASN.n29 0.00213636
R8671 VB.n12 VB.t10 34.0237
R8672 VB.n5 VB.t14 34.0237
R8673 VB.n12 VB.t8 33.763
R8674 VB.n5 VB.t12 33.763
R8675 VB.n27 VB.n26 6.43271
R8676 VB VB.n19 5.70007
R8677 VB.n23 VB.n22 4.61117
R8678 VB.n20 VB.t16 4.61117
R8679 VB.n14 VB.n12 4.0005
R8680 VB.n6 VB.n5 4.0005
R8681 VB.n19 VB.n1 3.93939
R8682 VB.n18 VB.n17 3.79764
R8683 VB.n15 VB.n11 3.56311
R8684 VB.n7 VB.n3 3.56311
R8685 VB.n18 VB.n10 3.36643
R8686 VB.n23 VB.n21 3.20717
R8687 VB.n20 VB.t18 3.20717
R8688 VB.n19 VB.n18 2.7315
R8689 VB.n27 VB.n24 2.55712
R8690 VB VB.n27 1.84653
R8691 VB.n24 VB.n20 1.53452
R8692 VB.n17 VB.n16 1.17148
R8693 VB.n10 VB.n9 1.17069
R8694 VB.n10 VB.n7 1.02459
R8695 VB.n17 VB.n15 1.02286
R8696 VB.n24 VB.n23 0.997286
R8697 VB.n26 VB.t2 0.607167
R8698 VB.n26 VB.n25 0.607167
R8699 VB.n16 VB.t0 0.607167
R8700 VB.n16 VB.t11 0.607167
R8701 VB.n11 VB.t7 0.607167
R8702 VB.n11 VB.t9 0.607167
R8703 VB.n9 VB.t15 0.607167
R8704 VB.n9 VB.n8 0.607167
R8705 VB.n3 VB.t13 0.607167
R8706 VB.n3 VB.n2 0.607167
R8707 VB.n1 VB.t4 0.607167
R8708 VB.n1 VB.n0 0.607167
R8709 VB.n7 VB.n6 0.198147
R8710 VB.n14 VB.n13 0.194618
R8711 VB.n15 VB.n14 0.187559
R8712 VB.n6 VB.n4 0.184029
R8713 IBIAS2.n18 IBIAS2.n17 21.2802
R8714 IBIAS2.n4 IBIAS2.t5 20.3847
R8715 IBIAS2.n6 IBIAS2.t10 20.3847
R8716 IBIAS2.n24 IBIAS2.t14 20.3482
R8717 IBIAS2.n28 IBIAS2.t9 20.3482
R8718 IBIAS2.n17 IBIAS2.n16 15.9126
R8719 IBIAS2.n7 IBIAS2.n6 13.7257
R8720 IBIAS2.n25 IBIAS2.n24 13.7257
R8721 IBIAS2.n29 IBIAS2.n28 12.1514
R8722 IBIAS2.n5 IBIAS2.n4 12.1514
R8723 IBIAS2.t14 IBIAS2.n23 9.746
R8724 IBIAS2.n28 IBIAS2.t12 7.3005
R8725 IBIAS2.n4 IBIAS2.t8 7.3005
R8726 IBIAS2.n6 IBIAS2.t7 7.3005
R8727 IBIAS2.n24 IBIAS2.t11 7.3005
R8728 IBIAS2.t11 IBIAS2.n22 7.3005
R8729 IBIAS2.n27 IBIAS2.t3 7.3005
R8730 IBIAS2.n3 IBIAS2.t1 7.3005
R8731 IBIAS2.n2 IBIAS2.n1 4.68528
R8732 IBIAS2.n20 IBIAS2.n19 4.13787
R8733 IBIAS2.n8 IBIAS2.n5 4.13405
R8734 IBIAS2 IBIAS2.n29 4.07405
R8735 IBIAS2.n8 IBIAS2.n7 4.0005
R8736 IBIAS2.n26 IBIAS2.n25 4.0005
R8737 IBIAS2.n21 IBIAS2.n0 3.5105
R8738 IBIAS2.n19 IBIAS2.n18 1.77182
R8739 IBIAS2.n14 IBIAS2.n2 1.21038
R8740 IBIAS2.n13 IBIAS2.n12 1.18612
R8741 IBIAS2.n12 IBIAS2.n11 0.9105
R8742 IBIAS2.n26 IBIAS2.n21 0.38117
R8743 IBIAS2.n21 IBIAS2.n20 0.323938
R8744 IBIAS2.n5 IBIAS2.n3 0.222835
R8745 IBIAS2.n29 IBIAS2.n27 0.222835
R8746 IBIAS2.n9 IBIAS2.n8 0.206795
R8747 IBIAS2.n20 IBIAS2.n15 0.125656
R8748 IBIAS2.n10 IBIAS2.n9 0.0952117
R8749 IBIAS2.n15 IBIAS2.n14 0.0862668
R8750 IBIAS2 IBIAS2.n26 0.0605
R8751 IBIAS2.n14 IBIAS2.n13 0.0562224
R8752 IBIAS2.n13 IBIAS2.n10 0.0541071
C0 m3_9877_n5042# m3_10208_n5041# 0.0187f
C1 VP VA 0.00427f
C2 VDD VINN 4.21f
C3 IBIAS VB 1.21f
C4 m3_10209_n7335# OUT 0.0426f
C5 m3_9883_n7335# OUT 0.0417f
C6 VD VBS2 0.0152f
C7 IBIAS3 c_mid 0.00271f
C8 VINP OUT 1.49e-20
C9 VC VX 4.68f
C10 m3_9246_n5046# IBIAS3 9.48e-20
C11 m3_9560_n5045# m3_9877_n5042# 0.019f
C12 m3_9573_n7334# OUT 0.0419f
C13 IBIAS2 VBIASN2 1.26f
C14 m3_9245_n7337# OUT 0.0332f
C15 VP VINN 1.42f
C16 IBIAS VC 8.68e-20
C17 VA VB 4.07f
C18 VDD VINP 2.43f
C19 m3_9246_n5046# m3_9560_n5045# 0.0196f
C20 m3_10527_n5042# OUT 0.0562f
C21 VD VX 3.33f
C22 IBIAS3 OUT 0.00672f
C23 m3_10208_n5041# OUT 0.0424f
C24 m3_9877_n5042# OUT 0.0425f
C25 VB VINN 7.18e-19
C26 IBIAS VD 1.91e-19
C27 VA VC 0.00682f
C28 VP VINP 1.39f
C29 VDD IBIAS3 40.9f
C30 m3_9560_n5045# OUT 0.042f
C31 m3_10524_n10331# OUTo 0.00211f
C32 c_mid OUT 4.11f
C33 VD VBIASN 9.8e-19
C34 m3_9246_n5046# OUT 0.0325f
C35 m3_10209_n10335# OUTo 0.00209f
C36 m3_9883_n10335# OUTo 0.00211f
C37 VA VD 3.72e-19
C38 VDD c_mid 1.69f
C39 VINN VC 0.975f
C40 IBIAS OUTo 0.0368f
C41 m3_9573_n10334# OUTo 0.00211f
C42 VBS2 VX 0.357f
C43 IBIAS3 IBIAS2 0.163f
C44 m3_9245_n10337# OUTo 0.0021f
C45 m3_10527_n8042# OUTo 0.0107f
C46 VC VINP 1.39f
C47 VA OUTo 0.0015f
C48 IBIAS VBS2 0.155f
C49 VDD OUT 3.1f
C50 VB IBIAS3 0.00629f
C51 VINN VD 1.54f
C52 m3_10208_n8041# OUTo 0.0107f
C53 OUT VBS3 0.917f
C54 VBS2 VBIASN 1.09f
C55 OUTo VBIASN2 0.0245f
C56 m3_9877_n8042# OUTo 0.0103f
C57 m3_10209_n10335# m3_10524_n10331# 0.0189f
C58 m3_9560_n8045# OUTo 0.0108f
C59 VP OUT 5.32e-19
C60 VDD VBS3 1.37f
C61 IBIAS VX 4.44e-20
C62 VINP VD 0.924f
C63 VA VBS2 0.392f
C64 m3_9246_n8046# OUTo 0.0119f
C65 m3_9573_n10334# m3_10524_n10331# 7.35e-20
C66 m3_9883_n10335# m3_10209_n10335# 0.0191f
C67 m3_10524_n7331# OUTo 0.0112f
C68 VBS2 VBIASN2 7.02e-21
C69 VDD VP 7.52f
C70 m3_10209_n7335# OUTo 0.011f
C71 m3_9573_n10334# m3_9883_n10335# 0.0199f
C72 m3_9883_n7335# OUTo 0.0112f
C73 VDD IBIAS2 7.02f
C74 VB OUT 1.44f
C75 IBIAS VBIASN 0.5f
C76 VINN VBS2 0.00594f
C77 VA VX 1.4f
C78 m3_9245_n10337# m3_9883_n10335# 1.09e-19
C79 m3_9573_n7334# OUTo 0.0114f
C80 m3_9245_n10337# m3_9573_n10334# 0.0184f
C81 VBS3 IBIAS2 0.00224f
C82 m3_9245_n7337# OUTo 0.012f
C83 VDD VB 7.1f
C84 IBIAS VA 3.14f
C85 m3_10527_n5042# OUTo 0.0156f
C86 IBIAS VBIASN2 9.61e-19
C87 VINP VBS2 4.79e-19
C88 VINN VX 0.0406f
C89 VC OUT 0.634f
C90 IBIAS3 OUTo 16.3f
C91 m3_10208_n5041# OUTo 0.0156f
C92 m3_9877_n5042# OUTo 0.0153f
C93 m3_10208_n8041# m3_10527_n8042# 0.0193f
C94 VP VB 0.00311f
C95 VDD VC 2.64f
C96 IBIAS VINN 0.0199f
C97 m3_9560_n5045# OUTo 0.0155f
C98 m3_9877_n8042# m3_10527_n8042# 1.07e-19
C99 VD OUT 4.89f
C100 IBIAS3 VBS2 3.04e-19
C101 VINP VX 0.00441f
C102 OUTo c_mid 0.168f
C103 VC VBS3 0.735f
C104 m3_9246_n5046# OUTo 0.0168f
C105 m3_9877_n8042# m3_10208_n8041# 0.0187f
C106 VDD VD 2.48f
C107 VA VINN 0.00975f
C108 VP VC 6.6f
C109 IBIAS VINP 0.00116f
C110 m3_10524_n7331# m3_10527_n8042# 0.00854f
C111 m3_9560_n8045# m3_9877_n8042# 0.019f
C112 OUTo OUT 6.64f
C113 VD VBS3 0.637f
C114 m3_9246_n8046# m3_9560_n8045# 0.0196f
C115 m3_10209_n7335# m3_10208_n8041# 0.0088f
C116 VDD OUTo 56.2f
C117 IBIAS IBIAS3 1.9e-20
C118 VB VC 9.06e-20
C119 VP VD 6.79f
C120 VA VINP 4.07e-19
C121 m3_10524_n10331# c_mid 4.88e-20
C122 m3_9883_n7335# m3_9877_n8042# 0.00829f
C123 OUTo VBS3 0.0125f
C124 IBIAS3 VBIASN 4.45e-19
C125 VBS2 OUT 0.814f
C126 m3_10209_n7335# m3_10524_n7331# 0.0189f
C127 m3_9573_n7334# m3_9560_n8045# 0.00756f
C128 VDD VBS2 4.17f
C129 VINN VINP 1.74f
C130 VA IBIAS3 5.49e-19
C131 VB VD 0.00394f
C132 m3_10524_n10331# OUT 0.0709f
C133 OUTo IBIAS2 0.0417f
C134 VBS2 VBS3 0.611f
C135 OUT VX 3.18f
C136 IBIAS3 VBIASN2 3.06f
C137 m3_9573_n7334# m3_10524_n7331# 7.35e-20
C138 m3_9245_n7337# m3_9246_n8046# 0.00876f
C139 m3_9883_n7335# m3_10209_n7335# 0.0191f
C140 m3_10209_n10335# OUT 0.0641f
C141 m3_9883_n10335# OUT 0.0634f
C142 IBIAS OUT 0.0035f
C143 VC VD 10.2f
C144 VB OUTo 0.172f
C145 VP VBS2 4.99e-19
C146 VDD VX 0.441f
C147 m3_9573_n7334# m3_9883_n7335# 0.0199f
C148 m3_9573_n10334# OUT 0.0637f
C149 VBS2 IBIAS2 0.153f
C150 VX VBS3 0.874f
C151 m3_9245_n7337# m3_9883_n7335# 1.09e-19
C152 m3_9245_n10337# OUT 0.0548f
C153 VDD IBIAS 22.9f
C154 m3_9245_n7337# m3_9573_n7334# 0.0184f
C155 m3_10527_n8042# OUT 0.0564f
C156 VDD VBIASN 0.921f
C157 VA OUT 0.014f
C158 VP VX 0.00165f
C159 VB VBS2 0.488f
C160 IBIAS VBS3 0.501f
C161 m3_10208_n8041# OUT 0.0426f
C162 OUT VBIASN2 0.038f
C163 VBS3 VBIASN 0.272f
C164 m3_9877_n8042# OUT 0.0429f
C165 VDD VA 6.26f
C166 IBIAS VP 4.97f
C167 m3_9560_n8045# OUT 0.0423f
C168 m3_10208_n5041# m3_10527_n5042# 0.0193f
C169 VA VBS3 1.29e-19
C170 VINN OUT 0.00979f
C171 VDD VBIASN2 1.56f
C172 IBIAS IBIAS2 0.00103f
C173 VB VX 1.71f
C174 VC VBS2 0.00166f
C175 m3_9246_n8046# OUT 0.0326f
C176 m3_9877_n5042# m3_10527_n5042# 1.07e-19
C177 m3_10524_n7331# OUT 0.0565f
C178 VBIASN IBIAS2 0.0279f
.ends

