magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2278 -4528 2278 4528
<< nwell >>
rect -278 -2528 278 2528
<< nsubdiff >>
rect -195 2423 195 2445
rect -195 -2423 -173 2423
rect 173 -2423 195 2423
rect -195 -2445 195 -2423
<< nsubdiffcont >>
rect -173 -2423 173 2423
<< metal1 >>
rect -184 2423 184 2434
rect -184 -2423 -173 2423
rect 173 -2423 184 2423
rect -184 -2434 184 -2423
<< end >>
