* NGSPICE file created from AWG_MUX_MAGIC.ext - technology: gf180mcuC

.subckt pmos_3p3_ME7U2H a_28_n313# a_n28_n357# a_n116_n313# w_n202_n443#
X0 a_28_n313# a_n28_n357# a_n116_n313# w_n202_n443# pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
.ends

.subckt pmos_3p3_MA2VAR w_n202_n430# a_28_n300# a_n28_n344# a_n116_n300#
X0 a_28_n300# a_n28_n344# a_n116_n300# w_n202_n430# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt nmos_3p3_876RT2 a_n196_n100# a_n52_n100# a_108_n100# a_52_n144# a_n108_n144#
+ VSUBS
X0 a_n52_n100# a_n108_n144# a_n196_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_108_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_3A6RT2 a_28_n100# a_n28_n144# a_n116_n100# VSUBS
X0 a_28_n100# a_n28_n144# a_n116_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt nmos_3p3_7WQWW2 a_108_n288# a_n196_n288# a_52_n332# a_n52_n288# a_n108_n332#
+ VSUBS
X0 a_108_n288# a_52_n332# a_n52_n288# VSUBS nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1 a_n52_n288# a_n108_n332# a_n196_n288# VSUBS nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
.ends

.subckt pmos_3p3_M22VAR a_52_n344# a_108_n300# a_n108_n344# a_n196_n300# a_n52_n300#
+ w_n282_n430#
X0 a_108_n300# a_52_n344# a_n52_n300# w_n282_n430# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1 a_n52_n300# a_n108_n344# a_n196_n300# w_n282_n430# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt pmos_3p3_MNS6FR w_n282_n505# a_108_n375# a_n196_n375# a_52_n419# a_n108_n419#
+ a_n52_n375#
X0 a_108_n375# a_52_n419# a_n52_n375# w_n282_n505# pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X1 a_n52_n375# a_n108_n419# a_n196_n375# w_n282_n505# pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
.ends

.subckt nmos_3p3_M86RTJ a_28_n300# a_n28_n344# a_n116_n300# VSUBS
X0 a_28_n300# a_n28_n344# a_n116_n300# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt nmos_3p3_276RTJ a_52_n344# a_108_n300# a_n108_n344# a_n196_n300# a_n52_n300#
+ VSUBS
X0 a_108_n300# a_52_n344# a_n52_n300# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1 a_n52_n300# a_n108_n344# a_n196_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt nmos_3p3_2F3WC4 a_n796_n468# a_100_n468# a_n708_24# a_508_n512# a_n508_n468#
+ a_508_24# a_404_68# a_204_n512# a_n204_n468# a_n508_68# a_n100_24# a_n708_n512#
+ a_708_68# a_n796_68# a_n404_n512# a_n100_n512# a_n404_24# a_204_24# a_708_n468#
+ a_100_68# a_404_n468# a_n204_68# VSUBS
X0 a_n204_n468# a_n404_n512# a_n508_n468# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1 a_n508_n468# a_n708_n512# a_n796_n468# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X2 a_100_68# a_n100_24# a_n204_68# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X3 a_404_n468# a_204_n512# a_100_n468# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X4 a_100_n468# a_n100_n512# a_n204_n468# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X5 a_708_n468# a_508_n512# a_404_n468# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X6 a_404_68# a_204_24# a_100_68# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X7 a_n204_68# a_n404_24# a_n508_68# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X8 a_708_68# a_508_24# a_404_68# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X9 a_n508_68# a_n708_24# a_n796_68# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
.ends

.subckt nmos_3p3_NE3WC4 a_100_n200# a_n100_n244# a_n188_n200# VSUBS
X0 a_100_n200# a_n100_n244# a_n188_n200# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=1u
.ends

.subckt ppolyf_u_2VJWHK a_n100_500# a_n100_n602# w_n284_n786#
X0 a_n100_500# a_n100_n602# w_n284_n786# ppolyf_u r_width=1u r_length=5u
.ends

.subckt nmos_3p3_EA6RT2 a_212_n144# a_268_n100# a_n268_n144# a_n356_n100# a_n52_n100#
+ a_n212_n100# a_108_n100# a_52_n144# a_n108_n144# VSUBS
X0 a_n52_n100# a_n108_n144# a_n212_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n212_n100# a_n268_n144# a_n356_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 a_108_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_268_n100# a_212_n144# a_108_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt pmos_3p3_5L6RD7 w_n230_n530# a_56_n400# a_n56_n444# a_n144_n400#
X0 a_56_n400# a_n56_n444# a_n144_n400# w_n230_n530# pfet_03v3 ad=1.76p pd=8.88u as=1.76p ps=8.88u w=4u l=0.56u
.ends

.subckt nmos_3p3_S75EG7 a_212_n144# a_n908_n144# a_268_n100# a_n1068_n144# a_1012_n144#
+ a_1068_n100# a_n1156_n100# a_n692_n100# a_n268_n144# a_372_n144# a_428_n100# a_n52_n100#
+ a_n852_n100# a_n428_n144# a_n1012_n100# a_532_n144# a_588_n100# a_n212_n100# a_n588_n144#
+ a_692_n144# a_748_n100# a_n372_n100# a_n748_n144# a_852_n144# a_108_n100# a_52_n144#
+ a_908_n100# a_n532_n100# a_n108_n144# VSUBS
X0 a_n52_n100# a_n108_n144# a_n212_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_588_n100# a_532_n144# a_428_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n212_n100# a_n268_n144# a_n372_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_n692_n100# a_n748_n144# a_n852_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_1068_n100# a_1012_n144# a_908_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_748_n100# a_692_n144# a_588_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_108_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_268_n100# a_212_n144# a_108_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 a_n372_n100# a_n428_n144# a_n532_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_n852_n100# a_n908_n144# a_n1012_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X10 a_428_n100# a_372_n144# a_268_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X11 a_n1012_n100# a_n1068_n144# a_n1156_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X12 a_908_n100# a_852_n144# a_748_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X13 a_n532_n100# a_n588_n144# a_n692_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_5J7TC4 a_252_n100# a_n252_n144# a_n340_n100# a_n52_n100# a_52_n144#
+ VSUBS
X0 a_n52_n100# a_n252_n144# a_n340_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=1u
X1 a_252_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=1u
.ends

.subckt pmos_3p3_MYZUAR w_n202_n530# a_28_n400# a_n28_n444# a_n116_n400#
X0 a_28_n400# a_n28_n444# a_n116_n400# w_n202_n530# pfet_03v3 ad=1.76p pd=8.88u as=1.76p ps=8.88u w=4u l=0.28u
.ends

.subckt nfet_03v3_DNL5WS a_n196_n100# a_n52_n100# a_108_n100# a_52_n144# a_n108_n144#
+ VSUBS
X0 a_n52_n100# a_n108_n144# a_n196_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_108_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt pfet_03v3_6DZECV a_n196_n100# a_n52_n100# w_n282_n230# a_108_n100# a_52_n144#
+ a_n108_n144#
X0 a_n52_n100# a_n108_n144# a_n196_n100# w_n282_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_108_n100# a_52_n144# a_n52_n100# w_n282_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nfet_03v3_DNQ7WS a_28_n100# a_n28_n144# a_n116_n100# VSUBS
X0 a_28_n100# a_n28_n144# a_n116_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt TGATE_PGA_MAGIC VDD VSS B CLK A
Xnfet_03v3_DNL5WS_0 A B A CLK CLK VSS nfet_03v3_DNL5WS
Xpfet_03v3_6DZECV_0 VDD a_n36_13# VDD VDD CLK CLK pfet_03v3_6DZECV
Xpfet_03v3_6DZECV_1 A B VDD A a_n36_13# a_n36_13# pfet_03v3_6DZECV
Xnfet_03v3_DNQ7WS_0 a_n36_13# CLK VSS VSS nfet_03v3_DNQ7WS
.ends

.subckt ppolyf_u_VRC5QE a_2280_n202# a_4240_100# a_1720_n202# a_2560_100# a_n2200_n202#
+ a_n1640_n202# a_n4160_100# a_3120_n202# a_n2480_100# a_2560_n202# a_n3040_n202#
+ a_880_100# a_n2480_n202# a_n1920_n202# a_n2200_100# a_600_100# a_3680_100# w_n4904_n386#
+ a_3400_n202# a_2840_n202# a_n3320_n202# a_n520_100# a_n2760_n202# a_3400_100# a_1720_100#
+ a_4240_n202# a_3680_n202# a_n4160_n202# a_n3320_100# a_n1640_100# a_n3600_n202#
+ a_40_n202# a_4520_100# a_4520_n202# a_2840_100# a_3960_n202# a_320_n202# a_n4440_n202#
+ a_n3880_n202# a_n4440_100# a_1160_100# a_40_100# a_n2760_100# a_600_n202# a_n1080_100#
+ a_n4720_n202# a_3960_100# a_n800_100# a_880_n202# a_2280_100# a_n240_n202# a_n3880_100#
+ a_2000_100# a_n3600_100# a_n1920_100# a_n520_n202# a_1160_n202# a_320_100# a_n1080_n202#
+ a_n240_100# a_3120_100# a_n4720_100# a_1440_100# a_n800_n202# a_2000_n202# a_1440_n202#
+ a_n1360_n202# a_n3040_100# a_n1360_100#
X0 a_600_100# a_600_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X1 a_2280_100# a_2280_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X2 a_n800_100# a_n800_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X3 a_1160_100# a_1160_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X4 a_n4160_100# a_n4160_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X5 a_n240_100# a_n240_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X6 a_n3600_100# a_n3600_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X7 a_40_100# a_40_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X8 a_n3040_100# a_n3040_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X9 a_4520_100# a_4520_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X10 a_n2480_100# a_n2480_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X11 a_3960_100# a_3960_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X12 a_n1360_100# a_n1360_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X13 a_3400_100# a_3400_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X14 a_2840_100# a_2840_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X15 a_1720_100# a_1720_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X16 a_n4720_100# a_n4720_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X17 a_880_100# a_880_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X18 a_320_100# a_320_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X19 a_n1920_100# a_n1920_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X20 a_4240_100# a_4240_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X21 a_n2200_100# a_n2200_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X22 a_3680_100# a_3680_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X23 a_3120_100# a_3120_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X24 a_n1080_100# a_n1080_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X25 a_2560_100# a_2560_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X26 a_2000_100# a_2000_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X27 a_1440_100# a_1440_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X28 a_n4440_100# a_n4440_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X29 a_n520_100# a_n520_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X30 a_n3880_100# a_n3880_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X31 a_n3320_100# a_n3320_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X32 a_n2760_100# a_n2760_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
X33 a_n1640_100# a_n1640_n202# w_n4904_n386# ppolyf_u r_width=1u r_length=1u
.ends

.subckt pag_res_magic A B G E C H F D VDD
Xppolyf_u_VRC5QE_0 m1_7017_3724# F m1_5335_5023# m1_7297_4056# m1_2973_3724# m1_6642_3724#
+ m1_577_3724# m1_8322_3724# m1_2680_4056# m1_7575_3720# C m1_5335_4371# m1_2973_3724#
+ m1_3095_3720# m1_2973_4056# m1_6642_4376# m1_8882_4056# VDD H D m1_3842_3724# m1_3095_5024#
+ m1_855_5023# m1_8415_4029# m1_6737_4056# m1_8977_3724# F m1_577_3724# m1_1695_4029#
+ m1_3512_4056# G m1_5057_3724# VDD VDD m1_7992_4056# m1_8977_3724# m1_5057_3724#
+ m1_577_3724# G E m1_6175_4029# m1_5242_4056# m1_2680_4056# m1_5802_3724# m1_3935_4029#
+ VDD m1_7575_5024# m1_4402_4056# m1_6082_3724# m1_7297_4056# m1_4497_3724# m1_2162_4376#
+ m1_6737_4056# G m1_2973_4056# m1_4497_3724# m1_8322_3724# m1_5335_4029# m1_6082_3724#
+ m1_5242_4056# m1_7575_4371# VDD m1_6642_4056# m1_5802_3724# m1_7017_3724# m1_6642_3724#
+ m1_3842_3724# m1_2162_4056# m1_3095_4371# ppolyf_u_VRC5QE
Xppolyf_u_VRC5QE_1 m1_7017_5028# m1_8966_5360# m1_5335_4029# m1_7297_5360# m1_2537_5028#
+ m1_3512_4920# E m1_7575_4677# m1_2257_5360# m1_7575_5024# m1_2162_5028# m1_6036_5360#
+ m1_2537_5028# m1_3095_5024# m1_2817_5360# m1_8882_5360# m1_8882_5360# VDD m1_9442_4708#
+ m1_7992_4920# m1_1695_5024# m1_4486_5360# m1_577_3724# m1_8602_5360# m1_6737_5360#
+ D m1_8882_5028# m1_855_5023# G m1_3562_5360# m1_714_4708# m1_5242_5028# VDD VDD
+ m1_8042_5360# m1_7575_3720# m1_5335_5023# E m1_2162_4708# E a_5435_4665# m1_5057_5360#
+ m1_2257_5360# m1_6642_4708# m1_4122_5360# VDD m1_8966_5360# m1_4402_5360# m1_5194_4708#
+ m1_7297_5360# m1_5242_5028# m1_4402_5360# m1_6737_5360# m1_4122_5360# m1_2817_5360#
+ m1_3095_3720# m1_6175_5024# m1_5057_5360# m1_4962_4708# m1_4486_5360# m1_8135_5333#
+ VDD m1_8042_5360# m1_4402_5028# m1_7017_5028# m1_6642_5028# m1_3095_4677# m1_3562_5360#
+ m1_3655_5333# ppolyf_u_VRC5QE
Xppolyf_u_VRC5QE_2 m1_7017_4376# m1_9442_4708# m1_6175_4029# m1_7575_4677# m1_4122_5360#
+ m1_4402_4056# G m1_8137_4376# m1_4122_5360# m1_7575_4371# m1_2162_4376# m1_6082_4708#
+ m1_4122_5360# m1_3095_4371# m1_4122_5360# m1_6642_5028# m1_7992_4920# VDD m1_8137_4376#
+ m1_8882_4056# m1_1417_4376# m1_3655_5333# m1_1695_4029# B m1_6175_5024# B m1_7992_4056#
+ G m1_3842_4708# m1_4402_5028# m1_1417_4376# m1_5242_4376# VDD VDD m1_8882_5028#
+ m1_8415_4029# m1_5335_4371# A m1_2162_4056# m1_714_4708# m1_8322_4708# m1_5194_4708#
+ m1_1695_5024# m1_6642_4056# m1_6082_4708# VDD m1_8135_5333# m1_3512_4920# m1_5897_4376#
+ m1_8602_5360# m1_5242_4376# m1_2162_5028# m1_6036_5360# C m1_3095_4677# m1_3935_4029#
+ m1_5897_4376# a_5435_4665# m1_3657_4376# m1_4962_4708# m1_8322_4708# VDD m1_6642_4708#
+ m1_3512_4056# m1_7017_4376# m1_6642_4376# m1_3657_4376# m1_2162_4708# m1_3842_4708#
+ ppolyf_u_VRC5QE
.ends

.subckt pga_res_magice_parallel VDD C B D H G E F A
Xpag_res_magic_0 A B G E C H F D VDD pag_res_magic
Xpag_res_magic_1 A B G E C H F D VDD pag_res_magic
.ends

.subckt pmos_3p3_MAEVAR a_28_n668# a_n116_n668# a_28_68# a_n28_n712# a_n28_24# w_n202_n798#
+ a_n116_68#
X0 a_28_68# a_n28_24# a_n116_68# w_n202_n798# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X1 a_28_n668# a_n28_n712# a_n116_n668# w_n202_n798# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt pmos_3p3_MES6FR w_n202_n505# a_28_n375# a_n116_n375# a_n28_n419#
X0 a_28_n375# a_n28_n419# a_n116_n375# w_n202_n505# pfet_03v3 ad=1.65p pd=8.38u as=1.65p ps=8.38u w=3.75u l=0.28u
.ends

.subckt pmos_3p3_RKK9DS a_n52_n50# a_n1172_n50# a_428_n50# a_908_n50# a_588_n50# a_1068_n50#
+ a_n428_n94# a_n588_n94# a_n908_n94# a_n1068_n94# a_n212_n50# a_532_n94# a_n372_n50#
+ a_1012_n94# a_n852_n50# a_1172_n94# a_692_n94# a_52_n94# w_n1402_n180# a_108_n50#
+ a_268_n50# a_748_n50# a_1228_n50# a_n1316_n50# a_n108_n94# a_n268_n94# a_n748_n94#
+ a_n1228_n94# a_212_n94# a_372_n94# a_n532_n50# a_n692_n50# a_n1012_n50# a_852_n94#
X0 a_1228_n50# a_1172_n94# a_1068_n50# w_n1402_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 a_108_n50# a_52_n94# a_n52_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 a_268_n50# a_212_n94# a_108_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X3 a_n372_n50# a_n428_n94# a_n532_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 a_n852_n50# a_n908_n94# a_n1012_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 a_428_n50# a_372_n94# a_268_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X6 a_n1012_n50# a_n1068_n94# a_n1172_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X7 a_908_n50# a_852_n94# a_748_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X8 a_n532_n50# a_n588_n94# a_n692_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X9 a_n52_n50# a_n108_n94# a_n212_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X10 a_588_n50# a_532_n94# a_428_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X11 a_n1172_n50# a_n1228_n94# a_n1316_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X12 a_n212_n50# a_n268_n94# a_n372_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X13 a_n692_n50# a_n748_n94# a_n852_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X14 a_1068_n50# a_1012_n94# a_908_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X15 a_748_n50# a_692_n94# a_588_n50# w_n1402_n180# pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
.ends

.subckt cap_mim_2p0fF_3FUNHB m4_n2340_n4500# m4_n2220_n4380#
X0 m4_n2220_n4380# m4_n2340_n4500# cap_mim_2f0_m4m5_noshield c_width=21u c_length=21u
X1 m4_n2220_n4380# m4_n2340_n4500# cap_mim_2f0_m4m5_noshield c_width=21u c_length=21u
.ends

.subckt pmos_3p3_5UYQD7 a_n52_n400# a_164_n400# a_n164_n444# a_n252_n400# a_52_n444#
+ w_n338_n530#
X0 a_n52_n400# a_n164_n444# a_n252_n400# w_n338_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
X1 a_164_n400# a_52_n444# a_n52_n400# w_n338_n530# pfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.56u
.ends

.subckt pmos_3p3_5LZQD7 a_488_n400# a_n488_n444# a_n160_n400# a_376_n444# a_n576_n400#
+ a_272_n400# a_56_n400# a_n56_n444# a_n272_n444# a_160_n444# a_n376_n400# w_n662_n530#
X0 a_56_n400# a_n56_n444# a_n160_n400# w_n662_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1 a_272_n400# a_160_n444# a_56_n400# w_n662_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X2 a_n160_n400# a_n272_n444# a_n376_n400# w_n662_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X3 a_488_n400# a_376_n444# a_272_n400# w_n662_n530# pfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.56u
X4 a_n376_n400# a_n488_n444# a_n576_n400# w_n662_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
.ends

.subckt pmos_3p3_5C3RD7 a_268_n444# a_n52_n400# a_n468_n400# a_380_n400# a_164_n400#
+ a_n164_n444# a_n380_n444# a_52_n444# a_n268_n400# w_n554_n530#
X0 a_n52_n400# a_n164_n444# a_n268_n400# w_n554_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1 a_164_n400# a_52_n444# a_n52_n400# w_n554_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X2 a_380_n400# a_268_n444# a_164_n400# w_n554_n530# pfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.56u
X3 a_n268_n400# a_n380_n444# a_n468_n400# w_n554_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
.ends

.subckt pmos_3p3_HMY8L7 a_812_68# a_n268_68# a_n700_830# a_268_786# a_n484_830# w_n986_n1586#
+ a_164_n1456# a_n596_24# a_n596_n1500# a_n268_n694# a_n484_n694# a_n52_68# a_52_24#
+ a_n484_n1456# a_n700_n694# a_n52_830# a_n164_n738# a_n380_n738# a_380_830# a_n380_786#
+ a_812_n1456# a_484_n1500# a_n268_n1456# a_n900_n1456# a_52_n738# a_380_68# a_484_24#
+ a_n380_n1500# a_52_n1500# a_n484_68# a_n164_24# a_n52_n1456# a_596_n694# a_700_786#
+ a_268_n1500# a_n164_n1500# a_812_n694# a_n812_24# a_484_786# a_596_68# a_n52_n694#
+ a_n268_830# a_52_786# a_n900_830# a_n812_n1500# a_n900_n694# a_812_830# a_596_n1456#
+ a_n700_n1456# a_700_24# a_596_830# a_164_830# a_n812_786# a_n164_786# a_268_n738#
+ a_n596_n738# a_n596_786# a_484_n738# a_700_n1500# a_700_n738# a_n812_n738# a_n700_68#
+ a_268_24# a_164_n694# a_164_68# a_n380_24# a_380_n1456# a_380_n694# a_n900_68#
X0 a_n700_830# a_n812_786# a_n900_830# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.56u
X1 a_n700_68# a_n812_24# a_n900_68# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.56u
X2 a_n700_n1456# a_n812_n1500# a_n900_n1456# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.56u
X3 a_n484_68# a_n596_24# a_n700_68# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X4 a_n268_68# a_n380_24# a_n484_68# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X5 a_n484_n1456# a_n596_n1500# a_n700_n1456# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X6 a_n52_n694# a_n164_n738# a_n268_n694# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X7 a_n52_830# a_n164_786# a_n268_830# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X8 a_380_n1456# a_268_n1500# a_164_n1456# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X9 a_812_830# a_700_786# a_596_830# w_n986_n1586# pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.56u
X10 a_812_n694# a_700_n738# a_596_n694# w_n986_n1586# pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.56u
X11 a_n268_830# a_n380_786# a_n484_830# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X12 a_164_68# a_52_24# a_n52_68# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X13 a_n700_n694# a_n812_n738# a_n900_n694# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.56u
X14 a_n484_830# a_n596_786# a_n700_830# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X15 a_812_68# a_700_24# a_596_68# w_n986_n1586# pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.56u
X16 a_n268_n1456# a_n380_n1500# a_n484_n1456# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X17 a_n52_68# a_n164_24# a_n268_68# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X18 a_812_n1456# a_700_n1500# a_596_n1456# w_n986_n1586# pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.56u
X19 a_380_68# a_268_24# a_164_68# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X20 a_596_68# a_484_24# a_380_68# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X21 a_596_n694# a_484_n738# a_380_n694# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X22 a_380_830# a_268_786# a_164_830# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X23 a_164_n694# a_52_n738# a_n52_n694# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X24 a_380_n694# a_268_n738# a_164_n694# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X25 a_596_n1456# a_484_n1500# a_380_n1456# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X26 a_n484_n694# a_n596_n738# a_n700_n694# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X27 a_n52_n1456# a_n164_n1500# a_n268_n1456# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X28 a_164_n1456# a_52_n1500# a_n52_n1456# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X29 a_164_830# a_52_786# a_n52_830# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X30 a_n268_n694# a_n380_n738# a_n484_n694# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X31 a_596_830# a_484_786# a_380_830# w_n986_n1586# pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
.ends

.subckt pmos_3p3_K823KY a_100_n50# a_n100_n94# a_n188_n50# w_n274_n180#
X0 a_100_n50# a_n100_n94# a_n188_n50# w_n274_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=1u
.ends

.subckt nmos_3p3_U56RT2 a_212_n144# a_268_n100# a_n268_n144# a_372_n144# a_428_n100#
+ a_n52_n100# a_n428_n144# a_n516_n100# a_n212_n100# a_n372_n100# a_108_n100# a_52_n144#
+ a_n108_n144# VSUBS
X0 a_n52_n100# a_n108_n144# a_n212_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n212_n100# a_n268_n144# a_n372_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_108_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_268_n100# a_212_n144# a_108_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_n372_n100# a_n428_n144# a_n516_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X5 a_428_n100# a_372_n144# a_268_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_JE3WC4 a_708_n200# a_404_n200# a_n708_n244# a_n796_n200# a_100_n200#
+ a_n404_n244# a_n100_n244# a_n508_n200# a_n204_n200# a_508_n244# a_204_n244# VSUBS
X0 a_n508_n200# a_n708_n244# a_n796_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X1 a_404_n200# a_204_n244# a_100_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X2 a_100_n200# a_n100_n244# a_n204_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X3 a_708_n200# a_508_n244# a_404_n200# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X4 a_n204_n200# a_n404_n244# a_n508_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
.ends

.subckt ppolyf_u_2V2ZHK a_40_n602# a_40_500# a_n240_n602# w_n424_n786# a_n240_500#
X0 a_40_500# a_40_n602# w_n424_n786# ppolyf_u r_width=1u r_length=5u
X1 a_n240_500# a_n240_n602# w_n424_n786# ppolyf_u r_width=1u r_length=5u
.ends

.subckt nmos_3p3_UUQWW2 a_n28_n332# a_28_n288# a_n116_n288# VSUBS
X0 a_28_n288# a_n28_n332# a_n116_n288# VSUBS nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
.ends

.subckt pmos_3p3_M2NNAR a_n108_n1448# a_52_n712# a_108_n1404# a_n52_n668# a_52_n1448#
+ a_n52_68# a_52_24# a_n108_n712# a_108_804# a_108_68# a_n196_68# a_52_760# a_n196_n1404#
+ a_n108_760# a_108_n668# a_n52_804# a_n52_n1404# a_n196_n668# a_n196_804# a_n108_24#
+ w_n282_n1534#
X0 a_n52_n1404# a_n108_n1448# a_n196_n1404# w_n282_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1 a_108_n668# a_52_n712# a_n52_n668# w_n282_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X2 a_108_804# a_52_760# a_n52_804# w_n282_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X3 a_n52_n668# a_n108_n712# a_n196_n668# w_n282_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X4 a_n52_68# a_n108_24# a_n196_68# w_n282_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X5 a_108_68# a_52_24# a_n52_68# w_n282_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X6 a_n52_804# a_n108_760# a_n196_804# w_n282_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X7 a_108_n1404# a_52_n1448# a_n52_n1404# w_n282_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
.ends

.subckt pmos_3p3_MGRCNG a_n204_n36# a_56_n69# a_112_n25# a_n112_n69# w_n290_n161#
+ a_n56_n25#
X0 a_n56_n25# a_n112_n69# a_n204_n36# w_n290_n161# pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X1 a_112_n25# a_56_n69# a_n56_n25# w_n290_n161# pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
.ends

.subckt nmos_3p3_H9QVWA a_n120_n36# a_28_n25# a_n28_n69# VSUBS
X0 a_28_n25# a_n28_n69# a_n120_n36# VSUBS nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
.ends

.subckt INVERTER_magic IN OUT VDD VSS
Xpmos_3p3_MGRCNG_0 OUT IN OUT IN VDD VDD pmos_3p3_MGRCNG
Xnmos_3p3_H9QVWA_0 VSS OUT IN VSS nmos_3p3_H9QVWA
Xnmos_3p3_H9QVWA_1 VSS VSS VSS VSS nmos_3p3_H9QVWA
.ends

.subckt nmos_3p3_49QVWA a_n204_n36# a_56_n69# a_112_n25# a_n112_n69# a_n56_n25# VSUBS
X0 a_n56_n25# a_n112_n69# a_n204_n36# VSUBS nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X1 a_112_n25# a_56_n69# a_n56_n25# VSUBS nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
.ends

.subckt pmos_3p3_M8RWPS a_n28_n94# w_n202_n180# a_n116_n50# a_28_n50#
X0 a_28_n50# a_n28_n94# a_n116_n50# w_n202_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt AND A B OUT VDD VSS
Xnmos_3p3_H9QVWA_0 VSS OUT a_571_376# VSS nmos_3p3_H9QVWA
Xnmos_3p3_49QVWA_0 m1_41_62# B m1_41_62# B VSS VSS nmos_3p3_49QVWA
Xnmos_3p3_49QVWA_1 m1_41_62# A m1_41_62# A a_571_376# VSS nmos_3p3_49QVWA
Xpmos_3p3_M8RWPS_0 a_571_376# VDD VDD OUT pmos_3p3_M8RWPS
Xpmos_3p3_M8RWPS_1 A VDD VDD a_571_376# pmos_3p3_M8RWPS
Xpmos_3p3_M8RWPS_2 B VDD a_571_376# VDD pmos_3p3_M8RWPS
.ends

.subckt pmos_3p3_M8RCNG a_n120_n36# w_n206_n161# a_28_n25# a_n28_n69#
X0 a_28_n25# a_n28_n69# a_n120_n36# w_n206_n161# pfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
.ends

.subckt OR_magic A B OUT VDD VSS
Xnmos_3p3_H9QVWA_0 a_607_n374# VSS A VSS nmos_3p3_H9QVWA
Xnmos_3p3_H9QVWA_1 VSS a_607_n374# B VSS nmos_3p3_H9QVWA
Xnmos_3p3_H9QVWA_2 VSS OUT a_607_n374# VSS nmos_3p3_H9QVWA
Xpmos_3p3_M8RCNG_11 m1_267_n209# VDD a_607_n374# B pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_10 m1_267_n209# VDD a_607_n374# B pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_0 VDD VDD OUT a_607_n374# pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_1 VDD VDD m1_267_n209# A pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_2 VDD VDD OUT a_607_n374# pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_3 VDD VDD m1_267_n209# A pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_4 VDD VDD m1_267_n209# A pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_6 VDD VDD VDD VDD pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_7 VDD VDD m1_267_n209# A pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_8 m1_267_n209# VDD a_607_n374# B pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_9 m1_267_n209# VDD a_607_n374# B pmos_3p3_M8RCNG
.ends

.subckt nmos_3p3_F9QVWA a_140_n69# a_28_n25# a_n28_n69# a_n140_n25# a_n288_n36# a_196_n25#
+ a_n196_n69# VSUBS
X0 a_28_n25# a_n28_n69# a_n140_n25# VSUBS nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X1 a_196_n25# a_140_n69# a_28_n25# VSUBS nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X2 a_n140_n25# a_n196_n69# a_n288_n36# VSUBS nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
.ends

.subckt AND_3_magic B C OUT VDD VSS A
Xpmos_3p3_MGRCNG_0 VDD A VDD A VDD a_1469_n10# pmos_3p3_MGRCNG
Xpmos_3p3_MGRCNG_1 VDD a_1469_n10# VDD a_1469_n10# VDD OUT pmos_3p3_MGRCNG
Xnmos_3p3_H9QVWA_0 VSS OUT a_1469_n10# VSS nmos_3p3_H9QVWA
Xpmos_3p3_MGRCNG_2 VDD B VDD B VDD a_1469_n10# pmos_3p3_MGRCNG
Xpmos_3p3_MGRCNG_4 VDD C VDD C VDD a_1469_n10# pmos_3p3_MGRCNG
Xpmos_3p3_M8RCNG_0 VDD VDD VDD VDD pmos_3p3_M8RCNG
Xpmos_3p3_M8RCNG_1 VDD VDD VDD VDD pmos_3p3_M8RCNG
Xnmos_3p3_F9QVWA_0 B m1_603_n148# B m1_771_n286# m1_603_n148# m1_771_n286# B VSS nmos_3p3_F9QVWA
Xnmos_3p3_F9QVWA_2 C m1_771_n286# C VSS m1_771_n286# VSS C VSS nmos_3p3_F9QVWA
Xnmos_3p3_F9QVWA_1 A a_1469_n10# A m1_603_n148# a_1469_n10# m1_603_n148# A VSS nmos_3p3_F9QVWA
.ends

.subckt PGA_DECODER_magic A B C VDD S1 S2 S3 S4 S5 S6 AND_3_magic_5/C AND_3_magic_3/A
+ AND_3_magic_5/B VSS
XINVERTER_magic_0 A AND_3_magic_3/A VDD VSS INVERTER_magic
XAND_1 AND_1/A A S6 VDD VSS AND
XINVERTER_magic_1 C AND_3_magic_5/C VDD VSS INVERTER_magic
XINVERTER_magic_2 B AND_3_magic_5/B VDD VSS INVERTER_magic
XOR_magic_1 B C AND_1/A VDD VSS OR_magic
XAND_3_magic_0 AND_3_magic_5/B C S2 VDD VSS AND_3_magic_3/A AND_3_magic
XAND_3_magic_1 AND_3_magic_5/B AND_3_magic_5/C S1 VDD VSS AND_3_magic_3/A AND_3_magic
XAND_3_magic_2 B C S4 VDD VSS AND_3_magic_3/A AND_3_magic
XAND_3_magic_3 B AND_3_magic_5/C S3 VDD VSS AND_3_magic_3/A AND_3_magic
XAND_3_magic_5 AND_3_magic_5/B AND_3_magic_5/C S5 VDD VSS A AND_3_magic
.ends

.subckt pmos_3p3_MQ2VAR a_n52_n400# w_n282_n530# a_52_n444# a_108_n400# a_n108_n444#
+ a_n196_n400#
X0 a_108_n400# a_52_n444# a_n52_n400# w_n282_n530# pfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.28u
X1 a_n52_n400# a_n108_n444# a_n196_n400# w_n282_n530# pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.28u
.ends

.subckt pmos_3p3_MN7U2H a_n52_n313# w_n282_n443# a_52_n357# a_108_n313# a_n108_n357#
+ a_n196_n313#
X0 a_n52_n313# a_n108_n357# a_n196_n313# w_n282_n443# pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X1 a_108_n313# a_52_n357# a_n52_n313# w_n282_n443# pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
.ends

.subckt ppolyf_u_RRG95T a_n240_n722# a_n520_n722# a_320_620# a_n240_620# w_n704_n906#
+ a_n520_620# a_40_n722# a_320_n722# a_40_620#
X0 a_320_620# a_320_n722# w_n704_n906# ppolyf_u r_width=1u r_length=6.2u
X1 a_n520_620# a_n520_n722# w_n704_n906# ppolyf_u r_width=1u r_length=6.2u
X2 a_n240_620# a_n240_n722# w_n704_n906# ppolyf_u r_width=1u r_length=6.2u
X3 a_40_620# a_40_n722# w_n704_n906# ppolyf_u r_width=1u r_length=6.2u
.ends

.subckt nmos_3p3_FSHHD6 a_n52_n100# a_164_n100# a_n164_n144# a_n252_n100# a_52_n144#
+ VSUBS
X0 a_164_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X1 a_n52_n100# a_n164_n144# a_n252_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
.ends

.subckt nmos_3p3_V56RT2 a_n508_n144# a_n596_n100# a_n292_n100# a_28_n100# a_n452_n100#
+ a_n28_n144# a_132_n144# a_188_n100# a_n188_n144# a_292_n144# a_348_n100# a_n348_n144#
+ a_452_n144# a_508_n100# a_n132_n100# VSUBS
X0 a_n132_n100# a_n188_n144# a_n292_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_188_n100# a_132_n144# a_28_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n292_n100# a_n348_n144# a_n452_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_348_n100# a_292_n144# a_188_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_28_n100# a_n28_n144# a_n132_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_n452_n100# a_n508_n144# a_n596_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 a_508_n100# a_452_n144# a_348_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt pmos_3p3_HDY8L7 a_56_n694# a_n144_n694# a_n56_24# a_n144_68# a_n144_n1456#
+ a_n56_n738# a_n144_830# a_n56_n1500# a_56_830# a_56_68# a_n56_786# w_n230_n1586#
+ a_56_n1456#
X0 a_56_830# a_n56_786# a_n144_830# w_n230_n1586# pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.56u
X1 a_56_n694# a_n56_n738# a_n144_n694# w_n230_n1586# pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.56u
X2 a_56_n1456# a_n56_n1500# a_n144_n1456# w_n230_n1586# pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.56u
X3 a_56_68# a_n56_24# a_n144_68# w_n230_n1586# pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.56u
.ends

.subckt pmos_3p3_Q3NTJU a_428_68# a_428_n668# a_n1068_n1448# a_212_n1448# a_n748_n712#
+ a_n108_n1448# a_n852_68# a_n212_804# a_852_n712# a_52_n712# a_n428_760# a_692_24#
+ a_n908_24# a_108_n1404# a_n372_804# a_n52_n668# a_n852_n668# a_1012_24# a_n588_760#
+ a_n908_760# a_n1156_n1404# a_52_24# a_n52_68# a_n852_804# a_1068_n1404# a_268_68#
+ a_52_n1448# a_n1068_760# a_n1012_n668# a_n852_n1404# a_n372_n1404# a_532_24# a_n108_n712#
+ a_588_n668# a_n692_68# a_n1012_68# a_1012_n1448# a_212_n712# a_108_804# a_n908_n712#
+ a_n748_24# a_692_n1448# a_108_68# a_n1068_n712# a_n588_n1448# a_268_804# a_532_760#
+ a_n212_n668# a_1012_n712# a_1012_760# a_748_804# a_n1068_24# a_692_760# a_n532_68#
+ a_588_n1404# a_52_760# a_372_24# a_n212_n1404# a_n268_n712# a_n588_24# a_n908_n1448#
+ a_532_n1448# a_372_n712# a_748_n668# a_n428_n1448# a_212_24# a_n372_n668# a_n372_68#
+ a_908_n1404# a_428_n1404# a_n1012_n1404# a_n428_24# a_908_68# a_n108_760# a_n268_760#
+ a_n212_68# a_n532_804# a_108_n668# a_n692_n1404# a_n428_n712# a_n748_760# a_n692_804#
+ a_n1012_804# a_532_n712# a_908_n668# a_n52_804# a_n268_24# a_n532_n668# a_n52_n1404#
+ w_n1242_n1534# a_748_68# a_n1156_68# a_212_760# a_n532_n1404# a_372_760# a_428_804#
+ a_268_n668# a_1068_68# a_n588_n712# a_n108_24# a_588_804# a_908_804# a_852_760#
+ a_852_n1448# a_n1156_804# a_1068_804# a_692_n712# a_n748_n1448# a_372_n1448# a_1068_n668#
+ a_n1156_n668# a_n268_n1448# a_588_68# a_n692_n668# a_748_n1404# a_852_24# a_268_n1404#
X0 a_748_804# a_692_760# a_588_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1 a_n52_n1404# a_n108_n1448# a_n212_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X2 a_268_68# a_212_24# a_108_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X3 a_n372_68# a_n428_24# a_n532_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X4 a_108_n668# a_52_n712# a_n52_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X5 a_428_n668# a_372_n712# a_268_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X6 a_268_n668# a_212_n712# a_108_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X7 a_1068_n668# a_1012_n712# a_908_n668# w_n1242_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X8 a_268_n1404# a_212_n1448# a_108_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X9 a_108_804# a_52_760# a_n52_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X10 a_908_68# a_852_24# a_748_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X11 a_n212_n668# a_n268_n712# a_n372_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X12 a_n372_n1404# a_n428_n1448# a_n532_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X13 a_268_804# a_212_760# a_108_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X14 a_n852_n1404# a_n908_n1448# a_n1012_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X15 a_1068_n1404# a_1012_n1448# a_908_n1404# w_n1242_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X16 a_n212_68# a_n268_24# a_n372_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X17 a_n52_n668# a_n108_n712# a_n212_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X18 a_n852_n668# a_n908_n712# a_n1012_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X19 a_n372_804# a_n428_760# a_n532_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X20 a_n1012_n668# a_n1068_n712# a_n1156_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X21 a_n852_804# a_n908_760# a_n1012_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X22 a_428_804# a_372_760# a_268_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X23 a_588_n1404# a_532_n1448# a_428_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X24 a_908_804# a_852_760# a_748_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X25 a_n852_68# a_n908_24# a_n1012_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X26 a_748_68# a_692_24# a_588_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X27 a_908_n668# a_852_n712# a_748_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X28 a_n212_n1404# a_n268_n1448# a_n372_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X29 a_n1012_804# a_n1068_760# a_n1156_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X30 a_n52_68# a_n108_24# a_n212_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X31 a_n692_n1404# a_n748_n1448# a_n852_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X32 a_n532_804# a_n588_760# a_n692_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X33 a_108_68# a_52_24# a_n52_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X34 a_588_68# a_532_24# a_428_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X35 a_n692_n668# a_n748_n712# a_n852_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X36 a_428_n1404# a_372_n1448# a_268_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X37 a_n1012_68# a_n1068_24# a_n1156_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X38 a_n692_68# a_n748_24# a_n852_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X39 a_908_n1404# a_852_n1448# a_748_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X40 a_n1012_n1404# a_n1068_n1448# a_n1156_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X41 a_n532_n1404# a_n588_n1448# a_n692_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X42 a_748_n668# a_692_n712# a_588_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X43 a_n52_804# a_n108_760# a_n212_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X44 a_108_n1404# a_52_n1448# a_n52_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X45 a_588_n668# a_532_n712# a_428_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X46 a_588_804# a_532_760# a_428_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X47 a_428_68# a_372_24# a_268_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X48 a_748_n1404# a_692_n1448# a_588_n1404# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X49 a_n532_68# a_n588_24# a_n692_68# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X50 a_1068_68# a_1012_24# a_908_68# w_n1242_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X51 a_n532_n668# a_n588_n712# a_n692_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X52 a_n692_804# a_n748_760# a_n852_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X53 a_n212_804# a_n268_760# a_n372_804# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X54 a_1068_804# a_1012_760# a_908_804# w_n1242_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X55 a_n372_n668# a_n428_n712# a_n532_n668# w_n1242_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
.ends

.subckt nmos_3p3_QNHHD6 a_56_n100# a_n56_n144# a_n144_n100# VSUBS
X0 a_56_n100# a_n56_n144# a_n144_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.56u
.ends

.subckt pfet_03v3_6DHECV w_n202_n530# a_28_n400# a_n28_n444# a_n116_n400#
X0 a_28_n400# a_n28_n444# a_n116_n400# w_n202_n530# pfet_03v3 ad=1.76p pd=8.88u as=1.76p ps=8.88u w=4u l=0.28u
.ends

.subckt nmos_3p3_6F3WC4 a_100_n468# a_n100_24# a_n188_68# a_n100_n512# a_n188_n468#
+ a_100_68# VSUBS
X0 a_100_68# a_n100_24# a_n188_68# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=1u
X1 a_100_n468# a_n100_n512# a_n188_n468# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=1u
.ends

.subckt ppolyf_u_RKG95T a_n100_620# a_n100_n722# w_n284_n906#
X0 a_n100_620# a_n100_n722# w_n284_n906# ppolyf_u r_width=1u r_length=6.2u
.ends

.subckt nmos_3p3_BSHHD6 a_596_n100# a_268_n144# a_n596_n144# a_n52_n100# a_484_n144#
+ a_n684_n100# a_164_n100# a_380_n100# a_n164_n144# a_n380_n144# a_52_n144# a_n268_n100#
+ a_n484_n100# VSUBS
X0 a_n268_n100# a_n380_n144# a_n484_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X1 a_n484_n100# a_n596_n144# a_n684_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X2 a_380_n100# a_268_n144# a_164_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X3 a_164_n100# a_52_n144# a_n52_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X4 a_596_n100# a_484_n144# a_380_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X5 a_n52_n100# a_n164_n144# a_n268_n100# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
.ends

.subckt pmos_3p3_MANNAR a_28_n1404# a_28_n668# a_n28_n1448# a_n116_n668# a_n116_n1404#
+ a_28_68# a_n116_804# a_28_804# a_n28_n712# a_n28_24# a_n116_68# w_n202_n1534# a_n28_760#
X0 a_28_68# a_n28_24# a_n116_68# w_n202_n1534# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X1 a_28_804# a_n28_760# a_n116_804# w_n202_n1534# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X2 a_28_n668# a_n28_n712# a_n116_n668# w_n202_n1534# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X3 a_28_n1404# a_n28_n1448# a_n116_n1404# w_n202_n1534# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt pmos_3p3_MEKUKR w_n202_n380# a_28_n250# a_n28_n294# a_n116_n250#
X0 a_28_n250# a_n28_n294# a_n116_n250# w_n202_n380# pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
.ends

.subckt nmos_3p3_3AEFT2 a_56_n100# a_n56_n144# a_n144_n100# VSUBS
X0 a_56_n100# a_n56_n144# a_n144_n100# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.56u
.ends

.subckt pmos_3p3_M82RNG a_n28_n94# w_n202_n180# a_n116_n50# a_28_n50#
X0 a_28_n50# a_n28_n94# a_n116_n50# w_n202_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt PGA_MAGIC BD IND IPD VSS VB4 VB2 VB3 VB1 VND VPD IBIAS1 VBIASN VOUT VBM VCD
+ IBIAS4 IBIAS3 IBS OUT_P OUT_N IBIAS2 IBIAS VCM IVS IB4 IB2 IB3 IB5 IN_P IN_N OUT1
+ OUT2 VIN_P VIN_N S_PGA_1 S_PGA_2 S_PGA_3 VDD
Xpmos_3p3_ME7U2H_2 VND VB1 VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_1 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_876RT2_10 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xnmos_3p3_3A6RT2_7 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_4 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_71 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_82 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_93 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_60 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_6 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_MA2VAR_106 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_67 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_45 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_56 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_15 VDD VB1 VND VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_26 OUT2 VB2 VPD VDD pmos_3p3_ME7U2H
Xnmos_3p3_276RTJ_3 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_12 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_23 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_34 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xnmos_3p3_2F3WC4_1 VSS IVS IVS IVS IVS IVS VSS IVS VSS IVS IVS IVS IVS VSS IVS IVS
+ IVS IVS IVS IVS VSS VSS VSS nmos_3p3_2F3WC4
Xpmos_3p3_MA2VAR_28 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_17 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_39 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xnmos_3p3_NE3WC4_0 VSS VSS VSS VSS nmos_3p3_NE3WC4
Xppolyf_u_2VJWHK_7 VDD VDD VDD ppolyf_u_2VJWHK
Xnmos_3p3_EA6RT2_0 IB5 VB4 IB5 VB4 VB4 IB5 IB5 IB5 IB5 VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_3 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_2 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_876RT2_11 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xpmos_3p3_5L6RD7_1 VDD IBIAS1 IBIAS1 VDD pmos_3p3_5L6RD7
Xnmos_3p3_3A6RT2_8 VCD VOUT VB1 VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_5 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_50 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_72 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_94 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_61 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_83 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_20 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_S75EG7_0 VB4 VB4 VSS VB4 VB4 VB4 VB4 VSS VB4 VB4 VB4 VSS VB4 VB4 VSS VB4
+ VSS VB4 VB4 VB4 VB4 VSS VB4 VB4 VB4 VB4 VSS VB4 VB4 VSS nmos_3p3_S75EG7
Xpmos_3p3_MNS6FR_7 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_MA2VAR_107 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_4 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_ME7U2H_16 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_68 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_46 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_24 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_57 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_27 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_13 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_35 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_NE3WC4_1 VSS VSS VSS VSS nmos_3p3_NE3WC4
Xpmos_3p3_MA2VAR_29 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_18 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_EA6RT2_1 VCM VCD VCM VCD VCD VBM VBM VCM VCM VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_4 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_3 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_876RT2_0 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_5L6RD7_2 VDD VDD IBIAS1 VBIASN pmos_3p3_5L6RD7
Xnmos_3p3_3A6RT2_9 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_6 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_51 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_40 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_73 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_84 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_95 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_62 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xnmos_3p3_5J7TC4_0 VSS IBS VSS IBIAS IBS VSS nmos_3p3_5J7TC4
Xpmos_3p3_MNS6FR_8 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_MA2VAR_108 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_3A6RT2_21 VBM VCM VCD VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_10 VB1 VOUT VCD VSS nmos_3p3_3A6RT2
Xnmos_3p3_276RTJ_5 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_69 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_47 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_25 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_17 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_14 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_28 VND VB2 OUT1 VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_36 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_58 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_19 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xnmos_3p3_NE3WC4_2 VSS VBIASN IBIAS4 VSS nmos_3p3_NE3WC4
Xnmos_3p3_EA6RT2_2 VOUT VCD VOUT VCD VCD VB1 VB1 VOUT VOUT VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_5 VPD VB1 VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_4 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MYZUAR_0 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xnmos_3p3_876RT2_1 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xnmos_3p3_7WQWW2_7 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_52 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_41 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_30 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_74 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_85 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_96 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_63 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_5J7TC4_1 VSS IBS VSS IBS IBS VSS nmos_3p3_5J7TC4
Xpmos_3p3_MNS6FR_9 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xnmos_3p3_3A6RT2_22 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_11 VCD VCM VBM VSS nmos_3p3_3A6RT2
Xnmos_3p3_276RTJ_6 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_MA2VAR_109 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_48 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_26 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_59 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_18 VPD VB2 OUT2 VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_15 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_29 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_37 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
XTGATE_PGA_MAGIC_0 VDD VSS IN_P TGATE_PGA_MAGIC_0/CLK TGATE_PGA_MAGIC_0/A TGATE_PGA_MAGIC
Xnmos_3p3_EA6RT2_3 VOUT VCD VOUT VCD VCD VB1 VB1 VOUT VOUT VSS nmos_3p3_EA6RT2
Xpga_res_magice_parallel_0 VDD TGATE_PGA_MAGIC_1/A TGATE_PGA_MAGIC_0/A TGATE_PGA_MAGIC_3/A
+ OUT_N TGATE_PGA_MAGIC_2/A TGATE_PGA_MAGIC_4/A TGATE_PGA_MAGIC_5/A VIN_P pga_res_magice_parallel
Xpmos_3p3_ME7U2H_6 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_5 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MYZUAR_1 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xpmos_3p3_MAEVAR_0 VDD VDD VDD VDD VDD VDD VDD pmos_3p3_MAEVAR
Xnmos_3p3_876RT2_2 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xnmos_3p3_7WQWW2_8 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_53 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_20 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_42 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_31 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_75 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_86 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_64 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_97 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_23 VCD VOUT VB1 VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_12 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_276RTJ_7 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_27 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_49 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_19 OUT2 VB2 VPD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_16 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_38 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
XTGATE_PGA_MAGIC_1 VDD VSS IN_P TGATE_PGA_MAGIC_9/CLK TGATE_PGA_MAGIC_1/A TGATE_PGA_MAGIC
Xnmos_3p3_EA6RT2_4 VCM VCD VCM VCD VCD VBM VBM VCM VCM VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_7 VND VB1 VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_6 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MYZUAR_2 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xpga_res_magice_parallel_1 VDD TGATE_PGA_MAGIC_9/A TGATE_PGA_MAGIC_10/A TGATE_PGA_MAGIC_8/A
+ OUT_P TGATE_PGA_MAGIC_11/A TGATE_PGA_MAGIC_7/A TGATE_PGA_MAGIC_6/A VIN_N pga_res_magice_parallel
Xnmos_3p3_876RT2_3 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xnmos_3p3_7WQWW2_9 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_21 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_54 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_43 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_10 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_32 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_76 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_87 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_65 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_98 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_24 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_13 VB1 VOUT VCD VSS nmos_3p3_3A6RT2
Xnmos_3p3_M86RTJ_28 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_276RTJ_8 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_17 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_39 VSS VSS VSS VSS nmos_3p3_M86RTJ
XTGATE_PGA_MAGIC_2 VDD VSS IN_P TGATE_PGA_MAGIC_2/CLK TGATE_PGA_MAGIC_2/A TGATE_PGA_MAGIC
Xnmos_3p3_EA6RT2_5 VCM VCD VCM VCD VCD VBM VBM VCM VCM VSS nmos_3p3_EA6RT2
Xpmos_3p3_MES6FR_0 VDD IND BD IN_N pmos_3p3_MES6FR
Xpmos_3p3_MYZUAR_3 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xpmos_3p3_ME7U2H_8 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_7 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_RKK9DS_0 IB2 VB2 VB2 IB2 IB2 VB2 VB2 VB2 VB2 VB2 VB2 VB2 IB2 VB2 VB2 VB2
+ VB2 VB2 VDD VB2 IB2 VB2 IB2 IB2 VB2 VB2 VB2 VB2 VB2 VB2 VB2 IB2 IB2 VB2 pmos_3p3_RKK9DS
Xnmos_3p3_876RT2_4 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_22 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_55 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_44 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_11 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_33 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_77 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_88 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_66 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_99 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_25 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_14 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_276RTJ_9 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_29 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_18 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xcap_mim_2p0fF_3FUNHB_0 OUT_P m1_29250_n5500# cap_mim_2p0fF_3FUNHB
XTGATE_PGA_MAGIC_3 VDD VSS IN_P TGATE_PGA_MAGIC_8/CLK TGATE_PGA_MAGIC_3/A TGATE_PGA_MAGIC
Xnmos_3p3_EA6RT2_6 VOUT VCD VOUT VCD VCD VB1 VB1 VOUT VOUT VSS nmos_3p3_EA6RT2
Xpmos_3p3_5UYQD7_0 VB3 VDD IBIAS1 VDD IBIAS1 VDD pmos_3p3_5UYQD7
Xpmos_3p3_MYZUAR_4 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xpmos_3p3_MES6FR_1 VDD BD IND IN_N pmos_3p3_MES6FR
Xpmos_3p3_ME7U2H_9 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_8 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xnmos_3p3_876RT2_5 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_23 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_45 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_12 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_34 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_78 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_89 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_67 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_56 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_5LZQD7_0 VDD IBIAS1 IBS IBIAS1 IBS IBS VDD IBIAS1 IBIAS1 IBIAS1 VDD VDD
+ pmos_3p3_5LZQD7
Xnmos_3p3_3A6RT2_26 VB1 VOUT VCD VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_15 VCD VOUT VB1 VSS nmos_3p3_3A6RT2
Xnmos_3p3_M86RTJ_19 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xcap_mim_2p0fF_3FUNHB_1 OUT_N m1_29250_n7512# cap_mim_2p0fF_3FUNHB
XTGATE_PGA_MAGIC_4 VDD VSS IN_P TGATE_PGA_MAGIC_7/CLK TGATE_PGA_MAGIC_4/A TGATE_PGA_MAGIC
Xpmos_3p3_MES6FR_2 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MA2VAR_9 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MYZUAR_5 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xnmos_3p3_876RT2_6 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_24 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_46 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_35 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_13 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_79 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_57 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_68 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_5LZQD7_1 VDD IBIAS IBIAS IBIAS IBIAS IBIAS VDD IBIAS IBIAS IBIAS VDD VDD
+ pmos_3p3_5LZQD7
Xnmos_3p3_3A6RT2_16 VSS VSS VSS VSS nmos_3p3_3A6RT2
XTGATE_PGA_MAGIC_5 VDD VSS IN_P TGATE_PGA_MAGIC_6/CLK TGATE_PGA_MAGIC_5/A TGATE_PGA_MAGIC
Xpmos_3p3_MES6FR_3 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MYZUAR_6 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xpmos_3p3_5C3RD7_0 IBIAS1 VDD VDD VDD IB5 IBIAS1 IBIAS1 IBIAS1 IB5 VDD pmos_3p3_5C3RD7
Xnmos_3p3_876RT2_7 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_HMY8L7_0 VDD BD BD IBIAS VDD VDD BD IBIAS IBIAS BD VDD VDD IBIAS VDD BD
+ VDD IBIAS IBIAS VDD IBIAS VDD IBIAS BD VDD IBIAS VDD IBIAS IBIAS IBIAS VDD IBIAS
+ VDD BD IBIAS IBIAS IBIAS VDD IBIAS IBIAS BD VDD BD IBIAS VDD IBIAS VDD VDD BD BD
+ IBIAS BD BD IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS BD IBIAS BD BD
+ IBIAS VDD VDD VDD pmos_3p3_HMY8L7
Xpmos_3p3_M22VAR_25 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_47 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_14 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_36 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_58 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_69 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_17 VBM VCM VCD VSS nmos_3p3_3A6RT2
Xpmos_3p3_K823KY_0 VDD VB2 IB2 VDD pmos_3p3_K823KY
XTGATE_PGA_MAGIC_6 VDD VSS IN_N TGATE_PGA_MAGIC_6/CLK TGATE_PGA_MAGIC_6/A TGATE_PGA_MAGIC
Xpmos_3p3_MES6FR_4 VDD BD IPD IN_P pmos_3p3_MES6FR
Xnmos_3p3_876RT2_8 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_26 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_48 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_15 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_37 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_59 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_18 VSS VSS VSS VSS nmos_3p3_3A6RT2
XTGATE_PGA_MAGIC_7 VDD VSS IN_N TGATE_PGA_MAGIC_7/CLK TGATE_PGA_MAGIC_7/A TGATE_PGA_MAGIC
Xpmos_3p3_MES6FR_5 VDD IPD BD IN_P pmos_3p3_MES6FR
Xnmos_3p3_U56RT2_0 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS nmos_3p3_U56RT2
Xnmos_3p3_JE3WC4_0 VSS IBIAS3 IB4 IBIAS3 VSS IB4 IB4 VSS IBIAS3 IB4 IB4 VSS nmos_3p3_JE3WC4
Xppolyf_u_2V2ZHK_0 m1_26256_n7401# m1_26536_n6269# m1_26256_n7401# VDD m1_25080_n6269#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_MNS6FR_10 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xnmos_3p3_876RT2_9 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_27 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_49 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_16 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_38 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_19 VCD VCM VBM VSS nmos_3p3_3A6RT2
Xnmos_3p3_UUQWW2_0 VB3 OUT1 IND VSS nmos_3p3_UUQWW2
Xpmos_3p3_M2NNAR_0 IBIAS4 IBIAS4 VDD IB4 IBIAS4 IB4 IBIAS4 IBIAS4 VDD VDD VDD IBIAS4
+ VDD IBIAS4 VDD IB4 IB4 VDD VDD IBIAS4 VDD pmos_3p3_M2NNAR
XTGATE_PGA_MAGIC_8 VDD VSS IN_N TGATE_PGA_MAGIC_8/CLK TGATE_PGA_MAGIC_8/A TGATE_PGA_MAGIC
Xnmos_3p3_JE3WC4_1 IB4 VSS IB4 VSS IB4 IB4 IB4 IB4 VSS IB4 IB4 VSS nmos_3p3_JE3WC4
Xpmos_3p3_MES6FR_6 VDD IND BD IN_N pmos_3p3_MES6FR
Xppolyf_u_2V2ZHK_1 m1_24352_n7688# m1_24072_n6269# OUT_N VDD m1_24072_n6269# ppolyf_u_2V2ZHK
Xpmos_3p3_MNS6FR_11 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_M22VAR_17 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_39 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_28 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_UUQWW2_1 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_M2NNAR_1 IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD
+ IBIAS3 VDD IBIAS3 VDD IBIAS3 IBIAS3 VDD VDD IBIAS3 VDD pmos_3p3_M2NNAR
XTGATE_PGA_MAGIC_9 VDD VSS IN_N TGATE_PGA_MAGIC_9/CLK TGATE_PGA_MAGIC_9/A TGATE_PGA_MAGIC
Xpmos_3p3_MES6FR_7 VDD BD IND IN_N pmos_3p3_MES6FR
Xppolyf_u_2V2ZHK_2 m1_24800_n7401# m1_25080_n6269# m1_24800_n7401# VDD m1_23624_n6269#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_MNS6FR_12 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_M22VAR_18 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
XPGA_DECODER_magic_0 PGA_DECODER_magic_0/A PGA_DECODER_magic_0/B PGA_DECODER_magic_0/C
+ VDD TGATE_PGA_MAGIC_2/CLK TGATE_PGA_MAGIC_6/CLK TGATE_PGA_MAGIC_7/CLK TGATE_PGA_MAGIC_8/CLK
+ TGATE_PGA_MAGIC_9/CLK TGATE_PGA_MAGIC_0/CLK S_PGA_1 S_PGA_3 S_PGA_2 VSS PGA_DECODER_magic
Xpmos_3p3_M22VAR_29 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_UUQWW2_2 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MES6FR_8 VDD IND BD IN_N pmos_3p3_MES6FR
Xppolyf_u_2V2ZHK_3 m1_25808_n7688# m1_25528_n6269# m1_24352_n7688# VDD m1_25528_n6269#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_MNS6FR_13 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_M22VAR_19 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_UUQWW2_3 VB3 IND OUT1 VSS nmos_3p3_UUQWW2
Xpmos_3p3_MQ2VAR_0 VBM VDD VBM VDD VBM VDD pmos_3p3_MQ2VAR
Xpmos_3p3_MES6FR_9 VDD BD IND IN_N pmos_3p3_MES6FR
Xppolyf_u_2V2ZHK_4 m1_26536_n5429# m1_26256_n4297# m1_25080_n5716# VDD m1_26256_n4297#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_MNS6FR_14 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xnmos_3p3_UUQWW2_40 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MQ2VAR_1 VB1 VDD VB1 VDD VB1 VDD pmos_3p3_MQ2VAR
Xnmos_3p3_UUQWW2_4 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_M22VAR_190 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xppolyf_u_2V2ZHK_5 m1_25528_n5429# m1_25808_n4297# m1_25528_n5429# VDD m1_24352_n4297#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_MNS6FR_15 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_MN7U2H_20 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xppolyf_u_RRG95T_0 m1_29250_n7512# m1_29250_n7512# OUT1 OUT1 VDD OUT1 m1_29250_n7512#
+ m1_29250_n7512# OUT1 ppolyf_u_RRG95T
Xnmos_3p3_UUQWW2_30 VB4 IPD VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_41 VB4 VSS IPD VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_5 VB3 IND OUT1 VSS nmos_3p3_UUQWW2
Xpmos_3p3_M22VAR_180 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_191 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_FSHHD6_0 VBIASN VSS VBIASN VSS VBIASN VSS nmos_3p3_FSHHD6
Xppolyf_u_2V2ZHK_6 m1_25080_n5716# m1_24800_n4297# m1_23624_n5716# VDD m1_24800_n4297#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_MNS6FR_16 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_MN7U2H_21 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xpmos_3p3_MN7U2H_10 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_V56RT2_0 VB3 IB3 IB3 IB3 VB3 VB3 VB3 VB3 VB3 VB3 IB3 VB3 VB3 VB3 VB3 VSS
+ nmos_3p3_V56RT2
Xppolyf_u_RRG95T_1 m1_29250_n5500# m1_29250_n5500# OUT2 OUT2 VDD OUT2 m1_29250_n5500#
+ m1_29250_n5500# OUT2 ppolyf_u_RRG95T
Xnmos_3p3_UUQWW2_20 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_31 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_42 VB4 IPD VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_6 VB3 OUT1 IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_30 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_181 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_192 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_170 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xppolyf_u_2V2ZHK_7 m1_24072_n5429# m1_24352_n4297# m1_24072_n5429# VDD VOUT ppolyf_u_2V2ZHK
Xpmos_3p3_MNS6FR_17 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_M22VAR_0 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_22 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xpmos_3p3_MN7U2H_11 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_21 VB4 IND VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_10 VB3 IPD OUT2 VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_32 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_43 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_7 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_20 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_31 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_160 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_193 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_171 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_182 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_1 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_12 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xpmos_3p3_MN7U2H_23 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_44 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_22 VB4 VSS IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_8 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_11 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_33 VB4 VSS IPD VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_21 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_10 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_32 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_161 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_150 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_194 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_172 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_183 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_2 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_13 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_45 VB4 VSS IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_23 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_12 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_34 VB4 IPD VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_9 VB3 OUT2 IPD VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_33 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_22 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_11 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_162 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_173 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_140 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_151 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_195 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_184 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_HDY8L7_0 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pmos_3p3_HDY8L7
Xnmos_3p3_276RTJ_50 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_Q3NTJU_0 VDD VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD VDD IBIAS3 IBIAS3 IBIAS3
+ IBIAS3 IBIAS3 VDD IVS IVS VDD IBIAS3 IBIAS3 IBIAS3 VDD IBIAS3 IVS VDD VDD IVS IBIAS3
+ IBIAS3 IVS VDD IVS IBIAS3 IBIAS3 IVS IVS IVS IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3
+ VDD IBIAS3 IBIAS3 IVS IBIAS3 VDD IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 VDD IVS IBIAS3
+ IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IVS IVS IVS VDD
+ IVS IBIAS3 IVS IBIAS3 IBIAS3 VDD VDD VDD IVS IBIAS3 IBIAS3 IVS IVS IBIAS3 IVS IVS
+ IBIAS3 VDD IVS VDD VDD VDD IBIAS3 VDD IBIAS3 VDD IVS VDD IBIAS3 IBIAS3 IVS IVS IBIAS3
+ IBIAS3 VDD VDD IBIAS3 IBIAS3 IBIAS3 VDD VDD IBIAS3 IVS IVS VDD IBIAS3 IVS pmos_3p3_Q3NTJU
Xpmos_3p3_M22VAR_3 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_14 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_46 VB4 IND VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_24 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_35 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_13 VB3 OUT2 IPD VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_34 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_12 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_23 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_163 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_174 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_141 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_152 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_185 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_130 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_HDY8L7_1 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pmos_3p3_HDY8L7
Xpmos_3p3_MA2VAR_90 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_51 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_40 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_QNHHD6_0 VSS VBIASN VB2 VSS nmos_3p3_QNHHD6
Xpmos_3p3_M22VAR_4 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_15 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_47 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_25 VB4 VSS IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_36 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_14 VB3 IPD OUT2 VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_0 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_35 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_13 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_24 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_164 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_142 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_120 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_153 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_131 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_175 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_91 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_80 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_186 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_30 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_52 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_41 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_M22VAR_5 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_16 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_37 VB4 VSS IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_26 VB4 IND VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_15 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_1 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_14 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_25 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_110 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_70 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_165 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_143 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_81 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_121 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_187 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_132 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_154 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_92 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_176 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_31 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_53 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_20 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_42 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_M22VAR_6 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MES6FR_20 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MN7U2H_17 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_16 VB4 VSS IPD VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_2 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_27 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_38 VB4 IND VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_15 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_26 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_111 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_60 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_71 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_100 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_133 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_166 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_144 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_122 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_82 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_188 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_155 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_177 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_93 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_32 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_21 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_10 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_43 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpfet_03v3_6DHECV_0 VDD VDD VDD VDD pfet_03v3_6DHECV
Xpmos_3p3_M22VAR_7 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_6F3WC4_0 VSS VSS VSS VSS VSS VSS VSS nmos_3p3_6F3WC4
Xpmos_3p3_MES6FR_21 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MES6FR_10 VDD BD IPD IN_P pmos_3p3_MES6FR
Xpmos_3p3_MN7U2H_18 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xppolyf_u_RKG95T_0 VDD VDD VDD ppolyf_u_RKG95T
Xnmos_3p3_UUQWW2_17 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_28 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_39 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_3 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_16 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_27 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_M86RTJ_0 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_61 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_50 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_101 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_72 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_134 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_167 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_112 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_145 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_178 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_123 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_83 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_156 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_94 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_189 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_33 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_22 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_11 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_44 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_M22VAR_8 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_6F3WC4_1 VSS VSS VSS VSS VSS VSS VSS nmos_3p3_6F3WC4
Xpmos_3p3_MES6FR_22 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MES6FR_11 VDD IPD BD IN_P pmos_3p3_MES6FR
Xpmos_3p3_MN7U2H_19 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xppolyf_u_RKG95T_1 VDD VDD VDD ppolyf_u_RKG95T
Xnmos_3p3_UUQWW2_18 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_29 VB4 VSS IPD VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_4 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_17 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_28 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_M86RTJ_1 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_40 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_102 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_135 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_168 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_113 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_146 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_179 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_124 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_157 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_62 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_51 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_73 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_84 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_95 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_34 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_23 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_12 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_45 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_BSHHD6_0 VSS VBIASN VBIASN VCD VBIASN VSS VSS VCD VBIASN VBIASN VBIASN VSS
+ VCD VSS nmos_3p3_BSHHD6
Xpmos_3p3_M22VAR_9 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_6F3WC4_2 VSS VSS VSS VSS VSS VSS VSS nmos_3p3_6F3WC4
Xpmos_3p3_MES6FR_12 VDD IND BD IN_N pmos_3p3_MES6FR
Xpmos_3p3_MES6FR_23 VDD VDD VDD VDD pmos_3p3_MES6FR
Xppolyf_u_RKG95T_2 VDD VDD VDD ppolyf_u_RKG95T
Xnmos_3p3_UUQWW2_19 VB4 IPD VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_5 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_18 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_29 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_M86RTJ_2 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_M22VAR_103 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_136 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_169 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_114 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_125 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_147 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_158 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_30 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_41 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_63 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_52 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_74 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_85 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_96 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_35 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_13 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_46 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_24 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_MES6FR_13 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MANNAR_0 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pmos_3p3_MANNAR
Xppolyf_u_RKG95T_3 VDD VDD VDD ppolyf_u_RKG95T
Xpmos_3p3_MN7U2H_6 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_M86RTJ_70 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_7WQWW2_19 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_M86RTJ_3 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_31 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_20 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_42 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_64 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_104 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_53 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_137 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_97 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_115 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_86 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_75 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_148 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_126 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_159 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_36 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_14 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_47 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_25 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_3A6RT2_0 VSS VSS VSS VSS nmos_3p3_3A6RT2
XTGATE_PGA_MAGIC_10 VDD VSS IN_N TGATE_PGA_MAGIC_0/CLK TGATE_PGA_MAGIC_10/A TGATE_PGA_MAGIC
Xpmos_3p3_MES6FR_14 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MANNAR_1 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pmos_3p3_MANNAR
Xpmos_3p3_MN7U2H_7 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xpmos_3p3_MEKUKR_0 VDD VDD IBIAS4 IBIAS4 pmos_3p3_MEKUKR
Xpmos_3p3_MA2VAR_110 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_71 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_30 OUT1 VB2 VND VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_60 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_4 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_10 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_21 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_105 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_76 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_43 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_54 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_65 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_32 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_138 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_98 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_116 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_149 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_127 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_87 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_0 m1_23624_n6269# OUT_P VDD ppolyf_u_2VJWHK
Xnmos_3p3_276RTJ_48 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_37 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_15 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_26 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_3A6RT2_1 VSS VSS VSS VSS nmos_3p3_3A6RT2
XTGATE_PGA_MAGIC_11 VDD VSS IN_N TGATE_PGA_MAGIC_2/CLK TGATE_PGA_MAGIC_11/A TGATE_PGA_MAGIC
Xpmos_3p3_MES6FR_15 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MNS6FR_0 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_MN7U2H_8 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xpmos_3p3_MA2VAR_111 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MEKUKR_1 VDD VDD IBIAS4 IBIAS4 pmos_3p3_MEKUKR
Xpmos_3p3_ME7U2H_20 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_31 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_61 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_100 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_50 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_5 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_11 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_22 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_106 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_55 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_33 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_44 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_66 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_139 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_77 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_117 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_88 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_128 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_99 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_1 VDD VDD VDD ppolyf_u_2VJWHK
Xnmos_3p3_276RTJ_49 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_38 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_16 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_27 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_3AEFT2_0 IB3 VB3 VSS VSS nmos_3p3_3AEFT2
Xnmos_3p3_3A6RT2_2 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_16 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MNS6FR_1 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_MN7U2H_9 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_M86RTJ_40 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_101 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_ME7U2H_21 VND VB2 OUT1 VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_10 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_51 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_62 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_6 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_12 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_23 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_107 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_34 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_45 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_56 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_118 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_129 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xppolyf_u_2VJWHK_2 m1_25808_n4297# m1_26536_n6269# VDD ppolyf_u_2VJWHK
Xpmos_3p3_MA2VAR_78 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_89 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_67 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_39 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_17 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_28 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_3A6RT2_3 VCD VCM VBM VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_0 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_MES6FR_17 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MNS6FR_2 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_MA2VAR_102 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_ME7U2H_11 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_41 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_52 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_30 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_22 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_7 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_63 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_M22VAR_108 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_119 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xppolyf_u_2VJWHK_3 VOUT m1_23624_n5716# VDD ppolyf_u_2VJWHK
Xpmos_3p3_MA2VAR_13 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_24 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_35 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_46 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_57 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_79 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_68 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_18 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_29 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_M82RNG_0 VDD VDD VDD VDD pmos_3p3_M82RNG
Xnmos_3p3_3A6RT2_4 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_18 VDD BD IND IN_N pmos_3p3_MES6FR
Xnmos_3p3_7WQWW2_1 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_90 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_3 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_MA2VAR_103 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_0 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_64 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_42 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_53 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_31 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_23 OUT1 VB2 VND VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_8 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_12 VDD VB1 VND VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_20 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_14 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_25 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_109 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_36 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_47 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_58 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_69 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_4 m1_26536_n5429# m1_25808_n7688# VDD ppolyf_u_2VJWHK
Xnmos_3p3_276RTJ_19 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_ME7U2H_0 VPD VB1 VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_M82RNG_1 VDD VDD VDD VDD pmos_3p3_M82RNG
Xnmos_3p3_3A6RT2_5 VBM VCM VCD VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_19 VDD VDD VDD VDD pmos_3p3_MES6FR
Xnmos_3p3_7WQWW2_2 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_80 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_91 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_4 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xnmos_3p3_276RTJ_1 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_MA2VAR_104 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_43 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_65 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_54 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_24 VPD VB2 OUT2 VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_10 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_13 VDD VB1 VPD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_21 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_32 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_9 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_15 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_26 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_37 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_48 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_59 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_5 VDD VDD VDD ppolyf_u_2VJWHK
Xpmos_3p3_ME7U2H_1 VDD VB1 VPD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_0 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xnmos_3p3_3A6RT2_6 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_3 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_70 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_81 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_92 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_5 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xnmos_3p3_276RTJ_2 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_MA2VAR_105 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_66 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_44 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_55 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_2F3WC4_0 IBIAS2 VSS IVS IVS VSS IVS IBIAS2 IVS IBIAS2 VSS IVS IVS VSS IBIAS2
+ IVS IVS IVS IVS VSS VSS IBIAS2 IBIAS2 VSS nmos_3p3_2F3WC4
Xpmos_3p3_ME7U2H_25 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_11 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_14 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_22 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_33 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_27 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_16 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_38 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_49 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_6 VDD VDD VDD ppolyf_u_2VJWHK
.ends

.subckt ppolyf_u_3VY3SR w_n1124_n1136# a_460_850# a_n380_850# a_180_n952# a_n100_850#
+ a_460_n952# a_740_n952# a_n100_n952# a_740_850# a_n380_n952# a_n660_850# a_n660_n952#
+ a_180_850# a_n940_n952# a_n940_850#
X0 a_460_850# a_460_n952# w_n1124_n1136# ppolyf_u r_width=1u r_length=8.5u
X1 a_180_850# a_180_n952# w_n1124_n1136# ppolyf_u r_width=1u r_length=8.5u
X2 a_n940_850# a_n940_n952# w_n1124_n1136# ppolyf_u r_width=1u r_length=8.5u
X3 a_n660_850# a_n660_n952# w_n1124_n1136# ppolyf_u r_width=1u r_length=8.5u
X4 a_n100_850# a_n100_n952# w_n1124_n1136# ppolyf_u r_width=1u r_length=8.5u
X5 a_n380_850# a_n380_n952# w_n1124_n1136# ppolyf_u r_width=1u r_length=8.5u
X6 a_740_850# a_740_n952# w_n1124_n1136# ppolyf_u r_width=1u r_length=8.5u
.ends

.subckt VCM_1.3V_magic VDD VSS VCM_1.3
Xppolyf_u_3VY3SR_0 VDD m1_905_2023# m1_626_1599# VCM_1.3 m1_905_2023# VCM_1.3 VDD
+ m1_345_n120# VDD VSS VDD m1_345_n120# m1_626_1599# VDD VDD ppolyf_u_3VY3SR
.ends

.subckt pmos_3p3_9K6RD7 a_56_n300# a_n56_n344# a_n144_n300# w_n230_n430#
X0 a_56_n300# a_n56_n344# a_n144_n300# w_n230_n430# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.56u
.ends

.subckt pmos_3p3_VK6RD7 w_n230_n330# a_56_n200# a_n56_n244# a_n144_n200#
X0 a_56_n200# a_n56_n244# a_n144_n200# w_n230_n330# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.56u
.ends

.subckt pmos_3p3_HWZ2RY a_100_n468# w_n274_n598# a_n100_24# a_n188_68# a_n100_n512#
+ a_n188_n468# a_100_68#
X0 a_100_68# a_n100_24# a_n188_68# w_n274_n598# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=1u
X1 a_100_n468# a_n100_n512# a_n188_n468# w_n274_n598# pfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=1u
.ends

.subckt pmos_3p3_MAJNAR a_n28_392# a_n116_n1772# a_n28_n1816# a_28_n1036# a_n116_n1036#
+ a_28_1172# a_n28_n1080# a_n116_436# a_n116_1172# a_28_n300# a_28_436# a_n28_1128#
+ a_n28_n344# a_n116_n300# a_28_n1772# w_n202_n1902#
X0 a_28_1172# a_n28_1128# a_n116_1172# w_n202_n1902# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X1 a_28_n1772# a_n28_n1816# a_n116_n1772# w_n202_n1902# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X2 a_28_436# a_n28_392# a_n116_436# w_n202_n1902# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X3 a_28_n300# a_n28_n344# a_n116_n300# w_n202_n1902# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X4 a_28_n1036# a_n28_n1080# a_n116_n1036# w_n202_n1902# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt pmos_3p3_VTYQD7 a_n52_n200# a_164_n200# a_n164_n244# a_n252_n200# a_52_n244#
+ w_n338_n330#
X0 a_164_n200# a_52_n244# a_n52_n200# w_n338_n330# pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.56u
X1 a_n52_n200# a_n164_n244# a_n252_n200# w_n338_n330# pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.56u
.ends

.subckt cap_mim_2p0fF_XHV85N m4_n2640_n3400# m4_n2520_n3280#
X0 m4_n2520_n3280# m4_n2640_n3400# cap_mim_2f0_m4m5_noshield c_width=24u c_length=15.5u
X1 m4_n2520_n3280# m4_n2640_n3400# cap_mim_2f0_m4m5_noshield c_width=24u c_length=15.5u
.ends

.subckt nmos_3p3_NQ5EG7 a_748_n1036# a_748_n300# a_268_n1036# a_n836_n1036# a_n372_n300#
+ a_n748_n344# a_52_n344# a_n212_436# a_n428_392# a_108_n1036# a_372_n1080# a_n748_n1080#
+ a_108_n300# a_n836_n300# a_n372_436# a_n268_n1080# a_n588_392# a_n372_n1036# a_n532_n300#
+ a_n108_n344# a_212_n344# a_268_n300# a_108_436# a_212_n1080# a_n108_n1080# a_268_436#
+ a_n836_436# a_532_392# a_748_436# a_692_392# a_588_n1036# a_n212_n1036# a_52_392#
+ a_n692_n300# a_n268_n344# a_52_n1080# a_372_n344# a_428_n1036# a_692_n1080# a_428_n300#
+ a_n588_n1080# a_n108_392# a_n268_392# a_n692_n1036# a_n52_n300# a_n428_n344# a_n532_436#
+ a_n692_436# a_n748_392# a_532_n344# a_n52_n1036# a_532_n1080# a_n428_n1080# a_588_n300#
+ a_n52_436# a_n532_n1036# a_212_392# a_n212_n300# a_n588_n344# a_428_436# a_372_392#
+ a_692_n344# a_588_436# VSUBS
X0 a_748_436# a_692_392# a_588_436# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1 a_n52_n1036# a_n108_n1080# a_n212_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X2 a_108_n300# a_52_n344# a_n52_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X3 a_428_n300# a_372_n344# a_268_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X4 a_268_n300# a_212_n344# a_108_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X5 a_268_n1036# a_212_n1080# a_108_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X6 a_108_436# a_52_392# a_n52_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X7 a_n212_n300# a_n268_n344# a_n372_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X8 a_n372_n1036# a_n428_n1080# a_n532_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X9 a_268_436# a_212_392# a_108_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X10 a_n52_n300# a_n108_n344# a_n212_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X11 a_n372_436# a_n428_392# a_n532_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X12 a_428_436# a_372_392# a_268_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X13 a_588_n1036# a_532_n1080# a_428_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X14 a_n212_n1036# a_n268_n1080# a_n372_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X15 a_n692_n1036# a_n748_n1080# a_n836_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X16 a_n532_436# a_n588_392# a_n692_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X17 a_n692_n300# a_n748_n344# a_n836_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X18 a_428_n1036# a_372_n1080# a_268_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X19 a_n532_n1036# a_n588_n1080# a_n692_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X20 a_748_n300# a_692_n344# a_588_n300# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X21 a_108_n1036# a_52_n1080# a_n52_n1036# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X22 a_n52_436# a_n108_392# a_n212_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X23 a_588_n300# a_532_n344# a_428_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X24 a_588_436# a_532_392# a_428_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X25 a_748_n1036# a_692_n1080# a_588_n1036# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X26 a_n532_n300# a_n588_n344# a_n692_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X27 a_n692_436# a_n748_392# a_n836_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X28 a_n212_436# a_n268_392# a_n372_436# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X29 a_n372_n300# a_n428_n344# a_n532_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
.ends

.subckt nmos_3p3_QNHHV5 a_56_n200# a_n56_n244# a_n144_n200# VSUBS
X0 a_56_n200# a_n56_n244# a_n144_n200# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.56u
.ends

.subckt nmos_3p3_4F3WC4 a_n204_336# a_404_n200# a_100_336# a_100_n200# a_n404_292#
+ a_404_n736# a_n404_n244# a_204_n780# a_n492_n200# a_100_n736# a_n100_n244# a_n492_n736#
+ a_n492_336# a_n204_n200# a_n100_292# a_n204_n736# a_n404_n780# a_n100_n780# a_204_292#
+ a_204_n244# a_404_336# VSUBS
X0 a_100_n736# a_n100_n780# a_n204_n736# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1 a_404_336# a_204_292# a_100_336# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X2 a_404_n200# a_204_n244# a_100_n200# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X3 a_100_336# a_n100_292# a_n204_336# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X4 a_100_n200# a_n100_n244# a_n204_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X5 a_n204_336# a_n404_292# a_n492_336# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X6 a_n204_n736# a_n404_n780# a_n492_n736# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X7 a_404_n736# a_204_n780# a_100_n736# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X8 a_n204_n200# a_n404_n244# a_n492_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
.ends

.subckt pmos_3p3_H6V2RY a_n340_68# a_252_68# a_n252_n512# a_n52_68# a_52_24# a_252_n468#
+ a_n252_24# a_n340_n468# a_52_n512# w_n426_n598# a_n52_n468#
X0 a_n52_68# a_n252_24# a_n340_68# w_n426_n598# pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X1 a_252_68# a_52_24# a_n52_68# w_n426_n598# pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X2 a_252_n468# a_52_n512# a_n52_n468# w_n426_n598# pfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X3 a_n52_n468# a_n252_n512# a_n340_n468# w_n426_n598# pfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
.ends

.subckt pmos_3p3_M22VUP a_n164_n344# a_n252_n300# a_52_n344# w_n338_n430# a_n52_n300#
+ a_164_n300#
X0 a_164_n300# a_52_n344# a_n52_n300# w_n338_n430# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.56u
X1 a_n52_n300# a_n164_n344# a_n252_n300# w_n338_n430# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.56u
.ends

.subckt nmos_3p3_5F3WC4 a_n52_n200# a_n52_n736# a_n52_336# a_n252_292# a_n252_n780#
+ a_52_n244# a_252_n200# a_252_n736# a_n252_n244# a_n340_336# a_52_292# a_252_336#
+ a_n340_n200# a_52_n780# a_n340_n736# VSUBS
X0 a_n52_n736# a_n252_n780# a_n340_n736# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X1 a_252_n736# a_52_n780# a_n52_n736# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X2 a_252_n200# a_52_n244# a_n52_n200# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X3 a_n52_n200# a_n252_n244# a_n340_n200# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X4 a_n52_336# a_n252_292# a_n340_336# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X5 a_252_336# a_52_292# a_n52_336# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
.ends

.subckt pmos_3p3_M2JNAR a_n108_n1816# a_108_1172# a_52_1128# a_n196_n1772# a_52_n1816#
+ a_52_n344# a_n196_1172# a_108_n1036# a_108_n300# a_n108_n344# a_n108_1128# a_n196_n300#
+ a_108_436# a_n108_n1080# a_52_392# a_n52_n1772# a_n196_n1036# a_52_n1080# a_n52_1172#
+ a_n108_392# a_n52_n300# a_n52_n1036# a_n52_436# a_n196_436# a_108_n1772# w_n282_n1902#
X0 a_n52_n1036# a_n108_n1080# a_n196_n1036# w_n282_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1 a_108_n1772# a_52_n1816# a_n52_n1772# w_n282_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X2 a_108_n300# a_52_n344# a_n52_n300# w_n282_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X3 a_108_436# a_52_392# a_n52_436# w_n282_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X4 a_n52_n300# a_n108_n344# a_n196_n300# w_n282_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X5 a_n52_n1772# a_n108_n1816# a_n196_n1772# w_n282_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X6 a_108_1172# a_52_1128# a_n52_1172# w_n282_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X7 a_n52_1172# a_n108_1128# a_n196_1172# w_n282_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X8 a_108_n1036# a_52_n1080# a_n52_n1036# w_n282_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X9 a_n52_436# a_n108_392# a_n196_436# w_n282_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt pmos_3p3_MJGNAR a_212_n1816# a_n108_n1816# a_108_1172# a_268_n1036# a_n356_n1036#
+ a_n212_n1772# a_52_1128# a_52_n1816# a_52_n344# a_n212_436# a_108_n1036# a_108_n300#
+ a_268_1172# a_n268_n1080# a_n108_n344# a_n108_1128# a_212_n344# a_212_1128# a_268_n300#
+ a_108_436# a_n356_436# a_212_n1080# a_n108_n1080# a_268_436# a_n356_1172# a_n212_n1036#
+ a_52_392# a_n52_n1772# a_n268_n344# a_n268_1128# a_52_n1080# a_n52_1172# w_n442_n1902#
+ a_n356_n300# a_n108_392# a_n268_392# a_n52_n300# a_n212_1172# a_268_n1772# a_n356_n1772#
+ a_n52_n1036# a_n52_436# a_n268_n1816# a_212_392# a_108_n1772# a_n212_n300#
X0 a_n52_n1036# a_n108_n1080# a_n212_n1036# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1 a_108_n1772# a_52_n1816# a_n52_n1772# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X2 a_108_n300# a_52_n344# a_n52_n300# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X3 a_268_n300# a_212_n344# a_108_n300# w_n442_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X4 a_268_n1036# a_212_n1080# a_108_n1036# w_n442_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X5 a_108_436# a_52_392# a_n52_436# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X6 a_n212_n300# a_n268_n344# a_n356_n300# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X7 a_268_436# a_212_392# a_108_436# w_n442_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X8 a_n52_n300# a_n108_n344# a_n212_n300# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X9 a_n52_n1772# a_n108_n1816# a_n212_n1772# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X10 a_268_n1772# a_212_n1816# a_108_n1772# w_n442_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X11 a_108_1172# a_52_1128# a_n52_1172# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X12 a_n212_n1036# a_n268_n1080# a_n356_n1036# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X13 a_268_1172# a_212_1128# a_108_1172# w_n442_n1902# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X14 a_n212_1172# a_n268_1128# a_n356_1172# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X15 a_n52_1172# a_n108_1128# a_n212_1172# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X16 a_n212_n1772# a_n268_n1816# a_n356_n1772# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X17 a_108_n1036# a_52_n1080# a_n52_n1036# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X18 a_n52_436# a_n108_392# a_n212_436# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X19 a_n212_436# a_n268_392# a_n356_436# w_n442_n1902# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt nmos_3p3_676RTJ a_n372_n300# a_52_n344# a_108_n300# a_n108_n344# a_212_n344#
+ a_268_n300# a_n268_n344# a_372_n344# a_428_n300# a_n52_n300# a_n428_n344# a_n516_n300#
+ a_n212_n300# VSUBS
X0 a_108_n300# a_52_n344# a_n52_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1 a_428_n300# a_372_n344# a_268_n300# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X2 a_268_n300# a_212_n344# a_108_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X3 a_n212_n300# a_n268_n344# a_n372_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X4 a_n52_n300# a_n108_n344# a_n212_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X5 a_n372_n300# a_n428_n344# a_n516_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt ppolyf_u_WRMTN3 a_40_n748# a_n200_n748# a_520_646# a_40_646# a_n440_646# w_n864_n932#
+ a_n200_646# a_520_n748# a_n680_n748# a_280_n748# a_n440_n748# a_280_646# a_n680_646#
X0 a_n680_646# a_n680_n748# w_n864_n932# ppolyf_u r_width=0.8u r_length=6.46u
X1 a_280_646# a_280_n748# w_n864_n932# ppolyf_u r_width=0.8u r_length=6.46u
X2 a_520_646# a_520_n748# w_n864_n932# ppolyf_u r_width=0.8u r_length=6.46u
X3 a_40_646# a_40_n748# w_n864_n932# ppolyf_u r_width=0.8u r_length=6.46u
X4 a_n200_646# a_n200_n748# w_n864_n932# ppolyf_u r_width=0.8u r_length=6.46u
X5 a_n440_646# a_n440_n748# w_n864_n932# ppolyf_u r_width=0.8u r_length=6.46u
.ends

.subckt nmos_3p3_M56RTJ a_n28_392# a_28_n1036# a_n116_n1036# a_n28_n1080# a_n116_436#
+ a_28_n300# a_28_436# a_n28_n344# a_n116_n300# VSUBS
X0 a_28_436# a_n28_392# a_n116_436# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X1 a_28_n300# a_n28_n344# a_n116_n300# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
X2 a_28_n1036# a_n28_n1080# a_n116_n1036# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.28u
.ends

.subckt pmos_3p3_9BLZD7 a_n164_n712# a_n380_n712# a_n268_68# a_n380_760# a_52_n712#
+ a_n468_68# a_n380_n1448# a_n268_804# a_n52_n668# a_n468_n668# a_52_n1448# a_n52_68#
+ a_52_24# a_380_n1404# a_n468_n1404# a_268_n1448# a_164_804# a_n164_n1448# a_164_n1404#
+ a_380_68# a_52_760# a_380_n668# a_164_n668# a_n164_24# a_n164_760# a_n268_n1404#
+ a_268_n712# a_n268_n668# a_n52_804# a_n52_n1404# a_380_804# w_n554_n1534# a_n468_804#
+ a_268_760# a_268_24# a_164_68# a_n380_24#
X0 a_380_804# a_268_760# a_164_804# w_n554_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.56u
X1 a_164_n668# a_52_n712# a_n52_n668# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X2 a_380_n668# a_268_n712# a_164_n668# w_n554_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.56u
X3 a_n268_68# a_n380_24# a_n468_68# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.56u
X4 a_380_n1404# a_268_n1448# a_164_n1404# w_n554_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.56u
X5 a_164_804# a_52_760# a_n52_804# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X6 a_n268_n668# a_n380_n712# a_n468_n668# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.56u
X7 a_n52_804# a_n164_760# a_n268_804# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X8 a_n52_n668# a_n164_n712# a_n268_n668# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X9 a_n268_n1404# a_n380_n1448# a_n468_n1404# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.56u
X10 a_164_68# a_52_24# a_n52_68# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X11 a_n52_68# a_n164_24# a_n268_68# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X12 a_n268_804# a_n380_760# a_n468_804# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.56u
X13 a_380_68# a_268_24# a_164_68# w_n554_n1534# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.56u
X14 a_n52_n1404# a_n164_n1448# a_n268_n1404# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
X15 a_164_n1404# a_52_n1448# a_n52_n1404# w_n554_n1534# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.56u
.ends

.subckt nmos_3p3_N3WVC4 a_n188_n736# a_100_336# a_100_n200# a_100_n736# a_n100_n244#
+ a_n100_292# a_n100_n780# a_n188_336# a_n188_n200# VSUBS
X0 a_100_n736# a_n100_n780# a_n188_n736# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=1u
X1 a_100_336# a_n100_292# a_n188_336# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=1u
X2 a_100_n200# a_n100_n244# a_n188_n200# VSUBS nfet_03v3 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=1u
.ends

.subckt fold_cascode_opamp_mag VDD VSS VINP VINN OUT VC VD VX VA VB VBS2 VBS3 VBIASN
+ IBIAS2 VBIASN2 IBIAS3 IBIAS OUTo VP c_mid
Xpmos_3p3_9K6RD7_9 VB IBIAS VDD VDD pmos_3p3_9K6RD7
Xpmos_3p3_MA2VAR_1 VDD OUT OUT OUT pmos_3p3_MA2VAR
Xpmos_3p3_VK6RD7_3 VDD VBIASN IBIAS VDD pmos_3p3_VK6RD7
Xpmos_3p3_HWZ2RY_2 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD IBIAS2 pmos_3p3_HWZ2RY
Xpmos_3p3_MA2VAR_28 VDD VD VD VD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_3 VX VSS VX VSS VD VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_12 VD VX VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_34 VX VX VX VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_17 VDD VD VD VD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_23 VC VC VC VSS nmos_3p3_M86RTJ
Xpmos_3p3_MAJNAR_0 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ pmos_3p3_MAJNAR
Xpmos_3p3_MA2VAR_2 VDD OUT OUT OUT pmos_3p3_MA2VAR
Xpmos_3p3_VK6RD7_4 VDD VDD VBS2 VBS2 pmos_3p3_VK6RD7
Xnmos_3p3_276RTJ_4 VX VSS VX VSS VC VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_13 VSS VX VD VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_35 VC VBS3 VX VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_24 VD VBS3 OUT VSS nmos_3p3_M86RTJ
Xpmos_3p3_MAJNAR_1 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ pmos_3p3_MAJNAR
Xpmos_3p3_MA2VAR_29 VDD VC VC VC pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_18 VDD VD VINP VP pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_3 VDD OUT VBS2 VB pmos_3p3_MA2VAR
Xpmos_3p3_VK6RD7_5 VDD VBIASN IBIAS VDD pmos_3p3_VK6RD7
Xnmos_3p3_M86RTJ_14 VD VD VD VSS nmos_3p3_M86RTJ
Xnmos_3p3_276RTJ_5 VX VSS VX VSS VC VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_25 OUT OUT OUT VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_36 OUT OUT OUT VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_19 VDD VD VINP VP pmos_3p3_MA2VAR
Xpmos_3p3_MAJNAR_2 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ pmos_3p3_MAJNAR
Xpmos_3p3_MA2VAR_4 VDD OUT OUT OUT pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_15 VD VD VD VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_26 OUT OUT OUT VSS nmos_3p3_M86RTJ
Xnmos_3p3_276RTJ_6 VX VSS VX VSS VD VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_37 OUT VBS3 VD VSS nmos_3p3_M86RTJ
Xpmos_3p3_VK6RD7_6 VDD VDD VDD VDD pmos_3p3_VK6RD7
Xpmos_3p3_MAJNAR_3 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ pmos_3p3_MAJNAR
Xpmos_3p3_MA2VAR_5 VDD VB VBS2 OUT pmos_3p3_MA2VAR
Xpmos_3p3_VK6RD7_7 VDD VDD VDD VDD pmos_3p3_VK6RD7
Xpmos_3p3_VTYQD7_0 VBS3 VDD IBIAS VDD IBIAS VDD pmos_3p3_VTYQD7
Xnmos_3p3_M86RTJ_16 VSS VX VD VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_27 OUT VBS3 VD VSS nmos_3p3_M86RTJ
Xnmos_3p3_276RTJ_7 VX VSS VX VSS VD VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_38 OUT OUT OUT VSS nmos_3p3_M86RTJ
Xpmos_3p3_MAJNAR_4 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ pmos_3p3_MAJNAR
Xpmos_3p3_VTYQD7_1 VBS3 VDD IBIAS VDD IBIAS VDD pmos_3p3_VTYQD7
Xpmos_3p3_MA2VAR_6 VDD OUT OUT OUT pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_17 VD VX VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_276RTJ_8 VBS3 VC VBS3 VC VX VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_28 VX VX VX VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_39 VD VBS3 OUT VSS nmos_3p3_M86RTJ
Xpmos_3p3_MAJNAR_5 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ pmos_3p3_MAJNAR
Xpmos_3p3_MA2VAR_7 VDD OUT VBS2 VB pmos_3p3_MA2VAR
Xcap_mim_2p0fF_XHV85N_0 OUT c_mid cap_mim_2p0fF_XHV85N
Xpmos_3p3_VTYQD7_2 IBIAS VDD IBIAS VDD IBIAS VDD pmos_3p3_VTYQD7
Xnmos_3p3_276RTJ_9 VBS3 VD VBS3 VD OUT VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_29 VC VBS3 VX VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_18 VC VX VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_8 VDD VD VD VD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_19 VC VC VC VSS nmos_3p3_M86RTJ
Xnmos_3p3_NQ5EG7_0 VSS VSS OUTo VSS OUTo OUT OUT VSS OUT VSS OUT OUT VSS VSS OUTo
+ OUT OUT OUTo VSS OUT OUT OUTo VSS OUT OUT OUTo VSS OUT VSS OUT OUTo VSS OUT OUTo
+ OUT OUT OUT VSS OUT VSS OUT OUT OUT OUTo OUTo OUT VSS OUTo OUT OUT OUTo OUT OUT
+ OUTo OUTo VSS OUT VSS OUT VSS OUT OUT OUTo VSS nmos_3p3_NQ5EG7
Xpmos_3p3_MA2VAR_9 VDD VP VINP VD pmos_3p3_MA2VAR
Xnmos_3p3_NQ5EG7_1 VSS VSS OUTo VSS OUTo OUT OUT VSS OUT VSS OUT OUT VSS VSS OUTo
+ OUT OUT OUTo VSS OUT OUT OUTo VSS OUT OUT OUTo VSS OUT VSS OUT OUTo VSS OUT OUTo
+ OUT OUT OUT VSS OUT VSS OUT OUT OUT OUTo OUTo OUT VSS OUTo OUT OUT OUTo OUT OUT
+ OUTo OUTo VSS OUT VSS OUT VSS OUT OUT OUTo VSS nmos_3p3_NQ5EG7
Xnmos_3p3_QNHHV5_0 VSS VBS3 VBS3 VSS nmos_3p3_QNHHV5
Xnmos_3p3_QNHHV5_1 VSS VSS VSS VSS nmos_3p3_QNHHV5
Xnmos_3p3_QNHHV5_2 VBS3 VBS3 VSS VSS nmos_3p3_QNHHV5
Xnmos_3p3_QNHHV5_3 IBIAS2 VBIASN VSS VSS nmos_3p3_QNHHV5
Xnmos_3p3_4F3WC4_0 VSS VSS IBIAS3 IBIAS3 VBIASN2 VSS VBIASN2 VBIASN2 IBIAS3 IBIAS3
+ VBIASN2 IBIAS3 IBIAS3 VSS VBIASN2 VSS VBIASN2 VBIASN2 VBIASN2 VBIASN2 VSS VSS nmos_3p3_4F3WC4
Xnmos_3p3_4F3WC4_1 IBIAS3 IBIAS3 VSS VSS VBIASN2 IBIAS3 VBIASN2 VBIASN2 VSS VSS VBIASN2
+ VSS VSS IBIAS3 VBIASN2 IBIAS3 VBIASN2 VBIASN2 VBIASN2 VBIASN2 IBIAS3 VSS nmos_3p3_4F3WC4
Xpmos_3p3_H6V2RY_0 VDD VDD IBIAS2 VBIASN2 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD VBIASN2
+ pmos_3p3_H6V2RY
Xnmos_3p3_QNHHV5_4 VBS2 VBIASN VSS VSS nmos_3p3_QNHHV5
Xpmos_3p3_M22VUP_0 IBIAS VDD IBIAS VDD VA VDD pmos_3p3_M22VUP
Xpmos_3p3_H6V2RY_1 VDD VDD IBIAS2 VBIASN2 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD VBIASN2
+ pmos_3p3_H6V2RY
Xnmos_3p3_QNHHV5_5 VBIASN VBIASN VSS VSS nmos_3p3_QNHHV5
Xpmos_3p3_M22VUP_1 IBIAS VDD IBIAS VDD VB VDD pmos_3p3_M22VUP
Xnmos_3p3_QNHHV5_6 VSS VBIASN VBS2 VSS nmos_3p3_QNHHV5
Xpmos_3p3_M22VUP_2 IBIAS VDD IBIAS VDD VA VDD pmos_3p3_M22VUP
Xpmos_3p3_M22VUP_3 IBIAS VDD IBIAS VDD VB VDD pmos_3p3_M22VUP
Xnmos_3p3_QNHHV5_8 VSS VSS VSS VSS nmos_3p3_QNHHV5
Xpmos_3p3_M22VAR_0 VBS2 VX VBS2 VX VA VDD pmos_3p3_M22VAR
Xnmos_3p3_5F3WC4_0 VBIASN2 VBIASN2 VBIASN2 VBIASN2 VBIASN2 VBIASN2 VSS VSS VBIASN2
+ VSS VBIASN2 VSS VSS VBIASN2 VSS VSS nmos_3p3_5F3WC4
Xpmos_3p3_M22VAR_1 VBS2 VX VBS2 VX VA VDD pmos_3p3_M22VAR
Xpmos_3p3_M2JNAR_0 IBIAS3 VDD IBIAS3 VDD IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD
+ VDD IBIAS3 IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD
+ pmos_3p3_M2JNAR
Xpmos_3p3_M22VAR_2 VINN VP VINN VP VC VDD pmos_3p3_M22VAR
Xpmos_3p3_M2JNAR_1 IBIAS3 VDD IBIAS3 VDD IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD
+ VDD IBIAS3 IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD
+ pmos_3p3_M2JNAR
Xpmos_3p3_M22VAR_3 VINP VP VINP VP VD VDD pmos_3p3_M22VAR
Xpmos_3p3_M2JNAR_2 IBIAS3 VDD IBIAS3 VDD IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD
+ VDD IBIAS3 IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD
+ pmos_3p3_M2JNAR
Xpmos_3p3_M22VAR_4 VINN VP VINN VP VC VDD pmos_3p3_M22VAR
Xpmos_3p3_MJGNAR_0 IBIAS3 IBIAS3 OUTo VDD VDD OUTo IBIAS3 IBIAS3 IBIAS3 OUTo OUTo
+ OUTo VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD OUTo VDD IBIAS3 IBIAS3 VDD VDD OUTo
+ IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD OUTo VDD VDD VDD VDD
+ IBIAS3 IBIAS3 OUTo OUTo pmos_3p3_MJGNAR
Xnmos_3p3_676RTJ_0 VD VD VSS VD VD VD VD VD VSS VD VD VSS VSS VSS nmos_3p3_676RTJ
Xpmos_3p3_M22VAR_5 VINP VP VINP VP VD VDD pmos_3p3_M22VAR
Xppolyf_u_WRMTN3_0 OUTo OUTo VDD c_mid c_mid VDD c_mid VDD VDD OUTo OUTo c_mid VDD
+ ppolyf_u_WRMTN3
Xpmos_3p3_MJGNAR_1 IBIAS3 IBIAS3 OUTo VDD VDD OUTo IBIAS3 IBIAS3 IBIAS3 OUTo OUTo
+ OUTo VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD OUTo VDD IBIAS3 IBIAS3 VDD VDD OUTo
+ IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD OUTo VDD VDD VDD VDD
+ IBIAS3 IBIAS3 OUTo OUTo pmos_3p3_MJGNAR
Xnmos_3p3_676RTJ_1 VC VC VSS VC VC VC VC VC VSS VC VC VSS VSS VSS nmos_3p3_676RTJ
Xpmos_3p3_M22VAR_6 VINN VP VINN VP VC VDD pmos_3p3_M22VAR
Xpmos_3p3_MJGNAR_2 IBIAS3 IBIAS3 OUTo VDD VDD OUTo IBIAS3 IBIAS3 IBIAS3 OUTo OUTo
+ OUTo VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD OUTo VDD IBIAS3 IBIAS3 VDD VDD OUTo
+ IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD OUTo VDD VDD VDD VDD
+ IBIAS3 IBIAS3 OUTo OUTo pmos_3p3_MJGNAR
Xnmos_3p3_276RTJ_10 VBS3 VD VBS3 VD OUT VSS nmos_3p3_276RTJ
Xpmos_3p3_9K6RD7_20 VP VP VP VDD pmos_3p3_9K6RD7
Xpmos_3p3_M22VAR_7 VINN VP VINN VP VC VDD pmos_3p3_M22VAR
Xpmos_3p3_MJGNAR_3 IBIAS3 IBIAS3 OUTo VDD VDD OUTo IBIAS3 IBIAS3 IBIAS3 OUTo OUTo
+ OUTo VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD OUTo VDD IBIAS3 IBIAS3 VDD VDD OUTo
+ IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD OUTo VDD VDD VDD VDD
+ IBIAS3 IBIAS3 OUTo OUTo pmos_3p3_MJGNAR
Xnmos_3p3_M86RTJ_0 VD VD VD VSS nmos_3p3_M86RTJ
Xnmos_3p3_276RTJ_11 VBS3 VC VBS3 VC VX VSS nmos_3p3_276RTJ
Xpmos_3p3_9K6RD7_10 VA IBIAS VDD VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_21 VP VP VP VDD pmos_3p3_9K6RD7
Xpmos_3p3_M22VAR_8 VINP VP VINP VP VD VDD pmos_3p3_M22VAR
Xpmos_3p3_MJGNAR_4 IBIAS3 IBIAS3 OUTo VDD VDD OUTo IBIAS3 IBIAS3 IBIAS3 OUTo OUTo
+ OUTo VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD OUTo VDD IBIAS3 IBIAS3 VDD VDD OUTo
+ IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD OUTo VDD VDD VDD VDD
+ IBIAS3 IBIAS3 OUTo OUTo pmos_3p3_MJGNAR
Xnmos_3p3_M86RTJ_1 VD VX VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_9K6RD7_0 VB VB VB VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_11 VA VA VA VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_22 VP VP VP VDD pmos_3p3_9K6RD7
Xpmos_3p3_M22VAR_9 VINP VP VINP VP VD VDD pmos_3p3_M22VAR
Xpmos_3p3_MJGNAR_5 IBIAS3 IBIAS3 OUTo VDD VDD OUTo IBIAS3 IBIAS3 IBIAS3 OUTo OUTo
+ OUTo VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD OUTo VDD IBIAS3 IBIAS3 VDD VDD OUTo
+ IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD IBIAS3 IBIAS3 VDD OUTo VDD VDD VDD VDD
+ IBIAS3 IBIAS3 OUTo OUTo pmos_3p3_MJGNAR
Xpmos_3p3_MA2VAR_30 VDD VP VINN VC pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_2 VSS VX VD VSS nmos_3p3_M86RTJ
Xpmos_3p3_9K6RD7_12 VDD IBIAS VB VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_23 VP VP VP VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_1 VA VA VA VDD pmos_3p3_9K6RD7
Xpmos_3p3_MA2VAR_31 VDD VC VINN VP pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_3 VC VX VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_20 VDD VP VINN VC pmos_3p3_MA2VAR
Xpmos_3p3_9K6RD7_13 VB VB VB VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_2 VDD IBIAS VA VDD pmos_3p3_9K6RD7
Xnmos_3p3_M56RTJ_0 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS nmos_3p3_M56RTJ
Xnmos_3p3_M86RTJ_4 VC VC VC VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_21 VDD VC VC VC pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_10 VDD VD VINP VP pmos_3p3_MA2VAR
Xpmos_3p3_9BLZD7_0 IBIAS IBIAS VDD IBIAS IBIAS VP IBIAS VDD VP VP IBIAS VP IBIAS VP
+ VP IBIAS VDD IBIAS VDD VP IBIAS VP VDD IBIAS IBIAS VDD IBIAS VDD VP VP VP VDD VP
+ IBIAS IBIAS VDD IBIAS pmos_3p3_9BLZD7
Xpmos_3p3_9K6RD7_14 VA VA VA VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_3 VB IBIAS VDD VDD pmos_3p3_9K6RD7
Xnmos_3p3_M56RTJ_1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS nmos_3p3_M56RTJ
Xnmos_3p3_M86RTJ_5 VSS VX VC VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_22 VDD VC VINN VP pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_11 VDD VP VINN VC pmos_3p3_MA2VAR
Xnmos_3p3_N3WVC4_0 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS nmos_3p3_N3WVC4
Xpmos_3p3_9K6RD7_15 VDD IBIAS VA VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_4 VA VA VA VDD pmos_3p3_9K6RD7
Xnmos_3p3_M56RTJ_2 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS nmos_3p3_M56RTJ
Xnmos_3p3_M86RTJ_6 VD VX VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_12 VDD VC VC VC pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_23 VDD VD VINP VP pmos_3p3_MA2VAR
Xnmos_3p3_N3WVC4_1 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS nmos_3p3_N3WVC4
Xpmos_3p3_9K6RD7_16 VP VP VP VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_5 VA IBIAS VDD VDD pmos_3p3_9K6RD7
Xnmos_3p3_M56RTJ_3 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS nmos_3p3_M56RTJ
Xnmos_3p3_M86RTJ_7 VSS VX VD VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_30 VX VX VX VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_13 VDD VC VINN VP pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_24 VDD VP VINN VC pmos_3p3_MA2VAR
Xpmos_3p3_9K6RD7_17 VP VP VP VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_6 VB VB VB VDD pmos_3p3_9K6RD7
Xnmos_3p3_276RTJ_0 VX VSS VX VSS VC VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_8 VD VD VD VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_31 VX VBS3 VC VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_20 VSS VX VC VSS nmos_3p3_M86RTJ
Xpmos_3p3_VK6RD7_0 VDD VDD VDD VDD pmos_3p3_VK6RD7
Xpmos_3p3_MA2VAR_14 VDD VP VINP VD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_25 VDD VC VC VC pmos_3p3_MA2VAR
Xpmos_3p3_9K6RD7_7 VDD IBIAS VB VDD pmos_3p3_9K6RD7
Xpmos_3p3_VK6RD7_1 VDD VDD VDD VDD pmos_3p3_VK6RD7
Xpmos_3p3_9K6RD7_18 VP VP VP VDD pmos_3p3_9K6RD7
Xnmos_3p3_276RTJ_1 VX VSS VX VSS VD VSS nmos_3p3_276RTJ
Xpmos_3p3_HWZ2RY_0 VDD VDD VDD VDD VDD VDD VDD pmos_3p3_HWZ2RY
Xpmos_3p3_MA2VAR_26 VDD VC VINN VP pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_9 VC VX VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_10 VC VC VC VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_32 VX VBS3 VC VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_21 VC VX VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_15 VDD VD VD VD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_0 VDD VB VBS2 OUT pmos_3p3_MA2VAR
Xpmos_3p3_9K6RD7_8 VB VB VB VDD pmos_3p3_9K6RD7
Xpmos_3p3_9K6RD7_19 VP VP VP VDD pmos_3p3_9K6RD7
Xpmos_3p3_VK6RD7_2 VDD VDD IBIAS IBIAS pmos_3p3_VK6RD7
Xnmos_3p3_276RTJ_2 VX VSS VX VSS VC VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_11 VSS VX VC VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_33 VX VX VX VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_22 VSS VX VC VSS nmos_3p3_M86RTJ
Xpmos_3p3_HWZ2RY_1 VDD VDD VDD VDD VDD VDD VDD pmos_3p3_HWZ2RY
Xpmos_3p3_MA2VAR_27 VDD VP VINP VD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_16 VDD VP VINP VD pmos_3p3_MA2VAR
.ends

.subckt ppolyf_u_PVCJS8 a_880_700# a_600_700# a_n520_700# a_40_n802# a_320_n802# w_n1264_n986#
+ a_40_700# a_600_n802# a_n1080_700# a_n800_700# a_880_n802# a_n240_n802# a_320_700#
+ a_n520_n802# a_n1080_n802# a_n240_700# a_n800_n802#
X0 a_n520_700# a_n520_n802# w_n1264_n986# ppolyf_u r_width=1u r_length=7u
X1 a_n1080_700# a_n1080_n802# w_n1264_n986# ppolyf_u r_width=1u r_length=7u
X2 a_n800_700# a_n800_n802# w_n1264_n986# ppolyf_u r_width=1u r_length=7u
X3 a_n240_700# a_n240_n802# w_n1264_n986# ppolyf_u r_width=1u r_length=7u
X4 a_40_700# a_40_n802# w_n1264_n986# ppolyf_u r_width=1u r_length=7u
X5 a_600_700# a_600_n802# w_n1264_n986# ppolyf_u r_width=1u r_length=7u
X6 a_880_700# a_880_n802# w_n1264_n986# ppolyf_u r_width=1u r_length=7u
X7 a_320_700# a_320_n802# w_n1264_n986# ppolyf_u r_width=1u r_length=7u
.ends

.subckt VCM_1.6_MAGIC VDD VSS VCM_1.6
Xppolyf_u_PVCJS8_0 VDD m1_1247_1427# VSS m1_689_136# VCM_1.6 VDD m1_1247_1427# VCM_1.6
+ VDD VDD VDD m1_406_n84# m1_966_1668# m1_689_136# VDD m1_966_1668# m1_406_n84# ppolyf_u_PVCJS8
.ends

.subckt nfet_03v3_CT75PZ a_n52_n240# a_152_n240# a_52_n284# a_n152_n284# a_n240_n240#
+ VSUBS
X0 a_n52_n240# a_n152_n284# a_n240_n240# VSUBS nfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.5u
X1 a_152_n240# a_52_n284# a_n52_n240# VSUBS nfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.5u
.ends

.subckt nfet_03v3_CTB5PZ a_50_n240# a_n50_n284# a_n138_n240# VSUBS
X0 a_50_n240# a_n50_n284# a_n138_n240# VSUBS nfet_03v3 ad=1.06p pd=5.68u as=1.06p ps=5.68u w=2.4u l=0.5u
.ends

.subckt BIASING_CURRENT_MAGIC IBIAS_BUF1 IBIAS_BUF2 IBIAS_FILTER IBIAS_PGA G_SINK_UP
+ G_SINK_DOWN VSS
Xnfet_03v3_CT75PZ_1 m1_1867_n835# IBIAS_PGA G_SINK_UP G_SINK_UP IBIAS_PGA VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_0 m1_1867_n835# VSS G_SINK_DOWN G_SINK_DOWN VSS VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_2 m1_214_n835# IBIAS_BUF1 G_SINK_UP G_SINK_UP IBIAS_BUF1 VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_3 m1_214_n835# VSS G_SINK_DOWN G_SINK_DOWN VSS VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_4 m1_765_n835# VSS G_SINK_DOWN G_SINK_DOWN VSS VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_5 m1_765_n835# IBIAS_BUF2 G_SINK_UP G_SINK_UP IBIAS_BUF2 VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_6 m1_1316_n835# VSS G_SINK_DOWN G_SINK_DOWN VSS VSS nfet_03v3_CT75PZ
Xnfet_03v3_CT75PZ_7 m1_1316_n835# IBIAS_FILTER G_SINK_UP G_SINK_UP IBIAS_FILTER VSS
+ nfet_03v3_CT75PZ
Xnfet_03v3_CTB5PZ_0 VSS VSS VSS VSS nfet_03v3_CTB5PZ
Xnfet_03v3_CTB5PZ_1 VSS VSS VSS VSS nfet_03v3_CTB5PZ
Xnfet_03v3_CTB5PZ_2 VSS VSS VSS VSS nfet_03v3_CTB5PZ
Xnfet_03v3_CTB5PZ_3 VSS VSS VSS VSS nfet_03v3_CTB5PZ
.ends

.subckt Folded_Diff_Op_Amp_Layout VDD BD IND IPD VSS VB4 VB2 VB3 VB1 VND VPD IBIAS1
+ VBIASN VOUT VBM VCD IBIAS4 IBIAS3 IBS OUT_P OUT_N IBIAS2 IBIAS VCM IVS IB4 IB2 IB3
+ IB5 IN_P IN_N OUT1 OUT2 m1_29250_n7512# m1_29250_n5500#
Xpmos_3p3_ME7U2H_2 VND VB1 VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_1 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_876RT2_10 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xnmos_3p3_3A6RT2_7 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_4 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_71 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_82 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_93 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_60 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_6 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xnmos_3p3_M86RTJ_67 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_45 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_23 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_15 VDD VB1 VND VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_26 OUT2 VB2 VPD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_12 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_276RTJ_3 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_34 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_106 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_56 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_2F3WC4_1 VSS IVS IVS IVS IVS IVS VSS IVS VSS IVS IVS IVS IVS VSS IVS IVS
+ IVS IVS IVS IVS VSS VSS VSS nmos_3p3_2F3WC4
Xpmos_3p3_MA2VAR_28 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_39 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_17 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_7 VDD VDD VDD ppolyf_u_2VJWHK
Xnmos_3p3_NE3WC4_0 VSS VSS VSS VSS nmos_3p3_NE3WC4
Xnmos_3p3_EA6RT2_0 IB5 VB4 IB5 VB4 VB4 IB5 IB5 IB5 IB5 VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_3 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_2 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_876RT2_11 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xpmos_3p3_5L6RD7_1 VDD IBIAS1 IBIAS1 VDD pmos_3p3_5L6RD7
Xnmos_3p3_3A6RT2_8 VCD VOUT VB1 VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_5 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_50 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_72 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_94 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_61 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_83 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_20 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_S75EG7_0 VB4 VB4 VSS VB4 VB4 VB4 VB4 VSS VB4 VB4 VB4 VSS VB4 VB4 VSS VB4
+ VSS VB4 VB4 VB4 VB4 VSS VB4 VB4 VB4 VB4 VSS VB4 VB4 VSS nmos_3p3_S75EG7
Xpmos_3p3_MNS6FR_7 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_ME7U2H_16 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_276RTJ_4 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_MA2VAR_107 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_68 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_46 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_27 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_13 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_35 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_57 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_24 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_NE3WC4_1 VSS VSS VSS VSS nmos_3p3_NE3WC4
Xpmos_3p3_MA2VAR_29 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_18 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_EA6RT2_1 VCM VCD VCM VCD VCD VBM VBM VCM VCM VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_4 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_3 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_876RT2_0 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_5L6RD7_2 VDD VDD IBIAS1 VBIASN pmos_3p3_5L6RD7
Xnmos_3p3_3A6RT2_9 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_6 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_51 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_40 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_73 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_84 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_95 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_62 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xnmos_3p3_5J7TC4_0 VSS IBS VSS IBIAS IBS VSS nmos_3p3_5J7TC4
Xpmos_3p3_MNS6FR_8 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_MA2VAR_108 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_3A6RT2_21 VBM VCM VCD VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_10 VB1 VOUT VCD VSS nmos_3p3_3A6RT2
Xnmos_3p3_276RTJ_5 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_69 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_47 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_17 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_28 VND VB2 OUT1 VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_36 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_14 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_25 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_58 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_19 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xnmos_3p3_NE3WC4_2 VSS VBIASN IBIAS4 VSS nmos_3p3_NE3WC4
Xnmos_3p3_EA6RT2_2 VOUT VCD VOUT VCD VCD VB1 VB1 VOUT VOUT VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_5 VPD VB1 VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_4 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MYZUAR_0 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xnmos_3p3_876RT2_1 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xnmos_3p3_7WQWW2_7 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_52 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_74 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_9 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_M22VAR_41 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_30 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_85 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_96 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_63 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_5J7TC4_1 VSS IBS VSS IBS IBS VSS nmos_3p3_5J7TC4
Xnmos_3p3_3A6RT2_22 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_11 VCD VCM VBM VSS nmos_3p3_3A6RT2
Xnmos_3p3_276RTJ_6 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_MA2VAR_109 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_ME7U2H_18 VPD VB2 OUT2 VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_29 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_37 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_15 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_26 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_48 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_59 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_EA6RT2_3 VOUT VCD VOUT VCD VCD VB1 VB1 VOUT VOUT VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_6 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_5 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MAEVAR_0 VDD VDD VDD VDD VDD VDD VDD pmos_3p3_MAEVAR
Xpmos_3p3_MYZUAR_1 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xnmos_3p3_876RT2_2 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xnmos_3p3_7WQWW2_8 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_53 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_75 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_20 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_42 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_31 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_86 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_64 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_97 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_23 VCD VOUT VB1 VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_12 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_276RTJ_7 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_16 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_19 OUT2 VB2 VPD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_38 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_49 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_27 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_EA6RT2_4 VCM VCD VCM VCD VCD VBM VBM VCM VCM VSS nmos_3p3_EA6RT2
Xpmos_3p3_ME7U2H_7 VND VB1 VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_6 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MYZUAR_2 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xnmos_3p3_876RT2_3 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xnmos_3p3_7WQWW2_9 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_21 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_54 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_76 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_43 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_10 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_32 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_87 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_65 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_98 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_24 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_13 VB1 VOUT VCD VSS nmos_3p3_3A6RT2
Xnmos_3p3_M86RTJ_17 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_39 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_276RTJ_8 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_28 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_EA6RT2_5 VCM VCD VCM VCD VCD VBM VBM VCM VCM VSS nmos_3p3_EA6RT2
Xpmos_3p3_MES6FR_0 VDD IND BD IN_N pmos_3p3_MES6FR
Xpmos_3p3_MYZUAR_3 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xpmos_3p3_ME7U2H_8 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_7 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_RKK9DS_0 IB2 VB2 VB2 IB2 IB2 VB2 VB2 VB2 VB2 VB2 VB2 VB2 IB2 VB2 VB2 VB2
+ VB2 VB2 VDD VB2 IB2 VB2 IB2 IB2 VB2 VB2 VB2 VB2 VB2 VB2 VB2 IB2 IB2 VB2 pmos_3p3_RKK9DS
Xnmos_3p3_876RT2_4 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_22 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_55 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_77 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_44 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_11 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_33 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_88 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_66 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_99 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_25 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_14 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_276RTJ_9 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_18 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_29 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xcap_mim_2p0fF_3FUNHB_0 OUT_P m1_29250_n5500# cap_mim_2p0fF_3FUNHB
Xnmos_3p3_EA6RT2_6 VOUT VCD VOUT VCD VCD VB1 VB1 VOUT VOUT VSS nmos_3p3_EA6RT2
Xpmos_3p3_5UYQD7_0 VB3 VDD IBIAS1 VDD IBIAS1 VDD pmos_3p3_5UYQD7
Xpmos_3p3_MYZUAR_4 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xpmos_3p3_MES6FR_1 VDD BD IND IN_N pmos_3p3_MES6FR
Xpmos_3p3_ME7U2H_9 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_8 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xnmos_3p3_876RT2_5 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_23 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_78 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_45 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_12 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_34 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_89 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_67 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_56 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_5LZQD7_0 VDD IBIAS1 IBS IBIAS1 IBS IBS VDD IBIAS1 IBIAS1 IBIAS1 VDD VDD
+ pmos_3p3_5LZQD7
Xnmos_3p3_3A6RT2_26 VB1 VOUT VCD VSS nmos_3p3_3A6RT2
Xnmos_3p3_3A6RT2_15 VCD VOUT VB1 VSS nmos_3p3_3A6RT2
Xnmos_3p3_M86RTJ_19 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xcap_mim_2p0fF_3FUNHB_1 OUT_N m1_29250_n7512# cap_mim_2p0fF_3FUNHB
Xpmos_3p3_MES6FR_2 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MA2VAR_9 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MYZUAR_5 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xnmos_3p3_876RT2_6 VCD VBM VCD VCM VCM VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_24 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_79 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_46 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_35 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_13 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_57 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_68 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_5LZQD7_1 VDD IBIAS IBIAS IBIAS IBIAS IBIAS VDD IBIAS IBIAS IBIAS VDD VDD
+ pmos_3p3_5LZQD7
Xnmos_3p3_3A6RT2_16 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_3 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MYZUAR_6 VDD VDD VDD VDD pmos_3p3_MYZUAR
Xpmos_3p3_5C3RD7_0 IBIAS1 VDD VDD VDD IB5 IBIAS1 IBIAS1 IBIAS1 IB5 VDD pmos_3p3_5C3RD7
Xnmos_3p3_876RT2_7 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_HMY8L7_0 VDD BD BD IBIAS VDD VDD BD IBIAS IBIAS BD VDD VDD IBIAS VDD BD
+ VDD IBIAS IBIAS VDD IBIAS VDD IBIAS BD VDD IBIAS VDD IBIAS IBIAS IBIAS VDD IBIAS
+ VDD BD IBIAS IBIAS IBIAS VDD IBIAS IBIAS BD VDD BD IBIAS VDD IBIAS VDD VDD BD BD
+ IBIAS BD BD IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS IBIAS BD IBIAS BD BD
+ IBIAS VDD VDD VDD pmos_3p3_HMY8L7
Xpmos_3p3_M22VAR_25 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_47 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_14 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_36 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_58 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_69 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_17 VBM VCM VCD VSS nmos_3p3_3A6RT2
Xpmos_3p3_K823KY_0 VDD VB2 IB2 VDD pmos_3p3_K823KY
Xpmos_3p3_MES6FR_4 VDD BD IPD IN_P pmos_3p3_MES6FR
Xnmos_3p3_876RT2_8 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_26 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_48 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_15 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_37 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_59 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_18 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_5 VDD IPD BD IN_P pmos_3p3_MES6FR
Xnmos_3p3_JE3WC4_0 VSS IBIAS3 IB4 IBIAS3 VSS IB4 IB4 VSS IBIAS3 IB4 IB4 VSS nmos_3p3_JE3WC4
Xnmos_3p3_U56RT2_0 VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS VSS nmos_3p3_U56RT2
Xpmos_3p3_MNS6FR_10 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xppolyf_u_2V2ZHK_0 m1_26256_n7401# m1_26536_n6269# m1_26256_n7401# VDD m1_25080_n6269#
+ ppolyf_u_2V2ZHK
Xnmos_3p3_876RT2_9 VCD VB1 VCD VOUT VOUT VSS nmos_3p3_876RT2
Xpmos_3p3_M22VAR_27 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_49 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_16 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_38 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_3A6RT2_19 VCD VCM VBM VSS nmos_3p3_3A6RT2
Xnmos_3p3_UUQWW2_0 VB3 OUT1 IND VSS nmos_3p3_UUQWW2
Xpmos_3p3_M2NNAR_0 IBIAS4 IBIAS4 VDD IB4 IBIAS4 IB4 IBIAS4 IBIAS4 VDD VDD VDD IBIAS4
+ VDD IBIAS4 VDD IB4 IB4 VDD VDD IBIAS4 VDD pmos_3p3_M2NNAR
Xpmos_3p3_MES6FR_6 VDD IND BD IN_N pmos_3p3_MES6FR
Xnmos_3p3_JE3WC4_1 IB4 VSS IB4 VSS IB4 IB4 IB4 IB4 VSS IB4 IB4 VSS nmos_3p3_JE3WC4
Xpmos_3p3_MNS6FR_11 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xppolyf_u_2V2ZHK_1 m1_24352_n7688# m1_24072_n6269# OUT_N VDD m1_24072_n6269# ppolyf_u_2V2ZHK
Xpmos_3p3_M22VAR_17 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_39 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_28 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_UUQWW2_1 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_M2NNAR_1 IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD VDD VDD
+ IBIAS3 VDD IBIAS3 VDD IBIAS3 IBIAS3 VDD VDD IBIAS3 VDD pmos_3p3_M2NNAR
Xpmos_3p3_MES6FR_7 VDD BD IND IN_N pmos_3p3_MES6FR
Xpmos_3p3_MNS6FR_12 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xppolyf_u_2V2ZHK_2 m1_24800_n7401# m1_25080_n6269# m1_24800_n7401# VDD m1_23624_n6269#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_M22VAR_18 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_29 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_UUQWW2_2 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MES6FR_8 VDD IND BD IN_N pmos_3p3_MES6FR
Xpmos_3p3_MNS6FR_13 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xppolyf_u_2V2ZHK_3 m1_25808_n7688# m1_25528_n6269# m1_24352_n7688# VDD m1_25528_n6269#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_M22VAR_19 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_UUQWW2_3 VB3 IND OUT1 VSS nmos_3p3_UUQWW2
Xpmos_3p3_MQ2VAR_0 VBM VDD VBM VDD VBM VDD pmos_3p3_MQ2VAR
Xpmos_3p3_MES6FR_9 VDD BD IND IN_N pmos_3p3_MES6FR
Xpmos_3p3_MNS6FR_14 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xppolyf_u_2V2ZHK_4 m1_26536_n5429# m1_26256_n4297# m1_25080_n5716# VDD m1_26256_n4297#
+ ppolyf_u_2V2ZHK
Xnmos_3p3_UUQWW2_40 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MQ2VAR_1 VB1 VDD VB1 VDD VB1 VDD pmos_3p3_MQ2VAR
Xnmos_3p3_UUQWW2_4 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_M22VAR_190 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_15 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xppolyf_u_2V2ZHK_5 m1_25528_n5429# m1_25808_n4297# m1_25528_n5429# VDD m1_24352_n4297#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_MN7U2H_20 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_41 VB4 VSS IPD VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_30 VB4 IPD VSS VSS nmos_3p3_UUQWW2
Xppolyf_u_RRG95T_0 m1_29250_n7512# m1_29250_n7512# OUT1 OUT1 VDD OUT1 m1_29250_n7512#
+ m1_29250_n7512# OUT1 ppolyf_u_RRG95T
Xnmos_3p3_UUQWW2_5 VB3 IND OUT1 VSS nmos_3p3_UUQWW2
Xpmos_3p3_M22VAR_191 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_180 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_FSHHD6_0 VBIASN VSS VBIASN VSS VBIASN VSS nmos_3p3_FSHHD6
Xpmos_3p3_MNS6FR_16 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xppolyf_u_2V2ZHK_6 m1_25080_n5716# m1_24800_n4297# m1_23624_n5716# VDD m1_24800_n4297#
+ ppolyf_u_2V2ZHK
Xpmos_3p3_MN7U2H_21 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xpmos_3p3_MN7U2H_10 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_42 VB4 IPD VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_31 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_V56RT2_0 VB3 IB3 IB3 IB3 VB3 VB3 VB3 VB3 VB3 VB3 IB3 VB3 VB3 VB3 VB3 VSS
+ nmos_3p3_V56RT2
Xppolyf_u_RRG95T_1 m1_29250_n5500# m1_29250_n5500# OUT2 OUT2 VDD OUT2 m1_29250_n5500#
+ m1_29250_n5500# OUT2 ppolyf_u_RRG95T
Xnmos_3p3_UUQWW2_20 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_6 VB3 OUT1 IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_30 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_170 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_192 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_181 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_17 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xppolyf_u_2V2ZHK_7 m1_24072_n5429# m1_24352_n4297# m1_24072_n5429# VDD VOUT ppolyf_u_2V2ZHK
Xpmos_3p3_M22VAR_0 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_22 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xpmos_3p3_MN7U2H_11 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_43 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_32 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_21 VB4 IND VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_10 VB3 IPD OUT2 VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_7 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_31 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_20 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_171 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_193 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_182 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_160 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_1 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_12 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xpmos_3p3_MN7U2H_23 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_44 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_22 VB4 VSS IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_33 VB4 VSS IPD VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_8 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_11 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_32 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_21 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_10 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_161 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_172 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_150 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_194 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_183 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_2 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_13 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_45 VB4 VSS IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_23 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_12 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_34 VB4 IPD VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_9 VB3 OUT2 IPD VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_33 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_22 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_11 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_162 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_173 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_140 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_151 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_HDY8L7_0 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pmos_3p3_HDY8L7
Xpmos_3p3_M22VAR_195 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_184 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_50 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_Q3NTJU_0 VDD VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD VDD IBIAS3 IBIAS3 IBIAS3
+ IBIAS3 IBIAS3 VDD IVS IVS VDD IBIAS3 IBIAS3 IBIAS3 VDD IBIAS3 IVS VDD VDD IVS IBIAS3
+ IBIAS3 IVS VDD IVS IBIAS3 IBIAS3 IVS IVS IVS IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3
+ VDD IBIAS3 IBIAS3 IVS IBIAS3 VDD IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 VDD IVS IBIAS3
+ IBIAS3 VDD IBIAS3 IBIAS3 IBIAS3 IBIAS3 IBIAS3 VDD IBIAS3 IBIAS3 IVS IVS IVS VDD
+ IVS IBIAS3 IVS IBIAS3 IBIAS3 VDD VDD VDD IVS IBIAS3 IBIAS3 IVS IVS IBIAS3 IVS IVS
+ IBIAS3 VDD IVS VDD VDD VDD IBIAS3 VDD IBIAS3 VDD IVS VDD IBIAS3 IBIAS3 IVS IVS IBIAS3
+ IBIAS3 VDD VDD IBIAS3 IBIAS3 IBIAS3 VDD VDD IBIAS3 IVS IVS VDD IBIAS3 IVS pmos_3p3_Q3NTJU
Xpmos_3p3_M22VAR_3 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_14 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_46 VB4 IND VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_24 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_35 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_13 VB3 OUT2 IPD VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_34 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_23 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_12 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_163 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_174 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_141 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_152 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_130 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_HDY8L7_1 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pmos_3p3_HDY8L7
Xpmos_3p3_M22VAR_185 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_90 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_51 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_40 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_QNHHD6_0 VSS VBIASN VB2 VSS nmos_3p3_QNHHD6
Xpmos_3p3_M22VAR_4 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_15 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_47 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_36 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_25 VB4 VSS IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_14 VB3 IPD OUT2 VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_0 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_35 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_13 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_24 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_164 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_142 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_120 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_153 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_131 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_175 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_91 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_80 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_186 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_52 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_30 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_41 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_M22VAR_5 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MN7U2H_16 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_37 VB4 VSS IND VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_26 VB4 IND VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_1 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_15 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_14 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_25 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_110 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_165 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_92 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_70 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_143 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_121 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_132 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_187 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_176 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_81 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_154 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_53 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_31 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_20 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_42 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_M22VAR_6 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MES6FR_20 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MN7U2H_17 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_16 VB4 VSS IPD VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_2 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_38 VB4 IND VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_27 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_7WQWW2_15 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_26 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_111 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_60 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_133 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_166 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_100 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_144 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_71 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_122 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_82 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_188 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_93 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_177 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_155 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_32 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_21 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_10 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_43 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpfet_03v3_6DHECV_0 VDD VDD VDD VDD pfet_03v3_6DHECV
Xpmos_3p3_M22VAR_7 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_6F3WC4_0 VSS VSS VSS VSS VSS VSS VSS nmos_3p3_6F3WC4
Xpmos_3p3_MES6FR_10 VDD BD IPD IN_P pmos_3p3_MES6FR
Xpmos_3p3_MES6FR_21 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MN7U2H_18 OUT1 VDD VB2 VND VB2 VND pmos_3p3_MN7U2H
Xppolyf_u_RKG95T_0 VDD VDD VDD ppolyf_u_RKG95T
Xnmos_3p3_UUQWW2_39 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_28 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xnmos_3p3_UUQWW2_17 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_3 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_27 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_16 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_M86RTJ_0 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_61 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_134 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_167 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_50 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_101 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_112 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_145 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_123 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_72 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_94 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_189 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_83 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_178 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_156 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_33 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_22 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_11 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_44 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_M22VAR_8 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_6F3WC4_1 VSS VSS VSS VSS VSS VSS VSS nmos_3p3_6F3WC4
Xpmos_3p3_MES6FR_11 VDD IPD BD IN_P pmos_3p3_MES6FR
Xpmos_3p3_MES6FR_22 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MN7U2H_19 OUT2 VDD VB2 VPD VB2 VPD pmos_3p3_MN7U2H
Xnmos_3p3_UUQWW2_29 VB4 VSS IPD VSS nmos_3p3_UUQWW2
Xppolyf_u_RKG95T_1 VDD VDD VDD ppolyf_u_RKG95T
Xnmos_3p3_UUQWW2_18 VSS VSS VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_4 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_28 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_17 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_M86RTJ_1 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_40 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_135 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_168 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_102 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_113 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_146 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_124 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_179 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_157 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_62 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_51 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_73 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_84 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_95 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_12 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_34 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_23 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_45 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_BSHHD6_0 VSS VBIASN VBIASN VCD VBIASN VSS VSS VCD VBIASN VBIASN VBIASN VSS
+ VCD VSS nmos_3p3_BSHHD6
Xpmos_3p3_M22VAR_9 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xnmos_3p3_6F3WC4_2 VSS VSS VSS VSS VSS VSS VSS nmos_3p3_6F3WC4
Xpmos_3p3_MES6FR_23 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MES6FR_12 VDD IND BD IN_N pmos_3p3_MES6FR
Xppolyf_u_RKG95T_2 VDD VDD VDD ppolyf_u_RKG95T
Xnmos_3p3_UUQWW2_19 VB4 IPD VSS VSS nmos_3p3_UUQWW2
Xpmos_3p3_MN7U2H_5 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_7WQWW2_29 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_7WQWW2_18 VSS VSS VB4 IPD VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_M86RTJ_2 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_M22VAR_136 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_169 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_103 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_114 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_125 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_147 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_158 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_30 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_41 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_63 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_96 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_52 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_85 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_74 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_13 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_35 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_24 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_46 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xpmos_3p3_MES6FR_13 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MANNAR_0 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pmos_3p3_MANNAR
Xppolyf_u_RKG95T_3 VDD VDD VDD ppolyf_u_RKG95T
Xpmos_3p3_MN7U2H_6 VPD VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_M86RTJ_70 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_7WQWW2_19 VSS VSS VB4 IND VB4 VSS nmos_3p3_7WQWW2
Xnmos_3p3_M86RTJ_3 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_31 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_137 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_97 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_20 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_42 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_104 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_53 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_64 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_115 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_86 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_75 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_148 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_126 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_159 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xnmos_3p3_276RTJ_14 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_25 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_47 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_36 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_3A6RT2_0 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_14 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MANNAR_1 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pmos_3p3_MANNAR
Xpmos_3p3_MN7U2H_7 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xpmos_3p3_MEKUKR_0 VDD VDD IBIAS4 IBIAS4 pmos_3p3_MEKUKR
Xnmos_3p3_M86RTJ_71 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_30 OUT1 VB2 VND VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_60 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_110 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_4 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_M22VAR_105 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_138 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_76 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_98 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_10 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_21 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_43 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_54 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_32 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_116 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_65 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_149 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_127 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xppolyf_u_2VJWHK_0 m1_23624_n6269# OUT_P VDD ppolyf_u_2VJWHK
Xpmos_3p3_MA2VAR_87 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_48 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_15 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_26 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_37 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_3A6RT2_1 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_15 VDD VDD VDD VDD pmos_3p3_MES6FR
Xpmos_3p3_MNS6FR_0 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_MN7U2H_8 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xpmos_3p3_MA2VAR_111 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MEKUKR_1 VDD VDD IBIAS4 IBIAS4 pmos_3p3_MEKUKR
Xpmos_3p3_ME7U2H_20 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_31 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_50 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_61 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_100 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_5 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_M22VAR_106 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_139 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_77 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_11 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_22 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_55 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_33 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_44 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_117 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_88 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_66 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_128 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xppolyf_u_2VJWHK_1 VDD VDD VDD ppolyf_u_2VJWHK
Xpmos_3p3_MA2VAR_99 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_49 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_16 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_27 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_38 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_3AEFT2_0 IB3 VB3 VSS VSS nmos_3p3_3AEFT2
Xpmos_3p3_MES6FR_16 VDD VDD VDD VDD pmos_3p3_MES6FR
Xnmos_3p3_3A6RT2_2 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xpmos_3p3_MNS6FR_1 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xpmos_3p3_MN7U2H_9 VND VDD VB1 VDD VB1 VDD pmos_3p3_MN7U2H
Xnmos_3p3_M86RTJ_40 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_21 VND VB2 OUT1 VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_10 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_51 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_62 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_101 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_6 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_12 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_107 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_23 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_34 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_45 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_56 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_118 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_129 IBIAS2 VDD IBIAS2 VDD IBIAS2 VDD pmos_3p3_M22VAR
Xppolyf_u_2VJWHK_2 m1_25808_n4297# m1_26536_n6269# VDD ppolyf_u_2VJWHK
Xpmos_3p3_MA2VAR_78 VDD VDD IBIAS2 OUT_N pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_89 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_67 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_17 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_28 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_39 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_MES6FR_17 VDD VDD VDD VDD pmos_3p3_MES6FR
Xnmos_3p3_3A6RT2_3 VCD VCM VBM VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_0 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_MNS6FR_2 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xpmos_3p3_ME7U2H_11 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_102 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_41 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_22 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_7 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_63 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_30 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_52 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_M22VAR_108 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_119 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xppolyf_u_2VJWHK_3 VOUT m1_23624_n5716# VDD ppolyf_u_2VJWHK
Xpmos_3p3_MA2VAR_13 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_79 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_24 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_35 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_46 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_57 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_68 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xnmos_3p3_276RTJ_29 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_276RTJ_18 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_M82RNG_0 VDD VDD VDD VDD pmos_3p3_M82RNG
Xnmos_3p3_3A6RT2_4 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_18 VDD BD IND IN_N pmos_3p3_MES6FR
Xnmos_3p3_7WQWW2_1 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_90 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_3 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xnmos_3p3_276RTJ_0 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_MA2VAR_103 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_64 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_42 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_20 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_23 OUT1 VB2 VND VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_8 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_12 VDD VB1 VND VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_31 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_53 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_14 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_M22VAR_109 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MA2VAR_25 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_36 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_47 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_58 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_69 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_4 m1_26536_n5429# m1_25808_n7688# VDD ppolyf_u_2VJWHK
Xnmos_3p3_276RTJ_19 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xpmos_3p3_ME7U2H_0 VPD VB1 VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_M82RNG_1 VDD VDD VDD VDD pmos_3p3_M82RNG
Xnmos_3p3_3A6RT2_5 VBM VCM VCD VSS nmos_3p3_3A6RT2
Xpmos_3p3_MES6FR_19 VDD VDD VDD VDD pmos_3p3_MES6FR
Xnmos_3p3_7WQWW2_2 OUT1 OUT1 VB3 IND VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_80 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_91 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_4 VDD BD BD IN_N IN_N IND pmos_3p3_MNS6FR
Xnmos_3p3_276RTJ_1 OUT2 VSS OUT2 VSS OUT_P VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_43 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_65 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_21 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xpmos_3p3_ME7U2H_24 VPD VB2 OUT2 VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_13 VDD VB1 VPD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_10 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_32 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_54 VSS OUT1 OUT_N VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_104 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_9 VSS OUT2 OUT_P VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_15 VDD OUT_N IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_26 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_37 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_48 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_59 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_5 VDD VDD VDD ppolyf_u_2VJWHK
Xpmos_3p3_ME7U2H_1 VDD VB1 VPD VDD pmos_3p3_ME7U2H
Xpmos_3p3_MA2VAR_0 VDD VDD IBIAS2 OUT_P pmos_3p3_MA2VAR
Xnmos_3p3_3A6RT2_6 VSS VSS VSS VSS nmos_3p3_3A6RT2
Xnmos_3p3_7WQWW2_3 OUT2 OUT2 VB3 IPD VB3 VSS nmos_3p3_7WQWW2
Xpmos_3p3_M22VAR_70 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_81 IBIAS2 VDD IBIAS2 VDD OUT_N VDD pmos_3p3_M22VAR
Xpmos_3p3_M22VAR_92 IBIAS2 VDD IBIAS2 VDD OUT_P VDD pmos_3p3_M22VAR
Xpmos_3p3_MNS6FR_5 VDD BD BD IN_P IN_P IPD pmos_3p3_MNS6FR
Xnmos_3p3_276RTJ_2 OUT1 VSS OUT1 VSS OUT_N VSS nmos_3p3_276RTJ
Xnmos_3p3_M86RTJ_66 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_44 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_22 OUT_P OUT2 VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_2F3WC4_0 IBIAS2 VSS IVS IVS VSS IVS IBIAS2 IVS IBIAS2 VSS IVS IVS VSS IBIAS2
+ IVS IVS IVS IVS VSS VSS IBIAS2 IBIAS2 VSS nmos_3p3_2F3WC4
Xpmos_3p3_ME7U2H_25 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xpmos_3p3_ME7U2H_14 VDD VDD VDD VDD pmos_3p3_ME7U2H
Xnmos_3p3_M86RTJ_11 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xnmos_3p3_M86RTJ_33 VSS VSS VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_105 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xnmos_3p3_M86RTJ_55 OUT_N OUT1 VSS VSS nmos_3p3_M86RTJ
Xpmos_3p3_MA2VAR_38 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_27 VDD OUT_P IBIAS2 VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_16 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xpmos_3p3_MA2VAR_49 VDD VDD VDD VDD pmos_3p3_MA2VAR
Xppolyf_u_2VJWHK_6 VDD VDD VDD ppolyf_u_2VJWHK
.ends

.subckt cap_mim_2p0fF_NEQE26 m4_n1840_n3340# m4_n1720_n3220#
X0 m4_n1720_n3220# m4_n1840_n3340# cap_mim_2f0_m4m5_noshield c_width=16u c_length=15.2u
X1 m4_n1720_n3220# m4_n1840_n3340# cap_mim_2f0_m4m5_noshield c_width=16u c_length=15.2u
.ends

.subckt ppolyf_u_6V6NLJ a_n520_n332# a_1160_n332# a_320_230# a_n1080_n332# a_n240_230#
+ a_1440_230# a_n800_n332# w_n1824_n516# a_1440_n332# a_n1360_n332# a_n1360_230# a_n1640_n332#
+ a_880_230# a_600_230# a_n520_230# a_40_n332# a_n1640_230# a_320_n332# a_1160_230#
+ a_40_230# a_600_n332# a_n1080_230# a_880_n332# a_n240_n332# a_n800_230#
X0 a_n1640_230# a_n1640_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X1 a_n1360_230# a_n1360_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X2 a_n520_230# a_n520_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X3 a_n1080_230# a_n1080_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X4 a_n800_230# a_n800_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X5 a_n240_230# a_n240_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X6 a_1440_230# a_1440_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X7 a_40_230# a_40_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X8 a_1160_230# a_1160_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X9 a_600_230# a_600_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X10 a_880_230# a_880_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
X11 a_320_230# a_320_n332# w_n1824_n516# ppolyf_u r_width=1u r_length=2.3u
.ends

.subckt filter_res_magic R7_R8_R10_C R3_R7 INN_P VDD OP_AMP_IN_P OP_AMP_IN_N m1_387_n1103#
+ m1_2627_n3434# m1_387_n186# m1_387_n4916# m1_387_731#
Xcap_mim_2p0fF_NEQE26_0 OP_AMP_IN_N m1_387_n4916# cap_mim_2p0fF_NEQE26
Xcap_mim_2p0fF_NEQE26_1 R3_R7 m1_387_n186# cap_mim_2p0fF_NEQE26
Xcap_mim_2p0fF_NEQE26_2 OP_AMP_IN_P m1_387_731# cap_mim_2p0fF_NEQE26
Xcap_mim_2p0fF_NEQE26_3 R3_R7 m1_387_n186# cap_mim_2p0fF_NEQE26
Xcap_mim_2p0fF_NEQE26_4 R3_R7 m1_387_n186# cap_mim_2p0fF_NEQE26
Xcap_mim_2p0fF_NEQE26_5 m1_387_n1103# R7_R8_R10_C cap_mim_2p0fF_NEQE26
Xppolyf_u_6V6NLJ_1 m1_767_n4438# m1_2067_n3999# m1_2167_n5030# m1_767_n4438# m1_1047_n5030#
+ VDD m1_486_n4324# VDD VDD m1_486_n4324# m1_387_n4916# VDD m1_2167_n5030# m1_2446_n4916#
+ m1_1326_n4916# m1_1887_n4438# VDD m1_1607_n4324# m1_2446_n4916# m1_1326_n4916# m1_1887_n4438#
+ R3_R7 m1_2704_n4323# m1_1607_n4324# m1_1047_n5030# ppolyf_u_6V6NLJ
Xppolyf_u_6V6NLJ_0 m1_946_n2582# OP_AMP_IN_N m1_1789_n3097# m1_384_n2588# m1_1227_n3094#
+ VDD m1_946_n2582# VDD VDD m1_384_n2588# R7_R8_R10_C VDD OP_AMP_IN_N OP_AMP_IN_N
+ m1_1227_n3094# m1_1506_n2582# VDD m1_2066_n2585# OP_AMP_IN_N m1_1789_n3097# m1_2066_n2585#
+ m1_667_n3094# OP_AMP_IN_N m1_1506_n2582# m1_667_n3094# ppolyf_u_6V6NLJ
Xppolyf_u_6V6NLJ_2 m1_1327_n3521# m1_2447_n3407# m1_2067_n3999# R7_R8_R10_C m1_1607_n3999#
+ VDD m1_1047_n3636# VDD VDD m1_488_n3407# R3_R7 VDD m1_1607_n3999# m1_1887_n4113#
+ m1_767_n4113# m1_1327_n3521# VDD m1_1047_n3636# m1_2704_n4323# m1_1887_n4113# m1_2447_n3407#
+ m1_767_n4113# m1_2627_n3434# m1_488_n3407# R7_R8_R10_C ppolyf_u_6V6NLJ
Xppolyf_u_6V6NLJ_3 m1_945_n1681# OP_AMP_IN_P m1_1783_n1186# m1_387_n1682# m1_1225_n1159#
+ VDD m1_945_n1681# VDD VDD m1_387_n1682# m1_387_n1103# VDD OP_AMP_IN_P OP_AMP_IN_P
+ m1_1225_n1159# m1_1506_n1677# VDD m1_2064_n1679# OP_AMP_IN_P m1_1783_n1186# m1_2064_n1679#
+ m1_665_n1170# OP_AMP_IN_P m1_1506_n1677# m1_665_n1170# ppolyf_u_6V6NLJ
Xppolyf_u_6V6NLJ_4 m1_767_166# m1_2067_n186# m1_2167_758# m1_767_166# m1_1047_758#
+ VDD m1_486_52# VDD VDD m1_486_52# m1_387_731# VDD m1_2167_758# m1_2446_644# m1_1326_644#
+ m1_1887_166# VDD m1_1607_52# m1_2446_644# m1_1326_644# m1_1887_166# m1_387_n186#
+ m1_2704_51# m1_1607_52# m1_1047_758# ppolyf_u_6V6NLJ
Xppolyf_u_6V6NLJ_5 m1_1327_n751# m1_2447_n865# m1_2067_n186# m1_387_n1103# m1_1607_n300#
+ VDD m1_1047_n751# VDD VDD m1_488_n865# m1_387_n186# VDD m1_1607_n300# m1_1887_n159#
+ m1_767_n159# m1_1327_n751# VDD m1_1047_n751# m1_2704_51# m1_1887_n159# m1_2447_n865#
+ m1_767_n159# INN_P m1_488_n865# m1_387_n1103# ppolyf_u_6V6NLJ
.ends

.subckt Filter_magic VIN_N1 VOUT_N VDD VSS VOUT_OPAMP_P VOUT_OPAMP_N VIN_P1 R3_R7_1
+ R7_R8_R10_C1 IB21 IBIAS11 VBM1 VBIASN1 IB31 IBS1 VB21 VB31 VB41 VCD1 IND1 IPD1 OUT2_1
+ OUT1_1 IBIAS3_1 IB4_1 IBIAS4_1 IVS_1 IBIAS2_1 VB1_1 BD_1 R_1 R11_1 OPAMP_C_1 OPAMP_C1_1
+ VOUT_1_1 VOUT_P VCM1
XFolded_Diff_Op_Amp_Layout_0 VDD BD_1 IND1 IPD1 VSS VB41 VB21 VB31 VB1_1 Folded_Diff_Op_Amp_Layout_0/VND
+ Folded_Diff_Op_Amp_Layout_0/VPD IBIAS11 VBIASN1 VOUT_1_1 VBM1 VCD1 IBIAS4_1 IBIAS3_1
+ IBS1 VOUT_P VOUT_N IBIAS2_1 Folded_Diff_Op_Amp_Layout_0/IBIAS VCM1 IVS_1 IB4_1 IB21
+ IB31 Folded_Diff_Op_Amp_Layout_0/IB5 VOUT_OPAMP_P VOUT_OPAMP_N OUT1_1 OUT2_1 OPAMP_C_1
+ OPAMP_C1_1 Folded_Diff_Op_Amp_Layout
Xfilter_res_magic_0 R7_R8_R10_C1 R3_R7_1 VIN_P1 VDD VOUT_OPAMP_P VOUT_OPAMP_N R_1
+ VIN_N1 R11_1 VOUT_P VOUT_N filter_res_magic
.ends

.subckt ppolyf_u_S2N82J a_1160_n492# a_320_390# a_n520_n492# w_n1544_n676# a_n1080_n492#
+ a_n240_390# a_n800_n492# a_n1360_n492# a_n1360_390# a_880_390# a_600_390# a_n520_390#
+ a_40_n492# a_320_n492# a_1160_390# a_40_390# a_600_n492# a_n1080_390# a_880_n492#
+ a_n240_n492# a_n800_390#
X0 a_n1360_390# a_n1360_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X1 a_n520_390# a_n520_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X2 a_n1080_390# a_n1080_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X3 a_n800_390# a_n800_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X4 a_n240_390# a_n240_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X5 a_40_390# a_40_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X6 a_1160_390# a_1160_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X7 a_600_390# a_600_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X8 a_320_390# a_320_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
X9 a_880_390# a_880_n492# w_n1544_n676# ppolyf_u r_width=1u r_length=3.9u
.ends

.subckt x200_ohm_magic R1_IN R2_IN COMMON VDD
Xppolyf_u_S2N82J_0 VDD COMMON R2_IN VDD R2_IN COMMON R1_IN VDD VDD COMMON COMMON COMMON
+ R2_IN R1_IN VDD COMMON R2_IN COMMON R1_IN R1_IN COMMON ppolyf_u_S2N82J
Xppolyf_u_S2N82J_1 VDD R2_IN COMMON VDD COMMON R2_IN COMMON VDD VDD R2_IN R1_IN R1_IN
+ COMMON COMMON VDD R1_IN COMMON R1_IN COMMON COMMON R2_IN ppolyf_u_S2N82J
.ends

.subckt pfet_03v3_GKYWHF a_n1100_n1036# a_n404_n1080# a_n100_n344# a_1012_n1036# a_n508_n1036#
+ a_n508_n300# a_n1012_n344# a_n812_436# a_1012_n300# a_n1100_n300# a_n204_n300# a_508_392#
+ a_812_n1080# a_n708_n1080# a_n1012_n1080# a_n100_392# a_n1012_392# a_n812_n1036#
+ a_708_436# a_n812_n300# a_204_392# a_n508_436# a_508_n344# a_204_n344# a_404_436#
+ a_n708_392# a_100_n1036# a_708_n300# a_n204_436# a_204_n1080# a_812_392# a_404_n1036#
+ w_n1186_n1166# a_n100_n1080# a_404_n300# a_n708_n344# a_n204_n1036# a_100_n300#
+ a_812_n344# a_100_436# a_n1100_436# a_n404_392# a_n404_n344# a_1012_436# a_508_n1080#
+ a_708_n1036#
X0 a_n508_436# a_n708_392# a_n812_436# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X1 a_100_n300# a_n100_n344# a_n204_n300# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X2 a_708_n300# a_508_n344# a_404_n300# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X3 a_n204_436# a_n404_392# a_n508_436# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X4 a_708_n1036# a_508_n1080# a_404_n1036# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X5 a_n812_n300# a_n1012_n344# a_n1100_n300# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=1u
X6 a_1012_436# a_812_392# a_708_436# w_n1186_n1166# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=1u
X7 a_n508_n1036# a_n708_n1080# a_n812_n1036# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X8 a_n204_n300# a_n404_n344# a_n508_n300# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X9 a_100_n1036# a_n100_n1080# a_n204_n1036# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X10 a_1012_n1036# a_812_n1080# a_708_n1036# w_n1186_n1166# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=1u
X11 a_1012_n300# a_812_n344# a_708_n300# w_n1186_n1166# pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=1u
X12 a_n812_436# a_n1012_392# a_n1100_436# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=1u
X13 a_708_436# a_508_392# a_404_436# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X14 a_n812_n1036# a_n1012_n1080# a_n1100_n1036# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=1u
X15 a_n508_n300# a_n708_n344# a_n812_n300# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X16 a_404_n1036# a_204_n1080# a_100_n1036# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X17 a_404_436# a_204_392# a_100_436# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X18 a_404_n300# a_204_n344# a_100_n300# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X19 a_n204_n1036# a_n404_n1080# a_n508_n1036# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
X20 a_100_436# a_n100_392# a_n204_436# w_n1186_n1166# pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=1u
.ends

.subckt pfet_03v3_GKYJHF a_n100_n344# a_n100_392# w_n274_n1166# a_n188_436# a_n188_n300#
+ a_100_n1036# a_n100_n1080# a_n188_n1036# a_100_n300# a_100_436#
X0 a_100_n300# a_n100_n344# a_n188_n300# w_n274_n1166# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=1u
X1 a_100_n1036# a_n100_n1080# a_n188_n1036# w_n274_n1166# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=1u
X2 a_100_436# a_n100_392# a_n188_436# w_n274_n1166# pfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=1u
.ends

.subckt nfet_03v3_U5DXAV a_458_n300# a_358_n344# a_662_n300# a_n458_n344# a_562_n344#
+ a_n662_n344# a_254_n300# a_n766_n300# a_154_n344# a_n970_n300# a_n1158_n300# a_n254_n344#
+ a_n358_n300# a_n562_n300# a_50_n300# a_866_n300# a_766_n344# a_n1070_n344# a_n50_n344#
+ a_n866_n344# a_1070_n300# a_n154_n300# a_970_n344# VSUBS
X0 a_n358_n300# a_n458_n344# a_n562_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_1070_n300# a_970_n344# a_866_n300# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.5u
X2 a_458_n300# a_358_n344# a_254_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
X3 a_n766_n300# a_n866_n344# a_n970_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
X4 a_866_n300# a_766_n344# a_662_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
X5 a_n154_n300# a_n254_n344# a_n358_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
X6 a_50_n300# a_n50_n344# a_n154_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
X7 a_254_n300# a_154_n344# a_50_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
X8 a_n562_n300# a_n662_n344# a_n766_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
X9 a_n970_n300# a_n1070_n344# a_n1158_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.5u
X10 a_662_n300# a_562_n344# a_458_n300# VSUBS nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.5u
.ends

.subckt nfet_03v3_8Z2ENZ a_n138_n300# a_50_n300# a_n50_n344# VSUBS
X0 a_50_n300# a_n50_n344# a_n138_n300# VSUBS nfet_03v3 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.5u
.ends

.subckt BIASING_1m_MAGIC VDD IOUT G_SINK_UP G_SINK_DOWN VSS
Xpfet_03v3_GKYWHF_0 VDD a_207_1485# a_207_1485# IOUT VDD VDD a_207_1485# IOUT IOUT
+ VDD IOUT a_207_1485# a_207_1485# a_207_1485# a_207_1485# a_207_1485# a_207_1485#
+ IOUT VDD IOUT a_207_1485# VDD a_207_1485# a_207_1485# IOUT a_207_1485# VDD VDD IOUT
+ a_207_1485# a_207_1485# IOUT VDD a_207_1485# IOUT a_207_1485# IOUT VDD a_207_1485#
+ VDD VDD a_207_1485# a_207_1485# IOUT a_207_1485# VDD pfet_03v3_GKYWHF
Xpfet_03v3_GKYJHF_0 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pfet_03v3_GKYJHF
Xpfet_03v3_GKYJHF_1 a_207_1485# a_207_1485# VDD a_207_1485# a_207_1485# VDD a_207_1485#
+ a_207_1485# VDD VDD pfet_03v3_GKYJHF
Xpfet_03v3_GKYJHF_2 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD pfet_03v3_GKYJHF
Xnfet_03v3_U5DXAV_0 a_207_1485# G_SINK_UP m1_221_n1033# G_SINK_UP G_SINK_UP G_SINK_UP
+ m1_221_n1033# a_207_1485# G_SINK_UP m1_221_n1033# a_207_1485# G_SINK_UP a_207_1485#
+ m1_221_n1033# a_207_1485# a_207_1485# G_SINK_UP G_SINK_UP G_SINK_UP G_SINK_UP m1_221_n1033#
+ m1_221_n1033# G_SINK_UP VSS nfet_03v3_U5DXAV
Xnfet_03v3_U5DXAV_1 VSS G_SINK_DOWN m1_221_n1033# G_SINK_DOWN G_SINK_DOWN G_SINK_DOWN
+ m1_221_n1033# VSS G_SINK_DOWN m1_221_n1033# VSS G_SINK_DOWN VSS m1_221_n1033# VSS
+ VSS G_SINK_DOWN G_SINK_DOWN G_SINK_DOWN G_SINK_DOWN m1_221_n1033# m1_221_n1033#
+ G_SINK_DOWN VSS nfet_03v3_U5DXAV
Xnfet_03v3_8Z2ENZ_0 VSS VSS VSS VSS nfet_03v3_8Z2ENZ
Xnfet_03v3_8Z2ENZ_1 m1_221_n1033# a_207_1485# G_SINK_UP VSS nfet_03v3_8Z2ENZ
Xnfet_03v3_8Z2ENZ_2 VSS VSS VSS VSS nfet_03v3_8Z2ENZ
Xnfet_03v3_8Z2ENZ_3 VSS VSS VSS VSS nfet_03v3_8Z2ENZ
Xnfet_03v3_8Z2ENZ_4 m1_221_n1033# VSS G_SINK_DOWN VSS nfet_03v3_8Z2ENZ
Xnfet_03v3_8Z2ENZ_5 VSS VSS VSS VSS nfet_03v3_8Z2ENZ
.ends

.subckt pmos_3p3_MNHNAR a_28_404# a_n28_n312# a_n28_360# a_28_68# a_28_n268# w_n202_n734#
+ a_n116_n268# a_28_n604# a_n28_n648# a_n28_24# a_n116_n604# a_n116_68# a_n116_404#
X0 a_28_n268# a_n28_n312# a_n116_n268# w_n202_n734# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_28_n604# a_n28_n648# a_n116_n604# w_n202_n734# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X2 a_28_68# a_n28_24# a_n116_68# w_n202_n734# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X3 a_28_404# a_n28_360# a_n116_404# w_n202_n734# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt nmos_3p3_K66RT2 a_n28_n312# a_28_68# a_28_n268# a_n116_n268# a_n28_24# a_n116_68#
+ VSUBS
X0 a_28_68# a_n28_24# a_n116_68# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_28_n268# a_n28_n312# a_n116_n268# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt nmos_3p3_CU6RT2 a_108_n268# a_n428_n312# a_428_68# a_268_n268# a_268_68# a_n52_68#
+ a_52_24# a_108_68# a_428_n268# a_372_24# a_52_n312# a_n52_n268# a_n372_68# a_212_24#
+ a_n428_24# a_n516_n268# a_n108_n312# a_212_n312# a_n212_68# a_n212_n268# a_n268_24#
+ a_n268_n312# a_372_n312# a_n108_24# a_n372_n268# a_n516_68# VSUBS
X0 a_268_68# a_212_24# a_108_68# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n372_68# a_n428_24# a_n516_68# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 a_n372_n268# a_n428_n312# a_n516_n268# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 a_n212_68# a_n268_24# a_n372_68# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_108_n268# a_52_n312# a_n52_n268# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_428_n268# a_372_n312# a_268_n268# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_268_n268# a_212_n312# a_108_n268# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_n52_68# a_n108_24# a_n212_68# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 a_n212_n268# a_n268_n312# a_n372_n268# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_n52_n268# a_n108_n312# a_n212_n268# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X10 a_108_68# a_52_24# a_n52_68# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X11 a_428_68# a_372_24# a_268_68# VSUBS nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt pmos_3p3_MENMAR a_108_n268# a_n428_n312# a_428_68# a_n52_404# a_n372_n604#
+ a_n516_404# a_212_360# a_268_n268# a_268_68# a_n52_68# a_52_24# a_428_404# a_372_360#
+ a_52_n648# a_108_n604# a_108_68# a_n108_n648# a_212_n648# a_428_n268# a_372_24#
+ a_268_n604# w_n602_n734# a_52_n312# a_n212_404# a_n428_360# a_n52_n268# a_n372_404#
+ a_n372_68# a_212_24# a_n268_n648# a_n428_24# a_372_n648# a_n516_n268# a_n108_n312#
+ a_212_n312# a_n212_68# a_108_404# a_428_n604# a_n212_n268# a_268_404# a_n268_24#
+ a_52_360# a_n52_n604# a_n428_n648# a_n268_n312# a_372_n312# a_n108_24# a_n516_n604#
+ a_n372_n268# a_n108_360# a_n212_n604# a_n516_68# a_n268_360#
X0 a_n52_404# a_n108_360# a_n212_404# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_268_68# a_212_24# a_108_68# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n372_68# a_n428_24# a_n516_68# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 a_n212_404# a_n268_360# a_n372_404# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_n372_n268# a_n428_n312# a_n516_n268# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X5 a_n212_68# a_n268_24# a_n372_68# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_108_n268# a_52_n312# a_n52_n268# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_428_n268# a_372_n312# a_268_n268# w_n602_n734# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X8 a_268_n268# a_212_n312# a_108_n268# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_108_404# a_52_360# a_n52_404# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X10 a_n372_n604# a_n428_n648# a_n516_n604# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X11 a_n52_68# a_n108_24# a_n212_68# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X12 a_n212_n268# a_n268_n312# a_n372_n268# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X13 a_268_404# a_212_360# a_108_404# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X14 a_n52_n268# a_n108_n312# a_n212_n268# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X15 a_108_68# a_52_24# a_n52_68# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X16 a_108_n604# a_52_n648# a_n52_n604# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X17 a_428_n604# a_372_n648# a_268_n604# w_n602_n734# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X18 a_n372_404# a_n428_360# a_n516_404# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X19 a_268_n604# a_212_n648# a_108_n604# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X20 a_428_404# a_372_360# a_268_404# w_n602_n734# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X21 a_n212_n604# a_n268_n648# a_n372_n604# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X22 a_n52_n604# a_n108_n648# a_n212_n604# w_n602_n734# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X23 a_428_68# a_372_24# a_268_68# w_n602_n734# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt TG_magic B VSS CLK A VDD
Xpmos_3p3_MNHNAR_0 a_614_229# CLK CLK a_614_229# a_614_229# VDD VDD a_614_229# CLK
+ CLK VDD VDD VDD pmos_3p3_MNHNAR
Xnmos_3p3_K66RT2_0 CLK a_614_229# a_614_229# VSS CLK VSS VSS nmos_3p3_K66RT2
Xnmos_3p3_CU6RT2_0 A CLK A B B B CLK A A CLK CLK B B CLK CLK A CLK CLK A A CLK CLK
+ CLK CLK B A VSS nmos_3p3_CU6RT2
Xpmos_3p3_MENMAR_0 A a_614_229# A B B A a_614_229# B B B a_614_229# A a_614_229# a_614_229#
+ A A a_614_229# a_614_229# A a_614_229# B VDD a_614_229# A a_614_229# B B B a_614_229#
+ a_614_229# a_614_229# a_614_229# A a_614_229# a_614_229# A A A A B a_614_229# a_614_229#
+ B a_614_229# a_614_229# a_614_229# a_614_229# A B a_614_229# A A a_614_229# pmos_3p3_MENMAR
.ends

.subckt pmos_3p3_MWBYAR a_108_n268# a_n356_68# a_268_n268# a_268_68# a_n52_68# a_52_24#
+ a_108_68# a_n356_n268# a_52_n312# a_n52_n268# a_212_24# a_n108_n312# a_212_n312#
+ a_n212_68# a_n212_n268# a_n268_24# a_n268_n312# a_n108_24# w_n442_n398#
X0 a_268_68# a_212_24# a_108_68# w_n442_n398# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_n212_68# a_n268_24# a_n356_68# w_n442_n398# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 a_108_n268# a_52_n312# a_n52_n268# w_n442_n398# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_268_n268# a_212_n312# a_108_n268# w_n442_n398# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_n52_68# a_n108_24# a_n212_68# w_n442_n398# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_n212_n268# a_n268_n312# a_n356_n268# w_n442_n398# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X6 a_n52_n268# a_n108_n312# a_n212_n268# w_n442_n398# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_108_68# a_52_24# a_n52_68# w_n442_n398# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_MEGST2 a_n212_n168# a_n268_n212# a_n356_68# a_268_68# a_n52_68# a_52_24#
+ a_108_68# a_108_n168# a_268_n168# a_212_24# a_n212_68# a_n356_n168# a_n268_24# a_52_n212#
+ a_n52_n168# a_n108_24# a_n108_n212# a_212_n212# VSUBS
X0 a_268_68# a_212_24# a_108_68# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 a_n212_68# a_n268_24# a_n356_68# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 a_n52_68# a_n108_24# a_n212_68# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X3 a_108_68# a_52_24# a_n52_68# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 a_108_n168# a_52_n212# a_n52_n168# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 a_268_n168# a_212_n212# a_108_n168# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X6 a_n212_n168# a_n268_n212# a_n356_n168# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X7 a_n52_n168# a_n108_n212# a_n212_n168# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
.ends

.subckt INVERTER_MUX VDD VSS IN OUT
Xpmos_3p3_MWBYAR_0 OUT VDD VDD VDD VDD IN OUT VDD IN VDD IN IN IN OUT OUT IN IN IN
+ VDD pmos_3p3_MWBYAR
Xnmos_3p3_MEGST2_0 OUT IN VSS VSS VSS IN OUT OUT VSS IN OUT VSS IN IN VSS IN IN IN
+ VSS nmos_3p3_MEGST2
.ends

.subckt TG_GATE_SWITCH_magic B VDD VSS A CLK
Xpmos_3p3_MNHNAR_0 a_42_9# CLK CLK a_42_9# a_42_9# VDD VDD a_42_9# CLK CLK VDD VDD
+ VDD pmos_3p3_MNHNAR
Xpmos_3p3_MNHNAR_1 a_614_229# a_42_9# a_42_9# a_614_229# a_614_229# VDD VDD a_614_229#
+ a_42_9# a_42_9# VDD VDD VDD pmos_3p3_MNHNAR
Xnmos_3p3_K66RT2_1 a_42_9# a_614_229# a_614_229# VSS a_42_9# VSS VSS nmos_3p3_K66RT2
Xnmos_3p3_K66RT2_2 CLK a_42_9# a_42_9# VSS CLK VSS VSS nmos_3p3_K66RT2
Xnmos_3p3_CU6RT2_0 A a_42_9# A B B B a_42_9# A A a_42_9# a_42_9# B B a_42_9# a_42_9#
+ A a_42_9# a_42_9# A A a_42_9# a_42_9# a_42_9# a_42_9# B A VSS nmos_3p3_CU6RT2
Xpmos_3p3_MENMAR_0 A a_614_229# A B B A a_614_229# B B B a_614_229# A a_614_229# a_614_229#
+ A A a_614_229# a_614_229# A a_614_229# B VDD a_614_229# A a_614_229# B B B a_614_229#
+ a_614_229# a_614_229# a_614_229# A a_614_229# a_614_229# A A A A B a_614_229# a_614_229#
+ B a_614_229# a_614_229# a_614_229# a_614_229# A B a_614_229# A A a_614_229# pmos_3p3_MENMAR
.ends

.subckt MUX_1x8 S0 A0 A2 A6 A4 S2 S1 A3 A7 ENA A5 A1 Vout VSS VDD
XTG_magic_13 TG_magic_7/A VSS S0 TG_magic_13/A VDD TG_magic
XINVERTER_MUX_0 VDD VSS S0 TG_magic_6/CLK INVERTER_MUX
XINVERTER_MUX_1 VDD VSS S2 TG_magic_8/CLK INVERTER_MUX
XTG_GATE_SWITCH_magic_0 TG_magic_6/A VDD VSS A0 ENA TG_GATE_SWITCH_magic
XINVERTER_MUX_2 VDD VSS S1 TG_magic_7/CLK INVERTER_MUX
XTG_GATE_SWITCH_magic_1 TG_magic_1/A VDD VSS A3 ENA TG_GATE_SWITCH_magic
XTG_magic_0 TG_magic_8/A VSS TG_magic_7/CLK TG_magic_6/B VDD TG_magic
XTG_GATE_SWITCH_magic_2 TG_magic_13/A VDD VSS A5 ENA TG_GATE_SWITCH_magic
XTG_GATE_SWITCH_magic_3 TG_magic_3/A VDD VSS A6 ENA TG_GATE_SWITCH_magic
XTG_magic_1 TG_magic_9/A VSS TG_magic_6/CLK TG_magic_1/A VDD TG_magic
XTG_magic_2 TG_magic_7/A VSS TG_magic_6/CLK TG_magic_2/A VDD TG_magic
XTG_GATE_SWITCH_magic_4 TG_magic_2/A VDD VSS A1 ENA TG_GATE_SWITCH_magic
XTG_magic_3 TG_magic_5/A VSS S0 TG_magic_3/A VDD TG_magic
XTG_GATE_SWITCH_magic_5 TG_magic_4/A VDD VSS A7 ENA TG_GATE_SWITCH_magic
XTG_GATE_SWITCH_magic_7 TG_magic_11/A VDD VSS A2 ENA TG_GATE_SWITCH_magic
XTG_GATE_SWITCH_magic_6 TG_magic_10/A VDD VSS A4 ENA TG_GATE_SWITCH_magic
XTG_magic_4 TG_magic_9/A VSS S0 TG_magic_4/A VDD TG_magic
XTG_magic_5 TG_magic_8/A VSS S1 TG_magic_5/A VDD TG_magic
XTG_magic_6 TG_magic_6/B VSS TG_magic_6/CLK TG_magic_6/A VDD TG_magic
XTG_magic_10 TG_magic_6/B VSS S0 TG_magic_10/A VDD TG_magic
XTG_magic_8 Vout VSS TG_magic_8/CLK TG_magic_8/A VDD TG_magic
XTG_magic_7 TG_magic_9/B VSS TG_magic_7/CLK TG_magic_7/A VDD TG_magic
XTG_magic_11 TG_magic_5/A VSS TG_magic_6/CLK TG_magic_11/A VDD TG_magic
XTG_magic_9 TG_magic_9/B VSS S1 TG_magic_9/A VDD TG_magic
XTG_magic_12 Vout VSS S2 TG_magic_9/B VDD TG_magic
.ends

.subckt AWG_MUX_MAGIC A0 A1 A5 A3 A7 A4 A2 A6 A6_B A2_B A0_B A4_B A7_B A3_B A1_B A5_B
+ S2 S1 S0 ENA IN_P IN_N IBIAS VDD VSS G_SINK_UP G_SINK_DOWN S_PGA_1 S_PGA_2 S_PGA_3
+ PGA_P_T PGA_N_T FIL_P_T FIL_N_T IV_P_T IV_N_T
XPGA_MAGIC_0 PGA_MAGIC_0/BD PGA_MAGIC_0/IND PGA_MAGIC_0/IPD VSS PGA_MAGIC_0/VB4 PGA_MAGIC_0/VB2
+ PGA_MAGIC_0/VB3 PGA_MAGIC_0/VB1 PGA_MAGIC_0/VND PGA_MAGIC_0/VPD PGA_MAGIC_0/IBIAS1
+ PGA_MAGIC_0/VBIASN PGA_MAGIC_0/VOUT PGA_MAGIC_0/VBM PGA_MAGIC_0/VCD PGA_MAGIC_0/IBIAS4
+ PGA_MAGIC_0/IBIAS3 PGA_MAGIC_0/IBS PGA_P_T PGA_N_T PGA_MAGIC_0/IBIAS2 PGA_MAGIC_0/IBIAS
+ PGA_MAGIC_0/VCM PGA_MAGIC_0/IVS PGA_MAGIC_0/IB4 PGA_MAGIC_0/IB2 PGA_MAGIC_0/IB3
+ PGA_MAGIC_0/IB5 PGA_MAGIC_0/IN_P PGA_MAGIC_0/IN_N PGA_MAGIC_0/OUT1 PGA_MAGIC_0/OUT2
+ FIL_N_T FIL_P_T S_PGA_1 S_PGA_2 S_PGA_3 VDD PGA_MAGIC
XVCM_1.3V_magic_0 VDD VSS Filter_magic_0/VCM1 VCM_1.3V_magic
Xfold_cascode_opamp_mag_0 VDD VSS IN_N IV_N_T fold_cascode_opamp_mag_0/OUT fold_cascode_opamp_mag_0/VC
+ fold_cascode_opamp_mag_0/VD fold_cascode_opamp_mag_0/VX fold_cascode_opamp_mag_0/VA
+ fold_cascode_opamp_mag_0/VB fold_cascode_opamp_mag_0/VBS2 fold_cascode_opamp_mag_0/VBS3
+ fold_cascode_opamp_mag_0/VBIASN fold_cascode_opamp_mag_0/IBIAS2 fold_cascode_opamp_mag_0/VBIASN2
+ fold_cascode_opamp_mag_0/IBIAS3 fold_cascode_opamp_mag_0/IBIAS IV_N_T fold_cascode_opamp_mag_0/VP
+ fold_cascode_opamp_mag_0/c_mid fold_cascode_opamp_mag
Xfold_cascode_opamp_mag_1 VDD VSS IN_P IV_P_T fold_cascode_opamp_mag_1/OUT fold_cascode_opamp_mag_1/VC
+ fold_cascode_opamp_mag_1/VD fold_cascode_opamp_mag_1/VX fold_cascode_opamp_mag_1/VA
+ fold_cascode_opamp_mag_1/VB fold_cascode_opamp_mag_1/VBS2 fold_cascode_opamp_mag_1/VBS3
+ fold_cascode_opamp_mag_1/VBIASN fold_cascode_opamp_mag_1/IBIAS2 fold_cascode_opamp_mag_1/VBIASN2
+ fold_cascode_opamp_mag_1/IBIAS3 IBIAS IV_P_T fold_cascode_opamp_mag_1/VP fold_cascode_opamp_mag_1/c_mid
+ fold_cascode_opamp_mag
XVCM_1.6_MAGIC_0 VDD VSS PGA_MAGIC_0/VCM VCM_1.6_MAGIC
XBIASING_CURRENT_MAGIC_0 IBIAS fold_cascode_opamp_mag_0/IBIAS Filter_magic_0/IBIAS11
+ PGA_MAGIC_0/IBIAS1 G_SINK_UP G_SINK_DOWN VSS BIASING_CURRENT_MAGIC
XFilter_magic_0 IV_N_T FIL_N_T VDD VSS Filter_magic_0/VOUT_OPAMP_P Filter_magic_0/VOUT_OPAMP_N
+ IV_P_T Filter_magic_0/R3_R7_1 Filter_magic_0/R7_R8_R10_C1 Filter_magic_0/IB21 Filter_magic_0/IBIAS11
+ Filter_magic_0/VBM1 Filter_magic_0/VBIASN1 Filter_magic_0/IB31 Filter_magic_0/IBS1
+ Filter_magic_0/VB21 Filter_magic_0/VB31 Filter_magic_0/VB41 Filter_magic_0/VCD1
+ Filter_magic_0/IND1 Filter_magic_0/IPD1 Filter_magic_0/OUT2_1 Filter_magic_0/OUT1_1
+ Filter_magic_0/IBIAS3_1 Filter_magic_0/IB4_1 Filter_magic_0/IBIAS4_1 Filter_magic_0/IVS_1
+ Filter_magic_0/IBIAS2_1 Filter_magic_0/VB1_1 Filter_magic_0/BD_1 Filter_magic_0/R_1
+ Filter_magic_0/R11_1 Filter_magic_0/OPAMP_C_1 Filter_magic_0/OPAMP_C1_1 Filter_magic_0/VOUT_1_1
+ FIL_P_T Filter_magic_0/VCM1 Filter_magic
X200_ohm_magic_0 IN_P IN_N VSS VDD x200_ohm_magic
XBIASING_1m_MAGIC_0 VDD IN_N G_SINK_UP G_SINK_DOWN VSS BIASING_1m_MAGIC
XMUX_1x8_0 S0 A0_B A2_B A6_B A4_B S2 S1 A3_B A7_B ENA A5_B A1_B PGA_P_T VSS VDD MUX_1x8
XBIASING_1m_MAGIC_1 VDD IN_P G_SINK_UP G_SINK_DOWN VSS BIASING_1m_MAGIC
XMUX_1x8_1 S0 A0 A2 A6 A4 S2 S1 A3 A7 ENA A5 A1 PGA_N_T VSS VDD MUX_1x8
.ends

