magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1047 -1075 1047 1075
<< metal2 >>
rect -47 70 47 75
rect -47 42 -42 70
rect -14 42 14 70
rect 42 42 47 70
rect -47 14 47 42
rect -47 -14 -42 14
rect -14 -14 14 14
rect 42 -14 47 14
rect -47 -42 47 -14
rect -47 -70 -42 -42
rect -14 -70 14 -42
rect 42 -70 47 -42
rect -47 -75 47 -70
<< via2 >>
rect -42 42 -14 70
rect 14 42 42 70
rect -42 -14 -14 14
rect 14 -14 42 14
rect -42 -70 -14 -42
rect 14 -70 42 -42
<< metal3 >>
rect -47 70 47 75
rect -47 42 -42 70
rect -14 42 14 70
rect 42 42 47 70
rect -47 14 47 42
rect -47 -14 -42 14
rect -14 -14 14 14
rect 42 -14 47 14
rect -47 -42 47 -14
rect -47 -70 -42 -42
rect -14 -70 14 -42
rect 42 -70 47 -42
rect -47 -75 47 -70
<< end >>
