* NGSPICE file created from folded_single_check5_flat.ext - technology: gf180mcuC

.subckt folded_single_check5_flat
R0 a_n2777_n5169.t0 a_n2777_n5169.n0 1.21383
R1 a_n2617_n5169.n0 a_n2617_n5169.t1 1.21383
R2 a_n3086_n6147.t1 a_n3086_n6147.t0 59.8509
R3 a_n2937_n6021.t0 a_n2937_n6021.n0 1.21383
R4 a_n1817_n6021.t0 a_n1817_n6021.n0 1.21383
R5 a_n1657_n6021.t0 a_n1657_n6021.n0 1.21383
R6 a_n3083_n5296.t1 a_n3083_n5296.t0 59.7671
R7 a_n2937_n5169.t0 a_n2937_n5169.n0 1.21383
R8 a_n2137_n6021.n0 a_n2137_n6021.t1 1.21383
R9 a_n1977_n6021.t0 a_n1977_n6021.n0 1.21383
R10 a_n2617_n6021.t0 a_n2617_n6021.n0 1.21383
R11 a_n2457_n6021.t0 a_n2457_n6021.n0 1.21383
R12 a_n1817_n5169.n0 a_n1817_n5169.t1 1.21383
R13 a_n1657_n5169.n0 a_n1657_n5169.t1 1.21383
R14 a_n1553_n6152.n0 a_n1553_n6152.t0 59.4488
R15 a_n2137_n5169.t0 a_n2137_n5169.n0 1.21383
R16 a_n1977_n5169.t0 a_n1977_n5169.n0 1.21383
R17 a_n2457_n5169.n0 a_n2457_n5169.t1 1.21383
R18 a_n2297_n6021.n0 a_n2297_n6021.t1 1.21383
R19 a_n2777_n6021.n0 a_n2777_n6021.t1 1.21383
R20 a_n1553_n5305.n0 a_n1553_n5305.t0 59.084
R21 a_n2297_n5169.t0 a_n2297_n5169.n0 1.21383
C0 a_n2845_n5323# a_n2849_n6153# 0.213f
C1 a_n2849_n6153# a_n2688_n4484# 2.58e-22
C2 a_n2845_n5323# w_n3327_n6363# 1.09f
C3 w_n3327_n6363# a_n2688_n4484# 0.735f
C4 w_n3327_n6363# a_n3086_n4453# 0.196f
C5 a_n2845_n5323# a_n2688_n4484# 0.192f
C6 w_n3327_n6363# a_n1553_n4448# 0.204f
C7 a_n3086_n4453# a_n2688_n4484# 0.0102f
C8 a_n1553_n4448# a_n2688_n4484# 0.0219f
C9 a_n1553_n4448# a_n3086_n4453# 0.00192f
C10 w_n3327_n6363# a_n2849_n6153# 1.21f
C11 a_n2849_n6153# VSUBS 0.138f $ **FLOATING
C12 a_n2845_n5323# VSUBS 0.26f $ **FLOATING
C13 a_n1553_n4448# VSUBS 0.0379f $ **FLOATING
C14 a_n2688_n4484# VSUBS 0.312f $ **FLOATING
C15 a_n3086_n4453# VSUBS 0.0363f $ **FLOATING
C16 w_n3327_n6363# VSUBS 14.6f $ **FLOATING
.ends

