* NGSPICE file created from Stage_INV_flat.ext - technology: gf180mcuC

.subckt GF_INV_STAGE_PEX VSS VDD OUT IN
X0 VDD IN.t0 OUT.t7 VDD.t7 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X1 VSS IN.t1 OUT.t1 VSS.t7 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X2 OUT IN.t2 VSS.t6 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X3 OUT IN.t3 VDD.t6 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X4 VSS IN.t4 OUT.t0 VSS.t2 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X5 VDD IN.t5 OUT.t6 VDD.t2 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X6 OUT IN.t6 VDD.t1 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X7 OUT IN.t7 VSS.t1 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
R0 IN.n0 IN.t1 19.1891
R1 IN.n1 IN.t2 19.1891
R2 IN.n2 IN.t4 19.1891
R3 IN.n3 IN.t7 18.6676
R4 IN.n1 IN.n0 16.9365
R5 IN.n2 IN.n1 16.9365
R6 IN.n3 IN.n2 16.6457
R7 IN.n0 IN.t5 11.6805
R8 IN.n1 IN.t6 11.6805
R9 IN.n2 IN.t0 11.6805
R10 IN.n3 IN.t3 11.4719
R11 IN IN.n3 9.89085
R12 OUT.n1 OUT.t6 3.6405
R13 OUT.n1 OUT.n0 3.6405
R14 OUT.n5 OUT.t7 3.6405
R15 OUT.n5 OUT.n4 3.6405
R16 OUT.n9 OUT.n3 3.48898
R17 OUT.n8 OUT.n7 3.48898
R18 OUT.n9 OUT.n1 2.89789
R19 OUT.n8 OUT.n5 2.89789
R20 OUT.n3 OUT.t1 1.6385
R21 OUT.n3 OUT.n2 1.6385
R22 OUT.n7 OUT.t0 1.6385
R23 OUT.n7 OUT.n6 1.6385
R24 OUT.n9 OUT.n8 0.68137
R25 OUT OUT.n9 0.370283
R26 VDD.n3 VDD.t2 179.427
R27 VDD.n9 VDD.t7 112.441
R28 VDD.n6 VDD.t0 52.6321
R29 VDD.n11 VDD.t5 23.9239
R30 VDD.n5 VDD.n2 6.66125
R31 VDD.n13 VDD.t6 6.58259
R32 VDD.n1 VDD.t1 3.6405
R33 VDD.n1 VDD.n0 3.6405
R34 VDD.n17 VDD.n10 3.1505
R35 VDD.n10 VDD.n9 3.1505
R36 VDD.n16 VDD.n15 3.1505
R37 VDD.n15 VDD.n14 3.1505
R38 VDD.n5 VDD.n4 3.1505
R39 VDD.n4 VDD.n3 3.1505
R40 VDD.n8 VDD.n7 3.1505
R41 VDD.n7 VDD.n6 3.1505
R42 VDD.n13 VDD.n12 3.1505
R43 VDD.n12 VDD.n11 3.1505
R44 VDD VDD.n1 2.82941
R45 VDD.n8 VDD.n5 0.143789
R46 VDD.n17 VDD.n16 0.127211
R47 VDD.n16 VDD.n13 0.123658
R48 VDD VDD.n8 0.0774737
R49 VDD VDD.n17 0.0478684
R50 VSS.n60 VSS.n59 317.899
R51 VSS.n7 VSS.n6 313.262
R52 VSS.n41 VSS.t0 141.304
R53 VSS.n31 VSS.t7 134.239
R54 VSS.n38 VSS.t2 49.457
R55 VSS.n34 VSS.t5 42.3918
R56 VSS.n69 VSS.n68 24.2542
R57 VSS.n16 VSS.n15 23.8976
R58 VSS.n30 VSS.n2 5.15437
R59 VSS VSS.t1 5.11524
R60 VSS.n37 VSS.n1 3.51637
R61 VSS.n11 VSS.n10 2.6005
R62 VSS.n10 VSS.n9 2.6005
R63 VSS.n23 VSS.n22 2.6005
R64 VSS.n20 VSS.n19 2.6005
R65 VSS.n18 VSS.n17 2.6005
R66 VSS.n17 VSS.n16 2.6005
R67 VSS.n14 VSS.n13 2.6005
R68 VSS.n13 VSS.n12 2.6005
R69 VSS.n8 VSS.n7 2.6005
R70 VSS.n5 VSS.n4 2.6005
R71 VSS.n4 VSS.n3 2.6005
R72 VSS.n46 VSS.n45 2.6005
R73 VSS.n45 VSS.n44 2.6005
R74 VSS.n49 VSS.n48 2.6005
R75 VSS.n48 VSS.n47 2.6005
R76 VSS.n52 VSS.n51 2.6005
R77 VSS.n51 VSS.n50 2.6005
R78 VSS.n55 VSS.n54 2.6005
R79 VSS.n54 VSS.n53 2.6005
R80 VSS.n58 VSS.n57 2.6005
R81 VSS.n57 VSS.n56 2.6005
R82 VSS.n61 VSS.n60 2.6005
R83 VSS.n67 VSS.n66 2.6005
R84 VSS.n66 VSS.n65 2.6005
R85 VSS.n71 VSS.n70 2.6005
R86 VSS.n70 VSS.n69 2.6005
R87 VSS.n73 VSS.n72 2.6005
R88 VSS.n76 VSS.n75 2.6005
R89 VSS.n64 VSS.n63 2.6005
R90 VSS.n63 VSS.n62 2.6005
R91 VSS.n29 VSS.n28 2.6005
R92 VSS.n28 VSS.n27 2.6005
R93 VSS.n33 VSS.n32 2.6005
R94 VSS.n32 VSS.n31 2.6005
R95 VSS.n36 VSS.n35 2.6005
R96 VSS.n35 VSS.n34 2.6005
R97 VSS.n40 VSS.n39 2.6005
R98 VSS.n39 VSS.n38 2.6005
R99 VSS.n43 VSS.n42 2.6005
R100 VSS.n42 VSS.n41 2.6005
R101 VSS.n82 VSS.n81 2.6005
R102 VSS.n81 VSS.n80 2.6005
R103 VSS.n79 VSS.n78 2.6005
R104 VSS.n78 VSS.n77 2.6005
R105 VSS.n26 VSS.n25 2.6005
R106 VSS.n25 VSS.n24 2.6005
R107 VSS.n22 VSS.n21 1.90397
R108 VSS.n75 VSS.n74 1.90335
R109 VSS.n1 VSS.t6 1.6385
R110 VSS.n1 VSS.n0 1.6385
R111 VSS.n14 VSS.n11 0.183918
R112 VSS.n18 VSS.n14 0.183918
R113 VSS.n20 VSS.n18 0.183918
R114 VSS.n67 VSS.n64 0.183918
R115 VSS.n71 VSS.n67 0.183918
R116 VSS.n73 VSS.n71 0.183918
R117 VSS.n23 VSS.n20 0.182778
R118 VSS.n76 VSS.n73 0.182778
R119 VSS.n8 VSS.n5 0.177207
R120 VSS.n49 VSS.n46 0.177207
R121 VSS.n52 VSS.n49 0.177207
R122 VSS.n55 VSS.n52 0.177207
R123 VSS.n58 VSS.n55 0.177207
R124 VSS.n61 VSS.n58 0.177207
R125 VSS.n29 VSS.n26 0.177207
R126 VSS.n36 VSS.n33 0.177207
R127 VSS.n43 VSS.n40 0.177207
R128 VSS.n82 VSS.n79 0.177207
R129 VSS.n11 VSS.n8 0.139362
R130 VSS.n64 VSS.n61 0.137167
R131 VSS.n83 VSS.n43 0.117939
R132 VSS.n33 VSS.n30 0.116841
R133 VSS.n37 VSS.n36 0.0894024
R134 VSS.n40 VSS.n37 0.0883049
R135 VSS.n26 VSS.n23 0.0687711
R136 VSS.n79 VSS.n76 0.0687711
R137 VSS.n30 VSS.n29 0.0608659
R138 VSS.n83 VSS.n82 0.0597683
R139 VSS VSS.n83 0.0396304
C0 VDD IN 0.604f
C1 OUT VDD 0.343f
C2 OUT IN 0.209f
.ends

