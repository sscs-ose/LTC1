magic
tech gf180mcuC
magscale 1 10
timestamp 1691673501
<< nwell >>
rect 0 770 1172 901
<< psubdiff >>
rect 251 -161 793 -148
rect 251 -207 264 -161
rect 310 -207 358 -161
rect 404 -207 452 -161
rect 498 -207 546 -161
rect 592 -207 640 -161
rect 686 -207 734 -161
rect 780 -207 793 -161
rect 251 -220 793 -207
<< nsubdiff >>
rect 24 855 1143 868
rect 24 809 37 855
rect 83 809 131 855
rect 177 809 225 855
rect 271 809 319 855
rect 365 809 413 855
rect 459 809 507 855
rect 553 809 601 855
rect 647 809 708 855
rect 754 809 802 855
rect 848 809 896 855
rect 942 809 990 855
rect 1036 809 1084 855
rect 1130 809 1143 855
rect 24 796 1143 809
<< psubdiffcont >>
rect 264 -207 310 -161
rect 358 -207 404 -161
rect 452 -207 498 -161
rect 546 -207 592 -161
rect 640 -207 686 -161
rect 734 -207 780 -161
<< nsubdiffcont >>
rect 37 809 83 855
rect 131 809 177 855
rect 225 809 271 855
rect 319 809 365 855
rect 413 809 459 855
rect 507 809 553 855
rect 601 809 647 855
rect 708 809 754 855
rect 802 809 848 855
rect 896 809 942 855
rect 990 809 1036 855
rect 1084 809 1130 855
<< polysilicon >>
rect 174 364 390 420
rect 178 297 250 305
rect 334 297 390 364
rect 178 292 390 297
rect 178 246 191 292
rect 237 246 390 292
rect 178 241 390 246
rect 178 233 250 241
rect 334 162 390 241
rect 494 364 710 420
rect 494 162 550 364
rect 622 276 694 284
rect 942 276 998 446
rect 622 271 998 276
rect 622 225 635 271
rect 681 225 998 271
rect 622 220 998 225
rect 622 212 710 220
rect 654 166 710 212
rect 132 -24 204 -16
rect 494 -24 550 74
rect 132 -29 550 -24
rect 132 -75 145 -29
rect 191 -75 550 -29
rect 132 -80 550 -75
rect 132 -88 204 -80
<< polycontact >>
rect 191 246 237 292
rect 635 225 681 271
rect 145 -75 191 -29
<< metal1 >>
rect 0 855 1172 888
rect 0 809 37 855
rect 83 809 131 855
rect 177 809 225 855
rect 271 809 319 855
rect 365 809 413 855
rect 459 809 507 855
rect 553 809 601 855
rect 647 809 708 855
rect 754 809 802 855
rect 848 809 896 855
rect 942 809 990 855
rect 1036 809 1084 855
rect 1130 809 1172 855
rect 0 776 1172 809
rect 259 609 305 776
rect 419 684 785 730
rect 419 609 465 684
rect 739 584 785 684
rect 1027 609 1073 776
rect 99 396 145 470
rect 419 396 465 464
rect 99 350 465 396
rect 180 297 248 303
rect 97 292 248 297
rect 97 246 191 292
rect 237 246 248 292
rect 579 282 625 470
rect 867 344 913 470
rect 867 298 1087 344
rect 579 271 692 282
rect 579 258 635 271
rect 97 241 248 246
rect 180 235 248 241
rect 419 225 635 258
rect 681 225 692 271
rect 867 228 913 298
rect 419 214 692 225
rect 419 212 625 214
rect 419 124 465 212
rect 739 182 913 228
rect 134 -29 202 -18
rect 100 -75 145 -29
rect 191 -75 202 -29
rect 134 -86 202 -75
rect 259 -128 305 98
rect 579 -128 625 98
rect 739 93 785 182
rect 222 -161 822 -128
rect 222 -207 264 -161
rect 310 -207 358 -161
rect 404 -207 452 -161
rect 498 -207 546 -161
rect 592 -207 640 -161
rect 686 -207 734 -161
rect 780 -207 822 -161
rect 222 -240 822 -207
use nmos_3p3_GGGST2#3  nmos_3p3_GGGST2_0
timestamp 1691670445
transform 1 0 682 0 1 118
box -140 -118 140 118
use nmos_3p3_GGGST2#3  nmos_3p3_GGGST2_1
timestamp 1691670445
transform 1 0 362 0 1 118
box -140 -118 140 118
use nmos_3p3_GGGST2#3  nmos_3p3_GGGST2_2
timestamp 1691670445
transform 1 0 522 0 1 118
box -140 -118 140 118
use pmos_3p3_MEVUAR#0  pmos_3p3_MEVUAR_0
timestamp 1691247348
transform 1 0 602 0 1 540
box -282 -230 282 230
use pmos_3p3_MEVUAR#0  pmos_3p3_MEVUAR_1
timestamp 1691247348
transform 1 0 282 0 1 540
box -282 -230 282 230
use pmos_3p3_MNVUAR#3  pmos_3p3_MNVUAR_0
timestamp 1691670445
transform 1 0 970 0 1 540
box -202 -230 202 230
<< labels >>
flabel metal1 577 832 577 832 0 FreeSans 320 0 0 0 VDD
port 5 nsew
flabel metal1 530 -184 530 -184 0 FreeSans 320 0 0 0 VSS
port 6 nsew
flabel polycontact 214 269 214 269 0 FreeSans 320 0 0 0 A
port 7 nsew
flabel polycontact 168 -52 168 -52 0 FreeSans 320 0 0 0 B
port 8 nsew
flabel metal1 1064 322 1064 322 0 FreeSans 320 0 0 0 OUT
port 4 nsew
<< end >>
