magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2201 -8945 2201 8945
<< psubdiff >>
rect -201 6885 201 6945
rect -201 -6885 -179 6885
rect -133 -6885 -75 6885
rect -29 -6885 29 6885
rect 75 -6885 133 6885
rect 179 -6885 201 6885
rect -201 -6945 201 -6885
<< psubdiffcont >>
rect -179 -6885 -133 6885
rect -75 -6885 -29 6885
rect 29 -6885 75 6885
rect 133 -6885 179 6885
<< metal1 >>
rect -190 6885 190 6934
rect -190 -6885 -179 6885
rect -133 -6885 -75 6885
rect -29 -6885 29 6885
rect 75 -6885 133 6885
rect 179 -6885 190 6885
rect -190 -6934 190 -6885
<< end >>
