magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2280 -2045 2280 2045
<< psubdiff >>
rect -280 23 280 45
rect -280 -23 -258 23
rect 258 -23 280 23
rect -280 -45 280 -23
<< psubdiffcont >>
rect -258 -23 258 23
<< metal1 >>
rect -269 23 269 34
rect -269 -23 -258 23
rect 258 -23 269 23
rect -269 -34 269 -23
<< end >>
