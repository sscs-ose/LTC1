magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2645 -2128 2645 2128
<< nwell >>
rect -645 -128 645 128
<< nsubdiff >>
rect -562 23 562 45
rect -562 -23 -540 23
rect 540 -23 562 23
rect -562 -45 562 -23
<< nsubdiffcont >>
rect -540 -23 540 23
<< metal1 >>
rect -551 23 551 34
rect -551 -23 -540 23
rect 540 -23 551 23
rect -551 -34 551 -23
<< end >>
