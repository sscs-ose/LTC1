magic
tech gf180mcuC
magscale 1 10
timestamp 1695127730
<< metal1 >>
rect 687 1389 4520 1596
rect 570 1321 672 1329
rect 570 1243 578 1321
rect 662 1243 672 1321
rect 570 1233 672 1243
rect 564 1119 661 1137
rect 564 1053 577 1119
rect 649 1053 661 1119
rect 564 1048 661 1053
rect 2025 1085 2096 1088
rect 1596 1007 1714 1037
rect 2091 1033 2096 1085
rect 573 953 818 1000
rect 1596 979 1759 1007
rect 1656 949 1759 979
rect 2542 974 2656 1032
rect 2598 937 2656 974
rect 3493 1020 3621 1021
rect 3493 1004 3633 1020
rect 3493 963 3685 1004
rect 4457 974 4617 1032
rect 3580 948 3685 963
rect 566 901 686 906
rect 566 846 579 901
rect 674 846 686 901
rect 566 832 686 846
rect 565 770 696 776
rect 565 710 578 770
rect 683 710 696 770
rect 565 697 696 710
rect 1366 622 1653 679
rect 2313 622 2600 679
rect 3147 622 3162 671
rect 3254 622 3551 678
rect 4228 622 4515 678
rect 665 619 4515 622
rect 665 403 4507 619
<< via1 >>
rect 578 1243 662 1321
rect 577 1053 649 1119
rect 1071 1040 1137 1092
rect 2025 1033 2091 1085
rect 2969 1023 3038 1076
rect 3935 1033 4004 1086
rect 579 846 674 901
rect 578 710 683 770
<< metal2 >>
rect 570 1321 672 1329
rect 570 1243 578 1321
rect 662 1256 672 1321
rect 662 1243 767 1256
rect 570 1238 767 1243
rect 570 1233 3995 1238
rect 571 1232 3995 1233
rect 587 1199 3995 1232
rect 718 1164 3995 1199
rect 564 1119 661 1137
rect 564 1053 577 1119
rect 649 1094 661 1119
rect 649 1092 1186 1094
rect 649 1053 1071 1092
rect 564 1040 1071 1053
rect 1137 1040 1186 1092
rect 3921 1088 3995 1164
rect 564 1038 1186 1040
rect 2005 1085 2132 1088
rect 2005 1033 2025 1085
rect 2091 1033 2132 1085
rect 3919 1086 4047 1088
rect 2005 1030 2132 1033
rect 2956 1076 3083 1079
rect 566 901 686 906
rect 566 846 579 901
rect 674 897 686 901
rect 2040 897 2096 1030
rect 2956 1023 2969 1076
rect 3038 1023 3083 1076
rect 3919 1033 3935 1086
rect 4004 1033 4047 1086
rect 3919 1031 4047 1033
rect 2956 1019 3083 1023
rect 3921 1021 3995 1031
rect 674 846 2100 897
rect 566 841 2100 846
rect 566 832 686 841
rect 565 770 696 776
rect 565 710 578 770
rect 683 767 696 770
rect 2964 767 3020 1019
rect 683 711 3020 767
rect 683 710 696 711
rect 565 697 696 710
use and2_mag  and2_mag_0
timestamp 1695127730
transform 1 0 748 0 1 675
box -70 -188 1009 863
use and2_mag  and2_mag_1
timestamp 1695127730
transform 1 0 1694 0 1 670
box -70 -188 1009 863
use and2_mag  and2_mag_2
timestamp 1695127730
transform 1 0 2645 0 1 659
box -70 -188 1009 863
use and2_mag  and2_mag_3
timestamp 1695127730
transform 1 0 3609 0 1 670
box -70 -188 1009 863
<< labels >>
flabel via1 610 1084 610 1084 0 FreeSans 480 0 0 0 A
port 0 nsew
flabel metal1 598 976 598 976 0 FreeSans 480 0 0 0 B
port 1 nsew
flabel via1 610 868 612 870 0 FreeSans 480 0 0 0 C
port 2 nsew
flabel via1 617 741 617 741 0 FreeSans 480 0 0 0 D
port 3 nsew
flabel via1 607 1288 607 1288 0 FreeSans 480 0 0 0 E
port 4 nsew
flabel metal1 1463 1540 1463 1540 0 FreeSans 480 0 0 0 VDD
port 5 nsew
flabel metal1 1496 540 1496 540 0 FreeSans 480 0 0 0 VSS
port 6 nsew
flabel metal1 4584 1007 4584 1007 0 FreeSans 480 0 0 0 VOUT
port 7 nsew
<< end >>
