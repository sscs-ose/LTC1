magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2876 -2348 2876 2348
<< pwell >>
rect -876 -348 876 348
<< nmos >>
rect -764 -280 -664 280
rect -560 -280 -460 280
rect -356 -280 -256 280
rect -152 -280 -52 280
rect 52 -280 152 280
rect 256 -280 356 280
rect 460 -280 560 280
rect 664 -280 764 280
<< ndiff >>
rect -852 258 -764 280
rect -852 -258 -839 258
rect -793 -258 -764 258
rect -852 -280 -764 -258
rect -664 258 -560 280
rect -664 -258 -635 258
rect -589 -258 -560 258
rect -664 -280 -560 -258
rect -460 258 -356 280
rect -460 -258 -431 258
rect -385 -258 -356 258
rect -460 -280 -356 -258
rect -256 258 -152 280
rect -256 -258 -227 258
rect -181 -258 -152 258
rect -256 -280 -152 -258
rect -52 258 52 280
rect -52 -258 -23 258
rect 23 -258 52 258
rect -52 -280 52 -258
rect 152 258 256 280
rect 152 -258 181 258
rect 227 -258 256 258
rect 152 -280 256 -258
rect 356 258 460 280
rect 356 -258 385 258
rect 431 -258 460 258
rect 356 -280 460 -258
rect 560 258 664 280
rect 560 -258 589 258
rect 635 -258 664 258
rect 560 -280 664 -258
rect 764 258 852 280
rect 764 -258 793 258
rect 839 -258 852 258
rect 764 -280 852 -258
<< ndiffc >>
rect -839 -258 -793 258
rect -635 -258 -589 258
rect -431 -258 -385 258
rect -227 -258 -181 258
rect -23 -258 23 258
rect 181 -258 227 258
rect 385 -258 431 258
rect 589 -258 635 258
rect 793 -258 839 258
<< polysilicon >>
rect -764 280 -664 324
rect -560 280 -460 324
rect -356 280 -256 324
rect -152 280 -52 324
rect 52 280 152 324
rect 256 280 356 324
rect 460 280 560 324
rect 664 280 764 324
rect -764 -324 -664 -280
rect -560 -324 -460 -280
rect -356 -324 -256 -280
rect -152 -324 -52 -280
rect 52 -324 152 -280
rect 256 -324 356 -280
rect 460 -324 560 -280
rect 664 -324 764 -280
<< metal1 >>
rect -839 258 -793 278
rect -839 -278 -793 -258
rect -635 258 -589 278
rect -635 -278 -589 -258
rect -431 258 -385 278
rect -431 -278 -385 -258
rect -227 258 -181 278
rect -227 -278 -181 -258
rect -23 258 23 278
rect -23 -278 23 -258
rect 181 258 227 278
rect 181 -278 227 -258
rect 385 258 431 278
rect 385 -278 431 -258
rect 589 258 635 278
rect 589 -278 635 -258
rect 793 258 839 278
rect 793 -278 839 -258
<< end >>
