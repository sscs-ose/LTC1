magic
tech gf180mcuC
magscale 1 10
timestamp 1694155832
<< nwell >>
rect -864 -933 864 933
<< nsubdiff >>
rect -840 896 840 909
rect -840 850 -724 896
rect 724 850 840 896
rect -840 837 840 850
rect -840 793 -768 837
rect -840 -793 -827 793
rect -781 -793 -768 793
rect 768 793 840 837
rect -840 -837 -768 -793
rect 768 -793 781 793
rect 827 -793 840 793
rect 768 -837 840 -793
rect -840 -850 840 -837
rect -840 -896 -724 -850
rect 724 -896 840 -850
rect -840 -909 840 -896
<< nsubdiffcont >>
rect -724 850 724 896
rect -827 -793 -781 793
rect 781 -793 827 793
rect -724 -896 724 -850
<< polysilicon >>
rect -680 736 -520 749
rect -680 690 -667 736
rect -533 690 -520 736
rect -680 646 -520 690
rect -680 -690 -520 -646
rect -680 -736 -667 -690
rect -533 -736 -520 -690
rect -680 -749 -520 -736
rect -440 736 -280 749
rect -440 690 -427 736
rect -293 690 -280 736
rect -440 646 -280 690
rect -440 -690 -280 -646
rect -440 -736 -427 -690
rect -293 -736 -280 -690
rect -440 -749 -280 -736
rect -200 736 -40 749
rect -200 690 -187 736
rect -53 690 -40 736
rect -200 646 -40 690
rect -200 -690 -40 -646
rect -200 -736 -187 -690
rect -53 -736 -40 -690
rect -200 -749 -40 -736
rect 40 736 200 749
rect 40 690 53 736
rect 187 690 200 736
rect 40 646 200 690
rect 40 -690 200 -646
rect 40 -736 53 -690
rect 187 -736 200 -690
rect 40 -749 200 -736
rect 280 736 440 749
rect 280 690 293 736
rect 427 690 440 736
rect 280 646 440 690
rect 280 -690 440 -646
rect 280 -736 293 -690
rect 427 -736 440 -690
rect 280 -749 440 -736
rect 520 736 680 749
rect 520 690 533 736
rect 667 690 680 736
rect 520 646 680 690
rect 520 -690 680 -646
rect 520 -736 533 -690
rect 667 -736 680 -690
rect 520 -749 680 -736
<< polycontact >>
rect -667 690 -533 736
rect -667 -736 -533 -690
rect -427 690 -293 736
rect -427 -736 -293 -690
rect -187 690 -53 736
rect -187 -736 -53 -690
rect 53 690 187 736
rect 53 -736 187 -690
rect 293 690 427 736
rect 293 -736 427 -690
rect 533 690 667 736
rect 533 -736 667 -690
<< ppolyres >>
rect -680 -646 -520 646
rect -440 -646 -280 646
rect -200 -646 -40 646
rect 40 -646 200 646
rect 280 -646 440 646
rect 520 -646 680 646
<< metal1 >>
rect -827 850 -724 896
rect 724 850 827 896
rect -827 793 -781 850
rect 781 793 827 850
rect -678 690 -667 736
rect -533 690 -522 736
rect -438 690 -427 736
rect -293 690 -282 736
rect -198 690 -187 736
rect -53 690 -42 736
rect 42 690 53 736
rect 187 690 198 736
rect 282 690 293 736
rect 427 690 438 736
rect 522 690 533 736
rect 667 690 678 736
rect -678 -736 -667 -690
rect -533 -736 -522 -690
rect -438 -736 -427 -690
rect -293 -736 -282 -690
rect -198 -736 -187 -690
rect -53 -736 -42 -690
rect 42 -736 53 -690
rect 187 -736 198 -690
rect 282 -736 293 -690
rect 427 -736 438 -690
rect 522 -736 533 -690
rect 667 -736 678 -690
rect -827 -850 -781 -793
rect 781 -850 827 -793
rect -827 -896 -724 -850
rect 724 -896 827 -850
<< properties >>
string FIXED_BBOX -804 -873 804 873
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 6.459 m 1 nx 6 wmin 0.80 lmin 1.00 rho 315 val 2.787k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1
<< end >>
