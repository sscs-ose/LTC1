magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1316 1019 1316
<< metal1 >>
rect -19 310 19 316
rect -19 284 -13 310
rect 13 284 19 310
rect -19 256 19 284
rect -19 230 -13 256
rect 13 230 19 256
rect -19 202 19 230
rect -19 176 -13 202
rect 13 176 19 202
rect -19 148 19 176
rect -19 122 -13 148
rect 13 122 19 148
rect -19 94 19 122
rect -19 68 -13 94
rect 13 68 19 94
rect -19 40 19 68
rect -19 14 -13 40
rect 13 14 19 40
rect -19 -14 19 14
rect -19 -40 -13 -14
rect 13 -40 19 -14
rect -19 -68 19 -40
rect -19 -94 -13 -68
rect 13 -94 19 -68
rect -19 -122 19 -94
rect -19 -148 -13 -122
rect 13 -148 19 -122
rect -19 -176 19 -148
rect -19 -202 -13 -176
rect 13 -202 19 -176
rect -19 -230 19 -202
rect -19 -256 -13 -230
rect 13 -256 19 -230
rect -19 -284 19 -256
rect -19 -310 -13 -284
rect 13 -310 19 -284
rect -19 -316 19 -310
<< via1 >>
rect -13 284 13 310
rect -13 230 13 256
rect -13 176 13 202
rect -13 122 13 148
rect -13 68 13 94
rect -13 14 13 40
rect -13 -40 13 -14
rect -13 -94 13 -68
rect -13 -148 13 -122
rect -13 -202 13 -176
rect -13 -256 13 -230
rect -13 -310 13 -284
<< metal2 >>
rect -19 310 19 316
rect -19 284 -13 310
rect 13 284 19 310
rect -19 256 19 284
rect -19 230 -13 256
rect 13 230 19 256
rect -19 202 19 230
rect -19 176 -13 202
rect 13 176 19 202
rect -19 148 19 176
rect -19 122 -13 148
rect 13 122 19 148
rect -19 94 19 122
rect -19 68 -13 94
rect 13 68 19 94
rect -19 40 19 68
rect -19 14 -13 40
rect 13 14 19 40
rect -19 -14 19 14
rect -19 -40 -13 -14
rect 13 -40 19 -14
rect -19 -68 19 -40
rect -19 -94 -13 -68
rect 13 -94 19 -68
rect -19 -122 19 -94
rect -19 -148 -13 -122
rect 13 -148 19 -122
rect -19 -176 19 -148
rect -19 -202 -13 -176
rect 13 -202 19 -176
rect -19 -230 19 -202
rect -19 -256 -13 -230
rect 13 -256 19 -230
rect -19 -284 19 -256
rect -19 -310 -13 -284
rect 13 -310 19 -284
rect -19 -316 19 -310
<< end >>
