magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2845 -2345 2845 2345
<< psubdiff >>
rect -845 323 845 345
rect -845 -323 -823 323
rect 823 -323 845 323
rect -845 -345 845 -323
<< psubdiffcont >>
rect -823 -323 823 323
<< metal1 >>
rect -834 323 834 334
rect -834 -323 -823 323
rect 823 -323 834 323
rect -834 -334 834 -323
<< end >>
