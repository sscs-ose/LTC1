magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1721 1019 1721
<< metal2 >>
rect -19 716 19 721
rect -19 -716 -14 716
rect 14 -716 19 716
rect -19 -721 19 -716
<< via2 >>
rect -14 -716 14 716
<< metal3 >>
rect -19 716 19 721
rect -19 -716 -14 716
rect 14 -716 19 716
rect -19 -721 19 -716
<< end >>
