magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1097 1019 1097
<< metal1 >>
rect -19 91 19 97
rect -19 -91 -13 91
rect 13 -91 19 91
rect -19 -97 19 -91
<< via1 >>
rect -13 -91 13 91
<< metal2 >>
rect -19 91 19 97
rect -19 -91 -13 91
rect 13 -91 19 91
rect -19 -97 19 -91
<< end >>
