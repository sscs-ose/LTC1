magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -3961 2128 3961
<< nwell >>
rect -128 -1961 128 1961
<< nsubdiff >>
rect -45 1856 45 1878
rect -45 -1856 -23 1856
rect 23 -1856 45 1856
rect -45 -1878 45 -1856
<< nsubdiffcont >>
rect -23 -1856 23 1856
<< metal1 >>
rect -34 1856 34 1867
rect -34 -1856 -23 1856
rect 23 -1856 34 1856
rect -34 -1867 34 -1856
<< end >>
