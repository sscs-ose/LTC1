** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/4x1_mux_test_ibr..sch
**.subckt 4x1_mux_test_ibr.
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V4 S0 VSS pulse(3.3 0 0 100p 100p 200n 400n)
.save i(v4)
V6 I0 VSS pulse(0 3.3 0 100p 100p 100n 200n)3.3
.save i(v6)
V7 I1 VSS pulse(0 3.3 0 100p 100p 200n 400n)
.save i(v7)
V5 S1 VSS pulse(3.3 0 0 100p 100p 400n 800n)
.save i(v5)
V13 I2 VSS pulse(0 3.3 0 100p 100p 400n 800n)3.3
.save i(v13)
V14 I3 VSS pulse(0 3.3 0 100p 100p 800n 1600n)3.3
.save i(v14)
x1 VDD S1 VSS I2 I3 S0 I0 I1 OUT 4x1_mux_ibr.
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical




.control
save all
tran 50p 800n
plot v(S0) v(S1)+4  v(I0)+8 v(I1)+12 i2+16 i3+20  v(OUT)+24


*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  4x1_mux_ibr..sym # of pins=9
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/4x1_mux_ibr..sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/4x1_mux_ibr..sch
.subckt 4x1_mux_ibr. VDD S1 VSS I2 I3 S0 I0 I1 OUT
*.iopin VDD
*.iopin VSS
*.ipin S1
*.opin OUT
*.ipin I2
*.ipin I3
*.ipin S0
*.ipin I0
*.ipin I1
x1 VSS S0 net1 I0 I1 VDD 2x1_mux_ibr
x2 VSS S0 net2 I2 I3 VDD 2x1_mux_ibr
x3 VSS S1 OUT net1 net2 VDD 2x1_mux_ibr
.ends


* expanding   symbol:  2x1_mux_ibr.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/2x1_mux_ibr.sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/2x1_mux_ibr.sch
.subckt 2x1_mux_ibr VSS Sel OUT I0 I1 VDD
*.iopin VDD
*.iopin VSS
*.ipin Sel
*.opin OUT
*.ipin I0
*.ipin I1
x4 VSS Sel net1 VDD inv_my_ibr
x1 I0 VSS VDD net2 net1 NAND_ibr_mx2
x2 Sel VSS VDD net3 I1 NAND_ibr_mx2
x3 net2 VSS VDD OUT net3 NAND_ibr_mx2
.ends


* expanding   symbol:  inv_my_ibr.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/inv_my_ibr.sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/inv_my_ibr.sch
.subckt inv_my_ibr VSS IN OUT VDD
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  NAND_ibr_mx2.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/NAND_ibr_mx2.sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/NAND_ibr_mx2.sch
.subckt NAND_ibr_mx2 IN1 VSS VDD OUT IN2
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin OUT
XM3 net1 IN2 VSS VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 OUT IN1 net1 VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 OUT IN1 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN2 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
