magic
tech gf180mcuD
magscale 1 10
timestamp 1713275964
<< checkpaint >>
rect -2028 -2113 6062 5793
<< nwell >>
rect 133 3540 3680 3793
rect 2958 1781 3381 1813
rect 133 -113 3682 205
<< pwell >>
rect 194 2188 2495 2679
rect 196 1049 2496 1539
<< psubdiff >>
rect 2956 2634 3396 2675
rect 677 1906 1770 1958
rect 677 1860 909 1906
rect 1707 1860 1770 1906
rect 677 1801 1770 1860
rect 2964 963 2968 970
rect 2964 930 3375 963
rect 2968 929 3375 930
<< nsubdiff >>
rect 2958 1781 3381 1813
rect 705 46 2004 112
rect 705 0 911 46
rect 1803 0 2004 46
rect 705 -72 2004 0
<< psubdiffcont >>
rect 909 1860 1707 1906
<< nsubdiffcont >>
rect 911 0 1803 46
<< polysilicon >>
rect 253 2748 339 2776
rect 253 2702 272 2748
rect 318 2702 339 2748
rect 253 2684 339 2702
rect 239 1026 349 1062
rect 239 980 271 1026
rect 317 980 349 1026
rect 239 955 349 980
rect 239 950 350 955
<< polycontact >>
rect 272 2702 318 2748
rect 271 980 317 1026
<< metal1 >>
rect 133 3739 3680 3793
rect 133 3540 3900 3739
rect 3508 3529 3900 3540
rect 3634 3158 3712 3178
rect 2744 3129 2835 3142
rect 2744 3077 2770 3129
rect 2822 3077 2835 3129
rect 3634 3106 3649 3158
rect 3701 3106 3712 3158
rect 3634 3088 3712 3106
rect 2744 3062 2835 3077
rect 1536 3040 1624 3045
rect 1536 2988 1554 3040
rect 1606 2988 1624 3040
rect 1536 2975 1624 2988
rect 1984 2985 1988 2989
rect 259 2756 337 2770
rect 42 2748 337 2756
rect 42 2702 272 2748
rect 318 2702 337 2748
rect 42 2691 337 2702
rect 259 2685 337 2691
rect 520 2195 603 2210
rect 520 2143 535 2195
rect 587 2143 603 2195
rect 520 2125 603 2143
rect 2291 2198 2361 2205
rect 2291 2146 2302 2198
rect 2354 2146 2361 2198
rect 2291 2134 2361 2146
rect 2697 2044 2788 2804
rect 2956 2634 3396 2675
rect 3012 2243 3107 2265
rect 3012 2191 3035 2243
rect 3087 2191 3107 2243
rect 3012 2175 3107 2191
rect 3489 2262 3575 2283
rect 3489 2210 3502 2262
rect 3554 2210 3575 2262
rect 3489 2188 3575 2210
rect 515 1924 1770 1999
rect 2440 1955 2788 2044
rect 3758 1955 3900 3529
rect 2439 1924 2788 1955
rect 163 1906 2501 1924
rect 163 1860 909 1906
rect 1707 1860 2501 1906
rect 3410 1899 3900 1955
rect 163 1825 2501 1860
rect 163 1734 2647 1825
rect 2958 1781 3381 1813
rect 3437 1745 3900 1899
rect 163 1695 2501 1734
rect 2279 1581 2360 1599
rect 2279 1529 2298 1581
rect 2350 1529 2360 1581
rect 2279 1510 2360 1529
rect 2556 1341 2647 1734
rect 3020 1391 3109 1407
rect 2556 1250 2803 1341
rect 3020 1339 3037 1391
rect 3089 1339 3109 1391
rect 3517 1388 3615 1415
rect 3020 1325 3109 1339
rect 3467 1385 3615 1388
rect 3467 1333 3535 1385
rect 3587 1333 3615 1385
rect 3467 1319 3615 1333
rect 3517 1299 3615 1319
rect 249 1031 336 1054
rect -28 1026 336 1031
rect -28 980 271 1026
rect 317 980 336 1026
rect -28 958 336 980
rect 2712 967 2803 1250
rect 249 951 336 958
rect 2964 963 2968 970
rect 2964 930 3375 963
rect 2968 929 3375 930
rect 1548 750 1618 754
rect 1548 739 1619 750
rect 1548 687 1557 739
rect 1609 687 1619 739
rect 1548 680 1619 687
rect 3593 549 3700 578
rect 2743 519 2843 546
rect 2743 467 2766 519
rect 2818 467 2843 519
rect 2743 453 2843 467
rect 3593 497 3619 549
rect 3671 514 3700 549
rect 3671 497 3712 514
rect 3593 463 3712 497
rect 3663 427 3712 463
rect 133 141 3682 205
rect 3758 141 3900 1745
rect 133 46 3900 141
rect 133 0 911 46
rect 1803 0 3900 46
rect 133 -69 3900 0
rect 133 -113 3682 -69
<< via1 >>
rect 2770 3077 2822 3129
rect 3649 3106 3701 3158
rect 1554 2988 1606 3040
rect 535 2143 587 2195
rect 2302 2146 2354 2198
rect 3035 2191 3087 2243
rect 3502 2210 3554 2262
rect 2298 1529 2350 1581
rect 3037 1339 3089 1391
rect 3535 1333 3587 1385
rect 1557 687 1609 739
rect 2766 467 2818 519
rect 3619 497 3671 549
<< metal2 >>
rect 3634 3176 3720 3178
rect 3634 3158 3981 3176
rect 2744 3132 2835 3142
rect 2598 3129 2835 3132
rect 2598 3077 2770 3129
rect 2822 3077 2835 3129
rect 3634 3106 3649 3158
rect 3701 3106 3981 3158
rect 3634 3090 3981 3106
rect 3634 3088 3720 3090
rect 2598 3075 2835 3077
rect 1538 3045 1625 3053
rect 1536 3042 1625 3045
rect 1536 2986 1553 3042
rect 1609 2986 1625 3042
rect 1536 2975 1625 2986
rect 1979 3046 2062 3061
rect 1979 2990 1994 3046
rect 2050 2990 2062 3046
rect 1979 2977 2062 2990
rect 2598 2590 2655 3075
rect 2744 3062 2835 3075
rect 2472 2533 2655 2590
rect 2736 2396 3900 2488
rect 520 2195 598 2211
rect 2291 2207 2367 2211
rect 2736 2207 2828 2396
rect 520 2143 535 2195
rect 587 2143 598 2195
rect 520 2125 598 2143
rect 2286 2200 2828 2207
rect 2286 2144 2301 2200
rect 2357 2144 2828 2200
rect 3012 2247 3107 2265
rect 3012 2191 3034 2247
rect 3090 2191 3107 2247
rect 3012 2175 3107 2191
rect 3489 2262 3575 2283
rect 3489 2210 3502 2262
rect 3554 2210 3575 2262
rect 3489 2188 3575 2210
rect 534 1901 590 2125
rect 2286 2115 2828 2144
rect 3511 1790 3569 2188
rect 2579 1732 3569 1790
rect 2278 1583 2372 1603
rect 2278 1527 2296 1583
rect 2352 1527 2372 1583
rect 2278 1517 2372 1527
rect 3015 1395 3116 1415
rect 3015 1339 3036 1395
rect 3092 1339 3116 1395
rect 3015 1321 3116 1339
rect 3517 1408 3615 1415
rect 3822 1408 3900 2396
rect 3517 1385 3900 1408
rect 3517 1333 3535 1385
rect 3587 1333 3900 1385
rect 3517 1316 3900 1333
rect 3517 1299 3615 1316
rect 1541 741 1626 755
rect 1541 685 1555 741
rect 1611 685 1626 741
rect 1541 676 1626 685
rect 1985 740 2065 752
rect 1985 684 1997 740
rect 2053 684 2065 740
rect 1985 675 2065 684
rect 2722 580 2836 645
rect 2741 546 2836 580
rect 3593 549 4062 578
rect 2741 543 2843 546
rect 2743 519 2843 543
rect 2743 467 2766 519
rect 2818 467 2843 519
rect 2743 453 2843 467
rect 3593 497 3619 549
rect 3671 497 4062 549
rect 3593 463 4062 497
<< via2 >>
rect 1553 3040 1609 3042
rect 1553 2988 1554 3040
rect 1554 2988 1606 3040
rect 1606 2988 1609 3040
rect 1553 2986 1609 2988
rect 1994 2990 2050 3046
rect 2301 2198 2357 2200
rect 2301 2146 2302 2198
rect 2302 2146 2354 2198
rect 2354 2146 2357 2198
rect 2301 2144 2357 2146
rect 3034 2243 3090 2247
rect 3034 2191 3035 2243
rect 3035 2191 3087 2243
rect 3087 2191 3090 2243
rect 2296 1581 2352 1583
rect 2296 1529 2298 1581
rect 2298 1529 2350 1581
rect 2350 1529 2352 1581
rect 2296 1527 2352 1529
rect 3036 1391 3092 1395
rect 3036 1339 3037 1391
rect 3037 1339 3089 1391
rect 3089 1339 3092 1391
rect 1555 739 1611 741
rect 1555 687 1557 739
rect 1557 687 1609 739
rect 1609 687 1611 739
rect 1555 685 1611 687
rect 1997 684 2053 740
<< metal3 >>
rect 1245 3187 2041 3255
rect 1245 1176 1313 3187
rect 1973 3061 2041 3187
rect 1538 3042 1625 3053
rect 1538 2986 1553 3042
rect 1609 2986 1625 3042
rect 1973 3046 2062 3061
rect 1973 2990 1994 3046
rect 2050 2990 2062 3046
rect 1538 2975 1625 2986
rect 1979 2977 2062 2990
rect 1546 2348 1618 2975
rect 1546 2276 3107 2348
rect 1546 1623 1618 2276
rect 2988 2247 3107 2276
rect 2287 2200 2374 2214
rect 2287 2181 2301 2200
rect 2278 2144 2301 2181
rect 2357 2144 2374 2200
rect 2988 2191 3034 2247
rect 3090 2191 3107 2247
rect 2988 2164 3107 2191
rect 2278 2133 2374 2144
rect 1546 1551 2043 1623
rect 2278 1608 2372 2133
rect 1245 1108 1619 1176
rect 1551 755 1619 1108
rect 1971 755 2043 1551
rect 2274 1583 2372 1608
rect 2274 1527 2296 1583
rect 2352 1527 2372 1583
rect 2274 1517 2372 1527
rect 2274 1503 2370 1517
rect 2436 1415 3053 1418
rect 2436 1395 3116 1415
rect 2436 1350 3036 1395
rect 1541 741 1626 755
rect 1541 685 1555 741
rect 1611 685 1626 741
rect 1541 676 1626 685
rect 1971 740 2067 755
rect 1971 684 1997 740
rect 2053 684 2067 740
rect 1551 614 1623 676
rect 1971 671 2067 684
rect 1971 664 2043 671
rect 1551 468 1619 614
rect 2436 468 2504 1350
rect 3015 1339 3036 1350
rect 3092 1339 3116 1395
rect 3015 1321 3116 1339
rect 1551 400 2504 468
use Buffer_V_2  Buffer_V_2_0
timestamp 1713185578
transform 1 0 2622 0 -1 532
box -8 -438 1070 535
use Buffer_V_2  Buffer_V_2_1
timestamp 1713185578
transform 1 0 2621 0 1 3070
box -8 -438 1070 535
use INV_mag  INV_mag_0
timestamp 1713185578
transform 1 0 2855 0 -1 2261
box 0 -400 652 485
use INV_mag  INV_mag_1
timestamp 1713185578
transform 1 0 2855 0 1 1321
box 0 -400 652 485
use PFD_2  PFD_2_0
timestamp 1713185578
transform 1 0 133 0 1 3063
box -45 -1176 2616 545
use PFD_2_down  PFD_2_down_0
timestamp 1713185578
transform 1 0 134 0 -1 664
box -45 -1251 2616 545
<< labels >>
flabel nsubdiffcont 1357 24 1357 24 0 FreeSans 2500 0 0 0 VDD
flabel psubdiffcont 1308 1883 1308 1883 0 FreeSans 2500 0 0 0 VSS
flabel metal1 s 57 2733 57 2733 0 FreeSans 2500 0 0 0 FIN
port 1 nsew
flabel metal1 s 20 1007 20 1007 0 FreeSans 2500 0 0 0 FDIV
port 2 nsew
flabel metal1 s 3702 3130 3702 3130 0 FreeSans 2500 0 0 0 UP
port 3 nsew
flabel metal1 s 3692 488 3692 488 0 FreeSans 2500 0 0 0 DOWN
port 4 nsew
<< end >>
