** sch_path: /home/shahid/GF180Projects/CP_PFD_dff_inv_nand_/Xschem/RES/pex_res_sch_test.sch
**.subckt pex_res_sch_test
x1 A B VDD pex_res_sch48new
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
* .lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_statistical



vp a 0 0
vm b 0 0
vb vdd 0 3.3
.include pex_res_48k_lay.spice
.control
save all
dc vp 0 3.3 0.01
write pex_res_sch_test.raw
.endc


**** end user architecture code
**.ends
.end
