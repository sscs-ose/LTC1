magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2180 -2535 2180 2535
<< metal2 >>
rect -180 525 180 535
rect -180 469 -170 525
rect -114 469 -28 525
rect 28 469 114 525
rect 170 469 180 525
rect -180 383 180 469
rect -180 327 -170 383
rect -114 327 -28 383
rect 28 327 114 383
rect 170 327 180 383
rect -180 241 180 327
rect -180 185 -170 241
rect -114 185 -28 241
rect 28 185 114 241
rect 170 185 180 241
rect -180 99 180 185
rect -180 43 -170 99
rect -114 43 -28 99
rect 28 43 114 99
rect 170 43 180 99
rect -180 -43 180 43
rect -180 -99 -170 -43
rect -114 -99 -28 -43
rect 28 -99 114 -43
rect 170 -99 180 -43
rect -180 -185 180 -99
rect -180 -241 -170 -185
rect -114 -241 -28 -185
rect 28 -241 114 -185
rect 170 -241 180 -185
rect -180 -327 180 -241
rect -180 -383 -170 -327
rect -114 -383 -28 -327
rect 28 -383 114 -327
rect 170 -383 180 -327
rect -180 -469 180 -383
rect -180 -525 -170 -469
rect -114 -525 -28 -469
rect 28 -525 114 -469
rect 170 -525 180 -469
rect -180 -535 180 -525
<< via2 >>
rect -170 469 -114 525
rect -28 469 28 525
rect 114 469 170 525
rect -170 327 -114 383
rect -28 327 28 383
rect 114 327 170 383
rect -170 185 -114 241
rect -28 185 28 241
rect 114 185 170 241
rect -170 43 -114 99
rect -28 43 28 99
rect 114 43 170 99
rect -170 -99 -114 -43
rect -28 -99 28 -43
rect 114 -99 170 -43
rect -170 -241 -114 -185
rect -28 -241 28 -185
rect 114 -241 170 -185
rect -170 -383 -114 -327
rect -28 -383 28 -327
rect 114 -383 170 -327
rect -170 -525 -114 -469
rect -28 -525 28 -469
rect 114 -525 170 -469
<< metal3 >>
rect -180 525 180 535
rect -180 469 -170 525
rect -114 469 -28 525
rect 28 469 114 525
rect 170 469 180 525
rect -180 383 180 469
rect -180 327 -170 383
rect -114 327 -28 383
rect 28 327 114 383
rect 170 327 180 383
rect -180 241 180 327
rect -180 185 -170 241
rect -114 185 -28 241
rect 28 185 114 241
rect 170 185 180 241
rect -180 99 180 185
rect -180 43 -170 99
rect -114 43 -28 99
rect 28 43 114 99
rect 170 43 180 99
rect -180 -43 180 43
rect -180 -99 -170 -43
rect -114 -99 -28 -43
rect 28 -99 114 -43
rect 170 -99 180 -43
rect -180 -185 180 -99
rect -180 -241 -170 -185
rect -114 -241 -28 -185
rect 28 -241 114 -185
rect 170 -241 180 -185
rect -180 -327 180 -241
rect -180 -383 -170 -327
rect -114 -383 -28 -327
rect 28 -383 114 -327
rect 170 -383 180 -327
rect -180 -469 180 -383
rect -180 -525 -170 -469
rect -114 -525 -28 -469
rect 28 -525 114 -469
rect 170 -525 180 -469
rect -180 -535 180 -525
<< end >>
