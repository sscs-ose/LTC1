magic
tech gf180mcuC
magscale 1 10
timestamp 1693483190
<< metal1 >>
rect 228 2374 4815 2538
rect 426 2113 482 2181
rect 412 2100 491 2113
rect 412 2048 425 2100
rect 478 2048 491 2100
rect -2788 2036 -2701 2044
rect 412 2036 491 2048
rect -2788 1964 -2546 2036
rect -2156 1975 -2079 1985
rect -2788 -181 -2701 1964
rect -2156 1918 -2145 1975
rect -2089 1918 -2079 1975
rect 2348 1935 2394 2089
rect -2156 1906 -2079 1918
rect 795 1908 865 1920
rect 795 1856 807 1908
rect 859 1856 865 1908
rect 4869 1914 5030 1929
rect 620 1839 693 1855
rect 795 1851 865 1856
rect 1440 1862 1508 1876
rect 620 1787 634 1839
rect 686 1787 693 1839
rect 1440 1806 1443 1862
rect 1495 1806 1508 1862
rect 4869 1862 4873 1914
rect 4926 1862 5030 1914
rect 4869 1847 5030 1862
rect 1440 1791 1508 1806
rect 620 1776 693 1787
rect 1441 1612 1882 1716
rect 1441 1501 1545 1612
rect 1595 1524 1686 1543
rect 1595 1468 1611 1524
rect 1669 1468 1686 1524
rect 1595 1453 1686 1468
rect 430 1417 512 1427
rect 919 1417 1001 1432
rect 430 1412 945 1417
rect -2636 1363 -2483 1367
rect -2636 1308 -2552 1363
rect -2498 1308 -2483 1363
rect 430 1358 456 1412
rect 508 1363 945 1412
rect 997 1363 1001 1417
rect 508 1358 1001 1363
rect 430 1353 1001 1358
rect 1947 1423 2024 1439
rect 1947 1367 1958 1423
rect 2014 1367 2024 1423
rect 1947 1356 2024 1367
rect 430 1345 512 1353
rect 919 1350 1001 1353
rect -2636 1303 -2483 1308
rect -2636 193 -2572 1303
rect 231 1259 968 1277
rect 208 1202 968 1259
rect 231 1183 968 1202
rect -1145 986 -1061 987
rect -1145 984 -1045 986
rect -1145 926 -1128 984
rect -1072 926 -1045 984
rect -2507 886 -2429 902
rect -2507 839 -2494 886
rect -2509 833 -2494 839
rect -2441 833 -2429 886
rect -2509 823 -2429 833
rect -2162 885 -2060 897
rect -2162 833 -2150 885
rect -2097 833 -2060 885
rect 381 884 463 899
rect 381 880 396 884
rect -2509 363 -2438 823
rect -2162 821 -2060 833
rect 356 829 396 880
rect 451 880 463 884
rect 451 829 471 880
rect 356 825 471 829
rect 381 823 463 825
rect 1197 702 1310 712
rect 624 648 712 658
rect 1197 650 1210 702
rect 1262 650 1310 702
rect 1197 649 1310 650
rect 624 640 1064 648
rect 624 586 644 640
rect 696 586 1064 640
rect 624 577 1064 586
rect 624 566 712 577
rect 341 399 608 487
rect 1849 452 1902 465
rect 1849 438 1850 452
rect 1836 400 1850 438
rect 341 368 929 399
rect 1836 387 1902 400
rect -2522 343 -2438 363
rect -2522 291 -2509 343
rect -2456 291 -2438 343
rect -2522 286 -2438 291
rect 489 280 929 368
rect 1948 273 2017 1356
rect 3318 934 3418 937
rect 3318 876 3337 934
rect 3393 876 3418 934
rect 2301 844 2412 856
rect 2301 792 2314 844
rect 2366 792 2412 844
rect 4949 830 5025 836
rect 2301 780 2412 792
rect 4823 824 5025 830
rect 4823 775 4961 824
rect 4949 772 4961 775
rect 5013 772 5025 824
rect 4949 760 5025 772
rect 4743 331 5463 450
rect 1948 207 3156 273
rect 463 195 535 205
rect 1197 195 1274 206
rect 463 193 1274 195
rect 463 189 1210 193
rect 463 136 475 189
rect 528 140 1210 189
rect 1263 140 1274 193
rect 528 136 1274 140
rect 463 130 1274 136
rect 463 124 535 130
rect 1197 127 1274 130
rect 1692 -58 1918 76
rect 609 -141 688 -133
rect 1379 -141 1461 -135
rect 517 -148 1461 -141
rect -3248 -268 -2565 -181
rect 517 -203 623 -148
rect 677 -149 1461 -148
rect 677 -202 1393 -149
rect 1446 -202 1461 -149
rect 677 -203 1461 -202
rect 517 -211 1461 -203
rect 517 -225 773 -211
rect 1379 -215 1461 -211
rect -2159 -248 -2094 -243
rect -2159 -300 -2147 -248
rect -2095 -300 -2094 -248
rect -2159 -322 -2094 -300
rect -2914 -488 -2631 -466
rect -2914 -542 -2897 -488
rect -2842 -542 -2631 -488
rect -2914 -556 -2631 -542
rect -2755 -1226 -2598 -1211
rect -2755 -1285 -2670 -1226
rect -2612 -1285 -2598 -1226
rect -2755 -1297 -2598 -1285
rect -1161 -1243 -1062 -1241
rect -1161 -1301 -1141 -1243
rect -1085 -1301 -1062 -1243
rect 517 -1328 584 -225
rect 653 -718 901 -679
rect 653 -770 682 -718
rect 734 -770 901 -718
rect 653 -801 901 -770
rect 1692 -970 1826 -58
rect 3090 -177 3156 207
rect 3748 105 4355 258
rect 4237 85 4355 105
rect 4237 22 4356 85
rect 5344 41 5463 331
rect 3090 -243 3410 -177
rect 3746 -240 4043 -182
rect 2850 -435 3089 -427
rect 1982 -469 2081 -467
rect 1982 -521 1995 -469
rect 2047 -521 2081 -469
rect 2850 -487 3025 -435
rect 3077 -487 3089 -435
rect 2850 -488 3089 -487
rect 1982 -530 2081 -521
rect 3173 -550 3409 -441
rect 3985 -537 4043 -240
rect 4955 -537 5021 -359
rect 3173 -683 3282 -550
rect 3985 -595 5022 -537
rect 4955 -599 5021 -595
rect 2813 -792 3282 -683
rect 1163 -1263 1253 -1262
rect 1163 -1316 1182 -1263
rect 1237 -1316 1253 -1263
rect 1163 -1320 1253 -1316
rect -2176 -1335 -2030 -1330
rect -2176 -1388 -2164 -1335
rect -2111 -1388 -2030 -1335
rect 363 -1346 442 -1333
rect 363 -1348 375 -1346
rect -2176 -1400 -2030 -1388
rect 342 -1400 375 -1348
rect 430 -1400 442 -1346
rect 517 -1395 1068 -1328
rect 1787 -1367 1978 -1310
rect 342 -1403 442 -1400
rect 363 -1412 442 -1403
rect 2122 -1565 2231 -890
rect 854 -1740 1005 -1635
rect 1805 -1674 2231 -1565
rect 2708 -1258 2726 -1204
rect 2780 -1258 2797 -1204
rect 257 -1848 1006 -1740
rect 2708 -1825 2797 -1258
rect 2967 -1644 3076 -792
rect 3212 -1230 3294 -1221
rect 3212 -1236 3615 -1230
rect 3212 -1288 3227 -1236
rect 3280 -1288 3615 -1236
rect 4286 -1271 4533 -1182
rect 3212 -1302 3615 -1288
rect 2967 -1753 3452 -1644
rect 4444 -1825 4533 -1271
rect 2708 -1914 4533 -1825
<< via1 >>
rect 425 2048 478 2100
rect -2145 1918 -2089 1975
rect 807 1856 859 1908
rect 634 1787 686 1839
rect 1443 1806 1495 1862
rect 4873 1862 4926 1914
rect -2359 1508 -2304 1564
rect 1611 1468 1669 1524
rect -2552 1308 -2498 1363
rect -2193 1309 -2139 1364
rect 456 1358 508 1412
rect 945 1363 997 1417
rect 1958 1367 2014 1423
rect -1128 926 -1072 984
rect -2494 833 -2441 886
rect -2150 833 -2097 885
rect 396 829 451 884
rect 1210 650 1262 702
rect 644 586 696 640
rect 1803 607 1855 659
rect 1850 400 1902 452
rect -2509 291 -2456 343
rect 3337 876 3393 934
rect 2314 792 2366 844
rect 4961 772 5013 824
rect 2116 400 2168 452
rect 475 136 528 189
rect 1210 140 1263 193
rect 623 -203 677 -148
rect 1393 -202 1446 -149
rect -2147 -300 -2095 -248
rect -2897 -542 -2842 -488
rect 281 -775 333 -723
rect -2670 -1285 -2612 -1226
rect -1141 -1301 -1085 -1243
rect 682 -770 734 -718
rect 2799 -61 2852 -8
rect 3372 177 3425 230
rect 5105 62 5158 115
rect 4959 -59 5011 -7
rect 4959 -199 5011 -147
rect 2310 -430 2362 -378
rect 1995 -521 2047 -469
rect 3025 -487 3077 -435
rect 1182 -1316 1237 -1263
rect -2164 -1388 -2111 -1335
rect 375 -1400 430 -1346
rect 2726 -1258 2780 -1204
rect 3429 -825 3486 -768
rect 3799 -1201 3852 -1148
rect 3227 -1288 3280 -1236
<< metal2 >>
rect -2610 2317 1695 2399
rect -2610 2099 -2528 2317
rect 412 2100 491 2113
rect -2610 2049 -2455 2099
rect -2610 1967 -2418 2049
rect 412 2048 425 2100
rect 478 2048 491 2100
rect 412 2036 491 2048
rect -2156 1975 -2079 1985
rect -2156 1918 -2145 1975
rect -2089 1918 -2079 1975
rect 420 1966 483 2036
rect -2156 1906 -2079 1918
rect 170 1903 483 1966
rect 1613 1996 1695 2317
rect 795 1908 865 1920
rect 1613 1915 2032 1996
rect 4856 1918 4939 1929
rect -2914 1574 -2824 1583
rect -2368 1574 -2295 1580
rect -2914 1564 -2295 1574
rect -2914 1508 -2359 1564
rect -2304 1508 -2295 1564
rect -2914 1502 -2295 1508
rect -2914 -488 -2824 1502
rect -2368 1497 -2295 1502
rect 311 1419 374 1903
rect 795 1856 807 1908
rect 859 1856 865 1908
rect 4637 1914 4939 1918
rect 620 1839 693 1855
rect 795 1851 865 1856
rect 1433 1862 1515 1880
rect 620 1787 634 1839
rect 686 1815 693 1839
rect 686 1787 702 1815
rect 620 1776 702 1787
rect 430 1419 512 1428
rect 311 1412 512 1419
rect -2215 1383 -2118 1384
rect -2559 1364 -2118 1383
rect -2559 1363 -2193 1364
rect -2559 1308 -2552 1363
rect -2498 1309 -2193 1363
rect -2139 1309 -2118 1364
rect 311 1358 456 1412
rect 508 1358 512 1412
rect 311 1356 512 1358
rect 430 1345 512 1356
rect -2498 1308 -2118 1309
rect -2559 1287 -2118 1308
rect -2559 1283 -2200 1287
rect -1145 984 -1054 994
rect -1145 926 -1128 984
rect -1072 926 -1054 984
rect -1145 914 -1054 926
rect -2507 897 -2430 901
rect -2507 886 -2060 897
rect 381 890 463 899
rect 635 890 702 1776
rect -2507 833 -2494 886
rect -2441 885 -2060 886
rect -2441 833 -2150 885
rect -2097 833 -2060 885
rect -2507 824 -2060 833
rect -2507 823 -2430 824
rect -2171 821 -2060 824
rect 328 884 702 890
rect 328 829 396 884
rect 451 829 702 884
rect 328 823 702 829
rect -2171 820 -2061 821
rect -2767 588 -1469 646
rect 624 640 712 658
rect -2767 -321 -2709 588
rect 624 586 644 640
rect 696 586 712 640
rect 624 566 712 586
rect 623 431 681 566
rect -2522 351 -2438 356
rect -2522 343 286 351
rect -2522 291 -2509 343
rect -2456 291 286 343
rect -2522 285 286 291
rect -2522 279 -2438 285
rect 220 194 286 285
rect 463 194 535 205
rect 220 189 535 194
rect 220 136 475 189
rect 528 136 535 189
rect 220 128 535 136
rect 463 124 535 128
rect 624 -133 680 431
rect 609 -148 688 -133
rect 609 -203 623 -148
rect 677 -203 688 -148
rect 609 -216 688 -203
rect -2116 -243 -2051 -242
rect -2181 -248 -2051 -243
rect -2181 -300 -2147 -248
rect -2095 -300 -2051 -248
rect 609 -266 680 -216
rect -2181 -321 -2051 -300
rect -2767 -379 -2093 -321
rect 102 -322 680 -266
rect -2914 -542 -2897 -488
rect -2842 -542 -2824 -488
rect -2914 -554 -2824 -542
rect 266 -712 336 -711
rect 653 -712 740 -697
rect 266 -718 740 -712
rect 266 -723 682 -718
rect 266 -775 281 -723
rect 333 -770 682 -723
rect 734 -770 740 -718
rect 333 -775 740 -770
rect 266 -786 336 -775
rect 653 -792 740 -775
rect -2686 -1226 -2597 -1190
rect -2686 -1285 -2670 -1226
rect -2612 -1285 -2597 -1226
rect -1144 -1229 -1072 -1223
rect -2686 -1306 -2597 -1285
rect -1161 -1243 -1072 -1229
rect -1161 -1301 -1141 -1243
rect -1085 -1301 -1072 -1243
rect -1161 -1314 -1072 -1301
rect -2385 -1335 -2030 -1329
rect -2385 -1388 -2164 -1335
rect -2111 -1388 -2030 -1335
rect 363 -1341 442 -1333
rect 796 -1341 859 1851
rect 1433 1806 1443 1862
rect 1495 1858 1515 1862
rect 4637 1862 4873 1914
rect 4926 1862 4939 1914
rect 1808 1858 1878 1859
rect 1495 1806 1878 1858
rect 4637 1855 4939 1862
rect 4856 1847 4939 1855
rect 1433 1788 1878 1806
rect 1595 1524 1686 1543
rect 1595 1468 1611 1524
rect 1669 1468 1686 1524
rect 1595 1453 1686 1468
rect 919 1417 1001 1433
rect 919 1363 945 1417
rect 997 1363 1001 1417
rect 919 1350 1001 1363
rect 926 1302 996 1350
rect 927 -587 995 1302
rect 1595 1139 1659 1453
rect 1808 1287 1878 1788
rect 1947 1435 2025 1440
rect 1947 1423 2666 1435
rect 1947 1367 1958 1423
rect 2014 1367 2666 1423
rect 1947 1362 2666 1367
rect 1947 1356 2025 1362
rect 1808 1217 2305 1287
rect 1595 1075 1861 1139
rect 1189 702 1274 722
rect 1189 650 1210 702
rect 1262 650 1274 702
rect 1797 682 1861 1075
rect 2235 856 2305 1217
rect 3327 934 3404 945
rect 3327 876 3337 934
rect 3393 876 3404 934
rect 3327 864 3404 876
rect 2235 844 2412 856
rect 2235 792 2314 844
rect 2366 792 2412 844
rect 2235 782 2412 792
rect 2301 780 2412 782
rect 4949 824 5025 836
rect 4949 772 4961 824
rect 5013 772 5025 824
rect 4949 760 5025 772
rect 1189 629 1274 650
rect 1782 659 1873 682
rect 1194 616 1269 629
rect 1206 335 1269 616
rect 1782 607 1803 659
rect 1855 607 1873 659
rect 1782 591 1873 607
rect 1838 452 2177 465
rect 1838 400 1850 452
rect 1902 400 2116 452
rect 2168 400 2177 452
rect 1838 392 2177 400
rect 2942 335 3008 594
rect 1206 269 3008 335
rect 1206 206 1269 269
rect 3366 233 3435 251
rect 1197 193 1274 206
rect 1197 140 1210 193
rect 1263 140 1274 193
rect 1197 127 1274 140
rect 3366 177 3370 233
rect 3426 177 3435 233
rect 1206 -466 1269 127
rect 3366 1 3435 177
rect 4957 9 5016 760
rect 5091 115 5171 124
rect 5091 62 5105 115
rect 5158 62 5171 115
rect 2786 -8 3435 1
rect 2786 -61 2799 -8
rect 2852 -61 3435 -8
rect 2786 -68 3435 -61
rect 4946 -7 5024 9
rect 4946 -59 4959 -7
rect 5011 -59 5024 -7
rect 2786 -70 2906 -68
rect 4946 -73 5024 -59
rect 1379 -141 1461 -135
rect 4947 -141 5022 -134
rect 1379 -147 5022 -141
rect 1379 -149 4959 -147
rect 1379 -202 1393 -149
rect 1446 -199 4959 -149
rect 5011 -199 5022 -147
rect 1446 -202 5022 -199
rect 1379 -210 5022 -202
rect 1379 -215 1461 -210
rect 4947 -215 5022 -210
rect 2439 -347 3295 -270
rect 2294 -370 2376 -366
rect 2439 -370 2517 -347
rect 2294 -378 2517 -370
rect 2294 -430 2310 -378
rect 2362 -430 2517 -378
rect 2294 -442 2517 -430
rect 2301 -448 2517 -442
rect 2964 -427 3031 -425
rect 2964 -435 3089 -427
rect 1206 -467 2079 -466
rect 1206 -469 2081 -467
rect 1206 -521 1995 -469
rect 2047 -521 2081 -469
rect 1206 -529 2081 -521
rect 1982 -530 2081 -529
rect 2301 -587 2369 -448
rect 927 -655 2369 -587
rect 2964 -487 3025 -435
rect 3077 -487 3089 -435
rect 2964 -488 3089 -487
rect 1164 -1204 2797 -1189
rect 1164 -1249 2726 -1204
rect 1162 -1250 2726 -1249
rect 1162 -1263 1254 -1250
rect 2708 -1258 2726 -1250
rect 2780 -1258 2797 -1204
rect 2708 -1261 2797 -1258
rect 1162 -1316 1182 -1263
rect 1237 -1316 1254 -1263
rect 1162 -1326 1254 -1316
rect -2385 -1412 -2030 -1388
rect 319 -1346 859 -1341
rect 319 -1400 375 -1346
rect 430 -1400 859 -1346
rect 319 -1404 859 -1400
rect 363 -1412 442 -1404
rect -2385 -1802 -2261 -1412
rect 2964 -1802 3085 -488
rect 3212 -1224 3295 -347
rect 5091 -589 5171 62
rect 3783 -669 5171 -589
rect 3405 -768 3505 -755
rect 3405 -825 3429 -768
rect 3486 -825 3505 -768
rect 3405 -845 3505 -825
rect 3783 -1130 3863 -669
rect 3783 -1148 3868 -1130
rect 3783 -1201 3799 -1148
rect 3852 -1201 3868 -1148
rect 3783 -1218 3868 -1201
rect 3212 -1236 3294 -1224
rect 3212 -1288 3227 -1236
rect 3280 -1288 3294 -1236
rect 3212 -1302 3294 -1288
rect -2385 -1944 3085 -1802
rect -2385 -1946 -2261 -1944
<< via2 >>
rect -2145 1918 -2089 1975
rect -1128 926 -1072 984
rect -2670 -1285 -2612 -1226
rect -1141 -1301 -1085 -1243
rect 1611 1468 1669 1524
rect 3337 876 3393 934
rect 3370 230 3426 233
rect 3370 177 3372 230
rect 3372 177 3425 230
rect 3425 177 3426 230
rect 3429 -825 3486 -768
<< metal3 >>
rect -2156 1975 1695 2001
rect -2156 1918 -2145 1975
rect -2089 1918 1695 1975
rect -2156 1892 1695 1918
rect 1586 1524 1695 1892
rect 1586 1468 1611 1524
rect 1669 1468 1695 1524
rect 1586 1447 1695 1468
rect -1140 984 -1045 994
rect -1140 926 -1128 984
rect -1072 953 -1045 984
rect -1072 945 3339 953
rect -1072 934 3404 945
rect -1072 926 3337 934
rect -1140 876 3337 926
rect 3393 876 3404 934
rect -1140 866 3404 876
rect -1144 864 3404 866
rect -1144 852 3339 864
rect -1144 -1189 -1042 852
rect 3352 233 3442 251
rect 3352 177 3370 233
rect 3426 207 3442 233
rect 3426 177 3443 207
rect 3352 154 3443 177
rect 3353 -755 3443 154
rect 3353 -768 3505 -755
rect 3353 -825 3429 -768
rect 3486 -825 3505 -768
rect 3353 -845 3505 -825
rect -2680 -1190 -1042 -1189
rect -2686 -1226 -1042 -1190
rect -2686 -1285 -2670 -1226
rect -2612 -1243 -1042 -1226
rect -2612 -1285 -1141 -1243
rect -2686 -1301 -1141 -1285
rect -1085 -1301 -1042 -1243
rect -2686 -1306 -1042 -1301
rect -2680 -1307 -1042 -1306
rect -1144 -1314 -1042 -1307
use and2_mag  and2_mag_0
timestamp 1692973937
transform 1 0 3471 0 1 -1564
box -70 -188 906 863
use and2_mag  and2_mag_1
timestamp 1692973937
transform 1 0 1950 0 1 -792
box -70 -188 906 863
use GF_INV_MAG  GF_INV_MAG_0
timestamp 1692973937
transform 1 0 3480 0 1 -371
box -118 -175 286 631
use JK_FF_mag  JK_FF_mag_0
timestamp 1692973937
transform 1 0 -2244 0 1 -1850
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_1
timestamp 1692973937
transform 1 0 2235 0 1 328
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_2
timestamp 1692973937
transform 1 0 -2228 0 1 378
box -390 0 2603 2148
use nor_3_mag  nor_3_mag_0
timestamp 1692973937
transform 0 -1 5902 1 0 -856
box 329 440 1054 1778
use or_2_mag  or_2_mag_1
timestamp 1692973937
transform 1 0 174 0 1 968
box 330 510 1298 1521
use or_2_mag  or_2_mag_2
timestamp 1692973937
transform 1 0 590 0 1 -230
box 330 510 1298 1521
use or_2_mag  or_2_mag_3
timestamp 1692973937
transform 1 0 527 0 1 -2204
box 330 510 1298 1521
<< labels >>
flabel metal1 604 -1771 604 -1771 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal1 1152 2472 1152 2472 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 4983 1886 4983 1886 0 FreeSans 1600 0 0 0 Q0
port 2 nsew
flabel metal1 452 2166 452 2166 0 FreeSans 1600 0 0 0 Q1
port 3 nsew
flabel metal1 539 -197 539 -197 0 FreeSans 1600 0 0 0 Q2
port 4 nsew
flabel metal1 -2723 -1252 -2723 -1252 0 FreeSans 1600 0 0 0 RST
port 5 nsew
flabel metal1 -3205 -230 -3205 -230 0 FreeSans 1600 0 0 0 CLK
port 10 nsew
flabel metal1 1930 -1340 1930 -1340 0 FreeSans 1600 0 0 0 Vdiv7
port 11 nsew
<< end >>
