magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1217 -1910 1217 1910
<< metal1 >>
rect -217 904 217 910
rect -217 878 -211 904
rect -185 878 -145 904
rect -119 878 -79 904
rect -53 878 -13 904
rect 13 878 53 904
rect 79 878 119 904
rect 145 878 185 904
rect 211 878 217 904
rect -217 838 217 878
rect -217 812 -211 838
rect -185 812 -145 838
rect -119 812 -79 838
rect -53 812 -13 838
rect 13 812 53 838
rect 79 812 119 838
rect 145 812 185 838
rect 211 812 217 838
rect -217 772 217 812
rect -217 746 -211 772
rect -185 746 -145 772
rect -119 746 -79 772
rect -53 746 -13 772
rect 13 746 53 772
rect 79 746 119 772
rect 145 746 185 772
rect 211 746 217 772
rect -217 706 217 746
rect -217 680 -211 706
rect -185 680 -145 706
rect -119 680 -79 706
rect -53 680 -13 706
rect 13 680 53 706
rect 79 680 119 706
rect 145 680 185 706
rect 211 680 217 706
rect -217 640 217 680
rect -217 614 -211 640
rect -185 614 -145 640
rect -119 614 -79 640
rect -53 614 -13 640
rect 13 614 53 640
rect 79 614 119 640
rect 145 614 185 640
rect 211 614 217 640
rect -217 574 217 614
rect -217 548 -211 574
rect -185 548 -145 574
rect -119 548 -79 574
rect -53 548 -13 574
rect 13 548 53 574
rect 79 548 119 574
rect 145 548 185 574
rect 211 548 217 574
rect -217 508 217 548
rect -217 482 -211 508
rect -185 482 -145 508
rect -119 482 -79 508
rect -53 482 -13 508
rect 13 482 53 508
rect 79 482 119 508
rect 145 482 185 508
rect 211 482 217 508
rect -217 442 217 482
rect -217 416 -211 442
rect -185 416 -145 442
rect -119 416 -79 442
rect -53 416 -13 442
rect 13 416 53 442
rect 79 416 119 442
rect 145 416 185 442
rect 211 416 217 442
rect -217 376 217 416
rect -217 350 -211 376
rect -185 350 -145 376
rect -119 350 -79 376
rect -53 350 -13 376
rect 13 350 53 376
rect 79 350 119 376
rect 145 350 185 376
rect 211 350 217 376
rect -217 310 217 350
rect -217 284 -211 310
rect -185 284 -145 310
rect -119 284 -79 310
rect -53 284 -13 310
rect 13 284 53 310
rect 79 284 119 310
rect 145 284 185 310
rect 211 284 217 310
rect -217 244 217 284
rect -217 218 -211 244
rect -185 218 -145 244
rect -119 218 -79 244
rect -53 218 -13 244
rect 13 218 53 244
rect 79 218 119 244
rect 145 218 185 244
rect 211 218 217 244
rect -217 178 217 218
rect -217 152 -211 178
rect -185 152 -145 178
rect -119 152 -79 178
rect -53 152 -13 178
rect 13 152 53 178
rect 79 152 119 178
rect 145 152 185 178
rect 211 152 217 178
rect -217 112 217 152
rect -217 86 -211 112
rect -185 86 -145 112
rect -119 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 119 112
rect 145 86 185 112
rect 211 86 217 112
rect -217 46 217 86
rect -217 20 -211 46
rect -185 20 -145 46
rect -119 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 119 46
rect 145 20 185 46
rect 211 20 217 46
rect -217 -20 217 20
rect -217 -46 -211 -20
rect -185 -46 -145 -20
rect -119 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 119 -20
rect 145 -46 185 -20
rect 211 -46 217 -20
rect -217 -86 217 -46
rect -217 -112 -211 -86
rect -185 -112 -145 -86
rect -119 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 119 -86
rect 145 -112 185 -86
rect 211 -112 217 -86
rect -217 -152 217 -112
rect -217 -178 -211 -152
rect -185 -178 -145 -152
rect -119 -178 -79 -152
rect -53 -178 -13 -152
rect 13 -178 53 -152
rect 79 -178 119 -152
rect 145 -178 185 -152
rect 211 -178 217 -152
rect -217 -218 217 -178
rect -217 -244 -211 -218
rect -185 -244 -145 -218
rect -119 -244 -79 -218
rect -53 -244 -13 -218
rect 13 -244 53 -218
rect 79 -244 119 -218
rect 145 -244 185 -218
rect 211 -244 217 -218
rect -217 -284 217 -244
rect -217 -310 -211 -284
rect -185 -310 -145 -284
rect -119 -310 -79 -284
rect -53 -310 -13 -284
rect 13 -310 53 -284
rect 79 -310 119 -284
rect 145 -310 185 -284
rect 211 -310 217 -284
rect -217 -350 217 -310
rect -217 -376 -211 -350
rect -185 -376 -145 -350
rect -119 -376 -79 -350
rect -53 -376 -13 -350
rect 13 -376 53 -350
rect 79 -376 119 -350
rect 145 -376 185 -350
rect 211 -376 217 -350
rect -217 -416 217 -376
rect -217 -442 -211 -416
rect -185 -442 -145 -416
rect -119 -442 -79 -416
rect -53 -442 -13 -416
rect 13 -442 53 -416
rect 79 -442 119 -416
rect 145 -442 185 -416
rect 211 -442 217 -416
rect -217 -482 217 -442
rect -217 -508 -211 -482
rect -185 -508 -145 -482
rect -119 -508 -79 -482
rect -53 -508 -13 -482
rect 13 -508 53 -482
rect 79 -508 119 -482
rect 145 -508 185 -482
rect 211 -508 217 -482
rect -217 -548 217 -508
rect -217 -574 -211 -548
rect -185 -574 -145 -548
rect -119 -574 -79 -548
rect -53 -574 -13 -548
rect 13 -574 53 -548
rect 79 -574 119 -548
rect 145 -574 185 -548
rect 211 -574 217 -548
rect -217 -614 217 -574
rect -217 -640 -211 -614
rect -185 -640 -145 -614
rect -119 -640 -79 -614
rect -53 -640 -13 -614
rect 13 -640 53 -614
rect 79 -640 119 -614
rect 145 -640 185 -614
rect 211 -640 217 -614
rect -217 -680 217 -640
rect -217 -706 -211 -680
rect -185 -706 -145 -680
rect -119 -706 -79 -680
rect -53 -706 -13 -680
rect 13 -706 53 -680
rect 79 -706 119 -680
rect 145 -706 185 -680
rect 211 -706 217 -680
rect -217 -746 217 -706
rect -217 -772 -211 -746
rect -185 -772 -145 -746
rect -119 -772 -79 -746
rect -53 -772 -13 -746
rect 13 -772 53 -746
rect 79 -772 119 -746
rect 145 -772 185 -746
rect 211 -772 217 -746
rect -217 -812 217 -772
rect -217 -838 -211 -812
rect -185 -838 -145 -812
rect -119 -838 -79 -812
rect -53 -838 -13 -812
rect 13 -838 53 -812
rect 79 -838 119 -812
rect 145 -838 185 -812
rect 211 -838 217 -812
rect -217 -878 217 -838
rect -217 -904 -211 -878
rect -185 -904 -145 -878
rect -119 -904 -79 -878
rect -53 -904 -13 -878
rect 13 -904 53 -878
rect 79 -904 119 -878
rect 145 -904 185 -878
rect 211 -904 217 -878
rect -217 -910 217 -904
<< via1 >>
rect -211 878 -185 904
rect -145 878 -119 904
rect -79 878 -53 904
rect -13 878 13 904
rect 53 878 79 904
rect 119 878 145 904
rect 185 878 211 904
rect -211 812 -185 838
rect -145 812 -119 838
rect -79 812 -53 838
rect -13 812 13 838
rect 53 812 79 838
rect 119 812 145 838
rect 185 812 211 838
rect -211 746 -185 772
rect -145 746 -119 772
rect -79 746 -53 772
rect -13 746 13 772
rect 53 746 79 772
rect 119 746 145 772
rect 185 746 211 772
rect -211 680 -185 706
rect -145 680 -119 706
rect -79 680 -53 706
rect -13 680 13 706
rect 53 680 79 706
rect 119 680 145 706
rect 185 680 211 706
rect -211 614 -185 640
rect -145 614 -119 640
rect -79 614 -53 640
rect -13 614 13 640
rect 53 614 79 640
rect 119 614 145 640
rect 185 614 211 640
rect -211 548 -185 574
rect -145 548 -119 574
rect -79 548 -53 574
rect -13 548 13 574
rect 53 548 79 574
rect 119 548 145 574
rect 185 548 211 574
rect -211 482 -185 508
rect -145 482 -119 508
rect -79 482 -53 508
rect -13 482 13 508
rect 53 482 79 508
rect 119 482 145 508
rect 185 482 211 508
rect -211 416 -185 442
rect -145 416 -119 442
rect -79 416 -53 442
rect -13 416 13 442
rect 53 416 79 442
rect 119 416 145 442
rect 185 416 211 442
rect -211 350 -185 376
rect -145 350 -119 376
rect -79 350 -53 376
rect -13 350 13 376
rect 53 350 79 376
rect 119 350 145 376
rect 185 350 211 376
rect -211 284 -185 310
rect -145 284 -119 310
rect -79 284 -53 310
rect -13 284 13 310
rect 53 284 79 310
rect 119 284 145 310
rect 185 284 211 310
rect -211 218 -185 244
rect -145 218 -119 244
rect -79 218 -53 244
rect -13 218 13 244
rect 53 218 79 244
rect 119 218 145 244
rect 185 218 211 244
rect -211 152 -185 178
rect -145 152 -119 178
rect -79 152 -53 178
rect -13 152 13 178
rect 53 152 79 178
rect 119 152 145 178
rect 185 152 211 178
rect -211 86 -185 112
rect -145 86 -119 112
rect -79 86 -53 112
rect -13 86 13 112
rect 53 86 79 112
rect 119 86 145 112
rect 185 86 211 112
rect -211 20 -185 46
rect -145 20 -119 46
rect -79 20 -53 46
rect -13 20 13 46
rect 53 20 79 46
rect 119 20 145 46
rect 185 20 211 46
rect -211 -46 -185 -20
rect -145 -46 -119 -20
rect -79 -46 -53 -20
rect -13 -46 13 -20
rect 53 -46 79 -20
rect 119 -46 145 -20
rect 185 -46 211 -20
rect -211 -112 -185 -86
rect -145 -112 -119 -86
rect -79 -112 -53 -86
rect -13 -112 13 -86
rect 53 -112 79 -86
rect 119 -112 145 -86
rect 185 -112 211 -86
rect -211 -178 -185 -152
rect -145 -178 -119 -152
rect -79 -178 -53 -152
rect -13 -178 13 -152
rect 53 -178 79 -152
rect 119 -178 145 -152
rect 185 -178 211 -152
rect -211 -244 -185 -218
rect -145 -244 -119 -218
rect -79 -244 -53 -218
rect -13 -244 13 -218
rect 53 -244 79 -218
rect 119 -244 145 -218
rect 185 -244 211 -218
rect -211 -310 -185 -284
rect -145 -310 -119 -284
rect -79 -310 -53 -284
rect -13 -310 13 -284
rect 53 -310 79 -284
rect 119 -310 145 -284
rect 185 -310 211 -284
rect -211 -376 -185 -350
rect -145 -376 -119 -350
rect -79 -376 -53 -350
rect -13 -376 13 -350
rect 53 -376 79 -350
rect 119 -376 145 -350
rect 185 -376 211 -350
rect -211 -442 -185 -416
rect -145 -442 -119 -416
rect -79 -442 -53 -416
rect -13 -442 13 -416
rect 53 -442 79 -416
rect 119 -442 145 -416
rect 185 -442 211 -416
rect -211 -508 -185 -482
rect -145 -508 -119 -482
rect -79 -508 -53 -482
rect -13 -508 13 -482
rect 53 -508 79 -482
rect 119 -508 145 -482
rect 185 -508 211 -482
rect -211 -574 -185 -548
rect -145 -574 -119 -548
rect -79 -574 -53 -548
rect -13 -574 13 -548
rect 53 -574 79 -548
rect 119 -574 145 -548
rect 185 -574 211 -548
rect -211 -640 -185 -614
rect -145 -640 -119 -614
rect -79 -640 -53 -614
rect -13 -640 13 -614
rect 53 -640 79 -614
rect 119 -640 145 -614
rect 185 -640 211 -614
rect -211 -706 -185 -680
rect -145 -706 -119 -680
rect -79 -706 -53 -680
rect -13 -706 13 -680
rect 53 -706 79 -680
rect 119 -706 145 -680
rect 185 -706 211 -680
rect -211 -772 -185 -746
rect -145 -772 -119 -746
rect -79 -772 -53 -746
rect -13 -772 13 -746
rect 53 -772 79 -746
rect 119 -772 145 -746
rect 185 -772 211 -746
rect -211 -838 -185 -812
rect -145 -838 -119 -812
rect -79 -838 -53 -812
rect -13 -838 13 -812
rect 53 -838 79 -812
rect 119 -838 145 -812
rect 185 -838 211 -812
rect -211 -904 -185 -878
rect -145 -904 -119 -878
rect -79 -904 -53 -878
rect -13 -904 13 -878
rect 53 -904 79 -878
rect 119 -904 145 -878
rect 185 -904 211 -878
<< metal2 >>
rect -217 904 217 910
rect -217 878 -211 904
rect -185 878 -145 904
rect -119 878 -79 904
rect -53 878 -13 904
rect 13 878 53 904
rect 79 878 119 904
rect 145 878 185 904
rect 211 878 217 904
rect -217 838 217 878
rect -217 812 -211 838
rect -185 812 -145 838
rect -119 812 -79 838
rect -53 812 -13 838
rect 13 812 53 838
rect 79 812 119 838
rect 145 812 185 838
rect 211 812 217 838
rect -217 772 217 812
rect -217 746 -211 772
rect -185 746 -145 772
rect -119 746 -79 772
rect -53 746 -13 772
rect 13 746 53 772
rect 79 746 119 772
rect 145 746 185 772
rect 211 746 217 772
rect -217 706 217 746
rect -217 680 -211 706
rect -185 680 -145 706
rect -119 680 -79 706
rect -53 680 -13 706
rect 13 680 53 706
rect 79 680 119 706
rect 145 680 185 706
rect 211 680 217 706
rect -217 640 217 680
rect -217 614 -211 640
rect -185 614 -145 640
rect -119 614 -79 640
rect -53 614 -13 640
rect 13 614 53 640
rect 79 614 119 640
rect 145 614 185 640
rect 211 614 217 640
rect -217 574 217 614
rect -217 548 -211 574
rect -185 548 -145 574
rect -119 548 -79 574
rect -53 548 -13 574
rect 13 548 53 574
rect 79 548 119 574
rect 145 548 185 574
rect 211 548 217 574
rect -217 508 217 548
rect -217 482 -211 508
rect -185 482 -145 508
rect -119 482 -79 508
rect -53 482 -13 508
rect 13 482 53 508
rect 79 482 119 508
rect 145 482 185 508
rect 211 482 217 508
rect -217 442 217 482
rect -217 416 -211 442
rect -185 416 -145 442
rect -119 416 -79 442
rect -53 416 -13 442
rect 13 416 53 442
rect 79 416 119 442
rect 145 416 185 442
rect 211 416 217 442
rect -217 376 217 416
rect -217 350 -211 376
rect -185 350 -145 376
rect -119 350 -79 376
rect -53 350 -13 376
rect 13 350 53 376
rect 79 350 119 376
rect 145 350 185 376
rect 211 350 217 376
rect -217 310 217 350
rect -217 284 -211 310
rect -185 284 -145 310
rect -119 284 -79 310
rect -53 284 -13 310
rect 13 284 53 310
rect 79 284 119 310
rect 145 284 185 310
rect 211 284 217 310
rect -217 244 217 284
rect -217 218 -211 244
rect -185 218 -145 244
rect -119 218 -79 244
rect -53 218 -13 244
rect 13 218 53 244
rect 79 218 119 244
rect 145 218 185 244
rect 211 218 217 244
rect -217 178 217 218
rect -217 152 -211 178
rect -185 152 -145 178
rect -119 152 -79 178
rect -53 152 -13 178
rect 13 152 53 178
rect 79 152 119 178
rect 145 152 185 178
rect 211 152 217 178
rect -217 112 217 152
rect -217 86 -211 112
rect -185 86 -145 112
rect -119 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 119 112
rect 145 86 185 112
rect 211 86 217 112
rect -217 46 217 86
rect -217 20 -211 46
rect -185 20 -145 46
rect -119 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 119 46
rect 145 20 185 46
rect 211 20 217 46
rect -217 -20 217 20
rect -217 -46 -211 -20
rect -185 -46 -145 -20
rect -119 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 119 -20
rect 145 -46 185 -20
rect 211 -46 217 -20
rect -217 -86 217 -46
rect -217 -112 -211 -86
rect -185 -112 -145 -86
rect -119 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 119 -86
rect 145 -112 185 -86
rect 211 -112 217 -86
rect -217 -152 217 -112
rect -217 -178 -211 -152
rect -185 -178 -145 -152
rect -119 -178 -79 -152
rect -53 -178 -13 -152
rect 13 -178 53 -152
rect 79 -178 119 -152
rect 145 -178 185 -152
rect 211 -178 217 -152
rect -217 -218 217 -178
rect -217 -244 -211 -218
rect -185 -244 -145 -218
rect -119 -244 -79 -218
rect -53 -244 -13 -218
rect 13 -244 53 -218
rect 79 -244 119 -218
rect 145 -244 185 -218
rect 211 -244 217 -218
rect -217 -284 217 -244
rect -217 -310 -211 -284
rect -185 -310 -145 -284
rect -119 -310 -79 -284
rect -53 -310 -13 -284
rect 13 -310 53 -284
rect 79 -310 119 -284
rect 145 -310 185 -284
rect 211 -310 217 -284
rect -217 -350 217 -310
rect -217 -376 -211 -350
rect -185 -376 -145 -350
rect -119 -376 -79 -350
rect -53 -376 -13 -350
rect 13 -376 53 -350
rect 79 -376 119 -350
rect 145 -376 185 -350
rect 211 -376 217 -350
rect -217 -416 217 -376
rect -217 -442 -211 -416
rect -185 -442 -145 -416
rect -119 -442 -79 -416
rect -53 -442 -13 -416
rect 13 -442 53 -416
rect 79 -442 119 -416
rect 145 -442 185 -416
rect 211 -442 217 -416
rect -217 -482 217 -442
rect -217 -508 -211 -482
rect -185 -508 -145 -482
rect -119 -508 -79 -482
rect -53 -508 -13 -482
rect 13 -508 53 -482
rect 79 -508 119 -482
rect 145 -508 185 -482
rect 211 -508 217 -482
rect -217 -548 217 -508
rect -217 -574 -211 -548
rect -185 -574 -145 -548
rect -119 -574 -79 -548
rect -53 -574 -13 -548
rect 13 -574 53 -548
rect 79 -574 119 -548
rect 145 -574 185 -548
rect 211 -574 217 -548
rect -217 -614 217 -574
rect -217 -640 -211 -614
rect -185 -640 -145 -614
rect -119 -640 -79 -614
rect -53 -640 -13 -614
rect 13 -640 53 -614
rect 79 -640 119 -614
rect 145 -640 185 -614
rect 211 -640 217 -614
rect -217 -680 217 -640
rect -217 -706 -211 -680
rect -185 -706 -145 -680
rect -119 -706 -79 -680
rect -53 -706 -13 -680
rect 13 -706 53 -680
rect 79 -706 119 -680
rect 145 -706 185 -680
rect 211 -706 217 -680
rect -217 -746 217 -706
rect -217 -772 -211 -746
rect -185 -772 -145 -746
rect -119 -772 -79 -746
rect -53 -772 -13 -746
rect 13 -772 53 -746
rect 79 -772 119 -746
rect 145 -772 185 -746
rect 211 -772 217 -746
rect -217 -812 217 -772
rect -217 -838 -211 -812
rect -185 -838 -145 -812
rect -119 -838 -79 -812
rect -53 -838 -13 -812
rect 13 -838 53 -812
rect 79 -838 119 -812
rect 145 -838 185 -812
rect 211 -838 217 -812
rect -217 -878 217 -838
rect -217 -904 -211 -878
rect -185 -904 -145 -878
rect -119 -904 -79 -878
rect -53 -904 -13 -878
rect 13 -904 53 -878
rect 79 -904 119 -878
rect 145 -904 185 -878
rect 211 -904 217 -878
rect -217 -910 217 -904
<< end >>
