magic
tech gf180mcuC
magscale 1 10
timestamp 1695127730
<< nwell >>
rect 3729 -609 3828 -532
<< ndiff >>
rect 994 -400 1050 -344
rect 3242 -409 3298 -353
rect 4773 -407 4825 -355
<< psubdiff >>
rect 75 -21 464 26
rect 1201 -21 1590 26
rect 2327 -21 2716 26
rect 3453 -21 3842 26
rect 4484 -241 4527 -162
<< nsubdiff >>
rect 4482 -1020 4538 -948
<< polysilicon >>
rect 1488 554 1540 606
rect 2616 545 2672 601
rect 3729 546 3809 608
rect 3575 438 3577 512
rect 569 -607 572 -548
rect 1482 -606 1506 -538
rect 1556 -606 1559 -538
rect 2603 -548 2605 -538
rect 2616 -595 2668 -542
rect 2842 -607 2843 -538
rect 3740 -602 3796 -545
<< metal1 >>
rect 1243 917 1572 1011
rect 4474 913 4536 1050
rect 247 725 314 827
rect 1375 813 1437 825
rect 813 641 870 800
rect 1375 660 1439 813
rect 1375 659 1437 660
rect 1541 657 1598 816
rect 1699 655 1761 821
rect 1945 635 2002 794
rect 2099 638 2161 804
rect 2342 657 2404 823
rect 2506 661 2568 827
rect 2662 657 2724 823
rect 2825 661 2887 827
rect 3229 633 3291 799
rect 3630 660 3692 826
rect 3788 657 3850 823
rect 3953 656 4015 822
rect 4190 639 4252 805
rect 4357 636 4419 802
rect 351 606 431 609
rect 1478 606 1557 607
rect 351 552 363 606
rect 415 552 431 606
rect 351 549 431 552
rect 496 603 589 606
rect 496 551 509 603
rect 561 551 589 603
rect 351 548 442 549
rect 496 548 589 551
rect 1478 554 1489 606
rect 1541 554 1557 606
rect 1478 549 1557 554
rect 1623 605 1717 607
rect 1623 551 1635 605
rect 1687 551 1717 605
rect 1623 548 1717 551
rect 2604 593 2684 608
rect -380 525 -196 540
rect 2604 537 2616 593
rect 2672 537 2684 593
rect 2749 553 2762 606
rect 2814 553 2844 606
rect 2749 548 2844 553
rect 3729 601 3812 608
rect 3729 546 3741 601
rect 3797 546 3812 601
rect 3874 604 3971 607
rect 3874 551 3893 604
rect 3946 551 3971 604
rect 3874 548 3971 551
rect 3729 538 3812 546
rect 2604 530 2683 537
rect -380 471 -267 525
rect -213 471 -196 525
rect 2371 522 2459 523
rect -96 471 207 521
rect -380 459 -196 471
rect -279 456 -196 459
rect 63 457 207 471
rect 63 403 101 457
rect 154 403 207 457
rect 865 453 919 518
rect 1201 485 1312 511
rect 1201 429 1229 485
rect 1287 429 1312 485
rect 1992 455 2057 519
rect 2370 507 2459 522
rect 2370 455 2395 507
rect 2447 455 2459 507
rect 2370 443 2459 455
rect 3496 505 3581 517
rect 3496 449 3509 505
rect 3569 449 3581 505
rect 4474 449 4537 913
rect 2370 442 2458 443
rect 3496 442 3581 449
rect 63 388 207 403
rect 973 411 1062 428
rect 1201 412 1312 429
rect 2209 415 2293 429
rect 2209 413 2222 415
rect 973 354 986 411
rect 1042 354 1062 411
rect 973 340 1062 354
rect 2104 359 2222 413
rect 2278 359 2293 415
rect 2104 352 2293 359
rect 2209 345 2293 352
rect 3227 415 3313 423
rect 3227 351 3239 415
rect 3300 351 3313 415
rect 3227 346 3313 351
rect 4319 386 4419 406
rect 4319 329 4335 386
rect 4393 329 4419 386
rect 4319 315 4419 329
rect 4475 354 4537 449
rect 4475 338 4637 354
rect 4475 312 4638 338
rect 4476 306 4638 312
rect -86 142 1 143
rect -86 109 2 142
rect 1053 109 1128 146
rect 2192 110 2254 141
rect 2192 109 2348 110
rect 3334 109 3380 152
rect -86 94 63 109
rect -86 61 64 94
rect 1053 61 1182 109
rect 1681 107 1850 109
rect 2192 68 2292 109
rect 1298 26 1473 68
rect 2192 64 2291 68
rect 3334 62 3423 109
rect 4581 26 4638 306
rect 4866 26 5092 27
rect 75 -21 464 26
rect 553 -7 773 8
rect 1201 -21 1590 26
rect 1679 -7 1899 8
rect 2327 -21 2716 26
rect 2805 -8 3025 7
rect 3453 -21 3842 26
rect 4564 23 5092 26
rect 3931 -6 4151 9
rect -84 -109 72 -51
rect 1055 -109 1192 -52
rect 1298 -60 1473 -21
rect 4564 -56 5095 23
rect 2187 -109 2318 -64
rect 3321 -72 3423 -56
rect 4581 -57 4638 -56
rect 3321 -109 3422 -72
rect -84 -154 2 -109
rect 1055 -141 1128 -109
rect 2187 -110 2348 -109
rect 2187 -143 2254 -110
rect 3321 -143 3380 -109
rect 3321 -144 3340 -143
rect 4484 -241 4527 -162
rect 979 -344 1065 -328
rect -151 -349 -75 -344
rect -151 -401 -139 -349
rect -87 -401 -75 -349
rect -151 -407 -75 -401
rect 979 -400 994 -344
rect 1050 -400 1065 -344
rect 2102 -343 2192 -327
rect 979 -415 1065 -400
rect 1180 -404 1302 -389
rect 2102 -404 2110 -343
rect 2169 -404 2192 -343
rect 1180 -434 1305 -404
rect 2102 -414 2192 -404
rect 3230 -352 3312 -332
rect 3230 -409 3242 -352
rect 3298 -409 3312 -352
rect 3230 -414 3312 -409
rect 4357 -336 4456 -322
rect 4357 -340 4367 -336
rect 4357 -398 4366 -340
rect 4428 -397 4456 -336
rect 4426 -398 4456 -397
rect 4357 -414 4456 -398
rect 4760 -355 4834 -343
rect 5002 -353 5095 -56
rect 4760 -407 4773 -355
rect 4825 -407 4834 -355
rect 4760 -417 4834 -407
rect -259 -461 -194 -454
rect -380 -473 -194 -461
rect 111 -463 204 -437
rect -380 -535 -253 -473
rect -201 -535 -194 -473
rect -136 -510 204 -463
rect 1180 -486 1213 -434
rect 1183 -492 1213 -486
rect 1277 -492 1305 -434
rect 4905 -429 5095 -353
rect 1183 -498 1305 -492
rect 2377 -453 2457 -442
rect 2377 -510 2389 -453
rect 2445 -510 2457 -453
rect 2377 -521 2457 -510
rect 3500 -454 3582 -442
rect 3500 -508 3518 -454
rect 3571 -508 3582 -454
rect 4618 -457 4714 -453
rect 3500 -522 3582 -508
rect 4567 -474 4714 -457
rect 4567 -528 4640 -474
rect 4694 -528 4714 -474
rect -380 -542 -194 -535
rect 1636 -536 1713 -535
rect -259 -543 -194 -542
rect 1482 -547 1559 -538
rect 359 -550 433 -548
rect 496 -550 572 -548
rect 359 -551 450 -550
rect 359 -605 367 -551
rect 419 -605 450 -551
rect 359 -608 450 -605
rect 496 -602 508 -550
rect 560 -602 572 -550
rect 496 -607 572 -602
rect 1482 -600 1495 -547
rect 1547 -600 1559 -547
rect 1482 -606 1559 -600
rect 1636 -546 1724 -536
rect 1636 -598 1648 -546
rect 1704 -598 1724 -546
rect 2603 -542 2683 -538
rect 2603 -548 2616 -542
rect 1636 -602 1724 -598
rect 2605 -595 2616 -548
rect 2668 -595 2683 -542
rect 2605 -605 2683 -595
rect 2756 -543 2843 -538
rect 2756 -602 2776 -543
rect 2831 -602 2843 -543
rect 2756 -607 2843 -602
rect 3729 -545 3828 -532
rect 3729 -602 3742 -545
rect 3798 -602 3828 -545
rect 3729 -609 3828 -602
rect 3881 -544 3968 -538
rect 3881 -605 3896 -544
rect 3952 -605 3968 -544
rect 4567 -542 4714 -528
rect 4567 -545 4703 -542
rect 3881 -607 3968 -605
rect 4482 -1020 4538 -948
rect 4905 -1045 5002 -429
<< via1 >>
rect 363 552 415 606
rect 509 551 561 603
rect 1489 554 1541 606
rect 1635 551 1687 605
rect 2616 537 2672 593
rect 2762 553 2814 606
rect 3741 546 3797 601
rect 3893 551 3946 604
rect -267 471 -213 525
rect 101 403 154 457
rect 1229 429 1287 485
rect 2395 455 2447 507
rect 3509 449 3569 505
rect 986 354 1042 411
rect 2222 359 2278 415
rect 3239 351 3300 415
rect 4335 329 4393 386
rect -139 -401 -87 -349
rect 994 -400 1050 -344
rect 2110 -404 2169 -343
rect 3242 -409 3298 -352
rect 4367 -340 4428 -336
rect 4366 -397 4428 -340
rect 4366 -398 4426 -397
rect 4773 -407 4825 -355
rect -253 -535 -201 -473
rect 1213 -492 1277 -434
rect 2389 -510 2445 -453
rect 3518 -508 3571 -454
rect 4640 -528 4694 -474
rect 367 -605 419 -551
rect 508 -602 560 -550
rect 1495 -600 1547 -547
rect 1648 -598 1704 -546
rect 2616 -595 2668 -542
rect 2776 -602 2831 -543
rect 3742 -602 3798 -545
rect 3896 -605 3952 -544
<< metal2 >>
rect 2598 898 2675 907
rect -276 894 2675 898
rect -276 838 2608 894
rect 2665 838 2675 894
rect -276 835 2675 838
rect -276 541 -205 835
rect 2598 828 2675 835
rect 496 697 4539 763
rect 496 674 589 697
rect -288 525 -205 541
rect -288 471 -267 525
rect -213 471 -205 525
rect -288 457 -205 471
rect -147 606 428 613
rect -147 603 363 606
rect 415 603 428 606
rect -147 547 361 603
rect 417 547 428 603
rect 493 603 589 674
rect 493 551 509 603
rect 561 551 589 603
rect 645 626 1144 627
rect 645 568 665 626
rect 721 620 1144 626
rect 721 568 1080 620
rect 645 567 1080 568
rect 1067 564 1080 567
rect 1136 566 1144 620
rect 1476 606 1557 615
rect 1136 564 1141 566
rect 1067 554 1141 564
rect 1476 554 1489 606
rect 1541 554 1557 606
rect 493 550 589 551
rect 496 548 589 550
rect 1476 549 1557 554
rect 1618 605 1714 697
rect 1618 551 1635 605
rect 1687 551 1714 605
rect -147 535 428 547
rect -147 -344 -91 535
rect 1201 485 1312 511
rect 63 473 203 477
rect 1201 473 1229 485
rect 63 457 783 473
rect 63 403 101 457
rect 154 407 783 457
rect 1199 429 1229 473
rect 1287 473 1312 485
rect 1287 429 1315 473
rect 973 412 1062 428
rect 154 403 203 407
rect 63 388 203 403
rect 725 210 782 407
rect 973 354 985 412
rect 1042 354 1062 412
rect 1199 407 1315 429
rect 973 340 1062 354
rect 1241 210 1308 407
rect 725 145 1308 210
rect 726 144 1308 145
rect 1241 -165 1308 144
rect 783 -225 1308 -165
rect -151 -349 -75 -344
rect -151 -401 -139 -349
rect -87 -401 -75 -349
rect 783 -388 847 -225
rect -151 -407 -75 -401
rect 359 -448 847 -388
rect 979 -344 1065 -328
rect 979 -400 994 -344
rect 1050 -400 1065 -344
rect 1241 -388 1308 -225
rect 979 -415 1065 -400
rect 1180 -434 1308 -388
rect 359 -449 811 -448
rect 1180 -449 1213 -434
rect -259 -473 -194 -454
rect -259 -535 -253 -473
rect -201 -535 -194 -473
rect -259 -543 -194 -535
rect -255 -629 -196 -543
rect 359 -549 433 -449
rect 1183 -492 1213 -449
rect 1277 -492 1308 -434
rect 1183 -516 1308 -492
rect 1183 -520 1262 -516
rect 1486 -530 1545 549
rect 1618 548 1714 551
rect 1817 616 2449 626
rect 1817 560 1832 616
rect 1888 566 2449 616
rect 1888 560 1901 566
rect 1817 549 1901 560
rect 2371 522 2449 566
rect 2604 608 2683 615
rect 2604 601 2684 608
rect 2604 537 2616 601
rect 2672 537 2684 601
rect 2745 606 2841 697
rect 2745 553 2762 606
rect 2814 553 2841 606
rect 2745 547 2841 553
rect 3729 601 3812 608
rect 3729 546 3741 601
rect 3797 546 3812 601
rect 3871 604 3968 697
rect 3871 551 3893 604
rect 3946 551 3968 604
rect 3871 548 3968 551
rect 3729 538 3812 546
rect 2371 507 2458 522
rect 2371 455 2395 507
rect 2447 455 2458 507
rect 2371 442 2458 455
rect 2606 443 2683 537
rect 3496 505 3581 517
rect 3496 449 3509 505
rect 3569 449 3581 505
rect 2999 443 3058 444
rect 2209 415 2293 429
rect 2209 359 2222 415
rect 2278 359 2293 415
rect 2209 345 2293 359
rect 2102 -343 2192 -327
rect 2102 -404 2110 -343
rect 2169 -404 2192 -343
rect 2102 -414 2192 -404
rect 2378 -415 2447 442
rect 2606 385 3061 443
rect 3496 442 3581 449
rect 3227 415 3313 423
rect 2999 207 3058 385
rect 3227 351 3239 415
rect 3300 351 3313 415
rect 3227 346 3313 351
rect 3505 385 3577 442
rect 3505 207 3571 385
rect 2999 145 3571 207
rect 2999 141 3058 145
rect 3505 -218 3571 145
rect 2997 -274 3571 -218
rect 2997 -415 3056 -274
rect 3230 -352 3312 -332
rect 3230 -409 3242 -352
rect 3298 -409 3312 -352
rect 3230 -414 3312 -409
rect 2377 -453 2458 -415
rect 2377 -510 2389 -453
rect 2445 -510 2458 -453
rect 2377 -512 2458 -510
rect 2612 -471 3056 -415
rect 3505 -442 3571 -274
rect 3500 -454 3582 -442
rect 2612 -472 3055 -471
rect 2377 -521 2457 -512
rect 2378 -523 2447 -521
rect 1477 -532 1545 -530
rect 1477 -538 1554 -532
rect 1636 -536 1713 -535
rect 1477 -546 1559 -538
rect 353 -550 433 -549
rect 496 -550 572 -548
rect 353 -551 439 -550
rect 353 -605 367 -551
rect 419 -605 439 -551
rect 353 -608 439 -605
rect 496 -602 508 -550
rect 560 -602 572 -550
rect 496 -607 572 -602
rect 1477 -603 1488 -546
rect 1544 -547 1559 -546
rect 1547 -600 1559 -547
rect 1544 -603 1559 -600
rect 1636 -546 1724 -536
rect 2612 -538 2671 -472
rect 3500 -508 3518 -454
rect 3571 -508 3582 -454
rect 3500 -522 3582 -508
rect 3734 -532 3794 538
rect 4330 406 4416 419
rect 4319 386 4419 406
rect 4319 329 4335 386
rect 4393 329 4419 386
rect 4319 315 4419 329
rect 4477 -60 4538 697
rect 4477 -61 4815 -60
rect 4477 -65 4816 -61
rect 4477 -123 4817 -65
rect 4477 -125 4538 -123
rect 4357 -336 4456 -322
rect 4357 -340 4367 -336
rect 4357 -398 4366 -340
rect 4428 -397 4456 -336
rect 4761 -343 4817 -123
rect 4426 -398 4456 -397
rect 4357 -414 4456 -398
rect 4760 -355 4834 -343
rect 4760 -407 4773 -355
rect 4825 -407 4834 -355
rect 4760 -417 4834 -407
rect 4618 -474 4714 -453
rect 4618 -528 4640 -474
rect 4694 -528 4714 -474
rect 1636 -598 1648 -546
rect 1704 -598 1724 -546
rect 1636 -602 1724 -598
rect 2605 -542 2683 -538
rect 2605 -595 2616 -542
rect 2668 -595 2683 -542
rect 1477 -606 1559 -603
rect -255 -830 -197 -629
rect 505 -685 562 -607
rect 1477 -608 1554 -606
rect 1647 -685 1709 -602
rect 2605 -605 2683 -595
rect 2756 -543 2843 -538
rect 2756 -602 2776 -543
rect 2831 -602 2843 -543
rect 2612 -606 2671 -605
rect 2756 -607 2843 -602
rect 3729 -545 3825 -532
rect 3729 -602 3740 -545
rect 3798 -602 3825 -545
rect 2768 -685 2825 -607
rect 3729 -609 3825 -602
rect 3881 -544 3968 -538
rect 4618 -542 4714 -528
rect 3881 -605 3896 -544
rect 3952 -605 3968 -544
rect 3881 -607 3968 -605
rect 3729 -614 3808 -609
rect 3891 -685 3947 -607
rect 4651 -685 4711 -542
rect 502 -748 4711 -685
rect 4651 -750 4711 -748
rect 1481 -830 1556 -823
rect 3725 -829 3806 -819
rect 3725 -830 3737 -829
rect -255 -833 3737 -830
rect -255 -890 1491 -833
rect 1547 -885 3737 -833
rect 3794 -885 3806 -829
rect 1547 -890 3806 -885
rect -255 -893 3806 -890
rect 1481 -899 1556 -893
rect 3725 -896 3806 -893
<< via2 >>
rect 2608 838 2665 894
rect 361 552 363 603
rect 363 552 415 603
rect 415 552 417 603
rect 361 547 417 552
rect 665 568 721 626
rect 1080 564 1136 620
rect 985 411 1042 412
rect 985 354 986 411
rect 986 354 1042 411
rect 994 -400 1050 -344
rect 1832 560 1888 616
rect 2616 593 2672 601
rect 2616 545 2672 593
rect 2222 359 2278 415
rect 2110 -404 2169 -343
rect 3239 351 3300 415
rect 3242 -409 3298 -353
rect 1488 -547 1544 -546
rect 1488 -600 1495 -547
rect 1495 -600 1544 -547
rect 1488 -603 1544 -600
rect 4336 330 4393 386
rect 4366 -398 4426 -340
rect 3740 -602 3742 -545
rect 3742 -602 3796 -545
rect 1491 -890 1547 -833
rect 3737 -885 3794 -829
<< metal3 >>
rect 796 797 862 1015
rect 796 679 863 797
rect 362 626 741 627
rect 362 612 665 626
rect 350 603 665 612
rect 350 547 361 603
rect 417 568 665 603
rect 721 568 741 626
rect 417 567 741 568
rect 417 547 429 567
rect 350 536 429 547
rect 797 240 863 679
rect 919 428 990 1007
rect 1141 626 1878 627
rect 1067 620 1901 626
rect 1067 564 1080 620
rect 1136 616 1901 620
rect 1136 566 1832 616
rect 1136 564 1141 566
rect 1067 554 1141 564
rect 1817 560 1832 566
rect 1888 560 1901 616
rect 1817 549 1901 560
rect 919 412 1062 428
rect 919 354 985 412
rect 1042 354 1062 412
rect 919 342 1062 354
rect 973 340 1062 342
rect 796 -22 863 240
rect 1999 290 2087 986
rect 2224 429 2311 982
rect 3019 977 3079 993
rect 2598 894 2675 907
rect 2598 838 2608 894
rect 2665 838 2675 894
rect 2598 828 2675 838
rect 2605 615 2672 828
rect 2604 601 2683 615
rect 2604 545 2616 601
rect 2672 545 2683 601
rect 2604 537 2683 545
rect 2209 415 2293 429
rect 2209 359 2222 415
rect 2278 359 2293 415
rect 2209 345 2293 359
rect 1999 288 2189 290
rect 1999 211 2190 288
rect 796 -289 862 -22
rect 796 -344 1065 -289
rect 2104 -327 2190 211
rect 796 -347 994 -344
rect 979 -400 994 -347
rect 1050 -400 1065 -344
rect 979 -415 1065 -400
rect 2102 -343 2192 -327
rect 2102 -404 2110 -343
rect 2169 -404 2192 -343
rect 3016 -342 3102 977
rect 3236 423 3294 990
rect 3227 415 3313 423
rect 3227 351 3239 415
rect 3300 351 3313 415
rect 3227 346 3313 351
rect 3230 -342 3312 -332
rect 3016 -353 3312 -342
rect 3016 -397 3242 -353
rect 3018 -398 3242 -397
rect 2102 -414 2192 -404
rect 3230 -409 3242 -398
rect 3298 -409 3312 -353
rect 4074 -338 4160 970
rect 4336 406 4396 958
rect 4319 386 4419 406
rect 4319 330 4336 386
rect 4393 330 4419 386
rect 4319 315 4419 330
rect 4357 -338 4456 -322
rect 4074 -340 4456 -338
rect 4074 -398 4366 -340
rect 4426 -398 4456 -340
rect 4074 -404 4456 -398
rect 4086 -405 4456 -404
rect 3230 -414 3312 -409
rect 4357 -414 4456 -405
rect 1477 -532 1544 -530
rect 1477 -546 1554 -532
rect 1477 -603 1488 -546
rect 1544 -603 1554 -546
rect 1477 -608 1554 -603
rect 3729 -545 3828 -532
rect 3729 -602 3740 -545
rect 3796 -602 3828 -545
rect 1487 -823 1544 -608
rect 3729 -609 3828 -602
rect 3729 -614 3808 -609
rect 3734 -819 3797 -614
rect 1481 -833 1556 -823
rect 1481 -890 1491 -833
rect 1547 -890 1556 -833
rect 1481 -899 1556 -890
rect 3725 -829 3806 -819
rect 3725 -885 3737 -829
rect 3794 -885 3806 -829
rect 3725 -896 3806 -885
use and_3_ibr  and_3_ibr_0
timestamp 1695127730
transform 1 0 -8 0 1 0
box 8 0 1136 1051
use and_3_ibr  and_3_ibr_1
timestamp 1695127730
transform 1 0 1118 0 1 0
box 8 0 1136 1051
use and_3_ibr  and_3_ibr_2
timestamp 1695127730
transform 1 0 2244 0 1 0
box 8 0 1136 1051
use and_3_ibr  and_3_ibr_3
timestamp 1695127730
transform 1 0 3370 0 1 0
box 8 0 1136 1051
use and_3_ibr  and_3_ibr_4
timestamp 1695127730
transform 1 0 -8 0 -1 0
box 8 0 1136 1051
use and_3_ibr  and_3_ibr_5
timestamp 1695127730
transform 1 0 1118 0 -1 0
box 8 0 1136 1051
use and_3_ibr  and_3_ibr_6
timestamp 1695127730
transform 1 0 2244 0 -1 0
box 8 0 1136 1051
use and_3_ibr  and_3_ibr_7
timestamp 1695127730
transform 1 0 3370 0 -1 0
box 8 0 1136 1051
use nverterlayout_ibr  nverterlayout_ibr_0
timestamp 1695109904
transform 1 0 4593 0 -1 79
box -88 220 316 1130
use nverterlayout_ibr  nverterlayout_ibr_1
timestamp 1695109904
transform 1 0 -314 0 -1 79
box -88 220 316 1130
use nverterlayout_ibr  nverterlayout_ibr_2
timestamp 1695109904
transform 1 0 -314 0 1 -78
box -88 220 316 1130
<< labels >>
flabel via1 -248 499 -248 499 0 FreeSans 480 0 0 0 IN1
port 0 nsew
flabel via1 -244 -501 -244 -501 0 FreeSans 480 0 0 0 IN2
port 1 nsew
flabel via1 4648 -509 4648 -509 0 FreeSans 480 0 0 0 IN3
port 2 nsew
flabel metal3 953 979 953 979 0 FreeSans 480 0 0 0 D0
port 3 nsew
flabel metal3 820 981 820 981 0 FreeSans 480 0 0 0 D1
port 4 nsew
flabel metal3 2252 947 2252 947 0 FreeSans 480 0 0 0 D2
port 5 nsew
flabel metal3 2052 949 2052 949 0 FreeSans 480 0 0 0 D3
port 6 nsew
flabel metal3 3259 941 3259 941 0 FreeSans 480 0 0 0 D4
port 7 nsew
flabel metal3 3044 955 3044 955 0 FreeSans 480 0 0 0 D5
port 8 nsew
flabel metal3 4366 933 4366 933 0 FreeSans 480 0 0 0 D6
port 9 nsew
flabel metal3 4116 935 4116 935 0 FreeSans 480 0 0 0 D7
port 10 nsew
flabel metal1 1383 960 1383 960 0 FreeSans 480 0 0 0 VDD
port 11 nsew
flabel metal1 1381 2 1381 2 0 FreeSans 480 0 0 0 VSS
port 12 nsew
<< end >>
