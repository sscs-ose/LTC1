* NGSPICE file created from INVERTER_magic.ext - technology: gf180mcuC

.subckt pmos_3p3_MGRCNG a_n204_n36# a_56_n69# a_112_n25# a_n112_n69# w_n290_n161#
+ a_n56_n25#
X0 a_n56_n25# a_n112_n69# a_n204_n36# w_n290_n161# pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X1 a_112_n25# a_56_n69# a_n56_n25# w_n290_n161# pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
.ends

.subckt nmos_3p3_H9QVWA a_n120_n36# a_28_n25# a_n28_n69# VSUBS
X0 a_28_n25# a_n28_n69# a_n120_n36# VSUBS nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
.ends

.subckt INVERTER_magic IN OUT VDD VSS
Xpmos_3p3_MGRCNG_0 OUT IN OUT IN VDD VDD pmos_3p3_MGRCNG
Xnmos_3p3_H9QVWA_0 VSS OUT IN VSS nmos_3p3_H9QVWA
Xnmos_3p3_H9QVWA_1 VSS VSS VSS VSS nmos_3p3_H9QVWA
.ends

