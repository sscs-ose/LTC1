* NGSPICE file created from 200_ohm_magic_flat.ext - technology: gf180mcuC

.subckt x200_ohm_magic_flat R1_IN R2_IN COMMON VDD
X0 VDD.t3 VDD.t4 VDD.t2 ppolyf_u r_width=1u r_length=3.9u
X1 VDD.t6 VDD.t7 VDD.t5 ppolyf_u r_width=1u r_length=3.9u
X2 VDD.t9 VDD.t10 VDD.t2 ppolyf_u r_width=1u r_length=3.9u
X3 COMMON.t4 R1_IN.t1 VDD.t1 ppolyf_u r_width=1u r_length=3.9u
X4 R1_IN.t3 COMMON.t6 VDD.t12 ppolyf_u r_width=1u r_length=3.9u
X5 R2_IN.t1 COMMON.t1 VDD.t1 ppolyf_u r_width=1u r_length=3.9u
X6 COMMON.t14 R2_IN.t6 VDD.t13 ppolyf_u r_width=1u r_length=3.9u
X7 VDD.t16 VDD.t17 VDD.t5 ppolyf_u r_width=1u r_length=3.9u
X8 COMMON.t3 R2_IN.t2 VDD.t8 ppolyf_u r_width=1u r_length=3.9u
X9 COMMON.t13 R1_IN.t7 VDD.t14 ppolyf_u r_width=1u r_length=3.9u
X10 R2_IN.t5 COMMON.t11 VDD.t15 ppolyf_u r_width=1u r_length=3.9u
X11 R2_IN.t4 COMMON.t10 VDD.t14 ppolyf_u r_width=1u r_length=3.9u
X12 COMMON.t15 R2_IN.t7 VDD.t11 ppolyf_u r_width=1u r_length=3.9u
X13 COMMON.t9 R2_IN.t3 VDD.t12 ppolyf_u r_width=1u r_length=3.9u
X14 COMMON.t12 R1_IN.t6 VDD.t15 ppolyf_u r_width=1u r_length=3.9u
X15 R2_IN.t0 COMMON.t0 VDD.t0 ppolyf_u r_width=1u r_length=3.9u
X16 COMMON.t2 R1_IN.t0 VDD.t0 ppolyf_u r_width=1u r_length=3.9u
X17 R1_IN.t4 COMMON.t7 VDD.t8 ppolyf_u r_width=1u r_length=3.9u
X18 R1_IN.t5 COMMON.t8 VDD.t13 ppolyf_u r_width=1u r_length=3.9u
X19 R1_IN.t2 COMMON.t5 VDD.t11 ppolyf_u r_width=1u r_length=3.9u
R0 VDD.n343 VDD.t14 13.6736
R1 VDD.n335 VDD.t8 12.4306
R2 VDD.n177 VDD.t12 9.32306
R3 VDD.n138 VDD.t2 8.08005
R4 VDD.n326 VDD.t1 8.08005
R5 VDD.n100 VDD.t9 6.90863
R6 VDD.n59 VDD.t3 6.90726
R7 VDD.n69 VDD.t10 6.90243
R8 VDD.n39 VDD.t4 6.89072
R9 VDD.n274 VDD.t16 6.85823
R10 VDD.n250 VDD.t17 6.85823
R11 VDD.n243 VDD.t6 6.85823
R12 VDD.n224 VDD.t7 6.85823
R13 VDD.n165 VDD.t0 4.97253
R14 VDD.n147 VDD.t15 3.72952
R15 VDD.n317 VDD.t13 3.72952
R16 VDD.n217 VDD.n184 3.1505
R17 VDD.n282 VDD.n281 3.1505
R18 VDD.n279 VDD.n278 3.1505
R19 VDD.n277 VDD.n276 3.1505
R20 VDD.n273 VDD.n272 3.1505
R21 VDD.n271 VDD.n270 3.1505
R22 VDD.n268 VDD.n267 3.1505
R23 VDD.n266 VDD.n265 3.1505
R24 VDD.n263 VDD.n262 3.1505
R25 VDD.n261 VDD.n260 3.1505
R26 VDD.n258 VDD.n257 3.1505
R27 VDD.n256 VDD.n255 3.1505
R28 VDD.n254 VDD.n253 3.1505
R29 VDD.n252 VDD.n251 3.1505
R30 VDD.n249 VDD.n248 3.1505
R31 VDD.n247 VDD.n246 3.1505
R32 VDD.n245 VDD.n244 3.1505
R33 VDD.n242 VDD.n241 3.1505
R34 VDD.n240 VDD.n239 3.1505
R35 VDD.n238 VDD.n237 3.1505
R36 VDD.n236 VDD.n235 3.1505
R37 VDD.n234 VDD.n233 3.1505
R38 VDD.n232 VDD.n231 3.1505
R39 VDD.n230 VDD.n229 3.1505
R40 VDD.n228 VDD.n227 3.1505
R41 VDD.n226 VDD.n225 3.1505
R42 VDD.n223 VDD.n222 3.1505
R43 VDD.n221 VDD.n220 3.1505
R44 VDD.n219 VDD.n218 3.1505
R45 VDD.n284 VDD.n283 3.1505
R46 VDD.n216 VDD.n215 3.1505
R47 VDD.n28 VDD.n27 3.1505
R48 VDD.n26 VDD.n25 3.1505
R49 VDD.n24 VDD.n23 3.1505
R50 VDD.n22 VDD.n21 3.1505
R51 VDD.n20 VDD.n19 3.1505
R52 VDD.n18 VDD.n17 3.1505
R53 VDD.n16 VDD.n15 3.1505
R54 VDD.n14 VDD.n13 3.1505
R55 VDD.n12 VDD.n11 3.1505
R56 VDD.n10 VDD.n9 3.1505
R57 VDD.n8 VDD.n7 3.1505
R58 VDD.n6 VDD.n5 3.1505
R59 VDD.n4 VDD.n3 3.1505
R60 VDD.n169 VDD.n168 3.1505
R61 VDD.n173 VDD.n172 3.1505
R62 VDD.n177 VDD.n176 3.1505
R63 VDD.n181 VDD.n180 3.1505
R64 VDD.n347 VDD.n346 3.1505
R65 VDD.n343 VDD.n342 3.1505
R66 VDD.n339 VDD.n338 3.1505
R67 VDD.n190 VDD.n189 3.1505
R68 VDD.n192 VDD.n191 3.1505
R69 VDD.n194 VDD.n193 3.1505
R70 VDD.n196 VDD.n195 3.1505
R71 VDD.n198 VDD.n197 3.1505
R72 VDD.n200 VDD.n199 3.1505
R73 VDD.n202 VDD.n201 3.1505
R74 VDD.n204 VDD.n203 3.1505
R75 VDD.n206 VDD.n205 3.1505
R76 VDD.n208 VDD.n207 3.1505
R77 VDD.n210 VDD.n209 3.1505
R78 VDD.n212 VDD.n211 3.1505
R79 VDD.n214 VDD.n213 3.1505
R80 VDD.n30 VDD.n29 3.1505
R81 VDD.n32 VDD.n31 3.1505
R82 VDD.n34 VDD.n33 3.1505
R83 VDD.n36 VDD.n35 3.1505
R84 VDD.n38 VDD.n37 3.1505
R85 VDD.n41 VDD.n40 3.1505
R86 VDD.n43 VDD.n42 3.1505
R87 VDD.n45 VDD.n44 3.1505
R88 VDD.n47 VDD.n46 3.1505
R89 VDD.n49 VDD.n48 3.1505
R90 VDD.n51 VDD.n50 3.1505
R91 VDD.n53 VDD.n52 3.1505
R92 VDD.n55 VDD.n54 3.1505
R93 VDD.n58 VDD.n57 3.1505
R94 VDD.n62 VDD.n61 3.1505
R95 VDD.n65 VDD.n64 3.1505
R96 VDD.n68 VDD.n67 3.1505
R97 VDD.n72 VDD.n71 3.1505
R98 VDD.n75 VDD.n74 3.1505
R99 VDD.n78 VDD.n77 3.1505
R100 VDD.n81 VDD.n80 3.1505
R101 VDD.n84 VDD.n83 3.1505
R102 VDD.n87 VDD.n86 3.1505
R103 VDD.n90 VDD.n89 3.1505
R104 VDD.n93 VDD.n92 3.1505
R105 VDD.n96 VDD.n95 3.1505
R106 VDD.n99 VDD.n98 3.1505
R107 VDD.n103 VDD.n102 3.1505
R108 VDD.n106 VDD.n105 3.1505
R109 VDD.n109 VDD.n108 3.1505
R110 VDD.n112 VDD.n111 3.1505
R111 VDD.n128 VDD.n127 3.1505
R112 VDD.n131 VDD.n130 3.1505
R113 VDD.n130 VDD.n129 3.1505
R114 VDD.n134 VDD.n133 3.1505
R115 VDD.n133 VDD.n132 3.1505
R116 VDD.n137 VDD.n136 3.1505
R117 VDD.n136 VDD.n135 3.1505
R118 VDD.n140 VDD.n139 3.1505
R119 VDD.n139 VDD.n138 3.1505
R120 VDD.n143 VDD.n142 3.1505
R121 VDD.n142 VDD.n141 3.1505
R122 VDD.n146 VDD.n145 3.1505
R123 VDD.n145 VDD.n144 3.1505
R124 VDD.n149 VDD.n148 3.1505
R125 VDD.n148 VDD.n147 3.1505
R126 VDD.n152 VDD.n151 3.1505
R127 VDD.n151 VDD.n150 3.1505
R128 VDD.n155 VDD.n154 3.1505
R129 VDD.n154 VDD.n153 3.1505
R130 VDD.n158 VDD.n157 3.1505
R131 VDD.n157 VDD.n156 3.1505
R132 VDD.n161 VDD.n160 3.1505
R133 VDD.n160 VDD.n159 3.1505
R134 VDD.n164 VDD.n163 3.1505
R135 VDD.n163 VDD.n162 3.1505
R136 VDD.n167 VDD.n166 3.1505
R137 VDD.n166 VDD.n165 3.1505
R138 VDD.n171 VDD.n170 3.1505
R139 VDD.n170 VDD.n169 3.1505
R140 VDD.n175 VDD.n174 3.1505
R141 VDD.n174 VDD.n173 3.1505
R142 VDD.n179 VDD.n178 3.1505
R143 VDD.n178 VDD.n177 3.1505
R144 VDD.n183 VDD.n182 3.1505
R145 VDD.n182 VDD.n181 3.1505
R146 VDD.n349 VDD.n348 3.1505
R147 VDD.n348 VDD.n347 3.1505
R148 VDD.n345 VDD.n344 3.1505
R149 VDD.n344 VDD.n343 3.1505
R150 VDD.n341 VDD.n340 3.1505
R151 VDD.n340 VDD.n339 3.1505
R152 VDD.n337 VDD.n336 3.1505
R153 VDD.n336 VDD.n335 3.1505
R154 VDD.n334 VDD.n333 3.1505
R155 VDD.n333 VDD.n332 3.1505
R156 VDD.n331 VDD.n330 3.1505
R157 VDD.n330 VDD.n329 3.1505
R158 VDD.n328 VDD.n327 3.1505
R159 VDD.n327 VDD.n326 3.1505
R160 VDD.n325 VDD.n324 3.1505
R161 VDD.n324 VDD.n323 3.1505
R162 VDD.n322 VDD.n321 3.1505
R163 VDD.n321 VDD.n320 3.1505
R164 VDD.n319 VDD.n318 3.1505
R165 VDD.n318 VDD.n317 3.1505
R166 VDD.n316 VDD.n315 3.1505
R167 VDD.n315 VDD.n314 3.1505
R168 VDD.n313 VDD.n312 3.1505
R169 VDD.n312 VDD.n311 3.1505
R170 VDD.n310 VDD.n309 3.1505
R171 VDD.n309 VDD.n308 3.1505
R172 VDD.n307 VDD.n306 3.1505
R173 VDD.n306 VDD.n305 3.1505
R174 VDD.n304 VDD.n303 3.1505
R175 VDD.n303 VDD.n302 3.1505
R176 VDD.n301 VDD.n300 3.1505
R177 VDD.n300 VDD.n299 3.1505
R178 VDD.n298 VDD.n297 3.1505
R179 VDD.n111 VDD.n110 2.39402
R180 VDD.n108 VDD.n107 2.39402
R181 VDD.n105 VDD.n104 2.39402
R182 VDD.n102 VDD.n101 2.39402
R183 VDD.n98 VDD.n97 2.39402
R184 VDD.n95 VDD.n94 2.39402
R185 VDD.n92 VDD.n91 2.39402
R186 VDD.n89 VDD.n88 2.39402
R187 VDD.n86 VDD.n85 2.39402
R188 VDD.n83 VDD.n82 2.39402
R189 VDD.n80 VDD.n79 2.39402
R190 VDD.n77 VDD.n76 2.39402
R191 VDD.n74 VDD.n73 2.39402
R192 VDD.n71 VDD.n70 2.39402
R193 VDD.n67 VDD.n66 2.39402
R194 VDD.n64 VDD.n63 2.39402
R195 VDD.n61 VDD.n60 2.39402
R196 VDD.n57 VDD.n56 2.39402
R197 VDD.n125 VDD.n114 1.95449
R198 VDD.n125 VDD.n115 1.95449
R199 VDD.n125 VDD.n116 1.95449
R200 VDD.n125 VDD.n117 1.95449
R201 VDD.n125 VDD.n118 1.95449
R202 VDD.n125 VDD.n119 1.95449
R203 VDD.n125 VDD.n120 1.95449
R204 VDD.n125 VDD.n121 1.95449
R205 VDD.n125 VDD.n122 1.95449
R206 VDD.n125 VDD.n123 1.95449
R207 VDD.n125 VDD.n124 1.95449
R208 VDD.n281 VDD.n280 1.73527
R209 VDD.n276 VDD.n275 1.73527
R210 VDD.n270 VDD.n269 1.73527
R211 VDD.n265 VDD.n264 1.73527
R212 VDD.n260 VDD.n259 1.73527
R213 VDD.n126 VDD.n125 1.4169
R214 VDD.n125 VDD.n113 1.41673
R215 VDD.n297 VDD.n296 1.32491
R216 VDD.n127 VDD.n126 1.02761
R217 VDD.n295 VDD.n294 0.914044
R218 VDD.n296 VDD.n295 0.914044
R219 VDD.n295 VDD.n293 0.708865
R220 VDD.n295 VDD.n292 0.708865
R221 VDD.n295 VDD.n291 0.708865
R222 VDD.n295 VDD.n290 0.708865
R223 VDD.n295 VDD.n289 0.708865
R224 VDD.n295 VDD.n288 0.708865
R225 VDD.n295 VDD.n287 0.708865
R226 VDD.n295 VDD.n286 0.708865
R227 VDD.n295 VDD.n285 0.708865
R228 VDD.n156 VDD.t11 0.622004
R229 VDD.n308 VDD.t5 0.622004
R230 VDD.n112 VDD.n109 0.11075
R231 VDD.n109 VDD.n106 0.11075
R232 VDD.n106 VDD.n103 0.11075
R233 VDD.n99 VDD.n96 0.11075
R234 VDD.n96 VDD.n93 0.11075
R235 VDD.n93 VDD.n90 0.11075
R236 VDD.n90 VDD.n87 0.11075
R237 VDD.n87 VDD.n84 0.11075
R238 VDD.n84 VDD.n81 0.11075
R239 VDD.n81 VDD.n78 0.11075
R240 VDD.n78 VDD.n75 0.11075
R241 VDD.n75 VDD.n72 0.11075
R242 VDD.n68 VDD.n65 0.11075
R243 VDD.n65 VDD.n62 0.11075
R244 VDD.n58 VDD.n55 0.11075
R245 VDD.n55 VDD.n53 0.11075
R246 VDD.n53 VDD.n51 0.11075
R247 VDD.n51 VDD.n49 0.11075
R248 VDD.n49 VDD.n47 0.11075
R249 VDD.n47 VDD.n45 0.11075
R250 VDD.n45 VDD.n43 0.11075
R251 VDD.n43 VDD.n41 0.11075
R252 VDD.n38 VDD.n36 0.11075
R253 VDD.n36 VDD.n34 0.11075
R254 VDD.n34 VDD.n32 0.11075
R255 VDD.n30 VDD.n28 0.11075
R256 VDD.n28 VDD.n26 0.11075
R257 VDD.n26 VDD.n24 0.11075
R258 VDD.n24 VDD.n22 0.11075
R259 VDD.n22 VDD.n20 0.11075
R260 VDD.n20 VDD.n18 0.11075
R261 VDD.n18 VDD.n16 0.11075
R262 VDD.n16 VDD.n14 0.11075
R263 VDD.n14 VDD.n12 0.11075
R264 VDD.n12 VDD.n10 0.11075
R265 VDD.n10 VDD.n8 0.11075
R266 VDD.n8 VDD.n6 0.11075
R267 VDD.n6 VDD.n4 0.11075
R268 VDD.n4 VDD.n2 0.11075
R269 VDD.n2 VDD.n1 0.11075
R270 VDD.n1 VDD.n0 0.11075
R271 VDD.n186 VDD.n185 0.11075
R272 VDD.n187 VDD.n186 0.11075
R273 VDD.n188 VDD.n187 0.11075
R274 VDD.n190 VDD.n188 0.11075
R275 VDD.n192 VDD.n190 0.11075
R276 VDD.n194 VDD.n192 0.11075
R277 VDD.n196 VDD.n194 0.11075
R278 VDD.n198 VDD.n196 0.11075
R279 VDD.n200 VDD.n198 0.11075
R280 VDD.n202 VDD.n200 0.11075
R281 VDD.n204 VDD.n202 0.11075
R282 VDD.n206 VDD.n204 0.11075
R283 VDD.n208 VDD.n206 0.11075
R284 VDD.n210 VDD.n208 0.11075
R285 VDD.n212 VDD.n210 0.11075
R286 VDD.n214 VDD.n212 0.11075
R287 VDD.n284 VDD.n282 0.11075
R288 VDD.n282 VDD.n279 0.11075
R289 VDD.n279 VDD.n277 0.11075
R290 VDD.n273 VDD.n271 0.11075
R291 VDD.n271 VDD.n268 0.11075
R292 VDD.n268 VDD.n266 0.11075
R293 VDD.n266 VDD.n263 0.11075
R294 VDD.n263 VDD.n261 0.11075
R295 VDD.n261 VDD.n258 0.11075
R296 VDD.n258 VDD.n256 0.11075
R297 VDD.n256 VDD.n254 0.11075
R298 VDD.n254 VDD.n252 0.11075
R299 VDD.n249 VDD.n247 0.11075
R300 VDD.n247 VDD.n245 0.11075
R301 VDD.n242 VDD.n240 0.11075
R302 VDD.n240 VDD.n238 0.11075
R303 VDD.n238 VDD.n236 0.11075
R304 VDD.n236 VDD.n234 0.11075
R305 VDD.n234 VDD.n232 0.11075
R306 VDD.n232 VDD.n230 0.11075
R307 VDD.n230 VDD.n228 0.11075
R308 VDD.n228 VDD.n226 0.11075
R309 VDD.n223 VDD.n221 0.11075
R310 VDD.n221 VDD.n219 0.11075
R311 VDD.n219 VDD.n217 0.11075
R312 VDD.n217 VDD.n216 0.11075
R313 VDD.n131 VDD.n128 0.11075
R314 VDD.n134 VDD.n131 0.11075
R315 VDD.n137 VDD.n134 0.11075
R316 VDD.n140 VDD.n137 0.11075
R317 VDD.n143 VDD.n140 0.11075
R318 VDD.n146 VDD.n143 0.11075
R319 VDD.n149 VDD.n146 0.11075
R320 VDD.n152 VDD.n149 0.11075
R321 VDD.n155 VDD.n152 0.11075
R322 VDD.n158 VDD.n155 0.11075
R323 VDD.n161 VDD.n158 0.11075
R324 VDD.n164 VDD.n161 0.11075
R325 VDD.n167 VDD.n164 0.11075
R326 VDD.n171 VDD.n167 0.11075
R327 VDD.n175 VDD.n171 0.11075
R328 VDD.n179 VDD.n175 0.11075
R329 VDD.n183 VDD.n179 0.11075
R330 VDD.n349 VDD.n345 0.11075
R331 VDD.n345 VDD.n341 0.11075
R332 VDD.n341 VDD.n337 0.11075
R333 VDD.n337 VDD.n334 0.11075
R334 VDD.n334 VDD.n331 0.11075
R335 VDD.n331 VDD.n328 0.11075
R336 VDD.n328 VDD.n325 0.11075
R337 VDD.n325 VDD.n322 0.11075
R338 VDD.n322 VDD.n319 0.11075
R339 VDD.n319 VDD.n316 0.11075
R340 VDD.n316 VDD.n313 0.11075
R341 VDD.n313 VDD.n310 0.11075
R342 VDD.n310 VDD.n307 0.11075
R343 VDD.n307 VDD.n304 0.11075
R344 VDD.n304 VDD.n301 0.11075
R345 VDD.n301 VDD.n298 0.11075
R346 VDD.n69 VDD.n68 0.1085
R347 VDD.n250 VDD.n249 0.107375
R348 VDD.n103 VDD.n100 0.089375
R349 VDD.n277 VDD.n274 0.087125
R350 VDD VDD.n183 0.0815
R351 VDD.n243 VDD.n242 0.071375
R352 VDD.n59 VDD.n58 0.07025
R353 VDD.n226 VDD.n224 0.066875
R354 VDD.n128 VDD.n112 0.06575
R355 VDD.n32 VDD.n30 0.06575
R356 VDD.n216 VDD.n214 0.06575
R357 VDD.n298 VDD.n284 0.06575
R358 VDD.n41 VDD.n39 0.0635
R359 VDD.n39 VDD.n38 0.04775
R360 VDD.n224 VDD.n223 0.044375
R361 VDD.n62 VDD.n59 0.041
R362 VDD.n245 VDD.n243 0.039875
R363 VDD VDD.n349 0.02975
R364 VDD.n274 VDD.n273 0.024125
R365 VDD.n100 VDD.n99 0.021875
R366 VDD.n252 VDD.n250 0.003875
R367 VDD.n72 VDD.n69 0.00275
R368 COMMON.n0 COMMON.t11 6.48297
R369 COMMON.n0 COMMON.t12 6.48297
R370 COMMON.n1 COMMON.t5 6.48297
R371 COMMON.n1 COMMON.t15 6.48297
R372 COMMON.n2 COMMON.t0 6.48297
R373 COMMON.n2 COMMON.t2 6.48297
R374 COMMON.n4 COMMON.t10 6.48297
R375 COMMON.n4 COMMON.t13 6.48297
R376 COMMON.n5 COMMON.t7 6.48297
R377 COMMON.n5 COMMON.t3 6.48297
R378 COMMON.n6 COMMON.t1 6.48297
R379 COMMON.n6 COMMON.t4 6.48297
R380 COMMON.n3 COMMON.t9 6.48265
R381 COMMON.n3 COMMON.t6 6.48265
R382 COMMON.n8 COMMON.t8 3.35666
R383 COMMON.n9 COMMON.t14 3.1864
R384 COMMON COMMON.n8 0.484053
R385 COMMON COMMON.n9 0.48098
R386 COMMON.n1 COMMON.n0 0.0465976
R387 COMMON.n2 COMMON.n1 0.0465976
R388 COMMON.n4 COMMON.n3 0.0465976
R389 COMMON.n5 COMMON.n4 0.0465976
R390 COMMON.n6 COMMON.n5 0.0465976
R391 COMMON.n7 COMMON.n6 0.0465976
R392 COMMON.n8 COMMON.n7 0.0464286
R393 COMMON.n3 COMMON.n2 0.0460488
R394 R1_IN.n1 R1_IN.t6 6.66964
R395 R1_IN.n0 R1_IN.t2 6.66964
R396 R1_IN.n3 R1_IN.t1 6.50903
R397 R1_IN R1_IN.t5 6.45911
R398 R1_IN.n2 R1_IN.t7 6.44761
R399 R1_IN.n1 R1_IN.t0 6.44761
R400 R1_IN.n8 R1_IN.t4 6.44761
R401 R1_IN.n0 R1_IN.t3 6.44761
R402 R1_IN.n4 R1_IN.n3 0.992758
R403 R1_IN.n7 R1_IN.n6 0.607189
R404 R1_IN.n2 R1_IN.n1 0.222526
R405 R1_IN.n7 R1_IN.n0 0.20072
R406 R1_IN.n3 R1_IN.n2 0.153317
R407 R1_IN R1_IN.n11 0.0813811
R408 R1_IN.n6 R1_IN.n5 0.0441123
R409 R1_IN.n10 R1_IN.n9 0.0441123
R410 R1_IN.n11 R1_IN.n10 0.0441123
R411 R1_IN.n9 R1_IN.n8 0.0429229
R412 R1_IN.n8 R1_IN.n7 0.0234786
R413 R1_IN.n5 R1_IN.n4 0.0195308
R414 R2_IN.n1 R2_IN.t1 6.66924
R415 R2_IN.n11 R2_IN.t7 6.51899
R416 R2_IN.n0 R2_IN.t5 6.49915
R417 R2_IN.n3 R2_IN.t0 6.44775
R418 R2_IN.n1 R2_IN.t4 6.44775
R419 R2_IN.n12 R2_IN.t3 6.44761
R420 R2_IN.n13 R2_IN.t2 6.44761
R421 R2_IN.n14 R2_IN.t6 6.44761
R422 R2_IN.n5 R2_IN.n2 1.16911
R423 R2_IN.n10 R2_IN.n0 1.15365
R424 R2_IN.n9 R2_IN.n8 1.1255
R425 R2_IN.n7 R2_IN.n6 1.1255
R426 R2_IN.n5 R2_IN.n4 1.1255
R427 R2_IN.n11 R2_IN.n10 0.997873
R428 R2_IN.n13 R2_IN.n12 0.222526
R429 R2_IN.n14 R2_IN.n13 0.222526
R430 R2_IN.n2 R2_IN.n1 0.181293
R431 R2_IN.n12 R2_IN.n11 0.141548
R432 R2_IN.n9 R2_IN.n7 0.0441123
R433 R2_IN.n7 R2_IN.n5 0.0441123
R434 R2_IN R2_IN.n14 0.0183414
R435 R2_IN.n10 R2_IN.n9 0.0159626
R436 R2_IN.n4 R2_IN.n3 0.00287885
C0 VDD COMMON 2.88f
C1 R1_IN R2_IN 3.53f
C2 VDD R1_IN 3.03f
C3 R1_IN COMMON 0.531f
C4 VDD R2_IN 3.42f
C5 COMMON R2_IN 0.419f
C6 R2_IN VSUBS 1.23f
C7 COMMON VSUBS 1.52f
C8 R1_IN VSUBS 1.44f
C9 VDD VSUBS 36.6f
C10 R2_IN.t6 VSUBS 0.0565f
C11 R2_IN.t2 VSUBS 0.0565f
C12 R2_IN.t3 VSUBS 0.0565f
C13 R2_IN.t5 VSUBS 0.0598f
C14 R2_IN.n0 VSUBS 0.409f
C15 R2_IN.t4 VSUBS 0.0565f
C16 R2_IN.t1 VSUBS 0.0702f
C17 R2_IN.n1 VSUBS 0.918f
C18 R2_IN.n2 VSUBS 0.238f
C19 R2_IN.t0 VSUBS 0.0565f
C20 R2_IN.n3 VSUBS 0.141f
C21 R2_IN.n4 VSUBS 0.0486f
C22 R2_IN.n5 VSUBS 0.173f
C23 R2_IN.n6 VSUBS 0.0921f
C24 R2_IN.n7 VSUBS 0.0921f
C25 R2_IN.n8 VSUBS 0.0921f
C26 R2_IN.n9 VSUBS 0.0624f
C27 R2_IN.n10 VSUBS 1.2f
C28 R2_IN.t7 VSUBS 0.0599f
C29 R2_IN.n11 VSUBS 1.45f
C30 R2_IN.n12 VSUBS 0.528f
C31 R2_IN.n13 VSUBS 0.564f
C32 R2_IN.n14 VSUBS 0.349f
C33 R1_IN.t4 VSUBS 0.0532f
C34 R1_IN.t3 VSUBS 0.0532f
C35 R1_IN.t2 VSUBS 0.0662f
C36 R1_IN.n0 VSUBS 0.888f
C37 R1_IN.t7 VSUBS 0.0532f
C38 R1_IN.t0 VSUBS 0.0532f
C39 R1_IN.t6 VSUBS 0.0662f
C40 R1_IN.n1 VSUBS 0.907f
C41 R1_IN.n2 VSUBS 0.497f
C42 R1_IN.t1 VSUBS 0.0559f
C43 R1_IN.n3 VSUBS 1.33f
C44 R1_IN.n4 VSUBS 1.12f
C45 R1_IN.n5 VSUBS 0.0623f
C46 R1_IN.n6 VSUBS 0.279f
C47 R1_IN.n7 VSUBS 0.216f
C48 R1_IN.n8 VSUBS 0.176f
C49 R1_IN.n9 VSUBS 0.0856f
C50 R1_IN.n10 VSUBS 0.0868f
C51 R1_IN.n11 VSUBS 0.125f
C52 R1_IN.t5 VSUBS 0.0536f
C53 COMMON.t11 VSUBS 0.0414f
C54 COMMON.t12 VSUBS 0.0414f
C55 COMMON.n0 VSUBS 0.236f
C56 COMMON.t5 VSUBS 0.0414f
C57 COMMON.t15 VSUBS 0.0414f
C58 COMMON.n1 VSUBS 0.254f
C59 COMMON.t0 VSUBS 0.0414f
C60 COMMON.t2 VSUBS 0.0414f
C61 COMMON.n2 VSUBS 0.254f
C62 COMMON.t6 VSUBS 0.0414f
C63 COMMON.t9 VSUBS 0.0414f
C64 COMMON.n3 VSUBS 0.255f
C65 COMMON.t10 VSUBS 0.0414f
C66 COMMON.t13 VSUBS 0.0414f
C67 COMMON.n4 VSUBS 0.254f
C68 COMMON.t7 VSUBS 0.0414f
C69 COMMON.t3 VSUBS 0.0414f
C70 COMMON.n5 VSUBS 0.254f
C71 COMMON.t1 VSUBS 0.0414f
C72 COMMON.t4 VSUBS 0.0414f
C73 COMMON.n6 VSUBS 0.254f
C74 COMMON.n7 VSUBS 0.0905f
C75 COMMON.t8 VSUBS 0.0289f
C76 COMMON.n8 VSUBS 0.096f
C77 COMMON.t14 VSUBS 0.0283f
C78 COMMON.n9 VSUBS 0.114f
C79 VDD.t9 VSUBS 0.0114f
C80 VDD.t10 VSUBS 0.0114f
C81 VDD.t3 VSUBS 0.0114f
C82 VDD.t4 VSUBS 0.0114f
C83 VDD.n0 VSUBS 0.00532f
C84 VDD.n1 VSUBS 0.00532f
C85 VDD.n2 VSUBS 0.00532f
C86 VDD.n3 VSUBS 0.00532f
C87 VDD.n4 VSUBS 0.00532f
C88 VDD.n5 VSUBS 0.00532f
C89 VDD.n6 VSUBS 0.00532f
C90 VDD.n7 VSUBS 0.00532f
C91 VDD.n8 VSUBS 0.00532f
C92 VDD.n9 VSUBS 0.00532f
C93 VDD.n10 VSUBS 0.00532f
C94 VDD.n11 VSUBS 0.00532f
C95 VDD.n12 VSUBS 0.00532f
C96 VDD.n13 VSUBS 0.00532f
C97 VDD.n14 VSUBS 0.00532f
C98 VDD.n15 VSUBS 0.00532f
C99 VDD.n16 VSUBS 0.00532f
C100 VDD.n17 VSUBS 0.00532f
C101 VDD.n18 VSUBS 0.00532f
C102 VDD.n19 VSUBS 0.00532f
C103 VDD.n20 VSUBS 0.00532f
C104 VDD.n21 VSUBS 0.00532f
C105 VDD.n22 VSUBS 0.00532f
C106 VDD.n23 VSUBS 0.00532f
C107 VDD.n24 VSUBS 0.00532f
C108 VDD.n25 VSUBS 0.00532f
C109 VDD.n26 VSUBS 0.00532f
C110 VDD.n27 VSUBS 0.00532f
C111 VDD.n28 VSUBS 0.00532f
C112 VDD.n29 VSUBS 0.0064f
C113 VDD.n30 VSUBS 0.0064f
C114 VDD.n31 VSUBS 0.00423f
C115 VDD.n32 VSUBS 0.00423f
C116 VDD.n33 VSUBS 0.00532f
C117 VDD.n34 VSUBS 0.00532f
C118 VDD.n35 VSUBS 0.00532f
C119 VDD.n36 VSUBS 0.00532f
C120 VDD.n37 VSUBS 0.00532f
C121 VDD.n38 VSUBS 0.0038f
C122 VDD.n39 VSUBS 0.0263f
C123 VDD.n40 VSUBS 0.00532f
C124 VDD.n41 VSUBS 0.00418f
C125 VDD.n42 VSUBS 0.00532f
C126 VDD.n43 VSUBS 0.00532f
C127 VDD.n44 VSUBS 0.00532f
C128 VDD.n45 VSUBS 0.00532f
C129 VDD.n46 VSUBS 0.00532f
C130 VDD.n47 VSUBS 0.00532f
C131 VDD.n48 VSUBS 0.00532f
C132 VDD.n49 VSUBS 0.00532f
C133 VDD.n50 VSUBS 0.00532f
C134 VDD.n51 VSUBS 0.00532f
C135 VDD.n52 VSUBS 0.00532f
C136 VDD.n53 VSUBS 0.00532f
C137 VDD.n54 VSUBS 0.00532f
C138 VDD.n55 VSUBS 0.00532f
C139 VDD.n57 VSUBS 0.00532f
C140 VDD.n58 VSUBS 0.00434f
C141 VDD.n59 VSUBS 0.0259f
C142 VDD.n61 VSUBS 0.00532f
C143 VDD.n62 VSUBS 0.00363f
C144 VDD.n64 VSUBS 0.00532f
C145 VDD.n65 VSUBS 0.00532f
C146 VDD.n67 VSUBS 0.00532f
C147 VDD.n68 VSUBS 0.00526f
C148 VDD.n69 VSUBS 0.026f
C149 VDD.n71 VSUBS 0.00532f
C150 VDD.n72 VSUBS 0.00271f
C151 VDD.n74 VSUBS 0.00532f
C152 VDD.n75 VSUBS 0.00532f
C153 VDD.n77 VSUBS 0.00532f
C154 VDD.n78 VSUBS 0.00532f
C155 VDD.n80 VSUBS 0.00532f
C156 VDD.n81 VSUBS 0.00532f
C157 VDD.n83 VSUBS 0.00532f
C158 VDD.n84 VSUBS 0.00532f
C159 VDD.n86 VSUBS 0.00532f
C160 VDD.n87 VSUBS 0.00532f
C161 VDD.n89 VSUBS 0.00532f
C162 VDD.n90 VSUBS 0.00532f
C163 VDD.n92 VSUBS 0.00532f
C164 VDD.n93 VSUBS 0.00532f
C165 VDD.n95 VSUBS 0.00532f
C166 VDD.n96 VSUBS 0.00532f
C167 VDD.n98 VSUBS 0.00532f
C168 VDD.n99 VSUBS 0.00317f
C169 VDD.n100 VSUBS 0.0259f
C170 VDD.n102 VSUBS 0.00532f
C171 VDD.n103 VSUBS 0.0048f
C172 VDD.n105 VSUBS 0.00532f
C173 VDD.n106 VSUBS 0.00532f
C174 VDD.n108 VSUBS 0.00532f
C175 VDD.n109 VSUBS 0.00532f
C176 VDD.n111 VSUBS 0.00423f
C177 VDD.n112 VSUBS 0.00423f
C178 VDD.n125 VSUBS 0.303f
C179 VDD.n127 VSUBS 0.0064f
C180 VDD.n128 VSUBS 0.0064f
C181 VDD.n129 VSUBS 0.214f
C182 VDD.n130 VSUBS 0.00532f
C183 VDD.n131 VSUBS 0.00532f
C184 VDD.n132 VSUBS 0.214f
C185 VDD.n133 VSUBS 0.00532f
C186 VDD.n134 VSUBS 0.00532f
C187 VDD.n135 VSUBS 0.214f
C188 VDD.n136 VSUBS 0.00532f
C189 VDD.n137 VSUBS 0.00532f
C190 VDD.t2 VSUBS 0.107f
C191 VDD.n138 VSUBS 0.135f
C192 VDD.n139 VSUBS 0.00532f
C193 VDD.n140 VSUBS 0.00532f
C194 VDD.n141 VSUBS 0.185f
C195 VDD.n142 VSUBS 0.00532f
C196 VDD.n143 VSUBS 0.00532f
C197 VDD.n144 VSUBS 0.214f
C198 VDD.n145 VSUBS 0.00532f
C199 VDD.n146 VSUBS 0.00532f
C200 VDD.t15 VSUBS 0.107f
C201 VDD.n147 VSUBS 0.12f
C202 VDD.n148 VSUBS 0.00532f
C203 VDD.n149 VSUBS 0.00532f
C204 VDD.n150 VSUBS 0.201f
C205 VDD.n151 VSUBS 0.00532f
C206 VDD.n152 VSUBS 0.00532f
C207 VDD.n153 VSUBS 0.212f
C208 VDD.n154 VSUBS 0.00532f
C209 VDD.n155 VSUBS 0.00532f
C210 VDD.t11 VSUBS 0.107f
C211 VDD.n156 VSUBS 0.109f
C212 VDD.n157 VSUBS 0.00532f
C213 VDD.n158 VSUBS 0.00532f
C214 VDD.n159 VSUBS 0.214f
C215 VDD.n160 VSUBS 0.00532f
C216 VDD.n161 VSUBS 0.00532f
C217 VDD.n162 VSUBS 0.196f
C218 VDD.n163 VSUBS 0.00532f
C219 VDD.n164 VSUBS 0.00532f
C220 VDD.t0 VSUBS 0.107f
C221 VDD.n165 VSUBS 0.124f
C222 VDD.n166 VSUBS 0.00532f
C223 VDD.n167 VSUBS 0.00532f
C224 VDD.n168 VSUBS 0.00532f
C225 VDD.n169 VSUBS 0.214f
C226 VDD.n170 VSUBS 0.00532f
C227 VDD.n171 VSUBS 0.00532f
C228 VDD.n172 VSUBS 0.00532f
C229 VDD.n173 VSUBS 0.181f
C230 VDD.n174 VSUBS 0.00532f
C231 VDD.n175 VSUBS 0.00532f
C232 VDD.t12 VSUBS 0.107f
C233 VDD.n176 VSUBS 0.00532f
C234 VDD.n177 VSUBS 0.14f
C235 VDD.n178 VSUBS 0.00532f
C236 VDD.n179 VSUBS 0.00532f
C237 VDD.n180 VSUBS 0.00532f
C238 VDD.n181 VSUBS 0.214f
C239 VDD.n182 VSUBS 0.00532f
C240 VDD.n183 VSUBS 0.00461f
C241 VDD.t16 VSUBS 0.011f
C242 VDD.t17 VSUBS 0.0109f
C243 VDD.t6 VSUBS 0.011f
C244 VDD.t7 VSUBS 0.011f
C245 VDD.n184 VSUBS 0.00423f
C246 VDD.n185 VSUBS 0.00532f
C247 VDD.n186 VSUBS 0.00532f
C248 VDD.n187 VSUBS 0.00532f
C249 VDD.n188 VSUBS 0.00532f
C250 VDD.n189 VSUBS 0.00532f
C251 VDD.n190 VSUBS 0.00532f
C252 VDD.n191 VSUBS 0.00532f
C253 VDD.n192 VSUBS 0.00532f
C254 VDD.n193 VSUBS 0.00532f
C255 VDD.n194 VSUBS 0.00532f
C256 VDD.n195 VSUBS 0.00532f
C257 VDD.n196 VSUBS 0.00532f
C258 VDD.n197 VSUBS 0.00532f
C259 VDD.n198 VSUBS 0.00532f
C260 VDD.n199 VSUBS 0.00532f
C261 VDD.n200 VSUBS 0.00532f
C262 VDD.n201 VSUBS 0.00532f
C263 VDD.n202 VSUBS 0.00532f
C264 VDD.n203 VSUBS 0.00532f
C265 VDD.n204 VSUBS 0.00532f
C266 VDD.n205 VSUBS 0.00532f
C267 VDD.n206 VSUBS 0.00532f
C268 VDD.n207 VSUBS 0.00532f
C269 VDD.n208 VSUBS 0.00532f
C270 VDD.n209 VSUBS 0.00532f
C271 VDD.n210 VSUBS 0.00532f
C272 VDD.n211 VSUBS 0.00532f
C273 VDD.n212 VSUBS 0.00532f
C274 VDD.n213 VSUBS 0.00532f
C275 VDD.n214 VSUBS 0.00423f
C276 VDD.n215 VSUBS 0.0064f
C277 VDD.n216 VSUBS 0.0064f
C278 VDD.n217 VSUBS 0.00532f
C279 VDD.n218 VSUBS 0.00532f
C280 VDD.n219 VSUBS 0.00532f
C281 VDD.n220 VSUBS 0.00532f
C282 VDD.n221 VSUBS 0.00532f
C283 VDD.n222 VSUBS 0.00532f
C284 VDD.n223 VSUBS 0.00372f
C285 VDD.n224 VSUBS 0.0203f
C286 VDD.n225 VSUBS 0.00532f
C287 VDD.n226 VSUBS 0.00426f
C288 VDD.n227 VSUBS 0.00532f
C289 VDD.n228 VSUBS 0.00532f
C290 VDD.n229 VSUBS 0.00532f
C291 VDD.n230 VSUBS 0.00532f
C292 VDD.n231 VSUBS 0.00532f
C293 VDD.n232 VSUBS 0.00532f
C294 VDD.n233 VSUBS 0.00532f
C295 VDD.n234 VSUBS 0.00532f
C296 VDD.n235 VSUBS 0.00532f
C297 VDD.n236 VSUBS 0.00532f
C298 VDD.n237 VSUBS 0.00532f
C299 VDD.n238 VSUBS 0.00532f
C300 VDD.n239 VSUBS 0.00532f
C301 VDD.n240 VSUBS 0.00532f
C302 VDD.n241 VSUBS 0.00532f
C303 VDD.n242 VSUBS 0.00437f
C304 VDD.n243 VSUBS 0.0206f
C305 VDD.n244 VSUBS 0.00532f
C306 VDD.n245 VSUBS 0.00361f
C307 VDD.n246 VSUBS 0.00532f
C308 VDD.n247 VSUBS 0.00532f
C309 VDD.n248 VSUBS 0.00532f
C310 VDD.n249 VSUBS 0.00524f
C311 VDD.n250 VSUBS 0.0199f
C312 VDD.n251 VSUBS 0.00532f
C313 VDD.n252 VSUBS 0.00274f
C314 VDD.n253 VSUBS 0.00532f
C315 VDD.n254 VSUBS 0.00532f
C316 VDD.n255 VSUBS 0.00532f
C317 VDD.n256 VSUBS 0.00532f
C318 VDD.n257 VSUBS 0.00532f
C319 VDD.n258 VSUBS 0.00532f
C320 VDD.n260 VSUBS 0.00532f
C321 VDD.n261 VSUBS 0.00532f
C322 VDD.n262 VSUBS 0.00532f
C323 VDD.n263 VSUBS 0.00532f
C324 VDD.n265 VSUBS 0.00532f
C325 VDD.n266 VSUBS 0.00532f
C326 VDD.n267 VSUBS 0.00532f
C327 VDD.n268 VSUBS 0.00532f
C328 VDD.n270 VSUBS 0.00532f
C329 VDD.n271 VSUBS 0.00532f
C330 VDD.n272 VSUBS 0.00532f
C331 VDD.n273 VSUBS 0.00323f
C332 VDD.n274 VSUBS 0.0208f
C333 VDD.n276 VSUBS 0.00532f
C334 VDD.n277 VSUBS 0.00475f
C335 VDD.n278 VSUBS 0.00532f
C336 VDD.n279 VSUBS 0.00532f
C337 VDD.n281 VSUBS 0.00532f
C338 VDD.n282 VSUBS 0.00532f
C339 VDD.n283 VSUBS 0.00423f
C340 VDD.n284 VSUBS 0.00423f
C341 VDD.n295 VSUBS 0.303f
C342 VDD.n297 VSUBS 0.0064f
C343 VDD.n298 VSUBS 0.0064f
C344 VDD.n299 VSUBS 0.214f
C345 VDD.n300 VSUBS 0.00532f
C346 VDD.n301 VSUBS 0.00532f
C347 VDD.n302 VSUBS 0.214f
C348 VDD.n303 VSUBS 0.00532f
C349 VDD.n304 VSUBS 0.00532f
C350 VDD.n305 VSUBS 0.214f
C351 VDD.n306 VSUBS 0.00532f
C352 VDD.n307 VSUBS 0.00532f
C353 VDD.t5 VSUBS 0.107f
C354 VDD.n308 VSUBS 0.109f
C355 VDD.n309 VSUBS 0.00532f
C356 VDD.n310 VSUBS 0.00532f
C357 VDD.n311 VSUBS 0.212f
C358 VDD.n312 VSUBS 0.00532f
C359 VDD.n313 VSUBS 0.00532f
C360 VDD.n314 VSUBS 0.201f
C361 VDD.n315 VSUBS 0.00532f
C362 VDD.n316 VSUBS 0.00532f
C363 VDD.t13 VSUBS 0.107f
C364 VDD.n317 VSUBS 0.12f
C365 VDD.n318 VSUBS 0.00532f
C366 VDD.n319 VSUBS 0.00532f
C367 VDD.n320 VSUBS 0.214f
C368 VDD.n321 VSUBS 0.00532f
C369 VDD.n322 VSUBS 0.00532f
C370 VDD.n323 VSUBS 0.185f
C371 VDD.n324 VSUBS 0.00532f
C372 VDD.n325 VSUBS 0.00532f
C373 VDD.t1 VSUBS 0.107f
C374 VDD.n326 VSUBS 0.135f
C375 VDD.n327 VSUBS 0.00532f
C376 VDD.n328 VSUBS 0.00532f
C377 VDD.n329 VSUBS 0.214f
C378 VDD.n330 VSUBS 0.00532f
C379 VDD.n331 VSUBS 0.00532f
C380 VDD.n332 VSUBS 0.17f
C381 VDD.n333 VSUBS 0.00532f
C382 VDD.n334 VSUBS 0.00532f
C383 VDD.t8 VSUBS 0.107f
C384 VDD.n335 VSUBS 0.151f
C385 VDD.n336 VSUBS 0.00532f
C386 VDD.n337 VSUBS 0.00532f
C387 VDD.n338 VSUBS 0.00532f
C388 VDD.n339 VSUBS 0.214f
C389 VDD.n340 VSUBS 0.00532f
C390 VDD.n341 VSUBS 0.00532f
C391 VDD.t14 VSUBS 0.107f
C392 VDD.n342 VSUBS 0.00532f
C393 VDD.n343 VSUBS 0.155f
C394 VDD.n344 VSUBS 0.00532f
C395 VDD.n345 VSUBS 0.00532f
C396 VDD.n346 VSUBS 0.00532f
C397 VDD.n347 VSUBS 0.166f
C398 VDD.n348 VSUBS 0.00532f
C399 VDD.n349 VSUBS 0.00336f
.ends

