magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1435 1019 1435
<< metal2 >>
rect -19 430 19 435
rect -19 -430 -14 430
rect 14 -430 19 430
rect -19 -435 19 -430
<< via2 >>
rect -14 -430 14 430
<< metal3 >>
rect -19 430 19 435
rect -19 -430 -14 430
rect 14 -430 19 430
rect -19 -435 19 -430
<< end >>
