magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -3844 2128 3844
<< nwell >>
rect -128 -1844 128 1844
<< nsubdiff >>
rect -45 1739 45 1761
rect -45 1693 -23 1739
rect 23 1693 45 1739
rect -45 1635 45 1693
rect -45 1589 -23 1635
rect 23 1589 45 1635
rect -45 1531 45 1589
rect -45 1485 -23 1531
rect 23 1485 45 1531
rect -45 1427 45 1485
rect -45 1381 -23 1427
rect 23 1381 45 1427
rect -45 1323 45 1381
rect -45 1277 -23 1323
rect 23 1277 45 1323
rect -45 1219 45 1277
rect -45 1173 -23 1219
rect 23 1173 45 1219
rect -45 1115 45 1173
rect -45 1069 -23 1115
rect 23 1069 45 1115
rect -45 1011 45 1069
rect -45 965 -23 1011
rect 23 965 45 1011
rect -45 907 45 965
rect -45 861 -23 907
rect 23 861 45 907
rect -45 803 45 861
rect -45 757 -23 803
rect 23 757 45 803
rect -45 699 45 757
rect -45 653 -23 699
rect 23 653 45 699
rect -45 595 45 653
rect -45 549 -23 595
rect 23 549 45 595
rect -45 491 45 549
rect -45 445 -23 491
rect 23 445 45 491
rect -45 387 45 445
rect -45 341 -23 387
rect 23 341 45 387
rect -45 283 45 341
rect -45 237 -23 283
rect 23 237 45 283
rect -45 179 45 237
rect -45 133 -23 179
rect 23 133 45 179
rect -45 75 45 133
rect -45 29 -23 75
rect 23 29 45 75
rect -45 -29 45 29
rect -45 -75 -23 -29
rect 23 -75 45 -29
rect -45 -133 45 -75
rect -45 -179 -23 -133
rect 23 -179 45 -133
rect -45 -237 45 -179
rect -45 -283 -23 -237
rect 23 -283 45 -237
rect -45 -341 45 -283
rect -45 -387 -23 -341
rect 23 -387 45 -341
rect -45 -445 45 -387
rect -45 -491 -23 -445
rect 23 -491 45 -445
rect -45 -549 45 -491
rect -45 -595 -23 -549
rect 23 -595 45 -549
rect -45 -653 45 -595
rect -45 -699 -23 -653
rect 23 -699 45 -653
rect -45 -757 45 -699
rect -45 -803 -23 -757
rect 23 -803 45 -757
rect -45 -861 45 -803
rect -45 -907 -23 -861
rect 23 -907 45 -861
rect -45 -965 45 -907
rect -45 -1011 -23 -965
rect 23 -1011 45 -965
rect -45 -1069 45 -1011
rect -45 -1115 -23 -1069
rect 23 -1115 45 -1069
rect -45 -1173 45 -1115
rect -45 -1219 -23 -1173
rect 23 -1219 45 -1173
rect -45 -1277 45 -1219
rect -45 -1323 -23 -1277
rect 23 -1323 45 -1277
rect -45 -1381 45 -1323
rect -45 -1427 -23 -1381
rect 23 -1427 45 -1381
rect -45 -1485 45 -1427
rect -45 -1531 -23 -1485
rect 23 -1531 45 -1485
rect -45 -1589 45 -1531
rect -45 -1635 -23 -1589
rect 23 -1635 45 -1589
rect -45 -1693 45 -1635
rect -45 -1739 -23 -1693
rect 23 -1739 45 -1693
rect -45 -1761 45 -1739
<< nsubdiffcont >>
rect -23 1693 23 1739
rect -23 1589 23 1635
rect -23 1485 23 1531
rect -23 1381 23 1427
rect -23 1277 23 1323
rect -23 1173 23 1219
rect -23 1069 23 1115
rect -23 965 23 1011
rect -23 861 23 907
rect -23 757 23 803
rect -23 653 23 699
rect -23 549 23 595
rect -23 445 23 491
rect -23 341 23 387
rect -23 237 23 283
rect -23 133 23 179
rect -23 29 23 75
rect -23 -75 23 -29
rect -23 -179 23 -133
rect -23 -283 23 -237
rect -23 -387 23 -341
rect -23 -491 23 -445
rect -23 -595 23 -549
rect -23 -699 23 -653
rect -23 -803 23 -757
rect -23 -907 23 -861
rect -23 -1011 23 -965
rect -23 -1115 23 -1069
rect -23 -1219 23 -1173
rect -23 -1323 23 -1277
rect -23 -1427 23 -1381
rect -23 -1531 23 -1485
rect -23 -1635 23 -1589
rect -23 -1739 23 -1693
<< metal1 >>
rect -34 1739 34 1750
rect -34 1693 -23 1739
rect 23 1693 34 1739
rect -34 1635 34 1693
rect -34 1589 -23 1635
rect 23 1589 34 1635
rect -34 1531 34 1589
rect -34 1485 -23 1531
rect 23 1485 34 1531
rect -34 1427 34 1485
rect -34 1381 -23 1427
rect 23 1381 34 1427
rect -34 1323 34 1381
rect -34 1277 -23 1323
rect 23 1277 34 1323
rect -34 1219 34 1277
rect -34 1173 -23 1219
rect 23 1173 34 1219
rect -34 1115 34 1173
rect -34 1069 -23 1115
rect 23 1069 34 1115
rect -34 1011 34 1069
rect -34 965 -23 1011
rect 23 965 34 1011
rect -34 907 34 965
rect -34 861 -23 907
rect 23 861 34 907
rect -34 803 34 861
rect -34 757 -23 803
rect 23 757 34 803
rect -34 699 34 757
rect -34 653 -23 699
rect 23 653 34 699
rect -34 595 34 653
rect -34 549 -23 595
rect 23 549 34 595
rect -34 491 34 549
rect -34 445 -23 491
rect 23 445 34 491
rect -34 387 34 445
rect -34 341 -23 387
rect 23 341 34 387
rect -34 283 34 341
rect -34 237 -23 283
rect 23 237 34 283
rect -34 179 34 237
rect -34 133 -23 179
rect 23 133 34 179
rect -34 75 34 133
rect -34 29 -23 75
rect 23 29 34 75
rect -34 -29 34 29
rect -34 -75 -23 -29
rect 23 -75 34 -29
rect -34 -133 34 -75
rect -34 -179 -23 -133
rect 23 -179 34 -133
rect -34 -237 34 -179
rect -34 -283 -23 -237
rect 23 -283 34 -237
rect -34 -341 34 -283
rect -34 -387 -23 -341
rect 23 -387 34 -341
rect -34 -445 34 -387
rect -34 -491 -23 -445
rect 23 -491 34 -445
rect -34 -549 34 -491
rect -34 -595 -23 -549
rect 23 -595 34 -549
rect -34 -653 34 -595
rect -34 -699 -23 -653
rect 23 -699 34 -653
rect -34 -757 34 -699
rect -34 -803 -23 -757
rect 23 -803 34 -757
rect -34 -861 34 -803
rect -34 -907 -23 -861
rect 23 -907 34 -861
rect -34 -965 34 -907
rect -34 -1011 -23 -965
rect 23 -1011 34 -965
rect -34 -1069 34 -1011
rect -34 -1115 -23 -1069
rect 23 -1115 34 -1069
rect -34 -1173 34 -1115
rect -34 -1219 -23 -1173
rect 23 -1219 34 -1173
rect -34 -1277 34 -1219
rect -34 -1323 -23 -1277
rect 23 -1323 34 -1277
rect -34 -1381 34 -1323
rect -34 -1427 -23 -1381
rect 23 -1427 34 -1381
rect -34 -1485 34 -1427
rect -34 -1531 -23 -1485
rect 23 -1531 34 -1485
rect -34 -1589 34 -1531
rect -34 -1635 -23 -1589
rect 23 -1635 34 -1589
rect -34 -1693 34 -1635
rect -34 -1739 -23 -1693
rect 23 -1739 34 -1693
rect -34 -1750 34 -1739
<< end >>
