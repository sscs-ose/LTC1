magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3470 -2083 8872 4575
<< isosubstrate >>
rect -1470 -83 6872 2575
<< nwell >>
rect 0 1281 6872 2575
<< psubdiff >>
rect 168 0 247 90
<< nsubdiff >>
rect 173 2402 247 2492
<< polysilicon >>
rect 1669 1560 1809 1771
rect 1913 1560 2053 1771
rect 2365 1644 2505 1768
rect 2609 1644 2749 1768
rect 2853 1644 2993 1768
rect 3315 1644 3455 1686
rect 3559 1644 3699 1686
rect 4183 1644 4323 1686
rect 4427 1644 4567 1686
rect 4815 1644 4955 1686
rect 5059 1644 5199 1686
rect 5831 1444 5971 1763
rect 6219 1444 6359 1763
rect 459 724 599 1291
rect 703 724 843 1291
rect 1170 963 1310 1101
rect 1747 963 1887 1101
rect 1991 963 2131 1101
rect 2235 963 2375 1101
rect 2479 963 2619 1101
rect 2723 963 2863 1101
rect 3203 912 3343 1106
rect 3447 912 3587 1106
rect 3691 912 3831 1106
rect 3935 912 4075 1106
rect 4323 912 4463 1120
rect 4567 912 4707 1120
rect 4811 912 4951 1120
rect 5055 912 5195 1120
rect 5831 913 5971 1232
rect 6219 913 6359 1232
rect 5443 477 5583 596
<< metal1 >>
rect 8 2413 148 2489
rect 162 2413 258 2481
rect 8 1581 106 2413
rect 384 2058 430 2419
rect 613 1224 689 2135
rect 872 2058 918 2419
rect 1594 2095 1640 2418
rect 2082 2095 2128 2418
rect 2290 1745 2346 2455
rect 2528 2301 3072 2357
rect 2528 1797 2584 2301
rect 2773 1745 2829 2197
rect 2290 1689 2829 1745
rect 3016 1740 3072 2301
rect 3227 1730 3303 2206
rect 3469 1730 3545 2430
rect 6624 2413 6710 2481
rect 4979 2285 6620 2341
rect 3751 2190 4171 2266
rect 4095 2110 4171 2190
rect 3751 1730 4171 2110
rect 4579 2110 4655 2206
rect 4579 1730 4764 2110
rect 4979 1766 5035 2285
rect 5203 1730 5279 2118
rect 5741 1637 5817 2037
rect 6042 1637 6144 2037
rect 1492 1568 1665 1636
rect 1775 1568 1916 1636
rect 2508 1568 2868 1636
rect 3434 1568 4420 1636
rect 4939 1568 5817 1636
rect 6564 1619 6620 2285
rect 1142 1224 1240 1442
rect 1492 1224 1560 1568
rect 5831 1508 6225 1520
rect 1658 1452 6472 1508
rect 2954 1280 6472 1396
rect 613 1168 1321 1224
rect 1492 1168 6472 1224
rect 8 11 94 1019
rect 495 876 811 1038
rect 905 826 981 1168
rect 1159 1112 1321 1168
rect 5831 1156 6225 1168
rect 615 750 981 826
rect 1508 1044 1740 1112
rect 1893 1044 2719 1112
rect 3247 1044 5044 1112
rect 152 11 259 79
rect 384 72 430 314
rect 615 280 687 750
rect 872 72 918 314
rect 1095 288 1141 623
rect 1339 77 1385 632
rect 1508 135 1576 1044
rect 1672 66 1718 282
rect 1901 217 1977 920
rect 2389 219 2465 920
rect 2877 918 3921 994
rect 2877 219 2953 918
rect 2389 217 2953 219
rect 1901 159 2953 217
rect 3113 235 3189 868
rect 3357 338 3433 918
rect 3601 235 3677 868
rect 3845 338 3921 918
rect 4233 948 5658 994
rect 4233 918 5285 948
rect 4233 868 4309 918
rect 4089 235 4311 868
rect 3113 233 4311 235
rect 4721 233 4797 918
rect 5209 233 5285 918
rect 5612 608 5658 948
rect 5741 751 5817 1031
rect 6042 731 6144 1031
rect 6373 505 6449 866
rect 5570 437 6449 505
rect 3113 159 4165 233
rect 6624 11 6710 79
<< metal2 >>
rect 3227 2190 3726 2266
rect 4095 2042 5279 2118
rect 1177 1442 1647 1518
rect 1150 1168 1672 1244
rect 1150 994 1330 1168
rect 1896 1029 1968 1977
rect 2611 1075 2791 1565
rect 3006 1396 3082 1733
rect 2954 1280 3134 1396
rect 3915 1044 4019 1590
rect 4326 1300 4435 1967
rect 826 918 1330 994
rect 1480 953 1968 1029
rect 1480 485 1556 953
rect 4477 842 4553 1376
rect 4965 842 5041 1353
rect 5364 1052 5468 2252
rect 5555 926 5631 2481
rect 5353 861 5631 926
rect 1719 574 2634 754
rect 5741 485 5817 1672
rect 6005 1006 6185 1637
rect 1480 409 5817 485
rect 6373 349 6449 1672
rect 1217 273 6449 349
rect 6554 15 6630 1632
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_0
timestamp 1713338890
transform 1 0 128 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_1
timestamp 1713338890
transform 1 0 6744 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145318  M1_NWELL_CDNS_40661953145318_0
timestamp 1713338890
transform 1 0 3441 0 1 2447
box -3277 -128 3277 128
use M1_NWELL_CDNS_40661953145320  M1_NWELL_CDNS_40661953145320_0
timestamp 1713338890
transform 1 0 -650 0 1 2031
box -752 -544 752 544
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_0
timestamp 1713338890
transform 1 0 1240 0 1 1078
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_1
timestamp 1713338890
transform 1 0 1817 0 1 1078
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_2
timestamp 1713338890
transform 1 0 2305 0 1 1078
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_3
timestamp 1713338890
transform 1 0 2061 0 1 1078
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_4
timestamp 1713338890
transform 1 0 2549 0 1 1078
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_5
timestamp 1713338890
transform 1 0 2793 0 1 1078
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_6
timestamp 1713338890
transform 1 0 5532 0 1 471
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform 1 0 773 0 -1 957
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform 1 0 529 0 -1 957
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_2
timestamp 1713338890
transform 0 -1 3517 1 0 1078
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_3
timestamp 1713338890
transform 0 -1 3273 1 0 1078
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_4
timestamp 1713338890
transform 0 -1 3761 1 0 1078
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_5
timestamp 1713338890
transform 0 -1 4393 1 0 1078
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_6
timestamp 1713338890
transform 0 -1 4637 1 0 1078
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_7
timestamp 1713338890
transform 0 -1 4005 1 0 1078
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_8
timestamp 1713338890
transform 0 -1 4881 1 0 1078
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_9
timestamp 1713338890
transform 0 -1 5125 1 0 1078
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_10
timestamp 1713338890
transform 0 1 5901 -1 0 1190
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_11
timestamp 1713338890
transform 0 1 6289 -1 0 1190
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_12
timestamp 1713338890
transform 0 -1 2435 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_13
timestamp 1713338890
transform 0 -1 2679 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_14
timestamp 1713338890
transform 0 -1 1739 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_15
timestamp 1713338890
transform 0 -1 1983 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_16
timestamp 1713338890
transform 0 -1 2923 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_17
timestamp 1713338890
transform 0 -1 3385 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_18
timestamp 1713338890
transform 0 -1 3629 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_19
timestamp 1713338890
transform 0 -1 4253 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_20
timestamp 1713338890
transform 0 -1 4497 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_21
timestamp 1713338890
transform 0 -1 4885 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_22
timestamp 1713338890
transform 0 -1 5129 1 0 1602
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_23
timestamp 1713338890
transform 0 1 5901 1 0 1486
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_24
timestamp 1713338890
transform 0 1 6289 1 0 1486
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 1 0 128 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 1 0 6744 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165616  M1_PSUB_CDNS_69033583165616_0
timestamp 1713338890
transform 1 0 -650 0 1 569
box -669 -461 669 461
use M1_PSUB_CDNS_69033583165617  M1_PSUB_CDNS_69033583165617_0
timestamp 1713338890
transform 1 0 3441 0 -1 45
box -3194 -45 3194 45
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_0
timestamp 1713338890
transform 1 0 1582 0 1 1206
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_1
timestamp 1713338890
transform 1 0 2701 0 1 1074
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_2
timestamp 1713338890
transform 1 0 4106 0 1 1082
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_3
timestamp 1713338890
transform 1 0 6540 0 1 49
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_4
timestamp 1713338890
transform 1 0 1232 0 1 1480
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_5
timestamp 1713338890
transform 1 0 2701 0 1 1598
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_6
timestamp 1713338890
transform 1 0 1730 0 1 1480
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_7
timestamp 1713338890
transform 1 0 3044 0 1 1337
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_8
timestamp 1713338890
transform 1 0 3691 0 1 2228
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_9
timestamp 1713338890
transform 1 0 3966 0 1 1606
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_10
timestamp 1713338890
transform 1 0 4951 0 1 1338
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_11
timestamp 1713338890
transform 1 0 4439 0 1 1338
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_12
timestamp 1713338890
transform 1 0 6095 0 1 1338
box -90 -38 90 38
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_0
timestamp 1713338890
transform 1 0 6095 0 1 941
box -90 -90 90 90
use M2_M1_CDNS_69033583165538  M2_M1_CDNS_69033583165538_1
timestamp 1713338890
transform 1 0 6095 0 1 1727
box -90 -90 90 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_0
timestamp 1713338890
transform 0 -1 708 1 0 956
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_1
timestamp 1713338890
transform 0 -1 1182 1 0 311
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_2
timestamp 1713338890
transform 1 0 2183 0 1 664
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_3
timestamp 1713338890
transform 1 0 1695 0 1 664
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_4
timestamp 1713338890
transform 1 0 2672 0 1 664
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_5
timestamp 1713338890
transform 1 0 4515 0 1 778
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_6
timestamp 1713338890
transform 1 0 5779 0 1 941
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_7
timestamp 1713338890
transform 1 0 5391 0 1 778
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_8
timestamp 1713338890
transform 1 0 5003 0 1 779
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_9
timestamp 1713338890
transform 1 0 6411 0 1 941
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_10
timestamp 1713338890
transform 1 0 1861 0 1 1887
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_11
timestamp 1713338890
transform 1 0 3044 0 1 1820
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_12
timestamp 1713338890
transform 1 0 3265 0 1 2132
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_13
timestamp 1713338890
transform 1 0 4133 0 1 2028
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_14
timestamp 1713338890
transform 1 0 4375 0 1 1820
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_15
timestamp 1713338890
transform 1 0 4617 0 1 2028
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_16
timestamp 1713338890
transform 1 0 5779 0 1 1726
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_17
timestamp 1713338890
transform 1 0 5241 0 1 2028
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_18
timestamp 1713338890
transform 1 0 6411 0 1 1727
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_19
timestamp 1713338890
transform 1 0 6592 0 1 1703
box -38 -90 38 90
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_0
timestamp 1713338890
transform 1 0 6219 0 1 731
box -88 -44 228 344
use nmos_6p0_CDNS_4066195314535  nmos_6p0_CDNS_4066195314535_0
timestamp 1713338890
transform 1 0 459 0 1 280
box -88 -44 472 444
use nmos_6p0_CDNS_4066195314536  nmos_6p0_CDNS_4066195314536_0
timestamp 1713338890
transform -1 0 1310 0 -1 920
box -88 -44 228 344
use nmos_6p0_CDNS_4066195314536  nmos_6p0_CDNS_4066195314536_1
timestamp 1713338890
transform 1 0 5831 0 1 731
box -88 -44 228 344
use nmos_6p0_CDNS_4066195314537  nmos_6p0_CDNS_4066195314537_0
timestamp 1713338890
transform 1 0 1747 0 1 280
box -88 -44 1204 684
use nmos_6p0_CDNS_4066195314540  nmos_6p0_CDNS_4066195314540_0
timestamp 1713338890
transform 1 0 5443 0 1 608
box -88 -44 228 304
use nmos_6p0_CDNS_4066195314541  nmos_6p0_CDNS_4066195314541_0
timestamp 1713338890
transform 1 0 3203 0 1 338
box -88 -44 960 574
use nmos_6p0_CDNS_4066195314542  nmos_6p0_CDNS_4066195314542_0
timestamp 1713338890
transform 1 0 4323 0 1 268
box -88 -44 960 644
use pmos_6p0_CDNS_4066195314534  pmos_6p0_CDNS_4066195314534_0
timestamp 1713338890
transform -1 0 2053 0 1 1797
box -208 -120 592 420
use pmos_6p0_CDNS_4066195314538  pmos_6p0_CDNS_4066195314538_0
timestamp 1713338890
transform 1 0 4183 0 1 1730
box -208 -120 592 550
use pmos_6p0_CDNS_4066195314539  pmos_6p0_CDNS_4066195314539_0
timestamp 1713338890
transform -1 0 5971 0 -1 2037
box -208 -120 348 520
use pmos_6p0_CDNS_4066195314539  pmos_6p0_CDNS_4066195314539_1
timestamp 1713338890
transform 1 0 6219 0 -1 2037
box -208 -120 348 520
use pmos_6p0_CDNS_4066195314543  pmos_6p0_CDNS_4066195314543_0
timestamp 1713338890
transform -1 0 2993 0 -1 2197
box -208 -120 836 520
use pmos_6p0_CDNS_4066195314544  pmos_6p0_CDNS_4066195314544_0
timestamp 1713338890
transform 1 0 3315 0 1 1730
box -208 -120 592 500
use pmos_6p0_CDNS_4066195314544  pmos_6p0_CDNS_4066195314544_1
timestamp 1713338890
transform 1 0 4815 0 1 1730
box -208 -120 592 500
use pmos_6p0_CDNS_4066195314545  pmos_6p0_CDNS_4066195314545_0
timestamp 1713338890
transform -1 0 843 0 1 1335
box -208 -120 592 920
<< labels >>
rlabel metal1 s 6269 1344 6269 1344 4 Z
port 1 nsew
rlabel metal1 s 320 39 320 39 4 DVSS
port 2 nsew
rlabel metal1 s 4228 1072 4228 1072 4 A
port 3 nsew
rlabel metal1 s 884 2452 884 2452 4 DVDD
port 4 nsew
rlabel metal2 s 855 960 855 960 4 CS
port 5 nsew
rlabel metal2 s 2695 1339 2695 1339 4 IE
port 6 nsew
<< end >>
