magic
tech gf180mcuC
magscale 1 10
timestamp 1691396512
<< pwell >>
rect -540 -772 540 772
<< nmos >>
rect -428 454 -372 704
rect -268 454 -212 704
rect -108 454 -52 704
rect 52 454 108 704
rect 212 454 268 704
rect 372 454 428 704
rect -428 68 -372 318
rect -268 68 -212 318
rect -108 68 -52 318
rect 52 68 108 318
rect 212 68 268 318
rect 372 68 428 318
rect -428 -318 -372 -68
rect -268 -318 -212 -68
rect -108 -318 -52 -68
rect 52 -318 108 -68
rect 212 -318 268 -68
rect 372 -318 428 -68
rect -428 -704 -372 -454
rect -268 -704 -212 -454
rect -108 -704 -52 -454
rect 52 -704 108 -454
rect 212 -704 268 -454
rect 372 -704 428 -454
<< ndiff >>
rect -516 691 -428 704
rect -516 467 -503 691
rect -457 467 -428 691
rect -516 454 -428 467
rect -372 691 -268 704
rect -372 467 -343 691
rect -297 467 -268 691
rect -372 454 -268 467
rect -212 691 -108 704
rect -212 467 -183 691
rect -137 467 -108 691
rect -212 454 -108 467
rect -52 691 52 704
rect -52 467 -23 691
rect 23 467 52 691
rect -52 454 52 467
rect 108 691 212 704
rect 108 467 137 691
rect 183 467 212 691
rect 108 454 212 467
rect 268 691 372 704
rect 268 467 297 691
rect 343 467 372 691
rect 268 454 372 467
rect 428 691 516 704
rect 428 467 457 691
rect 503 467 516 691
rect 428 454 516 467
rect -516 305 -428 318
rect -516 81 -503 305
rect -457 81 -428 305
rect -516 68 -428 81
rect -372 305 -268 318
rect -372 81 -343 305
rect -297 81 -268 305
rect -372 68 -268 81
rect -212 305 -108 318
rect -212 81 -183 305
rect -137 81 -108 305
rect -212 68 -108 81
rect -52 305 52 318
rect -52 81 -23 305
rect 23 81 52 305
rect -52 68 52 81
rect 108 305 212 318
rect 108 81 137 305
rect 183 81 212 305
rect 108 68 212 81
rect 268 305 372 318
rect 268 81 297 305
rect 343 81 372 305
rect 268 68 372 81
rect 428 305 516 318
rect 428 81 457 305
rect 503 81 516 305
rect 428 68 516 81
rect -516 -81 -428 -68
rect -516 -305 -503 -81
rect -457 -305 -428 -81
rect -516 -318 -428 -305
rect -372 -81 -268 -68
rect -372 -305 -343 -81
rect -297 -305 -268 -81
rect -372 -318 -268 -305
rect -212 -81 -108 -68
rect -212 -305 -183 -81
rect -137 -305 -108 -81
rect -212 -318 -108 -305
rect -52 -81 52 -68
rect -52 -305 -23 -81
rect 23 -305 52 -81
rect -52 -318 52 -305
rect 108 -81 212 -68
rect 108 -305 137 -81
rect 183 -305 212 -81
rect 108 -318 212 -305
rect 268 -81 372 -68
rect 268 -305 297 -81
rect 343 -305 372 -81
rect 268 -318 372 -305
rect 428 -81 516 -68
rect 428 -305 457 -81
rect 503 -305 516 -81
rect 428 -318 516 -305
rect -516 -467 -428 -454
rect -516 -691 -503 -467
rect -457 -691 -428 -467
rect -516 -704 -428 -691
rect -372 -467 -268 -454
rect -372 -691 -343 -467
rect -297 -691 -268 -467
rect -372 -704 -268 -691
rect -212 -467 -108 -454
rect -212 -691 -183 -467
rect -137 -691 -108 -467
rect -212 -704 -108 -691
rect -52 -467 52 -454
rect -52 -691 -23 -467
rect 23 -691 52 -467
rect -52 -704 52 -691
rect 108 -467 212 -454
rect 108 -691 137 -467
rect 183 -691 212 -467
rect 108 -704 212 -691
rect 268 -467 372 -454
rect 268 -691 297 -467
rect 343 -691 372 -467
rect 268 -704 372 -691
rect 428 -467 516 -454
rect 428 -691 457 -467
rect 503 -691 516 -467
rect 428 -704 516 -691
<< ndiffc >>
rect -503 467 -457 691
rect -343 467 -297 691
rect -183 467 -137 691
rect -23 467 23 691
rect 137 467 183 691
rect 297 467 343 691
rect 457 467 503 691
rect -503 81 -457 305
rect -343 81 -297 305
rect -183 81 -137 305
rect -23 81 23 305
rect 137 81 183 305
rect 297 81 343 305
rect 457 81 503 305
rect -503 -305 -457 -81
rect -343 -305 -297 -81
rect -183 -305 -137 -81
rect -23 -305 23 -81
rect 137 -305 183 -81
rect 297 -305 343 -81
rect 457 -305 503 -81
rect -503 -691 -457 -467
rect -343 -691 -297 -467
rect -183 -691 -137 -467
rect -23 -691 23 -467
rect 137 -691 183 -467
rect 297 -691 343 -467
rect 457 -691 503 -467
<< polysilicon >>
rect -428 704 -372 748
rect -268 704 -212 748
rect -108 704 -52 748
rect 52 704 108 748
rect 212 704 268 748
rect 372 704 428 748
rect -428 410 -372 454
rect -268 410 -212 454
rect -108 410 -52 454
rect 52 410 108 454
rect 212 410 268 454
rect 372 410 428 454
rect -428 318 -372 362
rect -268 318 -212 362
rect -108 318 -52 362
rect 52 318 108 362
rect 212 318 268 362
rect 372 318 428 362
rect -428 24 -372 68
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect 372 24 428 68
rect -428 -68 -372 -24
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect 372 -68 428 -24
rect -428 -362 -372 -318
rect -268 -362 -212 -318
rect -108 -362 -52 -318
rect 52 -362 108 -318
rect 212 -362 268 -318
rect 372 -362 428 -318
rect -428 -454 -372 -410
rect -268 -454 -212 -410
rect -108 -454 -52 -410
rect 52 -454 108 -410
rect 212 -454 268 -410
rect 372 -454 428 -410
rect -428 -748 -372 -704
rect -268 -748 -212 -704
rect -108 -748 -52 -704
rect 52 -748 108 -704
rect 212 -748 268 -704
rect 372 -748 428 -704
<< metal1 >>
rect -503 691 -457 702
rect -503 456 -457 467
rect -343 691 -297 702
rect -343 456 -297 467
rect -183 691 -137 702
rect -183 456 -137 467
rect -23 691 23 702
rect -23 456 23 467
rect 137 691 183 702
rect 137 456 183 467
rect 297 691 343 702
rect 297 456 343 467
rect 457 691 503 702
rect 457 456 503 467
rect -503 305 -457 316
rect -503 70 -457 81
rect -343 305 -297 316
rect -343 70 -297 81
rect -183 305 -137 316
rect -183 70 -137 81
rect -23 305 23 316
rect -23 70 23 81
rect 137 305 183 316
rect 137 70 183 81
rect 297 305 343 316
rect 297 70 343 81
rect 457 305 503 316
rect 457 70 503 81
rect -503 -81 -457 -70
rect -503 -316 -457 -305
rect -343 -81 -297 -70
rect -343 -316 -297 -305
rect -183 -81 -137 -70
rect -183 -316 -137 -305
rect -23 -81 23 -70
rect -23 -316 23 -305
rect 137 -81 183 -70
rect 137 -316 183 -305
rect 297 -81 343 -70
rect 297 -316 343 -305
rect 457 -81 503 -70
rect 457 -316 503 -305
rect -503 -467 -457 -456
rect -503 -702 -457 -691
rect -343 -467 -297 -456
rect -343 -702 -297 -691
rect -183 -467 -137 -456
rect -183 -702 -137 -691
rect -23 -467 23 -456
rect -23 -702 23 -691
rect 137 -467 183 -456
rect 137 -702 183 -691
rect 297 -467 343 -456
rect 297 -702 343 -691
rect 457 -467 503 -456
rect 457 -702 503 -691
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1.25 l 0.280 m 4 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
