* NGSPICE file created from DFF__flat.ext - technology: gf180mcuC

.subckt DFF__flat Q QB CLK RST D VSS VDD
X0 VDD nand2_2.IN1 nand2_3.IN2 VDD.t36 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1 a_3096_435# nand2_2.IN2 VSS.t16 VSS.t15 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2 a_2200_553# inv_0.OUT VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3 nand2_3.OUT nand2_3.IN2 VDD.t24 VDD.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 VDD nand2_5.OUT nand2_2.IN1 VDD.t15 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X5 nand2_2.IN1 nand2_5.OUT a_81_2165# VSS.t9 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X6 VDD QB.t3 Q.t1 VDD.t39 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X7 nand2_3.IN2 nand2_2.IN1 a_247_494# VSS.t23 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X8 VDD nand2_3.OUT nand2_5.OUT VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X9 VDD nand2_5.IN2 nand2_2.IN2 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X10 inv_0.OUT nand2_3.OUT VSS.t22 VSS.t21 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X11 nand2_5.OUT nand2_3.OUT a_2196_1932# VSS.t20 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X12 a_964_487# nand2_3.IN2 VSS.t12 VSS.t11 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X13 VDD RST.t0 nand2_3.OUT VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X14 Q QB.t4 a_3096_435# VSS.t10 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X15 VSS Q.t3 a_3092_1932# VSS.t24 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 VDD RST.t1 nand2_5.IN2 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X17 VDD Q.t4 QB.t2 VDD.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X18 a_3092_1932# nand2_5.OUT QB.t0 VSS.t8 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X19 QB nand2_5.OUT VDD.t14 VDD.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 nand2_2.IN2 nand2_5.IN2 a_2200_553# VSS.t7 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X21 nand2_5.IN2 RST.t2 a_967_2122# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X22 nand2_5.IN2 CLK.t0 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 nand2_3.OUT RST.t3 a_964_487# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X24 a_967_2122# CLK.t1 VSS.t4 VSS.t3 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X25 a_2196_1932# nand2_5.IN2 VSS.t6 VSS.t5 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X26 nand2_5.OUT nand2_5.IN2 VDD.t9 VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X27 nand2_3.IN2 nand2_2.IN2 VDD.t28 VDD.t27 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X28 Q nand2_2.IN2 VDD.t26 VDD.t25 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X29 nand2_2.IN1 D.t0 VDD.t4 VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X30 nand2_2.IN2 inv_0.OUT VDD.t30 VDD.t29 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 a_247_494# nand2_2.IN2 VSS.t14 VSS.t13 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X32 a_81_2165# D.t1 VSS.t2 VSS.t1 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X33 inv_0.OUT nand2_3.OUT VDD.t32 VDD.t31 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 VDD.t29 VDD.n26 354.539
R1 VDD.n26 VDD 285.887
R2 VDD.n26 VDD.t31 280.245
R3 VDD.n13 VDD.t39 232.809
R4 VDD.n16 VDD.t13 232.803
R5 VDD.n24 VDD.t33 230.548
R6 VDD.n24 VDD.t8 230.548
R7 VDD.n15 VDD.t18 227.667
R8 VDD.n14 VDD.t25 227.667
R9 VDD.n1 VDD.t36 193.183
R10 VDD.n46 VDD.t15 193.183
R11 VDD.n39 VDD.t5 193.183
R12 VDD.n35 VDD.t0 193.183
R13 VDD.n24 VDD.t10 143.345
R14 VDD.n1 VDD.t27 109.849
R15 VDD.n46 VDD.t3 109.849
R16 VDD.n39 VDD.t23 109.849
R17 VDD.n35 VDD.t21 109.849
R18 VDD.n27 VDD.t29 92.1507
R19 VDD.n17 VDD.n16 59.3792
R20 VDD.n13 VDD.n12 56.5869
R21 VDD.n25 VDD.n24 30.7172
R22 VDD.n42 VDD.n41 8.95925
R23 VDD.n27 VDD.n25 6.82644
R24 VDD.n2 VDD.t28 6.45146
R25 VDD.n47 VDD.n46 6.3005
R26 VDD.n36 VDD.n35 6.3005
R27 VDD.n40 VDD.n39 6.3005
R28 VDD.n51 VDD.n1 6.3005
R29 VDD.n15 VDD.n14 5.60274
R30 VDD.n38 VDD.n37 5.43849
R31 VDD.n33 VDD.t32 5.26145
R32 VDD.n47 VDD.t4 5.21701
R33 VDD.n45 VDD.n3 5.1806
R34 VDD.n31 VDD.t9 5.13746
R35 VDD.n5 VDD.t22 5.13746
R36 VDD.n41 VDD.t24 5.13746
R37 VDD.n11 VDD.n9 5.13586
R38 VDD.n18 VDD.t26 5.13586
R39 VDD.n11 VDD.n10 5.13334
R40 VDD.n21 VDD.n7 5.13287
R41 VDD.n34 VDD.n6 5.13287
R42 VDD.n43 VDD.n4 5.13287
R43 VDD.n19 VDD.t14 5.13129
R44 VDD.n30 VDD.t30 5.10854
R45 VDD.n20 VDD.n8 5.10445
R46 VDD.n20 VDD.n19 4.88931
R47 VDD.n44 VDD.n43 4.69819
R48 VDD.n34 VDD.n33 4.3827
R49 VDD.n42 VDD.n5 4.34898
R50 VDD.n29 VDD.n28 3.1505
R51 VDD.n28 VDD.n27 3.1505
R52 VDD.n23 VDD.n22 3.1505
R53 VDD.n25 VDD.n23 3.1505
R54 VDD.n45 VDD.n44 0.783866
R55 VDD.n50 VDD.n2 0.7205
R56 VDD.n41 VDD.n40 0.257375
R57 VDD.n49 VDD 0.256289
R58 VDD.n43 VDD.n42 0.238698
R59 VDD.n49 VDD.n48 0.147138
R60 VDD.n50 VDD.n49 0.143395
R61 VDD.n28 VDD.n23 0.138205
R62 VDD.n32 VDD.n31 0.134086
R63 VDD.n16 VDD.n15 0.117546
R64 VDD.n14 VDD.n13 0.111412
R65 VDD VDD.n0 0.1055
R66 VDD VDD.n21 0.0786463
R67 VDD.n30 VDD.n29 0.0588902
R68 VDD.n48 VDD 0.0585645
R69 VDD.n51 VDD.n50 0.0573421
R70 VDD.n12 VDD.n11 0.040956
R71 VDD.n18 VDD.n17 0.0406629
R72 VDD.n38 VDD.n34 0.0383228
R73 VDD VDD.n38 0.036125
R74 VDD.n36 VDD.n5 0.0317152
R75 VDD.n32 VDD 0.00853834
R76 VDD.n40 VDD 0.00425
R77 VDD.n38 VDD 0.00414557
R78 VDD.n19 VDD.n18 0.00284528
R79 VDD.n21 VDD.n20 0.0022561
R80 VDD.n31 VDD.n30 0.0022561
R81 VDD.n33 VDD.n32 0.00213514
R82 VDD VDD.n51 0.00207895
R83 VDD VDD.n47 0.00166129
R84 VDD.n22 VDD 0.00137805
R85 VDD.n22 VDD 0.00137805
R86 VDD.n29 VDD 0.00137805
R87 VDD.n17 VDD 0.00108632
R88 VDD.n48 VDD.n45 0.00102847
R89 VDD VDD.n36 0.000955696
R90 VDD.n12 VDD 0.00079316
R91 VSS.n20 VSS.n16 12464.5
R92 VSS.t24 VSS.t10 12443.8
R93 VSS.n13 VSS.n12 9145.5
R94 VSS.t13 VSS.n21 7295.5
R95 VSS.n18 VSS.n17 5903.67
R96 VSS.n8 VSS.n5 5863.4
R97 VSS.n13 VSS.t15 1981.2
R98 VSS.t19 VSS.n18 1806.74
R99 VSS.n8 VSS.t9 1797.09
R100 VSS.t7 VSS.n13 1774.48
R101 VSS.t3 VSS.n8 1504.67
R102 VSS.n20 VSS.t11 1486.68
R103 VSS.n10 VSS.t0 1474.19
R104 VSS.t23 VSS.n20 1469.11
R105 VSS.n12 VSS.t8 1422.12
R106 VSS.n12 VSS.t20 1422.12
R107 VSS.n15 VSS.t21 1013.61
R108 VSS.n15 VSS.t17 954.749
R109 VSS.t5 VSS.n10 788.294
R110 VSS.n18 VSS.n15 726.975
R111 VSS.n27 VSS.n15 600.497
R112 VSS.t10 VSS.n0 561.152
R113 VSS.t9 VSS.n7 513.159
R114 VSS.n19 VSS.t19 513.159
R115 VSS.n22 VSS.t23 507.317
R116 VSS.t0 VSS.n9 479.264
R117 VSS.n14 VSS.t7 462.909
R118 VSS.t15 VSS.n0 374.101
R119 VSS.t20 VSS.n11 370.988
R120 VSS.n7 VSS.t1 342.106
R121 VSS.t11 VSS.n19 342.106
R122 VSS.n22 VSS.t13 338.212
R123 VSS.n9 VSS.t3 319.509
R124 VSS.t17 VSS.n14 308.606
R125 VSS.n3 VSS.t24 247.326
R126 VSS.n11 VSS.t5 247.326
R127 VSS.n23 VSS.t14 13.7049
R128 VSS.n25 VSS.t22 9.38224
R129 VSS.n25 VSS.n24 8.91518
R130 VSS VSS.t2 7.20679
R131 VSS.n6 VSS.t4 7.19156
R132 VSS.n28 VSS.t18 7.19156
R133 VSS.n4 VSS.t6 7.18989
R134 VSS.n2 VSS.n1 7.18989
R135 VSS.n24 VSS.t12 7.12323
R136 VSS.n29 VSS.t16 7.03656
R137 VSS.n2 VSS 6.54995
R138 VSS.n7 VSS 5.2005
R139 VSS.n9 VSS 5.2005
R140 VSS VSS.n3 5.2005
R141 VSS.n11 VSS 5.2005
R142 VSS.n19 VSS 5.2005
R143 VSS VSS.n22 5.2005
R144 VSS VSS.n14 5.2005
R145 VSS VSS.n0 5.2005
R146 VSS.n24 VSS.n23 1.49675
R147 VSS VSS.n4 0.840934
R148 VSS VSS.n6 0.545498
R149 VSS.n26 VSS 0.283187
R150 VSS.n29 VSS 0.278241
R151 VSS.n23 VSS 0.175346
R152 VSS.n6 VSS 0.118573
R153 VSS.n28 VSS 0.114176
R154 VSS.n23 VSS 0.109927
R155 VSS VSS.n2 0.0874595
R156 VSS.n4 VSS 0.0874595
R157 VSS.n26 VSS.n25 0.0832857
R158 VSS VSS.n29 0.055266
R159 VSS VSS.n28 0.05
R160 VSS.n27 VSS.n26 0.0173321
R161 VSS VSS.n27 0.000843511
R162 QB.n4 QB.t4 31.528
R163 QB.n4 QB.t3 15.3826
R164 QB QB.n4 8.85715
R165 QB QB.t0 7.15141
R166 QB.n3 QB.n2 6.61429
R167 QB.n2 QB.n1 3.21115
R168 QB.n1 QB.t2 2.2755
R169 QB.n1 QB.n0 2.2755
R170 QB.n3 QB 0.667669
R171 QB QB.n3 0.0203305
R172 QB.n2 QB 0.0135909
R173 Q.n5 Q.t4 30.9379
R174 Q.n5 Q.t3 21.6422
R175 Q.n3 Q.n2 7.12686
R176 Q.n4 Q.n3 6.83791
R177 Q Q.n5 4.00612
R178 Q Q.n1 3.22776
R179 Q.n1 Q.t1 2.2755
R180 Q.n1 Q.n0 2.2755
R181 Q.n4 Q 0.539612
R182 Q Q.n4 0.385684
R183 Q.n3 Q 0.0250455
R184 RST.n0 RST.t2 31.528
R185 RST.n2 RST.t3 31.528
R186 RST.n0 RST.t1 15.3826
R187 RST.n2 RST.t0 15.3826
R188 RST RST.n0 8.85806
R189 RST RST.n2 8.85806
R190 RST.n1 RST 4.66096
R191 RST RST.n1 3.58511
R192 RST.n1 RST 2.45348
R193 CLK.n0 CLK.t0 30.9379
R194 CLK.n0 CLK.t1 21.6422
R195 CLK CLK.n0 4.005
R196 CLK CLK.n1 2.25153
R197 D.n0 D.t0 30.9379
R198 D.n0 D.t1 21.6422
R199 D D.n0 4.005
C0 nand2_2.IN2 nand2_5.OUT 0.0065f
C1 nand2_5.IN2 Q 0.0118f
C2 nand2_5.IN2 RST 0.487f
C3 nand2_5.IN2 a_3096_435# 1.63e-20
C4 nand2_5.IN2 nand2_2.IN1 0.00714f
C5 nand2_2.IN2 CLK 0.0318f
C6 nand2_5.IN2 a_2196_1932# 0.00376f
C7 a_81_2165# RST 8.75e-20
C8 a_81_2165# nand2_2.IN1 0.069f
C9 nand2_5.OUT VDD 0.742f
C10 nand2_5.OUT D 0.0475f
C11 Q a_2200_553# 1.06e-19
C12 nand2_5.OUT inv_0.OUT 1.02e-21
C13 VDD CLK 0.611f
C14 CLK D 0.0266f
C15 nand2_5.OUT a_967_2122# 3.83e-19
C16 nand2_2.IN2 nand2_3.OUT 0.0984f
C17 nand2_5.IN2 nand2_5.OUT 0.176f
C18 a_967_2122# CLK 0.00347f
C19 nand2_5.IN2 CLK 0.114f
C20 nand2_2.IN2 a_247_494# 0.0175f
C21 a_81_2165# nand2_5.OUT 0.00432f
C22 nand2_3.OUT VDD 0.886f
C23 VDD a_3092_1932# 3.15e-19
C24 nand2_2.IN2 QB 0.147f
C25 inv_0.OUT nand2_3.OUT 0.142f
C26 a_81_2165# CLK 9.59e-19
C27 a_247_494# VDD 3.14e-19
C28 QB VDD 1.07f
C29 nand2_5.IN2 nand2_3.OUT 0.39f
C30 QB inv_0.OUT 0.00316f
C31 nand2_2.IN2 nand2_3.IN2 0.159f
C32 nand2_3.OUT a_2200_553# 2.09e-19
C33 nand2_5.IN2 QB 0.273f
C34 a_964_487# RST 0.00348f
C35 a_3096_435# Q 0.069f
C36 a_964_487# nand2_2.IN1 9.39e-21
C37 nand2_3.IN2 VDD 0.39f
C38 nand2_2.IN1 RST 0.0963f
C39 RST a_2196_1932# 0.00168f
C40 nand2_5.OUT RST 0.355f
C41 nand2_5.OUT Q 0.0652f
C42 nand2_2.IN1 nand2_5.OUT 0.492f
C43 nand2_5.OUT a_2196_1932# 0.0703f
C44 RST CLK 0.0528f
C45 nand2_2.IN1 CLK 0.145f
C46 a_964_487# nand2_3.OUT 0.069f
C47 nand2_3.OUT Q 2.23e-19
C48 nand2_3.OUT RST 0.889f
C49 Q a_3092_1932# 0.00347f
C50 a_3096_435# nand2_3.OUT 9.07e-21
C51 nand2_2.IN1 nand2_3.OUT 0.0185f
C52 nand2_2.IN2 VDD 0.71f
C53 nand2_2.IN2 D 9.66e-20
C54 nand2_3.OUT a_2196_1932# 0.00594f
C55 nand2_2.IN2 inv_0.OUT 0.155f
C56 nand2_5.OUT CLK 0.115f
C57 nand2_2.IN1 a_247_494# 0.00348f
C58 QB Q 0.631f
C59 VDD D 0.183f
C60 nand2_2.IN2 a_967_2122# 2.82e-20
C61 a_3096_435# QB 0.00619f
C62 inv_0.OUT VDD 0.346f
C63 nand2_5.IN2 nand2_2.IN2 0.459f
C64 VDD a_967_2122# 3.14e-19
C65 nand2_5.OUT nand2_3.OUT 0.42f
C66 a_81_2165# nand2_2.IN2 1.16e-20
C67 nand2_5.OUT a_3092_1932# 0.00454f
C68 nand2_5.IN2 VDD 1.3f
C69 nand2_2.IN2 a_2200_553# 0.0769f
C70 nand2_5.IN2 inv_0.OUT 0.0551f
C71 a_964_487# nand2_3.IN2 0.00364f
C72 nand2_3.IN2 RST 0.0494f
C73 nand2_5.OUT a_247_494# 1.99e-20
C74 nand2_2.IN1 nand2_3.IN2 0.451f
C75 a_81_2165# VDD 3.14e-19
C76 a_81_2165# D 0.00347f
C77 nand2_5.OUT QB 0.581f
C78 a_247_494# CLK 1.27e-19
C79 VDD a_2200_553# 3.22e-19
C80 nand2_5.IN2 a_967_2122# 0.069f
C81 inv_0.OUT a_2200_553# 0.00372f
C82 nand2_5.IN2 a_2200_553# 0.00384f
C83 a_247_494# nand2_3.OUT 1.26e-20
C84 nand2_3.IN2 nand2_5.OUT 1.33e-19
C85 QB nand2_3.OUT 0.0138f
C86 QB a_3092_1932# 0.0692f
C87 nand2_3.IN2 CLK 0.00375f
C88 nand2_3.IN2 nand2_3.OUT 0.106f
C89 a_964_487# nand2_2.IN2 0.0144f
C90 nand2_2.IN2 RST 0.0259f
C91 nand2_2.IN2 Q 0.117f
C92 nand2_2.IN2 a_3096_435# 0.00411f
C93 nand2_2.IN1 nand2_2.IN2 0.0753f
C94 nand2_3.IN2 a_247_494# 0.069f
C95 a_964_487# VDD 3.14e-19
C96 VDD RST 0.727f
C97 VDD Q 0.507f
C98 RST D 1.99e-19
C99 a_3096_435# VDD 3.15e-19
C100 nand2_2.IN1 VDD 0.769f
C101 nand2_2.IN1 D 0.0995f
C102 VDD a_2196_1932# 3.14e-19
C103 a_964_487# inv_0.OUT 1.29e-20
C104 inv_0.OUT Q 5.29e-19
C105 inv_0.OUT RST 0.00685f
C106 nand2_2.IN1 inv_0.OUT 4.23e-20
C107 RST a_967_2122# 0.00519f
.ends

