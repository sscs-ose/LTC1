magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2109 -2251 2109 2251
<< metal2 >>
rect -109 241 109 251
rect -109 185 -99 241
rect -43 185 43 241
rect 99 185 109 241
rect -109 99 109 185
rect -109 43 -99 99
rect -43 43 43 99
rect 99 43 109 99
rect -109 -43 109 43
rect -109 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 109 -43
rect -109 -185 109 -99
rect -109 -241 -99 -185
rect -43 -241 43 -185
rect 99 -241 109 -185
rect -109 -251 109 -241
<< via2 >>
rect -99 185 -43 241
rect 43 185 99 241
rect -99 43 -43 99
rect 43 43 99 99
rect -99 -99 -43 -43
rect 43 -99 99 -43
rect -99 -241 -43 -185
rect 43 -241 99 -185
<< metal3 >>
rect -109 241 109 251
rect -109 185 -99 241
rect -43 185 43 241
rect 99 185 109 241
rect -109 99 109 185
rect -109 43 -99 99
rect -43 43 43 99
rect 99 43 109 99
rect -109 -43 109 43
rect -109 -99 -99 -43
rect -43 -99 43 -43
rect 99 -99 109 -43
rect -109 -185 109 -99
rect -109 -241 -99 -185
rect -43 -241 43 -185
rect 99 -241 109 -185
rect -109 -251 109 -241
<< end >>
