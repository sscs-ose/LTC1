magic
tech gf180mcuC
magscale 1 10
timestamp 1699938486
<< polysilicon >>
rect 1922 -2219 2195 -2192
rect 1922 -2269 1940 -2219
rect 1990 -2269 2195 -2219
rect 1922 -2292 2195 -2269
rect 4930 -2224 5203 -2197
rect 4930 -2274 4948 -2224
rect 4998 -2274 5203 -2224
rect 4930 -2297 5203 -2274
rect 7940 -2221 8213 -2194
rect 7940 -2271 7958 -2221
rect 8008 -2271 8213 -2221
rect 7940 -2294 8213 -2271
rect 10930 -2222 11203 -2195
rect 10930 -2272 10947 -2222
rect 10998 -2272 11203 -2222
rect 10930 -2295 11203 -2272
rect 13938 -2220 14211 -2193
rect 13938 -2270 13956 -2220
rect 14006 -2270 14211 -2220
rect 13938 -2293 14211 -2270
rect 16931 -2220 17204 -2193
rect 16931 -2270 16949 -2220
rect 16999 -2270 17204 -2220
rect 16931 -2293 17204 -2270
rect 29360 -2224 29633 -2197
rect 29360 -2274 29565 -2224
rect 29615 -2274 29633 -2224
rect 29360 -2297 29633 -2274
rect 32355 -2220 32628 -2193
rect 32355 -2270 32560 -2220
rect 32610 -2270 32628 -2220
rect 32355 -2293 32628 -2270
rect 35368 -2221 35641 -2194
rect 35368 -2271 35573 -2221
rect 35623 -2271 35641 -2221
rect 35368 -2294 35641 -2271
rect 38367 -2221 38640 -2194
rect 38367 -2271 38572 -2221
rect 38622 -2271 38640 -2221
rect 38367 -2294 38640 -2271
rect 41368 -2219 41641 -2192
rect 41368 -2269 41573 -2219
rect 41623 -2269 41641 -2219
rect 41368 -2292 41641 -2269
rect 44364 -2221 44637 -2194
rect 44364 -2271 44569 -2221
rect 44619 -2271 44637 -2221
rect 44364 -2294 44637 -2271
<< polycontact >>
rect 1940 -2269 1990 -2219
rect 4948 -2274 4998 -2224
rect 7958 -2271 8008 -2221
rect 10947 -2272 10998 -2222
rect 13956 -2270 14006 -2220
rect 16949 -2270 16999 -2220
rect 29565 -2274 29615 -2224
rect 32560 -2270 32610 -2220
rect 35573 -2271 35623 -2221
rect 38572 -2271 38622 -2221
rect 41573 -2269 41623 -2219
rect 44569 -2271 44619 -2221
<< metal1 >>
rect 1738 13337 2033 13381
rect 1738 13266 1770 13337
rect 1841 13334 2033 13337
rect 1841 13266 1913 13334
rect 1738 13263 1913 13266
rect 1984 13263 2033 13334
rect 1738 13205 2033 13263
rect 1738 13134 1770 13205
rect 1841 13134 1913 13205
rect 1984 13200 2033 13205
rect 1984 13134 2550 13200
rect 1738 13078 2550 13134
rect 1738 13007 1769 13078
rect 1840 13075 2550 13078
rect 1840 13007 1912 13075
rect 1738 13004 1912 13007
rect 1983 13040 2550 13075
rect 1983 13004 2033 13040
rect 1738 12946 2033 13004
rect 1738 12875 1769 12946
rect 1840 12875 1912 12946
rect 1983 12875 2033 12946
rect 1738 12857 2033 12875
rect 12903 12757 13223 14621
rect 15108 12757 15428 14642
rect 16747 12757 17067 14611
rect -428 7425 367 7585
rect 2564 6437 3090 7297
rect 4709 6437 5783 6736
rect -191 5911 5783 6437
rect -191 4272 335 5911
rect -191 3746 974 4272
rect -191 2853 335 3746
rect -191 2327 990 2853
rect -191 194 335 2327
rect 1021 194 1547 1498
rect 14192 1331 14476 1437
rect 16027 1331 16311 1408
rect 17235 1331 17519 1370
rect 14192 712 17542 1331
rect -191 -332 1547 194
rect -191 -3864 335 -332
rect 1021 -1330 1547 -332
rect 16923 177 17542 712
rect 16923 -442 19764 177
rect 1021 -1671 17438 -1330
rect 1021 -3864 1547 -1671
rect 19145 -1779 19764 -442
rect 20208 -191 20797 1200
rect 25804 31 26393 1101
rect 28356 31 28945 1200
rect 20208 -780 21909 -191
rect 21320 -1330 21909 -780
rect 25804 -558 28945 31
rect 25804 -1330 26393 -558
rect 21173 -1671 44832 -1330
rect 19145 -1829 19775 -1779
rect 19145 -1832 19518 -1829
rect 19145 -1900 19204 -1832
rect 19272 -1900 19324 -1832
rect 19392 -1897 19518 -1832
rect 19586 -1897 19638 -1829
rect 19706 -1897 19775 -1829
rect 19392 -1900 19775 -1897
rect 3504 -1952 3719 -1938
rect 3504 -2020 3518 -1952
rect 3586 -2020 3638 -1952
rect 3706 -2020 3719 -1952
rect 1733 -2094 1830 -2071
rect 1733 -2158 1748 -2094
rect 1813 -2158 1830 -2094
rect 3504 -2072 3719 -2020
rect 6504 -1952 6719 -1938
rect 6504 -2020 6518 -1952
rect 6586 -2020 6638 -1952
rect 6706 -2020 6719 -1952
rect 3504 -2107 3518 -2072
rect 3342 -2140 3518 -2107
rect 3586 -2140 3638 -2072
rect 3706 -2140 3719 -2072
rect 3342 -2153 3719 -2140
rect 4734 -2094 4831 -2071
rect 1733 -2192 1830 -2158
rect 4734 -2158 4749 -2094
rect 4814 -2158 4831 -2094
rect 6504 -2072 6719 -2020
rect 6504 -2107 6518 -2072
rect 6342 -2140 6518 -2107
rect 6586 -2140 6638 -2072
rect 6706 -2140 6719 -2072
rect 9504 -1952 9719 -1938
rect 9504 -2020 9518 -1952
rect 9586 -2020 9638 -1952
rect 9706 -2020 9719 -1952
rect 9504 -2072 9719 -2020
rect 12504 -1952 12719 -1938
rect 12504 -2020 12518 -1952
rect 12586 -2020 12638 -1952
rect 12706 -2020 12719 -1952
rect 6342 -2153 6719 -2140
rect 7750 -2097 7847 -2074
rect 4734 -2192 4831 -2158
rect 7750 -2161 7765 -2097
rect 7830 -2161 7847 -2097
rect 9504 -2107 9518 -2072
rect 9342 -2140 9518 -2107
rect 9586 -2140 9638 -2072
rect 9706 -2140 9719 -2072
rect 9342 -2153 9719 -2140
rect 10747 -2094 10844 -2071
rect 1733 -2214 2195 -2192
rect 1733 -2278 1748 -2214
rect 1813 -2278 1868 -2214
rect 1933 -2219 2195 -2214
rect 1933 -2269 1940 -2219
rect 1990 -2269 2195 -2219
rect 4734 -2197 4938 -2192
rect 7750 -2195 7847 -2161
rect 10747 -2158 10762 -2094
rect 10827 -2158 10844 -2094
rect 12504 -2072 12719 -2020
rect 15504 -1952 15719 -1938
rect 15504 -2020 15518 -1952
rect 15586 -2020 15638 -1952
rect 15706 -2020 15719 -1952
rect 12504 -2107 12518 -2072
rect 12342 -2140 12518 -2107
rect 12586 -2140 12638 -2072
rect 12706 -2140 12719 -2072
rect 12342 -2153 12719 -2140
rect 13776 -2092 13873 -2069
rect 10747 -2192 10844 -2158
rect 13776 -2156 13791 -2092
rect 13856 -2156 13873 -2092
rect 15504 -2072 15719 -2020
rect 18504 -1952 18719 -1938
rect 18504 -2020 18518 -1952
rect 18586 -2020 18638 -1952
rect 18706 -2020 18719 -1952
rect 15504 -2107 15518 -2072
rect 15342 -2140 15518 -2107
rect 15586 -2140 15638 -2072
rect 15706 -2140 15719 -2072
rect 15342 -2153 15719 -2140
rect 16807 -2094 16904 -2071
rect 13776 -2190 13873 -2156
rect 16807 -2158 16822 -2094
rect 16887 -2158 16904 -2094
rect 18504 -2072 18719 -2020
rect 18504 -2107 18518 -2072
rect 18342 -2140 18518 -2107
rect 18586 -2140 18638 -2072
rect 18706 -2140 18719 -2072
rect 18342 -2153 18719 -2140
rect 19145 -1949 19775 -1900
rect 19145 -1952 19518 -1949
rect 19145 -2020 19204 -1952
rect 19272 -2020 19324 -1952
rect 19392 -2017 19518 -1952
rect 19586 -2017 19638 -1949
rect 19706 -2017 19775 -1949
rect 19392 -2020 19775 -2017
rect 19145 -2075 19775 -2020
rect 19145 -2078 19520 -2075
rect 19145 -2146 19206 -2078
rect 19274 -2146 19326 -2078
rect 19394 -2143 19520 -2078
rect 19588 -2143 19640 -2075
rect 19708 -2143 19775 -2075
rect 19394 -2146 19775 -2143
rect 7940 -2195 8213 -2194
rect 4734 -2214 5203 -2197
rect 1933 -2278 2195 -2269
rect 1733 -2292 2195 -2278
rect 1733 -2297 1937 -2292
rect 3543 -2296 3734 -2250
rect 3598 -2318 3734 -2296
rect 4734 -2278 4749 -2214
rect 4814 -2278 4869 -2214
rect 4934 -2224 5203 -2214
rect 4934 -2274 4948 -2224
rect 4998 -2274 5203 -2224
rect 7750 -2217 8213 -2195
rect 4934 -2278 5203 -2274
rect 4734 -2297 5203 -2278
rect 6543 -2296 6734 -2250
rect 6598 -2318 6734 -2296
rect 7750 -2281 7765 -2217
rect 7830 -2281 7885 -2217
rect 7950 -2221 8213 -2217
rect 7950 -2271 7958 -2221
rect 8008 -2271 8213 -2221
rect 10747 -2195 10974 -2192
rect 13776 -2193 14003 -2190
rect 16807 -2192 16904 -2158
rect 16807 -2193 17034 -2192
rect 10747 -2214 11203 -2195
rect 7950 -2281 8213 -2271
rect 7750 -2294 8213 -2281
rect 7750 -2300 7977 -2294
rect 9543 -2296 9734 -2250
rect 9598 -2318 9734 -2296
rect 10747 -2278 10762 -2214
rect 10827 -2278 10882 -2214
rect 10947 -2222 11203 -2214
rect 10998 -2272 11203 -2222
rect 13776 -2212 14211 -2193
rect 10947 -2278 11203 -2272
rect 10747 -2295 11203 -2278
rect 10747 -2297 10974 -2295
rect 12543 -2296 12734 -2250
rect 13776 -2276 13791 -2212
rect 13856 -2276 13911 -2212
rect 13976 -2220 14211 -2212
rect 14006 -2270 14211 -2220
rect 16807 -2214 17204 -2193
rect 13976 -2276 14211 -2270
rect 13776 -2293 14211 -2276
rect 13776 -2295 14003 -2293
rect 15543 -2296 15734 -2250
rect 12598 -2318 12734 -2296
rect 15598 -2318 15734 -2296
rect 16807 -2278 16822 -2214
rect 16887 -2278 16942 -2214
rect 17007 -2278 17204 -2214
rect 19145 -2195 19775 -2146
rect 19145 -2198 19520 -2195
rect 16807 -2293 17204 -2278
rect 16807 -2297 17034 -2293
rect 18543 -2296 18734 -2250
rect 18598 -2318 18734 -2296
rect 19145 -2266 19206 -2198
rect 19274 -2266 19326 -2198
rect 19394 -2263 19520 -2198
rect 19588 -2263 19640 -2195
rect 19708 -2263 19775 -2195
rect 19394 -2266 19775 -2263
rect 3598 -2332 3864 -2318
rect 3598 -2400 3663 -2332
rect 3731 -2400 3783 -2332
rect 3851 -2400 3864 -2332
rect 3598 -2452 3864 -2400
rect 3598 -2479 3663 -2452
rect 3428 -2520 3663 -2479
rect 3731 -2520 3783 -2452
rect 3851 -2520 3864 -2452
rect 6598 -2332 6864 -2318
rect 6598 -2400 6663 -2332
rect 6731 -2400 6783 -2332
rect 6851 -2400 6864 -2332
rect 6598 -2452 6864 -2400
rect 6598 -2479 6663 -2452
rect 3428 -2525 3864 -2520
rect 6428 -2520 6663 -2479
rect 6731 -2520 6783 -2452
rect 6851 -2520 6864 -2452
rect 9598 -2332 9864 -2318
rect 9598 -2400 9663 -2332
rect 9731 -2400 9783 -2332
rect 9851 -2400 9864 -2332
rect 9598 -2452 9864 -2400
rect 9598 -2479 9663 -2452
rect 6428 -2525 6864 -2520
rect 9428 -2520 9663 -2479
rect 9731 -2520 9783 -2452
rect 9851 -2520 9864 -2452
rect 12598 -2332 12864 -2318
rect 12598 -2400 12663 -2332
rect 12731 -2400 12783 -2332
rect 12851 -2400 12864 -2332
rect 12598 -2452 12864 -2400
rect 12598 -2479 12663 -2452
rect 9428 -2525 9864 -2520
rect 12428 -2520 12663 -2479
rect 12731 -2520 12783 -2452
rect 12851 -2520 12864 -2452
rect 15598 -2332 15864 -2318
rect 15598 -2400 15663 -2332
rect 15731 -2400 15783 -2332
rect 15851 -2400 15864 -2332
rect 15598 -2452 15864 -2400
rect 15598 -2479 15663 -2452
rect 12428 -2525 12864 -2520
rect 15428 -2520 15663 -2479
rect 15731 -2520 15783 -2452
rect 15851 -2520 15864 -2452
rect 18598 -2332 18864 -2318
rect 18598 -2400 18663 -2332
rect 18731 -2400 18783 -2332
rect 18851 -2400 18864 -2332
rect 18598 -2452 18864 -2400
rect 18598 -2479 18663 -2452
rect 15428 -2525 15864 -2520
rect 18428 -2520 18663 -2479
rect 18731 -2520 18783 -2452
rect 18851 -2520 18864 -2452
rect 3649 -2533 3864 -2525
rect 6649 -2533 6864 -2525
rect 9649 -2533 9864 -2525
rect 12649 -2533 12864 -2525
rect 15649 -2533 15864 -2525
rect 2031 -2691 2315 -2543
rect 5038 -2691 5322 -2538
rect 8025 -2691 8309 -2541
rect 11066 -2691 11350 -2541
rect 14074 -2691 14358 -2543
rect 17049 -2691 17333 -2524
rect 18428 -2525 18864 -2520
rect 18649 -2533 18864 -2525
rect 19145 -2327 19775 -2266
rect 19145 -2691 19764 -2327
rect 2031 -2975 19764 -2691
rect 21320 -2388 26393 -1671
rect 21320 -3268 21909 -2388
rect 16771 -3857 21909 -3268
rect 25804 -3300 26393 -2388
rect 27160 -1990 27444 -1938
rect 27160 -2058 27207 -1990
rect 27275 -2058 27327 -1990
rect 27395 -2058 27444 -1990
rect 27160 -2110 27444 -2058
rect 27160 -2178 27207 -2110
rect 27275 -2178 27327 -2110
rect 27395 -2178 27444 -2110
rect 27842 -1952 28057 -1938
rect 27842 -2020 27855 -1952
rect 27923 -2020 27975 -1952
rect 28043 -2020 28057 -1952
rect 27842 -2072 28057 -2020
rect 30842 -1952 31057 -1938
rect 30842 -2020 30855 -1952
rect 30923 -2020 30975 -1952
rect 31043 -2020 31057 -1952
rect 27842 -2140 27855 -2072
rect 27923 -2140 27975 -2072
rect 28043 -2107 28057 -2072
rect 29703 -2094 29800 -2071
rect 28043 -2140 28219 -2107
rect 27842 -2153 28219 -2140
rect 27160 -2265 27444 -2178
rect 29703 -2158 29720 -2094
rect 29785 -2158 29800 -2094
rect 30842 -2072 31057 -2020
rect 33842 -1952 34057 -1938
rect 33842 -2020 33855 -1952
rect 33923 -2020 33975 -1952
rect 34043 -2020 34057 -1952
rect 30842 -2140 30855 -2072
rect 30923 -2140 30975 -2072
rect 31043 -2107 31057 -2072
rect 32737 -2090 32834 -2067
rect 31043 -2140 31219 -2107
rect 30842 -2153 31219 -2140
rect 29703 -2192 29800 -2158
rect 32737 -2154 32754 -2090
rect 32819 -2154 32834 -2090
rect 33842 -2072 34057 -2020
rect 36842 -1952 37057 -1938
rect 36842 -2020 36855 -1952
rect 36923 -2020 36975 -1952
rect 37043 -2020 37057 -1952
rect 33842 -2140 33855 -2072
rect 33923 -2140 33975 -2072
rect 34043 -2107 34057 -2072
rect 35723 -2091 35820 -2068
rect 34043 -2140 34219 -2107
rect 33842 -2153 34219 -2140
rect 32737 -2188 32834 -2154
rect 29573 -2197 29800 -2192
rect 32607 -2193 32834 -2188
rect 35723 -2155 35740 -2091
rect 35805 -2155 35820 -2091
rect 36842 -2072 37057 -2020
rect 39842 -1952 40057 -1938
rect 39842 -2020 39855 -1952
rect 39923 -2020 39975 -1952
rect 40043 -2020 40057 -1952
rect 36842 -2140 36855 -2072
rect 36923 -2140 36975 -2072
rect 37043 -2107 37057 -2072
rect 38721 -2091 38818 -2068
rect 37043 -2140 37219 -2107
rect 36842 -2153 37219 -2140
rect 35723 -2189 35820 -2155
rect 38721 -2155 38738 -2091
rect 38803 -2155 38818 -2091
rect 39842 -2072 40057 -2020
rect 42842 -1952 43057 -1938
rect 42842 -2020 42855 -1952
rect 42923 -2020 42975 -1952
rect 43043 -2020 43057 -1952
rect 39842 -2140 39855 -2072
rect 39923 -2140 39975 -2072
rect 40043 -2107 40057 -2072
rect 41721 -2089 41818 -2066
rect 40043 -2140 40219 -2107
rect 39842 -2153 40219 -2140
rect 41721 -2153 41738 -2089
rect 41803 -2153 41818 -2089
rect 42842 -2072 43057 -2020
rect 42842 -2140 42855 -2072
rect 42923 -2140 42975 -2072
rect 43043 -2107 43057 -2072
rect 44718 -2091 44815 -2068
rect 43043 -2140 43219 -2107
rect 42842 -2153 43219 -2140
rect 38721 -2189 38818 -2155
rect 41721 -2187 41818 -2153
rect 29360 -2214 29800 -2197
rect 29360 -2224 29600 -2214
rect 27160 -2333 27205 -2265
rect 27273 -2333 27325 -2265
rect 27393 -2333 27444 -2265
rect 27827 -2296 28018 -2250
rect 29360 -2274 29565 -2224
rect 29360 -2278 29600 -2274
rect 29665 -2278 29720 -2214
rect 29785 -2278 29800 -2214
rect 32355 -2210 32834 -2193
rect 35593 -2194 35820 -2189
rect 38591 -2194 38818 -2189
rect 41591 -2192 41818 -2187
rect 44718 -2155 44735 -2091
rect 44800 -2155 44815 -2091
rect 44718 -2189 44815 -2155
rect 32355 -2220 32634 -2210
rect 27827 -2318 27963 -2296
rect 29360 -2297 29800 -2278
rect 30827 -2296 31018 -2250
rect 32355 -2270 32560 -2220
rect 32610 -2270 32634 -2220
rect 32355 -2274 32634 -2270
rect 32699 -2274 32754 -2210
rect 32819 -2274 32834 -2210
rect 35368 -2211 35820 -2194
rect 35368 -2221 35620 -2211
rect 32355 -2293 32834 -2274
rect 33827 -2296 34018 -2250
rect 35368 -2271 35573 -2221
rect 35368 -2275 35620 -2271
rect 35685 -2275 35740 -2211
rect 35805 -2275 35820 -2211
rect 38367 -2211 38818 -2194
rect 38367 -2221 38618 -2211
rect 35368 -2294 35820 -2275
rect 36827 -2296 37018 -2250
rect 38367 -2271 38572 -2221
rect 38367 -2275 38618 -2271
rect 38683 -2275 38738 -2211
rect 38803 -2275 38818 -2211
rect 41368 -2209 41818 -2192
rect 44588 -2194 44815 -2189
rect 41368 -2219 41618 -2209
rect 38367 -2294 38818 -2275
rect 39827 -2296 40018 -2250
rect 41368 -2269 41573 -2219
rect 41368 -2273 41618 -2269
rect 41683 -2273 41738 -2209
rect 41803 -2273 41818 -2209
rect 44364 -2211 44815 -2194
rect 44364 -2221 44615 -2211
rect 41368 -2292 41818 -2273
rect 42827 -2296 43018 -2250
rect 44364 -2271 44569 -2221
rect 44364 -2275 44615 -2271
rect 44680 -2275 44735 -2211
rect 44800 -2275 44815 -2211
rect 44364 -2294 44815 -2275
rect 30827 -2318 30963 -2296
rect 33827 -2318 33963 -2296
rect 36827 -2318 36963 -2296
rect 39827 -2318 39963 -2296
rect 42827 -2318 42963 -2296
rect 27160 -2385 27444 -2333
rect 27160 -2453 27205 -2385
rect 27273 -2453 27325 -2385
rect 27393 -2453 27444 -2385
rect 27160 -2766 27444 -2453
rect 27697 -2332 27963 -2318
rect 27697 -2400 27710 -2332
rect 27778 -2400 27830 -2332
rect 27898 -2400 27963 -2332
rect 27697 -2452 27963 -2400
rect 27697 -2520 27710 -2452
rect 27778 -2520 27830 -2452
rect 27898 -2479 27963 -2452
rect 30697 -2332 30963 -2318
rect 30697 -2400 30710 -2332
rect 30778 -2400 30830 -2332
rect 30898 -2400 30963 -2332
rect 30697 -2452 30963 -2400
rect 27898 -2520 28133 -2479
rect 27697 -2525 28133 -2520
rect 30697 -2520 30710 -2452
rect 30778 -2520 30830 -2452
rect 30898 -2479 30963 -2452
rect 33697 -2332 33963 -2318
rect 33697 -2400 33710 -2332
rect 33778 -2400 33830 -2332
rect 33898 -2400 33963 -2332
rect 33697 -2452 33963 -2400
rect 30898 -2520 31133 -2479
rect 30697 -2525 31133 -2520
rect 33697 -2520 33710 -2452
rect 33778 -2520 33830 -2452
rect 33898 -2479 33963 -2452
rect 36697 -2332 36963 -2318
rect 36697 -2400 36710 -2332
rect 36778 -2400 36830 -2332
rect 36898 -2400 36963 -2332
rect 36697 -2452 36963 -2400
rect 33898 -2520 34133 -2479
rect 33697 -2525 34133 -2520
rect 36697 -2520 36710 -2452
rect 36778 -2520 36830 -2452
rect 36898 -2479 36963 -2452
rect 39697 -2332 39963 -2318
rect 39697 -2400 39710 -2332
rect 39778 -2400 39830 -2332
rect 39898 -2400 39963 -2332
rect 39697 -2452 39963 -2400
rect 36898 -2520 37133 -2479
rect 36697 -2525 37133 -2520
rect 39697 -2520 39710 -2452
rect 39778 -2520 39830 -2452
rect 39898 -2479 39963 -2452
rect 42697 -2332 42963 -2318
rect 42697 -2400 42710 -2332
rect 42778 -2400 42830 -2332
rect 42898 -2400 42963 -2332
rect 42697 -2452 42963 -2400
rect 39898 -2520 40133 -2479
rect 39697 -2525 40133 -2520
rect 42697 -2520 42710 -2452
rect 42778 -2520 42830 -2452
rect 42898 -2479 42963 -2452
rect 42898 -2520 43133 -2479
rect 42697 -2525 43133 -2520
rect 27697 -2533 27912 -2525
rect 30697 -2533 30912 -2525
rect 33697 -2533 33912 -2525
rect 36697 -2533 36912 -2525
rect 29208 -2766 29492 -2540
rect 32225 -2766 32509 -2541
rect 35206 -2766 35490 -2548
rect 38225 -2766 38509 -2530
rect 39697 -2533 39912 -2525
rect 42697 -2533 42912 -2525
rect 41211 -2766 41495 -2545
rect 44210 -2766 44494 -2544
rect 27079 -3050 44668 -2766
rect 16771 -3864 17360 -3857
rect -191 -4650 17360 -3864
rect -191 -7880 335 -4650
rect 16771 -6785 17360 -4650
rect 24358 -3889 29371 -3300
rect 24358 -4841 24947 -3889
rect 25524 -4708 25779 -4693
rect 25524 -4773 25549 -4708
rect 25615 -4773 25682 -4708
rect 25748 -4773 25779 -4708
rect 25524 -4832 25779 -4773
rect 25524 -4834 25683 -4832
rect 25524 -4899 25551 -4834
rect 25617 -4897 25683 -4834
rect 25749 -4897 25779 -4832
rect 25617 -4899 25779 -4897
rect 25524 -4914 25779 -4899
rect 25550 -5165 25730 -4914
rect 25887 -6311 26142 -6296
rect 25887 -6376 25912 -6311
rect 25978 -6376 26045 -6311
rect 26111 -6376 26142 -6311
rect 25887 -6435 26142 -6376
rect 25887 -6437 26046 -6435
rect 25887 -6467 25914 -6437
rect 25821 -6502 25914 -6467
rect 25980 -6500 26046 -6437
rect 26112 -6500 26142 -6435
rect 25980 -6502 26142 -6500
rect 25821 -6517 26142 -6502
rect 25821 -6623 26106 -6517
rect 28782 -6769 29371 -3889
rect 9037 -6978 9252 -6964
rect 1865 -7008 2080 -6994
rect 1865 -7076 1879 -7008
rect 1947 -7076 1999 -7008
rect 2067 -7076 2080 -7008
rect 1865 -7128 2080 -7076
rect 1865 -7196 1879 -7128
rect 1947 -7196 1999 -7128
rect 2067 -7196 2080 -7128
rect 1865 -7209 2080 -7196
rect 2191 -7007 2406 -6993
rect 2191 -7075 2205 -7007
rect 2273 -7075 2325 -7007
rect 2393 -7075 2406 -7007
rect 2191 -7127 2406 -7075
rect 2191 -7195 2205 -7127
rect 2273 -7195 2325 -7127
rect 2393 -7195 2406 -7127
rect 9037 -7046 9051 -6978
rect 9119 -7046 9171 -6978
rect 9239 -7046 9252 -6978
rect 10114 -7005 10796 -6892
rect 18637 -6978 18852 -6964
rect 9037 -7098 9252 -7046
rect 9037 -7166 9051 -7098
rect 9119 -7166 9171 -7098
rect 9239 -7166 9252 -7098
rect 9037 -7179 9252 -7166
rect 11465 -7008 11680 -6994
rect 11465 -7076 11479 -7008
rect 11547 -7076 11599 -7008
rect 11667 -7076 11680 -7008
rect 11465 -7128 11680 -7076
rect 2191 -7208 2406 -7195
rect 10113 -7298 10795 -7185
rect 11465 -7196 11479 -7128
rect 11547 -7196 11599 -7128
rect 11667 -7196 11680 -7128
rect 11465 -7209 11680 -7196
rect 11791 -7007 12006 -6993
rect 11791 -7075 11805 -7007
rect 11873 -7075 11925 -7007
rect 11993 -7075 12006 -7007
rect 11791 -7127 12006 -7075
rect 11791 -7195 11805 -7127
rect 11873 -7195 11925 -7127
rect 11993 -7195 12006 -7127
rect 18637 -7046 18651 -6978
rect 18719 -7046 18771 -6978
rect 18839 -7046 18852 -6978
rect 27709 -6978 27924 -6964
rect 18637 -7098 18852 -7046
rect 26271 -7021 26526 -7006
rect 26271 -7048 26296 -7021
rect 18637 -7166 18651 -7098
rect 18719 -7166 18771 -7098
rect 18839 -7166 18852 -7098
rect 18637 -7179 18852 -7166
rect 25865 -7086 26296 -7048
rect 26362 -7086 26429 -7021
rect 26495 -7086 26526 -7021
rect 25865 -7145 26526 -7086
rect 25865 -7147 26430 -7145
rect 11791 -7208 12006 -7195
rect 25865 -7208 26298 -7147
rect 26271 -7212 26298 -7208
rect 26364 -7210 26430 -7147
rect 26496 -7210 26526 -7145
rect 27709 -7046 27722 -6978
rect 27790 -7046 27842 -6978
rect 27910 -7046 27924 -6978
rect 27709 -7098 27924 -7046
rect 27709 -7166 27722 -7098
rect 27790 -7166 27842 -7098
rect 27910 -7166 27924 -7098
rect 27709 -7179 27924 -7166
rect 34555 -7007 34770 -6993
rect 34555 -7075 34568 -7007
rect 34636 -7075 34688 -7007
rect 34756 -7075 34770 -7007
rect 34555 -7127 34770 -7075
rect 34555 -7195 34568 -7127
rect 34636 -7195 34688 -7127
rect 34756 -7195 34770 -7127
rect 34555 -7208 34770 -7195
rect 34881 -7008 35096 -6994
rect 34881 -7076 34894 -7008
rect 34962 -7076 35014 -7008
rect 35082 -7076 35096 -7008
rect 35766 -7063 36448 -6950
rect 37309 -6978 37524 -6964
rect 37309 -7046 37322 -6978
rect 37390 -7046 37442 -6978
rect 37510 -7046 37524 -6978
rect 34881 -7128 35096 -7076
rect 34881 -7196 34894 -7128
rect 34962 -7196 35014 -7128
rect 35082 -7196 35096 -7128
rect 37309 -7098 37524 -7046
rect 37309 -7166 37322 -7098
rect 37390 -7166 37442 -7098
rect 37510 -7166 37524 -7098
rect 37309 -7179 37524 -7166
rect 44155 -7007 44370 -6993
rect 44155 -7075 44168 -7007
rect 44236 -7075 44288 -7007
rect 44356 -7075 44370 -7007
rect 44155 -7127 44370 -7075
rect 34881 -7209 35096 -7196
rect 44155 -7195 44168 -7127
rect 44236 -7195 44288 -7127
rect 44356 -7195 44370 -7127
rect 44155 -7208 44370 -7195
rect 44481 -7008 44696 -6994
rect 44481 -7076 44494 -7008
rect 44562 -7076 44614 -7008
rect 44682 -7076 44696 -7008
rect 44481 -7128 44696 -7076
rect 44481 -7196 44494 -7128
rect 44562 -7196 44614 -7128
rect 44682 -7196 44696 -7128
rect 44481 -7209 44696 -7196
rect 26364 -7212 26526 -7210
rect 26271 -7227 26526 -7212
rect 35769 -7395 36451 -7282
rect 20590 -7474 20757 -7424
rect 20590 -7487 20805 -7474
rect 20361 -7566 20470 -7539
rect 20361 -7593 20385 -7566
rect 10113 -7738 10795 -7625
rect 20327 -7632 20385 -7593
rect 20451 -7593 20470 -7566
rect 20590 -7593 20757 -7487
rect 20451 -7632 21045 -7593
rect 20327 -7696 21045 -7632
rect 20327 -7762 20385 -7696
rect 20451 -7760 21045 -7696
rect 35766 -7729 36448 -7616
rect 20451 -7762 20496 -7760
rect 20327 -7826 20496 -7762
rect -191 -8406 1202 -7880
rect 20327 -7892 20385 -7826
rect 20451 -7886 20496 -7826
rect 20590 -7886 20757 -7760
rect 20451 -7892 25877 -7886
rect 10112 -8024 10794 -7911
rect 20327 -7956 25877 -7892
rect 20327 -8022 20385 -7956
rect 20451 -8022 25877 -7956
rect 20327 -8053 25877 -8022
rect 35770 -8081 36452 -7968
rect 10115 -8273 10797 -8160
rect 35769 -8365 36451 -8252
rect -191 -9164 335 -8406
rect 10114 -8614 10796 -8501
rect 35770 -8666 36452 -8553
rect 2179 -8981 2394 -8967
rect 2179 -9049 2193 -8981
rect 2261 -9049 2313 -8981
rect 2381 -9049 2394 -8981
rect 2179 -9101 2394 -9049
rect -191 -9615 1202 -9164
rect 2179 -9169 2193 -9101
rect 2261 -9169 2313 -9101
rect 2381 -9169 2394 -9101
rect 2179 -9182 2394 -9169
rect 9225 -8990 9440 -8976
rect 9225 -9058 9239 -8990
rect 9307 -9058 9359 -8990
rect 9427 -9058 9440 -8990
rect 10112 -9006 10794 -8893
rect 11779 -8981 11994 -8967
rect 9225 -9110 9440 -9058
rect 9225 -9178 9239 -9110
rect 9307 -9178 9359 -9110
rect 9427 -9178 9440 -9110
rect 9225 -9191 9440 -9178
rect 11779 -9049 11793 -8981
rect 11861 -9049 11913 -8981
rect 11981 -9049 11994 -8981
rect 11779 -9101 11994 -9049
rect 11779 -9169 11793 -9101
rect 11861 -9169 11913 -9101
rect 11981 -9169 11994 -9101
rect 11779 -9182 11994 -9169
rect 18825 -8990 19040 -8976
rect 18825 -9058 18839 -8990
rect 18907 -9058 18959 -8990
rect 19027 -9058 19040 -8990
rect 18825 -9110 19040 -9058
rect 18825 -9178 18839 -9110
rect 18907 -9178 18959 -9110
rect 19027 -9178 19040 -9110
rect 18825 -9191 19040 -9178
rect 9356 -9256 9440 -9191
rect 18973 -9243 19040 -9191
rect 19671 -9194 26883 -8870
rect 27521 -8990 27736 -8976
rect 27521 -9058 27534 -8990
rect 27602 -9058 27654 -8990
rect 27722 -9058 27736 -8990
rect 27521 -9110 27736 -9058
rect 27521 -9178 27534 -9110
rect 27602 -9178 27654 -9110
rect 27722 -9178 27736 -9110
rect 27521 -9191 27736 -9178
rect 34567 -8981 34782 -8967
rect 34567 -9049 34580 -8981
rect 34648 -9049 34700 -8981
rect 34768 -9049 34782 -8981
rect 35767 -9041 36449 -8928
rect 37121 -8990 37336 -8976
rect 34567 -9101 34782 -9049
rect 34567 -9169 34580 -9101
rect 34648 -9169 34700 -9101
rect 34768 -9169 34782 -9101
rect 34567 -9182 34782 -9169
rect 37121 -9058 37134 -8990
rect 37202 -9058 37254 -8990
rect 37322 -9058 37336 -8990
rect 37121 -9110 37336 -9058
rect 37121 -9178 37134 -9110
rect 37202 -9178 37254 -9110
rect 37322 -9178 37336 -9110
rect 37121 -9191 37336 -9178
rect 44167 -8981 44382 -8967
rect 44167 -9049 44180 -8981
rect 44248 -9049 44300 -8981
rect 44368 -9049 44382 -8981
rect 44167 -9101 44382 -9049
rect 44167 -9169 44180 -9101
rect 44248 -9169 44300 -9101
rect 44368 -9169 44382 -9101
rect 44167 -9182 44382 -9169
rect 27521 -9243 27588 -9191
rect 37121 -9256 37205 -9191
rect 10112 -9410 10794 -9297
rect 35768 -9429 36450 -9316
rect -191 -9823 1251 -9615
rect 19686 -9625 26880 -9433
rect 19660 -9817 26905 -9625
rect 19660 -9823 20120 -9817
rect -191 -10061 20120 -9823
rect 26291 -9823 26905 -9817
rect 45311 -9823 45837 -6781
rect 26291 -10061 45837 -9823
rect -191 -10349 45837 -10061
<< via1 >>
rect 1770 13266 1841 13337
rect 1913 13263 1984 13334
rect 1770 13134 1841 13205
rect 1913 13134 1984 13205
rect 1769 13007 1840 13078
rect 1912 13004 1983 13075
rect 1769 12875 1840 12946
rect 1912 12875 1983 12946
rect 19204 -1900 19272 -1832
rect 19324 -1900 19392 -1832
rect 19518 -1897 19586 -1829
rect 19638 -1897 19706 -1829
rect 3518 -2020 3586 -1952
rect 3638 -2020 3706 -1952
rect 1748 -2158 1813 -2094
rect 6518 -2020 6586 -1952
rect 6638 -2020 6706 -1952
rect 3518 -2140 3586 -2072
rect 3638 -2140 3706 -2072
rect 4749 -2158 4814 -2094
rect 6518 -2140 6586 -2072
rect 6638 -2140 6706 -2072
rect 9518 -2020 9586 -1952
rect 9638 -2020 9706 -1952
rect 12518 -2020 12586 -1952
rect 12638 -2020 12706 -1952
rect 7765 -2161 7830 -2097
rect 9518 -2140 9586 -2072
rect 9638 -2140 9706 -2072
rect 1748 -2278 1813 -2214
rect 1868 -2278 1933 -2214
rect 10762 -2158 10827 -2094
rect 15518 -2020 15586 -1952
rect 15638 -2020 15706 -1952
rect 12518 -2140 12586 -2072
rect 12638 -2140 12706 -2072
rect 13791 -2156 13856 -2092
rect 18518 -2020 18586 -1952
rect 18638 -2020 18706 -1952
rect 15518 -2140 15586 -2072
rect 15638 -2140 15706 -2072
rect 16822 -2158 16887 -2094
rect 18518 -2140 18586 -2072
rect 18638 -2140 18706 -2072
rect 19204 -2020 19272 -1952
rect 19324 -2020 19392 -1952
rect 19518 -2017 19586 -1949
rect 19638 -2017 19706 -1949
rect 19206 -2146 19274 -2078
rect 19326 -2146 19394 -2078
rect 19520 -2143 19588 -2075
rect 19640 -2143 19708 -2075
rect 4749 -2278 4814 -2214
rect 4869 -2278 4934 -2214
rect 7765 -2281 7830 -2217
rect 7885 -2281 7950 -2217
rect 10762 -2278 10827 -2214
rect 10882 -2278 10947 -2214
rect 13791 -2276 13856 -2212
rect 13911 -2220 13976 -2212
rect 13911 -2270 13956 -2220
rect 13956 -2270 13976 -2220
rect 13911 -2276 13976 -2270
rect 16822 -2278 16887 -2214
rect 16942 -2220 17007 -2214
rect 16942 -2270 16949 -2220
rect 16949 -2270 16999 -2220
rect 16999 -2270 17007 -2220
rect 16942 -2278 17007 -2270
rect 19206 -2266 19274 -2198
rect 19326 -2266 19394 -2198
rect 19520 -2263 19588 -2195
rect 19640 -2263 19708 -2195
rect 3663 -2400 3731 -2332
rect 3783 -2400 3851 -2332
rect 3663 -2520 3731 -2452
rect 3783 -2520 3851 -2452
rect 6663 -2400 6731 -2332
rect 6783 -2400 6851 -2332
rect 6663 -2520 6731 -2452
rect 6783 -2520 6851 -2452
rect 9663 -2400 9731 -2332
rect 9783 -2400 9851 -2332
rect 9663 -2520 9731 -2452
rect 9783 -2520 9851 -2452
rect 12663 -2400 12731 -2332
rect 12783 -2400 12851 -2332
rect 12663 -2520 12731 -2452
rect 12783 -2520 12851 -2452
rect 15663 -2400 15731 -2332
rect 15783 -2400 15851 -2332
rect 15663 -2520 15731 -2452
rect 15783 -2520 15851 -2452
rect 18663 -2400 18731 -2332
rect 18783 -2400 18851 -2332
rect 18663 -2520 18731 -2452
rect 18783 -2520 18851 -2452
rect 27207 -2058 27275 -1990
rect 27327 -2058 27395 -1990
rect 27207 -2178 27275 -2110
rect 27327 -2178 27395 -2110
rect 27855 -2020 27923 -1952
rect 27975 -2020 28043 -1952
rect 30855 -2020 30923 -1952
rect 30975 -2020 31043 -1952
rect 27855 -2140 27923 -2072
rect 27975 -2140 28043 -2072
rect 29720 -2158 29785 -2094
rect 33855 -2020 33923 -1952
rect 33975 -2020 34043 -1952
rect 30855 -2140 30923 -2072
rect 30975 -2140 31043 -2072
rect 32754 -2154 32819 -2090
rect 36855 -2020 36923 -1952
rect 36975 -2020 37043 -1952
rect 33855 -2140 33923 -2072
rect 33975 -2140 34043 -2072
rect 35740 -2155 35805 -2091
rect 39855 -2020 39923 -1952
rect 39975 -2020 40043 -1952
rect 36855 -2140 36923 -2072
rect 36975 -2140 37043 -2072
rect 38738 -2155 38803 -2091
rect 42855 -2020 42923 -1952
rect 42975 -2020 43043 -1952
rect 39855 -2140 39923 -2072
rect 39975 -2140 40043 -2072
rect 41738 -2153 41803 -2089
rect 42855 -2140 42923 -2072
rect 42975 -2140 43043 -2072
rect 29600 -2224 29665 -2214
rect 27205 -2333 27273 -2265
rect 27325 -2333 27393 -2265
rect 29600 -2274 29615 -2224
rect 29615 -2274 29665 -2224
rect 29600 -2278 29665 -2274
rect 29720 -2278 29785 -2214
rect 44735 -2155 44800 -2091
rect 32634 -2274 32699 -2210
rect 32754 -2274 32819 -2210
rect 35620 -2221 35685 -2211
rect 35620 -2271 35623 -2221
rect 35623 -2271 35685 -2221
rect 35620 -2275 35685 -2271
rect 35740 -2275 35805 -2211
rect 38618 -2221 38683 -2211
rect 38618 -2271 38622 -2221
rect 38622 -2271 38683 -2221
rect 38618 -2275 38683 -2271
rect 38738 -2275 38803 -2211
rect 41618 -2219 41683 -2209
rect 41618 -2269 41623 -2219
rect 41623 -2269 41683 -2219
rect 41618 -2273 41683 -2269
rect 41738 -2273 41803 -2209
rect 44615 -2221 44680 -2211
rect 44615 -2271 44619 -2221
rect 44619 -2271 44680 -2221
rect 44615 -2275 44680 -2271
rect 44735 -2275 44800 -2211
rect 27205 -2453 27273 -2385
rect 27325 -2453 27393 -2385
rect 27710 -2400 27778 -2332
rect 27830 -2400 27898 -2332
rect 27710 -2520 27778 -2452
rect 27830 -2520 27898 -2452
rect 30710 -2400 30778 -2332
rect 30830 -2400 30898 -2332
rect 30710 -2520 30778 -2452
rect 30830 -2520 30898 -2452
rect 33710 -2400 33778 -2332
rect 33830 -2400 33898 -2332
rect 33710 -2520 33778 -2452
rect 33830 -2520 33898 -2452
rect 36710 -2400 36778 -2332
rect 36830 -2400 36898 -2332
rect 36710 -2520 36778 -2452
rect 36830 -2520 36898 -2452
rect 39710 -2400 39778 -2332
rect 39830 -2400 39898 -2332
rect 39710 -2520 39778 -2452
rect 39830 -2520 39898 -2452
rect 42710 -2400 42778 -2332
rect 42830 -2400 42898 -2332
rect 42710 -2520 42778 -2452
rect 42830 -2520 42898 -2452
rect 25549 -4773 25615 -4708
rect 25682 -4773 25748 -4708
rect 25551 -4899 25617 -4834
rect 25683 -4897 25749 -4832
rect 25912 -6376 25978 -6311
rect 26045 -6376 26111 -6311
rect 25914 -6502 25980 -6437
rect 26046 -6500 26112 -6435
rect 1879 -7076 1947 -7008
rect 1999 -7076 2067 -7008
rect 1879 -7196 1947 -7128
rect 1999 -7196 2067 -7128
rect 2205 -7075 2273 -7007
rect 2325 -7075 2393 -7007
rect 2205 -7195 2273 -7127
rect 2325 -7195 2393 -7127
rect 9051 -7046 9119 -6978
rect 9171 -7046 9239 -6978
rect 9051 -7166 9119 -7098
rect 9171 -7166 9239 -7098
rect 11479 -7076 11547 -7008
rect 11599 -7076 11667 -7008
rect 11479 -7196 11547 -7128
rect 11599 -7196 11667 -7128
rect 11805 -7075 11873 -7007
rect 11925 -7075 11993 -7007
rect 11805 -7195 11873 -7127
rect 11925 -7195 11993 -7127
rect 18651 -7046 18719 -6978
rect 18771 -7046 18839 -6978
rect 18651 -7166 18719 -7098
rect 18771 -7166 18839 -7098
rect 26296 -7086 26362 -7021
rect 26429 -7086 26495 -7021
rect 26298 -7212 26364 -7147
rect 26430 -7210 26496 -7145
rect 27722 -7046 27790 -6978
rect 27842 -7046 27910 -6978
rect 27722 -7166 27790 -7098
rect 27842 -7166 27910 -7098
rect 34568 -7075 34636 -7007
rect 34688 -7075 34756 -7007
rect 34568 -7195 34636 -7127
rect 34688 -7195 34756 -7127
rect 34894 -7076 34962 -7008
rect 35014 -7076 35082 -7008
rect 37322 -7046 37390 -6978
rect 37442 -7046 37510 -6978
rect 34894 -7196 34962 -7128
rect 35014 -7196 35082 -7128
rect 37322 -7166 37390 -7098
rect 37442 -7166 37510 -7098
rect 44168 -7075 44236 -7007
rect 44288 -7075 44356 -7007
rect 44168 -7195 44236 -7127
rect 44288 -7195 44356 -7127
rect 44494 -7076 44562 -7008
rect 44614 -7076 44682 -7008
rect 44494 -7196 44562 -7128
rect 44614 -7196 44682 -7128
rect 20385 -7632 20451 -7566
rect 20385 -7762 20451 -7696
rect 20385 -7892 20451 -7826
rect 20385 -8022 20451 -7956
rect 2193 -9049 2261 -8981
rect 2313 -9049 2381 -8981
rect 2193 -9169 2261 -9101
rect 2313 -9169 2381 -9101
rect 9239 -9058 9307 -8990
rect 9359 -9058 9427 -8990
rect 9239 -9178 9307 -9110
rect 9359 -9178 9427 -9110
rect 11793 -9049 11861 -8981
rect 11913 -9049 11981 -8981
rect 11793 -9169 11861 -9101
rect 11913 -9169 11981 -9101
rect 18839 -9058 18907 -8990
rect 18959 -9058 19027 -8990
rect 18839 -9178 18907 -9110
rect 18959 -9178 19027 -9110
rect 27534 -9058 27602 -8990
rect 27654 -9058 27722 -8990
rect 27534 -9178 27602 -9110
rect 27654 -9178 27722 -9110
rect 34580 -9049 34648 -8981
rect 34700 -9049 34768 -8981
rect 34580 -9169 34648 -9101
rect 34700 -9169 34768 -9101
rect 37134 -9058 37202 -8990
rect 37254 -9058 37322 -8990
rect 37134 -9178 37202 -9110
rect 37254 -9178 37322 -9110
rect 44180 -9049 44248 -8981
rect 44300 -9049 44368 -8981
rect 44180 -9169 44248 -9101
rect 44300 -9169 44368 -9101
<< metal2 >>
rect -2576 15008 3325 15050
rect -2576 14508 3331 15008
rect -2576 -887 -2034 14508
rect 2984 13990 3331 14508
rect -1676 13337 2140 13391
rect 2530 13366 2690 13791
rect 2984 13742 3277 13990
rect 2984 13582 3331 13742
rect -1676 13266 1770 13337
rect 1841 13334 2140 13337
rect 1841 13266 1913 13334
rect -1676 13263 1913 13266
rect 1984 13263 2140 13334
rect -1676 13205 2140 13263
rect -1676 13134 1770 13205
rect 1841 13134 1913 13205
rect 1984 13134 2140 13205
rect -1676 13078 2140 13134
rect -1676 13007 1769 13078
rect 1840 13075 2140 13078
rect 1840 13007 1912 13075
rect -1676 13004 1912 13007
rect 1983 13004 2140 13075
rect -1676 12946 2140 13004
rect -1676 12875 1769 12946
rect 1840 12875 1912 12946
rect 1983 12875 2140 12946
rect -1676 12849 2140 12875
rect -1676 -182 -1134 12849
rect -1676 -724 21718 -182
rect 21176 -779 21718 -724
rect -2576 -1429 19550 -887
rect 21176 -1321 45815 -779
rect 3538 -1938 3679 -1429
rect 6538 -1938 6679 -1429
rect 9538 -1938 9679 -1429
rect 12538 -1938 12679 -1429
rect 15538 -1938 15679 -1429
rect 18538 -1938 18679 -1429
rect 19168 -1829 19775 -1779
rect 19168 -1832 19518 -1829
rect 19168 -1900 19204 -1832
rect 19272 -1900 19324 -1832
rect 19392 -1897 19518 -1832
rect 19586 -1897 19638 -1829
rect 19706 -1830 19775 -1829
rect 19706 -1897 27465 -1830
rect 19392 -1900 27465 -1897
rect 3504 -1952 3719 -1938
rect 3504 -2020 3518 -1952
rect 3586 -2020 3638 -1952
rect 3706 -2020 3719 -1952
rect 1700 -2094 1856 -2061
rect 1700 -2158 1748 -2094
rect 1813 -2158 1856 -2094
rect 3504 -2072 3719 -2020
rect 6504 -1952 6719 -1938
rect 6504 -2020 6518 -1952
rect 6586 -2020 6638 -1952
rect 6706 -2020 6719 -1952
rect 9504 -1952 9719 -1938
rect 3504 -2140 3518 -2072
rect 3586 -2140 3638 -2072
rect 3706 -2140 3719 -2072
rect 3504 -2153 3719 -2140
rect 4714 -2094 4870 -2061
rect 1700 -2192 1856 -2158
rect 4714 -2158 4749 -2094
rect 4814 -2158 4870 -2094
rect 6504 -2072 6719 -2020
rect 6504 -2140 6518 -2072
rect 6586 -2140 6638 -2072
rect 6706 -2140 6719 -2072
rect 6504 -2153 6719 -2140
rect 7728 -2097 7884 -2014
rect 4714 -2192 4870 -2158
rect 7728 -2161 7765 -2097
rect 7830 -2161 7884 -2097
rect 9504 -2020 9518 -1952
rect 9586 -2020 9638 -1952
rect 9706 -2020 9719 -1952
rect 9504 -2072 9719 -2020
rect 12504 -1952 12719 -1938
rect 12504 -2020 12518 -1952
rect 12586 -2020 12638 -1952
rect 12706 -2020 12719 -1952
rect 15504 -1952 15719 -1938
rect 9504 -2140 9518 -2072
rect 9586 -2140 9638 -2072
rect 9706 -2140 9719 -2072
rect 9504 -2153 9719 -2140
rect 10695 -2094 10851 -2046
rect 1700 -2214 1937 -2192
rect 1700 -2278 1748 -2214
rect 1813 -2278 1868 -2214
rect 1933 -2278 1937 -2214
rect 1700 -2297 1937 -2278
rect 4714 -2214 4938 -2192
rect 4714 -2278 4749 -2214
rect 4814 -2278 4869 -2214
rect 4934 -2278 4938 -2214
rect 4714 -2297 4938 -2278
rect 7728 -2195 7884 -2161
rect 10695 -2158 10762 -2094
rect 10827 -2158 10851 -2094
rect 12504 -2072 12719 -2020
rect 12504 -2140 12518 -2072
rect 12586 -2140 12638 -2072
rect 12706 -2140 12719 -2072
rect 12504 -2153 12719 -2140
rect 13724 -2092 13880 -1998
rect 10695 -2192 10851 -2158
rect 13724 -2156 13791 -2092
rect 13856 -2156 13880 -2092
rect 15504 -2020 15518 -1952
rect 15586 -2020 15638 -1952
rect 15706 -2020 15719 -1952
rect 18504 -1952 18719 -1938
rect 15504 -2072 15719 -2020
rect 15504 -2140 15518 -2072
rect 15586 -2140 15638 -2072
rect 15706 -2140 15719 -2072
rect 15504 -2153 15719 -2140
rect 16754 -2094 16910 -1982
rect 13724 -2190 13880 -2156
rect 16754 -2158 16822 -2094
rect 16887 -2158 16910 -2094
rect 18504 -2020 18518 -1952
rect 18586 -2020 18638 -1952
rect 18706 -2020 18719 -1952
rect 18504 -2072 18719 -2020
rect 18504 -2140 18518 -2072
rect 18586 -2140 18638 -2072
rect 18706 -2140 18719 -2072
rect 18504 -2153 18719 -2140
rect 19168 -1949 27465 -1900
rect 27882 -1938 28023 -1321
rect 30882 -1938 31023 -1321
rect 33882 -1938 34023 -1321
rect 36882 -1938 37023 -1321
rect 39882 -1938 40023 -1321
rect 42882 -1938 43023 -1321
rect 19168 -1952 19518 -1949
rect 19168 -2020 19204 -1952
rect 19272 -2020 19324 -1952
rect 19392 -2017 19518 -1952
rect 19586 -2017 19638 -1949
rect 19706 -1962 27465 -1949
rect 19706 -1965 20570 -1962
rect 19706 -2017 20313 -1965
rect 19392 -2020 20313 -2017
rect 19168 -2033 20313 -2020
rect 20381 -2033 20433 -1965
rect 20501 -2030 20570 -1965
rect 20638 -2030 20690 -1962
rect 20758 -1990 27465 -1962
rect 20758 -2030 27207 -1990
rect 20501 -2033 27207 -2030
rect 19168 -2058 27207 -2033
rect 27275 -2058 27327 -1990
rect 27395 -2058 27465 -1990
rect 19168 -2075 27465 -2058
rect 19168 -2078 19520 -2075
rect 19168 -2146 19206 -2078
rect 19274 -2146 19326 -2078
rect 19394 -2143 19520 -2078
rect 19588 -2143 19640 -2075
rect 19708 -2082 27465 -2075
rect 19708 -2085 20570 -2082
rect 19708 -2143 20313 -2085
rect 19394 -2146 20313 -2143
rect 19168 -2153 20313 -2146
rect 20381 -2153 20433 -2085
rect 20501 -2150 20570 -2085
rect 20638 -2150 20690 -2082
rect 20758 -2110 27465 -2082
rect 20758 -2150 27207 -2110
rect 20501 -2153 27207 -2150
rect 7728 -2217 7977 -2195
rect 7728 -2281 7765 -2217
rect 7830 -2281 7885 -2217
rect 7950 -2281 7977 -2217
rect 1700 -3927 1856 -2297
rect 3649 -2332 3864 -2318
rect 3649 -2400 3663 -2332
rect 3731 -2400 3783 -2332
rect 3851 -2400 3864 -2332
rect 3649 -2452 3864 -2400
rect 3649 -2520 3663 -2452
rect 3731 -2520 3783 -2452
rect 3851 -2520 3864 -2452
rect 3649 -2533 3864 -2520
rect 4714 -3687 4870 -2297
rect 7728 -2300 7977 -2281
rect 10695 -2214 10974 -2192
rect 10695 -2278 10762 -2214
rect 10827 -2278 10882 -2214
rect 10947 -2278 10974 -2214
rect 10695 -2297 10974 -2278
rect 13724 -2212 14003 -2190
rect 13724 -2276 13791 -2212
rect 13856 -2276 13911 -2212
rect 13976 -2276 14003 -2212
rect 13724 -2295 14003 -2276
rect 16754 -2192 16910 -2158
rect 19168 -2178 27207 -2153
rect 27275 -2178 27327 -2110
rect 27395 -2178 27465 -2110
rect 27842 -1952 28057 -1938
rect 27842 -2020 27855 -1952
rect 27923 -2020 27975 -1952
rect 28043 -2020 28057 -1952
rect 27842 -2072 28057 -2020
rect 30842 -1952 31057 -1938
rect 30842 -2020 30855 -1952
rect 30923 -2020 30975 -1952
rect 31043 -2020 31057 -1952
rect 33842 -1952 34057 -1938
rect 27842 -2140 27855 -2072
rect 27923 -2140 27975 -2072
rect 28043 -2140 28057 -2072
rect 27842 -2153 28057 -2140
rect 29663 -2094 29819 -2030
rect 16754 -2214 17034 -2192
rect 16754 -2278 16822 -2214
rect 16887 -2278 16942 -2214
rect 17007 -2278 17034 -2214
rect 6649 -2332 6864 -2318
rect 6649 -2400 6663 -2332
rect 6731 -2400 6783 -2332
rect 6851 -2400 6864 -2332
rect 6649 -2452 6864 -2400
rect 6649 -2520 6663 -2452
rect 6731 -2520 6783 -2452
rect 6851 -2520 6864 -2452
rect 6649 -2533 6864 -2520
rect 7728 -3447 7884 -2300
rect 9649 -2332 9864 -2318
rect 9649 -2400 9663 -2332
rect 9731 -2400 9783 -2332
rect 9851 -2400 9864 -2332
rect 9649 -2452 9864 -2400
rect 9649 -2520 9663 -2452
rect 9731 -2520 9783 -2452
rect 9851 -2520 9864 -2452
rect 9649 -2533 9864 -2520
rect 10695 -3207 10851 -2297
rect 12649 -2332 12864 -2318
rect 12649 -2400 12663 -2332
rect 12731 -2400 12783 -2332
rect 12851 -2400 12864 -2332
rect 12649 -2452 12864 -2400
rect 12649 -2520 12663 -2452
rect 12731 -2520 12783 -2452
rect 12851 -2520 12864 -2452
rect 12649 -2533 12864 -2520
rect 13724 -2967 13880 -2295
rect 16754 -2297 17034 -2278
rect 19168 -2195 27465 -2178
rect 29663 -2158 29720 -2094
rect 29785 -2158 29819 -2094
rect 30842 -2072 31057 -2020
rect 30842 -2140 30855 -2072
rect 30923 -2140 30975 -2072
rect 31043 -2140 31057 -2072
rect 30842 -2153 31057 -2140
rect 32724 -2090 32880 -1998
rect 29663 -2192 29819 -2158
rect 32724 -2154 32754 -2090
rect 32819 -2154 32880 -2090
rect 33842 -2020 33855 -1952
rect 33923 -2020 33975 -1952
rect 34043 -2020 34057 -1952
rect 33842 -2072 34057 -2020
rect 36842 -1952 37057 -1938
rect 36842 -2020 36855 -1952
rect 36923 -2020 36975 -1952
rect 37043 -2020 37057 -1952
rect 33842 -2140 33855 -2072
rect 33923 -2140 33975 -2072
rect 34043 -2140 34057 -2072
rect 33842 -2153 34057 -2140
rect 35722 -2091 35878 -2046
rect 32724 -2188 32880 -2154
rect 19168 -2198 19520 -2195
rect 19168 -2266 19206 -2198
rect 19274 -2266 19326 -2198
rect 19394 -2263 19520 -2198
rect 19588 -2263 19640 -2195
rect 19708 -2263 27465 -2195
rect 19394 -2264 27465 -2263
rect 19394 -2266 19775 -2264
rect 15649 -2332 15864 -2318
rect 15649 -2400 15663 -2332
rect 15731 -2400 15783 -2332
rect 15851 -2400 15864 -2332
rect 15649 -2452 15864 -2400
rect 15649 -2520 15663 -2452
rect 15731 -2520 15783 -2452
rect 15851 -2520 15864 -2452
rect 15649 -2533 15864 -2520
rect 16754 -2727 16910 -2297
rect 18649 -2332 18864 -2318
rect 19168 -2327 19775 -2266
rect 27146 -2265 27465 -2264
rect 18649 -2400 18663 -2332
rect 18731 -2400 18783 -2332
rect 18851 -2400 18864 -2332
rect 18649 -2452 18864 -2400
rect 18649 -2520 18663 -2452
rect 18731 -2520 18783 -2452
rect 18851 -2520 18864 -2452
rect 27146 -2333 27205 -2265
rect 27273 -2333 27325 -2265
rect 27393 -2333 27465 -2265
rect 29573 -2214 29819 -2192
rect 29573 -2278 29600 -2214
rect 29665 -2278 29720 -2214
rect 29785 -2278 29819 -2214
rect 29573 -2297 29819 -2278
rect 32607 -2210 32880 -2188
rect 35722 -2155 35740 -2091
rect 35805 -2155 35878 -2091
rect 36842 -2072 37057 -2020
rect 39842 -1952 40057 -1938
rect 39842 -2020 39855 -1952
rect 39923 -2020 39975 -1952
rect 40043 -2020 40057 -1952
rect 36842 -2140 36855 -2072
rect 36923 -2140 36975 -2072
rect 37043 -2140 37057 -2072
rect 36842 -2153 37057 -2140
rect 38689 -2091 38845 -2046
rect 35722 -2189 35878 -2155
rect 38689 -2155 38738 -2091
rect 38803 -2155 38845 -2091
rect 39842 -2072 40057 -2020
rect 42842 -1952 43057 -1938
rect 42842 -2020 42855 -1952
rect 42923 -2020 42975 -1952
rect 43043 -2020 43057 -1952
rect 39842 -2140 39855 -2072
rect 39923 -2140 39975 -2072
rect 40043 -2140 40057 -2072
rect 39842 -2153 40057 -2140
rect 41703 -2089 41859 -2046
rect 41703 -2153 41738 -2089
rect 41803 -2153 41859 -2089
rect 42842 -2072 43057 -2020
rect 42842 -2140 42855 -2072
rect 42923 -2140 42975 -2072
rect 43043 -2140 43057 -2072
rect 42842 -2153 43057 -2140
rect 44685 -2091 44841 -1998
rect 38689 -2189 38845 -2155
rect 41703 -2187 41859 -2153
rect 32607 -2274 32634 -2210
rect 32699 -2274 32754 -2210
rect 32819 -2274 32880 -2210
rect 32607 -2293 32880 -2274
rect 27146 -2385 27465 -2333
rect 27146 -2453 27205 -2385
rect 27273 -2453 27325 -2385
rect 27393 -2453 27465 -2385
rect 27146 -2511 27465 -2453
rect 27697 -2332 27912 -2318
rect 27697 -2400 27710 -2332
rect 27778 -2400 27830 -2332
rect 27898 -2400 27912 -2332
rect 27697 -2452 27912 -2400
rect 18649 -2533 18864 -2520
rect 27697 -2520 27710 -2452
rect 27778 -2520 27830 -2452
rect 27898 -2520 27912 -2452
rect 27697 -2533 27912 -2520
rect 29663 -2727 29819 -2297
rect 30697 -2332 30912 -2318
rect 30697 -2400 30710 -2332
rect 30778 -2400 30830 -2332
rect 30898 -2400 30912 -2332
rect 30697 -2452 30912 -2400
rect 30697 -2520 30710 -2452
rect 30778 -2520 30830 -2452
rect 30898 -2520 30912 -2452
rect 30697 -2533 30912 -2520
rect 16754 -2773 29866 -2727
rect 16754 -2829 26445 -2773
rect 26501 -2775 29866 -2773
rect 26501 -2829 26574 -2775
rect 16754 -2831 26574 -2829
rect 26630 -2778 29866 -2775
rect 26630 -2831 26713 -2778
rect 16754 -2834 26713 -2831
rect 26769 -2834 29866 -2778
rect 16754 -2883 29866 -2834
rect 32724 -2967 32880 -2293
rect 35593 -2211 35878 -2189
rect 35593 -2275 35620 -2211
rect 35685 -2275 35740 -2211
rect 35805 -2275 35878 -2211
rect 35593 -2294 35878 -2275
rect 38591 -2211 38845 -2189
rect 38591 -2275 38618 -2211
rect 38683 -2275 38738 -2211
rect 38803 -2275 38845 -2211
rect 38591 -2294 38845 -2275
rect 41591 -2209 41859 -2187
rect 44685 -2155 44735 -2091
rect 44800 -2155 44841 -2091
rect 44685 -2189 44841 -2155
rect 41591 -2273 41618 -2209
rect 41683 -2273 41738 -2209
rect 41803 -2273 41859 -2209
rect 41591 -2292 41859 -2273
rect 33697 -2332 33912 -2318
rect 33697 -2400 33710 -2332
rect 33778 -2400 33830 -2332
rect 33898 -2400 33912 -2332
rect 33697 -2452 33912 -2400
rect 33697 -2520 33710 -2452
rect 33778 -2520 33830 -2452
rect 33898 -2520 33912 -2452
rect 33697 -2533 33912 -2520
rect 13677 -3005 32975 -2967
rect 13677 -3061 25434 -3005
rect 25490 -3007 32975 -3005
rect 25490 -3061 25563 -3007
rect 13677 -3063 25563 -3061
rect 25619 -3010 32975 -3007
rect 25619 -3063 25702 -3010
rect 13677 -3066 25702 -3063
rect 25758 -3066 32975 -3010
rect 13677 -3123 32975 -3066
rect 35722 -3207 35878 -2294
rect 36697 -2332 36912 -2318
rect 36697 -2400 36710 -2332
rect 36778 -2400 36830 -2332
rect 36898 -2400 36912 -2332
rect 36697 -2452 36912 -2400
rect 36697 -2520 36710 -2452
rect 36778 -2520 36830 -2452
rect 36898 -2520 36912 -2452
rect 36697 -2533 36912 -2520
rect 10600 -3256 35973 -3207
rect 10600 -3312 25905 -3256
rect 25961 -3258 35973 -3256
rect 25961 -3312 26034 -3258
rect 10600 -3314 26034 -3312
rect 26090 -3261 35973 -3258
rect 26090 -3314 26173 -3261
rect 10600 -3317 26173 -3314
rect 26229 -3317 35973 -3261
rect 10600 -3363 35973 -3317
rect 38689 -3447 38845 -2294
rect 39697 -2332 39912 -2318
rect 39697 -2400 39710 -2332
rect 39778 -2400 39830 -2332
rect 39898 -2400 39912 -2332
rect 39697 -2452 39912 -2400
rect 39697 -2520 39710 -2452
rect 39778 -2520 39830 -2452
rect 39898 -2520 39912 -2452
rect 39697 -2533 39912 -2520
rect 7633 -3495 38955 -3447
rect 7633 -3551 23649 -3495
rect 23705 -3497 38955 -3495
rect 23705 -3551 23778 -3497
rect 7633 -3553 23778 -3551
rect 23834 -3500 38955 -3497
rect 23834 -3553 23917 -3500
rect 7633 -3556 23917 -3553
rect 23973 -3556 38955 -3500
rect 7633 -3603 38955 -3556
rect 41703 -3687 41859 -2292
rect 44588 -2211 44841 -2189
rect 44588 -2275 44615 -2211
rect 44680 -2275 44735 -2211
rect 44800 -2275 44841 -2211
rect 44588 -2294 44841 -2275
rect 42697 -2332 42912 -2318
rect 42697 -2400 42710 -2332
rect 42778 -2400 42830 -2332
rect 42898 -2400 42912 -2332
rect 42697 -2452 42912 -2400
rect 42697 -2520 42710 -2452
rect 42778 -2520 42830 -2452
rect 42898 -2520 42912 -2452
rect 42697 -2533 42912 -2520
rect 4587 -3736 41859 -3687
rect 4587 -3792 23098 -3736
rect 23154 -3739 41859 -3736
rect 23154 -3792 23213 -3739
rect 4587 -3795 23213 -3792
rect 23269 -3795 23328 -3739
rect 23384 -3795 41859 -3739
rect 4587 -3843 41859 -3795
rect 44685 -3927 44841 -2294
rect 1700 -4083 45126 -3927
rect 9441 -4247 9656 -4233
rect 9441 -4251 9455 -4247
rect 836 -4315 9455 -4251
rect 9523 -4315 9575 -4247
rect 9643 -4251 9656 -4247
rect 19041 -4247 19256 -4233
rect 19041 -4251 19055 -4247
rect 9643 -4315 19055 -4251
rect 19123 -4315 19175 -4247
rect 19243 -4251 19256 -4247
rect 19243 -4292 20095 -4251
rect 19243 -4315 19331 -4292
rect 836 -4360 19331 -4315
rect 19399 -4360 19451 -4292
rect 19519 -4293 20095 -4292
rect 19519 -4296 19887 -4293
rect 19519 -4360 19579 -4296
rect 836 -4364 19579 -4360
rect 19647 -4364 19699 -4296
rect 19767 -4361 19887 -4296
rect 19955 -4361 20007 -4293
rect 20075 -4361 20095 -4293
rect 19767 -4364 20095 -4361
rect 836 -4367 20095 -4364
rect 836 -4435 9455 -4367
rect 9523 -4435 9575 -4367
rect 9643 -4435 19055 -4367
rect 19123 -4435 19175 -4367
rect 19243 -4435 20095 -4367
rect 836 -4451 20095 -4435
rect 20309 -4347 20812 -4328
rect 20309 -4350 20607 -4347
rect 20309 -4418 20350 -4350
rect 20418 -4418 20470 -4350
rect 20538 -4415 20607 -4350
rect 20675 -4415 20727 -4347
rect 20795 -4415 20812 -4347
rect 20538 -4418 20812 -4415
rect 20309 -4467 20812 -4418
rect 20309 -4470 20607 -4467
rect 1012 -4548 1227 -4534
rect 1012 -4551 1026 -4548
rect 836 -4616 1026 -4551
rect 1094 -4616 1146 -4548
rect 1214 -4551 1227 -4548
rect 10612 -4548 10827 -4534
rect 20309 -4538 20350 -4470
rect 20418 -4538 20470 -4470
rect 20538 -4535 20607 -4470
rect 20675 -4535 20727 -4467
rect 20795 -4535 20812 -4467
rect 22753 -4500 22903 -4083
rect 23098 -4229 23326 -4211
rect 22970 -4285 23126 -4229
rect 23182 -4230 23326 -4229
rect 23182 -4285 23244 -4230
rect 22753 -4503 22875 -4500
rect 20538 -4538 20812 -4535
rect 10612 -4551 10626 -4548
rect 1214 -4616 10626 -4551
rect 10694 -4616 10746 -4548
rect 10814 -4551 10827 -4548
rect 18288 -4551 18503 -4541
rect 10814 -4555 20097 -4551
rect 10814 -4616 18302 -4555
rect 836 -4623 18302 -4616
rect 18370 -4623 18422 -4555
rect 18490 -4623 20097 -4555
rect 20309 -4567 20812 -4538
rect 836 -4668 20097 -4623
rect 836 -4736 1026 -4668
rect 1094 -4736 1146 -4668
rect 1214 -4736 10626 -4668
rect 10694 -4736 10746 -4668
rect 10814 -4675 20097 -4668
rect 10814 -4736 18302 -4675
rect 836 -4743 18302 -4736
rect 18370 -4743 18422 -4675
rect 18490 -4743 20097 -4675
rect 836 -4751 20097 -4743
rect 18288 -4756 18503 -4751
rect 9862 -4851 10077 -4839
rect 15640 -4851 15855 -4841
rect 19462 -4851 19677 -4839
rect 836 -4853 20097 -4851
rect 836 -4921 9876 -4853
rect 9944 -4921 9996 -4853
rect 10064 -4855 19476 -4853
rect 10064 -4921 15654 -4855
rect 836 -4923 15654 -4921
rect 15722 -4923 15774 -4855
rect 15842 -4921 19476 -4855
rect 19544 -4921 19596 -4853
rect 19664 -4921 20097 -4853
rect 15842 -4923 20097 -4921
rect 836 -4973 20097 -4923
rect 836 -5041 9876 -4973
rect 9944 -5041 9996 -4973
rect 10064 -4975 19476 -4973
rect 10064 -5041 15654 -4975
rect 836 -5043 15654 -5041
rect 15722 -5043 15774 -4975
rect 15842 -5041 19476 -4975
rect 19544 -5041 19596 -4973
rect 19664 -5041 20097 -4973
rect 15842 -5043 20097 -5041
rect 836 -5051 20097 -5043
rect 9862 -5054 10077 -5051
rect 15640 -5056 15855 -5051
rect 19462 -5054 19677 -5051
rect 1407 -5151 1622 -5150
rect 11007 -5151 11222 -5150
rect 12639 -5151 12854 -5141
rect 836 -5155 20097 -5151
rect 836 -5164 12653 -5155
rect 836 -5232 1421 -5164
rect 1489 -5232 1541 -5164
rect 1609 -5232 11021 -5164
rect 11089 -5232 11141 -5164
rect 11209 -5223 12653 -5164
rect 12721 -5223 12773 -5155
rect 12841 -5223 20097 -5155
rect 11209 -5232 20097 -5223
rect 836 -5275 20097 -5232
rect 836 -5284 12653 -5275
rect 836 -5351 1421 -5284
rect 1407 -5352 1421 -5351
rect 1489 -5352 1541 -5284
rect 1609 -5351 11021 -5284
rect 1609 -5352 1622 -5351
rect 1407 -5365 1622 -5352
rect 11007 -5352 11021 -5351
rect 11089 -5352 11141 -5284
rect 11209 -5343 12653 -5284
rect 12721 -5343 12773 -5275
rect 12841 -5343 20097 -5275
rect 11209 -5351 20097 -5343
rect 11209 -5352 11222 -5351
rect 11007 -5365 11222 -5352
rect 12639 -5356 12854 -5351
rect 8569 -5444 8784 -5430
rect 8569 -5451 8583 -5444
rect 836 -5512 8583 -5451
rect 8651 -5512 8703 -5444
rect 8771 -5451 8784 -5444
rect 18169 -5444 18384 -5430
rect 18169 -5451 18183 -5444
rect 8771 -5512 18183 -5451
rect 18251 -5512 18303 -5444
rect 18371 -5451 18384 -5444
rect 18371 -5512 20097 -5451
rect 836 -5564 20097 -5512
rect 836 -5632 8583 -5564
rect 8651 -5632 8703 -5564
rect 8771 -5632 18183 -5564
rect 18251 -5632 18303 -5564
rect 18371 -5632 20097 -5564
rect 836 -5651 20097 -5632
rect 2184 -5751 2399 -5749
rect 6639 -5751 6854 -5739
rect 11784 -5751 11999 -5749
rect 836 -5753 20097 -5751
rect 836 -5763 6653 -5753
rect 836 -5831 2198 -5763
rect 2266 -5831 2318 -5763
rect 2386 -5821 6653 -5763
rect 6721 -5821 6773 -5753
rect 6841 -5763 20097 -5753
rect 6841 -5821 11798 -5763
rect 2386 -5831 11798 -5821
rect 11866 -5831 11918 -5763
rect 11986 -5831 20097 -5763
rect 836 -5873 20097 -5831
rect 836 -5883 6653 -5873
rect 836 -5951 2198 -5883
rect 2266 -5951 2318 -5883
rect 2386 -5941 6653 -5883
rect 6721 -5941 6773 -5873
rect 6841 -5883 20097 -5873
rect 6841 -5941 11798 -5883
rect 2386 -5951 11798 -5941
rect 11866 -5951 11918 -5883
rect 11986 -5951 20097 -5883
rect 2184 -5964 2399 -5951
rect 6639 -5954 6854 -5951
rect 11784 -5964 11999 -5951
rect 3637 -6051 3852 -6039
rect 9020 -6050 9235 -6036
rect 9020 -6051 9034 -6050
rect 836 -6053 9034 -6051
rect 836 -6121 3651 -6053
rect 3719 -6121 3771 -6053
rect 3839 -6118 9034 -6053
rect 9102 -6118 9154 -6050
rect 9222 -6051 9235 -6050
rect 18620 -6050 18835 -6036
rect 18620 -6051 18634 -6050
rect 9222 -6118 18634 -6051
rect 18702 -6118 18754 -6050
rect 18822 -6051 18835 -6050
rect 18822 -6118 20097 -6051
rect 3839 -6121 20097 -6118
rect 836 -6170 20097 -6121
rect 836 -6173 9034 -6170
rect 836 -6241 3651 -6173
rect 3719 -6241 3771 -6173
rect 3839 -6238 9034 -6173
rect 9102 -6238 9154 -6170
rect 9222 -6238 18634 -6170
rect 18702 -6238 18754 -6170
rect 18822 -6238 20097 -6170
rect 3839 -6241 20097 -6238
rect 836 -6251 20097 -6241
rect 3637 -6254 3852 -6251
rect 1860 -6351 2075 -6341
rect 11460 -6351 11675 -6341
rect -412 -6355 20097 -6351
rect -412 -6423 1874 -6355
rect 1942 -6423 1994 -6355
rect 2062 -6423 11474 -6355
rect 11542 -6423 11594 -6355
rect 11662 -6423 20097 -6355
rect -412 -6475 20097 -6423
rect -412 -6543 1874 -6475
rect 1942 -6543 1994 -6475
rect 2062 -6543 11474 -6475
rect 11542 -6543 11594 -6475
rect 11662 -6543 20097 -6475
rect -412 -6551 20097 -6543
rect 1860 -6556 2075 -6551
rect 11460 -6556 11675 -6551
rect 8580 -6883 8795 -6869
rect 8580 -6951 8594 -6883
rect 8662 -6951 8714 -6883
rect 8782 -6951 8795 -6883
rect 1865 -7008 2080 -6994
rect 1865 -7076 1879 -7008
rect 1947 -7076 1999 -7008
rect 2067 -7076 2080 -7008
rect 1865 -7128 2080 -7076
rect 1865 -7196 1879 -7128
rect 1947 -7196 1999 -7128
rect 2067 -7196 2080 -7128
rect 1865 -7209 2080 -7196
rect 2191 -7007 2406 -6993
rect 2191 -7075 2205 -7007
rect 2273 -7075 2325 -7007
rect 2393 -7075 2406 -7007
rect 2191 -7127 2406 -7075
rect 8580 -7003 8795 -6951
rect 18180 -6883 18395 -6869
rect 18180 -6951 18194 -6883
rect 18262 -6951 18314 -6883
rect 18382 -6951 18395 -6883
rect 8580 -7071 8594 -7003
rect 8662 -7071 8714 -7003
rect 8782 -7071 8795 -7003
rect 8580 -7084 8795 -7071
rect 9037 -6978 9252 -6964
rect 9037 -7046 9051 -6978
rect 9119 -7046 9171 -6978
rect 9239 -7046 9252 -6978
rect 2191 -7195 2205 -7127
rect 2273 -7195 2325 -7127
rect 2393 -7195 2406 -7127
rect 9037 -7098 9252 -7046
rect 9037 -7166 9051 -7098
rect 9119 -7166 9171 -7098
rect 9239 -7166 9252 -7098
rect 9037 -7179 9252 -7166
rect 11465 -7008 11680 -6994
rect 11465 -7076 11479 -7008
rect 11547 -7076 11599 -7008
rect 11667 -7076 11680 -7008
rect 11465 -7128 11680 -7076
rect 2191 -7208 2406 -7195
rect 11465 -7196 11479 -7128
rect 11547 -7196 11599 -7128
rect 11667 -7196 11680 -7128
rect 11465 -7209 11680 -7196
rect 11791 -7007 12006 -6993
rect 11791 -7075 11805 -7007
rect 11873 -7075 11925 -7007
rect 11993 -7075 12006 -7007
rect 11791 -7127 12006 -7075
rect 18180 -7003 18395 -6951
rect 18180 -7071 18194 -7003
rect 18262 -7071 18314 -7003
rect 18382 -7071 18395 -7003
rect 18180 -7084 18395 -7071
rect 18637 -6978 18852 -6964
rect 18637 -7046 18651 -6978
rect 18719 -7046 18771 -6978
rect 18839 -7046 18852 -6978
rect 11791 -7195 11805 -7127
rect 11873 -7195 11925 -7127
rect 11993 -7195 12006 -7127
rect 18637 -7098 18852 -7046
rect 18637 -7166 18651 -7098
rect 18719 -7166 18771 -7098
rect 18839 -7166 18852 -7098
rect 18637 -7179 18852 -7166
rect 11791 -7208 12006 -7195
rect 20327 -7566 20523 -4567
rect 22970 -4627 23026 -4285
rect 23098 -4286 23244 -4285
rect 23300 -4286 23326 -4230
rect 27305 -4247 27520 -4233
rect 27305 -4251 27318 -4247
rect 23098 -4303 23326 -4286
rect 26825 -4315 27318 -4251
rect 27386 -4315 27438 -4247
rect 27506 -4251 27520 -4247
rect 36905 -4247 37120 -4233
rect 36905 -4251 36918 -4247
rect 27506 -4291 36918 -4251
rect 27506 -4294 29847 -4291
rect 27506 -4315 29539 -4294
rect 26825 -4362 29539 -4315
rect 29607 -4362 29659 -4294
rect 29727 -4359 29847 -4294
rect 29915 -4359 29967 -4291
rect 30035 -4293 36918 -4291
rect 30035 -4359 30138 -4293
rect 29727 -4361 30138 -4359
rect 30206 -4361 30258 -4293
rect 30326 -4315 36918 -4293
rect 36986 -4315 37038 -4247
rect 37106 -4251 37120 -4247
rect 37106 -4315 45725 -4251
rect 30326 -4361 45725 -4315
rect 29727 -4362 45725 -4361
rect 26825 -4367 45725 -4362
rect 23659 -4449 23905 -4425
rect 23659 -4451 23686 -4449
rect 23093 -4505 23686 -4451
rect 23742 -4450 23905 -4449
rect 23742 -4505 23820 -4450
rect 23093 -4506 23820 -4505
rect 23876 -4506 23905 -4450
rect 26825 -4435 27318 -4367
rect 27386 -4435 27438 -4367
rect 27506 -4435 36918 -4367
rect 36986 -4435 37038 -4367
rect 37106 -4435 45725 -4367
rect 26825 -4451 45725 -4435
rect 23093 -4507 23905 -4506
rect 23093 -4719 23149 -4507
rect 23659 -4524 23905 -4507
rect 28058 -4551 28273 -4541
rect 35734 -4548 35949 -4534
rect 35734 -4551 35747 -4548
rect 26825 -4555 35747 -4551
rect 26825 -4623 28071 -4555
rect 28139 -4623 28191 -4555
rect 28259 -4616 35747 -4555
rect 35815 -4616 35867 -4548
rect 35935 -4551 35949 -4548
rect 45334 -4548 45549 -4534
rect 45334 -4551 45347 -4548
rect 35935 -4616 45347 -4551
rect 45415 -4616 45467 -4548
rect 45535 -4551 45549 -4548
rect 45535 -4616 45725 -4551
rect 28259 -4623 45725 -4616
rect 26825 -4668 45725 -4623
rect 26825 -4675 35747 -4668
rect 25524 -4708 25779 -4693
rect 25524 -4773 25549 -4708
rect 25615 -4773 25682 -4708
rect 25748 -4773 25779 -4708
rect 26825 -4743 28071 -4675
rect 28139 -4743 28191 -4675
rect 28259 -4736 35747 -4675
rect 35815 -4736 35867 -4668
rect 35935 -4736 45347 -4668
rect 45415 -4736 45467 -4668
rect 45535 -4736 45725 -4668
rect 28259 -4743 45725 -4736
rect 26825 -4751 45725 -4743
rect 28058 -4756 28273 -4751
rect 25524 -4832 25779 -4773
rect 25524 -4834 25683 -4832
rect 25524 -4899 25551 -4834
rect 25617 -4897 25683 -4834
rect 25749 -4897 25779 -4832
rect 26884 -4851 27099 -4839
rect 30706 -4851 30921 -4841
rect 36484 -4851 36699 -4839
rect 25617 -4899 25779 -4897
rect 25524 -4914 25779 -4899
rect 26825 -4853 45725 -4851
rect 26825 -4921 26897 -4853
rect 26965 -4921 27017 -4853
rect 27085 -4855 36497 -4853
rect 27085 -4921 30719 -4855
rect 26825 -4923 30719 -4921
rect 30787 -4923 30839 -4855
rect 30907 -4921 36497 -4855
rect 36565 -4921 36617 -4853
rect 36685 -4921 45725 -4853
rect 30907 -4923 45725 -4921
rect 26825 -4973 45725 -4923
rect 26825 -5041 26897 -4973
rect 26965 -5041 27017 -4973
rect 27085 -4975 36497 -4973
rect 27085 -5041 30719 -4975
rect 26825 -5043 30719 -5041
rect 30787 -5043 30839 -4975
rect 30907 -5041 36497 -4975
rect 36565 -5041 36617 -4973
rect 36685 -5041 45725 -4973
rect 30907 -5043 45725 -5041
rect 26825 -5051 45725 -5043
rect 26884 -5054 27099 -5051
rect 30706 -5056 30921 -5051
rect 36484 -5054 36699 -5051
rect 33707 -5151 33922 -5141
rect 35339 -5151 35554 -5150
rect 44939 -5151 45154 -5150
rect 26825 -5155 45725 -5151
rect 26825 -5223 33720 -5155
rect 33788 -5223 33840 -5155
rect 33908 -5164 45725 -5155
rect 33908 -5223 35352 -5164
rect 26825 -5232 35352 -5223
rect 35420 -5232 35472 -5164
rect 35540 -5232 44952 -5164
rect 45020 -5232 45072 -5164
rect 45140 -5232 45725 -5164
rect 26825 -5275 45725 -5232
rect 26825 -5343 33720 -5275
rect 33788 -5343 33840 -5275
rect 33908 -5284 45725 -5275
rect 33908 -5343 35352 -5284
rect 26825 -5351 35352 -5343
rect 33707 -5356 33922 -5351
rect 35339 -5352 35352 -5351
rect 35420 -5352 35472 -5284
rect 35540 -5351 44952 -5284
rect 35540 -5352 35554 -5351
rect 35339 -5365 35554 -5352
rect 44939 -5352 44952 -5351
rect 45020 -5352 45072 -5284
rect 45140 -5351 45725 -5284
rect 45140 -5352 45154 -5351
rect 44939 -5365 45154 -5352
rect 28177 -5444 28392 -5430
rect 28177 -5451 28190 -5444
rect 26825 -5512 28190 -5451
rect 28258 -5512 28310 -5444
rect 28378 -5451 28392 -5444
rect 37777 -5444 37992 -5430
rect 37777 -5451 37790 -5444
rect 28378 -5512 37790 -5451
rect 37858 -5512 37910 -5444
rect 37978 -5451 37992 -5444
rect 37978 -5512 45725 -5451
rect 26825 -5564 45725 -5512
rect 26825 -5632 28190 -5564
rect 28258 -5632 28310 -5564
rect 28378 -5632 37790 -5564
rect 37858 -5632 37910 -5564
rect 37978 -5632 45725 -5564
rect 26825 -5651 45725 -5632
rect 34562 -5751 34777 -5749
rect 39707 -5751 39922 -5739
rect 44162 -5751 44377 -5749
rect 26825 -5753 45725 -5751
rect 26825 -5763 39720 -5753
rect 26825 -5831 34575 -5763
rect 34643 -5831 34695 -5763
rect 34763 -5821 39720 -5763
rect 39788 -5821 39840 -5753
rect 39908 -5763 45725 -5753
rect 39908 -5821 44175 -5763
rect 34763 -5831 44175 -5821
rect 44243 -5831 44295 -5763
rect 44363 -5831 45725 -5763
rect 26825 -5873 45725 -5831
rect 26825 -5883 39720 -5873
rect 26825 -5951 34575 -5883
rect 34643 -5951 34695 -5883
rect 34763 -5941 39720 -5883
rect 39788 -5941 39840 -5873
rect 39908 -5883 45725 -5873
rect 39908 -5941 44175 -5883
rect 34763 -5951 44175 -5941
rect 44243 -5951 44295 -5883
rect 44363 -5951 45725 -5883
rect 34562 -5964 34777 -5951
rect 39707 -5954 39922 -5951
rect 44162 -5964 44377 -5951
rect 27726 -6050 27941 -6036
rect 27726 -6051 27739 -6050
rect 26825 -6118 27739 -6051
rect 27807 -6118 27859 -6050
rect 27927 -6051 27941 -6050
rect 37326 -6050 37541 -6036
rect 37326 -6051 37339 -6050
rect 27927 -6118 37339 -6051
rect 37407 -6118 37459 -6050
rect 37527 -6051 37541 -6050
rect 42709 -6051 42924 -6039
rect 37527 -6053 45725 -6051
rect 37527 -6118 42722 -6053
rect 26825 -6121 42722 -6118
rect 42790 -6121 42842 -6053
rect 42910 -6121 45725 -6053
rect 26825 -6170 45725 -6121
rect 26825 -6238 27739 -6170
rect 27807 -6238 27859 -6170
rect 27927 -6238 37339 -6170
rect 37407 -6238 37459 -6170
rect 37527 -6173 45725 -6170
rect 37527 -6238 42722 -6173
rect 26825 -6241 42722 -6238
rect 42790 -6241 42842 -6173
rect 42910 -6241 45725 -6173
rect 26825 -6251 45725 -6241
rect 42709 -6254 42924 -6251
rect 25887 -6311 26142 -6296
rect 25887 -6376 25912 -6311
rect 25978 -6376 26045 -6311
rect 26111 -6376 26142 -6311
rect 34886 -6351 35101 -6341
rect 44486 -6351 44701 -6341
rect 25887 -6435 26142 -6376
rect 25887 -6437 26046 -6435
rect 25887 -6502 25914 -6437
rect 25980 -6500 26046 -6437
rect 26112 -6500 26142 -6435
rect 25980 -6502 26142 -6500
rect 25887 -6517 26142 -6502
rect 26825 -6355 46780 -6351
rect 26825 -6423 34899 -6355
rect 34967 -6423 35019 -6355
rect 35087 -6423 44499 -6355
rect 44567 -6423 44619 -6355
rect 44687 -6423 46780 -6355
rect 26825 -6475 46780 -6423
rect 26825 -6543 34899 -6475
rect 34967 -6543 35019 -6475
rect 35087 -6543 44499 -6475
rect 44567 -6543 44619 -6475
rect 44687 -6543 46780 -6475
rect 26825 -6551 46780 -6543
rect 34886 -6556 35101 -6551
rect 44486 -6556 44701 -6551
rect 28166 -6883 28381 -6869
rect 28166 -6951 28179 -6883
rect 28247 -6951 28299 -6883
rect 28367 -6951 28381 -6883
rect 27709 -6978 27924 -6964
rect 26271 -7021 26526 -7006
rect 26271 -7086 26296 -7021
rect 26362 -7086 26429 -7021
rect 26495 -7086 26526 -7021
rect 26271 -7145 26526 -7086
rect 26271 -7147 26430 -7145
rect 26271 -7212 26298 -7147
rect 26364 -7210 26430 -7147
rect 26496 -7210 26526 -7145
rect 27709 -7046 27722 -6978
rect 27790 -7046 27842 -6978
rect 27910 -7046 27924 -6978
rect 27709 -7098 27924 -7046
rect 28166 -7003 28381 -6951
rect 37766 -6883 37981 -6869
rect 37766 -6951 37779 -6883
rect 37847 -6951 37899 -6883
rect 37967 -6951 37981 -6883
rect 37309 -6978 37524 -6964
rect 28166 -7071 28179 -7003
rect 28247 -7071 28299 -7003
rect 28367 -7071 28381 -7003
rect 28166 -7084 28381 -7071
rect 34555 -7007 34770 -6993
rect 34555 -7075 34568 -7007
rect 34636 -7075 34688 -7007
rect 34756 -7075 34770 -7007
rect 27709 -7166 27722 -7098
rect 27790 -7166 27842 -7098
rect 27910 -7166 27924 -7098
rect 27709 -7179 27924 -7166
rect 34555 -7127 34770 -7075
rect 34555 -7195 34568 -7127
rect 34636 -7195 34688 -7127
rect 34756 -7195 34770 -7127
rect 34555 -7208 34770 -7195
rect 34881 -7008 35096 -6994
rect 34881 -7076 34894 -7008
rect 34962 -7076 35014 -7008
rect 35082 -7076 35096 -7008
rect 34881 -7128 35096 -7076
rect 34881 -7196 34894 -7128
rect 34962 -7196 35014 -7128
rect 35082 -7196 35096 -7128
rect 37309 -7046 37322 -6978
rect 37390 -7046 37442 -6978
rect 37510 -7046 37524 -6978
rect 37309 -7098 37524 -7046
rect 37766 -7003 37981 -6951
rect 37766 -7071 37779 -7003
rect 37847 -7071 37899 -7003
rect 37967 -7071 37981 -7003
rect 37766 -7084 37981 -7071
rect 44155 -7007 44370 -6993
rect 44155 -7075 44168 -7007
rect 44236 -7075 44288 -7007
rect 44356 -7075 44370 -7007
rect 37309 -7166 37322 -7098
rect 37390 -7166 37442 -7098
rect 37510 -7166 37524 -7098
rect 37309 -7179 37524 -7166
rect 44155 -7127 44370 -7075
rect 34881 -7209 35096 -7196
rect 44155 -7195 44168 -7127
rect 44236 -7195 44288 -7127
rect 44356 -7195 44370 -7127
rect 44155 -7208 44370 -7195
rect 44481 -7008 44696 -6994
rect 44481 -7076 44494 -7008
rect 44562 -7076 44614 -7008
rect 44682 -7076 44696 -7008
rect 44481 -7128 44696 -7076
rect 44481 -7196 44494 -7128
rect 44562 -7196 44614 -7128
rect 44682 -7196 44696 -7128
rect 44481 -7209 44696 -7196
rect 26364 -7212 26526 -7210
rect 26271 -7227 26526 -7212
rect 20327 -7632 20385 -7566
rect 20451 -7632 20523 -7566
rect 20327 -7696 20523 -7632
rect 20327 -7762 20385 -7696
rect 20451 -7762 20523 -7696
rect 20327 -7826 20523 -7762
rect 9863 -7844 10078 -7830
rect 9863 -7912 9877 -7844
rect 9945 -7912 9997 -7844
rect 10065 -7912 10078 -7844
rect 9863 -7964 10078 -7912
rect 9863 -8032 9877 -7964
rect 9945 -8032 9997 -7964
rect 10065 -8032 10078 -7964
rect 9863 -8045 10078 -8032
rect 19463 -7844 19678 -7830
rect 19463 -7912 19477 -7844
rect 19545 -7912 19597 -7844
rect 19665 -7912 19678 -7844
rect 19463 -7964 19678 -7912
rect 19463 -8032 19477 -7964
rect 19545 -8032 19597 -7964
rect 19665 -8032 19678 -7964
rect 19463 -8045 19678 -8032
rect 20327 -7892 20385 -7826
rect 20451 -7892 20523 -7826
rect 20327 -7956 20523 -7892
rect 20327 -8022 20385 -7956
rect 20451 -8022 20523 -7956
rect 20327 -8049 20523 -8022
rect 26883 -7844 27098 -7830
rect 26883 -7912 26896 -7844
rect 26964 -7912 27016 -7844
rect 27084 -7912 27098 -7844
rect 26883 -7964 27098 -7912
rect 26883 -8032 26896 -7964
rect 26964 -8032 27016 -7964
rect 27084 -8032 27098 -7964
rect 26883 -8045 27098 -8032
rect 36483 -7844 36698 -7830
rect 36483 -7912 36496 -7844
rect 36564 -7912 36616 -7844
rect 36684 -7912 36698 -7844
rect 36483 -7964 36698 -7912
rect 36483 -8032 36496 -7964
rect 36564 -8032 36616 -7964
rect 36684 -8032 36698 -7964
rect 36483 -8045 36698 -8032
rect 1860 -8533 2075 -8519
rect 1860 -8601 1874 -8533
rect 1942 -8601 1994 -8533
rect 2062 -8601 2075 -8533
rect 1860 -8653 2075 -8601
rect 1860 -8721 1874 -8653
rect 1942 -8721 1994 -8653
rect 2062 -8721 2075 -8653
rect 1860 -8734 2075 -8721
rect 11460 -8533 11675 -8519
rect 11460 -8601 11474 -8533
rect 11542 -8601 11594 -8533
rect 11662 -8601 11675 -8533
rect 11460 -8653 11675 -8601
rect 11460 -8721 11474 -8653
rect 11542 -8721 11594 -8653
rect 11662 -8721 11675 -8653
rect 11460 -8734 11675 -8721
rect 34886 -8533 35101 -8519
rect 34886 -8601 34899 -8533
rect 34967 -8601 35019 -8533
rect 35087 -8601 35101 -8533
rect 34886 -8653 35101 -8601
rect 34886 -8721 34899 -8653
rect 34967 -8721 35019 -8653
rect 35087 -8721 35101 -8653
rect 34886 -8734 35101 -8721
rect 44486 -8533 44701 -8519
rect 44486 -8601 44499 -8533
rect 44567 -8601 44619 -8533
rect 44687 -8601 44701 -8533
rect 44486 -8653 44701 -8601
rect 44486 -8721 44499 -8653
rect 44567 -8721 44619 -8653
rect 44687 -8721 44701 -8653
rect 44486 -8734 44701 -8721
rect 2179 -8981 2394 -8967
rect 2179 -9049 2193 -8981
rect 2261 -9049 2313 -8981
rect 2381 -9049 2394 -8981
rect 2179 -9101 2394 -9049
rect 2179 -9169 2193 -9101
rect 2261 -9169 2313 -9101
rect 2381 -9169 2394 -9101
rect 2179 -9182 2394 -9169
rect 9225 -8990 9440 -8976
rect 9225 -9058 9239 -8990
rect 9307 -9058 9359 -8990
rect 9427 -9058 9440 -8990
rect 9225 -9110 9440 -9058
rect 9225 -9178 9239 -9110
rect 9307 -9178 9359 -9110
rect 9427 -9178 9440 -9110
rect 9225 -9191 9440 -9178
rect 11779 -8981 11994 -8967
rect 11779 -9049 11793 -8981
rect 11861 -9049 11913 -8981
rect 11981 -9049 11994 -8981
rect 11779 -9101 11994 -9049
rect 11779 -9169 11793 -9101
rect 11861 -9169 11913 -9101
rect 11981 -9169 11994 -9101
rect 11779 -9182 11994 -9169
rect 18825 -8990 19040 -8976
rect 18825 -9058 18839 -8990
rect 18907 -9058 18959 -8990
rect 19027 -9058 19040 -8990
rect 18825 -9110 19040 -9058
rect 18825 -9178 18839 -9110
rect 18907 -9178 18959 -9110
rect 19027 -9178 19040 -9110
rect 18825 -9191 19040 -9178
rect 27521 -8990 27736 -8976
rect 27521 -9058 27534 -8990
rect 27602 -9058 27654 -8990
rect 27722 -9058 27736 -8990
rect 27521 -9110 27736 -9058
rect 27521 -9178 27534 -9110
rect 27602 -9178 27654 -9110
rect 27722 -9178 27736 -9110
rect 27521 -9191 27736 -9178
rect 34567 -8981 34782 -8967
rect 34567 -9049 34580 -8981
rect 34648 -9049 34700 -8981
rect 34768 -9049 34782 -8981
rect 34567 -9101 34782 -9049
rect 34567 -9169 34580 -9101
rect 34648 -9169 34700 -9101
rect 34768 -9169 34782 -9101
rect 34567 -9182 34782 -9169
rect 37121 -8990 37336 -8976
rect 37121 -9058 37134 -8990
rect 37202 -9058 37254 -8990
rect 37322 -9058 37336 -8990
rect 37121 -9110 37336 -9058
rect 37121 -9178 37134 -9110
rect 37202 -9178 37254 -9110
rect 37322 -9178 37336 -9110
rect 37121 -9191 37336 -9178
rect 44167 -8981 44382 -8967
rect 44167 -9049 44180 -8981
rect 44248 -9049 44300 -8981
rect 44368 -9049 44382 -8981
rect 44167 -9101 44382 -9049
rect 44167 -9169 44180 -9101
rect 44248 -9169 44300 -9101
rect 44368 -9169 44382 -9101
rect 44167 -9182 44382 -9169
<< via2 >>
rect 20313 -2033 20381 -1965
rect 20433 -2033 20501 -1965
rect 20570 -2030 20638 -1962
rect 20690 -2030 20758 -1962
rect 20313 -2153 20381 -2085
rect 20433 -2153 20501 -2085
rect 20570 -2150 20638 -2082
rect 20690 -2150 20758 -2082
rect 3663 -2400 3731 -2332
rect 3783 -2400 3851 -2332
rect 3663 -2520 3731 -2452
rect 3783 -2520 3851 -2452
rect 6663 -2400 6731 -2332
rect 6783 -2400 6851 -2332
rect 6663 -2520 6731 -2452
rect 6783 -2520 6851 -2452
rect 9663 -2400 9731 -2332
rect 9783 -2400 9851 -2332
rect 9663 -2520 9731 -2452
rect 9783 -2520 9851 -2452
rect 12663 -2400 12731 -2332
rect 12783 -2400 12851 -2332
rect 12663 -2520 12731 -2452
rect 12783 -2520 12851 -2452
rect 15663 -2400 15731 -2332
rect 15783 -2400 15851 -2332
rect 15663 -2520 15731 -2452
rect 15783 -2520 15851 -2452
rect 18663 -2400 18731 -2332
rect 18783 -2400 18851 -2332
rect 18663 -2520 18731 -2452
rect 18783 -2520 18851 -2452
rect 27710 -2400 27778 -2332
rect 27830 -2400 27898 -2332
rect 27710 -2520 27778 -2452
rect 27830 -2520 27898 -2452
rect 30710 -2400 30778 -2332
rect 30830 -2400 30898 -2332
rect 30710 -2520 30778 -2452
rect 30830 -2520 30898 -2452
rect 26445 -2829 26501 -2773
rect 26574 -2831 26630 -2775
rect 26713 -2834 26769 -2778
rect 33710 -2400 33778 -2332
rect 33830 -2400 33898 -2332
rect 33710 -2520 33778 -2452
rect 33830 -2520 33898 -2452
rect 25434 -3061 25490 -3005
rect 25563 -3063 25619 -3007
rect 25702 -3066 25758 -3010
rect 36710 -2400 36778 -2332
rect 36830 -2400 36898 -2332
rect 36710 -2520 36778 -2452
rect 36830 -2520 36898 -2452
rect 25905 -3312 25961 -3256
rect 26034 -3314 26090 -3258
rect 26173 -3317 26229 -3261
rect 39710 -2400 39778 -2332
rect 39830 -2400 39898 -2332
rect 39710 -2520 39778 -2452
rect 39830 -2520 39898 -2452
rect 23649 -3551 23705 -3495
rect 23778 -3553 23834 -3497
rect 23917 -3556 23973 -3500
rect 42710 -2400 42778 -2332
rect 42830 -2400 42898 -2332
rect 42710 -2520 42778 -2452
rect 42830 -2520 42898 -2452
rect 23098 -3792 23154 -3736
rect 23213 -3795 23269 -3739
rect 23328 -3795 23384 -3739
rect 9455 -4315 9523 -4247
rect 9575 -4315 9643 -4247
rect 19055 -4315 19123 -4247
rect 19175 -4315 19243 -4247
rect 19331 -4360 19399 -4292
rect 19451 -4360 19519 -4292
rect 19579 -4364 19647 -4296
rect 19699 -4364 19767 -4296
rect 19887 -4361 19955 -4293
rect 20007 -4361 20075 -4293
rect 9455 -4435 9523 -4367
rect 9575 -4435 9643 -4367
rect 19055 -4435 19123 -4367
rect 19175 -4435 19243 -4367
rect 20350 -4418 20418 -4350
rect 20470 -4418 20538 -4350
rect 20607 -4415 20675 -4347
rect 20727 -4415 20795 -4347
rect 1026 -4616 1094 -4548
rect 1146 -4616 1214 -4548
rect 20350 -4538 20418 -4470
rect 20470 -4538 20538 -4470
rect 20607 -4535 20675 -4467
rect 20727 -4535 20795 -4467
rect 23126 -4285 23182 -4229
rect 10626 -4616 10694 -4548
rect 10746 -4616 10814 -4548
rect 18302 -4623 18370 -4555
rect 18422 -4623 18490 -4555
rect 1026 -4736 1094 -4668
rect 1146 -4736 1214 -4668
rect 10626 -4736 10694 -4668
rect 10746 -4736 10814 -4668
rect 18302 -4743 18370 -4675
rect 18422 -4743 18490 -4675
rect 9876 -4921 9944 -4853
rect 9996 -4921 10064 -4853
rect 15654 -4923 15722 -4855
rect 15774 -4923 15842 -4855
rect 19476 -4921 19544 -4853
rect 19596 -4921 19664 -4853
rect 9876 -5041 9944 -4973
rect 9996 -5041 10064 -4973
rect 15654 -5043 15722 -4975
rect 15774 -5043 15842 -4975
rect 19476 -5041 19544 -4973
rect 19596 -5041 19664 -4973
rect 1421 -5232 1489 -5164
rect 1541 -5232 1609 -5164
rect 11021 -5232 11089 -5164
rect 11141 -5232 11209 -5164
rect 12653 -5223 12721 -5155
rect 12773 -5223 12841 -5155
rect 1421 -5352 1489 -5284
rect 1541 -5352 1609 -5284
rect 11021 -5352 11089 -5284
rect 11141 -5352 11209 -5284
rect 12653 -5343 12721 -5275
rect 12773 -5343 12841 -5275
rect 8583 -5512 8651 -5444
rect 8703 -5512 8771 -5444
rect 18183 -5512 18251 -5444
rect 18303 -5512 18371 -5444
rect 8583 -5632 8651 -5564
rect 8703 -5632 8771 -5564
rect 18183 -5632 18251 -5564
rect 18303 -5632 18371 -5564
rect 2198 -5831 2266 -5763
rect 2318 -5831 2386 -5763
rect 6653 -5821 6721 -5753
rect 6773 -5821 6841 -5753
rect 11798 -5831 11866 -5763
rect 11918 -5831 11986 -5763
rect 2198 -5951 2266 -5883
rect 2318 -5951 2386 -5883
rect 6653 -5941 6721 -5873
rect 6773 -5941 6841 -5873
rect 11798 -5951 11866 -5883
rect 11918 -5951 11986 -5883
rect 3651 -6121 3719 -6053
rect 3771 -6121 3839 -6053
rect 9034 -6118 9102 -6050
rect 9154 -6118 9222 -6050
rect 18634 -6118 18702 -6050
rect 18754 -6118 18822 -6050
rect 3651 -6241 3719 -6173
rect 3771 -6241 3839 -6173
rect 9034 -6238 9102 -6170
rect 9154 -6238 9222 -6170
rect 18634 -6238 18702 -6170
rect 18754 -6238 18822 -6170
rect 1874 -6423 1942 -6355
rect 1994 -6423 2062 -6355
rect 11474 -6423 11542 -6355
rect 11594 -6423 11662 -6355
rect 1874 -6543 1942 -6475
rect 1994 -6543 2062 -6475
rect 11474 -6543 11542 -6475
rect 11594 -6543 11662 -6475
rect 8594 -6951 8662 -6883
rect 8714 -6951 8782 -6883
rect 1879 -7076 1947 -7008
rect 1999 -7076 2067 -7008
rect 1879 -7196 1947 -7128
rect 1999 -7196 2067 -7128
rect 2205 -7075 2273 -7007
rect 2325 -7075 2393 -7007
rect 18194 -6951 18262 -6883
rect 18314 -6951 18382 -6883
rect 8594 -7071 8662 -7003
rect 8714 -7071 8782 -7003
rect 9051 -7046 9119 -6978
rect 9171 -7046 9239 -6978
rect 2205 -7195 2273 -7127
rect 2325 -7195 2393 -7127
rect 9051 -7166 9119 -7098
rect 9171 -7166 9239 -7098
rect 11479 -7076 11547 -7008
rect 11599 -7076 11667 -7008
rect 11479 -7196 11547 -7128
rect 11599 -7196 11667 -7128
rect 11805 -7075 11873 -7007
rect 11925 -7075 11993 -7007
rect 18194 -7071 18262 -7003
rect 18314 -7071 18382 -7003
rect 18651 -7046 18719 -6978
rect 18771 -7046 18839 -6978
rect 11805 -7195 11873 -7127
rect 11925 -7195 11993 -7127
rect 18651 -7166 18719 -7098
rect 18771 -7166 18839 -7098
rect 23244 -4286 23300 -4230
rect 27318 -4315 27386 -4247
rect 27438 -4315 27506 -4247
rect 29539 -4362 29607 -4294
rect 29659 -4362 29727 -4294
rect 29847 -4359 29915 -4291
rect 29967 -4359 30035 -4291
rect 30138 -4361 30206 -4293
rect 30258 -4361 30326 -4293
rect 36918 -4315 36986 -4247
rect 37038 -4315 37106 -4247
rect 23686 -4505 23742 -4449
rect 23820 -4506 23876 -4450
rect 27318 -4435 27386 -4367
rect 27438 -4435 27506 -4367
rect 36918 -4435 36986 -4367
rect 37038 -4435 37106 -4367
rect 28071 -4623 28139 -4555
rect 28191 -4623 28259 -4555
rect 35747 -4616 35815 -4548
rect 35867 -4616 35935 -4548
rect 45347 -4616 45415 -4548
rect 45467 -4616 45535 -4548
rect 25549 -4773 25615 -4708
rect 25682 -4773 25748 -4708
rect 28071 -4743 28139 -4675
rect 28191 -4743 28259 -4675
rect 35747 -4736 35815 -4668
rect 35867 -4736 35935 -4668
rect 45347 -4736 45415 -4668
rect 45467 -4736 45535 -4668
rect 25551 -4899 25617 -4834
rect 25683 -4897 25749 -4832
rect 26897 -4921 26965 -4853
rect 27017 -4921 27085 -4853
rect 30719 -4923 30787 -4855
rect 30839 -4923 30907 -4855
rect 36497 -4921 36565 -4853
rect 36617 -4921 36685 -4853
rect 26897 -5041 26965 -4973
rect 27017 -5041 27085 -4973
rect 30719 -5043 30787 -4975
rect 30839 -5043 30907 -4975
rect 36497 -5041 36565 -4973
rect 36617 -5041 36685 -4973
rect 33720 -5223 33788 -5155
rect 33840 -5223 33908 -5155
rect 35352 -5232 35420 -5164
rect 35472 -5232 35540 -5164
rect 44952 -5232 45020 -5164
rect 45072 -5232 45140 -5164
rect 33720 -5343 33788 -5275
rect 33840 -5343 33908 -5275
rect 35352 -5352 35420 -5284
rect 35472 -5352 35540 -5284
rect 44952 -5352 45020 -5284
rect 45072 -5352 45140 -5284
rect 28190 -5512 28258 -5444
rect 28310 -5512 28378 -5444
rect 37790 -5512 37858 -5444
rect 37910 -5512 37978 -5444
rect 28190 -5632 28258 -5564
rect 28310 -5632 28378 -5564
rect 37790 -5632 37858 -5564
rect 37910 -5632 37978 -5564
rect 34575 -5831 34643 -5763
rect 34695 -5831 34763 -5763
rect 39720 -5821 39788 -5753
rect 39840 -5821 39908 -5753
rect 44175 -5831 44243 -5763
rect 44295 -5831 44363 -5763
rect 34575 -5951 34643 -5883
rect 34695 -5951 34763 -5883
rect 39720 -5941 39788 -5873
rect 39840 -5941 39908 -5873
rect 44175 -5951 44243 -5883
rect 44295 -5951 44363 -5883
rect 27739 -6118 27807 -6050
rect 27859 -6118 27927 -6050
rect 37339 -6118 37407 -6050
rect 37459 -6118 37527 -6050
rect 42722 -6121 42790 -6053
rect 42842 -6121 42910 -6053
rect 27739 -6238 27807 -6170
rect 27859 -6238 27927 -6170
rect 37339 -6238 37407 -6170
rect 37459 -6238 37527 -6170
rect 42722 -6241 42790 -6173
rect 42842 -6241 42910 -6173
rect 25912 -6376 25978 -6311
rect 26045 -6376 26111 -6311
rect 25914 -6502 25980 -6437
rect 26046 -6500 26112 -6435
rect 34899 -6423 34967 -6355
rect 35019 -6423 35087 -6355
rect 44499 -6423 44567 -6355
rect 44619 -6423 44687 -6355
rect 34899 -6543 34967 -6475
rect 35019 -6543 35087 -6475
rect 44499 -6543 44567 -6475
rect 44619 -6543 44687 -6475
rect 28179 -6951 28247 -6883
rect 28299 -6951 28367 -6883
rect 26296 -7086 26362 -7021
rect 26429 -7086 26495 -7021
rect 26298 -7212 26364 -7147
rect 26430 -7210 26496 -7145
rect 27722 -7046 27790 -6978
rect 27842 -7046 27910 -6978
rect 37779 -6951 37847 -6883
rect 37899 -6951 37967 -6883
rect 28179 -7071 28247 -7003
rect 28299 -7071 28367 -7003
rect 34568 -7075 34636 -7007
rect 34688 -7075 34756 -7007
rect 27722 -7166 27790 -7098
rect 27842 -7166 27910 -7098
rect 34568 -7195 34636 -7127
rect 34688 -7195 34756 -7127
rect 34894 -7076 34962 -7008
rect 35014 -7076 35082 -7008
rect 34894 -7196 34962 -7128
rect 35014 -7196 35082 -7128
rect 37322 -7046 37390 -6978
rect 37442 -7046 37510 -6978
rect 37779 -7071 37847 -7003
rect 37899 -7071 37967 -7003
rect 44168 -7075 44236 -7007
rect 44288 -7075 44356 -7007
rect 37322 -7166 37390 -7098
rect 37442 -7166 37510 -7098
rect 44168 -7195 44236 -7127
rect 44288 -7195 44356 -7127
rect 44494 -7076 44562 -7008
rect 44614 -7076 44682 -7008
rect 44494 -7196 44562 -7128
rect 44614 -7196 44682 -7128
rect 9877 -7912 9945 -7844
rect 9997 -7912 10065 -7844
rect 9877 -8032 9945 -7964
rect 9997 -8032 10065 -7964
rect 19477 -7912 19545 -7844
rect 19597 -7912 19665 -7844
rect 19477 -8032 19545 -7964
rect 19597 -8032 19665 -7964
rect 26896 -7912 26964 -7844
rect 27016 -7912 27084 -7844
rect 26896 -8032 26964 -7964
rect 27016 -8032 27084 -7964
rect 36496 -7912 36564 -7844
rect 36616 -7912 36684 -7844
rect 36496 -8032 36564 -7964
rect 36616 -8032 36684 -7964
rect 1874 -8601 1942 -8533
rect 1994 -8601 2062 -8533
rect 1874 -8721 1942 -8653
rect 1994 -8721 2062 -8653
rect 11474 -8601 11542 -8533
rect 11594 -8601 11662 -8533
rect 11474 -8721 11542 -8653
rect 11594 -8721 11662 -8653
rect 34899 -8601 34967 -8533
rect 35019 -8601 35087 -8533
rect 34899 -8721 34967 -8653
rect 35019 -8721 35087 -8653
rect 44499 -8601 44567 -8533
rect 44619 -8601 44687 -8533
rect 44499 -8721 44567 -8653
rect 44619 -8721 44687 -8653
rect 2193 -9049 2261 -8981
rect 2313 -9049 2381 -8981
rect 2193 -9169 2261 -9101
rect 2313 -9169 2381 -9101
rect 9239 -9058 9307 -8990
rect 9359 -9058 9427 -8990
rect 9239 -9178 9307 -9110
rect 9359 -9178 9427 -9110
rect 11793 -9049 11861 -8981
rect 11913 -9049 11981 -8981
rect 11793 -9169 11861 -9101
rect 11913 -9169 11981 -9101
rect 18839 -9058 18907 -8990
rect 18959 -9058 19027 -8990
rect 18839 -9178 18907 -9110
rect 18959 -9178 19027 -9110
rect 27534 -9058 27602 -8990
rect 27654 -9058 27722 -8990
rect 27534 -9178 27602 -9110
rect 27654 -9178 27722 -9110
rect 34580 -9049 34648 -8981
rect 34700 -9049 34768 -8981
rect 34580 -9169 34648 -9101
rect 34700 -9169 34768 -9101
rect 37134 -9058 37202 -8990
rect 37254 -9058 37322 -8990
rect 37134 -9178 37202 -9110
rect 37254 -9178 37322 -9110
rect 44180 -9049 44248 -8981
rect 44300 -9049 44368 -8981
rect 44180 -9169 44248 -9101
rect 44300 -9169 44368 -9101
<< metal3 >>
rect 56897 12776 57520 13060
rect 23282 513 25053 797
rect 23282 -914 23566 513
rect 19686 -1198 23566 -914
rect 3649 -2332 3864 -2318
rect 3649 -2400 3663 -2332
rect 3731 -2400 3783 -2332
rect 3851 -2400 3864 -2332
rect 3649 -2452 3864 -2400
rect 3649 -2520 3663 -2452
rect 3731 -2520 3783 -2452
rect 3851 -2520 3864 -2452
rect 3649 -2533 3864 -2520
rect 6649 -2332 6864 -2318
rect 6649 -2400 6663 -2332
rect 6731 -2400 6783 -2332
rect 6851 -2400 6864 -2332
rect 6649 -2452 6864 -2400
rect 6649 -2520 6663 -2452
rect 6731 -2520 6783 -2452
rect 6851 -2520 6864 -2452
rect 6649 -2533 6864 -2520
rect 9649 -2332 9864 -2318
rect 9649 -2400 9663 -2332
rect 9731 -2400 9783 -2332
rect 9851 -2400 9864 -2332
rect 9649 -2452 9864 -2400
rect 9649 -2520 9663 -2452
rect 9731 -2520 9783 -2452
rect 9851 -2520 9864 -2452
rect 9649 -2533 9864 -2520
rect 12649 -2332 12864 -2318
rect 12649 -2400 12663 -2332
rect 12731 -2400 12783 -2332
rect 12851 -2400 12864 -2332
rect 12649 -2452 12864 -2400
rect 12649 -2520 12663 -2452
rect 12731 -2520 12783 -2452
rect 12851 -2520 12864 -2452
rect 12649 -2533 12864 -2520
rect 15649 -2332 15864 -2318
rect 15649 -2400 15663 -2332
rect 15731 -2400 15783 -2332
rect 15851 -2400 15864 -2332
rect 15649 -2452 15864 -2400
rect 15649 -2520 15663 -2452
rect 15731 -2520 15783 -2452
rect 15851 -2520 15864 -2452
rect 15649 -2533 15864 -2520
rect 18649 -2332 18864 -2318
rect 18649 -2400 18663 -2332
rect 18731 -2400 18783 -2332
rect 18851 -2400 18864 -2332
rect 18649 -2452 18864 -2400
rect 18649 -2520 18663 -2452
rect 18731 -2520 18783 -2452
rect 18851 -2520 18864 -2452
rect 18649 -2533 18864 -2520
rect 1012 -4548 1227 -4534
rect 1012 -4616 1026 -4548
rect 1094 -4616 1146 -4548
rect 1214 -4616 1227 -4548
rect 1012 -4668 1227 -4616
rect 1012 -4736 1026 -4668
rect 1094 -4736 1146 -4668
rect 1214 -4736 1227 -4668
rect 1012 -4749 1227 -4736
rect 1043 -8997 1204 -4749
rect 1407 -5164 1622 -5150
rect 1407 -5232 1421 -5164
rect 1489 -5232 1541 -5164
rect 1609 -5232 1622 -5164
rect 1407 -5284 1622 -5232
rect 1407 -5352 1421 -5284
rect 1489 -5352 1541 -5284
rect 1609 -5352 1622 -5284
rect 1407 -5365 1622 -5352
rect 1438 -8547 1598 -5365
rect 2184 -5763 2399 -5749
rect 2184 -5831 2198 -5763
rect 2266 -5831 2318 -5763
rect 2386 -5831 2399 -5763
rect 2184 -5883 2399 -5831
rect 2184 -5951 2198 -5883
rect 2266 -5951 2318 -5883
rect 2386 -5951 2399 -5883
rect 2184 -5964 2399 -5951
rect 1860 -6355 2075 -6341
rect 1860 -6423 1874 -6355
rect 1942 -6423 1994 -6355
rect 2062 -6423 2075 -6355
rect 1860 -6475 2075 -6423
rect 1860 -6543 1874 -6475
rect 1942 -6543 1994 -6475
rect 2062 -6543 2075 -6475
rect 1860 -6556 2075 -6543
rect 1888 -6994 2050 -6556
rect 2216 -6993 2378 -5964
rect 3672 -6039 3834 -2533
rect 6672 -5739 6834 -2533
rect 9672 -2732 9834 -2533
rect 8603 -2894 9834 -2732
rect 8603 -5430 8765 -2894
rect 9441 -4247 9656 -4233
rect 9441 -4315 9455 -4247
rect 9523 -4315 9575 -4247
rect 9643 -4315 9656 -4247
rect 9441 -4367 9656 -4315
rect 9441 -4435 9455 -4367
rect 9523 -4435 9575 -4367
rect 9643 -4435 9656 -4367
rect 9441 -4448 9656 -4435
rect 8569 -5444 8784 -5430
rect 8569 -5512 8583 -5444
rect 8651 -5512 8703 -5444
rect 8771 -5512 8784 -5444
rect 8569 -5564 8784 -5512
rect 8569 -5632 8583 -5564
rect 8651 -5632 8703 -5564
rect 8771 -5632 8784 -5564
rect 8569 -5645 8784 -5632
rect 6639 -5753 6854 -5739
rect 6639 -5821 6653 -5753
rect 6721 -5821 6773 -5753
rect 6841 -5821 6854 -5753
rect 6639 -5873 6854 -5821
rect 6639 -5941 6653 -5873
rect 6721 -5941 6773 -5873
rect 6841 -5941 6854 -5873
rect 6639 -5954 6854 -5941
rect 3637 -6053 3852 -6039
rect 3637 -6121 3651 -6053
rect 3719 -6121 3771 -6053
rect 3839 -6121 3852 -6053
rect 3637 -6173 3852 -6121
rect 3637 -6241 3651 -6173
rect 3719 -6241 3771 -6173
rect 3839 -6241 3852 -6173
rect 3637 -6254 3852 -6241
rect 8603 -6869 8765 -5645
rect 9020 -6050 9235 -6036
rect 9020 -6118 9034 -6050
rect 9102 -6118 9154 -6050
rect 9222 -6118 9235 -6050
rect 9020 -6170 9235 -6118
rect 9020 -6238 9034 -6170
rect 9102 -6238 9154 -6170
rect 9222 -6238 9235 -6170
rect 9020 -6251 9235 -6238
rect 8580 -6883 8795 -6869
rect 8580 -6951 8594 -6883
rect 8662 -6951 8714 -6883
rect 8782 -6951 8795 -6883
rect 1865 -7008 2080 -6994
rect 1865 -7076 1879 -7008
rect 1947 -7076 1999 -7008
rect 2067 -7076 2080 -7008
rect 1865 -7128 2080 -7076
rect 1865 -7196 1879 -7128
rect 1947 -7196 1999 -7128
rect 2067 -7196 2080 -7128
rect 1865 -7209 2080 -7196
rect 2191 -7007 2406 -6993
rect 2191 -7075 2205 -7007
rect 2273 -7075 2325 -7007
rect 2393 -7075 2406 -7007
rect 2191 -7127 2406 -7075
rect 8580 -7003 8795 -6951
rect 9064 -6964 9226 -6251
rect 8580 -7071 8594 -7003
rect 8662 -7071 8714 -7003
rect 8782 -7071 8795 -7003
rect 8580 -7084 8795 -7071
rect 9037 -6978 9252 -6964
rect 9037 -7046 9051 -6978
rect 9119 -7046 9171 -6978
rect 9239 -7046 9252 -6978
rect 2191 -7195 2205 -7127
rect 2273 -7195 2325 -7127
rect 2393 -7195 2406 -7127
rect 9037 -7098 9252 -7046
rect 9037 -7166 9051 -7098
rect 9119 -7166 9171 -7098
rect 9239 -7166 9252 -7098
rect 9037 -7179 9252 -7166
rect 2191 -7208 2406 -7195
rect 9470 -8149 9632 -4448
rect 10612 -4548 10827 -4534
rect 10612 -4616 10626 -4548
rect 10694 -4616 10746 -4548
rect 10814 -4616 10827 -4548
rect 10612 -4668 10827 -4616
rect 10612 -4736 10626 -4668
rect 10694 -4736 10746 -4668
rect 10814 -4736 10827 -4668
rect 10612 -4749 10827 -4736
rect 9862 -4853 10077 -4839
rect 9862 -4921 9876 -4853
rect 9944 -4921 9996 -4853
rect 10064 -4921 10077 -4853
rect 9862 -4973 10077 -4921
rect 9862 -5041 9876 -4973
rect 9944 -5041 9996 -4973
rect 10064 -5041 10077 -4973
rect 9862 -5054 10077 -5041
rect 9888 -7830 10050 -5054
rect 9863 -7844 10078 -7830
rect 9863 -7912 9877 -7844
rect 9945 -7912 9997 -7844
rect 10065 -7912 10078 -7844
rect 9863 -7964 10078 -7912
rect 9863 -8032 9877 -7964
rect 9945 -8032 9997 -7964
rect 10065 -8032 10078 -7964
rect 9863 -8045 10078 -8032
rect 9254 -8311 9632 -8149
rect 1860 -8533 2075 -8519
rect 1860 -8547 1874 -8533
rect 1438 -8601 1874 -8547
rect 1942 -8601 1994 -8533
rect 2062 -8601 2075 -8533
rect 1438 -8653 2075 -8601
rect 1438 -8707 1874 -8653
rect 1860 -8721 1874 -8707
rect 1942 -8721 1994 -8653
rect 2062 -8721 2075 -8653
rect 1860 -8734 2075 -8721
rect 2179 -8981 2394 -8967
rect 9254 -8976 9416 -8311
rect 2179 -8997 2193 -8981
rect 1043 -9049 2193 -8997
rect 2261 -9049 2313 -8981
rect 2381 -9049 2394 -8981
rect 1043 -9101 2394 -9049
rect 1043 -9158 2193 -9101
rect 2179 -9169 2193 -9158
rect 2261 -9169 2313 -9101
rect 2381 -9169 2394 -9101
rect 2179 -9182 2394 -9169
rect 9225 -8990 9440 -8976
rect 9225 -9058 9239 -8990
rect 9307 -9058 9359 -8990
rect 9427 -9058 9440 -8990
rect 9225 -9110 9440 -9058
rect 9225 -9178 9239 -9110
rect 9307 -9178 9359 -9110
rect 9427 -9178 9440 -9110
rect 10643 -8997 10804 -4749
rect 12672 -5141 12834 -2533
rect 15672 -4841 15834 -2533
rect 18672 -2732 18834 -2533
rect 18305 -2894 18834 -2732
rect 18305 -4541 18467 -2894
rect 19686 -4222 19970 -1198
rect 20320 -1933 20773 -1868
rect 20267 -1962 20819 -1933
rect 20267 -1965 20570 -1962
rect 20267 -2033 20313 -1965
rect 20381 -2033 20433 -1965
rect 20501 -2030 20570 -1965
rect 20638 -2030 20690 -1962
rect 20758 -2030 20819 -1962
rect 20501 -2033 20819 -2030
rect 20267 -2082 20819 -2033
rect 20267 -2085 20570 -2082
rect 20267 -2153 20313 -2085
rect 20381 -2153 20433 -2085
rect 20501 -2150 20570 -2085
rect 20638 -2150 20690 -2082
rect 20758 -2150 20819 -2082
rect 20501 -2153 20819 -2150
rect 20267 -2180 20819 -2153
rect 19038 -4247 20094 -4222
rect 19038 -4315 19055 -4247
rect 19123 -4315 19175 -4247
rect 19243 -4259 20094 -4247
rect 19243 -4292 20095 -4259
rect 19243 -4315 19331 -4292
rect 19038 -4360 19331 -4315
rect 19399 -4360 19451 -4292
rect 19519 -4293 20095 -4292
rect 19519 -4296 19887 -4293
rect 19519 -4360 19579 -4296
rect 19038 -4364 19579 -4360
rect 19647 -4364 19699 -4296
rect 19767 -4361 19887 -4296
rect 19955 -4361 20007 -4293
rect 20075 -4361 20095 -4293
rect 20320 -4328 20773 -2180
rect 27697 -2332 27912 -2318
rect 27697 -2400 27710 -2332
rect 27778 -2400 27830 -2332
rect 27898 -2400 27912 -2332
rect 27697 -2452 27912 -2400
rect 27697 -2520 27710 -2452
rect 27778 -2520 27830 -2452
rect 27898 -2520 27912 -2452
rect 27697 -2533 27912 -2520
rect 27727 -2732 27889 -2533
rect 26415 -2773 26797 -2745
rect 26415 -2829 26445 -2773
rect 26501 -2775 26797 -2773
rect 26501 -2829 26574 -2775
rect 26415 -2831 26574 -2829
rect 26630 -2778 26797 -2775
rect 26630 -2831 26713 -2778
rect 26415 -2834 26713 -2831
rect 26769 -2834 26797 -2778
rect 26415 -2861 26797 -2834
rect 25404 -3005 25786 -2977
rect 25404 -3061 25434 -3005
rect 25490 -3007 25786 -3005
rect 25490 -3061 25563 -3007
rect 25404 -3063 25563 -3061
rect 25619 -3010 25786 -3007
rect 25619 -3063 25702 -3010
rect 25404 -3066 25702 -3063
rect 25758 -3066 25786 -3010
rect 25404 -3093 25786 -3066
rect 23619 -3495 24001 -3467
rect 23619 -3551 23649 -3495
rect 23705 -3497 24001 -3495
rect 23705 -3551 23778 -3497
rect 23619 -3553 23778 -3551
rect 23834 -3500 24001 -3497
rect 23834 -3553 23917 -3500
rect 23619 -3556 23917 -3553
rect 23973 -3556 24001 -3500
rect 23619 -3583 24001 -3556
rect 23071 -3736 23419 -3715
rect 23071 -3792 23098 -3736
rect 23154 -3739 23419 -3736
rect 23154 -3792 23213 -3739
rect 23071 -3795 23213 -3792
rect 23269 -3795 23328 -3739
rect 23384 -3795 23419 -3739
rect 23071 -3811 23419 -3795
rect 23118 -4211 23305 -3811
rect 23098 -4229 23326 -4211
rect 23098 -4285 23126 -4229
rect 23182 -4230 23326 -4229
rect 23182 -4285 23244 -4230
rect 23098 -4286 23244 -4285
rect 23300 -4286 23326 -4230
rect 23098 -4303 23326 -4286
rect 19767 -4364 20095 -4361
rect 19038 -4367 20095 -4364
rect 19038 -4435 19055 -4367
rect 19123 -4435 19175 -4367
rect 19243 -4433 20095 -4367
rect 20309 -4347 20812 -4328
rect 20309 -4350 20607 -4347
rect 20309 -4418 20350 -4350
rect 20418 -4418 20470 -4350
rect 20538 -4415 20607 -4350
rect 20675 -4415 20727 -4347
rect 20795 -4415 20812 -4347
rect 20538 -4418 20812 -4415
rect 19243 -4435 20094 -4433
rect 19038 -4451 20094 -4435
rect 18288 -4555 18503 -4541
rect 18288 -4623 18302 -4555
rect 18370 -4623 18422 -4555
rect 18490 -4623 18503 -4555
rect 18288 -4675 18503 -4623
rect 18288 -4743 18302 -4675
rect 18370 -4743 18422 -4675
rect 18490 -4743 18503 -4675
rect 18288 -4756 18503 -4743
rect 15640 -4855 15855 -4841
rect 15640 -4923 15654 -4855
rect 15722 -4923 15774 -4855
rect 15842 -4923 15855 -4855
rect 15640 -4975 15855 -4923
rect 15640 -5043 15654 -4975
rect 15722 -5043 15774 -4975
rect 15842 -5043 15855 -4975
rect 15640 -5056 15855 -5043
rect 11007 -5164 11222 -5150
rect 11007 -5232 11021 -5164
rect 11089 -5232 11141 -5164
rect 11209 -5232 11222 -5164
rect 11007 -5284 11222 -5232
rect 11007 -5352 11021 -5284
rect 11089 -5352 11141 -5284
rect 11209 -5352 11222 -5284
rect 11007 -5365 11222 -5352
rect 12639 -5155 12854 -5141
rect 12639 -5223 12653 -5155
rect 12721 -5223 12773 -5155
rect 12841 -5223 12854 -5155
rect 12639 -5275 12854 -5223
rect 12639 -5343 12653 -5275
rect 12721 -5343 12773 -5275
rect 12841 -5343 12854 -5275
rect 12639 -5356 12854 -5343
rect 11038 -8547 11198 -5365
rect 18169 -5444 18384 -5430
rect 18169 -5512 18183 -5444
rect 18251 -5512 18303 -5444
rect 18371 -5512 18384 -5444
rect 18169 -5564 18384 -5512
rect 18169 -5632 18183 -5564
rect 18251 -5632 18303 -5564
rect 18371 -5632 18384 -5564
rect 18169 -5645 18384 -5632
rect 11784 -5763 11999 -5749
rect 11784 -5831 11798 -5763
rect 11866 -5831 11918 -5763
rect 11986 -5831 11999 -5763
rect 11784 -5883 11999 -5831
rect 11784 -5951 11798 -5883
rect 11866 -5951 11918 -5883
rect 11986 -5951 11999 -5883
rect 11784 -5964 11999 -5951
rect 11460 -6355 11675 -6341
rect 11460 -6423 11474 -6355
rect 11542 -6423 11594 -6355
rect 11662 -6423 11675 -6355
rect 11460 -6475 11675 -6423
rect 11460 -6543 11474 -6475
rect 11542 -6543 11594 -6475
rect 11662 -6543 11675 -6475
rect 11460 -6556 11675 -6543
rect 11488 -6994 11650 -6556
rect 11816 -6993 11978 -5964
rect 18203 -6869 18365 -5645
rect 18620 -6050 18835 -6036
rect 18620 -6118 18634 -6050
rect 18702 -6118 18754 -6050
rect 18822 -6118 18835 -6050
rect 18620 -6170 18835 -6118
rect 18620 -6238 18634 -6170
rect 18702 -6238 18754 -6170
rect 18822 -6238 18835 -6170
rect 18620 -6251 18835 -6238
rect 18180 -6883 18395 -6869
rect 18180 -6951 18194 -6883
rect 18262 -6951 18314 -6883
rect 18382 -6951 18395 -6883
rect 11465 -7008 11680 -6994
rect 11465 -7076 11479 -7008
rect 11547 -7076 11599 -7008
rect 11667 -7076 11680 -7008
rect 11465 -7128 11680 -7076
rect 11465 -7196 11479 -7128
rect 11547 -7196 11599 -7128
rect 11667 -7196 11680 -7128
rect 11465 -7209 11680 -7196
rect 11791 -7007 12006 -6993
rect 11791 -7075 11805 -7007
rect 11873 -7075 11925 -7007
rect 11993 -7075 12006 -7007
rect 11791 -7127 12006 -7075
rect 18180 -7003 18395 -6951
rect 18664 -6964 18826 -6251
rect 18180 -7071 18194 -7003
rect 18262 -7071 18314 -7003
rect 18382 -7071 18395 -7003
rect 18180 -7084 18395 -7071
rect 18637 -6978 18852 -6964
rect 18637 -7046 18651 -6978
rect 18719 -7046 18771 -6978
rect 18839 -7046 18852 -6978
rect 11791 -7195 11805 -7127
rect 11873 -7195 11925 -7127
rect 11993 -7195 12006 -7127
rect 18637 -7098 18852 -7046
rect 18637 -7166 18651 -7098
rect 18719 -7166 18771 -7098
rect 18839 -7166 18852 -7098
rect 18637 -7179 18852 -7166
rect 11791 -7208 12006 -7195
rect 19070 -8149 19232 -4451
rect 20309 -4467 20812 -4418
rect 23684 -4425 23870 -3583
rect 20309 -4470 20607 -4467
rect 20309 -4538 20350 -4470
rect 20418 -4538 20470 -4470
rect 20538 -4535 20607 -4470
rect 20675 -4535 20727 -4467
rect 20795 -4535 20812 -4467
rect 23659 -4449 23905 -4425
rect 23659 -4505 23686 -4449
rect 23742 -4450 23905 -4449
rect 23742 -4505 23820 -4450
rect 23659 -4506 23820 -4505
rect 23876 -4506 23905 -4450
rect 23659 -4524 23905 -4506
rect 20538 -4538 20812 -4535
rect 20309 -4567 20812 -4538
rect 25552 -4693 25738 -3093
rect 25875 -3256 26257 -3228
rect 25875 -3312 25905 -3256
rect 25961 -3258 26257 -3256
rect 25961 -3312 26034 -3258
rect 25875 -3314 26034 -3312
rect 26090 -3261 26257 -3258
rect 26090 -3314 26173 -3261
rect 25875 -3317 26173 -3314
rect 26229 -3317 26257 -3261
rect 25875 -3344 26257 -3317
rect 25524 -4708 25779 -4693
rect 25524 -4773 25549 -4708
rect 25615 -4773 25682 -4708
rect 25748 -4773 25779 -4708
rect 25524 -4832 25779 -4773
rect 25524 -4834 25683 -4832
rect 19462 -4853 19677 -4839
rect 19462 -4921 19476 -4853
rect 19544 -4921 19596 -4853
rect 19664 -4921 19677 -4853
rect 25524 -4899 25551 -4834
rect 25617 -4897 25683 -4834
rect 25749 -4897 25779 -4832
rect 25617 -4899 25779 -4897
rect 25524 -4914 25779 -4899
rect 19462 -4973 19677 -4921
rect 19462 -5041 19476 -4973
rect 19544 -5041 19596 -4973
rect 19664 -5041 19677 -4973
rect 19462 -5054 19677 -5041
rect 19488 -7830 19650 -5054
rect 25915 -6296 26101 -3344
rect 26550 -3650 26736 -2861
rect 27727 -2894 28256 -2732
rect 26304 -3836 26736 -3650
rect 25887 -6311 26142 -6296
rect 25887 -6376 25912 -6311
rect 25978 -6376 26045 -6311
rect 26111 -6376 26142 -6311
rect 25887 -6435 26142 -6376
rect 25887 -6437 26046 -6435
rect 25887 -6502 25914 -6437
rect 25980 -6500 26046 -6437
rect 26112 -6500 26142 -6435
rect 25980 -6502 26142 -6500
rect 25887 -6517 26142 -6502
rect 26304 -7006 26490 -3836
rect 27305 -4247 27520 -4233
rect 27305 -4315 27318 -4247
rect 27386 -4315 27438 -4247
rect 27506 -4315 27520 -4247
rect 27305 -4367 27520 -4315
rect 27305 -4435 27318 -4367
rect 27386 -4435 27438 -4367
rect 27506 -4435 27520 -4367
rect 27305 -4448 27520 -4435
rect 26884 -4853 27099 -4839
rect 26884 -4921 26897 -4853
rect 26965 -4921 27017 -4853
rect 27085 -4921 27099 -4853
rect 26884 -4973 27099 -4921
rect 26884 -5041 26897 -4973
rect 26965 -5041 27017 -4973
rect 27085 -5041 27099 -4973
rect 26884 -5054 27099 -5041
rect 26271 -7021 26526 -7006
rect 26271 -7086 26296 -7021
rect 26362 -7086 26429 -7021
rect 26495 -7086 26526 -7021
rect 26271 -7145 26526 -7086
rect 26271 -7147 26430 -7145
rect 26271 -7212 26298 -7147
rect 26364 -7210 26430 -7147
rect 26496 -7210 26526 -7145
rect 26364 -7212 26526 -7210
rect 26271 -7227 26526 -7212
rect 26911 -7830 27073 -5054
rect 19463 -7844 19678 -7830
rect 19463 -7912 19477 -7844
rect 19545 -7912 19597 -7844
rect 19665 -7912 19678 -7844
rect 19463 -7964 19678 -7912
rect 19463 -8032 19477 -7964
rect 19545 -8032 19597 -7964
rect 19665 -8032 19678 -7964
rect 19463 -8045 19678 -8032
rect 26883 -7844 27098 -7830
rect 26883 -7912 26896 -7844
rect 26964 -7912 27016 -7844
rect 27084 -7912 27098 -7844
rect 26883 -7964 27098 -7912
rect 26883 -8032 26896 -7964
rect 26964 -8032 27016 -7964
rect 27084 -8032 27098 -7964
rect 26883 -8045 27098 -8032
rect 18854 -8311 19232 -8149
rect 27329 -8149 27491 -4448
rect 28094 -4541 28256 -2894
rect 29940 -4257 30224 396
rect 30697 -2332 30912 -2318
rect 30697 -2400 30710 -2332
rect 30778 -2400 30830 -2332
rect 30898 -2400 30912 -2332
rect 30697 -2452 30912 -2400
rect 30697 -2520 30710 -2452
rect 30778 -2520 30830 -2452
rect 30898 -2520 30912 -2452
rect 30697 -2533 30912 -2520
rect 33697 -2332 33912 -2318
rect 33697 -2400 33710 -2332
rect 33778 -2400 33830 -2332
rect 33898 -2400 33912 -2332
rect 33697 -2452 33912 -2400
rect 33697 -2520 33710 -2452
rect 33778 -2520 33830 -2452
rect 33898 -2520 33912 -2452
rect 33697 -2533 33912 -2520
rect 36697 -2332 36912 -2318
rect 36697 -2400 36710 -2332
rect 36778 -2400 36830 -2332
rect 36898 -2400 36912 -2332
rect 36697 -2452 36912 -2400
rect 36697 -2520 36710 -2452
rect 36778 -2520 36830 -2452
rect 36898 -2520 36912 -2452
rect 36697 -2533 36912 -2520
rect 39697 -2332 39912 -2318
rect 39697 -2400 39710 -2332
rect 39778 -2400 39830 -2332
rect 39898 -2400 39912 -2332
rect 39697 -2452 39912 -2400
rect 39697 -2520 39710 -2452
rect 39778 -2520 39830 -2452
rect 39898 -2520 39912 -2452
rect 39697 -2533 39912 -2520
rect 42697 -2332 42912 -2318
rect 42697 -2400 42710 -2332
rect 42778 -2400 42830 -2332
rect 42898 -2400 42912 -2332
rect 42697 -2452 42912 -2400
rect 42697 -2520 42710 -2452
rect 42778 -2520 42830 -2452
rect 42898 -2520 42912 -2452
rect 42697 -2533 42912 -2520
rect 29497 -4291 30383 -4257
rect 29497 -4294 29847 -4291
rect 29497 -4362 29539 -4294
rect 29607 -4362 29659 -4294
rect 29727 -4359 29847 -4294
rect 29915 -4359 29967 -4291
rect 30035 -4293 30383 -4291
rect 30035 -4359 30138 -4293
rect 29727 -4361 30138 -4359
rect 30206 -4361 30258 -4293
rect 30326 -4361 30383 -4293
rect 29727 -4362 30383 -4361
rect 29497 -4431 30383 -4362
rect 28058 -4555 28273 -4541
rect 28058 -4623 28071 -4555
rect 28139 -4623 28191 -4555
rect 28259 -4623 28273 -4555
rect 28058 -4675 28273 -4623
rect 28058 -4743 28071 -4675
rect 28139 -4743 28191 -4675
rect 28259 -4743 28273 -4675
rect 28058 -4756 28273 -4743
rect 30727 -4841 30889 -2533
rect 30706 -4855 30921 -4841
rect 30706 -4923 30719 -4855
rect 30787 -4923 30839 -4855
rect 30907 -4923 30921 -4855
rect 30706 -4975 30921 -4923
rect 30706 -5043 30719 -4975
rect 30787 -5043 30839 -4975
rect 30907 -5043 30921 -4975
rect 30706 -5056 30921 -5043
rect 33727 -5141 33889 -2533
rect 36727 -2732 36889 -2533
rect 36727 -2894 37958 -2732
rect 36905 -4247 37120 -4233
rect 36905 -4315 36918 -4247
rect 36986 -4315 37038 -4247
rect 37106 -4315 37120 -4247
rect 36905 -4367 37120 -4315
rect 36905 -4435 36918 -4367
rect 36986 -4435 37038 -4367
rect 37106 -4435 37120 -4367
rect 36905 -4448 37120 -4435
rect 35734 -4548 35949 -4534
rect 35734 -4616 35747 -4548
rect 35815 -4616 35867 -4548
rect 35935 -4616 35949 -4548
rect 35734 -4668 35949 -4616
rect 35734 -4736 35747 -4668
rect 35815 -4736 35867 -4668
rect 35935 -4736 35949 -4668
rect 35734 -4749 35949 -4736
rect 33707 -5155 33922 -5141
rect 33707 -5223 33720 -5155
rect 33788 -5223 33840 -5155
rect 33908 -5223 33922 -5155
rect 33707 -5275 33922 -5223
rect 33707 -5343 33720 -5275
rect 33788 -5343 33840 -5275
rect 33908 -5343 33922 -5275
rect 33707 -5356 33922 -5343
rect 35339 -5164 35554 -5150
rect 35339 -5232 35352 -5164
rect 35420 -5232 35472 -5164
rect 35540 -5232 35554 -5164
rect 35339 -5284 35554 -5232
rect 35339 -5352 35352 -5284
rect 35420 -5352 35472 -5284
rect 35540 -5352 35554 -5284
rect 35339 -5365 35554 -5352
rect 28177 -5444 28392 -5430
rect 28177 -5512 28190 -5444
rect 28258 -5512 28310 -5444
rect 28378 -5512 28392 -5444
rect 28177 -5564 28392 -5512
rect 28177 -5632 28190 -5564
rect 28258 -5632 28310 -5564
rect 28378 -5632 28392 -5564
rect 28177 -5645 28392 -5632
rect 27726 -6050 27941 -6036
rect 27726 -6118 27739 -6050
rect 27807 -6118 27859 -6050
rect 27927 -6118 27941 -6050
rect 27726 -6170 27941 -6118
rect 27726 -6238 27739 -6170
rect 27807 -6238 27859 -6170
rect 27927 -6238 27941 -6170
rect 27726 -6251 27941 -6238
rect 27735 -6964 27897 -6251
rect 28196 -6869 28358 -5645
rect 34562 -5763 34777 -5749
rect 34562 -5831 34575 -5763
rect 34643 -5831 34695 -5763
rect 34763 -5831 34777 -5763
rect 34562 -5883 34777 -5831
rect 34562 -5951 34575 -5883
rect 34643 -5951 34695 -5883
rect 34763 -5951 34777 -5883
rect 34562 -5964 34777 -5951
rect 28166 -6883 28381 -6869
rect 28166 -6951 28179 -6883
rect 28247 -6951 28299 -6883
rect 28367 -6951 28381 -6883
rect 27709 -6978 27924 -6964
rect 27709 -7046 27722 -6978
rect 27790 -7046 27842 -6978
rect 27910 -7046 27924 -6978
rect 27709 -7098 27924 -7046
rect 28166 -7003 28381 -6951
rect 34583 -6993 34745 -5964
rect 34886 -6355 35101 -6341
rect 34886 -6423 34899 -6355
rect 34967 -6423 35019 -6355
rect 35087 -6423 35101 -6355
rect 34886 -6475 35101 -6423
rect 34886 -6543 34899 -6475
rect 34967 -6543 35019 -6475
rect 35087 -6543 35101 -6475
rect 34886 -6556 35101 -6543
rect 28166 -7071 28179 -7003
rect 28247 -7071 28299 -7003
rect 28367 -7071 28381 -7003
rect 28166 -7084 28381 -7071
rect 34555 -7007 34770 -6993
rect 34911 -6994 35073 -6556
rect 34555 -7075 34568 -7007
rect 34636 -7075 34688 -7007
rect 34756 -7075 34770 -7007
rect 27709 -7166 27722 -7098
rect 27790 -7166 27842 -7098
rect 27910 -7166 27924 -7098
rect 27709 -7179 27924 -7166
rect 34555 -7127 34770 -7075
rect 34555 -7195 34568 -7127
rect 34636 -7195 34688 -7127
rect 34756 -7195 34770 -7127
rect 34555 -7208 34770 -7195
rect 34881 -7008 35096 -6994
rect 34881 -7076 34894 -7008
rect 34962 -7076 35014 -7008
rect 35082 -7076 35096 -7008
rect 34881 -7128 35096 -7076
rect 34881 -7196 34894 -7128
rect 34962 -7196 35014 -7128
rect 35082 -7196 35096 -7128
rect 34881 -7209 35096 -7196
rect 27329 -8311 27707 -8149
rect 11460 -8533 11675 -8519
rect 11460 -8547 11474 -8533
rect 11038 -8601 11474 -8547
rect 11542 -8601 11594 -8533
rect 11662 -8601 11675 -8533
rect 11038 -8653 11675 -8601
rect 11038 -8707 11474 -8653
rect 11460 -8721 11474 -8707
rect 11542 -8721 11594 -8653
rect 11662 -8721 11675 -8653
rect 11460 -8734 11675 -8721
rect 11779 -8981 11994 -8967
rect 18854 -8976 19016 -8311
rect 27545 -8976 27707 -8311
rect 34886 -8533 35101 -8519
rect 34886 -8601 34899 -8533
rect 34967 -8601 35019 -8533
rect 35087 -8547 35101 -8533
rect 35363 -8547 35523 -5365
rect 35087 -8601 35523 -8547
rect 34886 -8653 35523 -8601
rect 34886 -8721 34899 -8653
rect 34967 -8721 35019 -8653
rect 35087 -8707 35523 -8653
rect 35087 -8721 35101 -8707
rect 34886 -8734 35101 -8721
rect 11779 -8997 11793 -8981
rect 10643 -9049 11793 -8997
rect 11861 -9049 11913 -8981
rect 11981 -9049 11994 -8981
rect 10643 -9101 11994 -9049
rect 10643 -9158 11793 -9101
rect 9225 -9191 9440 -9178
rect 11779 -9169 11793 -9158
rect 11861 -9169 11913 -9101
rect 11981 -9169 11994 -9101
rect 11779 -9182 11994 -9169
rect 18825 -8990 19040 -8976
rect 18825 -9058 18839 -8990
rect 18907 -9058 18959 -8990
rect 19027 -9058 19040 -8990
rect 18825 -9110 19040 -9058
rect 18825 -9178 18839 -9110
rect 18907 -9178 18959 -9110
rect 19027 -9178 19040 -9110
rect 18825 -9191 19040 -9178
rect 27521 -8990 27736 -8976
rect 27521 -9058 27534 -8990
rect 27602 -9058 27654 -8990
rect 27722 -9058 27736 -8990
rect 27521 -9110 27736 -9058
rect 27521 -9178 27534 -9110
rect 27602 -9178 27654 -9110
rect 27722 -9178 27736 -9110
rect 27521 -9191 27736 -9178
rect 34567 -8981 34782 -8967
rect 34567 -9049 34580 -8981
rect 34648 -9049 34700 -8981
rect 34768 -8997 34782 -8981
rect 35757 -8997 35918 -4749
rect 36484 -4853 36699 -4839
rect 36484 -4921 36497 -4853
rect 36565 -4921 36617 -4853
rect 36685 -4921 36699 -4853
rect 36484 -4973 36699 -4921
rect 36484 -5041 36497 -4973
rect 36565 -5041 36617 -4973
rect 36685 -5041 36699 -4973
rect 36484 -5054 36699 -5041
rect 36511 -7830 36673 -5054
rect 36483 -7844 36698 -7830
rect 36483 -7912 36496 -7844
rect 36564 -7912 36616 -7844
rect 36684 -7912 36698 -7844
rect 36483 -7964 36698 -7912
rect 36483 -8032 36496 -7964
rect 36564 -8032 36616 -7964
rect 36684 -8032 36698 -7964
rect 36483 -8045 36698 -8032
rect 36929 -8149 37091 -4448
rect 37796 -5430 37958 -2894
rect 37777 -5444 37992 -5430
rect 37777 -5512 37790 -5444
rect 37858 -5512 37910 -5444
rect 37978 -5512 37992 -5444
rect 37777 -5564 37992 -5512
rect 37777 -5632 37790 -5564
rect 37858 -5632 37910 -5564
rect 37978 -5632 37992 -5564
rect 37777 -5645 37992 -5632
rect 37326 -6050 37541 -6036
rect 37326 -6118 37339 -6050
rect 37407 -6118 37459 -6050
rect 37527 -6118 37541 -6050
rect 37326 -6170 37541 -6118
rect 37326 -6238 37339 -6170
rect 37407 -6238 37459 -6170
rect 37527 -6238 37541 -6170
rect 37326 -6251 37541 -6238
rect 37335 -6964 37497 -6251
rect 37796 -6869 37958 -5645
rect 39727 -5739 39889 -2533
rect 39707 -5753 39922 -5739
rect 39707 -5821 39720 -5753
rect 39788 -5821 39840 -5753
rect 39908 -5821 39922 -5753
rect 39707 -5873 39922 -5821
rect 39707 -5941 39720 -5873
rect 39788 -5941 39840 -5873
rect 39908 -5941 39922 -5873
rect 39707 -5954 39922 -5941
rect 42727 -6039 42889 -2533
rect 45334 -4548 45549 -4534
rect 45334 -4616 45347 -4548
rect 45415 -4616 45467 -4548
rect 45535 -4616 45549 -4548
rect 45334 -4668 45549 -4616
rect 45334 -4736 45347 -4668
rect 45415 -4736 45467 -4668
rect 45535 -4736 45549 -4668
rect 45334 -4749 45549 -4736
rect 44939 -5164 45154 -5150
rect 44939 -5232 44952 -5164
rect 45020 -5232 45072 -5164
rect 45140 -5232 45154 -5164
rect 44939 -5284 45154 -5232
rect 44939 -5352 44952 -5284
rect 45020 -5352 45072 -5284
rect 45140 -5352 45154 -5284
rect 44939 -5365 45154 -5352
rect 44162 -5763 44377 -5749
rect 44162 -5831 44175 -5763
rect 44243 -5831 44295 -5763
rect 44363 -5831 44377 -5763
rect 44162 -5883 44377 -5831
rect 44162 -5951 44175 -5883
rect 44243 -5951 44295 -5883
rect 44363 -5951 44377 -5883
rect 44162 -5964 44377 -5951
rect 42709 -6053 42924 -6039
rect 42709 -6121 42722 -6053
rect 42790 -6121 42842 -6053
rect 42910 -6121 42924 -6053
rect 42709 -6173 42924 -6121
rect 42709 -6241 42722 -6173
rect 42790 -6241 42842 -6173
rect 42910 -6241 42924 -6173
rect 42709 -6254 42924 -6241
rect 37766 -6883 37981 -6869
rect 37766 -6951 37779 -6883
rect 37847 -6951 37899 -6883
rect 37967 -6951 37981 -6883
rect 37309 -6978 37524 -6964
rect 37309 -7046 37322 -6978
rect 37390 -7046 37442 -6978
rect 37510 -7046 37524 -6978
rect 37309 -7098 37524 -7046
rect 37766 -7003 37981 -6951
rect 44183 -6993 44345 -5964
rect 44486 -6355 44701 -6341
rect 44486 -6423 44499 -6355
rect 44567 -6423 44619 -6355
rect 44687 -6423 44701 -6355
rect 44486 -6475 44701 -6423
rect 44486 -6543 44499 -6475
rect 44567 -6543 44619 -6475
rect 44687 -6543 44701 -6475
rect 44486 -6556 44701 -6543
rect 37766 -7071 37779 -7003
rect 37847 -7071 37899 -7003
rect 37967 -7071 37981 -7003
rect 37766 -7084 37981 -7071
rect 44155 -7007 44370 -6993
rect 44511 -6994 44673 -6556
rect 44155 -7075 44168 -7007
rect 44236 -7075 44288 -7007
rect 44356 -7075 44370 -7007
rect 37309 -7166 37322 -7098
rect 37390 -7166 37442 -7098
rect 37510 -7166 37524 -7098
rect 37309 -7179 37524 -7166
rect 44155 -7127 44370 -7075
rect 44155 -7195 44168 -7127
rect 44236 -7195 44288 -7127
rect 44356 -7195 44370 -7127
rect 44155 -7208 44370 -7195
rect 44481 -7008 44696 -6994
rect 44481 -7076 44494 -7008
rect 44562 -7076 44614 -7008
rect 44682 -7076 44696 -7008
rect 44481 -7128 44696 -7076
rect 44481 -7196 44494 -7128
rect 44562 -7196 44614 -7128
rect 44682 -7196 44696 -7128
rect 44481 -7209 44696 -7196
rect 36929 -8311 37307 -8149
rect 37145 -8976 37307 -8311
rect 44486 -8533 44701 -8519
rect 44486 -8601 44499 -8533
rect 44567 -8601 44619 -8533
rect 44687 -8547 44701 -8533
rect 44963 -8547 45123 -5365
rect 44687 -8601 45123 -8547
rect 44486 -8653 45123 -8601
rect 44486 -8721 44499 -8653
rect 44567 -8721 44619 -8653
rect 44687 -8707 45123 -8653
rect 44687 -8721 44701 -8707
rect 44486 -8734 44701 -8721
rect 34768 -9049 35918 -8997
rect 34567 -9101 35918 -9049
rect 34567 -9169 34580 -9101
rect 34648 -9169 34700 -9101
rect 34768 -9158 35918 -9101
rect 37121 -8990 37336 -8976
rect 37121 -9058 37134 -8990
rect 37202 -9058 37254 -8990
rect 37322 -9058 37336 -8990
rect 37121 -9110 37336 -9058
rect 34768 -9169 34782 -9158
rect 34567 -9182 34782 -9169
rect 37121 -9178 37134 -9110
rect 37202 -9178 37254 -9110
rect 37322 -9178 37336 -9110
rect 37121 -9191 37336 -9178
rect 44167 -8981 44382 -8967
rect 44167 -9049 44180 -8981
rect 44248 -9049 44300 -8981
rect 44368 -8997 44382 -8981
rect 45357 -8997 45518 -4749
rect 44368 -9049 45518 -8997
rect 44167 -9101 45518 -9049
rect 44167 -9169 44180 -9101
rect 44248 -9169 44300 -9101
rect 44368 -9158 45518 -9101
rect 44368 -9169 44382 -9158
rect 44167 -9182 44382 -9169
use Folded_Diff_Op_Amp_Layout  Folded_Diff_Op_Amp_Layout_0 ~/GF180Projects/Tapeout/Magic/Op_Amp
timestamp 1699898304
transform 1 0 486 0 1 9157
box -486 -9157 66932 6239
use PGA_Dec_Layout  PGA_Dec_Layout_0 ~/GF180Projects/Tapeout/Magic/PGA_Decoder
timestamp 1699521709
transform 1 0 20565 0 1 -5932
box -99 -2026 5362 1565
use resistor_PGA_new  resistor_PGA_new_2 ~/GF180Projects/Tapeout/Magic/Resistor_divider
timestamp 1694518401
transform 1 0 -4292 0 1 -22418
box 5446 12554 14427 15705
use resistor_PGA_new  resistor_PGA_new_3
timestamp 1694518401
transform 1 0 5308 0 1 -22418
box 5446 12554 14427 15705
use resistor_PGA_new  resistor_PGA_new_4
timestamp 1694518401
transform -1 0 50853 0 1 -22418
box 5446 12554 14427 15705
use resistor_PGA_new  resistor_PGA_new_5
timestamp 1694518401
transform -1 0 41253 0 1 -22418
box 5446 12554 14427 15705
use TG_5x_Layout  TG_5x_Layout_6 ~/GF180Projects/Tapeout/Magic/Logic_Gates/5x_TG
timestamp 1699521709
transform 1 0 2107 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_7
timestamp 1699521709
transform 1 0 17107 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_8
timestamp 1699521709
transform 1 0 5107 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_9
timestamp 1699521709
transform 1 0 8107 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_10
timestamp 1699521709
transform 1 0 11107 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_11
timestamp 1699521709
transform 1 0 14107 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_12
timestamp 1699521709
transform -1 0 38454 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_13
timestamp 1699521709
transform -1 0 41454 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_14
timestamp 1699521709
transform -1 0 44454 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_15
timestamp 1699521709
transform -1 0 32454 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_16
timestamp 1699521709
transform -1 0 35454 0 1 -2600
box -112 -27 1482 953
use TG_5x_Layout  TG_5x_Layout_17
timestamp 1699521709
transform -1 0 29454 0 1 -2600
box -112 -27 1482 953
<< labels >>
flabel metal2 14231 -6149 14231 -6149 0 FreeSans 480 0 0 0 B1
port 9 nsew
flabel metal2 14398 -5857 14398 -5857 0 FreeSans 480 0 0 0 C1
port 10 nsew
flabel metal2 14174 -5561 14174 -5561 0 FreeSans 480 0 0 0 D1
port 11 nsew
flabel metal2 13981 -5254 13981 -5254 0 FreeSans 480 0 0 0 E1
port 12 nsew
flabel metal2 14288 -4958 14288 -4958 0 FreeSans 480 0 0 0 F1
port 13 nsew
flabel metal2 14131 -4676 14131 -4676 0 FreeSans 480 0 0 0 G1
port 14 nsew
flabel metal2 14145 -4352 14145 -4352 0 FreeSans 480 0 0 0 H1
port 15 nsew
flabel metal2 29482 -6170 29482 -6170 0 FreeSans 480 0 0 0 B2
port 17 nsew
flabel metal2 29650 -5860 29650 -5860 0 FreeSans 480 0 0 0 C2
port 18 nsew
flabel metal2 29422 -5568 29422 -5568 0 FreeSans 480 0 0 0 D2
port 19 nsew
flabel metal2 29183 -5272 29183 -5272 0 FreeSans 480 0 0 0 E2
port 20 nsew
flabel metal2 29568 -4965 29568 -4965 0 FreeSans 480 0 0 0 F2
port 21 nsew
flabel metal2 29272 -4673 29272 -4673 0 FreeSans 480 0 0 0 G2
port 22 nsew
flabel metal2 29614 -4334 29614 -4334 0 FreeSans 480 0 0 0 H2
port 23 nsew
flabel metal2 22511 -4008 22511 -4008 0 FreeSans 800 0 0 0 SS6
port 53 nsew
flabel metal2 22492 -3762 22492 -3762 0 FreeSans 800 0 0 0 SS5
port 54 nsew
flabel metal2 22492 -3524 22492 -3524 0 FreeSans 800 0 0 0 SS4
port 55 nsew
flabel metal2 22487 -3283 22487 -3283 0 FreeSans 800 0 0 0 SS3
port 56 nsew
flabel metal2 22476 -3049 22476 -3049 0 FreeSans 800 0 0 0 SS2
port 57 nsew
flabel metal2 22459 -2809 22459 -2809 0 FreeSans 800 0 0 0 SS1
port 58 nsew
flabel metal1 22811 -10288 22811 -10288 0 FreeSans 1600 0 0 0 VDD
port 59 nsew
flabel metal1 20705 -7967 20705 -7967 0 FreeSans 1600 0 0 0 VSS
port 60 nsew
flabel metal3 57212 12906 57212 12906 0 FreeSans 1600 0 0 0 IBS2
port 61 nsew
flabel metal2 44 14788 44 14788 0 FreeSans 1600 0 0 0 INN
port 64 nsew
flabel metal2 102 13097 102 13097 0 FreeSans 1600 0 0 0 INP
port 65 nsew
flabel metal2 2598 13608 2602 13608 0 FreeSans 1600 0 0 0 BD1
port 66 nsew
flabel metal1 -318 7493 -318 7493 0 FreeSans 1600 0 0 0 IBS
port 67 nsew
flabel space 31345 14870 31345 14870 0 FreeSans 1600 0 0 0 OUTP
port 70 nsew
flabel space 32240 14562 32240 14562 0 FreeSans 1600 0 0 0 OUTN
port 71 nsew
flabel metal2 -315 -6453 -315 -6453 0 FreeSans 1600 0 0 0 IN1
port 72 nsew
flabel metal2 46613 -6456 46613 -6456 0 FreeSans 1600 0 0 0 IN2
port 73 nsew
<< end >>
