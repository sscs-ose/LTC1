magic
tech gf180mcuC
magscale 1 10
timestamp 1695274000
<< mimcap >>
rect -1720 1440 1480 1520
rect -1720 -1440 -1640 1440
rect 1400 -1440 1480 1440
rect -1720 -1520 1480 -1440
<< mimcapcontact >>
rect -1640 -1440 1400 1440
<< metal4 >>
rect -1840 1573 1840 1640
rect -1840 1520 1690 1573
rect -1840 -1520 -1720 1520
rect 1480 -1520 1690 1520
rect -1840 -1573 1690 -1520
rect 1778 -1573 1840 1573
rect -1840 -1640 1840 -1573
<< via4 >>
rect 1690 -1573 1778 1573
<< metal5 >>
rect 1690 1573 1778 1583
rect 1690 -1583 1778 -1573
<< properties >>
string FIXED_BBOX -1840 -1640 1600 1640
string gencell cap_mim_2p0fF
string library gf180mcu
string parameters w 16 l 15.2 val 7.328k carea 25.00 cperi 20.00 nx 1 ny 1 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 1 tconnect 1
<< end >>
