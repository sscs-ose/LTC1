magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1316 -1316 1316 1316
<< metal1 >>
rect -316 310 316 316
rect -316 284 -310 310
rect -284 284 -244 310
rect -218 284 -178 310
rect -152 284 -112 310
rect -86 284 -46 310
rect -20 284 20 310
rect 46 284 86 310
rect 112 284 152 310
rect 178 284 218 310
rect 244 284 284 310
rect 310 284 316 310
rect -316 244 316 284
rect -316 218 -310 244
rect -284 218 -244 244
rect -218 218 -178 244
rect -152 218 -112 244
rect -86 218 -46 244
rect -20 218 20 244
rect 46 218 86 244
rect 112 218 152 244
rect 178 218 218 244
rect 244 218 284 244
rect 310 218 316 244
rect -316 178 316 218
rect -316 152 -310 178
rect -284 152 -244 178
rect -218 152 -178 178
rect -152 152 -112 178
rect -86 152 -46 178
rect -20 152 20 178
rect 46 152 86 178
rect 112 152 152 178
rect 178 152 218 178
rect 244 152 284 178
rect 310 152 316 178
rect -316 112 316 152
rect -316 86 -310 112
rect -284 86 -244 112
rect -218 86 -178 112
rect -152 86 -112 112
rect -86 86 -46 112
rect -20 86 20 112
rect 46 86 86 112
rect 112 86 152 112
rect 178 86 218 112
rect 244 86 284 112
rect 310 86 316 112
rect -316 46 316 86
rect -316 20 -310 46
rect -284 20 -244 46
rect -218 20 -178 46
rect -152 20 -112 46
rect -86 20 -46 46
rect -20 20 20 46
rect 46 20 86 46
rect 112 20 152 46
rect 178 20 218 46
rect 244 20 284 46
rect 310 20 316 46
rect -316 -20 316 20
rect -316 -46 -310 -20
rect -284 -46 -244 -20
rect -218 -46 -178 -20
rect -152 -46 -112 -20
rect -86 -46 -46 -20
rect -20 -46 20 -20
rect 46 -46 86 -20
rect 112 -46 152 -20
rect 178 -46 218 -20
rect 244 -46 284 -20
rect 310 -46 316 -20
rect -316 -86 316 -46
rect -316 -112 -310 -86
rect -284 -112 -244 -86
rect -218 -112 -178 -86
rect -152 -112 -112 -86
rect -86 -112 -46 -86
rect -20 -112 20 -86
rect 46 -112 86 -86
rect 112 -112 152 -86
rect 178 -112 218 -86
rect 244 -112 284 -86
rect 310 -112 316 -86
rect -316 -152 316 -112
rect -316 -178 -310 -152
rect -284 -178 -244 -152
rect -218 -178 -178 -152
rect -152 -178 -112 -152
rect -86 -178 -46 -152
rect -20 -178 20 -152
rect 46 -178 86 -152
rect 112 -178 152 -152
rect 178 -178 218 -152
rect 244 -178 284 -152
rect 310 -178 316 -152
rect -316 -218 316 -178
rect -316 -244 -310 -218
rect -284 -244 -244 -218
rect -218 -244 -178 -218
rect -152 -244 -112 -218
rect -86 -244 -46 -218
rect -20 -244 20 -218
rect 46 -244 86 -218
rect 112 -244 152 -218
rect 178 -244 218 -218
rect 244 -244 284 -218
rect 310 -244 316 -218
rect -316 -284 316 -244
rect -316 -310 -310 -284
rect -284 -310 -244 -284
rect -218 -310 -178 -284
rect -152 -310 -112 -284
rect -86 -310 -46 -284
rect -20 -310 20 -284
rect 46 -310 86 -284
rect 112 -310 152 -284
rect 178 -310 218 -284
rect 244 -310 284 -284
rect 310 -310 316 -284
rect -316 -316 316 -310
<< via1 >>
rect -310 284 -284 310
rect -244 284 -218 310
rect -178 284 -152 310
rect -112 284 -86 310
rect -46 284 -20 310
rect 20 284 46 310
rect 86 284 112 310
rect 152 284 178 310
rect 218 284 244 310
rect 284 284 310 310
rect -310 218 -284 244
rect -244 218 -218 244
rect -178 218 -152 244
rect -112 218 -86 244
rect -46 218 -20 244
rect 20 218 46 244
rect 86 218 112 244
rect 152 218 178 244
rect 218 218 244 244
rect 284 218 310 244
rect -310 152 -284 178
rect -244 152 -218 178
rect -178 152 -152 178
rect -112 152 -86 178
rect -46 152 -20 178
rect 20 152 46 178
rect 86 152 112 178
rect 152 152 178 178
rect 218 152 244 178
rect 284 152 310 178
rect -310 86 -284 112
rect -244 86 -218 112
rect -178 86 -152 112
rect -112 86 -86 112
rect -46 86 -20 112
rect 20 86 46 112
rect 86 86 112 112
rect 152 86 178 112
rect 218 86 244 112
rect 284 86 310 112
rect -310 20 -284 46
rect -244 20 -218 46
rect -178 20 -152 46
rect -112 20 -86 46
rect -46 20 -20 46
rect 20 20 46 46
rect 86 20 112 46
rect 152 20 178 46
rect 218 20 244 46
rect 284 20 310 46
rect -310 -46 -284 -20
rect -244 -46 -218 -20
rect -178 -46 -152 -20
rect -112 -46 -86 -20
rect -46 -46 -20 -20
rect 20 -46 46 -20
rect 86 -46 112 -20
rect 152 -46 178 -20
rect 218 -46 244 -20
rect 284 -46 310 -20
rect -310 -112 -284 -86
rect -244 -112 -218 -86
rect -178 -112 -152 -86
rect -112 -112 -86 -86
rect -46 -112 -20 -86
rect 20 -112 46 -86
rect 86 -112 112 -86
rect 152 -112 178 -86
rect 218 -112 244 -86
rect 284 -112 310 -86
rect -310 -178 -284 -152
rect -244 -178 -218 -152
rect -178 -178 -152 -152
rect -112 -178 -86 -152
rect -46 -178 -20 -152
rect 20 -178 46 -152
rect 86 -178 112 -152
rect 152 -178 178 -152
rect 218 -178 244 -152
rect 284 -178 310 -152
rect -310 -244 -284 -218
rect -244 -244 -218 -218
rect -178 -244 -152 -218
rect -112 -244 -86 -218
rect -46 -244 -20 -218
rect 20 -244 46 -218
rect 86 -244 112 -218
rect 152 -244 178 -218
rect 218 -244 244 -218
rect 284 -244 310 -218
rect -310 -310 -284 -284
rect -244 -310 -218 -284
rect -178 -310 -152 -284
rect -112 -310 -86 -284
rect -46 -310 -20 -284
rect 20 -310 46 -284
rect 86 -310 112 -284
rect 152 -310 178 -284
rect 218 -310 244 -284
rect 284 -310 310 -284
<< metal2 >>
rect -316 310 316 316
rect -316 284 -310 310
rect -284 284 -244 310
rect -218 284 -178 310
rect -152 284 -112 310
rect -86 284 -46 310
rect -20 284 20 310
rect 46 284 86 310
rect 112 284 152 310
rect 178 284 218 310
rect 244 284 284 310
rect 310 284 316 310
rect -316 244 316 284
rect -316 218 -310 244
rect -284 218 -244 244
rect -218 218 -178 244
rect -152 218 -112 244
rect -86 218 -46 244
rect -20 218 20 244
rect 46 218 86 244
rect 112 218 152 244
rect 178 218 218 244
rect 244 218 284 244
rect 310 218 316 244
rect -316 178 316 218
rect -316 152 -310 178
rect -284 152 -244 178
rect -218 152 -178 178
rect -152 152 -112 178
rect -86 152 -46 178
rect -20 152 20 178
rect 46 152 86 178
rect 112 152 152 178
rect 178 152 218 178
rect 244 152 284 178
rect 310 152 316 178
rect -316 112 316 152
rect -316 86 -310 112
rect -284 86 -244 112
rect -218 86 -178 112
rect -152 86 -112 112
rect -86 86 -46 112
rect -20 86 20 112
rect 46 86 86 112
rect 112 86 152 112
rect 178 86 218 112
rect 244 86 284 112
rect 310 86 316 112
rect -316 46 316 86
rect -316 20 -310 46
rect -284 20 -244 46
rect -218 20 -178 46
rect -152 20 -112 46
rect -86 20 -46 46
rect -20 20 20 46
rect 46 20 86 46
rect 112 20 152 46
rect 178 20 218 46
rect 244 20 284 46
rect 310 20 316 46
rect -316 -20 316 20
rect -316 -46 -310 -20
rect -284 -46 -244 -20
rect -218 -46 -178 -20
rect -152 -46 -112 -20
rect -86 -46 -46 -20
rect -20 -46 20 -20
rect 46 -46 86 -20
rect 112 -46 152 -20
rect 178 -46 218 -20
rect 244 -46 284 -20
rect 310 -46 316 -20
rect -316 -86 316 -46
rect -316 -112 -310 -86
rect -284 -112 -244 -86
rect -218 -112 -178 -86
rect -152 -112 -112 -86
rect -86 -112 -46 -86
rect -20 -112 20 -86
rect 46 -112 86 -86
rect 112 -112 152 -86
rect 178 -112 218 -86
rect 244 -112 284 -86
rect 310 -112 316 -86
rect -316 -152 316 -112
rect -316 -178 -310 -152
rect -284 -178 -244 -152
rect -218 -178 -178 -152
rect -152 -178 -112 -152
rect -86 -178 -46 -152
rect -20 -178 20 -152
rect 46 -178 86 -152
rect 112 -178 152 -152
rect 178 -178 218 -152
rect 244 -178 284 -152
rect 310 -178 316 -152
rect -316 -218 316 -178
rect -316 -244 -310 -218
rect -284 -244 -244 -218
rect -218 -244 -178 -218
rect -152 -244 -112 -218
rect -86 -244 -46 -218
rect -20 -244 20 -218
rect 46 -244 86 -218
rect 112 -244 152 -218
rect 178 -244 218 -218
rect 244 -244 284 -218
rect 310 -244 316 -218
rect -316 -284 316 -244
rect -316 -310 -310 -284
rect -284 -310 -244 -284
rect -218 -310 -178 -284
rect -152 -310 -112 -284
rect -86 -310 -46 -284
rect -20 -310 20 -284
rect 46 -310 86 -284
rect 112 -310 152 -284
rect 178 -310 218 -284
rect 244 -310 284 -284
rect 310 -310 316 -284
rect -316 -316 316 -310
<< end >>
