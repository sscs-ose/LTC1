magic
tech gf180mcuC
magscale 1 10
timestamp 1692680230
<< error_p >>
rect -3394 628 -3383 674
rect -3226 628 -3215 674
rect -3058 628 -3047 674
rect -2890 628 -2879 674
rect -2722 628 -2711 674
rect -2554 628 -2543 674
rect -2386 628 -2375 674
rect -2218 628 -2207 674
rect -2050 628 -2039 674
rect -1882 628 -1871 674
rect -1714 628 -1703 674
rect -1546 628 -1535 674
rect -1378 628 -1367 674
rect -1210 628 -1199 674
rect -1042 628 -1031 674
rect -874 628 -863 674
rect -706 628 -695 674
rect -538 628 -527 674
rect -370 628 -359 674
rect -202 628 -191 674
rect -34 628 -23 674
rect 134 628 145 674
rect 302 628 313 674
rect 470 628 481 674
rect 638 628 649 674
rect 806 628 817 674
rect 974 628 985 674
rect 1142 628 1153 674
rect 1310 628 1321 674
rect 1478 628 1489 674
rect 1646 628 1657 674
rect 1814 628 1825 674
rect 1982 628 1993 674
rect 2150 628 2161 674
rect 2318 628 2329 674
rect 2486 628 2497 674
rect 2654 628 2665 674
rect 2822 628 2833 674
rect 2990 628 3001 674
rect 3158 628 3169 674
rect 3326 628 3337 674
rect -3394 442 -3383 488
rect -3226 442 -3215 488
rect -3058 442 -3047 488
rect -2890 442 -2879 488
rect -2722 442 -2711 488
rect -2554 442 -2543 488
rect -2386 442 -2375 488
rect -2218 442 -2207 488
rect -2050 442 -2039 488
rect -1882 442 -1871 488
rect -1714 442 -1703 488
rect -1546 442 -1535 488
rect -1378 442 -1367 488
rect -1210 442 -1199 488
rect -1042 442 -1031 488
rect -874 442 -863 488
rect -706 442 -695 488
rect -538 442 -527 488
rect -370 442 -359 488
rect -202 442 -191 488
rect -34 442 -23 488
rect 134 442 145 488
rect 302 442 313 488
rect 470 442 481 488
rect 638 442 649 488
rect 806 442 817 488
rect 974 442 985 488
rect 1142 442 1153 488
rect 1310 442 1321 488
rect 1478 442 1489 488
rect 1646 442 1657 488
rect 1814 442 1825 488
rect 1982 442 1993 488
rect 2150 442 2161 488
rect 2318 442 2329 488
rect 2486 442 2497 488
rect 2654 442 2665 488
rect 2822 442 2833 488
rect 2990 442 3001 488
rect 3158 442 3169 488
rect 3326 442 3337 488
rect -3394 256 -3383 302
rect -3226 256 -3215 302
rect -3058 256 -3047 302
rect -2890 256 -2879 302
rect -2722 256 -2711 302
rect -2554 256 -2543 302
rect -2386 256 -2375 302
rect -2218 256 -2207 302
rect -2050 256 -2039 302
rect -1882 256 -1871 302
rect -1714 256 -1703 302
rect -1546 256 -1535 302
rect -1378 256 -1367 302
rect -1210 256 -1199 302
rect -1042 256 -1031 302
rect -874 256 -863 302
rect -706 256 -695 302
rect -538 256 -527 302
rect -370 256 -359 302
rect -202 256 -191 302
rect -34 256 -23 302
rect 134 256 145 302
rect 302 256 313 302
rect 470 256 481 302
rect 638 256 649 302
rect 806 256 817 302
rect 974 256 985 302
rect 1142 256 1153 302
rect 1310 256 1321 302
rect 1478 256 1489 302
rect 1646 256 1657 302
rect 1814 256 1825 302
rect 1982 256 1993 302
rect 2150 256 2161 302
rect 2318 256 2329 302
rect 2486 256 2497 302
rect 2654 256 2665 302
rect 2822 256 2833 302
rect 2990 256 3001 302
rect 3158 256 3169 302
rect 3326 256 3337 302
rect -3394 70 -3383 116
rect -3226 70 -3215 116
rect -3058 70 -3047 116
rect -2890 70 -2879 116
rect -2722 70 -2711 116
rect -2554 70 -2543 116
rect -2386 70 -2375 116
rect -2218 70 -2207 116
rect -2050 70 -2039 116
rect -1882 70 -1871 116
rect -1714 70 -1703 116
rect -1546 70 -1535 116
rect -1378 70 -1367 116
rect -1210 70 -1199 116
rect -1042 70 -1031 116
rect -874 70 -863 116
rect -706 70 -695 116
rect -538 70 -527 116
rect -370 70 -359 116
rect -202 70 -191 116
rect -34 70 -23 116
rect 134 70 145 116
rect 302 70 313 116
rect 470 70 481 116
rect 638 70 649 116
rect 806 70 817 116
rect 974 70 985 116
rect 1142 70 1153 116
rect 1310 70 1321 116
rect 1478 70 1489 116
rect 1646 70 1657 116
rect 1814 70 1825 116
rect 1982 70 1993 116
rect 2150 70 2161 116
rect 2318 70 2329 116
rect 2486 70 2497 116
rect 2654 70 2665 116
rect 2822 70 2833 116
rect 2990 70 3001 116
rect 3158 70 3169 116
rect 3326 70 3337 116
rect -3394 -116 -3383 -70
rect -3226 -116 -3215 -70
rect -3058 -116 -3047 -70
rect -2890 -116 -2879 -70
rect -2722 -116 -2711 -70
rect -2554 -116 -2543 -70
rect -2386 -116 -2375 -70
rect -2218 -116 -2207 -70
rect -2050 -116 -2039 -70
rect -1882 -116 -1871 -70
rect -1714 -116 -1703 -70
rect -1546 -116 -1535 -70
rect -1378 -116 -1367 -70
rect -1210 -116 -1199 -70
rect -1042 -116 -1031 -70
rect -874 -116 -863 -70
rect -706 -116 -695 -70
rect -538 -116 -527 -70
rect -370 -116 -359 -70
rect -202 -116 -191 -70
rect -34 -116 -23 -70
rect 134 -116 145 -70
rect 302 -116 313 -70
rect 470 -116 481 -70
rect 638 -116 649 -70
rect 806 -116 817 -70
rect 974 -116 985 -70
rect 1142 -116 1153 -70
rect 1310 -116 1321 -70
rect 1478 -116 1489 -70
rect 1646 -116 1657 -70
rect 1814 -116 1825 -70
rect 1982 -116 1993 -70
rect 2150 -116 2161 -70
rect 2318 -116 2329 -70
rect 2486 -116 2497 -70
rect 2654 -116 2665 -70
rect 2822 -116 2833 -70
rect 2990 -116 3001 -70
rect 3158 -116 3169 -70
rect 3326 -116 3337 -70
rect -3394 -302 -3383 -256
rect -3226 -302 -3215 -256
rect -3058 -302 -3047 -256
rect -2890 -302 -2879 -256
rect -2722 -302 -2711 -256
rect -2554 -302 -2543 -256
rect -2386 -302 -2375 -256
rect -2218 -302 -2207 -256
rect -2050 -302 -2039 -256
rect -1882 -302 -1871 -256
rect -1714 -302 -1703 -256
rect -1546 -302 -1535 -256
rect -1378 -302 -1367 -256
rect -1210 -302 -1199 -256
rect -1042 -302 -1031 -256
rect -874 -302 -863 -256
rect -706 -302 -695 -256
rect -538 -302 -527 -256
rect -370 -302 -359 -256
rect -202 -302 -191 -256
rect -34 -302 -23 -256
rect 134 -302 145 -256
rect 302 -302 313 -256
rect 470 -302 481 -256
rect 638 -302 649 -256
rect 806 -302 817 -256
rect 974 -302 985 -256
rect 1142 -302 1153 -256
rect 1310 -302 1321 -256
rect 1478 -302 1489 -256
rect 1646 -302 1657 -256
rect 1814 -302 1825 -256
rect 1982 -302 1993 -256
rect 2150 -302 2161 -256
rect 2318 -302 2329 -256
rect 2486 -302 2497 -256
rect 2654 -302 2665 -256
rect 2822 -302 2833 -256
rect 2990 -302 3001 -256
rect 3158 -302 3169 -256
rect 3326 -302 3337 -256
rect -3394 -488 -3383 -442
rect -3226 -488 -3215 -442
rect -3058 -488 -3047 -442
rect -2890 -488 -2879 -442
rect -2722 -488 -2711 -442
rect -2554 -488 -2543 -442
rect -2386 -488 -2375 -442
rect -2218 -488 -2207 -442
rect -2050 -488 -2039 -442
rect -1882 -488 -1871 -442
rect -1714 -488 -1703 -442
rect -1546 -488 -1535 -442
rect -1378 -488 -1367 -442
rect -1210 -488 -1199 -442
rect -1042 -488 -1031 -442
rect -874 -488 -863 -442
rect -706 -488 -695 -442
rect -538 -488 -527 -442
rect -370 -488 -359 -442
rect -202 -488 -191 -442
rect -34 -488 -23 -442
rect 134 -488 145 -442
rect 302 -488 313 -442
rect 470 -488 481 -442
rect 638 -488 649 -442
rect 806 -488 817 -442
rect 974 -488 985 -442
rect 1142 -488 1153 -442
rect 1310 -488 1321 -442
rect 1478 -488 1489 -442
rect 1646 -488 1657 -442
rect 1814 -488 1825 -442
rect 1982 -488 1993 -442
rect 2150 -488 2161 -442
rect 2318 -488 2329 -442
rect 2486 -488 2497 -442
rect 2654 -488 2665 -442
rect 2822 -488 2833 -442
rect 2990 -488 3001 -442
rect 3158 -488 3169 -442
rect 3326 -488 3337 -442
rect -3394 -674 -3383 -628
rect -3226 -674 -3215 -628
rect -3058 -674 -3047 -628
rect -2890 -674 -2879 -628
rect -2722 -674 -2711 -628
rect -2554 -674 -2543 -628
rect -2386 -674 -2375 -628
rect -2218 -674 -2207 -628
rect -2050 -674 -2039 -628
rect -1882 -674 -1871 -628
rect -1714 -674 -1703 -628
rect -1546 -674 -1535 -628
rect -1378 -674 -1367 -628
rect -1210 -674 -1199 -628
rect -1042 -674 -1031 -628
rect -874 -674 -863 -628
rect -706 -674 -695 -628
rect -538 -674 -527 -628
rect -370 -674 -359 -628
rect -202 -674 -191 -628
rect -34 -674 -23 -628
rect 134 -674 145 -628
rect 302 -674 313 -628
rect 470 -674 481 -628
rect 638 -674 649 -628
rect 806 -674 817 -628
rect 974 -674 985 -628
rect 1142 -674 1153 -628
rect 1310 -674 1321 -628
rect 1478 -674 1489 -628
rect 1646 -674 1657 -628
rect 1814 -674 1825 -628
rect 1982 -674 1993 -628
rect 2150 -674 2161 -628
rect 2318 -674 2329 -628
rect 2486 -674 2497 -628
rect 2654 -674 2665 -628
rect 2822 -674 2833 -628
rect 2990 -674 3001 -628
rect 3158 -674 3169 -628
rect 3326 -674 3337 -628
<< pwell >>
rect -3420 -750 3420 750
<< nmos >>
rect -3304 626 -3248 676
rect -3136 626 -3080 676
rect -2968 626 -2912 676
rect -2800 626 -2744 676
rect -2632 626 -2576 676
rect -2464 626 -2408 676
rect -2296 626 -2240 676
rect -2128 626 -2072 676
rect -1960 626 -1904 676
rect -1792 626 -1736 676
rect -1624 626 -1568 676
rect -1456 626 -1400 676
rect -1288 626 -1232 676
rect -1120 626 -1064 676
rect -952 626 -896 676
rect -784 626 -728 676
rect -616 626 -560 676
rect -448 626 -392 676
rect -280 626 -224 676
rect -112 626 -56 676
rect 56 626 112 676
rect 224 626 280 676
rect 392 626 448 676
rect 560 626 616 676
rect 728 626 784 676
rect 896 626 952 676
rect 1064 626 1120 676
rect 1232 626 1288 676
rect 1400 626 1456 676
rect 1568 626 1624 676
rect 1736 626 1792 676
rect 1904 626 1960 676
rect 2072 626 2128 676
rect 2240 626 2296 676
rect 2408 626 2464 676
rect 2576 626 2632 676
rect 2744 626 2800 676
rect 2912 626 2968 676
rect 3080 626 3136 676
rect 3248 626 3304 676
rect -3304 440 -3248 490
rect -3136 440 -3080 490
rect -2968 440 -2912 490
rect -2800 440 -2744 490
rect -2632 440 -2576 490
rect -2464 440 -2408 490
rect -2296 440 -2240 490
rect -2128 440 -2072 490
rect -1960 440 -1904 490
rect -1792 440 -1736 490
rect -1624 440 -1568 490
rect -1456 440 -1400 490
rect -1288 440 -1232 490
rect -1120 440 -1064 490
rect -952 440 -896 490
rect -784 440 -728 490
rect -616 440 -560 490
rect -448 440 -392 490
rect -280 440 -224 490
rect -112 440 -56 490
rect 56 440 112 490
rect 224 440 280 490
rect 392 440 448 490
rect 560 440 616 490
rect 728 440 784 490
rect 896 440 952 490
rect 1064 440 1120 490
rect 1232 440 1288 490
rect 1400 440 1456 490
rect 1568 440 1624 490
rect 1736 440 1792 490
rect 1904 440 1960 490
rect 2072 440 2128 490
rect 2240 440 2296 490
rect 2408 440 2464 490
rect 2576 440 2632 490
rect 2744 440 2800 490
rect 2912 440 2968 490
rect 3080 440 3136 490
rect 3248 440 3304 490
rect -3304 254 -3248 304
rect -3136 254 -3080 304
rect -2968 254 -2912 304
rect -2800 254 -2744 304
rect -2632 254 -2576 304
rect -2464 254 -2408 304
rect -2296 254 -2240 304
rect -2128 254 -2072 304
rect -1960 254 -1904 304
rect -1792 254 -1736 304
rect -1624 254 -1568 304
rect -1456 254 -1400 304
rect -1288 254 -1232 304
rect -1120 254 -1064 304
rect -952 254 -896 304
rect -784 254 -728 304
rect -616 254 -560 304
rect -448 254 -392 304
rect -280 254 -224 304
rect -112 254 -56 304
rect 56 254 112 304
rect 224 254 280 304
rect 392 254 448 304
rect 560 254 616 304
rect 728 254 784 304
rect 896 254 952 304
rect 1064 254 1120 304
rect 1232 254 1288 304
rect 1400 254 1456 304
rect 1568 254 1624 304
rect 1736 254 1792 304
rect 1904 254 1960 304
rect 2072 254 2128 304
rect 2240 254 2296 304
rect 2408 254 2464 304
rect 2576 254 2632 304
rect 2744 254 2800 304
rect 2912 254 2968 304
rect 3080 254 3136 304
rect 3248 254 3304 304
rect -3304 68 -3248 118
rect -3136 68 -3080 118
rect -2968 68 -2912 118
rect -2800 68 -2744 118
rect -2632 68 -2576 118
rect -2464 68 -2408 118
rect -2296 68 -2240 118
rect -2128 68 -2072 118
rect -1960 68 -1904 118
rect -1792 68 -1736 118
rect -1624 68 -1568 118
rect -1456 68 -1400 118
rect -1288 68 -1232 118
rect -1120 68 -1064 118
rect -952 68 -896 118
rect -784 68 -728 118
rect -616 68 -560 118
rect -448 68 -392 118
rect -280 68 -224 118
rect -112 68 -56 118
rect 56 68 112 118
rect 224 68 280 118
rect 392 68 448 118
rect 560 68 616 118
rect 728 68 784 118
rect 896 68 952 118
rect 1064 68 1120 118
rect 1232 68 1288 118
rect 1400 68 1456 118
rect 1568 68 1624 118
rect 1736 68 1792 118
rect 1904 68 1960 118
rect 2072 68 2128 118
rect 2240 68 2296 118
rect 2408 68 2464 118
rect 2576 68 2632 118
rect 2744 68 2800 118
rect 2912 68 2968 118
rect 3080 68 3136 118
rect 3248 68 3304 118
rect -3304 -118 -3248 -68
rect -3136 -118 -3080 -68
rect -2968 -118 -2912 -68
rect -2800 -118 -2744 -68
rect -2632 -118 -2576 -68
rect -2464 -118 -2408 -68
rect -2296 -118 -2240 -68
rect -2128 -118 -2072 -68
rect -1960 -118 -1904 -68
rect -1792 -118 -1736 -68
rect -1624 -118 -1568 -68
rect -1456 -118 -1400 -68
rect -1288 -118 -1232 -68
rect -1120 -118 -1064 -68
rect -952 -118 -896 -68
rect -784 -118 -728 -68
rect -616 -118 -560 -68
rect -448 -118 -392 -68
rect -280 -118 -224 -68
rect -112 -118 -56 -68
rect 56 -118 112 -68
rect 224 -118 280 -68
rect 392 -118 448 -68
rect 560 -118 616 -68
rect 728 -118 784 -68
rect 896 -118 952 -68
rect 1064 -118 1120 -68
rect 1232 -118 1288 -68
rect 1400 -118 1456 -68
rect 1568 -118 1624 -68
rect 1736 -118 1792 -68
rect 1904 -118 1960 -68
rect 2072 -118 2128 -68
rect 2240 -118 2296 -68
rect 2408 -118 2464 -68
rect 2576 -118 2632 -68
rect 2744 -118 2800 -68
rect 2912 -118 2968 -68
rect 3080 -118 3136 -68
rect 3248 -118 3304 -68
rect -3304 -304 -3248 -254
rect -3136 -304 -3080 -254
rect -2968 -304 -2912 -254
rect -2800 -304 -2744 -254
rect -2632 -304 -2576 -254
rect -2464 -304 -2408 -254
rect -2296 -304 -2240 -254
rect -2128 -304 -2072 -254
rect -1960 -304 -1904 -254
rect -1792 -304 -1736 -254
rect -1624 -304 -1568 -254
rect -1456 -304 -1400 -254
rect -1288 -304 -1232 -254
rect -1120 -304 -1064 -254
rect -952 -304 -896 -254
rect -784 -304 -728 -254
rect -616 -304 -560 -254
rect -448 -304 -392 -254
rect -280 -304 -224 -254
rect -112 -304 -56 -254
rect 56 -304 112 -254
rect 224 -304 280 -254
rect 392 -304 448 -254
rect 560 -304 616 -254
rect 728 -304 784 -254
rect 896 -304 952 -254
rect 1064 -304 1120 -254
rect 1232 -304 1288 -254
rect 1400 -304 1456 -254
rect 1568 -304 1624 -254
rect 1736 -304 1792 -254
rect 1904 -304 1960 -254
rect 2072 -304 2128 -254
rect 2240 -304 2296 -254
rect 2408 -304 2464 -254
rect 2576 -304 2632 -254
rect 2744 -304 2800 -254
rect 2912 -304 2968 -254
rect 3080 -304 3136 -254
rect 3248 -304 3304 -254
rect -3304 -490 -3248 -440
rect -3136 -490 -3080 -440
rect -2968 -490 -2912 -440
rect -2800 -490 -2744 -440
rect -2632 -490 -2576 -440
rect -2464 -490 -2408 -440
rect -2296 -490 -2240 -440
rect -2128 -490 -2072 -440
rect -1960 -490 -1904 -440
rect -1792 -490 -1736 -440
rect -1624 -490 -1568 -440
rect -1456 -490 -1400 -440
rect -1288 -490 -1232 -440
rect -1120 -490 -1064 -440
rect -952 -490 -896 -440
rect -784 -490 -728 -440
rect -616 -490 -560 -440
rect -448 -490 -392 -440
rect -280 -490 -224 -440
rect -112 -490 -56 -440
rect 56 -490 112 -440
rect 224 -490 280 -440
rect 392 -490 448 -440
rect 560 -490 616 -440
rect 728 -490 784 -440
rect 896 -490 952 -440
rect 1064 -490 1120 -440
rect 1232 -490 1288 -440
rect 1400 -490 1456 -440
rect 1568 -490 1624 -440
rect 1736 -490 1792 -440
rect 1904 -490 1960 -440
rect 2072 -490 2128 -440
rect 2240 -490 2296 -440
rect 2408 -490 2464 -440
rect 2576 -490 2632 -440
rect 2744 -490 2800 -440
rect 2912 -490 2968 -440
rect 3080 -490 3136 -440
rect 3248 -490 3304 -440
rect -3304 -676 -3248 -626
rect -3136 -676 -3080 -626
rect -2968 -676 -2912 -626
rect -2800 -676 -2744 -626
rect -2632 -676 -2576 -626
rect -2464 -676 -2408 -626
rect -2296 -676 -2240 -626
rect -2128 -676 -2072 -626
rect -1960 -676 -1904 -626
rect -1792 -676 -1736 -626
rect -1624 -676 -1568 -626
rect -1456 -676 -1400 -626
rect -1288 -676 -1232 -626
rect -1120 -676 -1064 -626
rect -952 -676 -896 -626
rect -784 -676 -728 -626
rect -616 -676 -560 -626
rect -448 -676 -392 -626
rect -280 -676 -224 -626
rect -112 -676 -56 -626
rect 56 -676 112 -626
rect 224 -676 280 -626
rect 392 -676 448 -626
rect 560 -676 616 -626
rect 728 -676 784 -626
rect 896 -676 952 -626
rect 1064 -676 1120 -626
rect 1232 -676 1288 -626
rect 1400 -676 1456 -626
rect 1568 -676 1624 -626
rect 1736 -676 1792 -626
rect 1904 -676 1960 -626
rect 2072 -676 2128 -626
rect 2240 -676 2296 -626
rect 2408 -676 2464 -626
rect 2576 -676 2632 -626
rect 2744 -676 2800 -626
rect 2912 -676 2968 -626
rect 3080 -676 3136 -626
rect 3248 -676 3304 -626
<< ndiff >>
rect -3396 676 -3324 687
rect -3228 676 -3156 687
rect -3060 676 -2988 687
rect -2892 676 -2820 687
rect -2724 676 -2652 687
rect -2556 676 -2484 687
rect -2388 676 -2316 687
rect -2220 676 -2148 687
rect -2052 676 -1980 687
rect -1884 676 -1812 687
rect -1716 676 -1644 687
rect -1548 676 -1476 687
rect -1380 676 -1308 687
rect -1212 676 -1140 687
rect -1044 676 -972 687
rect -876 676 -804 687
rect -708 676 -636 687
rect -540 676 -468 687
rect -372 676 -300 687
rect -204 676 -132 687
rect -36 676 36 687
rect 132 676 204 687
rect 300 676 372 687
rect 468 676 540 687
rect 636 676 708 687
rect 804 676 876 687
rect 972 676 1044 687
rect 1140 676 1212 687
rect 1308 676 1380 687
rect 1476 676 1548 687
rect 1644 676 1716 687
rect 1812 676 1884 687
rect 1980 676 2052 687
rect 2148 676 2220 687
rect 2316 676 2388 687
rect 2484 676 2556 687
rect 2652 676 2724 687
rect 2820 676 2892 687
rect 2988 676 3060 687
rect 3156 676 3228 687
rect 3324 676 3396 687
rect -3396 674 -3304 676
rect -3396 628 -3383 674
rect -3337 628 -3304 674
rect -3396 626 -3304 628
rect -3248 674 -3136 676
rect -3248 628 -3215 674
rect -3169 628 -3136 674
rect -3248 626 -3136 628
rect -3080 674 -2968 676
rect -3080 628 -3047 674
rect -3001 628 -2968 674
rect -3080 626 -2968 628
rect -2912 674 -2800 676
rect -2912 628 -2879 674
rect -2833 628 -2800 674
rect -2912 626 -2800 628
rect -2744 674 -2632 676
rect -2744 628 -2711 674
rect -2665 628 -2632 674
rect -2744 626 -2632 628
rect -2576 674 -2464 676
rect -2576 628 -2543 674
rect -2497 628 -2464 674
rect -2576 626 -2464 628
rect -2408 674 -2296 676
rect -2408 628 -2375 674
rect -2329 628 -2296 674
rect -2408 626 -2296 628
rect -2240 674 -2128 676
rect -2240 628 -2207 674
rect -2161 628 -2128 674
rect -2240 626 -2128 628
rect -2072 674 -1960 676
rect -2072 628 -2039 674
rect -1993 628 -1960 674
rect -2072 626 -1960 628
rect -1904 674 -1792 676
rect -1904 628 -1871 674
rect -1825 628 -1792 674
rect -1904 626 -1792 628
rect -1736 674 -1624 676
rect -1736 628 -1703 674
rect -1657 628 -1624 674
rect -1736 626 -1624 628
rect -1568 674 -1456 676
rect -1568 628 -1535 674
rect -1489 628 -1456 674
rect -1568 626 -1456 628
rect -1400 674 -1288 676
rect -1400 628 -1367 674
rect -1321 628 -1288 674
rect -1400 626 -1288 628
rect -1232 674 -1120 676
rect -1232 628 -1199 674
rect -1153 628 -1120 674
rect -1232 626 -1120 628
rect -1064 674 -952 676
rect -1064 628 -1031 674
rect -985 628 -952 674
rect -1064 626 -952 628
rect -896 674 -784 676
rect -896 628 -863 674
rect -817 628 -784 674
rect -896 626 -784 628
rect -728 674 -616 676
rect -728 628 -695 674
rect -649 628 -616 674
rect -728 626 -616 628
rect -560 674 -448 676
rect -560 628 -527 674
rect -481 628 -448 674
rect -560 626 -448 628
rect -392 674 -280 676
rect -392 628 -359 674
rect -313 628 -280 674
rect -392 626 -280 628
rect -224 674 -112 676
rect -224 628 -191 674
rect -145 628 -112 674
rect -224 626 -112 628
rect -56 674 56 676
rect -56 628 -23 674
rect 23 628 56 674
rect -56 626 56 628
rect 112 674 224 676
rect 112 628 145 674
rect 191 628 224 674
rect 112 626 224 628
rect 280 674 392 676
rect 280 628 313 674
rect 359 628 392 674
rect 280 626 392 628
rect 448 674 560 676
rect 448 628 481 674
rect 527 628 560 674
rect 448 626 560 628
rect 616 674 728 676
rect 616 628 649 674
rect 695 628 728 674
rect 616 626 728 628
rect 784 674 896 676
rect 784 628 817 674
rect 863 628 896 674
rect 784 626 896 628
rect 952 674 1064 676
rect 952 628 985 674
rect 1031 628 1064 674
rect 952 626 1064 628
rect 1120 674 1232 676
rect 1120 628 1153 674
rect 1199 628 1232 674
rect 1120 626 1232 628
rect 1288 674 1400 676
rect 1288 628 1321 674
rect 1367 628 1400 674
rect 1288 626 1400 628
rect 1456 674 1568 676
rect 1456 628 1489 674
rect 1535 628 1568 674
rect 1456 626 1568 628
rect 1624 674 1736 676
rect 1624 628 1657 674
rect 1703 628 1736 674
rect 1624 626 1736 628
rect 1792 674 1904 676
rect 1792 628 1825 674
rect 1871 628 1904 674
rect 1792 626 1904 628
rect 1960 674 2072 676
rect 1960 628 1993 674
rect 2039 628 2072 674
rect 1960 626 2072 628
rect 2128 674 2240 676
rect 2128 628 2161 674
rect 2207 628 2240 674
rect 2128 626 2240 628
rect 2296 674 2408 676
rect 2296 628 2329 674
rect 2375 628 2408 674
rect 2296 626 2408 628
rect 2464 674 2576 676
rect 2464 628 2497 674
rect 2543 628 2576 674
rect 2464 626 2576 628
rect 2632 674 2744 676
rect 2632 628 2665 674
rect 2711 628 2744 674
rect 2632 626 2744 628
rect 2800 674 2912 676
rect 2800 628 2833 674
rect 2879 628 2912 674
rect 2800 626 2912 628
rect 2968 674 3080 676
rect 2968 628 3001 674
rect 3047 628 3080 674
rect 2968 626 3080 628
rect 3136 674 3248 676
rect 3136 628 3169 674
rect 3215 628 3248 674
rect 3136 626 3248 628
rect 3304 674 3396 676
rect 3304 628 3337 674
rect 3383 628 3396 674
rect 3304 626 3396 628
rect -3396 615 -3324 626
rect -3228 615 -3156 626
rect -3060 615 -2988 626
rect -2892 615 -2820 626
rect -2724 615 -2652 626
rect -2556 615 -2484 626
rect -2388 615 -2316 626
rect -2220 615 -2148 626
rect -2052 615 -1980 626
rect -1884 615 -1812 626
rect -1716 615 -1644 626
rect -1548 615 -1476 626
rect -1380 615 -1308 626
rect -1212 615 -1140 626
rect -1044 615 -972 626
rect -876 615 -804 626
rect -708 615 -636 626
rect -540 615 -468 626
rect -372 615 -300 626
rect -204 615 -132 626
rect -36 615 36 626
rect 132 615 204 626
rect 300 615 372 626
rect 468 615 540 626
rect 636 615 708 626
rect 804 615 876 626
rect 972 615 1044 626
rect 1140 615 1212 626
rect 1308 615 1380 626
rect 1476 615 1548 626
rect 1644 615 1716 626
rect 1812 615 1884 626
rect 1980 615 2052 626
rect 2148 615 2220 626
rect 2316 615 2388 626
rect 2484 615 2556 626
rect 2652 615 2724 626
rect 2820 615 2892 626
rect 2988 615 3060 626
rect 3156 615 3228 626
rect 3324 615 3396 626
rect -3396 490 -3324 501
rect -3228 490 -3156 501
rect -3060 490 -2988 501
rect -2892 490 -2820 501
rect -2724 490 -2652 501
rect -2556 490 -2484 501
rect -2388 490 -2316 501
rect -2220 490 -2148 501
rect -2052 490 -1980 501
rect -1884 490 -1812 501
rect -1716 490 -1644 501
rect -1548 490 -1476 501
rect -1380 490 -1308 501
rect -1212 490 -1140 501
rect -1044 490 -972 501
rect -876 490 -804 501
rect -708 490 -636 501
rect -540 490 -468 501
rect -372 490 -300 501
rect -204 490 -132 501
rect -36 490 36 501
rect 132 490 204 501
rect 300 490 372 501
rect 468 490 540 501
rect 636 490 708 501
rect 804 490 876 501
rect 972 490 1044 501
rect 1140 490 1212 501
rect 1308 490 1380 501
rect 1476 490 1548 501
rect 1644 490 1716 501
rect 1812 490 1884 501
rect 1980 490 2052 501
rect 2148 490 2220 501
rect 2316 490 2388 501
rect 2484 490 2556 501
rect 2652 490 2724 501
rect 2820 490 2892 501
rect 2988 490 3060 501
rect 3156 490 3228 501
rect 3324 490 3396 501
rect -3396 488 -3304 490
rect -3396 442 -3383 488
rect -3337 442 -3304 488
rect -3396 440 -3304 442
rect -3248 488 -3136 490
rect -3248 442 -3215 488
rect -3169 442 -3136 488
rect -3248 440 -3136 442
rect -3080 488 -2968 490
rect -3080 442 -3047 488
rect -3001 442 -2968 488
rect -3080 440 -2968 442
rect -2912 488 -2800 490
rect -2912 442 -2879 488
rect -2833 442 -2800 488
rect -2912 440 -2800 442
rect -2744 488 -2632 490
rect -2744 442 -2711 488
rect -2665 442 -2632 488
rect -2744 440 -2632 442
rect -2576 488 -2464 490
rect -2576 442 -2543 488
rect -2497 442 -2464 488
rect -2576 440 -2464 442
rect -2408 488 -2296 490
rect -2408 442 -2375 488
rect -2329 442 -2296 488
rect -2408 440 -2296 442
rect -2240 488 -2128 490
rect -2240 442 -2207 488
rect -2161 442 -2128 488
rect -2240 440 -2128 442
rect -2072 488 -1960 490
rect -2072 442 -2039 488
rect -1993 442 -1960 488
rect -2072 440 -1960 442
rect -1904 488 -1792 490
rect -1904 442 -1871 488
rect -1825 442 -1792 488
rect -1904 440 -1792 442
rect -1736 488 -1624 490
rect -1736 442 -1703 488
rect -1657 442 -1624 488
rect -1736 440 -1624 442
rect -1568 488 -1456 490
rect -1568 442 -1535 488
rect -1489 442 -1456 488
rect -1568 440 -1456 442
rect -1400 488 -1288 490
rect -1400 442 -1367 488
rect -1321 442 -1288 488
rect -1400 440 -1288 442
rect -1232 488 -1120 490
rect -1232 442 -1199 488
rect -1153 442 -1120 488
rect -1232 440 -1120 442
rect -1064 488 -952 490
rect -1064 442 -1031 488
rect -985 442 -952 488
rect -1064 440 -952 442
rect -896 488 -784 490
rect -896 442 -863 488
rect -817 442 -784 488
rect -896 440 -784 442
rect -728 488 -616 490
rect -728 442 -695 488
rect -649 442 -616 488
rect -728 440 -616 442
rect -560 488 -448 490
rect -560 442 -527 488
rect -481 442 -448 488
rect -560 440 -448 442
rect -392 488 -280 490
rect -392 442 -359 488
rect -313 442 -280 488
rect -392 440 -280 442
rect -224 488 -112 490
rect -224 442 -191 488
rect -145 442 -112 488
rect -224 440 -112 442
rect -56 488 56 490
rect -56 442 -23 488
rect 23 442 56 488
rect -56 440 56 442
rect 112 488 224 490
rect 112 442 145 488
rect 191 442 224 488
rect 112 440 224 442
rect 280 488 392 490
rect 280 442 313 488
rect 359 442 392 488
rect 280 440 392 442
rect 448 488 560 490
rect 448 442 481 488
rect 527 442 560 488
rect 448 440 560 442
rect 616 488 728 490
rect 616 442 649 488
rect 695 442 728 488
rect 616 440 728 442
rect 784 488 896 490
rect 784 442 817 488
rect 863 442 896 488
rect 784 440 896 442
rect 952 488 1064 490
rect 952 442 985 488
rect 1031 442 1064 488
rect 952 440 1064 442
rect 1120 488 1232 490
rect 1120 442 1153 488
rect 1199 442 1232 488
rect 1120 440 1232 442
rect 1288 488 1400 490
rect 1288 442 1321 488
rect 1367 442 1400 488
rect 1288 440 1400 442
rect 1456 488 1568 490
rect 1456 442 1489 488
rect 1535 442 1568 488
rect 1456 440 1568 442
rect 1624 488 1736 490
rect 1624 442 1657 488
rect 1703 442 1736 488
rect 1624 440 1736 442
rect 1792 488 1904 490
rect 1792 442 1825 488
rect 1871 442 1904 488
rect 1792 440 1904 442
rect 1960 488 2072 490
rect 1960 442 1993 488
rect 2039 442 2072 488
rect 1960 440 2072 442
rect 2128 488 2240 490
rect 2128 442 2161 488
rect 2207 442 2240 488
rect 2128 440 2240 442
rect 2296 488 2408 490
rect 2296 442 2329 488
rect 2375 442 2408 488
rect 2296 440 2408 442
rect 2464 488 2576 490
rect 2464 442 2497 488
rect 2543 442 2576 488
rect 2464 440 2576 442
rect 2632 488 2744 490
rect 2632 442 2665 488
rect 2711 442 2744 488
rect 2632 440 2744 442
rect 2800 488 2912 490
rect 2800 442 2833 488
rect 2879 442 2912 488
rect 2800 440 2912 442
rect 2968 488 3080 490
rect 2968 442 3001 488
rect 3047 442 3080 488
rect 2968 440 3080 442
rect 3136 488 3248 490
rect 3136 442 3169 488
rect 3215 442 3248 488
rect 3136 440 3248 442
rect 3304 488 3396 490
rect 3304 442 3337 488
rect 3383 442 3396 488
rect 3304 440 3396 442
rect -3396 429 -3324 440
rect -3228 429 -3156 440
rect -3060 429 -2988 440
rect -2892 429 -2820 440
rect -2724 429 -2652 440
rect -2556 429 -2484 440
rect -2388 429 -2316 440
rect -2220 429 -2148 440
rect -2052 429 -1980 440
rect -1884 429 -1812 440
rect -1716 429 -1644 440
rect -1548 429 -1476 440
rect -1380 429 -1308 440
rect -1212 429 -1140 440
rect -1044 429 -972 440
rect -876 429 -804 440
rect -708 429 -636 440
rect -540 429 -468 440
rect -372 429 -300 440
rect -204 429 -132 440
rect -36 429 36 440
rect 132 429 204 440
rect 300 429 372 440
rect 468 429 540 440
rect 636 429 708 440
rect 804 429 876 440
rect 972 429 1044 440
rect 1140 429 1212 440
rect 1308 429 1380 440
rect 1476 429 1548 440
rect 1644 429 1716 440
rect 1812 429 1884 440
rect 1980 429 2052 440
rect 2148 429 2220 440
rect 2316 429 2388 440
rect 2484 429 2556 440
rect 2652 429 2724 440
rect 2820 429 2892 440
rect 2988 429 3060 440
rect 3156 429 3228 440
rect 3324 429 3396 440
rect -3396 304 -3324 315
rect -3228 304 -3156 315
rect -3060 304 -2988 315
rect -2892 304 -2820 315
rect -2724 304 -2652 315
rect -2556 304 -2484 315
rect -2388 304 -2316 315
rect -2220 304 -2148 315
rect -2052 304 -1980 315
rect -1884 304 -1812 315
rect -1716 304 -1644 315
rect -1548 304 -1476 315
rect -1380 304 -1308 315
rect -1212 304 -1140 315
rect -1044 304 -972 315
rect -876 304 -804 315
rect -708 304 -636 315
rect -540 304 -468 315
rect -372 304 -300 315
rect -204 304 -132 315
rect -36 304 36 315
rect 132 304 204 315
rect 300 304 372 315
rect 468 304 540 315
rect 636 304 708 315
rect 804 304 876 315
rect 972 304 1044 315
rect 1140 304 1212 315
rect 1308 304 1380 315
rect 1476 304 1548 315
rect 1644 304 1716 315
rect 1812 304 1884 315
rect 1980 304 2052 315
rect 2148 304 2220 315
rect 2316 304 2388 315
rect 2484 304 2556 315
rect 2652 304 2724 315
rect 2820 304 2892 315
rect 2988 304 3060 315
rect 3156 304 3228 315
rect 3324 304 3396 315
rect -3396 302 -3304 304
rect -3396 256 -3383 302
rect -3337 256 -3304 302
rect -3396 254 -3304 256
rect -3248 302 -3136 304
rect -3248 256 -3215 302
rect -3169 256 -3136 302
rect -3248 254 -3136 256
rect -3080 302 -2968 304
rect -3080 256 -3047 302
rect -3001 256 -2968 302
rect -3080 254 -2968 256
rect -2912 302 -2800 304
rect -2912 256 -2879 302
rect -2833 256 -2800 302
rect -2912 254 -2800 256
rect -2744 302 -2632 304
rect -2744 256 -2711 302
rect -2665 256 -2632 302
rect -2744 254 -2632 256
rect -2576 302 -2464 304
rect -2576 256 -2543 302
rect -2497 256 -2464 302
rect -2576 254 -2464 256
rect -2408 302 -2296 304
rect -2408 256 -2375 302
rect -2329 256 -2296 302
rect -2408 254 -2296 256
rect -2240 302 -2128 304
rect -2240 256 -2207 302
rect -2161 256 -2128 302
rect -2240 254 -2128 256
rect -2072 302 -1960 304
rect -2072 256 -2039 302
rect -1993 256 -1960 302
rect -2072 254 -1960 256
rect -1904 302 -1792 304
rect -1904 256 -1871 302
rect -1825 256 -1792 302
rect -1904 254 -1792 256
rect -1736 302 -1624 304
rect -1736 256 -1703 302
rect -1657 256 -1624 302
rect -1736 254 -1624 256
rect -1568 302 -1456 304
rect -1568 256 -1535 302
rect -1489 256 -1456 302
rect -1568 254 -1456 256
rect -1400 302 -1288 304
rect -1400 256 -1367 302
rect -1321 256 -1288 302
rect -1400 254 -1288 256
rect -1232 302 -1120 304
rect -1232 256 -1199 302
rect -1153 256 -1120 302
rect -1232 254 -1120 256
rect -1064 302 -952 304
rect -1064 256 -1031 302
rect -985 256 -952 302
rect -1064 254 -952 256
rect -896 302 -784 304
rect -896 256 -863 302
rect -817 256 -784 302
rect -896 254 -784 256
rect -728 302 -616 304
rect -728 256 -695 302
rect -649 256 -616 302
rect -728 254 -616 256
rect -560 302 -448 304
rect -560 256 -527 302
rect -481 256 -448 302
rect -560 254 -448 256
rect -392 302 -280 304
rect -392 256 -359 302
rect -313 256 -280 302
rect -392 254 -280 256
rect -224 302 -112 304
rect -224 256 -191 302
rect -145 256 -112 302
rect -224 254 -112 256
rect -56 302 56 304
rect -56 256 -23 302
rect 23 256 56 302
rect -56 254 56 256
rect 112 302 224 304
rect 112 256 145 302
rect 191 256 224 302
rect 112 254 224 256
rect 280 302 392 304
rect 280 256 313 302
rect 359 256 392 302
rect 280 254 392 256
rect 448 302 560 304
rect 448 256 481 302
rect 527 256 560 302
rect 448 254 560 256
rect 616 302 728 304
rect 616 256 649 302
rect 695 256 728 302
rect 616 254 728 256
rect 784 302 896 304
rect 784 256 817 302
rect 863 256 896 302
rect 784 254 896 256
rect 952 302 1064 304
rect 952 256 985 302
rect 1031 256 1064 302
rect 952 254 1064 256
rect 1120 302 1232 304
rect 1120 256 1153 302
rect 1199 256 1232 302
rect 1120 254 1232 256
rect 1288 302 1400 304
rect 1288 256 1321 302
rect 1367 256 1400 302
rect 1288 254 1400 256
rect 1456 302 1568 304
rect 1456 256 1489 302
rect 1535 256 1568 302
rect 1456 254 1568 256
rect 1624 302 1736 304
rect 1624 256 1657 302
rect 1703 256 1736 302
rect 1624 254 1736 256
rect 1792 302 1904 304
rect 1792 256 1825 302
rect 1871 256 1904 302
rect 1792 254 1904 256
rect 1960 302 2072 304
rect 1960 256 1993 302
rect 2039 256 2072 302
rect 1960 254 2072 256
rect 2128 302 2240 304
rect 2128 256 2161 302
rect 2207 256 2240 302
rect 2128 254 2240 256
rect 2296 302 2408 304
rect 2296 256 2329 302
rect 2375 256 2408 302
rect 2296 254 2408 256
rect 2464 302 2576 304
rect 2464 256 2497 302
rect 2543 256 2576 302
rect 2464 254 2576 256
rect 2632 302 2744 304
rect 2632 256 2665 302
rect 2711 256 2744 302
rect 2632 254 2744 256
rect 2800 302 2912 304
rect 2800 256 2833 302
rect 2879 256 2912 302
rect 2800 254 2912 256
rect 2968 302 3080 304
rect 2968 256 3001 302
rect 3047 256 3080 302
rect 2968 254 3080 256
rect 3136 302 3248 304
rect 3136 256 3169 302
rect 3215 256 3248 302
rect 3136 254 3248 256
rect 3304 302 3396 304
rect 3304 256 3337 302
rect 3383 256 3396 302
rect 3304 254 3396 256
rect -3396 243 -3324 254
rect -3228 243 -3156 254
rect -3060 243 -2988 254
rect -2892 243 -2820 254
rect -2724 243 -2652 254
rect -2556 243 -2484 254
rect -2388 243 -2316 254
rect -2220 243 -2148 254
rect -2052 243 -1980 254
rect -1884 243 -1812 254
rect -1716 243 -1644 254
rect -1548 243 -1476 254
rect -1380 243 -1308 254
rect -1212 243 -1140 254
rect -1044 243 -972 254
rect -876 243 -804 254
rect -708 243 -636 254
rect -540 243 -468 254
rect -372 243 -300 254
rect -204 243 -132 254
rect -36 243 36 254
rect 132 243 204 254
rect 300 243 372 254
rect 468 243 540 254
rect 636 243 708 254
rect 804 243 876 254
rect 972 243 1044 254
rect 1140 243 1212 254
rect 1308 243 1380 254
rect 1476 243 1548 254
rect 1644 243 1716 254
rect 1812 243 1884 254
rect 1980 243 2052 254
rect 2148 243 2220 254
rect 2316 243 2388 254
rect 2484 243 2556 254
rect 2652 243 2724 254
rect 2820 243 2892 254
rect 2988 243 3060 254
rect 3156 243 3228 254
rect 3324 243 3396 254
rect -3396 118 -3324 129
rect -3228 118 -3156 129
rect -3060 118 -2988 129
rect -2892 118 -2820 129
rect -2724 118 -2652 129
rect -2556 118 -2484 129
rect -2388 118 -2316 129
rect -2220 118 -2148 129
rect -2052 118 -1980 129
rect -1884 118 -1812 129
rect -1716 118 -1644 129
rect -1548 118 -1476 129
rect -1380 118 -1308 129
rect -1212 118 -1140 129
rect -1044 118 -972 129
rect -876 118 -804 129
rect -708 118 -636 129
rect -540 118 -468 129
rect -372 118 -300 129
rect -204 118 -132 129
rect -36 118 36 129
rect 132 118 204 129
rect 300 118 372 129
rect 468 118 540 129
rect 636 118 708 129
rect 804 118 876 129
rect 972 118 1044 129
rect 1140 118 1212 129
rect 1308 118 1380 129
rect 1476 118 1548 129
rect 1644 118 1716 129
rect 1812 118 1884 129
rect 1980 118 2052 129
rect 2148 118 2220 129
rect 2316 118 2388 129
rect 2484 118 2556 129
rect 2652 118 2724 129
rect 2820 118 2892 129
rect 2988 118 3060 129
rect 3156 118 3228 129
rect 3324 118 3396 129
rect -3396 116 -3304 118
rect -3396 70 -3383 116
rect -3337 70 -3304 116
rect -3396 68 -3304 70
rect -3248 116 -3136 118
rect -3248 70 -3215 116
rect -3169 70 -3136 116
rect -3248 68 -3136 70
rect -3080 116 -2968 118
rect -3080 70 -3047 116
rect -3001 70 -2968 116
rect -3080 68 -2968 70
rect -2912 116 -2800 118
rect -2912 70 -2879 116
rect -2833 70 -2800 116
rect -2912 68 -2800 70
rect -2744 116 -2632 118
rect -2744 70 -2711 116
rect -2665 70 -2632 116
rect -2744 68 -2632 70
rect -2576 116 -2464 118
rect -2576 70 -2543 116
rect -2497 70 -2464 116
rect -2576 68 -2464 70
rect -2408 116 -2296 118
rect -2408 70 -2375 116
rect -2329 70 -2296 116
rect -2408 68 -2296 70
rect -2240 116 -2128 118
rect -2240 70 -2207 116
rect -2161 70 -2128 116
rect -2240 68 -2128 70
rect -2072 116 -1960 118
rect -2072 70 -2039 116
rect -1993 70 -1960 116
rect -2072 68 -1960 70
rect -1904 116 -1792 118
rect -1904 70 -1871 116
rect -1825 70 -1792 116
rect -1904 68 -1792 70
rect -1736 116 -1624 118
rect -1736 70 -1703 116
rect -1657 70 -1624 116
rect -1736 68 -1624 70
rect -1568 116 -1456 118
rect -1568 70 -1535 116
rect -1489 70 -1456 116
rect -1568 68 -1456 70
rect -1400 116 -1288 118
rect -1400 70 -1367 116
rect -1321 70 -1288 116
rect -1400 68 -1288 70
rect -1232 116 -1120 118
rect -1232 70 -1199 116
rect -1153 70 -1120 116
rect -1232 68 -1120 70
rect -1064 116 -952 118
rect -1064 70 -1031 116
rect -985 70 -952 116
rect -1064 68 -952 70
rect -896 116 -784 118
rect -896 70 -863 116
rect -817 70 -784 116
rect -896 68 -784 70
rect -728 116 -616 118
rect -728 70 -695 116
rect -649 70 -616 116
rect -728 68 -616 70
rect -560 116 -448 118
rect -560 70 -527 116
rect -481 70 -448 116
rect -560 68 -448 70
rect -392 116 -280 118
rect -392 70 -359 116
rect -313 70 -280 116
rect -392 68 -280 70
rect -224 116 -112 118
rect -224 70 -191 116
rect -145 70 -112 116
rect -224 68 -112 70
rect -56 116 56 118
rect -56 70 -23 116
rect 23 70 56 116
rect -56 68 56 70
rect 112 116 224 118
rect 112 70 145 116
rect 191 70 224 116
rect 112 68 224 70
rect 280 116 392 118
rect 280 70 313 116
rect 359 70 392 116
rect 280 68 392 70
rect 448 116 560 118
rect 448 70 481 116
rect 527 70 560 116
rect 448 68 560 70
rect 616 116 728 118
rect 616 70 649 116
rect 695 70 728 116
rect 616 68 728 70
rect 784 116 896 118
rect 784 70 817 116
rect 863 70 896 116
rect 784 68 896 70
rect 952 116 1064 118
rect 952 70 985 116
rect 1031 70 1064 116
rect 952 68 1064 70
rect 1120 116 1232 118
rect 1120 70 1153 116
rect 1199 70 1232 116
rect 1120 68 1232 70
rect 1288 116 1400 118
rect 1288 70 1321 116
rect 1367 70 1400 116
rect 1288 68 1400 70
rect 1456 116 1568 118
rect 1456 70 1489 116
rect 1535 70 1568 116
rect 1456 68 1568 70
rect 1624 116 1736 118
rect 1624 70 1657 116
rect 1703 70 1736 116
rect 1624 68 1736 70
rect 1792 116 1904 118
rect 1792 70 1825 116
rect 1871 70 1904 116
rect 1792 68 1904 70
rect 1960 116 2072 118
rect 1960 70 1993 116
rect 2039 70 2072 116
rect 1960 68 2072 70
rect 2128 116 2240 118
rect 2128 70 2161 116
rect 2207 70 2240 116
rect 2128 68 2240 70
rect 2296 116 2408 118
rect 2296 70 2329 116
rect 2375 70 2408 116
rect 2296 68 2408 70
rect 2464 116 2576 118
rect 2464 70 2497 116
rect 2543 70 2576 116
rect 2464 68 2576 70
rect 2632 116 2744 118
rect 2632 70 2665 116
rect 2711 70 2744 116
rect 2632 68 2744 70
rect 2800 116 2912 118
rect 2800 70 2833 116
rect 2879 70 2912 116
rect 2800 68 2912 70
rect 2968 116 3080 118
rect 2968 70 3001 116
rect 3047 70 3080 116
rect 2968 68 3080 70
rect 3136 116 3248 118
rect 3136 70 3169 116
rect 3215 70 3248 116
rect 3136 68 3248 70
rect 3304 116 3396 118
rect 3304 70 3337 116
rect 3383 70 3396 116
rect 3304 68 3396 70
rect -3396 57 -3324 68
rect -3228 57 -3156 68
rect -3060 57 -2988 68
rect -2892 57 -2820 68
rect -2724 57 -2652 68
rect -2556 57 -2484 68
rect -2388 57 -2316 68
rect -2220 57 -2148 68
rect -2052 57 -1980 68
rect -1884 57 -1812 68
rect -1716 57 -1644 68
rect -1548 57 -1476 68
rect -1380 57 -1308 68
rect -1212 57 -1140 68
rect -1044 57 -972 68
rect -876 57 -804 68
rect -708 57 -636 68
rect -540 57 -468 68
rect -372 57 -300 68
rect -204 57 -132 68
rect -36 57 36 68
rect 132 57 204 68
rect 300 57 372 68
rect 468 57 540 68
rect 636 57 708 68
rect 804 57 876 68
rect 972 57 1044 68
rect 1140 57 1212 68
rect 1308 57 1380 68
rect 1476 57 1548 68
rect 1644 57 1716 68
rect 1812 57 1884 68
rect 1980 57 2052 68
rect 2148 57 2220 68
rect 2316 57 2388 68
rect 2484 57 2556 68
rect 2652 57 2724 68
rect 2820 57 2892 68
rect 2988 57 3060 68
rect 3156 57 3228 68
rect 3324 57 3396 68
rect -3396 -68 -3324 -57
rect -3228 -68 -3156 -57
rect -3060 -68 -2988 -57
rect -2892 -68 -2820 -57
rect -2724 -68 -2652 -57
rect -2556 -68 -2484 -57
rect -2388 -68 -2316 -57
rect -2220 -68 -2148 -57
rect -2052 -68 -1980 -57
rect -1884 -68 -1812 -57
rect -1716 -68 -1644 -57
rect -1548 -68 -1476 -57
rect -1380 -68 -1308 -57
rect -1212 -68 -1140 -57
rect -1044 -68 -972 -57
rect -876 -68 -804 -57
rect -708 -68 -636 -57
rect -540 -68 -468 -57
rect -372 -68 -300 -57
rect -204 -68 -132 -57
rect -36 -68 36 -57
rect 132 -68 204 -57
rect 300 -68 372 -57
rect 468 -68 540 -57
rect 636 -68 708 -57
rect 804 -68 876 -57
rect 972 -68 1044 -57
rect 1140 -68 1212 -57
rect 1308 -68 1380 -57
rect 1476 -68 1548 -57
rect 1644 -68 1716 -57
rect 1812 -68 1884 -57
rect 1980 -68 2052 -57
rect 2148 -68 2220 -57
rect 2316 -68 2388 -57
rect 2484 -68 2556 -57
rect 2652 -68 2724 -57
rect 2820 -68 2892 -57
rect 2988 -68 3060 -57
rect 3156 -68 3228 -57
rect 3324 -68 3396 -57
rect -3396 -70 -3304 -68
rect -3396 -116 -3383 -70
rect -3337 -116 -3304 -70
rect -3396 -118 -3304 -116
rect -3248 -70 -3136 -68
rect -3248 -116 -3215 -70
rect -3169 -116 -3136 -70
rect -3248 -118 -3136 -116
rect -3080 -70 -2968 -68
rect -3080 -116 -3047 -70
rect -3001 -116 -2968 -70
rect -3080 -118 -2968 -116
rect -2912 -70 -2800 -68
rect -2912 -116 -2879 -70
rect -2833 -116 -2800 -70
rect -2912 -118 -2800 -116
rect -2744 -70 -2632 -68
rect -2744 -116 -2711 -70
rect -2665 -116 -2632 -70
rect -2744 -118 -2632 -116
rect -2576 -70 -2464 -68
rect -2576 -116 -2543 -70
rect -2497 -116 -2464 -70
rect -2576 -118 -2464 -116
rect -2408 -70 -2296 -68
rect -2408 -116 -2375 -70
rect -2329 -116 -2296 -70
rect -2408 -118 -2296 -116
rect -2240 -70 -2128 -68
rect -2240 -116 -2207 -70
rect -2161 -116 -2128 -70
rect -2240 -118 -2128 -116
rect -2072 -70 -1960 -68
rect -2072 -116 -2039 -70
rect -1993 -116 -1960 -70
rect -2072 -118 -1960 -116
rect -1904 -70 -1792 -68
rect -1904 -116 -1871 -70
rect -1825 -116 -1792 -70
rect -1904 -118 -1792 -116
rect -1736 -70 -1624 -68
rect -1736 -116 -1703 -70
rect -1657 -116 -1624 -70
rect -1736 -118 -1624 -116
rect -1568 -70 -1456 -68
rect -1568 -116 -1535 -70
rect -1489 -116 -1456 -70
rect -1568 -118 -1456 -116
rect -1400 -70 -1288 -68
rect -1400 -116 -1367 -70
rect -1321 -116 -1288 -70
rect -1400 -118 -1288 -116
rect -1232 -70 -1120 -68
rect -1232 -116 -1199 -70
rect -1153 -116 -1120 -70
rect -1232 -118 -1120 -116
rect -1064 -70 -952 -68
rect -1064 -116 -1031 -70
rect -985 -116 -952 -70
rect -1064 -118 -952 -116
rect -896 -70 -784 -68
rect -896 -116 -863 -70
rect -817 -116 -784 -70
rect -896 -118 -784 -116
rect -728 -70 -616 -68
rect -728 -116 -695 -70
rect -649 -116 -616 -70
rect -728 -118 -616 -116
rect -560 -70 -448 -68
rect -560 -116 -527 -70
rect -481 -116 -448 -70
rect -560 -118 -448 -116
rect -392 -70 -280 -68
rect -392 -116 -359 -70
rect -313 -116 -280 -70
rect -392 -118 -280 -116
rect -224 -70 -112 -68
rect -224 -116 -191 -70
rect -145 -116 -112 -70
rect -224 -118 -112 -116
rect -56 -70 56 -68
rect -56 -116 -23 -70
rect 23 -116 56 -70
rect -56 -118 56 -116
rect 112 -70 224 -68
rect 112 -116 145 -70
rect 191 -116 224 -70
rect 112 -118 224 -116
rect 280 -70 392 -68
rect 280 -116 313 -70
rect 359 -116 392 -70
rect 280 -118 392 -116
rect 448 -70 560 -68
rect 448 -116 481 -70
rect 527 -116 560 -70
rect 448 -118 560 -116
rect 616 -70 728 -68
rect 616 -116 649 -70
rect 695 -116 728 -70
rect 616 -118 728 -116
rect 784 -70 896 -68
rect 784 -116 817 -70
rect 863 -116 896 -70
rect 784 -118 896 -116
rect 952 -70 1064 -68
rect 952 -116 985 -70
rect 1031 -116 1064 -70
rect 952 -118 1064 -116
rect 1120 -70 1232 -68
rect 1120 -116 1153 -70
rect 1199 -116 1232 -70
rect 1120 -118 1232 -116
rect 1288 -70 1400 -68
rect 1288 -116 1321 -70
rect 1367 -116 1400 -70
rect 1288 -118 1400 -116
rect 1456 -70 1568 -68
rect 1456 -116 1489 -70
rect 1535 -116 1568 -70
rect 1456 -118 1568 -116
rect 1624 -70 1736 -68
rect 1624 -116 1657 -70
rect 1703 -116 1736 -70
rect 1624 -118 1736 -116
rect 1792 -70 1904 -68
rect 1792 -116 1825 -70
rect 1871 -116 1904 -70
rect 1792 -118 1904 -116
rect 1960 -70 2072 -68
rect 1960 -116 1993 -70
rect 2039 -116 2072 -70
rect 1960 -118 2072 -116
rect 2128 -70 2240 -68
rect 2128 -116 2161 -70
rect 2207 -116 2240 -70
rect 2128 -118 2240 -116
rect 2296 -70 2408 -68
rect 2296 -116 2329 -70
rect 2375 -116 2408 -70
rect 2296 -118 2408 -116
rect 2464 -70 2576 -68
rect 2464 -116 2497 -70
rect 2543 -116 2576 -70
rect 2464 -118 2576 -116
rect 2632 -70 2744 -68
rect 2632 -116 2665 -70
rect 2711 -116 2744 -70
rect 2632 -118 2744 -116
rect 2800 -70 2912 -68
rect 2800 -116 2833 -70
rect 2879 -116 2912 -70
rect 2800 -118 2912 -116
rect 2968 -70 3080 -68
rect 2968 -116 3001 -70
rect 3047 -116 3080 -70
rect 2968 -118 3080 -116
rect 3136 -70 3248 -68
rect 3136 -116 3169 -70
rect 3215 -116 3248 -70
rect 3136 -118 3248 -116
rect 3304 -70 3396 -68
rect 3304 -116 3337 -70
rect 3383 -116 3396 -70
rect 3304 -118 3396 -116
rect -3396 -129 -3324 -118
rect -3228 -129 -3156 -118
rect -3060 -129 -2988 -118
rect -2892 -129 -2820 -118
rect -2724 -129 -2652 -118
rect -2556 -129 -2484 -118
rect -2388 -129 -2316 -118
rect -2220 -129 -2148 -118
rect -2052 -129 -1980 -118
rect -1884 -129 -1812 -118
rect -1716 -129 -1644 -118
rect -1548 -129 -1476 -118
rect -1380 -129 -1308 -118
rect -1212 -129 -1140 -118
rect -1044 -129 -972 -118
rect -876 -129 -804 -118
rect -708 -129 -636 -118
rect -540 -129 -468 -118
rect -372 -129 -300 -118
rect -204 -129 -132 -118
rect -36 -129 36 -118
rect 132 -129 204 -118
rect 300 -129 372 -118
rect 468 -129 540 -118
rect 636 -129 708 -118
rect 804 -129 876 -118
rect 972 -129 1044 -118
rect 1140 -129 1212 -118
rect 1308 -129 1380 -118
rect 1476 -129 1548 -118
rect 1644 -129 1716 -118
rect 1812 -129 1884 -118
rect 1980 -129 2052 -118
rect 2148 -129 2220 -118
rect 2316 -129 2388 -118
rect 2484 -129 2556 -118
rect 2652 -129 2724 -118
rect 2820 -129 2892 -118
rect 2988 -129 3060 -118
rect 3156 -129 3228 -118
rect 3324 -129 3396 -118
rect -3396 -254 -3324 -243
rect -3228 -254 -3156 -243
rect -3060 -254 -2988 -243
rect -2892 -254 -2820 -243
rect -2724 -254 -2652 -243
rect -2556 -254 -2484 -243
rect -2388 -254 -2316 -243
rect -2220 -254 -2148 -243
rect -2052 -254 -1980 -243
rect -1884 -254 -1812 -243
rect -1716 -254 -1644 -243
rect -1548 -254 -1476 -243
rect -1380 -254 -1308 -243
rect -1212 -254 -1140 -243
rect -1044 -254 -972 -243
rect -876 -254 -804 -243
rect -708 -254 -636 -243
rect -540 -254 -468 -243
rect -372 -254 -300 -243
rect -204 -254 -132 -243
rect -36 -254 36 -243
rect 132 -254 204 -243
rect 300 -254 372 -243
rect 468 -254 540 -243
rect 636 -254 708 -243
rect 804 -254 876 -243
rect 972 -254 1044 -243
rect 1140 -254 1212 -243
rect 1308 -254 1380 -243
rect 1476 -254 1548 -243
rect 1644 -254 1716 -243
rect 1812 -254 1884 -243
rect 1980 -254 2052 -243
rect 2148 -254 2220 -243
rect 2316 -254 2388 -243
rect 2484 -254 2556 -243
rect 2652 -254 2724 -243
rect 2820 -254 2892 -243
rect 2988 -254 3060 -243
rect 3156 -254 3228 -243
rect 3324 -254 3396 -243
rect -3396 -256 -3304 -254
rect -3396 -302 -3383 -256
rect -3337 -302 -3304 -256
rect -3396 -304 -3304 -302
rect -3248 -256 -3136 -254
rect -3248 -302 -3215 -256
rect -3169 -302 -3136 -256
rect -3248 -304 -3136 -302
rect -3080 -256 -2968 -254
rect -3080 -302 -3047 -256
rect -3001 -302 -2968 -256
rect -3080 -304 -2968 -302
rect -2912 -256 -2800 -254
rect -2912 -302 -2879 -256
rect -2833 -302 -2800 -256
rect -2912 -304 -2800 -302
rect -2744 -256 -2632 -254
rect -2744 -302 -2711 -256
rect -2665 -302 -2632 -256
rect -2744 -304 -2632 -302
rect -2576 -256 -2464 -254
rect -2576 -302 -2543 -256
rect -2497 -302 -2464 -256
rect -2576 -304 -2464 -302
rect -2408 -256 -2296 -254
rect -2408 -302 -2375 -256
rect -2329 -302 -2296 -256
rect -2408 -304 -2296 -302
rect -2240 -256 -2128 -254
rect -2240 -302 -2207 -256
rect -2161 -302 -2128 -256
rect -2240 -304 -2128 -302
rect -2072 -256 -1960 -254
rect -2072 -302 -2039 -256
rect -1993 -302 -1960 -256
rect -2072 -304 -1960 -302
rect -1904 -256 -1792 -254
rect -1904 -302 -1871 -256
rect -1825 -302 -1792 -256
rect -1904 -304 -1792 -302
rect -1736 -256 -1624 -254
rect -1736 -302 -1703 -256
rect -1657 -302 -1624 -256
rect -1736 -304 -1624 -302
rect -1568 -256 -1456 -254
rect -1568 -302 -1535 -256
rect -1489 -302 -1456 -256
rect -1568 -304 -1456 -302
rect -1400 -256 -1288 -254
rect -1400 -302 -1367 -256
rect -1321 -302 -1288 -256
rect -1400 -304 -1288 -302
rect -1232 -256 -1120 -254
rect -1232 -302 -1199 -256
rect -1153 -302 -1120 -256
rect -1232 -304 -1120 -302
rect -1064 -256 -952 -254
rect -1064 -302 -1031 -256
rect -985 -302 -952 -256
rect -1064 -304 -952 -302
rect -896 -256 -784 -254
rect -896 -302 -863 -256
rect -817 -302 -784 -256
rect -896 -304 -784 -302
rect -728 -256 -616 -254
rect -728 -302 -695 -256
rect -649 -302 -616 -256
rect -728 -304 -616 -302
rect -560 -256 -448 -254
rect -560 -302 -527 -256
rect -481 -302 -448 -256
rect -560 -304 -448 -302
rect -392 -256 -280 -254
rect -392 -302 -359 -256
rect -313 -302 -280 -256
rect -392 -304 -280 -302
rect -224 -256 -112 -254
rect -224 -302 -191 -256
rect -145 -302 -112 -256
rect -224 -304 -112 -302
rect -56 -256 56 -254
rect -56 -302 -23 -256
rect 23 -302 56 -256
rect -56 -304 56 -302
rect 112 -256 224 -254
rect 112 -302 145 -256
rect 191 -302 224 -256
rect 112 -304 224 -302
rect 280 -256 392 -254
rect 280 -302 313 -256
rect 359 -302 392 -256
rect 280 -304 392 -302
rect 448 -256 560 -254
rect 448 -302 481 -256
rect 527 -302 560 -256
rect 448 -304 560 -302
rect 616 -256 728 -254
rect 616 -302 649 -256
rect 695 -302 728 -256
rect 616 -304 728 -302
rect 784 -256 896 -254
rect 784 -302 817 -256
rect 863 -302 896 -256
rect 784 -304 896 -302
rect 952 -256 1064 -254
rect 952 -302 985 -256
rect 1031 -302 1064 -256
rect 952 -304 1064 -302
rect 1120 -256 1232 -254
rect 1120 -302 1153 -256
rect 1199 -302 1232 -256
rect 1120 -304 1232 -302
rect 1288 -256 1400 -254
rect 1288 -302 1321 -256
rect 1367 -302 1400 -256
rect 1288 -304 1400 -302
rect 1456 -256 1568 -254
rect 1456 -302 1489 -256
rect 1535 -302 1568 -256
rect 1456 -304 1568 -302
rect 1624 -256 1736 -254
rect 1624 -302 1657 -256
rect 1703 -302 1736 -256
rect 1624 -304 1736 -302
rect 1792 -256 1904 -254
rect 1792 -302 1825 -256
rect 1871 -302 1904 -256
rect 1792 -304 1904 -302
rect 1960 -256 2072 -254
rect 1960 -302 1993 -256
rect 2039 -302 2072 -256
rect 1960 -304 2072 -302
rect 2128 -256 2240 -254
rect 2128 -302 2161 -256
rect 2207 -302 2240 -256
rect 2128 -304 2240 -302
rect 2296 -256 2408 -254
rect 2296 -302 2329 -256
rect 2375 -302 2408 -256
rect 2296 -304 2408 -302
rect 2464 -256 2576 -254
rect 2464 -302 2497 -256
rect 2543 -302 2576 -256
rect 2464 -304 2576 -302
rect 2632 -256 2744 -254
rect 2632 -302 2665 -256
rect 2711 -302 2744 -256
rect 2632 -304 2744 -302
rect 2800 -256 2912 -254
rect 2800 -302 2833 -256
rect 2879 -302 2912 -256
rect 2800 -304 2912 -302
rect 2968 -256 3080 -254
rect 2968 -302 3001 -256
rect 3047 -302 3080 -256
rect 2968 -304 3080 -302
rect 3136 -256 3248 -254
rect 3136 -302 3169 -256
rect 3215 -302 3248 -256
rect 3136 -304 3248 -302
rect 3304 -256 3396 -254
rect 3304 -302 3337 -256
rect 3383 -302 3396 -256
rect 3304 -304 3396 -302
rect -3396 -315 -3324 -304
rect -3228 -315 -3156 -304
rect -3060 -315 -2988 -304
rect -2892 -315 -2820 -304
rect -2724 -315 -2652 -304
rect -2556 -315 -2484 -304
rect -2388 -315 -2316 -304
rect -2220 -315 -2148 -304
rect -2052 -315 -1980 -304
rect -1884 -315 -1812 -304
rect -1716 -315 -1644 -304
rect -1548 -315 -1476 -304
rect -1380 -315 -1308 -304
rect -1212 -315 -1140 -304
rect -1044 -315 -972 -304
rect -876 -315 -804 -304
rect -708 -315 -636 -304
rect -540 -315 -468 -304
rect -372 -315 -300 -304
rect -204 -315 -132 -304
rect -36 -315 36 -304
rect 132 -315 204 -304
rect 300 -315 372 -304
rect 468 -315 540 -304
rect 636 -315 708 -304
rect 804 -315 876 -304
rect 972 -315 1044 -304
rect 1140 -315 1212 -304
rect 1308 -315 1380 -304
rect 1476 -315 1548 -304
rect 1644 -315 1716 -304
rect 1812 -315 1884 -304
rect 1980 -315 2052 -304
rect 2148 -315 2220 -304
rect 2316 -315 2388 -304
rect 2484 -315 2556 -304
rect 2652 -315 2724 -304
rect 2820 -315 2892 -304
rect 2988 -315 3060 -304
rect 3156 -315 3228 -304
rect 3324 -315 3396 -304
rect -3396 -440 -3324 -429
rect -3228 -440 -3156 -429
rect -3060 -440 -2988 -429
rect -2892 -440 -2820 -429
rect -2724 -440 -2652 -429
rect -2556 -440 -2484 -429
rect -2388 -440 -2316 -429
rect -2220 -440 -2148 -429
rect -2052 -440 -1980 -429
rect -1884 -440 -1812 -429
rect -1716 -440 -1644 -429
rect -1548 -440 -1476 -429
rect -1380 -440 -1308 -429
rect -1212 -440 -1140 -429
rect -1044 -440 -972 -429
rect -876 -440 -804 -429
rect -708 -440 -636 -429
rect -540 -440 -468 -429
rect -372 -440 -300 -429
rect -204 -440 -132 -429
rect -36 -440 36 -429
rect 132 -440 204 -429
rect 300 -440 372 -429
rect 468 -440 540 -429
rect 636 -440 708 -429
rect 804 -440 876 -429
rect 972 -440 1044 -429
rect 1140 -440 1212 -429
rect 1308 -440 1380 -429
rect 1476 -440 1548 -429
rect 1644 -440 1716 -429
rect 1812 -440 1884 -429
rect 1980 -440 2052 -429
rect 2148 -440 2220 -429
rect 2316 -440 2388 -429
rect 2484 -440 2556 -429
rect 2652 -440 2724 -429
rect 2820 -440 2892 -429
rect 2988 -440 3060 -429
rect 3156 -440 3228 -429
rect 3324 -440 3396 -429
rect -3396 -442 -3304 -440
rect -3396 -488 -3383 -442
rect -3337 -488 -3304 -442
rect -3396 -490 -3304 -488
rect -3248 -442 -3136 -440
rect -3248 -488 -3215 -442
rect -3169 -488 -3136 -442
rect -3248 -490 -3136 -488
rect -3080 -442 -2968 -440
rect -3080 -488 -3047 -442
rect -3001 -488 -2968 -442
rect -3080 -490 -2968 -488
rect -2912 -442 -2800 -440
rect -2912 -488 -2879 -442
rect -2833 -488 -2800 -442
rect -2912 -490 -2800 -488
rect -2744 -442 -2632 -440
rect -2744 -488 -2711 -442
rect -2665 -488 -2632 -442
rect -2744 -490 -2632 -488
rect -2576 -442 -2464 -440
rect -2576 -488 -2543 -442
rect -2497 -488 -2464 -442
rect -2576 -490 -2464 -488
rect -2408 -442 -2296 -440
rect -2408 -488 -2375 -442
rect -2329 -488 -2296 -442
rect -2408 -490 -2296 -488
rect -2240 -442 -2128 -440
rect -2240 -488 -2207 -442
rect -2161 -488 -2128 -442
rect -2240 -490 -2128 -488
rect -2072 -442 -1960 -440
rect -2072 -488 -2039 -442
rect -1993 -488 -1960 -442
rect -2072 -490 -1960 -488
rect -1904 -442 -1792 -440
rect -1904 -488 -1871 -442
rect -1825 -488 -1792 -442
rect -1904 -490 -1792 -488
rect -1736 -442 -1624 -440
rect -1736 -488 -1703 -442
rect -1657 -488 -1624 -442
rect -1736 -490 -1624 -488
rect -1568 -442 -1456 -440
rect -1568 -488 -1535 -442
rect -1489 -488 -1456 -442
rect -1568 -490 -1456 -488
rect -1400 -442 -1288 -440
rect -1400 -488 -1367 -442
rect -1321 -488 -1288 -442
rect -1400 -490 -1288 -488
rect -1232 -442 -1120 -440
rect -1232 -488 -1199 -442
rect -1153 -488 -1120 -442
rect -1232 -490 -1120 -488
rect -1064 -442 -952 -440
rect -1064 -488 -1031 -442
rect -985 -488 -952 -442
rect -1064 -490 -952 -488
rect -896 -442 -784 -440
rect -896 -488 -863 -442
rect -817 -488 -784 -442
rect -896 -490 -784 -488
rect -728 -442 -616 -440
rect -728 -488 -695 -442
rect -649 -488 -616 -442
rect -728 -490 -616 -488
rect -560 -442 -448 -440
rect -560 -488 -527 -442
rect -481 -488 -448 -442
rect -560 -490 -448 -488
rect -392 -442 -280 -440
rect -392 -488 -359 -442
rect -313 -488 -280 -442
rect -392 -490 -280 -488
rect -224 -442 -112 -440
rect -224 -488 -191 -442
rect -145 -488 -112 -442
rect -224 -490 -112 -488
rect -56 -442 56 -440
rect -56 -488 -23 -442
rect 23 -488 56 -442
rect -56 -490 56 -488
rect 112 -442 224 -440
rect 112 -488 145 -442
rect 191 -488 224 -442
rect 112 -490 224 -488
rect 280 -442 392 -440
rect 280 -488 313 -442
rect 359 -488 392 -442
rect 280 -490 392 -488
rect 448 -442 560 -440
rect 448 -488 481 -442
rect 527 -488 560 -442
rect 448 -490 560 -488
rect 616 -442 728 -440
rect 616 -488 649 -442
rect 695 -488 728 -442
rect 616 -490 728 -488
rect 784 -442 896 -440
rect 784 -488 817 -442
rect 863 -488 896 -442
rect 784 -490 896 -488
rect 952 -442 1064 -440
rect 952 -488 985 -442
rect 1031 -488 1064 -442
rect 952 -490 1064 -488
rect 1120 -442 1232 -440
rect 1120 -488 1153 -442
rect 1199 -488 1232 -442
rect 1120 -490 1232 -488
rect 1288 -442 1400 -440
rect 1288 -488 1321 -442
rect 1367 -488 1400 -442
rect 1288 -490 1400 -488
rect 1456 -442 1568 -440
rect 1456 -488 1489 -442
rect 1535 -488 1568 -442
rect 1456 -490 1568 -488
rect 1624 -442 1736 -440
rect 1624 -488 1657 -442
rect 1703 -488 1736 -442
rect 1624 -490 1736 -488
rect 1792 -442 1904 -440
rect 1792 -488 1825 -442
rect 1871 -488 1904 -442
rect 1792 -490 1904 -488
rect 1960 -442 2072 -440
rect 1960 -488 1993 -442
rect 2039 -488 2072 -442
rect 1960 -490 2072 -488
rect 2128 -442 2240 -440
rect 2128 -488 2161 -442
rect 2207 -488 2240 -442
rect 2128 -490 2240 -488
rect 2296 -442 2408 -440
rect 2296 -488 2329 -442
rect 2375 -488 2408 -442
rect 2296 -490 2408 -488
rect 2464 -442 2576 -440
rect 2464 -488 2497 -442
rect 2543 -488 2576 -442
rect 2464 -490 2576 -488
rect 2632 -442 2744 -440
rect 2632 -488 2665 -442
rect 2711 -488 2744 -442
rect 2632 -490 2744 -488
rect 2800 -442 2912 -440
rect 2800 -488 2833 -442
rect 2879 -488 2912 -442
rect 2800 -490 2912 -488
rect 2968 -442 3080 -440
rect 2968 -488 3001 -442
rect 3047 -488 3080 -442
rect 2968 -490 3080 -488
rect 3136 -442 3248 -440
rect 3136 -488 3169 -442
rect 3215 -488 3248 -442
rect 3136 -490 3248 -488
rect 3304 -442 3396 -440
rect 3304 -488 3337 -442
rect 3383 -488 3396 -442
rect 3304 -490 3396 -488
rect -3396 -501 -3324 -490
rect -3228 -501 -3156 -490
rect -3060 -501 -2988 -490
rect -2892 -501 -2820 -490
rect -2724 -501 -2652 -490
rect -2556 -501 -2484 -490
rect -2388 -501 -2316 -490
rect -2220 -501 -2148 -490
rect -2052 -501 -1980 -490
rect -1884 -501 -1812 -490
rect -1716 -501 -1644 -490
rect -1548 -501 -1476 -490
rect -1380 -501 -1308 -490
rect -1212 -501 -1140 -490
rect -1044 -501 -972 -490
rect -876 -501 -804 -490
rect -708 -501 -636 -490
rect -540 -501 -468 -490
rect -372 -501 -300 -490
rect -204 -501 -132 -490
rect -36 -501 36 -490
rect 132 -501 204 -490
rect 300 -501 372 -490
rect 468 -501 540 -490
rect 636 -501 708 -490
rect 804 -501 876 -490
rect 972 -501 1044 -490
rect 1140 -501 1212 -490
rect 1308 -501 1380 -490
rect 1476 -501 1548 -490
rect 1644 -501 1716 -490
rect 1812 -501 1884 -490
rect 1980 -501 2052 -490
rect 2148 -501 2220 -490
rect 2316 -501 2388 -490
rect 2484 -501 2556 -490
rect 2652 -501 2724 -490
rect 2820 -501 2892 -490
rect 2988 -501 3060 -490
rect 3156 -501 3228 -490
rect 3324 -501 3396 -490
rect -3396 -626 -3324 -615
rect -3228 -626 -3156 -615
rect -3060 -626 -2988 -615
rect -2892 -626 -2820 -615
rect -2724 -626 -2652 -615
rect -2556 -626 -2484 -615
rect -2388 -626 -2316 -615
rect -2220 -626 -2148 -615
rect -2052 -626 -1980 -615
rect -1884 -626 -1812 -615
rect -1716 -626 -1644 -615
rect -1548 -626 -1476 -615
rect -1380 -626 -1308 -615
rect -1212 -626 -1140 -615
rect -1044 -626 -972 -615
rect -876 -626 -804 -615
rect -708 -626 -636 -615
rect -540 -626 -468 -615
rect -372 -626 -300 -615
rect -204 -626 -132 -615
rect -36 -626 36 -615
rect 132 -626 204 -615
rect 300 -626 372 -615
rect 468 -626 540 -615
rect 636 -626 708 -615
rect 804 -626 876 -615
rect 972 -626 1044 -615
rect 1140 -626 1212 -615
rect 1308 -626 1380 -615
rect 1476 -626 1548 -615
rect 1644 -626 1716 -615
rect 1812 -626 1884 -615
rect 1980 -626 2052 -615
rect 2148 -626 2220 -615
rect 2316 -626 2388 -615
rect 2484 -626 2556 -615
rect 2652 -626 2724 -615
rect 2820 -626 2892 -615
rect 2988 -626 3060 -615
rect 3156 -626 3228 -615
rect 3324 -626 3396 -615
rect -3396 -628 -3304 -626
rect -3396 -674 -3383 -628
rect -3337 -674 -3304 -628
rect -3396 -676 -3304 -674
rect -3248 -628 -3136 -626
rect -3248 -674 -3215 -628
rect -3169 -674 -3136 -628
rect -3248 -676 -3136 -674
rect -3080 -628 -2968 -626
rect -3080 -674 -3047 -628
rect -3001 -674 -2968 -628
rect -3080 -676 -2968 -674
rect -2912 -628 -2800 -626
rect -2912 -674 -2879 -628
rect -2833 -674 -2800 -628
rect -2912 -676 -2800 -674
rect -2744 -628 -2632 -626
rect -2744 -674 -2711 -628
rect -2665 -674 -2632 -628
rect -2744 -676 -2632 -674
rect -2576 -628 -2464 -626
rect -2576 -674 -2543 -628
rect -2497 -674 -2464 -628
rect -2576 -676 -2464 -674
rect -2408 -628 -2296 -626
rect -2408 -674 -2375 -628
rect -2329 -674 -2296 -628
rect -2408 -676 -2296 -674
rect -2240 -628 -2128 -626
rect -2240 -674 -2207 -628
rect -2161 -674 -2128 -628
rect -2240 -676 -2128 -674
rect -2072 -628 -1960 -626
rect -2072 -674 -2039 -628
rect -1993 -674 -1960 -628
rect -2072 -676 -1960 -674
rect -1904 -628 -1792 -626
rect -1904 -674 -1871 -628
rect -1825 -674 -1792 -628
rect -1904 -676 -1792 -674
rect -1736 -628 -1624 -626
rect -1736 -674 -1703 -628
rect -1657 -674 -1624 -628
rect -1736 -676 -1624 -674
rect -1568 -628 -1456 -626
rect -1568 -674 -1535 -628
rect -1489 -674 -1456 -628
rect -1568 -676 -1456 -674
rect -1400 -628 -1288 -626
rect -1400 -674 -1367 -628
rect -1321 -674 -1288 -628
rect -1400 -676 -1288 -674
rect -1232 -628 -1120 -626
rect -1232 -674 -1199 -628
rect -1153 -674 -1120 -628
rect -1232 -676 -1120 -674
rect -1064 -628 -952 -626
rect -1064 -674 -1031 -628
rect -985 -674 -952 -628
rect -1064 -676 -952 -674
rect -896 -628 -784 -626
rect -896 -674 -863 -628
rect -817 -674 -784 -628
rect -896 -676 -784 -674
rect -728 -628 -616 -626
rect -728 -674 -695 -628
rect -649 -674 -616 -628
rect -728 -676 -616 -674
rect -560 -628 -448 -626
rect -560 -674 -527 -628
rect -481 -674 -448 -628
rect -560 -676 -448 -674
rect -392 -628 -280 -626
rect -392 -674 -359 -628
rect -313 -674 -280 -628
rect -392 -676 -280 -674
rect -224 -628 -112 -626
rect -224 -674 -191 -628
rect -145 -674 -112 -628
rect -224 -676 -112 -674
rect -56 -628 56 -626
rect -56 -674 -23 -628
rect 23 -674 56 -628
rect -56 -676 56 -674
rect 112 -628 224 -626
rect 112 -674 145 -628
rect 191 -674 224 -628
rect 112 -676 224 -674
rect 280 -628 392 -626
rect 280 -674 313 -628
rect 359 -674 392 -628
rect 280 -676 392 -674
rect 448 -628 560 -626
rect 448 -674 481 -628
rect 527 -674 560 -628
rect 448 -676 560 -674
rect 616 -628 728 -626
rect 616 -674 649 -628
rect 695 -674 728 -628
rect 616 -676 728 -674
rect 784 -628 896 -626
rect 784 -674 817 -628
rect 863 -674 896 -628
rect 784 -676 896 -674
rect 952 -628 1064 -626
rect 952 -674 985 -628
rect 1031 -674 1064 -628
rect 952 -676 1064 -674
rect 1120 -628 1232 -626
rect 1120 -674 1153 -628
rect 1199 -674 1232 -628
rect 1120 -676 1232 -674
rect 1288 -628 1400 -626
rect 1288 -674 1321 -628
rect 1367 -674 1400 -628
rect 1288 -676 1400 -674
rect 1456 -628 1568 -626
rect 1456 -674 1489 -628
rect 1535 -674 1568 -628
rect 1456 -676 1568 -674
rect 1624 -628 1736 -626
rect 1624 -674 1657 -628
rect 1703 -674 1736 -628
rect 1624 -676 1736 -674
rect 1792 -628 1904 -626
rect 1792 -674 1825 -628
rect 1871 -674 1904 -628
rect 1792 -676 1904 -674
rect 1960 -628 2072 -626
rect 1960 -674 1993 -628
rect 2039 -674 2072 -628
rect 1960 -676 2072 -674
rect 2128 -628 2240 -626
rect 2128 -674 2161 -628
rect 2207 -674 2240 -628
rect 2128 -676 2240 -674
rect 2296 -628 2408 -626
rect 2296 -674 2329 -628
rect 2375 -674 2408 -628
rect 2296 -676 2408 -674
rect 2464 -628 2576 -626
rect 2464 -674 2497 -628
rect 2543 -674 2576 -628
rect 2464 -676 2576 -674
rect 2632 -628 2744 -626
rect 2632 -674 2665 -628
rect 2711 -674 2744 -628
rect 2632 -676 2744 -674
rect 2800 -628 2912 -626
rect 2800 -674 2833 -628
rect 2879 -674 2912 -628
rect 2800 -676 2912 -674
rect 2968 -628 3080 -626
rect 2968 -674 3001 -628
rect 3047 -674 3080 -628
rect 2968 -676 3080 -674
rect 3136 -628 3248 -626
rect 3136 -674 3169 -628
rect 3215 -674 3248 -628
rect 3136 -676 3248 -674
rect 3304 -628 3396 -626
rect 3304 -674 3337 -628
rect 3383 -674 3396 -628
rect 3304 -676 3396 -674
rect -3396 -687 -3324 -676
rect -3228 -687 -3156 -676
rect -3060 -687 -2988 -676
rect -2892 -687 -2820 -676
rect -2724 -687 -2652 -676
rect -2556 -687 -2484 -676
rect -2388 -687 -2316 -676
rect -2220 -687 -2148 -676
rect -2052 -687 -1980 -676
rect -1884 -687 -1812 -676
rect -1716 -687 -1644 -676
rect -1548 -687 -1476 -676
rect -1380 -687 -1308 -676
rect -1212 -687 -1140 -676
rect -1044 -687 -972 -676
rect -876 -687 -804 -676
rect -708 -687 -636 -676
rect -540 -687 -468 -676
rect -372 -687 -300 -676
rect -204 -687 -132 -676
rect -36 -687 36 -676
rect 132 -687 204 -676
rect 300 -687 372 -676
rect 468 -687 540 -676
rect 636 -687 708 -676
rect 804 -687 876 -676
rect 972 -687 1044 -676
rect 1140 -687 1212 -676
rect 1308 -687 1380 -676
rect 1476 -687 1548 -676
rect 1644 -687 1716 -676
rect 1812 -687 1884 -676
rect 1980 -687 2052 -676
rect 2148 -687 2220 -676
rect 2316 -687 2388 -676
rect 2484 -687 2556 -676
rect 2652 -687 2724 -676
rect 2820 -687 2892 -676
rect 2988 -687 3060 -676
rect 3156 -687 3228 -676
rect 3324 -687 3396 -676
<< ndiffc >>
rect -3383 628 -3337 674
rect -3215 628 -3169 674
rect -3047 628 -3001 674
rect -2879 628 -2833 674
rect -2711 628 -2665 674
rect -2543 628 -2497 674
rect -2375 628 -2329 674
rect -2207 628 -2161 674
rect -2039 628 -1993 674
rect -1871 628 -1825 674
rect -1703 628 -1657 674
rect -1535 628 -1489 674
rect -1367 628 -1321 674
rect -1199 628 -1153 674
rect -1031 628 -985 674
rect -863 628 -817 674
rect -695 628 -649 674
rect -527 628 -481 674
rect -359 628 -313 674
rect -191 628 -145 674
rect -23 628 23 674
rect 145 628 191 674
rect 313 628 359 674
rect 481 628 527 674
rect 649 628 695 674
rect 817 628 863 674
rect 985 628 1031 674
rect 1153 628 1199 674
rect 1321 628 1367 674
rect 1489 628 1535 674
rect 1657 628 1703 674
rect 1825 628 1871 674
rect 1993 628 2039 674
rect 2161 628 2207 674
rect 2329 628 2375 674
rect 2497 628 2543 674
rect 2665 628 2711 674
rect 2833 628 2879 674
rect 3001 628 3047 674
rect 3169 628 3215 674
rect 3337 628 3383 674
rect -3383 442 -3337 488
rect -3215 442 -3169 488
rect -3047 442 -3001 488
rect -2879 442 -2833 488
rect -2711 442 -2665 488
rect -2543 442 -2497 488
rect -2375 442 -2329 488
rect -2207 442 -2161 488
rect -2039 442 -1993 488
rect -1871 442 -1825 488
rect -1703 442 -1657 488
rect -1535 442 -1489 488
rect -1367 442 -1321 488
rect -1199 442 -1153 488
rect -1031 442 -985 488
rect -863 442 -817 488
rect -695 442 -649 488
rect -527 442 -481 488
rect -359 442 -313 488
rect -191 442 -145 488
rect -23 442 23 488
rect 145 442 191 488
rect 313 442 359 488
rect 481 442 527 488
rect 649 442 695 488
rect 817 442 863 488
rect 985 442 1031 488
rect 1153 442 1199 488
rect 1321 442 1367 488
rect 1489 442 1535 488
rect 1657 442 1703 488
rect 1825 442 1871 488
rect 1993 442 2039 488
rect 2161 442 2207 488
rect 2329 442 2375 488
rect 2497 442 2543 488
rect 2665 442 2711 488
rect 2833 442 2879 488
rect 3001 442 3047 488
rect 3169 442 3215 488
rect 3337 442 3383 488
rect -3383 256 -3337 302
rect -3215 256 -3169 302
rect -3047 256 -3001 302
rect -2879 256 -2833 302
rect -2711 256 -2665 302
rect -2543 256 -2497 302
rect -2375 256 -2329 302
rect -2207 256 -2161 302
rect -2039 256 -1993 302
rect -1871 256 -1825 302
rect -1703 256 -1657 302
rect -1535 256 -1489 302
rect -1367 256 -1321 302
rect -1199 256 -1153 302
rect -1031 256 -985 302
rect -863 256 -817 302
rect -695 256 -649 302
rect -527 256 -481 302
rect -359 256 -313 302
rect -191 256 -145 302
rect -23 256 23 302
rect 145 256 191 302
rect 313 256 359 302
rect 481 256 527 302
rect 649 256 695 302
rect 817 256 863 302
rect 985 256 1031 302
rect 1153 256 1199 302
rect 1321 256 1367 302
rect 1489 256 1535 302
rect 1657 256 1703 302
rect 1825 256 1871 302
rect 1993 256 2039 302
rect 2161 256 2207 302
rect 2329 256 2375 302
rect 2497 256 2543 302
rect 2665 256 2711 302
rect 2833 256 2879 302
rect 3001 256 3047 302
rect 3169 256 3215 302
rect 3337 256 3383 302
rect -3383 70 -3337 116
rect -3215 70 -3169 116
rect -3047 70 -3001 116
rect -2879 70 -2833 116
rect -2711 70 -2665 116
rect -2543 70 -2497 116
rect -2375 70 -2329 116
rect -2207 70 -2161 116
rect -2039 70 -1993 116
rect -1871 70 -1825 116
rect -1703 70 -1657 116
rect -1535 70 -1489 116
rect -1367 70 -1321 116
rect -1199 70 -1153 116
rect -1031 70 -985 116
rect -863 70 -817 116
rect -695 70 -649 116
rect -527 70 -481 116
rect -359 70 -313 116
rect -191 70 -145 116
rect -23 70 23 116
rect 145 70 191 116
rect 313 70 359 116
rect 481 70 527 116
rect 649 70 695 116
rect 817 70 863 116
rect 985 70 1031 116
rect 1153 70 1199 116
rect 1321 70 1367 116
rect 1489 70 1535 116
rect 1657 70 1703 116
rect 1825 70 1871 116
rect 1993 70 2039 116
rect 2161 70 2207 116
rect 2329 70 2375 116
rect 2497 70 2543 116
rect 2665 70 2711 116
rect 2833 70 2879 116
rect 3001 70 3047 116
rect 3169 70 3215 116
rect 3337 70 3383 116
rect -3383 -116 -3337 -70
rect -3215 -116 -3169 -70
rect -3047 -116 -3001 -70
rect -2879 -116 -2833 -70
rect -2711 -116 -2665 -70
rect -2543 -116 -2497 -70
rect -2375 -116 -2329 -70
rect -2207 -116 -2161 -70
rect -2039 -116 -1993 -70
rect -1871 -116 -1825 -70
rect -1703 -116 -1657 -70
rect -1535 -116 -1489 -70
rect -1367 -116 -1321 -70
rect -1199 -116 -1153 -70
rect -1031 -116 -985 -70
rect -863 -116 -817 -70
rect -695 -116 -649 -70
rect -527 -116 -481 -70
rect -359 -116 -313 -70
rect -191 -116 -145 -70
rect -23 -116 23 -70
rect 145 -116 191 -70
rect 313 -116 359 -70
rect 481 -116 527 -70
rect 649 -116 695 -70
rect 817 -116 863 -70
rect 985 -116 1031 -70
rect 1153 -116 1199 -70
rect 1321 -116 1367 -70
rect 1489 -116 1535 -70
rect 1657 -116 1703 -70
rect 1825 -116 1871 -70
rect 1993 -116 2039 -70
rect 2161 -116 2207 -70
rect 2329 -116 2375 -70
rect 2497 -116 2543 -70
rect 2665 -116 2711 -70
rect 2833 -116 2879 -70
rect 3001 -116 3047 -70
rect 3169 -116 3215 -70
rect 3337 -116 3383 -70
rect -3383 -302 -3337 -256
rect -3215 -302 -3169 -256
rect -3047 -302 -3001 -256
rect -2879 -302 -2833 -256
rect -2711 -302 -2665 -256
rect -2543 -302 -2497 -256
rect -2375 -302 -2329 -256
rect -2207 -302 -2161 -256
rect -2039 -302 -1993 -256
rect -1871 -302 -1825 -256
rect -1703 -302 -1657 -256
rect -1535 -302 -1489 -256
rect -1367 -302 -1321 -256
rect -1199 -302 -1153 -256
rect -1031 -302 -985 -256
rect -863 -302 -817 -256
rect -695 -302 -649 -256
rect -527 -302 -481 -256
rect -359 -302 -313 -256
rect -191 -302 -145 -256
rect -23 -302 23 -256
rect 145 -302 191 -256
rect 313 -302 359 -256
rect 481 -302 527 -256
rect 649 -302 695 -256
rect 817 -302 863 -256
rect 985 -302 1031 -256
rect 1153 -302 1199 -256
rect 1321 -302 1367 -256
rect 1489 -302 1535 -256
rect 1657 -302 1703 -256
rect 1825 -302 1871 -256
rect 1993 -302 2039 -256
rect 2161 -302 2207 -256
rect 2329 -302 2375 -256
rect 2497 -302 2543 -256
rect 2665 -302 2711 -256
rect 2833 -302 2879 -256
rect 3001 -302 3047 -256
rect 3169 -302 3215 -256
rect 3337 -302 3383 -256
rect -3383 -488 -3337 -442
rect -3215 -488 -3169 -442
rect -3047 -488 -3001 -442
rect -2879 -488 -2833 -442
rect -2711 -488 -2665 -442
rect -2543 -488 -2497 -442
rect -2375 -488 -2329 -442
rect -2207 -488 -2161 -442
rect -2039 -488 -1993 -442
rect -1871 -488 -1825 -442
rect -1703 -488 -1657 -442
rect -1535 -488 -1489 -442
rect -1367 -488 -1321 -442
rect -1199 -488 -1153 -442
rect -1031 -488 -985 -442
rect -863 -488 -817 -442
rect -695 -488 -649 -442
rect -527 -488 -481 -442
rect -359 -488 -313 -442
rect -191 -488 -145 -442
rect -23 -488 23 -442
rect 145 -488 191 -442
rect 313 -488 359 -442
rect 481 -488 527 -442
rect 649 -488 695 -442
rect 817 -488 863 -442
rect 985 -488 1031 -442
rect 1153 -488 1199 -442
rect 1321 -488 1367 -442
rect 1489 -488 1535 -442
rect 1657 -488 1703 -442
rect 1825 -488 1871 -442
rect 1993 -488 2039 -442
rect 2161 -488 2207 -442
rect 2329 -488 2375 -442
rect 2497 -488 2543 -442
rect 2665 -488 2711 -442
rect 2833 -488 2879 -442
rect 3001 -488 3047 -442
rect 3169 -488 3215 -442
rect 3337 -488 3383 -442
rect -3383 -674 -3337 -628
rect -3215 -674 -3169 -628
rect -3047 -674 -3001 -628
rect -2879 -674 -2833 -628
rect -2711 -674 -2665 -628
rect -2543 -674 -2497 -628
rect -2375 -674 -2329 -628
rect -2207 -674 -2161 -628
rect -2039 -674 -1993 -628
rect -1871 -674 -1825 -628
rect -1703 -674 -1657 -628
rect -1535 -674 -1489 -628
rect -1367 -674 -1321 -628
rect -1199 -674 -1153 -628
rect -1031 -674 -985 -628
rect -863 -674 -817 -628
rect -695 -674 -649 -628
rect -527 -674 -481 -628
rect -359 -674 -313 -628
rect -191 -674 -145 -628
rect -23 -674 23 -628
rect 145 -674 191 -628
rect 313 -674 359 -628
rect 481 -674 527 -628
rect 649 -674 695 -628
rect 817 -674 863 -628
rect 985 -674 1031 -628
rect 1153 -674 1199 -628
rect 1321 -674 1367 -628
rect 1489 -674 1535 -628
rect 1657 -674 1703 -628
rect 1825 -674 1871 -628
rect 1993 -674 2039 -628
rect 2161 -674 2207 -628
rect 2329 -674 2375 -628
rect 2497 -674 2543 -628
rect 2665 -674 2711 -628
rect 2833 -674 2879 -628
rect 3001 -674 3047 -628
rect 3169 -674 3215 -628
rect 3337 -674 3383 -628
<< polysilicon >>
rect -3304 676 -3248 720
rect -3136 676 -3080 720
rect -2968 676 -2912 720
rect -2800 676 -2744 720
rect -2632 676 -2576 720
rect -2464 676 -2408 720
rect -2296 676 -2240 720
rect -2128 676 -2072 720
rect -1960 676 -1904 720
rect -1792 676 -1736 720
rect -1624 676 -1568 720
rect -1456 676 -1400 720
rect -1288 676 -1232 720
rect -1120 676 -1064 720
rect -952 676 -896 720
rect -784 676 -728 720
rect -616 676 -560 720
rect -448 676 -392 720
rect -280 676 -224 720
rect -112 676 -56 720
rect 56 676 112 720
rect 224 676 280 720
rect 392 676 448 720
rect 560 676 616 720
rect 728 676 784 720
rect 896 676 952 720
rect 1064 676 1120 720
rect 1232 676 1288 720
rect 1400 676 1456 720
rect 1568 676 1624 720
rect 1736 676 1792 720
rect 1904 676 1960 720
rect 2072 676 2128 720
rect 2240 676 2296 720
rect 2408 676 2464 720
rect 2576 676 2632 720
rect 2744 676 2800 720
rect 2912 676 2968 720
rect 3080 676 3136 720
rect 3248 676 3304 720
rect -3304 582 -3248 626
rect -3136 582 -3080 626
rect -2968 582 -2912 626
rect -2800 582 -2744 626
rect -2632 582 -2576 626
rect -2464 582 -2408 626
rect -2296 582 -2240 626
rect -2128 582 -2072 626
rect -1960 582 -1904 626
rect -1792 582 -1736 626
rect -1624 582 -1568 626
rect -1456 582 -1400 626
rect -1288 582 -1232 626
rect -1120 582 -1064 626
rect -952 582 -896 626
rect -784 582 -728 626
rect -616 582 -560 626
rect -448 582 -392 626
rect -280 582 -224 626
rect -112 582 -56 626
rect 56 582 112 626
rect 224 582 280 626
rect 392 582 448 626
rect 560 582 616 626
rect 728 582 784 626
rect 896 582 952 626
rect 1064 582 1120 626
rect 1232 582 1288 626
rect 1400 582 1456 626
rect 1568 582 1624 626
rect 1736 582 1792 626
rect 1904 582 1960 626
rect 2072 582 2128 626
rect 2240 582 2296 626
rect 2408 582 2464 626
rect 2576 582 2632 626
rect 2744 582 2800 626
rect 2912 582 2968 626
rect 3080 582 3136 626
rect 3248 582 3304 626
rect -3304 490 -3248 534
rect -3136 490 -3080 534
rect -2968 490 -2912 534
rect -2800 490 -2744 534
rect -2632 490 -2576 534
rect -2464 490 -2408 534
rect -2296 490 -2240 534
rect -2128 490 -2072 534
rect -1960 490 -1904 534
rect -1792 490 -1736 534
rect -1624 490 -1568 534
rect -1456 490 -1400 534
rect -1288 490 -1232 534
rect -1120 490 -1064 534
rect -952 490 -896 534
rect -784 490 -728 534
rect -616 490 -560 534
rect -448 490 -392 534
rect -280 490 -224 534
rect -112 490 -56 534
rect 56 490 112 534
rect 224 490 280 534
rect 392 490 448 534
rect 560 490 616 534
rect 728 490 784 534
rect 896 490 952 534
rect 1064 490 1120 534
rect 1232 490 1288 534
rect 1400 490 1456 534
rect 1568 490 1624 534
rect 1736 490 1792 534
rect 1904 490 1960 534
rect 2072 490 2128 534
rect 2240 490 2296 534
rect 2408 490 2464 534
rect 2576 490 2632 534
rect 2744 490 2800 534
rect 2912 490 2968 534
rect 3080 490 3136 534
rect 3248 490 3304 534
rect -3304 396 -3248 440
rect -3136 396 -3080 440
rect -2968 396 -2912 440
rect -2800 396 -2744 440
rect -2632 396 -2576 440
rect -2464 396 -2408 440
rect -2296 396 -2240 440
rect -2128 396 -2072 440
rect -1960 396 -1904 440
rect -1792 396 -1736 440
rect -1624 396 -1568 440
rect -1456 396 -1400 440
rect -1288 396 -1232 440
rect -1120 396 -1064 440
rect -952 396 -896 440
rect -784 396 -728 440
rect -616 396 -560 440
rect -448 396 -392 440
rect -280 396 -224 440
rect -112 396 -56 440
rect 56 396 112 440
rect 224 396 280 440
rect 392 396 448 440
rect 560 396 616 440
rect 728 396 784 440
rect 896 396 952 440
rect 1064 396 1120 440
rect 1232 396 1288 440
rect 1400 396 1456 440
rect 1568 396 1624 440
rect 1736 396 1792 440
rect 1904 396 1960 440
rect 2072 396 2128 440
rect 2240 396 2296 440
rect 2408 396 2464 440
rect 2576 396 2632 440
rect 2744 396 2800 440
rect 2912 396 2968 440
rect 3080 396 3136 440
rect 3248 396 3304 440
rect -3304 304 -3248 348
rect -3136 304 -3080 348
rect -2968 304 -2912 348
rect -2800 304 -2744 348
rect -2632 304 -2576 348
rect -2464 304 -2408 348
rect -2296 304 -2240 348
rect -2128 304 -2072 348
rect -1960 304 -1904 348
rect -1792 304 -1736 348
rect -1624 304 -1568 348
rect -1456 304 -1400 348
rect -1288 304 -1232 348
rect -1120 304 -1064 348
rect -952 304 -896 348
rect -784 304 -728 348
rect -616 304 -560 348
rect -448 304 -392 348
rect -280 304 -224 348
rect -112 304 -56 348
rect 56 304 112 348
rect 224 304 280 348
rect 392 304 448 348
rect 560 304 616 348
rect 728 304 784 348
rect 896 304 952 348
rect 1064 304 1120 348
rect 1232 304 1288 348
rect 1400 304 1456 348
rect 1568 304 1624 348
rect 1736 304 1792 348
rect 1904 304 1960 348
rect 2072 304 2128 348
rect 2240 304 2296 348
rect 2408 304 2464 348
rect 2576 304 2632 348
rect 2744 304 2800 348
rect 2912 304 2968 348
rect 3080 304 3136 348
rect 3248 304 3304 348
rect -3304 210 -3248 254
rect -3136 210 -3080 254
rect -2968 210 -2912 254
rect -2800 210 -2744 254
rect -2632 210 -2576 254
rect -2464 210 -2408 254
rect -2296 210 -2240 254
rect -2128 210 -2072 254
rect -1960 210 -1904 254
rect -1792 210 -1736 254
rect -1624 210 -1568 254
rect -1456 210 -1400 254
rect -1288 210 -1232 254
rect -1120 210 -1064 254
rect -952 210 -896 254
rect -784 210 -728 254
rect -616 210 -560 254
rect -448 210 -392 254
rect -280 210 -224 254
rect -112 210 -56 254
rect 56 210 112 254
rect 224 210 280 254
rect 392 210 448 254
rect 560 210 616 254
rect 728 210 784 254
rect 896 210 952 254
rect 1064 210 1120 254
rect 1232 210 1288 254
rect 1400 210 1456 254
rect 1568 210 1624 254
rect 1736 210 1792 254
rect 1904 210 1960 254
rect 2072 210 2128 254
rect 2240 210 2296 254
rect 2408 210 2464 254
rect 2576 210 2632 254
rect 2744 210 2800 254
rect 2912 210 2968 254
rect 3080 210 3136 254
rect 3248 210 3304 254
rect -3304 118 -3248 162
rect -3136 118 -3080 162
rect -2968 118 -2912 162
rect -2800 118 -2744 162
rect -2632 118 -2576 162
rect -2464 118 -2408 162
rect -2296 118 -2240 162
rect -2128 118 -2072 162
rect -1960 118 -1904 162
rect -1792 118 -1736 162
rect -1624 118 -1568 162
rect -1456 118 -1400 162
rect -1288 118 -1232 162
rect -1120 118 -1064 162
rect -952 118 -896 162
rect -784 118 -728 162
rect -616 118 -560 162
rect -448 118 -392 162
rect -280 118 -224 162
rect -112 118 -56 162
rect 56 118 112 162
rect 224 118 280 162
rect 392 118 448 162
rect 560 118 616 162
rect 728 118 784 162
rect 896 118 952 162
rect 1064 118 1120 162
rect 1232 118 1288 162
rect 1400 118 1456 162
rect 1568 118 1624 162
rect 1736 118 1792 162
rect 1904 118 1960 162
rect 2072 118 2128 162
rect 2240 118 2296 162
rect 2408 118 2464 162
rect 2576 118 2632 162
rect 2744 118 2800 162
rect 2912 118 2968 162
rect 3080 118 3136 162
rect 3248 118 3304 162
rect -3304 24 -3248 68
rect -3136 24 -3080 68
rect -2968 24 -2912 68
rect -2800 24 -2744 68
rect -2632 24 -2576 68
rect -2464 24 -2408 68
rect -2296 24 -2240 68
rect -2128 24 -2072 68
rect -1960 24 -1904 68
rect -1792 24 -1736 68
rect -1624 24 -1568 68
rect -1456 24 -1400 68
rect -1288 24 -1232 68
rect -1120 24 -1064 68
rect -952 24 -896 68
rect -784 24 -728 68
rect -616 24 -560 68
rect -448 24 -392 68
rect -280 24 -224 68
rect -112 24 -56 68
rect 56 24 112 68
rect 224 24 280 68
rect 392 24 448 68
rect 560 24 616 68
rect 728 24 784 68
rect 896 24 952 68
rect 1064 24 1120 68
rect 1232 24 1288 68
rect 1400 24 1456 68
rect 1568 24 1624 68
rect 1736 24 1792 68
rect 1904 24 1960 68
rect 2072 24 2128 68
rect 2240 24 2296 68
rect 2408 24 2464 68
rect 2576 24 2632 68
rect 2744 24 2800 68
rect 2912 24 2968 68
rect 3080 24 3136 68
rect 3248 24 3304 68
rect -3304 -68 -3248 -24
rect -3136 -68 -3080 -24
rect -2968 -68 -2912 -24
rect -2800 -68 -2744 -24
rect -2632 -68 -2576 -24
rect -2464 -68 -2408 -24
rect -2296 -68 -2240 -24
rect -2128 -68 -2072 -24
rect -1960 -68 -1904 -24
rect -1792 -68 -1736 -24
rect -1624 -68 -1568 -24
rect -1456 -68 -1400 -24
rect -1288 -68 -1232 -24
rect -1120 -68 -1064 -24
rect -952 -68 -896 -24
rect -784 -68 -728 -24
rect -616 -68 -560 -24
rect -448 -68 -392 -24
rect -280 -68 -224 -24
rect -112 -68 -56 -24
rect 56 -68 112 -24
rect 224 -68 280 -24
rect 392 -68 448 -24
rect 560 -68 616 -24
rect 728 -68 784 -24
rect 896 -68 952 -24
rect 1064 -68 1120 -24
rect 1232 -68 1288 -24
rect 1400 -68 1456 -24
rect 1568 -68 1624 -24
rect 1736 -68 1792 -24
rect 1904 -68 1960 -24
rect 2072 -68 2128 -24
rect 2240 -68 2296 -24
rect 2408 -68 2464 -24
rect 2576 -68 2632 -24
rect 2744 -68 2800 -24
rect 2912 -68 2968 -24
rect 3080 -68 3136 -24
rect 3248 -68 3304 -24
rect -3304 -162 -3248 -118
rect -3136 -162 -3080 -118
rect -2968 -162 -2912 -118
rect -2800 -162 -2744 -118
rect -2632 -162 -2576 -118
rect -2464 -162 -2408 -118
rect -2296 -162 -2240 -118
rect -2128 -162 -2072 -118
rect -1960 -162 -1904 -118
rect -1792 -162 -1736 -118
rect -1624 -162 -1568 -118
rect -1456 -162 -1400 -118
rect -1288 -162 -1232 -118
rect -1120 -162 -1064 -118
rect -952 -162 -896 -118
rect -784 -162 -728 -118
rect -616 -162 -560 -118
rect -448 -162 -392 -118
rect -280 -162 -224 -118
rect -112 -162 -56 -118
rect 56 -162 112 -118
rect 224 -162 280 -118
rect 392 -162 448 -118
rect 560 -162 616 -118
rect 728 -162 784 -118
rect 896 -162 952 -118
rect 1064 -162 1120 -118
rect 1232 -162 1288 -118
rect 1400 -162 1456 -118
rect 1568 -162 1624 -118
rect 1736 -162 1792 -118
rect 1904 -162 1960 -118
rect 2072 -162 2128 -118
rect 2240 -162 2296 -118
rect 2408 -162 2464 -118
rect 2576 -162 2632 -118
rect 2744 -162 2800 -118
rect 2912 -162 2968 -118
rect 3080 -162 3136 -118
rect 3248 -162 3304 -118
rect -3304 -254 -3248 -210
rect -3136 -254 -3080 -210
rect -2968 -254 -2912 -210
rect -2800 -254 -2744 -210
rect -2632 -254 -2576 -210
rect -2464 -254 -2408 -210
rect -2296 -254 -2240 -210
rect -2128 -254 -2072 -210
rect -1960 -254 -1904 -210
rect -1792 -254 -1736 -210
rect -1624 -254 -1568 -210
rect -1456 -254 -1400 -210
rect -1288 -254 -1232 -210
rect -1120 -254 -1064 -210
rect -952 -254 -896 -210
rect -784 -254 -728 -210
rect -616 -254 -560 -210
rect -448 -254 -392 -210
rect -280 -254 -224 -210
rect -112 -254 -56 -210
rect 56 -254 112 -210
rect 224 -254 280 -210
rect 392 -254 448 -210
rect 560 -254 616 -210
rect 728 -254 784 -210
rect 896 -254 952 -210
rect 1064 -254 1120 -210
rect 1232 -254 1288 -210
rect 1400 -254 1456 -210
rect 1568 -254 1624 -210
rect 1736 -254 1792 -210
rect 1904 -254 1960 -210
rect 2072 -254 2128 -210
rect 2240 -254 2296 -210
rect 2408 -254 2464 -210
rect 2576 -254 2632 -210
rect 2744 -254 2800 -210
rect 2912 -254 2968 -210
rect 3080 -254 3136 -210
rect 3248 -254 3304 -210
rect -3304 -348 -3248 -304
rect -3136 -348 -3080 -304
rect -2968 -348 -2912 -304
rect -2800 -348 -2744 -304
rect -2632 -348 -2576 -304
rect -2464 -348 -2408 -304
rect -2296 -348 -2240 -304
rect -2128 -348 -2072 -304
rect -1960 -348 -1904 -304
rect -1792 -348 -1736 -304
rect -1624 -348 -1568 -304
rect -1456 -348 -1400 -304
rect -1288 -348 -1232 -304
rect -1120 -348 -1064 -304
rect -952 -348 -896 -304
rect -784 -348 -728 -304
rect -616 -348 -560 -304
rect -448 -348 -392 -304
rect -280 -348 -224 -304
rect -112 -348 -56 -304
rect 56 -348 112 -304
rect 224 -348 280 -304
rect 392 -348 448 -304
rect 560 -348 616 -304
rect 728 -348 784 -304
rect 896 -348 952 -304
rect 1064 -348 1120 -304
rect 1232 -348 1288 -304
rect 1400 -348 1456 -304
rect 1568 -348 1624 -304
rect 1736 -348 1792 -304
rect 1904 -348 1960 -304
rect 2072 -348 2128 -304
rect 2240 -348 2296 -304
rect 2408 -348 2464 -304
rect 2576 -348 2632 -304
rect 2744 -348 2800 -304
rect 2912 -348 2968 -304
rect 3080 -348 3136 -304
rect 3248 -348 3304 -304
rect -3304 -440 -3248 -396
rect -3136 -440 -3080 -396
rect -2968 -440 -2912 -396
rect -2800 -440 -2744 -396
rect -2632 -440 -2576 -396
rect -2464 -440 -2408 -396
rect -2296 -440 -2240 -396
rect -2128 -440 -2072 -396
rect -1960 -440 -1904 -396
rect -1792 -440 -1736 -396
rect -1624 -440 -1568 -396
rect -1456 -440 -1400 -396
rect -1288 -440 -1232 -396
rect -1120 -440 -1064 -396
rect -952 -440 -896 -396
rect -784 -440 -728 -396
rect -616 -440 -560 -396
rect -448 -440 -392 -396
rect -280 -440 -224 -396
rect -112 -440 -56 -396
rect 56 -440 112 -396
rect 224 -440 280 -396
rect 392 -440 448 -396
rect 560 -440 616 -396
rect 728 -440 784 -396
rect 896 -440 952 -396
rect 1064 -440 1120 -396
rect 1232 -440 1288 -396
rect 1400 -440 1456 -396
rect 1568 -440 1624 -396
rect 1736 -440 1792 -396
rect 1904 -440 1960 -396
rect 2072 -440 2128 -396
rect 2240 -440 2296 -396
rect 2408 -440 2464 -396
rect 2576 -440 2632 -396
rect 2744 -440 2800 -396
rect 2912 -440 2968 -396
rect 3080 -440 3136 -396
rect 3248 -440 3304 -396
rect -3304 -534 -3248 -490
rect -3136 -534 -3080 -490
rect -2968 -534 -2912 -490
rect -2800 -534 -2744 -490
rect -2632 -534 -2576 -490
rect -2464 -534 -2408 -490
rect -2296 -534 -2240 -490
rect -2128 -534 -2072 -490
rect -1960 -534 -1904 -490
rect -1792 -534 -1736 -490
rect -1624 -534 -1568 -490
rect -1456 -534 -1400 -490
rect -1288 -534 -1232 -490
rect -1120 -534 -1064 -490
rect -952 -534 -896 -490
rect -784 -534 -728 -490
rect -616 -534 -560 -490
rect -448 -534 -392 -490
rect -280 -534 -224 -490
rect -112 -534 -56 -490
rect 56 -534 112 -490
rect 224 -534 280 -490
rect 392 -534 448 -490
rect 560 -534 616 -490
rect 728 -534 784 -490
rect 896 -534 952 -490
rect 1064 -534 1120 -490
rect 1232 -534 1288 -490
rect 1400 -534 1456 -490
rect 1568 -534 1624 -490
rect 1736 -534 1792 -490
rect 1904 -534 1960 -490
rect 2072 -534 2128 -490
rect 2240 -534 2296 -490
rect 2408 -534 2464 -490
rect 2576 -534 2632 -490
rect 2744 -534 2800 -490
rect 2912 -534 2968 -490
rect 3080 -534 3136 -490
rect 3248 -534 3304 -490
rect -3304 -626 -3248 -582
rect -3136 -626 -3080 -582
rect -2968 -626 -2912 -582
rect -2800 -626 -2744 -582
rect -2632 -626 -2576 -582
rect -2464 -626 -2408 -582
rect -2296 -626 -2240 -582
rect -2128 -626 -2072 -582
rect -1960 -626 -1904 -582
rect -1792 -626 -1736 -582
rect -1624 -626 -1568 -582
rect -1456 -626 -1400 -582
rect -1288 -626 -1232 -582
rect -1120 -626 -1064 -582
rect -952 -626 -896 -582
rect -784 -626 -728 -582
rect -616 -626 -560 -582
rect -448 -626 -392 -582
rect -280 -626 -224 -582
rect -112 -626 -56 -582
rect 56 -626 112 -582
rect 224 -626 280 -582
rect 392 -626 448 -582
rect 560 -626 616 -582
rect 728 -626 784 -582
rect 896 -626 952 -582
rect 1064 -626 1120 -582
rect 1232 -626 1288 -582
rect 1400 -626 1456 -582
rect 1568 -626 1624 -582
rect 1736 -626 1792 -582
rect 1904 -626 1960 -582
rect 2072 -626 2128 -582
rect 2240 -626 2296 -582
rect 2408 -626 2464 -582
rect 2576 -626 2632 -582
rect 2744 -626 2800 -582
rect 2912 -626 2968 -582
rect 3080 -626 3136 -582
rect 3248 -626 3304 -582
rect -3304 -720 -3248 -676
rect -3136 -720 -3080 -676
rect -2968 -720 -2912 -676
rect -2800 -720 -2744 -676
rect -2632 -720 -2576 -676
rect -2464 -720 -2408 -676
rect -2296 -720 -2240 -676
rect -2128 -720 -2072 -676
rect -1960 -720 -1904 -676
rect -1792 -720 -1736 -676
rect -1624 -720 -1568 -676
rect -1456 -720 -1400 -676
rect -1288 -720 -1232 -676
rect -1120 -720 -1064 -676
rect -952 -720 -896 -676
rect -784 -720 -728 -676
rect -616 -720 -560 -676
rect -448 -720 -392 -676
rect -280 -720 -224 -676
rect -112 -720 -56 -676
rect 56 -720 112 -676
rect 224 -720 280 -676
rect 392 -720 448 -676
rect 560 -720 616 -676
rect 728 -720 784 -676
rect 896 -720 952 -676
rect 1064 -720 1120 -676
rect 1232 -720 1288 -676
rect 1400 -720 1456 -676
rect 1568 -720 1624 -676
rect 1736 -720 1792 -676
rect 1904 -720 1960 -676
rect 2072 -720 2128 -676
rect 2240 -720 2296 -676
rect 2408 -720 2464 -676
rect 2576 -720 2632 -676
rect 2744 -720 2800 -676
rect 2912 -720 2968 -676
rect 3080 -720 3136 -676
rect 3248 -720 3304 -676
<< metal1 >>
rect -3394 628 -3383 674
rect -3337 628 -3326 674
rect -3226 628 -3215 674
rect -3169 628 -3158 674
rect -3058 628 -3047 674
rect -3001 628 -2990 674
rect -2890 628 -2879 674
rect -2833 628 -2822 674
rect -2722 628 -2711 674
rect -2665 628 -2654 674
rect -2554 628 -2543 674
rect -2497 628 -2486 674
rect -2386 628 -2375 674
rect -2329 628 -2318 674
rect -2218 628 -2207 674
rect -2161 628 -2150 674
rect -2050 628 -2039 674
rect -1993 628 -1982 674
rect -1882 628 -1871 674
rect -1825 628 -1814 674
rect -1714 628 -1703 674
rect -1657 628 -1646 674
rect -1546 628 -1535 674
rect -1489 628 -1478 674
rect -1378 628 -1367 674
rect -1321 628 -1310 674
rect -1210 628 -1199 674
rect -1153 628 -1142 674
rect -1042 628 -1031 674
rect -985 628 -974 674
rect -874 628 -863 674
rect -817 628 -806 674
rect -706 628 -695 674
rect -649 628 -638 674
rect -538 628 -527 674
rect -481 628 -470 674
rect -370 628 -359 674
rect -313 628 -302 674
rect -202 628 -191 674
rect -145 628 -134 674
rect -34 628 -23 674
rect 23 628 34 674
rect 134 628 145 674
rect 191 628 202 674
rect 302 628 313 674
rect 359 628 370 674
rect 470 628 481 674
rect 527 628 538 674
rect 638 628 649 674
rect 695 628 706 674
rect 806 628 817 674
rect 863 628 874 674
rect 974 628 985 674
rect 1031 628 1042 674
rect 1142 628 1153 674
rect 1199 628 1210 674
rect 1310 628 1321 674
rect 1367 628 1378 674
rect 1478 628 1489 674
rect 1535 628 1546 674
rect 1646 628 1657 674
rect 1703 628 1714 674
rect 1814 628 1825 674
rect 1871 628 1882 674
rect 1982 628 1993 674
rect 2039 628 2050 674
rect 2150 628 2161 674
rect 2207 628 2218 674
rect 2318 628 2329 674
rect 2375 628 2386 674
rect 2486 628 2497 674
rect 2543 628 2554 674
rect 2654 628 2665 674
rect 2711 628 2722 674
rect 2822 628 2833 674
rect 2879 628 2890 674
rect 2990 628 3001 674
rect 3047 628 3058 674
rect 3158 628 3169 674
rect 3215 628 3226 674
rect 3326 628 3337 674
rect 3383 628 3394 674
rect -3394 442 -3383 488
rect -3337 442 -3326 488
rect -3226 442 -3215 488
rect -3169 442 -3158 488
rect -3058 442 -3047 488
rect -3001 442 -2990 488
rect -2890 442 -2879 488
rect -2833 442 -2822 488
rect -2722 442 -2711 488
rect -2665 442 -2654 488
rect -2554 442 -2543 488
rect -2497 442 -2486 488
rect -2386 442 -2375 488
rect -2329 442 -2318 488
rect -2218 442 -2207 488
rect -2161 442 -2150 488
rect -2050 442 -2039 488
rect -1993 442 -1982 488
rect -1882 442 -1871 488
rect -1825 442 -1814 488
rect -1714 442 -1703 488
rect -1657 442 -1646 488
rect -1546 442 -1535 488
rect -1489 442 -1478 488
rect -1378 442 -1367 488
rect -1321 442 -1310 488
rect -1210 442 -1199 488
rect -1153 442 -1142 488
rect -1042 442 -1031 488
rect -985 442 -974 488
rect -874 442 -863 488
rect -817 442 -806 488
rect -706 442 -695 488
rect -649 442 -638 488
rect -538 442 -527 488
rect -481 442 -470 488
rect -370 442 -359 488
rect -313 442 -302 488
rect -202 442 -191 488
rect -145 442 -134 488
rect -34 442 -23 488
rect 23 442 34 488
rect 134 442 145 488
rect 191 442 202 488
rect 302 442 313 488
rect 359 442 370 488
rect 470 442 481 488
rect 527 442 538 488
rect 638 442 649 488
rect 695 442 706 488
rect 806 442 817 488
rect 863 442 874 488
rect 974 442 985 488
rect 1031 442 1042 488
rect 1142 442 1153 488
rect 1199 442 1210 488
rect 1310 442 1321 488
rect 1367 442 1378 488
rect 1478 442 1489 488
rect 1535 442 1546 488
rect 1646 442 1657 488
rect 1703 442 1714 488
rect 1814 442 1825 488
rect 1871 442 1882 488
rect 1982 442 1993 488
rect 2039 442 2050 488
rect 2150 442 2161 488
rect 2207 442 2218 488
rect 2318 442 2329 488
rect 2375 442 2386 488
rect 2486 442 2497 488
rect 2543 442 2554 488
rect 2654 442 2665 488
rect 2711 442 2722 488
rect 2822 442 2833 488
rect 2879 442 2890 488
rect 2990 442 3001 488
rect 3047 442 3058 488
rect 3158 442 3169 488
rect 3215 442 3226 488
rect 3326 442 3337 488
rect 3383 442 3394 488
rect -3394 256 -3383 302
rect -3337 256 -3326 302
rect -3226 256 -3215 302
rect -3169 256 -3158 302
rect -3058 256 -3047 302
rect -3001 256 -2990 302
rect -2890 256 -2879 302
rect -2833 256 -2822 302
rect -2722 256 -2711 302
rect -2665 256 -2654 302
rect -2554 256 -2543 302
rect -2497 256 -2486 302
rect -2386 256 -2375 302
rect -2329 256 -2318 302
rect -2218 256 -2207 302
rect -2161 256 -2150 302
rect -2050 256 -2039 302
rect -1993 256 -1982 302
rect -1882 256 -1871 302
rect -1825 256 -1814 302
rect -1714 256 -1703 302
rect -1657 256 -1646 302
rect -1546 256 -1535 302
rect -1489 256 -1478 302
rect -1378 256 -1367 302
rect -1321 256 -1310 302
rect -1210 256 -1199 302
rect -1153 256 -1142 302
rect -1042 256 -1031 302
rect -985 256 -974 302
rect -874 256 -863 302
rect -817 256 -806 302
rect -706 256 -695 302
rect -649 256 -638 302
rect -538 256 -527 302
rect -481 256 -470 302
rect -370 256 -359 302
rect -313 256 -302 302
rect -202 256 -191 302
rect -145 256 -134 302
rect -34 256 -23 302
rect 23 256 34 302
rect 134 256 145 302
rect 191 256 202 302
rect 302 256 313 302
rect 359 256 370 302
rect 470 256 481 302
rect 527 256 538 302
rect 638 256 649 302
rect 695 256 706 302
rect 806 256 817 302
rect 863 256 874 302
rect 974 256 985 302
rect 1031 256 1042 302
rect 1142 256 1153 302
rect 1199 256 1210 302
rect 1310 256 1321 302
rect 1367 256 1378 302
rect 1478 256 1489 302
rect 1535 256 1546 302
rect 1646 256 1657 302
rect 1703 256 1714 302
rect 1814 256 1825 302
rect 1871 256 1882 302
rect 1982 256 1993 302
rect 2039 256 2050 302
rect 2150 256 2161 302
rect 2207 256 2218 302
rect 2318 256 2329 302
rect 2375 256 2386 302
rect 2486 256 2497 302
rect 2543 256 2554 302
rect 2654 256 2665 302
rect 2711 256 2722 302
rect 2822 256 2833 302
rect 2879 256 2890 302
rect 2990 256 3001 302
rect 3047 256 3058 302
rect 3158 256 3169 302
rect 3215 256 3226 302
rect 3326 256 3337 302
rect 3383 256 3394 302
rect -3394 70 -3383 116
rect -3337 70 -3326 116
rect -3226 70 -3215 116
rect -3169 70 -3158 116
rect -3058 70 -3047 116
rect -3001 70 -2990 116
rect -2890 70 -2879 116
rect -2833 70 -2822 116
rect -2722 70 -2711 116
rect -2665 70 -2654 116
rect -2554 70 -2543 116
rect -2497 70 -2486 116
rect -2386 70 -2375 116
rect -2329 70 -2318 116
rect -2218 70 -2207 116
rect -2161 70 -2150 116
rect -2050 70 -2039 116
rect -1993 70 -1982 116
rect -1882 70 -1871 116
rect -1825 70 -1814 116
rect -1714 70 -1703 116
rect -1657 70 -1646 116
rect -1546 70 -1535 116
rect -1489 70 -1478 116
rect -1378 70 -1367 116
rect -1321 70 -1310 116
rect -1210 70 -1199 116
rect -1153 70 -1142 116
rect -1042 70 -1031 116
rect -985 70 -974 116
rect -874 70 -863 116
rect -817 70 -806 116
rect -706 70 -695 116
rect -649 70 -638 116
rect -538 70 -527 116
rect -481 70 -470 116
rect -370 70 -359 116
rect -313 70 -302 116
rect -202 70 -191 116
rect -145 70 -134 116
rect -34 70 -23 116
rect 23 70 34 116
rect 134 70 145 116
rect 191 70 202 116
rect 302 70 313 116
rect 359 70 370 116
rect 470 70 481 116
rect 527 70 538 116
rect 638 70 649 116
rect 695 70 706 116
rect 806 70 817 116
rect 863 70 874 116
rect 974 70 985 116
rect 1031 70 1042 116
rect 1142 70 1153 116
rect 1199 70 1210 116
rect 1310 70 1321 116
rect 1367 70 1378 116
rect 1478 70 1489 116
rect 1535 70 1546 116
rect 1646 70 1657 116
rect 1703 70 1714 116
rect 1814 70 1825 116
rect 1871 70 1882 116
rect 1982 70 1993 116
rect 2039 70 2050 116
rect 2150 70 2161 116
rect 2207 70 2218 116
rect 2318 70 2329 116
rect 2375 70 2386 116
rect 2486 70 2497 116
rect 2543 70 2554 116
rect 2654 70 2665 116
rect 2711 70 2722 116
rect 2822 70 2833 116
rect 2879 70 2890 116
rect 2990 70 3001 116
rect 3047 70 3058 116
rect 3158 70 3169 116
rect 3215 70 3226 116
rect 3326 70 3337 116
rect 3383 70 3394 116
rect -3394 -116 -3383 -70
rect -3337 -116 -3326 -70
rect -3226 -116 -3215 -70
rect -3169 -116 -3158 -70
rect -3058 -116 -3047 -70
rect -3001 -116 -2990 -70
rect -2890 -116 -2879 -70
rect -2833 -116 -2822 -70
rect -2722 -116 -2711 -70
rect -2665 -116 -2654 -70
rect -2554 -116 -2543 -70
rect -2497 -116 -2486 -70
rect -2386 -116 -2375 -70
rect -2329 -116 -2318 -70
rect -2218 -116 -2207 -70
rect -2161 -116 -2150 -70
rect -2050 -116 -2039 -70
rect -1993 -116 -1982 -70
rect -1882 -116 -1871 -70
rect -1825 -116 -1814 -70
rect -1714 -116 -1703 -70
rect -1657 -116 -1646 -70
rect -1546 -116 -1535 -70
rect -1489 -116 -1478 -70
rect -1378 -116 -1367 -70
rect -1321 -116 -1310 -70
rect -1210 -116 -1199 -70
rect -1153 -116 -1142 -70
rect -1042 -116 -1031 -70
rect -985 -116 -974 -70
rect -874 -116 -863 -70
rect -817 -116 -806 -70
rect -706 -116 -695 -70
rect -649 -116 -638 -70
rect -538 -116 -527 -70
rect -481 -116 -470 -70
rect -370 -116 -359 -70
rect -313 -116 -302 -70
rect -202 -116 -191 -70
rect -145 -116 -134 -70
rect -34 -116 -23 -70
rect 23 -116 34 -70
rect 134 -116 145 -70
rect 191 -116 202 -70
rect 302 -116 313 -70
rect 359 -116 370 -70
rect 470 -116 481 -70
rect 527 -116 538 -70
rect 638 -116 649 -70
rect 695 -116 706 -70
rect 806 -116 817 -70
rect 863 -116 874 -70
rect 974 -116 985 -70
rect 1031 -116 1042 -70
rect 1142 -116 1153 -70
rect 1199 -116 1210 -70
rect 1310 -116 1321 -70
rect 1367 -116 1378 -70
rect 1478 -116 1489 -70
rect 1535 -116 1546 -70
rect 1646 -116 1657 -70
rect 1703 -116 1714 -70
rect 1814 -116 1825 -70
rect 1871 -116 1882 -70
rect 1982 -116 1993 -70
rect 2039 -116 2050 -70
rect 2150 -116 2161 -70
rect 2207 -116 2218 -70
rect 2318 -116 2329 -70
rect 2375 -116 2386 -70
rect 2486 -116 2497 -70
rect 2543 -116 2554 -70
rect 2654 -116 2665 -70
rect 2711 -116 2722 -70
rect 2822 -116 2833 -70
rect 2879 -116 2890 -70
rect 2990 -116 3001 -70
rect 3047 -116 3058 -70
rect 3158 -116 3169 -70
rect 3215 -116 3226 -70
rect 3326 -116 3337 -70
rect 3383 -116 3394 -70
rect -3394 -302 -3383 -256
rect -3337 -302 -3326 -256
rect -3226 -302 -3215 -256
rect -3169 -302 -3158 -256
rect -3058 -302 -3047 -256
rect -3001 -302 -2990 -256
rect -2890 -302 -2879 -256
rect -2833 -302 -2822 -256
rect -2722 -302 -2711 -256
rect -2665 -302 -2654 -256
rect -2554 -302 -2543 -256
rect -2497 -302 -2486 -256
rect -2386 -302 -2375 -256
rect -2329 -302 -2318 -256
rect -2218 -302 -2207 -256
rect -2161 -302 -2150 -256
rect -2050 -302 -2039 -256
rect -1993 -302 -1982 -256
rect -1882 -302 -1871 -256
rect -1825 -302 -1814 -256
rect -1714 -302 -1703 -256
rect -1657 -302 -1646 -256
rect -1546 -302 -1535 -256
rect -1489 -302 -1478 -256
rect -1378 -302 -1367 -256
rect -1321 -302 -1310 -256
rect -1210 -302 -1199 -256
rect -1153 -302 -1142 -256
rect -1042 -302 -1031 -256
rect -985 -302 -974 -256
rect -874 -302 -863 -256
rect -817 -302 -806 -256
rect -706 -302 -695 -256
rect -649 -302 -638 -256
rect -538 -302 -527 -256
rect -481 -302 -470 -256
rect -370 -302 -359 -256
rect -313 -302 -302 -256
rect -202 -302 -191 -256
rect -145 -302 -134 -256
rect -34 -302 -23 -256
rect 23 -302 34 -256
rect 134 -302 145 -256
rect 191 -302 202 -256
rect 302 -302 313 -256
rect 359 -302 370 -256
rect 470 -302 481 -256
rect 527 -302 538 -256
rect 638 -302 649 -256
rect 695 -302 706 -256
rect 806 -302 817 -256
rect 863 -302 874 -256
rect 974 -302 985 -256
rect 1031 -302 1042 -256
rect 1142 -302 1153 -256
rect 1199 -302 1210 -256
rect 1310 -302 1321 -256
rect 1367 -302 1378 -256
rect 1478 -302 1489 -256
rect 1535 -302 1546 -256
rect 1646 -302 1657 -256
rect 1703 -302 1714 -256
rect 1814 -302 1825 -256
rect 1871 -302 1882 -256
rect 1982 -302 1993 -256
rect 2039 -302 2050 -256
rect 2150 -302 2161 -256
rect 2207 -302 2218 -256
rect 2318 -302 2329 -256
rect 2375 -302 2386 -256
rect 2486 -302 2497 -256
rect 2543 -302 2554 -256
rect 2654 -302 2665 -256
rect 2711 -302 2722 -256
rect 2822 -302 2833 -256
rect 2879 -302 2890 -256
rect 2990 -302 3001 -256
rect 3047 -302 3058 -256
rect 3158 -302 3169 -256
rect 3215 -302 3226 -256
rect 3326 -302 3337 -256
rect 3383 -302 3394 -256
rect -3394 -488 -3383 -442
rect -3337 -488 -3326 -442
rect -3226 -488 -3215 -442
rect -3169 -488 -3158 -442
rect -3058 -488 -3047 -442
rect -3001 -488 -2990 -442
rect -2890 -488 -2879 -442
rect -2833 -488 -2822 -442
rect -2722 -488 -2711 -442
rect -2665 -488 -2654 -442
rect -2554 -488 -2543 -442
rect -2497 -488 -2486 -442
rect -2386 -488 -2375 -442
rect -2329 -488 -2318 -442
rect -2218 -488 -2207 -442
rect -2161 -488 -2150 -442
rect -2050 -488 -2039 -442
rect -1993 -488 -1982 -442
rect -1882 -488 -1871 -442
rect -1825 -488 -1814 -442
rect -1714 -488 -1703 -442
rect -1657 -488 -1646 -442
rect -1546 -488 -1535 -442
rect -1489 -488 -1478 -442
rect -1378 -488 -1367 -442
rect -1321 -488 -1310 -442
rect -1210 -488 -1199 -442
rect -1153 -488 -1142 -442
rect -1042 -488 -1031 -442
rect -985 -488 -974 -442
rect -874 -488 -863 -442
rect -817 -488 -806 -442
rect -706 -488 -695 -442
rect -649 -488 -638 -442
rect -538 -488 -527 -442
rect -481 -488 -470 -442
rect -370 -488 -359 -442
rect -313 -488 -302 -442
rect -202 -488 -191 -442
rect -145 -488 -134 -442
rect -34 -488 -23 -442
rect 23 -488 34 -442
rect 134 -488 145 -442
rect 191 -488 202 -442
rect 302 -488 313 -442
rect 359 -488 370 -442
rect 470 -488 481 -442
rect 527 -488 538 -442
rect 638 -488 649 -442
rect 695 -488 706 -442
rect 806 -488 817 -442
rect 863 -488 874 -442
rect 974 -488 985 -442
rect 1031 -488 1042 -442
rect 1142 -488 1153 -442
rect 1199 -488 1210 -442
rect 1310 -488 1321 -442
rect 1367 -488 1378 -442
rect 1478 -488 1489 -442
rect 1535 -488 1546 -442
rect 1646 -488 1657 -442
rect 1703 -488 1714 -442
rect 1814 -488 1825 -442
rect 1871 -488 1882 -442
rect 1982 -488 1993 -442
rect 2039 -488 2050 -442
rect 2150 -488 2161 -442
rect 2207 -488 2218 -442
rect 2318 -488 2329 -442
rect 2375 -488 2386 -442
rect 2486 -488 2497 -442
rect 2543 -488 2554 -442
rect 2654 -488 2665 -442
rect 2711 -488 2722 -442
rect 2822 -488 2833 -442
rect 2879 -488 2890 -442
rect 2990 -488 3001 -442
rect 3047 -488 3058 -442
rect 3158 -488 3169 -442
rect 3215 -488 3226 -442
rect 3326 -488 3337 -442
rect 3383 -488 3394 -442
rect -3394 -674 -3383 -628
rect -3337 -674 -3326 -628
rect -3226 -674 -3215 -628
rect -3169 -674 -3158 -628
rect -3058 -674 -3047 -628
rect -3001 -674 -2990 -628
rect -2890 -674 -2879 -628
rect -2833 -674 -2822 -628
rect -2722 -674 -2711 -628
rect -2665 -674 -2654 -628
rect -2554 -674 -2543 -628
rect -2497 -674 -2486 -628
rect -2386 -674 -2375 -628
rect -2329 -674 -2318 -628
rect -2218 -674 -2207 -628
rect -2161 -674 -2150 -628
rect -2050 -674 -2039 -628
rect -1993 -674 -1982 -628
rect -1882 -674 -1871 -628
rect -1825 -674 -1814 -628
rect -1714 -674 -1703 -628
rect -1657 -674 -1646 -628
rect -1546 -674 -1535 -628
rect -1489 -674 -1478 -628
rect -1378 -674 -1367 -628
rect -1321 -674 -1310 -628
rect -1210 -674 -1199 -628
rect -1153 -674 -1142 -628
rect -1042 -674 -1031 -628
rect -985 -674 -974 -628
rect -874 -674 -863 -628
rect -817 -674 -806 -628
rect -706 -674 -695 -628
rect -649 -674 -638 -628
rect -538 -674 -527 -628
rect -481 -674 -470 -628
rect -370 -674 -359 -628
rect -313 -674 -302 -628
rect -202 -674 -191 -628
rect -145 -674 -134 -628
rect -34 -674 -23 -628
rect 23 -674 34 -628
rect 134 -674 145 -628
rect 191 -674 202 -628
rect 302 -674 313 -628
rect 359 -674 370 -628
rect 470 -674 481 -628
rect 527 -674 538 -628
rect 638 -674 649 -628
rect 695 -674 706 -628
rect 806 -674 817 -628
rect 863 -674 874 -628
rect 974 -674 985 -628
rect 1031 -674 1042 -628
rect 1142 -674 1153 -628
rect 1199 -674 1210 -628
rect 1310 -674 1321 -628
rect 1367 -674 1378 -628
rect 1478 -674 1489 -628
rect 1535 -674 1546 -628
rect 1646 -674 1657 -628
rect 1703 -674 1714 -628
rect 1814 -674 1825 -628
rect 1871 -674 1882 -628
rect 1982 -674 1993 -628
rect 2039 -674 2050 -628
rect 2150 -674 2161 -628
rect 2207 -674 2218 -628
rect 2318 -674 2329 -628
rect 2375 -674 2386 -628
rect 2486 -674 2497 -628
rect 2543 -674 2554 -628
rect 2654 -674 2665 -628
rect 2711 -674 2722 -628
rect 2822 -674 2833 -628
rect 2879 -674 2890 -628
rect 2990 -674 3001 -628
rect 3047 -674 3058 -628
rect 3158 -674 3169 -628
rect 3215 -674 3226 -628
rect 3326 -674 3337 -628
rect 3383 -674 3394 -628
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.250 l 0.280 m 8 nf 40 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
