magic
tech gf180mcuC
magscale 1 10
timestamp 1714558667
<< error_s >>
rect 9563 4519 9573 4556
rect 9619 4475 9629 4519
rect 10612 2382 10641 2402
<< nwell >>
rect 2785 2433 3073 2794
rect 5745 2433 5861 2435
rect -19 2081 5861 2433
rect 10597 2382 10612 2510
rect 10685 2474 10686 2492
rect 11607 2289 11692 2348
rect -19 1969 6016 2081
rect 2705 1604 2945 1969
rect 5745 1613 6016 1969
<< nsubdiff >>
rect 10597 2474 10686 2510
rect 10597 2473 10685 2474
rect 10474 2428 10739 2473
rect 10597 2382 10612 2428
<< polysilicon >>
rect 11607 2289 11692 2348
<< metal1 >>
rect 10647 4650 11322 4666
rect -163 4415 5621 4513
rect -454 4396 5621 4415
rect -459 4313 5621 4396
rect 5739 4475 5871 4532
rect 10647 4477 11200 4650
rect 11309 4477 11322 4650
rect 5739 4473 6758 4475
rect 5739 4392 5750 4473
rect 5855 4398 6758 4473
rect 10647 4435 11322 4477
rect 5855 4392 5871 4398
rect 5739 4380 5871 4392
rect 6681 4388 6758 4398
rect 6681 4325 6788 4388
rect 6701 4323 6788 4325
rect -459 4306 -55 4313
rect -459 1301 -295 4306
rect 2452 4304 2970 4313
rect 6032 4215 6118 4224
rect 6032 4148 6044 4215
rect 6106 4198 6118 4215
rect 6106 4148 6774 4198
rect 6032 4138 6774 4148
rect 5871 4085 5947 4097
rect 10658 4095 13910 4131
rect 5871 4012 5881 4085
rect 5935 4071 5947 4085
rect 6413 4077 6502 4090
rect 6413 4071 6420 4077
rect 5935 4024 6420 4071
rect 5935 4012 5947 4024
rect 5871 3999 5947 4012
rect 6413 4016 6420 4024
rect 6487 4071 6502 4077
rect 6487 4024 6787 4071
rect 6487 4016 6502 4024
rect 6413 3999 6502 4016
rect 10658 4019 13783 4095
rect 13893 4019 13910 4095
rect 10658 3993 13910 4019
rect 2275 3967 2363 3977
rect 2275 3901 2285 3967
rect 2351 3901 2363 3967
rect 2275 3892 2363 3901
rect 5326 3940 5426 3954
rect 5326 3881 5338 3940
rect 5415 3881 5426 3940
rect 6225 3953 6312 3955
rect 6225 3946 6808 3953
rect 6225 3892 6235 3946
rect 6294 3898 6808 3946
rect 6294 3892 6312 3898
rect 6225 3891 6312 3892
rect 6225 3882 6311 3891
rect 5326 3869 5426 3881
rect 1248 3864 1328 3867
rect 1248 3812 1258 3864
rect 1315 3812 1328 3864
rect 1248 3809 1328 3812
rect 4288 3864 4388 3866
rect 4288 3812 4322 3864
rect 4374 3812 4388 3864
rect 4288 3808 4388 3812
rect 5905 3836 5971 3846
rect 5905 3832 6804 3836
rect 5905 3778 5912 3832
rect 5964 3778 6804 3832
rect 5905 3772 6804 3778
rect 5905 3765 5971 3772
rect 5587 3352 6843 3541
rect 11845 3236 12035 3262
rect 6230 3174 6312 3186
rect 6230 3172 6793 3174
rect 6230 3118 6241 3172
rect 6300 3118 6793 3172
rect 6230 3112 6793 3118
rect 6230 3109 6312 3112
rect 11845 3069 11867 3236
rect 12009 3069 12035 3236
rect 11845 3040 12035 3069
rect 6409 2936 6496 2943
rect 2264 2895 2352 2907
rect 13 2839 71 2872
rect 2264 2841 2276 2895
rect 2345 2841 2352 2895
rect 5328 2875 5407 2883
rect 2264 2838 2352 2841
rect 3073 2840 3131 2873
rect 2270 2810 2351 2838
rect 5328 2822 5337 2875
rect 5395 2822 5407 2875
rect 6409 2881 6425 2936
rect 6484 2925 6496 2936
rect 6484 2881 6811 2925
rect 6409 2878 6811 2881
rect 11028 2902 11155 2923
rect 6409 2868 6496 2878
rect 11028 2840 11047 2902
rect 11135 2840 11155 2902
rect 5328 2809 5407 2822
rect 5725 2835 5847 2836
rect 5725 2829 5848 2835
rect 5725 2765 5766 2829
rect 5832 2765 5848 2829
rect 11028 2821 11155 2840
rect 11212 2918 11315 2928
rect 11212 2842 11221 2918
rect 11300 2877 11315 2918
rect 11300 2842 11361 2877
rect 5725 2760 5848 2765
rect 11212 2816 11361 2842
rect 5725 2756 5847 2760
rect 6030 2644 6130 2658
rect 6030 2565 6036 2644
rect 6118 2629 6130 2644
rect 6118 2565 6778 2629
rect 6030 2561 6778 2565
rect 6030 2552 6130 2561
rect 11212 2440 11315 2816
rect -170 2073 8973 2344
rect 10981 2337 11315 2440
rect 11607 2345 11692 2348
rect 11607 2292 11622 2345
rect 11679 2292 11692 2345
rect 11607 2289 11692 2292
rect 11411 2277 11513 2283
rect 11411 2224 11423 2277
rect 11501 2224 11513 2277
rect 12200 2244 12576 2302
rect 11411 2214 11513 2224
rect 11863 1843 12268 1941
rect 9085 1619 9426 1755
rect 3386 1592 3490 1601
rect 349 1582 440 1589
rect 349 1529 364 1582
rect 428 1529 440 1582
rect 349 1523 440 1529
rect 2620 1520 2677 1576
rect 3386 1528 3395 1592
rect 3477 1528 3490 1592
rect 6464 1591 6553 1600
rect 5663 1530 5720 1586
rect 3386 1518 3490 1528
rect 6464 1527 6478 1591
rect 6543 1527 6553 1591
rect 8735 1528 8792 1584
rect 6464 1517 6553 1527
rect -459 1137 292 1301
rect -454 1081 292 1137
rect 4403 598 4501 600
rect 1361 588 1460 590
rect 1361 536 1374 588
rect 1439 536 1460 588
rect 4403 544 4415 598
rect 4477 544 4501 598
rect 4403 541 4501 544
rect 1361 532 1460 536
rect 349 500 440 513
rect 349 441 360 500
rect 414 441 440 500
rect 3387 510 3459 520
rect 3387 458 3396 510
rect 3449 458 3459 510
rect 3387 450 3459 458
rect 6464 506 6542 514
rect 349 426 440 441
rect 6464 446 6475 506
rect 6532 446 6542 506
rect 6464 437 6542 446
rect 9085 101 9156 1619
rect 13774 1476 13910 1487
rect 13774 1460 13783 1476
rect 13635 1399 13783 1460
rect 13901 1399 13910 1476
rect 13635 1388 13910 1399
rect 9347 985 9477 997
rect 9347 904 9376 985
rect 9444 904 9477 985
rect 9347 896 9477 904
rect 13587 494 13710 496
rect 13587 488 13711 494
rect 13587 410 13597 488
rect 13700 410 13711 488
rect 13587 400 13711 410
rect 128 -156 13617 101
<< via1 >>
rect 11200 4477 11309 4650
rect 5750 4392 5855 4473
rect 6044 4148 6106 4215
rect 5881 4012 5935 4085
rect 6420 4016 6487 4077
rect 13783 4019 13893 4095
rect 2285 3901 2351 3967
rect 5338 3881 5415 3940
rect 6235 3892 6294 3946
rect 1258 3812 1315 3864
rect 4322 3812 4374 3864
rect 5912 3778 5964 3832
rect 2286 3391 2352 3457
rect 5354 3423 5412 3476
rect 6241 3118 6300 3172
rect 11867 3069 12009 3236
rect 2276 2841 2345 2895
rect 5337 2822 5395 2875
rect 6425 2881 6484 2936
rect 11047 2840 11135 2902
rect 5766 2765 5832 2829
rect 11221 2842 11300 2918
rect 6036 2565 6118 2644
rect 11622 2292 11679 2345
rect 11423 2224 11501 2277
rect 364 1529 428 1582
rect 3395 1528 3477 1592
rect 6478 1527 6543 1591
rect 356 909 410 968
rect 3390 930 3445 1001
rect 6471 915 6536 979
rect 8899 908 8967 989
rect 1374 536 1439 588
rect 4415 544 4477 598
rect 7487 542 7553 594
rect 360 441 414 500
rect 3396 458 3449 510
rect 6475 446 6532 506
rect 13783 1399 13901 1476
rect 9376 904 9444 985
rect 13597 410 13700 488
<< metal2 >>
rect 11178 4650 11321 4665
rect 5739 4477 5871 4532
rect 5739 4387 5747 4477
rect 5860 4387 5871 4477
rect 11178 4477 11200 4650
rect 11309 4477 11321 4650
rect 11178 4448 11321 4477
rect 5739 4380 5871 4387
rect 2653 4264 6118 4322
rect 6638 4304 6758 4398
rect 2653 4205 2711 4264
rect 1672 4147 2711 4205
rect 6032 4215 6118 4264
rect 6032 4148 6044 4215
rect 6106 4148 6118 4215
rect 5871 4085 5947 4097
rect 5871 4076 5881 4085
rect 4920 4012 5881 4076
rect 5935 4012 5947 4085
rect 4920 4011 5947 4012
rect 5871 3999 5947 4011
rect 2275 3967 2363 3977
rect 2275 3901 2285 3967
rect 2351 3901 2363 3967
rect 2275 3892 2363 3901
rect 5326 3940 5426 3954
rect 1248 3874 1338 3884
rect 1248 3804 1258 3874
rect 1329 3804 1338 3874
rect 1248 3793 1338 3804
rect 2278 3457 2358 3892
rect 5326 3881 5338 3940
rect 5415 3881 5426 3940
rect 4308 3874 4400 3877
rect 4308 3866 4319 3874
rect 4298 3808 4319 3866
rect 4308 3804 4319 3808
rect 4390 3804 4400 3874
rect 5326 3869 5426 3881
rect 4308 3798 4400 3804
rect 2278 3391 2286 3457
rect 2352 3391 2358 3457
rect 1 2885 57 3015
rect 2278 2907 2358 3391
rect 5350 3476 5422 3869
rect 5905 3832 5971 3846
rect 5905 3778 5912 3832
rect 5964 3778 5971 3832
rect 5905 3765 5971 3778
rect 5350 3423 5354 3476
rect 5412 3423 5422 3476
rect -80 2824 57 2885
rect 2264 2895 2358 2907
rect 2264 2841 2276 2895
rect 2345 2841 2358 2895
rect 3061 2885 3117 2977
rect 2264 2838 2358 2841
rect -80 1705 14 2824
rect 2270 2810 2358 2838
rect 2745 2829 3117 2885
rect 5350 2883 5422 3423
rect 2278 2809 2358 2810
rect 2600 2828 3117 2829
rect 5328 2875 5422 2883
rect 2278 2808 2352 2809
rect 2600 2757 3061 2828
rect 5328 2822 5337 2875
rect 5395 2822 5422 2875
rect 5725 2835 5847 2836
rect 5328 2809 5422 2822
rect 5350 2807 5422 2809
rect 5659 2832 5848 2835
rect 5659 2762 5732 2832
rect 5836 2762 5848 2832
rect 5659 2760 5848 2762
rect 5659 2757 5847 2760
rect 5659 2693 5716 2757
rect 5909 2285 5966 3765
rect 6032 2658 6118 4148
rect 6413 4077 6502 4090
rect 6413 4076 6420 4077
rect 6405 4016 6420 4076
rect 6487 4016 6502 4077
rect 6405 4011 6502 4016
rect 6413 3999 6502 4011
rect 6222 3946 6309 3965
rect 6222 3892 6235 3946
rect 6294 3892 6309 3946
rect 6222 3172 6309 3892
rect 6222 3118 6241 3172
rect 6300 3118 6309 3172
rect 6030 2644 6130 2658
rect 6030 2565 6036 2644
rect 6118 2565 6130 2644
rect 6030 2552 6130 2565
rect 2656 2206 5966 2285
rect 2657 2171 5966 2206
rect -80 1648 297 1705
rect -80 1570 93 1648
rect 349 1582 440 1589
rect 349 1529 364 1582
rect 428 1529 440 1582
rect 349 1523 440 1529
rect 2657 1584 2770 2171
rect 6222 2095 6309 3118
rect 6421 2943 6486 3999
rect 6559 3778 6764 3834
rect 6559 3037 6615 3778
rect 6559 2981 6910 3037
rect 6409 2936 6496 2943
rect 6409 2881 6425 2936
rect 6484 2881 6496 2936
rect 6409 2868 6496 2881
rect 11028 2909 11155 2923
rect 6568 2796 6894 2840
rect 11028 2833 11039 2909
rect 11139 2833 11155 2909
rect 11028 2821 11155 2833
rect 11212 2918 11321 4448
rect 13774 4095 13910 4104
rect 13774 4019 13783 4095
rect 13893 4019 13910 4095
rect 11845 3245 12035 3262
rect 11845 3056 11862 3245
rect 12020 3056 12035 3245
rect 11845 3040 12035 3056
rect 11212 2842 11221 2918
rect 11300 2842 11321 2918
rect 11212 2831 11321 2842
rect 6523 2784 6894 2796
rect 6523 2738 6777 2784
rect 6523 2275 6624 2738
rect 11607 2345 11692 2348
rect 11607 2292 11622 2345
rect 11679 2343 11692 2345
rect 11679 2292 11694 2343
rect 11411 2277 11513 2283
rect 11411 2275 11423 2277
rect 6523 2224 11423 2275
rect 11501 2275 11513 2277
rect 11501 2224 11516 2275
rect 6523 2219 11516 2224
rect 6523 2214 11513 2219
rect 6523 2137 11471 2214
rect 6523 2133 9039 2137
rect 5916 2089 6309 2095
rect 5845 2008 6309 2089
rect 5845 2001 5972 2008
rect 5845 1732 5944 2001
rect 3076 1657 3374 1714
rect 5845 1713 6197 1732
rect 3076 1584 3133 1657
rect 5845 1656 6204 1713
rect 5845 1633 6197 1656
rect 349 968 417 1523
rect 2657 1475 3133 1584
rect 3386 1592 3490 1601
rect 3386 1528 3395 1592
rect 3477 1528 3490 1592
rect 3386 1518 3490 1528
rect 2638 1418 3133 1475
rect 349 909 356 968
rect 410 909 417 968
rect 349 513 417 909
rect 3387 1001 3451 1518
rect 5845 1515 5944 1633
rect 5674 1416 5944 1515
rect 6464 1591 6553 1600
rect 6464 1527 6478 1591
rect 6543 1527 6553 1591
rect 8939 1576 9039 2133
rect 6464 1517 6553 1527
rect 8799 1563 9039 1576
rect 3387 930 3390 1001
rect 3445 930 3451 1001
rect 1358 597 1451 607
rect 1358 532 1365 597
rect 1437 588 1451 597
rect 1439 536 1451 588
rect 1437 532 1451 536
rect 1358 523 1451 532
rect 3387 520 3451 930
rect 6464 979 6542 1517
rect 8799 1445 9034 1563
rect 6464 915 6471 979
rect 6536 915 6542 979
rect 4390 608 4483 611
rect 4390 605 4484 608
rect 4390 539 4398 605
rect 4470 598 4484 605
rect 4477 544 4484 598
rect 4470 539 4484 544
rect 4390 531 4484 539
rect 4390 530 4483 531
rect 349 500 440 513
rect 349 441 360 500
rect 414 441 440 500
rect 3387 510 3459 520
rect 3387 458 3396 510
rect 3449 458 3459 510
rect 3387 450 3459 458
rect 6464 506 6542 915
rect 8887 989 9478 998
rect 8887 908 8899 989
rect 8967 985 9478 989
rect 8967 908 9376 985
rect 8887 904 9376 908
rect 9444 904 9478 985
rect 8887 897 9478 904
rect 7470 601 7558 606
rect 7470 536 7480 601
rect 7548 594 7558 601
rect 7553 542 7558 594
rect 7548 536 7558 542
rect 7470 530 7558 536
rect 349 426 440 441
rect 6464 446 6475 506
rect 6532 446 6542 506
rect 6464 433 6542 446
rect 11607 496 11694 2292
rect 13774 1476 13910 4019
rect 13774 1399 13783 1476
rect 13901 1399 13910 1476
rect 13774 1388 13910 1399
rect 11607 488 13711 496
rect 11607 410 13597 488
rect 13700 410 13711 488
rect 11607 409 13711 410
rect 13587 400 13711 409
<< via2 >>
rect 5747 4473 5860 4477
rect 5747 4392 5750 4473
rect 5750 4392 5855 4473
rect 5855 4392 5860 4473
rect 5747 4387 5860 4392
rect 1258 3864 1329 3874
rect 1258 3812 1315 3864
rect 1315 3812 1329 3864
rect 1258 3804 1329 3812
rect 4319 3864 4390 3874
rect 4319 3812 4322 3864
rect 4322 3812 4374 3864
rect 4374 3812 4390 3864
rect 4319 3804 4390 3812
rect 5732 2829 5836 2832
rect 5732 2765 5766 2829
rect 5766 2765 5832 2829
rect 5832 2765 5836 2829
rect 5732 2762 5836 2765
rect 11039 2902 11139 2909
rect 11039 2840 11047 2902
rect 11047 2840 11135 2902
rect 11135 2840 11139 2902
rect 11039 2833 11139 2840
rect 11862 3236 12020 3245
rect 11862 3069 11867 3236
rect 11867 3069 12009 3236
rect 12009 3069 12020 3236
rect 11862 3056 12020 3069
rect 1365 588 1437 597
rect 1365 536 1374 588
rect 1374 536 1437 588
rect 1365 532 1437 536
rect 4398 598 4470 605
rect 4398 544 4415 598
rect 4415 544 4470 598
rect 4398 539 4470 544
rect 7480 594 7548 601
rect 7480 542 7487 594
rect 7487 542 7548 594
rect 7480 536 7548 542
<< metal3 >>
rect 5739 4477 5871 4532
rect 5739 4387 5747 4477
rect 5860 4387 5871 4477
rect 5739 4380 5871 4387
rect 1248 3881 1338 3884
rect 1248 3874 4401 3881
rect 1248 3804 1258 3874
rect 1329 3804 4319 3874
rect 4390 3804 4401 3874
rect 1248 3800 4401 3804
rect 1248 3793 1338 3800
rect 2679 3241 2755 3800
rect 2679 3165 3008 3241
rect 2932 2236 3008 3165
rect 5759 2836 5848 4380
rect 11845 3245 12035 3262
rect 11845 3161 11862 3245
rect 11031 3056 11862 3161
rect 12020 3056 12035 3245
rect 11031 3044 12035 3056
rect 11031 2923 11148 3044
rect 11845 3040 12035 3044
rect 5721 2832 5848 2836
rect 5721 2762 5732 2832
rect 5836 2762 5848 2832
rect 11028 2909 11155 2923
rect 11028 2833 11039 2909
rect 11139 2833 11155 2909
rect 11028 2821 11155 2833
rect 5721 2760 5848 2762
rect 5721 2757 5847 2760
rect 5721 2756 5838 2757
rect 11031 2236 11148 2821
rect 2932 2119 11148 2236
rect 1358 606 1451 607
rect 2932 606 3008 2119
rect 4389 606 4483 611
rect 1358 605 7568 606
rect 1358 597 4398 605
rect 1358 532 1365 597
rect 1437 539 4398 597
rect 4470 601 7568 605
rect 4470 539 7480 601
rect 1437 536 7480 539
rect 7548 536 7568 601
rect 1437 532 7568 536
rect 1358 530 7568 532
rect 1358 523 1451 530
use and_5_mag  and_5_mag_0
timestamp 1714558667
transform 1 0 6132 0 1 3071
box 564 403 4618 1596
use Buffer_Delayed1_mag  Buffer_Delayed1_mag_0
timestamp 1714534647
transform 1 0 9363 0 1 97
box -147 -111 4363 1747
use JK_FF_mag  JK_FF_mag_0
timestamp 1714558667
transform 1 0 278 0 1 -16
box -430 0 2603 2148
use JK_FF_mag  JK_FF_mag_1
timestamp 1714558667
transform 1 0 3320 0 1 -7
box -430 0 2603 2148
use JK_FF_mag  JK_FF_mag_2
timestamp 1714558667
transform -1 0 2411 0 -1 4415
box -430 0 2603 2148
use JK_FF_mag  JK_FF_mag_3
timestamp 1714558667
transform -1 0 5471 0 -1 4414
box -430 0 2603 2148
use JK_FF_mag  JK_FF_mag_4
timestamp 1714558667
transform 1 0 6392 0 1 -8
box -430 0 2603 2148
use nand_5_mag  nand_5_mag_0
timestamp 1714558667
transform 1 0 6695 0 -1 3475
box 0 -1 4454 1193
use or_2_mag  or_2_mag_0
timestamp 1714558667
transform 1 0 10970 0 1 1407
box 330 510 1401 1521
<< labels >>
flabel metal1 6001 -85 6001 -85 0 FreeSans 640 0 0 0 VSS
port 0 nsew
flabel metal1 10850 4562 10850 4562 0 FreeSans 640 0 0 0 VDD
port 1 nsew
flabel via2 11925 3147 11925 3147 0 FreeSans 640 0 0 0 RST
port 2 nsew
flabel metal1 12512 2277 12512 2277 0 FreeSans 640 0 0 0 Vdiv31
port 3 nsew
flabel via2 5797 4438 5797 4438 0 FreeSans 640 0 0 0 CLK
port 4 nsew
flabel metal2 3093 2853 3093 2853 0 FreeSans 640 0 0 0 Q0
port 5 nsew
flabel metal2 32 2854 32 2854 0 FreeSans 640 0 0 0 Q1
port 6 nsew
flabel metal2 2661 1549 2661 1549 0 FreeSans 640 0 0 0 Q2
port 7 nsew
flabel metal1 5686 1554 5686 1554 0 FreeSans 640 0 0 0 Q3
port 8 nsew
flabel metal1 8757 1552 8757 1552 0 FreeSans 640 0 0 0 Q4
port 9 nsew
<< end >>
