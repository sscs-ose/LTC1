magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2208 -2120 7960 3120
<< nwell >>
rect -208 -120 5960 1120
<< mvpmos >>
rect 0 0 140 1000
rect 244 0 384 1000
rect 488 0 628 1000
rect 732 0 872 1000
rect 976 0 1116 1000
rect 1220 0 1360 1000
rect 1464 0 1604 1000
rect 1708 0 1848 1000
rect 1952 0 2092 1000
rect 2196 0 2336 1000
rect 2440 0 2580 1000
rect 2684 0 2824 1000
rect 2928 0 3068 1000
rect 3172 0 3312 1000
rect 3416 0 3556 1000
rect 3660 0 3800 1000
rect 3904 0 4044 1000
rect 4148 0 4288 1000
rect 4392 0 4532 1000
rect 4636 0 4776 1000
rect 4880 0 5020 1000
rect 5124 0 5264 1000
rect 5368 0 5508 1000
rect 5612 0 5752 1000
<< mvpdiff >>
rect -88 987 0 1000
rect -88 941 -75 987
rect -29 941 0 987
rect -88 884 0 941
rect -88 838 -75 884
rect -29 838 0 884
rect -88 781 0 838
rect -88 735 -75 781
rect -29 735 0 781
rect -88 678 0 735
rect -88 632 -75 678
rect -29 632 0 678
rect -88 575 0 632
rect -88 529 -75 575
rect -29 529 0 575
rect -88 472 0 529
rect -88 426 -75 472
rect -29 426 0 472
rect -88 369 0 426
rect -88 323 -75 369
rect -29 323 0 369
rect -88 266 0 323
rect -88 220 -75 266
rect -29 220 0 266
rect -88 163 0 220
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 987 244 1000
rect 140 941 169 987
rect 215 941 244 987
rect 140 884 244 941
rect 140 838 169 884
rect 215 838 244 884
rect 140 781 244 838
rect 140 735 169 781
rect 215 735 244 781
rect 140 678 244 735
rect 140 632 169 678
rect 215 632 244 678
rect 140 575 244 632
rect 140 529 169 575
rect 215 529 244 575
rect 140 472 244 529
rect 140 426 169 472
rect 215 426 244 472
rect 140 369 244 426
rect 140 323 169 369
rect 215 323 244 369
rect 140 266 244 323
rect 140 220 169 266
rect 215 220 244 266
rect 140 163 244 220
rect 140 117 169 163
rect 215 117 244 163
rect 140 59 244 117
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 987 488 1000
rect 384 941 413 987
rect 459 941 488 987
rect 384 884 488 941
rect 384 838 413 884
rect 459 838 488 884
rect 384 781 488 838
rect 384 735 413 781
rect 459 735 488 781
rect 384 678 488 735
rect 384 632 413 678
rect 459 632 488 678
rect 384 575 488 632
rect 384 529 413 575
rect 459 529 488 575
rect 384 472 488 529
rect 384 426 413 472
rect 459 426 488 472
rect 384 369 488 426
rect 384 323 413 369
rect 459 323 488 369
rect 384 266 488 323
rect 384 220 413 266
rect 459 220 488 266
rect 384 163 488 220
rect 384 117 413 163
rect 459 117 488 163
rect 384 59 488 117
rect 384 13 413 59
rect 459 13 488 59
rect 384 0 488 13
rect 628 987 732 1000
rect 628 941 657 987
rect 703 941 732 987
rect 628 884 732 941
rect 628 838 657 884
rect 703 838 732 884
rect 628 781 732 838
rect 628 735 657 781
rect 703 735 732 781
rect 628 678 732 735
rect 628 632 657 678
rect 703 632 732 678
rect 628 575 732 632
rect 628 529 657 575
rect 703 529 732 575
rect 628 472 732 529
rect 628 426 657 472
rect 703 426 732 472
rect 628 369 732 426
rect 628 323 657 369
rect 703 323 732 369
rect 628 266 732 323
rect 628 220 657 266
rect 703 220 732 266
rect 628 163 732 220
rect 628 117 657 163
rect 703 117 732 163
rect 628 59 732 117
rect 628 13 657 59
rect 703 13 732 59
rect 628 0 732 13
rect 872 987 976 1000
rect 872 941 901 987
rect 947 941 976 987
rect 872 884 976 941
rect 872 838 901 884
rect 947 838 976 884
rect 872 781 976 838
rect 872 735 901 781
rect 947 735 976 781
rect 872 678 976 735
rect 872 632 901 678
rect 947 632 976 678
rect 872 575 976 632
rect 872 529 901 575
rect 947 529 976 575
rect 872 472 976 529
rect 872 426 901 472
rect 947 426 976 472
rect 872 369 976 426
rect 872 323 901 369
rect 947 323 976 369
rect 872 266 976 323
rect 872 220 901 266
rect 947 220 976 266
rect 872 163 976 220
rect 872 117 901 163
rect 947 117 976 163
rect 872 59 976 117
rect 872 13 901 59
rect 947 13 976 59
rect 872 0 976 13
rect 1116 987 1220 1000
rect 1116 941 1145 987
rect 1191 941 1220 987
rect 1116 884 1220 941
rect 1116 838 1145 884
rect 1191 838 1220 884
rect 1116 781 1220 838
rect 1116 735 1145 781
rect 1191 735 1220 781
rect 1116 678 1220 735
rect 1116 632 1145 678
rect 1191 632 1220 678
rect 1116 575 1220 632
rect 1116 529 1145 575
rect 1191 529 1220 575
rect 1116 472 1220 529
rect 1116 426 1145 472
rect 1191 426 1220 472
rect 1116 369 1220 426
rect 1116 323 1145 369
rect 1191 323 1220 369
rect 1116 266 1220 323
rect 1116 220 1145 266
rect 1191 220 1220 266
rect 1116 163 1220 220
rect 1116 117 1145 163
rect 1191 117 1220 163
rect 1116 59 1220 117
rect 1116 13 1145 59
rect 1191 13 1220 59
rect 1116 0 1220 13
rect 1360 987 1464 1000
rect 1360 941 1389 987
rect 1435 941 1464 987
rect 1360 884 1464 941
rect 1360 838 1389 884
rect 1435 838 1464 884
rect 1360 781 1464 838
rect 1360 735 1389 781
rect 1435 735 1464 781
rect 1360 678 1464 735
rect 1360 632 1389 678
rect 1435 632 1464 678
rect 1360 575 1464 632
rect 1360 529 1389 575
rect 1435 529 1464 575
rect 1360 472 1464 529
rect 1360 426 1389 472
rect 1435 426 1464 472
rect 1360 369 1464 426
rect 1360 323 1389 369
rect 1435 323 1464 369
rect 1360 266 1464 323
rect 1360 220 1389 266
rect 1435 220 1464 266
rect 1360 163 1464 220
rect 1360 117 1389 163
rect 1435 117 1464 163
rect 1360 59 1464 117
rect 1360 13 1389 59
rect 1435 13 1464 59
rect 1360 0 1464 13
rect 1604 987 1708 1000
rect 1604 941 1633 987
rect 1679 941 1708 987
rect 1604 884 1708 941
rect 1604 838 1633 884
rect 1679 838 1708 884
rect 1604 781 1708 838
rect 1604 735 1633 781
rect 1679 735 1708 781
rect 1604 678 1708 735
rect 1604 632 1633 678
rect 1679 632 1708 678
rect 1604 575 1708 632
rect 1604 529 1633 575
rect 1679 529 1708 575
rect 1604 472 1708 529
rect 1604 426 1633 472
rect 1679 426 1708 472
rect 1604 369 1708 426
rect 1604 323 1633 369
rect 1679 323 1708 369
rect 1604 266 1708 323
rect 1604 220 1633 266
rect 1679 220 1708 266
rect 1604 163 1708 220
rect 1604 117 1633 163
rect 1679 117 1708 163
rect 1604 59 1708 117
rect 1604 13 1633 59
rect 1679 13 1708 59
rect 1604 0 1708 13
rect 1848 987 1952 1000
rect 1848 941 1877 987
rect 1923 941 1952 987
rect 1848 884 1952 941
rect 1848 838 1877 884
rect 1923 838 1952 884
rect 1848 781 1952 838
rect 1848 735 1877 781
rect 1923 735 1952 781
rect 1848 678 1952 735
rect 1848 632 1877 678
rect 1923 632 1952 678
rect 1848 575 1952 632
rect 1848 529 1877 575
rect 1923 529 1952 575
rect 1848 472 1952 529
rect 1848 426 1877 472
rect 1923 426 1952 472
rect 1848 369 1952 426
rect 1848 323 1877 369
rect 1923 323 1952 369
rect 1848 266 1952 323
rect 1848 220 1877 266
rect 1923 220 1952 266
rect 1848 163 1952 220
rect 1848 117 1877 163
rect 1923 117 1952 163
rect 1848 59 1952 117
rect 1848 13 1877 59
rect 1923 13 1952 59
rect 1848 0 1952 13
rect 2092 987 2196 1000
rect 2092 941 2121 987
rect 2167 941 2196 987
rect 2092 884 2196 941
rect 2092 838 2121 884
rect 2167 838 2196 884
rect 2092 781 2196 838
rect 2092 735 2121 781
rect 2167 735 2196 781
rect 2092 678 2196 735
rect 2092 632 2121 678
rect 2167 632 2196 678
rect 2092 575 2196 632
rect 2092 529 2121 575
rect 2167 529 2196 575
rect 2092 472 2196 529
rect 2092 426 2121 472
rect 2167 426 2196 472
rect 2092 369 2196 426
rect 2092 323 2121 369
rect 2167 323 2196 369
rect 2092 266 2196 323
rect 2092 220 2121 266
rect 2167 220 2196 266
rect 2092 163 2196 220
rect 2092 117 2121 163
rect 2167 117 2196 163
rect 2092 59 2196 117
rect 2092 13 2121 59
rect 2167 13 2196 59
rect 2092 0 2196 13
rect 2336 987 2440 1000
rect 2336 941 2365 987
rect 2411 941 2440 987
rect 2336 884 2440 941
rect 2336 838 2365 884
rect 2411 838 2440 884
rect 2336 781 2440 838
rect 2336 735 2365 781
rect 2411 735 2440 781
rect 2336 678 2440 735
rect 2336 632 2365 678
rect 2411 632 2440 678
rect 2336 575 2440 632
rect 2336 529 2365 575
rect 2411 529 2440 575
rect 2336 472 2440 529
rect 2336 426 2365 472
rect 2411 426 2440 472
rect 2336 369 2440 426
rect 2336 323 2365 369
rect 2411 323 2440 369
rect 2336 266 2440 323
rect 2336 220 2365 266
rect 2411 220 2440 266
rect 2336 163 2440 220
rect 2336 117 2365 163
rect 2411 117 2440 163
rect 2336 59 2440 117
rect 2336 13 2365 59
rect 2411 13 2440 59
rect 2336 0 2440 13
rect 2580 987 2684 1000
rect 2580 941 2609 987
rect 2655 941 2684 987
rect 2580 884 2684 941
rect 2580 838 2609 884
rect 2655 838 2684 884
rect 2580 781 2684 838
rect 2580 735 2609 781
rect 2655 735 2684 781
rect 2580 678 2684 735
rect 2580 632 2609 678
rect 2655 632 2684 678
rect 2580 575 2684 632
rect 2580 529 2609 575
rect 2655 529 2684 575
rect 2580 472 2684 529
rect 2580 426 2609 472
rect 2655 426 2684 472
rect 2580 369 2684 426
rect 2580 323 2609 369
rect 2655 323 2684 369
rect 2580 266 2684 323
rect 2580 220 2609 266
rect 2655 220 2684 266
rect 2580 163 2684 220
rect 2580 117 2609 163
rect 2655 117 2684 163
rect 2580 59 2684 117
rect 2580 13 2609 59
rect 2655 13 2684 59
rect 2580 0 2684 13
rect 2824 987 2928 1000
rect 2824 941 2853 987
rect 2899 941 2928 987
rect 2824 884 2928 941
rect 2824 838 2853 884
rect 2899 838 2928 884
rect 2824 781 2928 838
rect 2824 735 2853 781
rect 2899 735 2928 781
rect 2824 678 2928 735
rect 2824 632 2853 678
rect 2899 632 2928 678
rect 2824 575 2928 632
rect 2824 529 2853 575
rect 2899 529 2928 575
rect 2824 472 2928 529
rect 2824 426 2853 472
rect 2899 426 2928 472
rect 2824 369 2928 426
rect 2824 323 2853 369
rect 2899 323 2928 369
rect 2824 266 2928 323
rect 2824 220 2853 266
rect 2899 220 2928 266
rect 2824 163 2928 220
rect 2824 117 2853 163
rect 2899 117 2928 163
rect 2824 59 2928 117
rect 2824 13 2853 59
rect 2899 13 2928 59
rect 2824 0 2928 13
rect 3068 987 3172 1000
rect 3068 941 3097 987
rect 3143 941 3172 987
rect 3068 884 3172 941
rect 3068 838 3097 884
rect 3143 838 3172 884
rect 3068 781 3172 838
rect 3068 735 3097 781
rect 3143 735 3172 781
rect 3068 678 3172 735
rect 3068 632 3097 678
rect 3143 632 3172 678
rect 3068 575 3172 632
rect 3068 529 3097 575
rect 3143 529 3172 575
rect 3068 472 3172 529
rect 3068 426 3097 472
rect 3143 426 3172 472
rect 3068 369 3172 426
rect 3068 323 3097 369
rect 3143 323 3172 369
rect 3068 266 3172 323
rect 3068 220 3097 266
rect 3143 220 3172 266
rect 3068 163 3172 220
rect 3068 117 3097 163
rect 3143 117 3172 163
rect 3068 59 3172 117
rect 3068 13 3097 59
rect 3143 13 3172 59
rect 3068 0 3172 13
rect 3312 987 3416 1000
rect 3312 941 3341 987
rect 3387 941 3416 987
rect 3312 884 3416 941
rect 3312 838 3341 884
rect 3387 838 3416 884
rect 3312 781 3416 838
rect 3312 735 3341 781
rect 3387 735 3416 781
rect 3312 678 3416 735
rect 3312 632 3341 678
rect 3387 632 3416 678
rect 3312 575 3416 632
rect 3312 529 3341 575
rect 3387 529 3416 575
rect 3312 472 3416 529
rect 3312 426 3341 472
rect 3387 426 3416 472
rect 3312 369 3416 426
rect 3312 323 3341 369
rect 3387 323 3416 369
rect 3312 266 3416 323
rect 3312 220 3341 266
rect 3387 220 3416 266
rect 3312 163 3416 220
rect 3312 117 3341 163
rect 3387 117 3416 163
rect 3312 59 3416 117
rect 3312 13 3341 59
rect 3387 13 3416 59
rect 3312 0 3416 13
rect 3556 987 3660 1000
rect 3556 941 3585 987
rect 3631 941 3660 987
rect 3556 884 3660 941
rect 3556 838 3585 884
rect 3631 838 3660 884
rect 3556 781 3660 838
rect 3556 735 3585 781
rect 3631 735 3660 781
rect 3556 678 3660 735
rect 3556 632 3585 678
rect 3631 632 3660 678
rect 3556 575 3660 632
rect 3556 529 3585 575
rect 3631 529 3660 575
rect 3556 472 3660 529
rect 3556 426 3585 472
rect 3631 426 3660 472
rect 3556 369 3660 426
rect 3556 323 3585 369
rect 3631 323 3660 369
rect 3556 266 3660 323
rect 3556 220 3585 266
rect 3631 220 3660 266
rect 3556 163 3660 220
rect 3556 117 3585 163
rect 3631 117 3660 163
rect 3556 59 3660 117
rect 3556 13 3585 59
rect 3631 13 3660 59
rect 3556 0 3660 13
rect 3800 987 3904 1000
rect 3800 941 3829 987
rect 3875 941 3904 987
rect 3800 884 3904 941
rect 3800 838 3829 884
rect 3875 838 3904 884
rect 3800 781 3904 838
rect 3800 735 3829 781
rect 3875 735 3904 781
rect 3800 678 3904 735
rect 3800 632 3829 678
rect 3875 632 3904 678
rect 3800 575 3904 632
rect 3800 529 3829 575
rect 3875 529 3904 575
rect 3800 472 3904 529
rect 3800 426 3829 472
rect 3875 426 3904 472
rect 3800 369 3904 426
rect 3800 323 3829 369
rect 3875 323 3904 369
rect 3800 266 3904 323
rect 3800 220 3829 266
rect 3875 220 3904 266
rect 3800 163 3904 220
rect 3800 117 3829 163
rect 3875 117 3904 163
rect 3800 59 3904 117
rect 3800 13 3829 59
rect 3875 13 3904 59
rect 3800 0 3904 13
rect 4044 987 4148 1000
rect 4044 941 4073 987
rect 4119 941 4148 987
rect 4044 884 4148 941
rect 4044 838 4073 884
rect 4119 838 4148 884
rect 4044 781 4148 838
rect 4044 735 4073 781
rect 4119 735 4148 781
rect 4044 678 4148 735
rect 4044 632 4073 678
rect 4119 632 4148 678
rect 4044 575 4148 632
rect 4044 529 4073 575
rect 4119 529 4148 575
rect 4044 472 4148 529
rect 4044 426 4073 472
rect 4119 426 4148 472
rect 4044 369 4148 426
rect 4044 323 4073 369
rect 4119 323 4148 369
rect 4044 266 4148 323
rect 4044 220 4073 266
rect 4119 220 4148 266
rect 4044 163 4148 220
rect 4044 117 4073 163
rect 4119 117 4148 163
rect 4044 59 4148 117
rect 4044 13 4073 59
rect 4119 13 4148 59
rect 4044 0 4148 13
rect 4288 987 4392 1000
rect 4288 941 4317 987
rect 4363 941 4392 987
rect 4288 884 4392 941
rect 4288 838 4317 884
rect 4363 838 4392 884
rect 4288 781 4392 838
rect 4288 735 4317 781
rect 4363 735 4392 781
rect 4288 678 4392 735
rect 4288 632 4317 678
rect 4363 632 4392 678
rect 4288 575 4392 632
rect 4288 529 4317 575
rect 4363 529 4392 575
rect 4288 472 4392 529
rect 4288 426 4317 472
rect 4363 426 4392 472
rect 4288 369 4392 426
rect 4288 323 4317 369
rect 4363 323 4392 369
rect 4288 266 4392 323
rect 4288 220 4317 266
rect 4363 220 4392 266
rect 4288 163 4392 220
rect 4288 117 4317 163
rect 4363 117 4392 163
rect 4288 59 4392 117
rect 4288 13 4317 59
rect 4363 13 4392 59
rect 4288 0 4392 13
rect 4532 987 4636 1000
rect 4532 941 4561 987
rect 4607 941 4636 987
rect 4532 884 4636 941
rect 4532 838 4561 884
rect 4607 838 4636 884
rect 4532 781 4636 838
rect 4532 735 4561 781
rect 4607 735 4636 781
rect 4532 678 4636 735
rect 4532 632 4561 678
rect 4607 632 4636 678
rect 4532 575 4636 632
rect 4532 529 4561 575
rect 4607 529 4636 575
rect 4532 472 4636 529
rect 4532 426 4561 472
rect 4607 426 4636 472
rect 4532 369 4636 426
rect 4532 323 4561 369
rect 4607 323 4636 369
rect 4532 266 4636 323
rect 4532 220 4561 266
rect 4607 220 4636 266
rect 4532 163 4636 220
rect 4532 117 4561 163
rect 4607 117 4636 163
rect 4532 59 4636 117
rect 4532 13 4561 59
rect 4607 13 4636 59
rect 4532 0 4636 13
rect 4776 987 4880 1000
rect 4776 941 4805 987
rect 4851 941 4880 987
rect 4776 884 4880 941
rect 4776 838 4805 884
rect 4851 838 4880 884
rect 4776 781 4880 838
rect 4776 735 4805 781
rect 4851 735 4880 781
rect 4776 678 4880 735
rect 4776 632 4805 678
rect 4851 632 4880 678
rect 4776 575 4880 632
rect 4776 529 4805 575
rect 4851 529 4880 575
rect 4776 472 4880 529
rect 4776 426 4805 472
rect 4851 426 4880 472
rect 4776 369 4880 426
rect 4776 323 4805 369
rect 4851 323 4880 369
rect 4776 266 4880 323
rect 4776 220 4805 266
rect 4851 220 4880 266
rect 4776 163 4880 220
rect 4776 117 4805 163
rect 4851 117 4880 163
rect 4776 59 4880 117
rect 4776 13 4805 59
rect 4851 13 4880 59
rect 4776 0 4880 13
rect 5020 987 5124 1000
rect 5020 941 5049 987
rect 5095 941 5124 987
rect 5020 884 5124 941
rect 5020 838 5049 884
rect 5095 838 5124 884
rect 5020 781 5124 838
rect 5020 735 5049 781
rect 5095 735 5124 781
rect 5020 678 5124 735
rect 5020 632 5049 678
rect 5095 632 5124 678
rect 5020 575 5124 632
rect 5020 529 5049 575
rect 5095 529 5124 575
rect 5020 472 5124 529
rect 5020 426 5049 472
rect 5095 426 5124 472
rect 5020 369 5124 426
rect 5020 323 5049 369
rect 5095 323 5124 369
rect 5020 266 5124 323
rect 5020 220 5049 266
rect 5095 220 5124 266
rect 5020 163 5124 220
rect 5020 117 5049 163
rect 5095 117 5124 163
rect 5020 59 5124 117
rect 5020 13 5049 59
rect 5095 13 5124 59
rect 5020 0 5124 13
rect 5264 987 5368 1000
rect 5264 941 5293 987
rect 5339 941 5368 987
rect 5264 884 5368 941
rect 5264 838 5293 884
rect 5339 838 5368 884
rect 5264 781 5368 838
rect 5264 735 5293 781
rect 5339 735 5368 781
rect 5264 678 5368 735
rect 5264 632 5293 678
rect 5339 632 5368 678
rect 5264 575 5368 632
rect 5264 529 5293 575
rect 5339 529 5368 575
rect 5264 472 5368 529
rect 5264 426 5293 472
rect 5339 426 5368 472
rect 5264 369 5368 426
rect 5264 323 5293 369
rect 5339 323 5368 369
rect 5264 266 5368 323
rect 5264 220 5293 266
rect 5339 220 5368 266
rect 5264 163 5368 220
rect 5264 117 5293 163
rect 5339 117 5368 163
rect 5264 59 5368 117
rect 5264 13 5293 59
rect 5339 13 5368 59
rect 5264 0 5368 13
rect 5508 987 5612 1000
rect 5508 941 5537 987
rect 5583 941 5612 987
rect 5508 884 5612 941
rect 5508 838 5537 884
rect 5583 838 5612 884
rect 5508 781 5612 838
rect 5508 735 5537 781
rect 5583 735 5612 781
rect 5508 678 5612 735
rect 5508 632 5537 678
rect 5583 632 5612 678
rect 5508 575 5612 632
rect 5508 529 5537 575
rect 5583 529 5612 575
rect 5508 472 5612 529
rect 5508 426 5537 472
rect 5583 426 5612 472
rect 5508 369 5612 426
rect 5508 323 5537 369
rect 5583 323 5612 369
rect 5508 266 5612 323
rect 5508 220 5537 266
rect 5583 220 5612 266
rect 5508 163 5612 220
rect 5508 117 5537 163
rect 5583 117 5612 163
rect 5508 59 5612 117
rect 5508 13 5537 59
rect 5583 13 5612 59
rect 5508 0 5612 13
rect 5752 987 5840 1000
rect 5752 941 5781 987
rect 5827 941 5840 987
rect 5752 884 5840 941
rect 5752 838 5781 884
rect 5827 838 5840 884
rect 5752 781 5840 838
rect 5752 735 5781 781
rect 5827 735 5840 781
rect 5752 678 5840 735
rect 5752 632 5781 678
rect 5827 632 5840 678
rect 5752 575 5840 632
rect 5752 529 5781 575
rect 5827 529 5840 575
rect 5752 472 5840 529
rect 5752 426 5781 472
rect 5827 426 5840 472
rect 5752 369 5840 426
rect 5752 323 5781 369
rect 5827 323 5840 369
rect 5752 266 5840 323
rect 5752 220 5781 266
rect 5827 220 5840 266
rect 5752 163 5840 220
rect 5752 117 5781 163
rect 5827 117 5840 163
rect 5752 59 5840 117
rect 5752 13 5781 59
rect 5827 13 5840 59
rect 5752 0 5840 13
<< mvpdiffc >>
rect -75 941 -29 987
rect -75 838 -29 884
rect -75 735 -29 781
rect -75 632 -29 678
rect -75 529 -29 575
rect -75 426 -29 472
rect -75 323 -29 369
rect -75 220 -29 266
rect -75 117 -29 163
rect -75 13 -29 59
rect 169 941 215 987
rect 169 838 215 884
rect 169 735 215 781
rect 169 632 215 678
rect 169 529 215 575
rect 169 426 215 472
rect 169 323 215 369
rect 169 220 215 266
rect 169 117 215 163
rect 169 13 215 59
rect 413 941 459 987
rect 413 838 459 884
rect 413 735 459 781
rect 413 632 459 678
rect 413 529 459 575
rect 413 426 459 472
rect 413 323 459 369
rect 413 220 459 266
rect 413 117 459 163
rect 413 13 459 59
rect 657 941 703 987
rect 657 838 703 884
rect 657 735 703 781
rect 657 632 703 678
rect 657 529 703 575
rect 657 426 703 472
rect 657 323 703 369
rect 657 220 703 266
rect 657 117 703 163
rect 657 13 703 59
rect 901 941 947 987
rect 901 838 947 884
rect 901 735 947 781
rect 901 632 947 678
rect 901 529 947 575
rect 901 426 947 472
rect 901 323 947 369
rect 901 220 947 266
rect 901 117 947 163
rect 901 13 947 59
rect 1145 941 1191 987
rect 1145 838 1191 884
rect 1145 735 1191 781
rect 1145 632 1191 678
rect 1145 529 1191 575
rect 1145 426 1191 472
rect 1145 323 1191 369
rect 1145 220 1191 266
rect 1145 117 1191 163
rect 1145 13 1191 59
rect 1389 941 1435 987
rect 1389 838 1435 884
rect 1389 735 1435 781
rect 1389 632 1435 678
rect 1389 529 1435 575
rect 1389 426 1435 472
rect 1389 323 1435 369
rect 1389 220 1435 266
rect 1389 117 1435 163
rect 1389 13 1435 59
rect 1633 941 1679 987
rect 1633 838 1679 884
rect 1633 735 1679 781
rect 1633 632 1679 678
rect 1633 529 1679 575
rect 1633 426 1679 472
rect 1633 323 1679 369
rect 1633 220 1679 266
rect 1633 117 1679 163
rect 1633 13 1679 59
rect 1877 941 1923 987
rect 1877 838 1923 884
rect 1877 735 1923 781
rect 1877 632 1923 678
rect 1877 529 1923 575
rect 1877 426 1923 472
rect 1877 323 1923 369
rect 1877 220 1923 266
rect 1877 117 1923 163
rect 1877 13 1923 59
rect 2121 941 2167 987
rect 2121 838 2167 884
rect 2121 735 2167 781
rect 2121 632 2167 678
rect 2121 529 2167 575
rect 2121 426 2167 472
rect 2121 323 2167 369
rect 2121 220 2167 266
rect 2121 117 2167 163
rect 2121 13 2167 59
rect 2365 941 2411 987
rect 2365 838 2411 884
rect 2365 735 2411 781
rect 2365 632 2411 678
rect 2365 529 2411 575
rect 2365 426 2411 472
rect 2365 323 2411 369
rect 2365 220 2411 266
rect 2365 117 2411 163
rect 2365 13 2411 59
rect 2609 941 2655 987
rect 2609 838 2655 884
rect 2609 735 2655 781
rect 2609 632 2655 678
rect 2609 529 2655 575
rect 2609 426 2655 472
rect 2609 323 2655 369
rect 2609 220 2655 266
rect 2609 117 2655 163
rect 2609 13 2655 59
rect 2853 941 2899 987
rect 2853 838 2899 884
rect 2853 735 2899 781
rect 2853 632 2899 678
rect 2853 529 2899 575
rect 2853 426 2899 472
rect 2853 323 2899 369
rect 2853 220 2899 266
rect 2853 117 2899 163
rect 2853 13 2899 59
rect 3097 941 3143 987
rect 3097 838 3143 884
rect 3097 735 3143 781
rect 3097 632 3143 678
rect 3097 529 3143 575
rect 3097 426 3143 472
rect 3097 323 3143 369
rect 3097 220 3143 266
rect 3097 117 3143 163
rect 3097 13 3143 59
rect 3341 941 3387 987
rect 3341 838 3387 884
rect 3341 735 3387 781
rect 3341 632 3387 678
rect 3341 529 3387 575
rect 3341 426 3387 472
rect 3341 323 3387 369
rect 3341 220 3387 266
rect 3341 117 3387 163
rect 3341 13 3387 59
rect 3585 941 3631 987
rect 3585 838 3631 884
rect 3585 735 3631 781
rect 3585 632 3631 678
rect 3585 529 3631 575
rect 3585 426 3631 472
rect 3585 323 3631 369
rect 3585 220 3631 266
rect 3585 117 3631 163
rect 3585 13 3631 59
rect 3829 941 3875 987
rect 3829 838 3875 884
rect 3829 735 3875 781
rect 3829 632 3875 678
rect 3829 529 3875 575
rect 3829 426 3875 472
rect 3829 323 3875 369
rect 3829 220 3875 266
rect 3829 117 3875 163
rect 3829 13 3875 59
rect 4073 941 4119 987
rect 4073 838 4119 884
rect 4073 735 4119 781
rect 4073 632 4119 678
rect 4073 529 4119 575
rect 4073 426 4119 472
rect 4073 323 4119 369
rect 4073 220 4119 266
rect 4073 117 4119 163
rect 4073 13 4119 59
rect 4317 941 4363 987
rect 4317 838 4363 884
rect 4317 735 4363 781
rect 4317 632 4363 678
rect 4317 529 4363 575
rect 4317 426 4363 472
rect 4317 323 4363 369
rect 4317 220 4363 266
rect 4317 117 4363 163
rect 4317 13 4363 59
rect 4561 941 4607 987
rect 4561 838 4607 884
rect 4561 735 4607 781
rect 4561 632 4607 678
rect 4561 529 4607 575
rect 4561 426 4607 472
rect 4561 323 4607 369
rect 4561 220 4607 266
rect 4561 117 4607 163
rect 4561 13 4607 59
rect 4805 941 4851 987
rect 4805 838 4851 884
rect 4805 735 4851 781
rect 4805 632 4851 678
rect 4805 529 4851 575
rect 4805 426 4851 472
rect 4805 323 4851 369
rect 4805 220 4851 266
rect 4805 117 4851 163
rect 4805 13 4851 59
rect 5049 941 5095 987
rect 5049 838 5095 884
rect 5049 735 5095 781
rect 5049 632 5095 678
rect 5049 529 5095 575
rect 5049 426 5095 472
rect 5049 323 5095 369
rect 5049 220 5095 266
rect 5049 117 5095 163
rect 5049 13 5095 59
rect 5293 941 5339 987
rect 5293 838 5339 884
rect 5293 735 5339 781
rect 5293 632 5339 678
rect 5293 529 5339 575
rect 5293 426 5339 472
rect 5293 323 5339 369
rect 5293 220 5339 266
rect 5293 117 5339 163
rect 5293 13 5339 59
rect 5537 941 5583 987
rect 5537 838 5583 884
rect 5537 735 5583 781
rect 5537 632 5583 678
rect 5537 529 5583 575
rect 5537 426 5583 472
rect 5537 323 5583 369
rect 5537 220 5583 266
rect 5537 117 5583 163
rect 5537 13 5583 59
rect 5781 941 5827 987
rect 5781 838 5827 884
rect 5781 735 5827 781
rect 5781 632 5827 678
rect 5781 529 5827 575
rect 5781 426 5827 472
rect 5781 323 5827 369
rect 5781 220 5827 266
rect 5781 117 5827 163
rect 5781 13 5827 59
<< polysilicon >>
rect 0 1000 140 1044
rect 244 1000 384 1044
rect 488 1000 628 1044
rect 732 1000 872 1044
rect 976 1000 1116 1044
rect 1220 1000 1360 1044
rect 1464 1000 1604 1044
rect 1708 1000 1848 1044
rect 1952 1000 2092 1044
rect 2196 1000 2336 1044
rect 2440 1000 2580 1044
rect 2684 1000 2824 1044
rect 2928 1000 3068 1044
rect 3172 1000 3312 1044
rect 3416 1000 3556 1044
rect 3660 1000 3800 1044
rect 3904 1000 4044 1044
rect 4148 1000 4288 1044
rect 4392 1000 4532 1044
rect 4636 1000 4776 1044
rect 4880 1000 5020 1044
rect 5124 1000 5264 1044
rect 5368 1000 5508 1044
rect 5612 1000 5752 1044
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
rect 976 -44 1116 0
rect 1220 -44 1360 0
rect 1464 -44 1604 0
rect 1708 -44 1848 0
rect 1952 -44 2092 0
rect 2196 -44 2336 0
rect 2440 -44 2580 0
rect 2684 -44 2824 0
rect 2928 -44 3068 0
rect 3172 -44 3312 0
rect 3416 -44 3556 0
rect 3660 -44 3800 0
rect 3904 -44 4044 0
rect 4148 -44 4288 0
rect 4392 -44 4532 0
rect 4636 -44 4776 0
rect 4880 -44 5020 0
rect 5124 -44 5264 0
rect 5368 -44 5508 0
rect 5612 -44 5752 0
<< metal1 >>
rect -75 987 -29 1000
rect -75 884 -29 941
rect -75 781 -29 838
rect -75 678 -29 735
rect -75 575 -29 632
rect -75 472 -29 529
rect -75 369 -29 426
rect -75 266 -29 323
rect -75 163 -29 220
rect -75 59 -29 117
rect -75 0 -29 13
rect 169 987 215 1000
rect 169 884 215 941
rect 169 781 215 838
rect 169 678 215 735
rect 169 575 215 632
rect 169 472 215 529
rect 169 369 215 426
rect 169 266 215 323
rect 169 163 215 220
rect 169 59 215 117
rect 169 0 215 13
rect 413 987 459 1000
rect 413 884 459 941
rect 413 781 459 838
rect 413 678 459 735
rect 413 575 459 632
rect 413 472 459 529
rect 413 369 459 426
rect 413 266 459 323
rect 413 163 459 220
rect 413 59 459 117
rect 413 0 459 13
rect 657 987 703 1000
rect 657 884 703 941
rect 657 781 703 838
rect 657 678 703 735
rect 657 575 703 632
rect 657 472 703 529
rect 657 369 703 426
rect 657 266 703 323
rect 657 163 703 220
rect 657 59 703 117
rect 657 0 703 13
rect 901 987 947 1000
rect 901 884 947 941
rect 901 781 947 838
rect 901 678 947 735
rect 901 575 947 632
rect 901 472 947 529
rect 901 369 947 426
rect 901 266 947 323
rect 901 163 947 220
rect 901 59 947 117
rect 901 0 947 13
rect 1145 987 1191 1000
rect 1145 884 1191 941
rect 1145 781 1191 838
rect 1145 678 1191 735
rect 1145 575 1191 632
rect 1145 472 1191 529
rect 1145 369 1191 426
rect 1145 266 1191 323
rect 1145 163 1191 220
rect 1145 59 1191 117
rect 1145 0 1191 13
rect 1389 987 1435 1000
rect 1389 884 1435 941
rect 1389 781 1435 838
rect 1389 678 1435 735
rect 1389 575 1435 632
rect 1389 472 1435 529
rect 1389 369 1435 426
rect 1389 266 1435 323
rect 1389 163 1435 220
rect 1389 59 1435 117
rect 1389 0 1435 13
rect 1633 987 1679 1000
rect 1633 884 1679 941
rect 1633 781 1679 838
rect 1633 678 1679 735
rect 1633 575 1679 632
rect 1633 472 1679 529
rect 1633 369 1679 426
rect 1633 266 1679 323
rect 1633 163 1679 220
rect 1633 59 1679 117
rect 1633 0 1679 13
rect 1877 987 1923 1000
rect 1877 884 1923 941
rect 1877 781 1923 838
rect 1877 678 1923 735
rect 1877 575 1923 632
rect 1877 472 1923 529
rect 1877 369 1923 426
rect 1877 266 1923 323
rect 1877 163 1923 220
rect 1877 59 1923 117
rect 1877 0 1923 13
rect 2121 987 2167 1000
rect 2121 884 2167 941
rect 2121 781 2167 838
rect 2121 678 2167 735
rect 2121 575 2167 632
rect 2121 472 2167 529
rect 2121 369 2167 426
rect 2121 266 2167 323
rect 2121 163 2167 220
rect 2121 59 2167 117
rect 2121 0 2167 13
rect 2365 987 2411 1000
rect 2365 884 2411 941
rect 2365 781 2411 838
rect 2365 678 2411 735
rect 2365 575 2411 632
rect 2365 472 2411 529
rect 2365 369 2411 426
rect 2365 266 2411 323
rect 2365 163 2411 220
rect 2365 59 2411 117
rect 2365 0 2411 13
rect 2609 987 2655 1000
rect 2609 884 2655 941
rect 2609 781 2655 838
rect 2609 678 2655 735
rect 2609 575 2655 632
rect 2609 472 2655 529
rect 2609 369 2655 426
rect 2609 266 2655 323
rect 2609 163 2655 220
rect 2609 59 2655 117
rect 2609 0 2655 13
rect 2853 987 2899 1000
rect 2853 884 2899 941
rect 2853 781 2899 838
rect 2853 678 2899 735
rect 2853 575 2899 632
rect 2853 472 2899 529
rect 2853 369 2899 426
rect 2853 266 2899 323
rect 2853 163 2899 220
rect 2853 59 2899 117
rect 2853 0 2899 13
rect 3097 987 3143 1000
rect 3097 884 3143 941
rect 3097 781 3143 838
rect 3097 678 3143 735
rect 3097 575 3143 632
rect 3097 472 3143 529
rect 3097 369 3143 426
rect 3097 266 3143 323
rect 3097 163 3143 220
rect 3097 59 3143 117
rect 3097 0 3143 13
rect 3341 987 3387 1000
rect 3341 884 3387 941
rect 3341 781 3387 838
rect 3341 678 3387 735
rect 3341 575 3387 632
rect 3341 472 3387 529
rect 3341 369 3387 426
rect 3341 266 3387 323
rect 3341 163 3387 220
rect 3341 59 3387 117
rect 3341 0 3387 13
rect 3585 987 3631 1000
rect 3585 884 3631 941
rect 3585 781 3631 838
rect 3585 678 3631 735
rect 3585 575 3631 632
rect 3585 472 3631 529
rect 3585 369 3631 426
rect 3585 266 3631 323
rect 3585 163 3631 220
rect 3585 59 3631 117
rect 3585 0 3631 13
rect 3829 987 3875 1000
rect 3829 884 3875 941
rect 3829 781 3875 838
rect 3829 678 3875 735
rect 3829 575 3875 632
rect 3829 472 3875 529
rect 3829 369 3875 426
rect 3829 266 3875 323
rect 3829 163 3875 220
rect 3829 59 3875 117
rect 3829 0 3875 13
rect 4073 987 4119 1000
rect 4073 884 4119 941
rect 4073 781 4119 838
rect 4073 678 4119 735
rect 4073 575 4119 632
rect 4073 472 4119 529
rect 4073 369 4119 426
rect 4073 266 4119 323
rect 4073 163 4119 220
rect 4073 59 4119 117
rect 4073 0 4119 13
rect 4317 987 4363 1000
rect 4317 884 4363 941
rect 4317 781 4363 838
rect 4317 678 4363 735
rect 4317 575 4363 632
rect 4317 472 4363 529
rect 4317 369 4363 426
rect 4317 266 4363 323
rect 4317 163 4363 220
rect 4317 59 4363 117
rect 4317 0 4363 13
rect 4561 987 4607 1000
rect 4561 884 4607 941
rect 4561 781 4607 838
rect 4561 678 4607 735
rect 4561 575 4607 632
rect 4561 472 4607 529
rect 4561 369 4607 426
rect 4561 266 4607 323
rect 4561 163 4607 220
rect 4561 59 4607 117
rect 4561 0 4607 13
rect 4805 987 4851 1000
rect 4805 884 4851 941
rect 4805 781 4851 838
rect 4805 678 4851 735
rect 4805 575 4851 632
rect 4805 472 4851 529
rect 4805 369 4851 426
rect 4805 266 4851 323
rect 4805 163 4851 220
rect 4805 59 4851 117
rect 4805 0 4851 13
rect 5049 987 5095 1000
rect 5049 884 5095 941
rect 5049 781 5095 838
rect 5049 678 5095 735
rect 5049 575 5095 632
rect 5049 472 5095 529
rect 5049 369 5095 426
rect 5049 266 5095 323
rect 5049 163 5095 220
rect 5049 59 5095 117
rect 5049 0 5095 13
rect 5293 987 5339 1000
rect 5293 884 5339 941
rect 5293 781 5339 838
rect 5293 678 5339 735
rect 5293 575 5339 632
rect 5293 472 5339 529
rect 5293 369 5339 426
rect 5293 266 5339 323
rect 5293 163 5339 220
rect 5293 59 5339 117
rect 5293 0 5339 13
rect 5537 987 5583 1000
rect 5537 884 5583 941
rect 5537 781 5583 838
rect 5537 678 5583 735
rect 5537 575 5583 632
rect 5537 472 5583 529
rect 5537 369 5583 426
rect 5537 266 5583 323
rect 5537 163 5583 220
rect 5537 59 5583 117
rect 5537 0 5583 13
rect 5781 987 5827 1000
rect 5781 884 5827 941
rect 5781 781 5827 838
rect 5781 678 5827 735
rect 5781 575 5827 632
rect 5781 472 5827 529
rect 5781 369 5827 426
rect 5781 266 5827 323
rect 5781 163 5827 220
rect 5781 59 5827 117
rect 5781 0 5827 13
<< labels >>
rlabel metal1 5560 500 5560 500 4 D
rlabel metal1 5316 500 5316 500 4 S
rlabel metal1 5072 500 5072 500 4 D
rlabel metal1 4828 500 4828 500 4 S
rlabel metal1 4584 500 4584 500 4 D
rlabel metal1 4340 500 4340 500 4 S
rlabel metal1 4096 500 4096 500 4 D
rlabel metal1 3852 500 3852 500 4 S
rlabel metal1 3608 500 3608 500 4 D
rlabel metal1 3364 500 3364 500 4 S
rlabel metal1 3120 500 3120 500 4 D
rlabel metal1 2876 500 2876 500 4 S
rlabel metal1 2632 500 2632 500 4 D
rlabel metal1 2388 500 2388 500 4 S
rlabel metal1 2144 500 2144 500 4 D
rlabel metal1 1900 500 1900 500 4 S
rlabel metal1 1656 500 1656 500 4 D
rlabel metal1 1412 500 1412 500 4 S
rlabel metal1 1168 500 1168 500 4 D
rlabel metal1 924 500 924 500 4 S
rlabel metal1 680 500 680 500 4 D
rlabel metal1 436 500 436 500 4 S
rlabel metal1 192 500 192 500 4 D
rlabel metal1 5804 500 5804 500 4 S
rlabel metal1 -52 500 -52 500 4 S
<< end >>
