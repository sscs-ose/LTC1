magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1646 -1151 1646 1151
<< metal1 >>
rect -646 145 646 151
rect -646 119 -640 145
rect -614 119 -574 145
rect -548 119 -508 145
rect -482 119 -442 145
rect -416 119 -376 145
rect -350 119 -310 145
rect -284 119 -244 145
rect -218 119 -178 145
rect -152 119 -112 145
rect -86 119 -46 145
rect -20 119 20 145
rect 46 119 86 145
rect 112 119 152 145
rect 178 119 218 145
rect 244 119 284 145
rect 310 119 350 145
rect 376 119 416 145
rect 442 119 482 145
rect 508 119 548 145
rect 574 119 614 145
rect 640 119 646 145
rect -646 79 646 119
rect -646 53 -640 79
rect -614 53 -574 79
rect -548 53 -508 79
rect -482 53 -442 79
rect -416 53 -376 79
rect -350 53 -310 79
rect -284 53 -244 79
rect -218 53 -178 79
rect -152 53 -112 79
rect -86 53 -46 79
rect -20 53 20 79
rect 46 53 86 79
rect 112 53 152 79
rect 178 53 218 79
rect 244 53 284 79
rect 310 53 350 79
rect 376 53 416 79
rect 442 53 482 79
rect 508 53 548 79
rect 574 53 614 79
rect 640 53 646 79
rect -646 13 646 53
rect -646 -13 -640 13
rect -614 -13 -574 13
rect -548 -13 -508 13
rect -482 -13 -442 13
rect -416 -13 -376 13
rect -350 -13 -310 13
rect -284 -13 -244 13
rect -218 -13 -178 13
rect -152 -13 -112 13
rect -86 -13 -46 13
rect -20 -13 20 13
rect 46 -13 86 13
rect 112 -13 152 13
rect 178 -13 218 13
rect 244 -13 284 13
rect 310 -13 350 13
rect 376 -13 416 13
rect 442 -13 482 13
rect 508 -13 548 13
rect 574 -13 614 13
rect 640 -13 646 13
rect -646 -53 646 -13
rect -646 -79 -640 -53
rect -614 -79 -574 -53
rect -548 -79 -508 -53
rect -482 -79 -442 -53
rect -416 -79 -376 -53
rect -350 -79 -310 -53
rect -284 -79 -244 -53
rect -218 -79 -178 -53
rect -152 -79 -112 -53
rect -86 -79 -46 -53
rect -20 -79 20 -53
rect 46 -79 86 -53
rect 112 -79 152 -53
rect 178 -79 218 -53
rect 244 -79 284 -53
rect 310 -79 350 -53
rect 376 -79 416 -53
rect 442 -79 482 -53
rect 508 -79 548 -53
rect 574 -79 614 -53
rect 640 -79 646 -53
rect -646 -119 646 -79
rect -646 -145 -640 -119
rect -614 -145 -574 -119
rect -548 -145 -508 -119
rect -482 -145 -442 -119
rect -416 -145 -376 -119
rect -350 -145 -310 -119
rect -284 -145 -244 -119
rect -218 -145 -178 -119
rect -152 -145 -112 -119
rect -86 -145 -46 -119
rect -20 -145 20 -119
rect 46 -145 86 -119
rect 112 -145 152 -119
rect 178 -145 218 -119
rect 244 -145 284 -119
rect 310 -145 350 -119
rect 376 -145 416 -119
rect 442 -145 482 -119
rect 508 -145 548 -119
rect 574 -145 614 -119
rect 640 -145 646 -119
rect -646 -151 646 -145
<< via1 >>
rect -640 119 -614 145
rect -574 119 -548 145
rect -508 119 -482 145
rect -442 119 -416 145
rect -376 119 -350 145
rect -310 119 -284 145
rect -244 119 -218 145
rect -178 119 -152 145
rect -112 119 -86 145
rect -46 119 -20 145
rect 20 119 46 145
rect 86 119 112 145
rect 152 119 178 145
rect 218 119 244 145
rect 284 119 310 145
rect 350 119 376 145
rect 416 119 442 145
rect 482 119 508 145
rect 548 119 574 145
rect 614 119 640 145
rect -640 53 -614 79
rect -574 53 -548 79
rect -508 53 -482 79
rect -442 53 -416 79
rect -376 53 -350 79
rect -310 53 -284 79
rect -244 53 -218 79
rect -178 53 -152 79
rect -112 53 -86 79
rect -46 53 -20 79
rect 20 53 46 79
rect 86 53 112 79
rect 152 53 178 79
rect 218 53 244 79
rect 284 53 310 79
rect 350 53 376 79
rect 416 53 442 79
rect 482 53 508 79
rect 548 53 574 79
rect 614 53 640 79
rect -640 -13 -614 13
rect -574 -13 -548 13
rect -508 -13 -482 13
rect -442 -13 -416 13
rect -376 -13 -350 13
rect -310 -13 -284 13
rect -244 -13 -218 13
rect -178 -13 -152 13
rect -112 -13 -86 13
rect -46 -13 -20 13
rect 20 -13 46 13
rect 86 -13 112 13
rect 152 -13 178 13
rect 218 -13 244 13
rect 284 -13 310 13
rect 350 -13 376 13
rect 416 -13 442 13
rect 482 -13 508 13
rect 548 -13 574 13
rect 614 -13 640 13
rect -640 -79 -614 -53
rect -574 -79 -548 -53
rect -508 -79 -482 -53
rect -442 -79 -416 -53
rect -376 -79 -350 -53
rect -310 -79 -284 -53
rect -244 -79 -218 -53
rect -178 -79 -152 -53
rect -112 -79 -86 -53
rect -46 -79 -20 -53
rect 20 -79 46 -53
rect 86 -79 112 -53
rect 152 -79 178 -53
rect 218 -79 244 -53
rect 284 -79 310 -53
rect 350 -79 376 -53
rect 416 -79 442 -53
rect 482 -79 508 -53
rect 548 -79 574 -53
rect 614 -79 640 -53
rect -640 -145 -614 -119
rect -574 -145 -548 -119
rect -508 -145 -482 -119
rect -442 -145 -416 -119
rect -376 -145 -350 -119
rect -310 -145 -284 -119
rect -244 -145 -218 -119
rect -178 -145 -152 -119
rect -112 -145 -86 -119
rect -46 -145 -20 -119
rect 20 -145 46 -119
rect 86 -145 112 -119
rect 152 -145 178 -119
rect 218 -145 244 -119
rect 284 -145 310 -119
rect 350 -145 376 -119
rect 416 -145 442 -119
rect 482 -145 508 -119
rect 548 -145 574 -119
rect 614 -145 640 -119
<< metal2 >>
rect -646 145 646 151
rect -646 119 -640 145
rect -614 119 -574 145
rect -548 119 -508 145
rect -482 119 -442 145
rect -416 119 -376 145
rect -350 119 -310 145
rect -284 119 -244 145
rect -218 119 -178 145
rect -152 119 -112 145
rect -86 119 -46 145
rect -20 119 20 145
rect 46 119 86 145
rect 112 119 152 145
rect 178 119 218 145
rect 244 119 284 145
rect 310 119 350 145
rect 376 119 416 145
rect 442 119 482 145
rect 508 119 548 145
rect 574 119 614 145
rect 640 119 646 145
rect -646 79 646 119
rect -646 53 -640 79
rect -614 53 -574 79
rect -548 53 -508 79
rect -482 53 -442 79
rect -416 53 -376 79
rect -350 53 -310 79
rect -284 53 -244 79
rect -218 53 -178 79
rect -152 53 -112 79
rect -86 53 -46 79
rect -20 53 20 79
rect 46 53 86 79
rect 112 53 152 79
rect 178 53 218 79
rect 244 53 284 79
rect 310 53 350 79
rect 376 53 416 79
rect 442 53 482 79
rect 508 53 548 79
rect 574 53 614 79
rect 640 53 646 79
rect -646 13 646 53
rect -646 -13 -640 13
rect -614 -13 -574 13
rect -548 -13 -508 13
rect -482 -13 -442 13
rect -416 -13 -376 13
rect -350 -13 -310 13
rect -284 -13 -244 13
rect -218 -13 -178 13
rect -152 -13 -112 13
rect -86 -13 -46 13
rect -20 -13 20 13
rect 46 -13 86 13
rect 112 -13 152 13
rect 178 -13 218 13
rect 244 -13 284 13
rect 310 -13 350 13
rect 376 -13 416 13
rect 442 -13 482 13
rect 508 -13 548 13
rect 574 -13 614 13
rect 640 -13 646 13
rect -646 -53 646 -13
rect -646 -79 -640 -53
rect -614 -79 -574 -53
rect -548 -79 -508 -53
rect -482 -79 -442 -53
rect -416 -79 -376 -53
rect -350 -79 -310 -53
rect -284 -79 -244 -53
rect -218 -79 -178 -53
rect -152 -79 -112 -53
rect -86 -79 -46 -53
rect -20 -79 20 -53
rect 46 -79 86 -53
rect 112 -79 152 -53
rect 178 -79 218 -53
rect 244 -79 284 -53
rect 310 -79 350 -53
rect 376 -79 416 -53
rect 442 -79 482 -53
rect 508 -79 548 -53
rect 574 -79 614 -53
rect 640 -79 646 -53
rect -646 -119 646 -79
rect -646 -145 -640 -119
rect -614 -145 -574 -119
rect -548 -145 -508 -119
rect -482 -145 -442 -119
rect -416 -145 -376 -119
rect -350 -145 -310 -119
rect -284 -145 -244 -119
rect -218 -145 -178 -119
rect -152 -145 -112 -119
rect -86 -145 -46 -119
rect -20 -145 20 -119
rect 46 -145 86 -119
rect 112 -145 152 -119
rect 178 -145 218 -119
rect 244 -145 284 -119
rect 310 -145 350 -119
rect 376 -145 416 -119
rect 442 -145 482 -119
rect 508 -145 548 -119
rect 574 -145 614 -119
rect 640 -145 646 -119
rect -646 -151 646 -145
<< end >>
