magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 6864 12044
<< mvnmos >>
rect 0 0 140 10000
rect 244 0 384 10000
rect 488 0 628 10000
rect 732 0 872 10000
rect 976 0 1116 10000
rect 1220 0 1360 10000
rect 1464 0 1604 10000
rect 1708 0 1848 10000
rect 1952 0 2092 10000
rect 2196 0 2336 10000
rect 2440 0 2580 10000
rect 2684 0 2824 10000
rect 2928 0 3068 10000
rect 3172 0 3312 10000
rect 3416 0 3556 10000
rect 3660 0 3800 10000
rect 3904 0 4044 10000
rect 4148 0 4288 10000
rect 4392 0 4532 10000
rect 4636 0 4776 10000
<< mvndiff >>
rect -88 9958 0 10000
rect -88 42 -75 9958
rect -29 42 0 9958
rect -88 0 0 42
rect 140 9958 244 10000
rect 140 42 169 9958
rect 215 42 244 9958
rect 140 0 244 42
rect 384 9958 488 10000
rect 384 42 413 9958
rect 459 42 488 9958
rect 384 0 488 42
rect 628 9958 732 10000
rect 628 42 657 9958
rect 703 42 732 9958
rect 628 0 732 42
rect 872 9958 976 10000
rect 872 42 901 9958
rect 947 42 976 9958
rect 872 0 976 42
rect 1116 9958 1220 10000
rect 1116 42 1145 9958
rect 1191 42 1220 9958
rect 1116 0 1220 42
rect 1360 9958 1464 10000
rect 1360 42 1389 9958
rect 1435 42 1464 9958
rect 1360 0 1464 42
rect 1604 9958 1708 10000
rect 1604 42 1633 9958
rect 1679 42 1708 9958
rect 1604 0 1708 42
rect 1848 9958 1952 10000
rect 1848 42 1877 9958
rect 1923 42 1952 9958
rect 1848 0 1952 42
rect 2092 9958 2196 10000
rect 2092 42 2121 9958
rect 2167 42 2196 9958
rect 2092 0 2196 42
rect 2336 9958 2440 10000
rect 2336 42 2365 9958
rect 2411 42 2440 9958
rect 2336 0 2440 42
rect 2580 9958 2684 10000
rect 2580 42 2609 9958
rect 2655 42 2684 9958
rect 2580 0 2684 42
rect 2824 9958 2928 10000
rect 2824 42 2853 9958
rect 2899 42 2928 9958
rect 2824 0 2928 42
rect 3068 9958 3172 10000
rect 3068 42 3097 9958
rect 3143 42 3172 9958
rect 3068 0 3172 42
rect 3312 9958 3416 10000
rect 3312 42 3341 9958
rect 3387 42 3416 9958
rect 3312 0 3416 42
rect 3556 9958 3660 10000
rect 3556 42 3585 9958
rect 3631 42 3660 9958
rect 3556 0 3660 42
rect 3800 9958 3904 10000
rect 3800 42 3829 9958
rect 3875 42 3904 9958
rect 3800 0 3904 42
rect 4044 9958 4148 10000
rect 4044 42 4073 9958
rect 4119 42 4148 9958
rect 4044 0 4148 42
rect 4288 9958 4392 10000
rect 4288 42 4317 9958
rect 4363 42 4392 9958
rect 4288 0 4392 42
rect 4532 9958 4636 10000
rect 4532 42 4561 9958
rect 4607 42 4636 9958
rect 4532 0 4636 42
rect 4776 9958 4864 10000
rect 4776 42 4805 9958
rect 4851 42 4864 9958
rect 4776 0 4864 42
<< mvndiffc >>
rect -75 42 -29 9958
rect 169 42 215 9958
rect 413 42 459 9958
rect 657 42 703 9958
rect 901 42 947 9958
rect 1145 42 1191 9958
rect 1389 42 1435 9958
rect 1633 42 1679 9958
rect 1877 42 1923 9958
rect 2121 42 2167 9958
rect 2365 42 2411 9958
rect 2609 42 2655 9958
rect 2853 42 2899 9958
rect 3097 42 3143 9958
rect 3341 42 3387 9958
rect 3585 42 3631 9958
rect 3829 42 3875 9958
rect 4073 42 4119 9958
rect 4317 42 4363 9958
rect 4561 42 4607 9958
rect 4805 42 4851 9958
<< polysilicon >>
rect 0 10000 140 10044
rect 244 10000 384 10044
rect 488 10000 628 10044
rect 732 10000 872 10044
rect 976 10000 1116 10044
rect 1220 10000 1360 10044
rect 1464 10000 1604 10044
rect 1708 10000 1848 10044
rect 1952 10000 2092 10044
rect 2196 10000 2336 10044
rect 2440 10000 2580 10044
rect 2684 10000 2824 10044
rect 2928 10000 3068 10044
rect 3172 10000 3312 10044
rect 3416 10000 3556 10044
rect 3660 10000 3800 10044
rect 3904 10000 4044 10044
rect 4148 10000 4288 10044
rect 4392 10000 4532 10044
rect 4636 10000 4776 10044
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
rect 976 -44 1116 0
rect 1220 -44 1360 0
rect 1464 -44 1604 0
rect 1708 -44 1848 0
rect 1952 -44 2092 0
rect 2196 -44 2336 0
rect 2440 -44 2580 0
rect 2684 -44 2824 0
rect 2928 -44 3068 0
rect 3172 -44 3312 0
rect 3416 -44 3556 0
rect 3660 -44 3800 0
rect 3904 -44 4044 0
rect 4148 -44 4288 0
rect 4392 -44 4532 0
rect 4636 -44 4776 0
<< metal1 >>
rect -75 9958 -29 10000
rect -75 0 -29 42
rect 169 9958 215 10000
rect 169 0 215 42
rect 413 9958 459 10000
rect 413 0 459 42
rect 657 9958 703 10000
rect 657 0 703 42
rect 901 9958 947 10000
rect 901 0 947 42
rect 1145 9958 1191 10000
rect 1145 0 1191 42
rect 1389 9958 1435 10000
rect 1389 0 1435 42
rect 1633 9958 1679 10000
rect 1633 0 1679 42
rect 1877 9958 1923 10000
rect 1877 0 1923 42
rect 2121 9958 2167 10000
rect 2121 0 2167 42
rect 2365 9958 2411 10000
rect 2365 0 2411 42
rect 2609 9958 2655 10000
rect 2609 0 2655 42
rect 2853 9958 2899 10000
rect 2853 0 2899 42
rect 3097 9958 3143 10000
rect 3097 0 3143 42
rect 3341 9958 3387 10000
rect 3341 0 3387 42
rect 3585 9958 3631 10000
rect 3585 0 3631 42
rect 3829 9958 3875 10000
rect 3829 0 3875 42
rect 4073 9958 4119 10000
rect 4073 0 4119 42
rect 4317 9958 4363 10000
rect 4317 0 4363 42
rect 4561 9958 4607 10000
rect 4561 0 4607 42
rect 4805 9958 4851 10000
rect 4805 0 4851 42
<< labels >>
rlabel mvndiffc 4584 5000 4584 5000 4 D
rlabel mvndiffc 4340 5000 4340 5000 4 S
rlabel mvndiffc 4096 5000 4096 5000 4 D
rlabel mvndiffc 3852 5000 3852 5000 4 S
rlabel mvndiffc 3608 5000 3608 5000 4 D
rlabel mvndiffc 3364 5000 3364 5000 4 S
rlabel mvndiffc 3120 5000 3120 5000 4 D
rlabel mvndiffc 2876 5000 2876 5000 4 S
rlabel mvndiffc 2632 5000 2632 5000 4 D
rlabel mvndiffc 2388 5000 2388 5000 4 S
rlabel mvndiffc 2144 5000 2144 5000 4 D
rlabel mvndiffc 1900 5000 1900 5000 4 S
rlabel mvndiffc 1656 5000 1656 5000 4 D
rlabel mvndiffc 1412 5000 1412 5000 4 S
rlabel mvndiffc 1168 5000 1168 5000 4 D
rlabel mvndiffc 924 5000 924 5000 4 S
rlabel mvndiffc 680 5000 680 5000 4 D
rlabel mvndiffc 436 5000 436 5000 4 S
rlabel mvndiffc 192 5000 192 5000 4 D
rlabel mvndiffc 4828 5000 4828 5000 4 S
rlabel mvndiffc -52 5000 -52 5000 4 S
<< end >>
