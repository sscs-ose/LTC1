magic
tech gf180mcuC
magscale 1 10
timestamp 1694921777
<< nwell >>
rect -1242 -1534 1242 1534
<< pmos >>
rect -1068 804 -1012 1404
rect -908 804 -852 1404
rect -748 804 -692 1404
rect -588 804 -532 1404
rect -428 804 -372 1404
rect -268 804 -212 1404
rect -108 804 -52 1404
rect 52 804 108 1404
rect 212 804 268 1404
rect 372 804 428 1404
rect 532 804 588 1404
rect 692 804 748 1404
rect 852 804 908 1404
rect 1012 804 1068 1404
rect -1068 68 -1012 668
rect -908 68 -852 668
rect -748 68 -692 668
rect -588 68 -532 668
rect -428 68 -372 668
rect -268 68 -212 668
rect -108 68 -52 668
rect 52 68 108 668
rect 212 68 268 668
rect 372 68 428 668
rect 532 68 588 668
rect 692 68 748 668
rect 852 68 908 668
rect 1012 68 1068 668
rect -1068 -668 -1012 -68
rect -908 -668 -852 -68
rect -748 -668 -692 -68
rect -588 -668 -532 -68
rect -428 -668 -372 -68
rect -268 -668 -212 -68
rect -108 -668 -52 -68
rect 52 -668 108 -68
rect 212 -668 268 -68
rect 372 -668 428 -68
rect 532 -668 588 -68
rect 692 -668 748 -68
rect 852 -668 908 -68
rect 1012 -668 1068 -68
rect -1068 -1404 -1012 -804
rect -908 -1404 -852 -804
rect -748 -1404 -692 -804
rect -588 -1404 -532 -804
rect -428 -1404 -372 -804
rect -268 -1404 -212 -804
rect -108 -1404 -52 -804
rect 52 -1404 108 -804
rect 212 -1404 268 -804
rect 372 -1404 428 -804
rect 532 -1404 588 -804
rect 692 -1404 748 -804
rect 852 -1404 908 -804
rect 1012 -1404 1068 -804
<< pdiff >>
rect -1156 1391 -1068 1404
rect -1156 817 -1143 1391
rect -1097 817 -1068 1391
rect -1156 804 -1068 817
rect -1012 1391 -908 1404
rect -1012 817 -983 1391
rect -937 817 -908 1391
rect -1012 804 -908 817
rect -852 1391 -748 1404
rect -852 817 -823 1391
rect -777 817 -748 1391
rect -852 804 -748 817
rect -692 1391 -588 1404
rect -692 817 -663 1391
rect -617 817 -588 1391
rect -692 804 -588 817
rect -532 1391 -428 1404
rect -532 817 -503 1391
rect -457 817 -428 1391
rect -532 804 -428 817
rect -372 1391 -268 1404
rect -372 817 -343 1391
rect -297 817 -268 1391
rect -372 804 -268 817
rect -212 1391 -108 1404
rect -212 817 -183 1391
rect -137 817 -108 1391
rect -212 804 -108 817
rect -52 1391 52 1404
rect -52 817 -23 1391
rect 23 817 52 1391
rect -52 804 52 817
rect 108 1391 212 1404
rect 108 817 137 1391
rect 183 817 212 1391
rect 108 804 212 817
rect 268 1391 372 1404
rect 268 817 297 1391
rect 343 817 372 1391
rect 268 804 372 817
rect 428 1391 532 1404
rect 428 817 457 1391
rect 503 817 532 1391
rect 428 804 532 817
rect 588 1391 692 1404
rect 588 817 617 1391
rect 663 817 692 1391
rect 588 804 692 817
rect 748 1391 852 1404
rect 748 817 777 1391
rect 823 817 852 1391
rect 748 804 852 817
rect 908 1391 1012 1404
rect 908 817 937 1391
rect 983 817 1012 1391
rect 908 804 1012 817
rect 1068 1391 1156 1404
rect 1068 817 1097 1391
rect 1143 817 1156 1391
rect 1068 804 1156 817
rect -1156 655 -1068 668
rect -1156 81 -1143 655
rect -1097 81 -1068 655
rect -1156 68 -1068 81
rect -1012 655 -908 668
rect -1012 81 -983 655
rect -937 81 -908 655
rect -1012 68 -908 81
rect -852 655 -748 668
rect -852 81 -823 655
rect -777 81 -748 655
rect -852 68 -748 81
rect -692 655 -588 668
rect -692 81 -663 655
rect -617 81 -588 655
rect -692 68 -588 81
rect -532 655 -428 668
rect -532 81 -503 655
rect -457 81 -428 655
rect -532 68 -428 81
rect -372 655 -268 668
rect -372 81 -343 655
rect -297 81 -268 655
rect -372 68 -268 81
rect -212 655 -108 668
rect -212 81 -183 655
rect -137 81 -108 655
rect -212 68 -108 81
rect -52 655 52 668
rect -52 81 -23 655
rect 23 81 52 655
rect -52 68 52 81
rect 108 655 212 668
rect 108 81 137 655
rect 183 81 212 655
rect 108 68 212 81
rect 268 655 372 668
rect 268 81 297 655
rect 343 81 372 655
rect 268 68 372 81
rect 428 655 532 668
rect 428 81 457 655
rect 503 81 532 655
rect 428 68 532 81
rect 588 655 692 668
rect 588 81 617 655
rect 663 81 692 655
rect 588 68 692 81
rect 748 655 852 668
rect 748 81 777 655
rect 823 81 852 655
rect 748 68 852 81
rect 908 655 1012 668
rect 908 81 937 655
rect 983 81 1012 655
rect 908 68 1012 81
rect 1068 655 1156 668
rect 1068 81 1097 655
rect 1143 81 1156 655
rect 1068 68 1156 81
rect -1156 -81 -1068 -68
rect -1156 -655 -1143 -81
rect -1097 -655 -1068 -81
rect -1156 -668 -1068 -655
rect -1012 -81 -908 -68
rect -1012 -655 -983 -81
rect -937 -655 -908 -81
rect -1012 -668 -908 -655
rect -852 -81 -748 -68
rect -852 -655 -823 -81
rect -777 -655 -748 -81
rect -852 -668 -748 -655
rect -692 -81 -588 -68
rect -692 -655 -663 -81
rect -617 -655 -588 -81
rect -692 -668 -588 -655
rect -532 -81 -428 -68
rect -532 -655 -503 -81
rect -457 -655 -428 -81
rect -532 -668 -428 -655
rect -372 -81 -268 -68
rect -372 -655 -343 -81
rect -297 -655 -268 -81
rect -372 -668 -268 -655
rect -212 -81 -108 -68
rect -212 -655 -183 -81
rect -137 -655 -108 -81
rect -212 -668 -108 -655
rect -52 -81 52 -68
rect -52 -655 -23 -81
rect 23 -655 52 -81
rect -52 -668 52 -655
rect 108 -81 212 -68
rect 108 -655 137 -81
rect 183 -655 212 -81
rect 108 -668 212 -655
rect 268 -81 372 -68
rect 268 -655 297 -81
rect 343 -655 372 -81
rect 268 -668 372 -655
rect 428 -81 532 -68
rect 428 -655 457 -81
rect 503 -655 532 -81
rect 428 -668 532 -655
rect 588 -81 692 -68
rect 588 -655 617 -81
rect 663 -655 692 -81
rect 588 -668 692 -655
rect 748 -81 852 -68
rect 748 -655 777 -81
rect 823 -655 852 -81
rect 748 -668 852 -655
rect 908 -81 1012 -68
rect 908 -655 937 -81
rect 983 -655 1012 -81
rect 908 -668 1012 -655
rect 1068 -81 1156 -68
rect 1068 -655 1097 -81
rect 1143 -655 1156 -81
rect 1068 -668 1156 -655
rect -1156 -817 -1068 -804
rect -1156 -1391 -1143 -817
rect -1097 -1391 -1068 -817
rect -1156 -1404 -1068 -1391
rect -1012 -817 -908 -804
rect -1012 -1391 -983 -817
rect -937 -1391 -908 -817
rect -1012 -1404 -908 -1391
rect -852 -817 -748 -804
rect -852 -1391 -823 -817
rect -777 -1391 -748 -817
rect -852 -1404 -748 -1391
rect -692 -817 -588 -804
rect -692 -1391 -663 -817
rect -617 -1391 -588 -817
rect -692 -1404 -588 -1391
rect -532 -817 -428 -804
rect -532 -1391 -503 -817
rect -457 -1391 -428 -817
rect -532 -1404 -428 -1391
rect -372 -817 -268 -804
rect -372 -1391 -343 -817
rect -297 -1391 -268 -817
rect -372 -1404 -268 -1391
rect -212 -817 -108 -804
rect -212 -1391 -183 -817
rect -137 -1391 -108 -817
rect -212 -1404 -108 -1391
rect -52 -817 52 -804
rect -52 -1391 -23 -817
rect 23 -1391 52 -817
rect -52 -1404 52 -1391
rect 108 -817 212 -804
rect 108 -1391 137 -817
rect 183 -1391 212 -817
rect 108 -1404 212 -1391
rect 268 -817 372 -804
rect 268 -1391 297 -817
rect 343 -1391 372 -817
rect 268 -1404 372 -1391
rect 428 -817 532 -804
rect 428 -1391 457 -817
rect 503 -1391 532 -817
rect 428 -1404 532 -1391
rect 588 -817 692 -804
rect 588 -1391 617 -817
rect 663 -1391 692 -817
rect 588 -1404 692 -1391
rect 748 -817 852 -804
rect 748 -1391 777 -817
rect 823 -1391 852 -817
rect 748 -1404 852 -1391
rect 908 -817 1012 -804
rect 908 -1391 937 -817
rect 983 -1391 1012 -817
rect 908 -1404 1012 -1391
rect 1068 -817 1156 -804
rect 1068 -1391 1097 -817
rect 1143 -1391 1156 -817
rect 1068 -1404 1156 -1391
<< pdiffc >>
rect -1143 817 -1097 1391
rect -983 817 -937 1391
rect -823 817 -777 1391
rect -663 817 -617 1391
rect -503 817 -457 1391
rect -343 817 -297 1391
rect -183 817 -137 1391
rect -23 817 23 1391
rect 137 817 183 1391
rect 297 817 343 1391
rect 457 817 503 1391
rect 617 817 663 1391
rect 777 817 823 1391
rect 937 817 983 1391
rect 1097 817 1143 1391
rect -1143 81 -1097 655
rect -983 81 -937 655
rect -823 81 -777 655
rect -663 81 -617 655
rect -503 81 -457 655
rect -343 81 -297 655
rect -183 81 -137 655
rect -23 81 23 655
rect 137 81 183 655
rect 297 81 343 655
rect 457 81 503 655
rect 617 81 663 655
rect 777 81 823 655
rect 937 81 983 655
rect 1097 81 1143 655
rect -1143 -655 -1097 -81
rect -983 -655 -937 -81
rect -823 -655 -777 -81
rect -663 -655 -617 -81
rect -503 -655 -457 -81
rect -343 -655 -297 -81
rect -183 -655 -137 -81
rect -23 -655 23 -81
rect 137 -655 183 -81
rect 297 -655 343 -81
rect 457 -655 503 -81
rect 617 -655 663 -81
rect 777 -655 823 -81
rect 937 -655 983 -81
rect 1097 -655 1143 -81
rect -1143 -1391 -1097 -817
rect -983 -1391 -937 -817
rect -823 -1391 -777 -817
rect -663 -1391 -617 -817
rect -503 -1391 -457 -817
rect -343 -1391 -297 -817
rect -183 -1391 -137 -817
rect -23 -1391 23 -817
rect 137 -1391 183 -817
rect 297 -1391 343 -817
rect 457 -1391 503 -817
rect 617 -1391 663 -817
rect 777 -1391 823 -817
rect 937 -1391 983 -817
rect 1097 -1391 1143 -817
<< polysilicon >>
rect -1068 1404 -1012 1448
rect -908 1404 -852 1448
rect -748 1404 -692 1448
rect -588 1404 -532 1448
rect -428 1404 -372 1448
rect -268 1404 -212 1448
rect -108 1404 -52 1448
rect 52 1404 108 1448
rect 212 1404 268 1448
rect 372 1404 428 1448
rect 532 1404 588 1448
rect 692 1404 748 1448
rect 852 1404 908 1448
rect 1012 1404 1068 1448
rect -1068 760 -1012 804
rect -908 760 -852 804
rect -748 760 -692 804
rect -588 760 -532 804
rect -428 760 -372 804
rect -268 760 -212 804
rect -108 760 -52 804
rect 52 760 108 804
rect 212 760 268 804
rect 372 760 428 804
rect 532 760 588 804
rect 692 760 748 804
rect 852 760 908 804
rect 1012 760 1068 804
rect -1068 668 -1012 712
rect -908 668 -852 712
rect -748 668 -692 712
rect -588 668 -532 712
rect -428 668 -372 712
rect -268 668 -212 712
rect -108 668 -52 712
rect 52 668 108 712
rect 212 668 268 712
rect 372 668 428 712
rect 532 668 588 712
rect 692 668 748 712
rect 852 668 908 712
rect 1012 668 1068 712
rect -1068 24 -1012 68
rect -908 24 -852 68
rect -748 24 -692 68
rect -588 24 -532 68
rect -428 24 -372 68
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect 372 24 428 68
rect 532 24 588 68
rect 692 24 748 68
rect 852 24 908 68
rect 1012 24 1068 68
rect -1068 -68 -1012 -24
rect -908 -68 -852 -24
rect -748 -68 -692 -24
rect -588 -68 -532 -24
rect -428 -68 -372 -24
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect 372 -68 428 -24
rect 532 -68 588 -24
rect 692 -68 748 -24
rect 852 -68 908 -24
rect 1012 -68 1068 -24
rect -1068 -712 -1012 -668
rect -908 -712 -852 -668
rect -748 -712 -692 -668
rect -588 -712 -532 -668
rect -428 -712 -372 -668
rect -268 -712 -212 -668
rect -108 -712 -52 -668
rect 52 -712 108 -668
rect 212 -712 268 -668
rect 372 -712 428 -668
rect 532 -712 588 -668
rect 692 -712 748 -668
rect 852 -712 908 -668
rect 1012 -712 1068 -668
rect -1068 -804 -1012 -760
rect -908 -804 -852 -760
rect -748 -804 -692 -760
rect -588 -804 -532 -760
rect -428 -804 -372 -760
rect -268 -804 -212 -760
rect -108 -804 -52 -760
rect 52 -804 108 -760
rect 212 -804 268 -760
rect 372 -804 428 -760
rect 532 -804 588 -760
rect 692 -804 748 -760
rect 852 -804 908 -760
rect 1012 -804 1068 -760
rect -1068 -1448 -1012 -1404
rect -908 -1448 -852 -1404
rect -748 -1448 -692 -1404
rect -588 -1448 -532 -1404
rect -428 -1448 -372 -1404
rect -268 -1448 -212 -1404
rect -108 -1448 -52 -1404
rect 52 -1448 108 -1404
rect 212 -1448 268 -1404
rect 372 -1448 428 -1404
rect 532 -1448 588 -1404
rect 692 -1448 748 -1404
rect 852 -1448 908 -1404
rect 1012 -1448 1068 -1404
<< metal1 >>
rect -1143 1391 -1097 1402
rect -1143 806 -1097 817
rect -983 1391 -937 1402
rect -983 806 -937 817
rect -823 1391 -777 1402
rect -823 806 -777 817
rect -663 1391 -617 1402
rect -663 806 -617 817
rect -503 1391 -457 1402
rect -503 806 -457 817
rect -343 1391 -297 1402
rect -343 806 -297 817
rect -183 1391 -137 1402
rect -183 806 -137 817
rect -23 1391 23 1402
rect -23 806 23 817
rect 137 1391 183 1402
rect 137 806 183 817
rect 297 1391 343 1402
rect 297 806 343 817
rect 457 1391 503 1402
rect 457 806 503 817
rect 617 1391 663 1402
rect 617 806 663 817
rect 777 1391 823 1402
rect 777 806 823 817
rect 937 1391 983 1402
rect 937 806 983 817
rect 1097 1391 1143 1402
rect 1097 806 1143 817
rect -1143 655 -1097 666
rect -1143 70 -1097 81
rect -983 655 -937 666
rect -983 70 -937 81
rect -823 655 -777 666
rect -823 70 -777 81
rect -663 655 -617 666
rect -663 70 -617 81
rect -503 655 -457 666
rect -503 70 -457 81
rect -343 655 -297 666
rect -343 70 -297 81
rect -183 655 -137 666
rect -183 70 -137 81
rect -23 655 23 666
rect -23 70 23 81
rect 137 655 183 666
rect 137 70 183 81
rect 297 655 343 666
rect 297 70 343 81
rect 457 655 503 666
rect 457 70 503 81
rect 617 655 663 666
rect 617 70 663 81
rect 777 655 823 666
rect 777 70 823 81
rect 937 655 983 666
rect 937 70 983 81
rect 1097 655 1143 666
rect 1097 70 1143 81
rect -1143 -81 -1097 -70
rect -1143 -666 -1097 -655
rect -983 -81 -937 -70
rect -983 -666 -937 -655
rect -823 -81 -777 -70
rect -823 -666 -777 -655
rect -663 -81 -617 -70
rect -663 -666 -617 -655
rect -503 -81 -457 -70
rect -503 -666 -457 -655
rect -343 -81 -297 -70
rect -343 -666 -297 -655
rect -183 -81 -137 -70
rect -183 -666 -137 -655
rect -23 -81 23 -70
rect -23 -666 23 -655
rect 137 -81 183 -70
rect 137 -666 183 -655
rect 297 -81 343 -70
rect 297 -666 343 -655
rect 457 -81 503 -70
rect 457 -666 503 -655
rect 617 -81 663 -70
rect 617 -666 663 -655
rect 777 -81 823 -70
rect 777 -666 823 -655
rect 937 -81 983 -70
rect 937 -666 983 -655
rect 1097 -81 1143 -70
rect 1097 -666 1143 -655
rect -1143 -817 -1097 -806
rect -1143 -1402 -1097 -1391
rect -983 -817 -937 -806
rect -983 -1402 -937 -1391
rect -823 -817 -777 -806
rect -823 -1402 -777 -1391
rect -663 -817 -617 -806
rect -663 -1402 -617 -1391
rect -503 -817 -457 -806
rect -503 -1402 -457 -1391
rect -343 -817 -297 -806
rect -343 -1402 -297 -1391
rect -183 -817 -137 -806
rect -183 -1402 -137 -1391
rect -23 -817 23 -806
rect -23 -1402 23 -1391
rect 137 -817 183 -806
rect 137 -1402 183 -1391
rect 297 -817 343 -806
rect 297 -1402 343 -1391
rect 457 -817 503 -806
rect 457 -1402 503 -1391
rect 617 -817 663 -806
rect 617 -1402 663 -1391
rect 777 -817 823 -806
rect 777 -1402 823 -1391
rect 937 -817 983 -806
rect 937 -1402 983 -1391
rect 1097 -817 1143 -806
rect 1097 -1402 1143 -1391
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 4 nf 14 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
