magic
tech gf180mcuC
magscale 1 10
timestamp 1695119997
<< nwell >>
rect 4706 3910 4860 4149
rect 5178 3910 5332 4149
rect 5503 3910 5657 4149
rect 5806 3910 5960 4149
<< pwell >>
rect 4449 1071 4562 1078
rect 4820 1070 4906 1073
rect 5244 1069 5330 1072
rect 6012 1069 6098 1072
rect 5630 1056 5716 1059
<< metal1 >>
rect -447 5362 6494 5567
rect -447 5270 4370 5362
rect -447 5171 -313 5270
rect -237 5263 4370 5270
rect -237 5171 -63 5263
rect -447 5164 -63 5171
rect 13 5224 4370 5263
rect 4475 5359 6494 5362
rect 4475 5224 4742 5359
rect 13 5221 4742 5224
rect 4847 5221 5214 5359
rect 5319 5221 5539 5359
rect 5644 5221 5842 5359
rect 5947 5221 6494 5359
rect 13 5164 6494 5221
rect -447 5140 6494 5164
rect 3236 4420 3351 4467
rect -70 3890 24 3974
rect -70 3837 -58 3890
rect 9 3837 24 3890
rect -70 3806 24 3837
rect 3789 3833 4253 4038
rect 4706 4101 4860 4149
rect 4706 3963 4742 4101
rect 4847 3963 4860 4101
rect 4706 3911 4860 3963
rect 5178 4101 5332 4149
rect 5178 3963 5214 4101
rect 5319 3963 5332 4101
rect 5178 3911 5332 3963
rect 5503 4101 5657 4149
rect 5503 3963 5539 4101
rect 5644 3963 5657 4101
rect 5503 3911 5657 3963
rect 5806 4101 5960 4149
rect 5806 3963 5842 4101
rect 5947 3963 5960 4101
rect 5806 3911 5960 3963
rect 4712 3910 4772 3911
rect 5184 3910 5244 3911
rect 5509 3910 5569 3911
rect 5812 3910 5872 3911
rect -69 3804 24 3806
rect -521 3392 -370 3442
rect -60 3392 166 3492
rect 4170 3428 4322 3442
rect 4170 3376 4191 3428
rect -73 3325 63 3340
rect -73 3272 -60 3325
rect 7 3272 63 3325
rect 3648 3301 3772 3349
rect 4095 3324 4191 3376
rect 4269 3356 4322 3428
rect 5899 3389 6558 3441
rect 4269 3324 4290 3356
rect 4095 3301 4290 3324
rect -73 3261 63 3272
rect 16 3119 63 3261
rect -472 3104 -373 3118
rect -472 3025 -457 3104
rect -386 3025 -373 3104
rect 16 3109 97 3119
rect 16 3048 28 3109
rect 86 3048 97 3109
rect 16 3036 97 3048
rect -472 3004 -373 3025
rect 3982 2796 4268 3135
rect 5921 2867 6577 3135
rect 204 2732 310 2754
rect 204 2722 214 2732
rect -472 2705 214 2722
rect -472 2644 -454 2705
rect -393 2644 214 2705
rect -472 2624 214 2644
rect 204 2617 214 2624
rect 294 2617 310 2732
rect 204 2603 310 2617
rect 3265 2729 3347 2731
rect 3265 2718 4100 2729
rect 3265 2666 4024 2718
rect 4082 2666 4100 2718
rect 3265 2654 4100 2666
rect 3265 2549 3347 2654
rect 3265 2542 4108 2549
rect 3265 2524 4033 2542
rect 3266 2490 4033 2524
rect 4091 2490 4108 2542
rect 3266 2473 4108 2490
rect 6362 2523 6519 2535
rect 204 2357 311 2363
rect -475 2343 311 2357
rect -475 2340 215 2343
rect -475 2240 -460 2340
rect -390 2240 215 2340
rect -475 2228 215 2240
rect 295 2228 311 2343
rect 3266 2317 3347 2473
rect 6362 2468 6431 2523
rect 6495 2468 6519 2523
rect 6362 2454 6519 2468
rect 5972 2370 6098 2427
rect 5972 2325 6043 2370
rect 3265 2308 4099 2317
rect 3265 2256 4022 2308
rect 4080 2256 4099 2308
rect 3265 2242 4099 2256
rect 5972 2251 5987 2325
rect 6039 2251 6043 2325
rect 5972 2237 6043 2251
rect -475 2220 311 2228
rect 204 2211 311 2220
rect 4170 2106 6569 2108
rect -472 1940 -373 1956
rect -472 1861 -458 1940
rect -387 1861 -373 1940
rect 4170 1943 6570 2106
rect 17 1914 97 1918
rect -472 1846 -373 1861
rect 17 1860 29 1914
rect 85 1860 97 1914
rect 17 1850 97 1860
rect 4170 1866 4198 1943
rect 4259 1866 6570 1943
rect 17 1786 64 1850
rect 4170 1836 6570 1866
rect -91 1773 64 1786
rect -91 1716 -73 1773
rect -9 1716 64 1773
rect -91 1700 64 1716
rect 3662 1617 3774 1665
rect 4087 1617 4356 1665
rect -555 1522 -419 1572
rect -73 1474 94 1572
rect 4308 1411 4356 1617
rect 4308 1401 4590 1411
rect 4308 1301 4443 1401
rect 4557 1301 4590 1401
rect 6029 1340 6587 1392
rect 4308 1288 4590 1301
rect -91 1211 5 1224
rect -91 1154 -76 1211
rect -12 1154 5 1211
rect -91 1139 5 1154
rect 3789 1221 4284 1233
rect -67 990 0 1139
rect 3789 1087 4185 1221
rect 4271 1087 4284 1221
rect 3789 1058 4284 1087
rect 4479 1074 4535 1078
rect 4389 1053 4562 1074
rect 4389 918 4411 1053
rect 4512 918 4562 1053
rect 4389 895 4562 918
rect 4760 1052 4906 1073
rect 4760 917 4782 1052
rect 4883 917 4906 1052
rect 4389 894 4534 895
rect 4760 894 4906 917
rect 5184 1051 5330 1072
rect 5184 916 5206 1051
rect 5307 916 5330 1051
rect 4760 893 4905 894
rect 5184 893 5330 916
rect 5570 1038 5716 1059
rect 5570 903 5592 1038
rect 5693 903 5716 1038
rect 5184 892 5329 893
rect 5570 880 5716 903
rect 5952 1051 6098 1072
rect 5952 916 5974 1051
rect 6075 916 6098 1051
rect 5952 893 6098 916
rect 5952 892 6097 893
rect 5570 879 5715 880
rect 3208 499 3359 546
rect -470 242 -355 246
rect 6367 242 6511 245
rect -470 200 6511 242
rect -470 62 -453 200
rect -383 199 6511 200
rect -383 62 -253 199
rect -470 56 -253 62
rect -173 185 6511 199
rect -173 56 4404 185
rect -470 50 4404 56
rect 4505 184 6511 185
rect 4505 50 4775 184
rect -470 49 4775 50
rect 4876 183 6511 184
rect 4876 49 5199 183
rect -470 48 5199 49
rect 5300 170 5967 183
rect 5300 48 5585 170
rect -470 35 5585 48
rect 5686 48 5967 170
rect 6068 48 6511 183
rect 5686 35 6511 48
rect -470 -147 6511 35
rect -470 -148 6374 -147
<< via1 >>
rect -313 5171 -237 5270
rect -63 5164 13 5263
rect 4370 5224 4475 5362
rect 4742 5221 4847 5359
rect 5214 5221 5319 5359
rect 5539 5221 5644 5359
rect 5842 5221 5947 5359
rect -313 3869 -237 3968
rect -58 3837 9 3890
rect 4370 3966 4475 4104
rect 4742 3963 4847 4101
rect 5214 3963 5319 4101
rect 5539 3963 5644 4101
rect 5842 3963 5947 4101
rect -60 3272 7 3325
rect 4191 3324 4269 3428
rect -457 3025 -386 3104
rect -151 3025 -85 3095
rect 28 3048 86 3109
rect -454 2644 -393 2705
rect 214 2617 294 2732
rect 4024 2666 4082 2718
rect 4033 2490 4091 2542
rect -460 2240 -390 2340
rect 215 2228 295 2343
rect 6431 2468 6495 2523
rect 4022 2256 4080 2308
rect 5987 2251 6039 2325
rect -458 1861 -387 1940
rect -149 1866 -83 1936
rect 29 1860 85 1914
rect 4198 1866 4259 1943
rect -73 1716 -9 1773
rect 4443 1301 4557 1401
rect -76 1154 -12 1211
rect 4185 1087 4271 1221
rect 4411 918 4512 1053
rect 4782 917 4883 1052
rect 5206 916 5307 1051
rect 5592 903 5693 1038
rect 5974 916 6075 1051
rect -453 62 -383 200
rect -253 56 -173 199
rect 4404 50 4505 185
rect 4775 49 4876 184
rect 5199 48 5300 183
rect 5585 35 5686 170
rect 5967 48 6068 183
<< metal2 >>
rect 4355 5362 4491 5389
rect -326 5270 -227 5283
rect -326 5171 -313 5270
rect -237 5171 -227 5270
rect -326 3975 -227 5171
rect -75 5263 24 5287
rect -75 5164 -63 5263
rect 13 5164 24 5263
rect -340 3968 -214 3975
rect -340 3869 -313 3968
rect -237 3869 -214 3968
rect -75 3911 24 5164
rect 4355 5224 4370 5362
rect 4475 5224 4491 5362
rect 4355 4104 4491 5224
rect 4355 3966 4370 4104
rect 4475 3966 4491 4104
rect 4355 3914 4491 3966
rect 4727 5359 4860 5386
rect 4727 5221 4742 5359
rect 4847 5221 4860 5359
rect 4727 4101 4860 5221
rect 4727 3963 4742 4101
rect 4847 3963 4860 4101
rect 4727 3911 4860 3963
rect 5199 5359 5332 5386
rect 5199 5221 5214 5359
rect 5319 5221 5332 5359
rect 5199 4101 5332 5221
rect 5199 3963 5214 4101
rect 5319 3963 5332 4101
rect 5199 3911 5332 3963
rect 5524 5359 5657 5386
rect 5524 5221 5539 5359
rect 5644 5221 5657 5359
rect 5524 4101 5657 5221
rect 5524 3963 5539 4101
rect 5644 3963 5657 4101
rect 5524 3911 5657 3963
rect 5827 5359 5960 5386
rect 5827 5221 5842 5359
rect 5947 5221 5960 5359
rect 5827 4101 5960 5221
rect 5827 3963 5842 4101
rect 5947 3963 5960 4101
rect 5827 3911 5960 3963
rect -340 3849 -214 3869
rect -73 3890 21 3911
rect -73 3837 -58 3890
rect 9 3837 21 3890
rect -73 3325 21 3837
rect -73 3272 -60 3325
rect 7 3272 21 3325
rect 4170 3428 4289 3442
rect 4170 3324 4191 3428
rect 4269 3324 4289 3428
rect 4170 3301 4289 3324
rect -73 3261 21 3272
rect -472 3104 -373 3118
rect -472 3025 -457 3104
rect -386 3025 -373 3104
rect -472 2705 -373 3025
rect -472 2644 -454 2705
rect -393 2644 -373 2705
rect -472 2340 -373 2644
rect -472 2240 -460 2340
rect -390 2240 -373 2340
rect -472 1940 -373 2240
rect -179 3095 -65 3117
rect -179 3025 -151 3095
rect -85 3025 -65 3095
rect -179 1961 -65 3025
rect -472 1861 -458 1940
rect -387 1861 -373 1940
rect -472 1846 -373 1861
rect -269 1936 -65 1961
rect -269 1866 -149 1936
rect -83 1866 -65 1936
rect -269 1847 -65 1866
rect 17 3109 97 3117
rect 17 3048 28 3109
rect 86 3048 97 3109
rect 17 1914 97 3048
rect 204 2732 310 2754
rect 204 2617 214 2732
rect 294 2617 310 2732
rect 204 2603 310 2617
rect 4010 2731 4100 2732
rect 4010 2718 4101 2731
rect 4010 2666 4024 2718
rect 4082 2666 4101 2718
rect 204 2363 286 2603
rect 4010 2542 4101 2666
rect 4010 2490 4033 2542
rect 4091 2490 4101 2542
rect 204 2343 311 2363
rect 204 2228 215 2343
rect 295 2228 311 2343
rect 4010 2308 4101 2490
rect 4171 2456 4279 3301
rect 6362 2523 6519 2535
rect 6362 2468 6431 2523
rect 6495 2468 6519 2523
rect 4171 2347 6043 2456
rect 6362 2454 6519 2468
rect 4171 2346 4279 2347
rect 4010 2256 4022 2308
rect 4080 2256 4101 2308
rect 4010 2243 4101 2256
rect 5934 2325 6043 2347
rect 5934 2251 5987 2325
rect 6039 2251 6043 2325
rect 4010 2242 4100 2243
rect 5934 2237 6043 2251
rect 204 2211 311 2228
rect 6415 1988 6519 2454
rect 17 1860 29 1914
rect 85 1860 97 1914
rect 17 1851 97 1860
rect 4170 1943 4282 1965
rect 4170 1866 4198 1943
rect 4259 1866 4282 1943
rect -470 246 -374 1846
rect -470 200 -355 246
rect -470 62 -453 200
rect -383 62 -355 200
rect -470 -148 -355 62
rect -269 199 -160 1847
rect 4170 1839 4282 1866
rect 4388 1884 6519 1988
rect -91 1773 6 1786
rect -91 1716 -73 1773
rect -9 1716 6 1773
rect -91 1211 6 1716
rect -91 1154 -76 1211
rect -12 1154 6 1211
rect -91 1139 6 1154
rect 4170 1221 4284 1839
rect 4388 1412 4492 1884
rect 4388 1401 4590 1412
rect 4388 1301 4443 1401
rect 4557 1301 4590 1401
rect 4388 1288 4590 1301
rect 4170 1087 4185 1221
rect 4271 1087 4284 1221
rect 4170 1058 4284 1087
rect 4389 1053 4534 1074
rect 4389 918 4411 1053
rect 4512 918 4534 1053
rect 4389 894 4534 918
rect 4760 1052 4905 1073
rect 4760 917 4782 1052
rect 4883 917 4905 1052
rect -269 56 -253 199
rect -173 56 -160 199
rect -269 -146 -160 56
rect 4390 240 4524 894
rect 4760 893 4905 917
rect 5184 1051 5329 1072
rect 5184 916 5206 1051
rect 5307 916 5329 1051
rect 4390 185 4525 240
rect 4390 50 4404 185
rect 4505 50 4525 185
rect 4390 0 4525 50
rect 4761 239 4895 893
rect 5184 892 5329 916
rect 5570 1038 5715 1059
rect 5570 903 5592 1038
rect 5693 903 5715 1038
rect 4761 184 4896 239
rect 4761 49 4775 184
rect 4876 49 4896 184
rect 4761 5 4896 49
rect 5185 238 5319 892
rect 5570 879 5715 903
rect 5952 1051 6097 1072
rect 5952 916 5974 1051
rect 6075 916 6097 1051
rect 5952 892 6097 916
rect 5185 183 5320 238
rect 5185 48 5199 183
rect 5300 48 5320 183
rect 5185 4 5320 48
rect 5571 225 5705 879
rect 5953 238 6087 892
rect 5571 170 5706 225
rect 5571 35 5585 170
rect 5686 35 5706 170
rect 5571 -9 5706 35
rect 5953 183 6088 238
rect 5953 48 5967 183
rect 6068 48 6088 183
rect 5953 4 6088 48
use buffer_loading_mag  buffer_loading_mag_0
timestamp 1691670594
transform 1 0 4310 0 1 3120
box -64 -176 1693 1032
use buffer_loading_mag  buffer_loading_mag_1
timestamp 1691670594
transform 1 0 4449 0 1 1071
box -64 -176 1693 1032
use buffer_mag  buffer_mag_0
timestamp 1691809051
transform -1 0 6016 0 -1 3136
box -110 0 1928 1300
use DFF_  DFF__0
timestamp 1695119997
transform 1 0 364 0 1 -146
box -365 146 3828 2594
use DFF_  DFF__1
timestamp 1695119997
transform 1 0 363 0 -1 5112
box -365 146 3828 2594
use inv  inv_0
timestamp 1695119997
transform 1 0 -398 0 1 2946
box -61 58 345 1028
use inv  inv_1
timestamp 1695119997
transform 1 0 -411 0 -1 2018
box -61 58 345 1028
use inv_my_mag  inv_my_mag_0
timestamp 1695119997
transform 1 0 -398 0 1 2946
box -61 58 345 1028
use inv_my_mag  inv_my_mag_1
timestamp 1695119997
transform 1 0 -411 0 -1 2018
box -61 58 345 1028
use nand2  nand2_0
timestamp 1694691991
transform -1 0 6506 0 -1 2788
box -70 -188 502 863
<< labels >>
flabel metal1 6563 1364 6563 1364 0 FreeSans 640 0 0 0 PD
port 0 nsew
flabel metal1 6538 3418 6538 3418 0 FreeSans 640 0 0 0 PU
port 1 nsew
flabel metal1 2659 5365 2659 5365 0 FreeSans 640 0 0 0 VDD
port 2 nsew
flabel metal1 2686 -25 2686 -25 0 FreeSans 640 0 0 0 VSS
port 3 nsew
flabel metal1 -498 3417 -498 3417 0 FreeSans 640 0 0 0 VREF
port 4 nsew
flabel metal1 -535 1544 -535 1544 0 FreeSans 640 0 0 0 VDIV
port 5 nsew
<< end >>
