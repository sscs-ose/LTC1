magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -9351 -2606 9351 2606
<< metal3 >>
rect -7351 596 7351 606
rect -7351 540 -7341 596
rect -7285 540 -7199 596
rect -7143 540 -7057 596
rect -7001 540 -6915 596
rect -6859 540 -6773 596
rect -6717 540 -6631 596
rect -6575 540 -6489 596
rect -6433 540 -6347 596
rect -6291 540 -6205 596
rect -6149 540 -6063 596
rect -6007 540 -5921 596
rect -5865 540 -5779 596
rect -5723 540 -5637 596
rect -5581 540 -5495 596
rect -5439 540 -5353 596
rect -5297 540 -5211 596
rect -5155 540 -5069 596
rect -5013 540 -4927 596
rect -4871 540 -4785 596
rect -4729 540 -4643 596
rect -4587 540 -4501 596
rect -4445 540 -4359 596
rect -4303 540 -4217 596
rect -4161 540 -4075 596
rect -4019 540 -3933 596
rect -3877 540 -3791 596
rect -3735 540 -3649 596
rect -3593 540 -3507 596
rect -3451 540 -3365 596
rect -3309 540 -3223 596
rect -3167 540 -3081 596
rect -3025 540 -2939 596
rect -2883 540 -2797 596
rect -2741 540 -2655 596
rect -2599 540 -2513 596
rect -2457 540 -2371 596
rect -2315 540 -2229 596
rect -2173 540 -2087 596
rect -2031 540 -1945 596
rect -1889 540 -1803 596
rect -1747 540 -1661 596
rect -1605 540 -1519 596
rect -1463 540 -1377 596
rect -1321 540 -1235 596
rect -1179 540 -1093 596
rect -1037 540 -951 596
rect -895 540 -809 596
rect -753 540 -667 596
rect -611 540 -525 596
rect -469 540 -383 596
rect -327 540 -241 596
rect -185 540 -99 596
rect -43 540 43 596
rect 99 540 185 596
rect 241 540 327 596
rect 383 540 469 596
rect 525 540 611 596
rect 667 540 753 596
rect 809 540 895 596
rect 951 540 1037 596
rect 1093 540 1179 596
rect 1235 540 1321 596
rect 1377 540 1463 596
rect 1519 540 1605 596
rect 1661 540 1747 596
rect 1803 540 1889 596
rect 1945 540 2031 596
rect 2087 540 2173 596
rect 2229 540 2315 596
rect 2371 540 2457 596
rect 2513 540 2599 596
rect 2655 540 2741 596
rect 2797 540 2883 596
rect 2939 540 3025 596
rect 3081 540 3167 596
rect 3223 540 3309 596
rect 3365 540 3451 596
rect 3507 540 3593 596
rect 3649 540 3735 596
rect 3791 540 3877 596
rect 3933 540 4019 596
rect 4075 540 4161 596
rect 4217 540 4303 596
rect 4359 540 4445 596
rect 4501 540 4587 596
rect 4643 540 4729 596
rect 4785 540 4871 596
rect 4927 540 5013 596
rect 5069 540 5155 596
rect 5211 540 5297 596
rect 5353 540 5439 596
rect 5495 540 5581 596
rect 5637 540 5723 596
rect 5779 540 5865 596
rect 5921 540 6007 596
rect 6063 540 6149 596
rect 6205 540 6291 596
rect 6347 540 6433 596
rect 6489 540 6575 596
rect 6631 540 6717 596
rect 6773 540 6859 596
rect 6915 540 7001 596
rect 7057 540 7143 596
rect 7199 540 7285 596
rect 7341 540 7351 596
rect -7351 454 7351 540
rect -7351 398 -7341 454
rect -7285 398 -7199 454
rect -7143 398 -7057 454
rect -7001 398 -6915 454
rect -6859 398 -6773 454
rect -6717 398 -6631 454
rect -6575 398 -6489 454
rect -6433 398 -6347 454
rect -6291 398 -6205 454
rect -6149 398 -6063 454
rect -6007 398 -5921 454
rect -5865 398 -5779 454
rect -5723 398 -5637 454
rect -5581 398 -5495 454
rect -5439 398 -5353 454
rect -5297 398 -5211 454
rect -5155 398 -5069 454
rect -5013 398 -4927 454
rect -4871 398 -4785 454
rect -4729 398 -4643 454
rect -4587 398 -4501 454
rect -4445 398 -4359 454
rect -4303 398 -4217 454
rect -4161 398 -4075 454
rect -4019 398 -3933 454
rect -3877 398 -3791 454
rect -3735 398 -3649 454
rect -3593 398 -3507 454
rect -3451 398 -3365 454
rect -3309 398 -3223 454
rect -3167 398 -3081 454
rect -3025 398 -2939 454
rect -2883 398 -2797 454
rect -2741 398 -2655 454
rect -2599 398 -2513 454
rect -2457 398 -2371 454
rect -2315 398 -2229 454
rect -2173 398 -2087 454
rect -2031 398 -1945 454
rect -1889 398 -1803 454
rect -1747 398 -1661 454
rect -1605 398 -1519 454
rect -1463 398 -1377 454
rect -1321 398 -1235 454
rect -1179 398 -1093 454
rect -1037 398 -951 454
rect -895 398 -809 454
rect -753 398 -667 454
rect -611 398 -525 454
rect -469 398 -383 454
rect -327 398 -241 454
rect -185 398 -99 454
rect -43 398 43 454
rect 99 398 185 454
rect 241 398 327 454
rect 383 398 469 454
rect 525 398 611 454
rect 667 398 753 454
rect 809 398 895 454
rect 951 398 1037 454
rect 1093 398 1179 454
rect 1235 398 1321 454
rect 1377 398 1463 454
rect 1519 398 1605 454
rect 1661 398 1747 454
rect 1803 398 1889 454
rect 1945 398 2031 454
rect 2087 398 2173 454
rect 2229 398 2315 454
rect 2371 398 2457 454
rect 2513 398 2599 454
rect 2655 398 2741 454
rect 2797 398 2883 454
rect 2939 398 3025 454
rect 3081 398 3167 454
rect 3223 398 3309 454
rect 3365 398 3451 454
rect 3507 398 3593 454
rect 3649 398 3735 454
rect 3791 398 3877 454
rect 3933 398 4019 454
rect 4075 398 4161 454
rect 4217 398 4303 454
rect 4359 398 4445 454
rect 4501 398 4587 454
rect 4643 398 4729 454
rect 4785 398 4871 454
rect 4927 398 5013 454
rect 5069 398 5155 454
rect 5211 398 5297 454
rect 5353 398 5439 454
rect 5495 398 5581 454
rect 5637 398 5723 454
rect 5779 398 5865 454
rect 5921 398 6007 454
rect 6063 398 6149 454
rect 6205 398 6291 454
rect 6347 398 6433 454
rect 6489 398 6575 454
rect 6631 398 6717 454
rect 6773 398 6859 454
rect 6915 398 7001 454
rect 7057 398 7143 454
rect 7199 398 7285 454
rect 7341 398 7351 454
rect -7351 312 7351 398
rect -7351 256 -7341 312
rect -7285 256 -7199 312
rect -7143 256 -7057 312
rect -7001 256 -6915 312
rect -6859 256 -6773 312
rect -6717 256 -6631 312
rect -6575 256 -6489 312
rect -6433 256 -6347 312
rect -6291 256 -6205 312
rect -6149 256 -6063 312
rect -6007 256 -5921 312
rect -5865 256 -5779 312
rect -5723 256 -5637 312
rect -5581 256 -5495 312
rect -5439 256 -5353 312
rect -5297 256 -5211 312
rect -5155 256 -5069 312
rect -5013 256 -4927 312
rect -4871 256 -4785 312
rect -4729 256 -4643 312
rect -4587 256 -4501 312
rect -4445 256 -4359 312
rect -4303 256 -4217 312
rect -4161 256 -4075 312
rect -4019 256 -3933 312
rect -3877 256 -3791 312
rect -3735 256 -3649 312
rect -3593 256 -3507 312
rect -3451 256 -3365 312
rect -3309 256 -3223 312
rect -3167 256 -3081 312
rect -3025 256 -2939 312
rect -2883 256 -2797 312
rect -2741 256 -2655 312
rect -2599 256 -2513 312
rect -2457 256 -2371 312
rect -2315 256 -2229 312
rect -2173 256 -2087 312
rect -2031 256 -1945 312
rect -1889 256 -1803 312
rect -1747 256 -1661 312
rect -1605 256 -1519 312
rect -1463 256 -1377 312
rect -1321 256 -1235 312
rect -1179 256 -1093 312
rect -1037 256 -951 312
rect -895 256 -809 312
rect -753 256 -667 312
rect -611 256 -525 312
rect -469 256 -383 312
rect -327 256 -241 312
rect -185 256 -99 312
rect -43 256 43 312
rect 99 256 185 312
rect 241 256 327 312
rect 383 256 469 312
rect 525 256 611 312
rect 667 256 753 312
rect 809 256 895 312
rect 951 256 1037 312
rect 1093 256 1179 312
rect 1235 256 1321 312
rect 1377 256 1463 312
rect 1519 256 1605 312
rect 1661 256 1747 312
rect 1803 256 1889 312
rect 1945 256 2031 312
rect 2087 256 2173 312
rect 2229 256 2315 312
rect 2371 256 2457 312
rect 2513 256 2599 312
rect 2655 256 2741 312
rect 2797 256 2883 312
rect 2939 256 3025 312
rect 3081 256 3167 312
rect 3223 256 3309 312
rect 3365 256 3451 312
rect 3507 256 3593 312
rect 3649 256 3735 312
rect 3791 256 3877 312
rect 3933 256 4019 312
rect 4075 256 4161 312
rect 4217 256 4303 312
rect 4359 256 4445 312
rect 4501 256 4587 312
rect 4643 256 4729 312
rect 4785 256 4871 312
rect 4927 256 5013 312
rect 5069 256 5155 312
rect 5211 256 5297 312
rect 5353 256 5439 312
rect 5495 256 5581 312
rect 5637 256 5723 312
rect 5779 256 5865 312
rect 5921 256 6007 312
rect 6063 256 6149 312
rect 6205 256 6291 312
rect 6347 256 6433 312
rect 6489 256 6575 312
rect 6631 256 6717 312
rect 6773 256 6859 312
rect 6915 256 7001 312
rect 7057 256 7143 312
rect 7199 256 7285 312
rect 7341 256 7351 312
rect -7351 170 7351 256
rect -7351 114 -7341 170
rect -7285 114 -7199 170
rect -7143 114 -7057 170
rect -7001 114 -6915 170
rect -6859 114 -6773 170
rect -6717 114 -6631 170
rect -6575 114 -6489 170
rect -6433 114 -6347 170
rect -6291 114 -6205 170
rect -6149 114 -6063 170
rect -6007 114 -5921 170
rect -5865 114 -5779 170
rect -5723 114 -5637 170
rect -5581 114 -5495 170
rect -5439 114 -5353 170
rect -5297 114 -5211 170
rect -5155 114 -5069 170
rect -5013 114 -4927 170
rect -4871 114 -4785 170
rect -4729 114 -4643 170
rect -4587 114 -4501 170
rect -4445 114 -4359 170
rect -4303 114 -4217 170
rect -4161 114 -4075 170
rect -4019 114 -3933 170
rect -3877 114 -3791 170
rect -3735 114 -3649 170
rect -3593 114 -3507 170
rect -3451 114 -3365 170
rect -3309 114 -3223 170
rect -3167 114 -3081 170
rect -3025 114 -2939 170
rect -2883 114 -2797 170
rect -2741 114 -2655 170
rect -2599 114 -2513 170
rect -2457 114 -2371 170
rect -2315 114 -2229 170
rect -2173 114 -2087 170
rect -2031 114 -1945 170
rect -1889 114 -1803 170
rect -1747 114 -1661 170
rect -1605 114 -1519 170
rect -1463 114 -1377 170
rect -1321 114 -1235 170
rect -1179 114 -1093 170
rect -1037 114 -951 170
rect -895 114 -809 170
rect -753 114 -667 170
rect -611 114 -525 170
rect -469 114 -383 170
rect -327 114 -241 170
rect -185 114 -99 170
rect -43 114 43 170
rect 99 114 185 170
rect 241 114 327 170
rect 383 114 469 170
rect 525 114 611 170
rect 667 114 753 170
rect 809 114 895 170
rect 951 114 1037 170
rect 1093 114 1179 170
rect 1235 114 1321 170
rect 1377 114 1463 170
rect 1519 114 1605 170
rect 1661 114 1747 170
rect 1803 114 1889 170
rect 1945 114 2031 170
rect 2087 114 2173 170
rect 2229 114 2315 170
rect 2371 114 2457 170
rect 2513 114 2599 170
rect 2655 114 2741 170
rect 2797 114 2883 170
rect 2939 114 3025 170
rect 3081 114 3167 170
rect 3223 114 3309 170
rect 3365 114 3451 170
rect 3507 114 3593 170
rect 3649 114 3735 170
rect 3791 114 3877 170
rect 3933 114 4019 170
rect 4075 114 4161 170
rect 4217 114 4303 170
rect 4359 114 4445 170
rect 4501 114 4587 170
rect 4643 114 4729 170
rect 4785 114 4871 170
rect 4927 114 5013 170
rect 5069 114 5155 170
rect 5211 114 5297 170
rect 5353 114 5439 170
rect 5495 114 5581 170
rect 5637 114 5723 170
rect 5779 114 5865 170
rect 5921 114 6007 170
rect 6063 114 6149 170
rect 6205 114 6291 170
rect 6347 114 6433 170
rect 6489 114 6575 170
rect 6631 114 6717 170
rect 6773 114 6859 170
rect 6915 114 7001 170
rect 7057 114 7143 170
rect 7199 114 7285 170
rect 7341 114 7351 170
rect -7351 28 7351 114
rect -7351 -28 -7341 28
rect -7285 -28 -7199 28
rect -7143 -28 -7057 28
rect -7001 -28 -6915 28
rect -6859 -28 -6773 28
rect -6717 -28 -6631 28
rect -6575 -28 -6489 28
rect -6433 -28 -6347 28
rect -6291 -28 -6205 28
rect -6149 -28 -6063 28
rect -6007 -28 -5921 28
rect -5865 -28 -5779 28
rect -5723 -28 -5637 28
rect -5581 -28 -5495 28
rect -5439 -28 -5353 28
rect -5297 -28 -5211 28
rect -5155 -28 -5069 28
rect -5013 -28 -4927 28
rect -4871 -28 -4785 28
rect -4729 -28 -4643 28
rect -4587 -28 -4501 28
rect -4445 -28 -4359 28
rect -4303 -28 -4217 28
rect -4161 -28 -4075 28
rect -4019 -28 -3933 28
rect -3877 -28 -3791 28
rect -3735 -28 -3649 28
rect -3593 -28 -3507 28
rect -3451 -28 -3365 28
rect -3309 -28 -3223 28
rect -3167 -28 -3081 28
rect -3025 -28 -2939 28
rect -2883 -28 -2797 28
rect -2741 -28 -2655 28
rect -2599 -28 -2513 28
rect -2457 -28 -2371 28
rect -2315 -28 -2229 28
rect -2173 -28 -2087 28
rect -2031 -28 -1945 28
rect -1889 -28 -1803 28
rect -1747 -28 -1661 28
rect -1605 -28 -1519 28
rect -1463 -28 -1377 28
rect -1321 -28 -1235 28
rect -1179 -28 -1093 28
rect -1037 -28 -951 28
rect -895 -28 -809 28
rect -753 -28 -667 28
rect -611 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 611 28
rect 667 -28 753 28
rect 809 -28 895 28
rect 951 -28 1037 28
rect 1093 -28 1179 28
rect 1235 -28 1321 28
rect 1377 -28 1463 28
rect 1519 -28 1605 28
rect 1661 -28 1747 28
rect 1803 -28 1889 28
rect 1945 -28 2031 28
rect 2087 -28 2173 28
rect 2229 -28 2315 28
rect 2371 -28 2457 28
rect 2513 -28 2599 28
rect 2655 -28 2741 28
rect 2797 -28 2883 28
rect 2939 -28 3025 28
rect 3081 -28 3167 28
rect 3223 -28 3309 28
rect 3365 -28 3451 28
rect 3507 -28 3593 28
rect 3649 -28 3735 28
rect 3791 -28 3877 28
rect 3933 -28 4019 28
rect 4075 -28 4161 28
rect 4217 -28 4303 28
rect 4359 -28 4445 28
rect 4501 -28 4587 28
rect 4643 -28 4729 28
rect 4785 -28 4871 28
rect 4927 -28 5013 28
rect 5069 -28 5155 28
rect 5211 -28 5297 28
rect 5353 -28 5439 28
rect 5495 -28 5581 28
rect 5637 -28 5723 28
rect 5779 -28 5865 28
rect 5921 -28 6007 28
rect 6063 -28 6149 28
rect 6205 -28 6291 28
rect 6347 -28 6433 28
rect 6489 -28 6575 28
rect 6631 -28 6717 28
rect 6773 -28 6859 28
rect 6915 -28 7001 28
rect 7057 -28 7143 28
rect 7199 -28 7285 28
rect 7341 -28 7351 28
rect -7351 -114 7351 -28
rect -7351 -170 -7341 -114
rect -7285 -170 -7199 -114
rect -7143 -170 -7057 -114
rect -7001 -170 -6915 -114
rect -6859 -170 -6773 -114
rect -6717 -170 -6631 -114
rect -6575 -170 -6489 -114
rect -6433 -170 -6347 -114
rect -6291 -170 -6205 -114
rect -6149 -170 -6063 -114
rect -6007 -170 -5921 -114
rect -5865 -170 -5779 -114
rect -5723 -170 -5637 -114
rect -5581 -170 -5495 -114
rect -5439 -170 -5353 -114
rect -5297 -170 -5211 -114
rect -5155 -170 -5069 -114
rect -5013 -170 -4927 -114
rect -4871 -170 -4785 -114
rect -4729 -170 -4643 -114
rect -4587 -170 -4501 -114
rect -4445 -170 -4359 -114
rect -4303 -170 -4217 -114
rect -4161 -170 -4075 -114
rect -4019 -170 -3933 -114
rect -3877 -170 -3791 -114
rect -3735 -170 -3649 -114
rect -3593 -170 -3507 -114
rect -3451 -170 -3365 -114
rect -3309 -170 -3223 -114
rect -3167 -170 -3081 -114
rect -3025 -170 -2939 -114
rect -2883 -170 -2797 -114
rect -2741 -170 -2655 -114
rect -2599 -170 -2513 -114
rect -2457 -170 -2371 -114
rect -2315 -170 -2229 -114
rect -2173 -170 -2087 -114
rect -2031 -170 -1945 -114
rect -1889 -170 -1803 -114
rect -1747 -170 -1661 -114
rect -1605 -170 -1519 -114
rect -1463 -170 -1377 -114
rect -1321 -170 -1235 -114
rect -1179 -170 -1093 -114
rect -1037 -170 -951 -114
rect -895 -170 -809 -114
rect -753 -170 -667 -114
rect -611 -170 -525 -114
rect -469 -170 -383 -114
rect -327 -170 -241 -114
rect -185 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 185 -114
rect 241 -170 327 -114
rect 383 -170 469 -114
rect 525 -170 611 -114
rect 667 -170 753 -114
rect 809 -170 895 -114
rect 951 -170 1037 -114
rect 1093 -170 1179 -114
rect 1235 -170 1321 -114
rect 1377 -170 1463 -114
rect 1519 -170 1605 -114
rect 1661 -170 1747 -114
rect 1803 -170 1889 -114
rect 1945 -170 2031 -114
rect 2087 -170 2173 -114
rect 2229 -170 2315 -114
rect 2371 -170 2457 -114
rect 2513 -170 2599 -114
rect 2655 -170 2741 -114
rect 2797 -170 2883 -114
rect 2939 -170 3025 -114
rect 3081 -170 3167 -114
rect 3223 -170 3309 -114
rect 3365 -170 3451 -114
rect 3507 -170 3593 -114
rect 3649 -170 3735 -114
rect 3791 -170 3877 -114
rect 3933 -170 4019 -114
rect 4075 -170 4161 -114
rect 4217 -170 4303 -114
rect 4359 -170 4445 -114
rect 4501 -170 4587 -114
rect 4643 -170 4729 -114
rect 4785 -170 4871 -114
rect 4927 -170 5013 -114
rect 5069 -170 5155 -114
rect 5211 -170 5297 -114
rect 5353 -170 5439 -114
rect 5495 -170 5581 -114
rect 5637 -170 5723 -114
rect 5779 -170 5865 -114
rect 5921 -170 6007 -114
rect 6063 -170 6149 -114
rect 6205 -170 6291 -114
rect 6347 -170 6433 -114
rect 6489 -170 6575 -114
rect 6631 -170 6717 -114
rect 6773 -170 6859 -114
rect 6915 -170 7001 -114
rect 7057 -170 7143 -114
rect 7199 -170 7285 -114
rect 7341 -170 7351 -114
rect -7351 -256 7351 -170
rect -7351 -312 -7341 -256
rect -7285 -312 -7199 -256
rect -7143 -312 -7057 -256
rect -7001 -312 -6915 -256
rect -6859 -312 -6773 -256
rect -6717 -312 -6631 -256
rect -6575 -312 -6489 -256
rect -6433 -312 -6347 -256
rect -6291 -312 -6205 -256
rect -6149 -312 -6063 -256
rect -6007 -312 -5921 -256
rect -5865 -312 -5779 -256
rect -5723 -312 -5637 -256
rect -5581 -312 -5495 -256
rect -5439 -312 -5353 -256
rect -5297 -312 -5211 -256
rect -5155 -312 -5069 -256
rect -5013 -312 -4927 -256
rect -4871 -312 -4785 -256
rect -4729 -312 -4643 -256
rect -4587 -312 -4501 -256
rect -4445 -312 -4359 -256
rect -4303 -312 -4217 -256
rect -4161 -312 -4075 -256
rect -4019 -312 -3933 -256
rect -3877 -312 -3791 -256
rect -3735 -312 -3649 -256
rect -3593 -312 -3507 -256
rect -3451 -312 -3365 -256
rect -3309 -312 -3223 -256
rect -3167 -312 -3081 -256
rect -3025 -312 -2939 -256
rect -2883 -312 -2797 -256
rect -2741 -312 -2655 -256
rect -2599 -312 -2513 -256
rect -2457 -312 -2371 -256
rect -2315 -312 -2229 -256
rect -2173 -312 -2087 -256
rect -2031 -312 -1945 -256
rect -1889 -312 -1803 -256
rect -1747 -312 -1661 -256
rect -1605 -312 -1519 -256
rect -1463 -312 -1377 -256
rect -1321 -312 -1235 -256
rect -1179 -312 -1093 -256
rect -1037 -312 -951 -256
rect -895 -312 -809 -256
rect -753 -312 -667 -256
rect -611 -312 -525 -256
rect -469 -312 -383 -256
rect -327 -312 -241 -256
rect -185 -312 -99 -256
rect -43 -312 43 -256
rect 99 -312 185 -256
rect 241 -312 327 -256
rect 383 -312 469 -256
rect 525 -312 611 -256
rect 667 -312 753 -256
rect 809 -312 895 -256
rect 951 -312 1037 -256
rect 1093 -312 1179 -256
rect 1235 -312 1321 -256
rect 1377 -312 1463 -256
rect 1519 -312 1605 -256
rect 1661 -312 1747 -256
rect 1803 -312 1889 -256
rect 1945 -312 2031 -256
rect 2087 -312 2173 -256
rect 2229 -312 2315 -256
rect 2371 -312 2457 -256
rect 2513 -312 2599 -256
rect 2655 -312 2741 -256
rect 2797 -312 2883 -256
rect 2939 -312 3025 -256
rect 3081 -312 3167 -256
rect 3223 -312 3309 -256
rect 3365 -312 3451 -256
rect 3507 -312 3593 -256
rect 3649 -312 3735 -256
rect 3791 -312 3877 -256
rect 3933 -312 4019 -256
rect 4075 -312 4161 -256
rect 4217 -312 4303 -256
rect 4359 -312 4445 -256
rect 4501 -312 4587 -256
rect 4643 -312 4729 -256
rect 4785 -312 4871 -256
rect 4927 -312 5013 -256
rect 5069 -312 5155 -256
rect 5211 -312 5297 -256
rect 5353 -312 5439 -256
rect 5495 -312 5581 -256
rect 5637 -312 5723 -256
rect 5779 -312 5865 -256
rect 5921 -312 6007 -256
rect 6063 -312 6149 -256
rect 6205 -312 6291 -256
rect 6347 -312 6433 -256
rect 6489 -312 6575 -256
rect 6631 -312 6717 -256
rect 6773 -312 6859 -256
rect 6915 -312 7001 -256
rect 7057 -312 7143 -256
rect 7199 -312 7285 -256
rect 7341 -312 7351 -256
rect -7351 -398 7351 -312
rect -7351 -454 -7341 -398
rect -7285 -454 -7199 -398
rect -7143 -454 -7057 -398
rect -7001 -454 -6915 -398
rect -6859 -454 -6773 -398
rect -6717 -454 -6631 -398
rect -6575 -454 -6489 -398
rect -6433 -454 -6347 -398
rect -6291 -454 -6205 -398
rect -6149 -454 -6063 -398
rect -6007 -454 -5921 -398
rect -5865 -454 -5779 -398
rect -5723 -454 -5637 -398
rect -5581 -454 -5495 -398
rect -5439 -454 -5353 -398
rect -5297 -454 -5211 -398
rect -5155 -454 -5069 -398
rect -5013 -454 -4927 -398
rect -4871 -454 -4785 -398
rect -4729 -454 -4643 -398
rect -4587 -454 -4501 -398
rect -4445 -454 -4359 -398
rect -4303 -454 -4217 -398
rect -4161 -454 -4075 -398
rect -4019 -454 -3933 -398
rect -3877 -454 -3791 -398
rect -3735 -454 -3649 -398
rect -3593 -454 -3507 -398
rect -3451 -454 -3365 -398
rect -3309 -454 -3223 -398
rect -3167 -454 -3081 -398
rect -3025 -454 -2939 -398
rect -2883 -454 -2797 -398
rect -2741 -454 -2655 -398
rect -2599 -454 -2513 -398
rect -2457 -454 -2371 -398
rect -2315 -454 -2229 -398
rect -2173 -454 -2087 -398
rect -2031 -454 -1945 -398
rect -1889 -454 -1803 -398
rect -1747 -454 -1661 -398
rect -1605 -454 -1519 -398
rect -1463 -454 -1377 -398
rect -1321 -454 -1235 -398
rect -1179 -454 -1093 -398
rect -1037 -454 -951 -398
rect -895 -454 -809 -398
rect -753 -454 -667 -398
rect -611 -454 -525 -398
rect -469 -454 -383 -398
rect -327 -454 -241 -398
rect -185 -454 -99 -398
rect -43 -454 43 -398
rect 99 -454 185 -398
rect 241 -454 327 -398
rect 383 -454 469 -398
rect 525 -454 611 -398
rect 667 -454 753 -398
rect 809 -454 895 -398
rect 951 -454 1037 -398
rect 1093 -454 1179 -398
rect 1235 -454 1321 -398
rect 1377 -454 1463 -398
rect 1519 -454 1605 -398
rect 1661 -454 1747 -398
rect 1803 -454 1889 -398
rect 1945 -454 2031 -398
rect 2087 -454 2173 -398
rect 2229 -454 2315 -398
rect 2371 -454 2457 -398
rect 2513 -454 2599 -398
rect 2655 -454 2741 -398
rect 2797 -454 2883 -398
rect 2939 -454 3025 -398
rect 3081 -454 3167 -398
rect 3223 -454 3309 -398
rect 3365 -454 3451 -398
rect 3507 -454 3593 -398
rect 3649 -454 3735 -398
rect 3791 -454 3877 -398
rect 3933 -454 4019 -398
rect 4075 -454 4161 -398
rect 4217 -454 4303 -398
rect 4359 -454 4445 -398
rect 4501 -454 4587 -398
rect 4643 -454 4729 -398
rect 4785 -454 4871 -398
rect 4927 -454 5013 -398
rect 5069 -454 5155 -398
rect 5211 -454 5297 -398
rect 5353 -454 5439 -398
rect 5495 -454 5581 -398
rect 5637 -454 5723 -398
rect 5779 -454 5865 -398
rect 5921 -454 6007 -398
rect 6063 -454 6149 -398
rect 6205 -454 6291 -398
rect 6347 -454 6433 -398
rect 6489 -454 6575 -398
rect 6631 -454 6717 -398
rect 6773 -454 6859 -398
rect 6915 -454 7001 -398
rect 7057 -454 7143 -398
rect 7199 -454 7285 -398
rect 7341 -454 7351 -398
rect -7351 -540 7351 -454
rect -7351 -596 -7341 -540
rect -7285 -596 -7199 -540
rect -7143 -596 -7057 -540
rect -7001 -596 -6915 -540
rect -6859 -596 -6773 -540
rect -6717 -596 -6631 -540
rect -6575 -596 -6489 -540
rect -6433 -596 -6347 -540
rect -6291 -596 -6205 -540
rect -6149 -596 -6063 -540
rect -6007 -596 -5921 -540
rect -5865 -596 -5779 -540
rect -5723 -596 -5637 -540
rect -5581 -596 -5495 -540
rect -5439 -596 -5353 -540
rect -5297 -596 -5211 -540
rect -5155 -596 -5069 -540
rect -5013 -596 -4927 -540
rect -4871 -596 -4785 -540
rect -4729 -596 -4643 -540
rect -4587 -596 -4501 -540
rect -4445 -596 -4359 -540
rect -4303 -596 -4217 -540
rect -4161 -596 -4075 -540
rect -4019 -596 -3933 -540
rect -3877 -596 -3791 -540
rect -3735 -596 -3649 -540
rect -3593 -596 -3507 -540
rect -3451 -596 -3365 -540
rect -3309 -596 -3223 -540
rect -3167 -596 -3081 -540
rect -3025 -596 -2939 -540
rect -2883 -596 -2797 -540
rect -2741 -596 -2655 -540
rect -2599 -596 -2513 -540
rect -2457 -596 -2371 -540
rect -2315 -596 -2229 -540
rect -2173 -596 -2087 -540
rect -2031 -596 -1945 -540
rect -1889 -596 -1803 -540
rect -1747 -596 -1661 -540
rect -1605 -596 -1519 -540
rect -1463 -596 -1377 -540
rect -1321 -596 -1235 -540
rect -1179 -596 -1093 -540
rect -1037 -596 -951 -540
rect -895 -596 -809 -540
rect -753 -596 -667 -540
rect -611 -596 -525 -540
rect -469 -596 -383 -540
rect -327 -596 -241 -540
rect -185 -596 -99 -540
rect -43 -596 43 -540
rect 99 -596 185 -540
rect 241 -596 327 -540
rect 383 -596 469 -540
rect 525 -596 611 -540
rect 667 -596 753 -540
rect 809 -596 895 -540
rect 951 -596 1037 -540
rect 1093 -596 1179 -540
rect 1235 -596 1321 -540
rect 1377 -596 1463 -540
rect 1519 -596 1605 -540
rect 1661 -596 1747 -540
rect 1803 -596 1889 -540
rect 1945 -596 2031 -540
rect 2087 -596 2173 -540
rect 2229 -596 2315 -540
rect 2371 -596 2457 -540
rect 2513 -596 2599 -540
rect 2655 -596 2741 -540
rect 2797 -596 2883 -540
rect 2939 -596 3025 -540
rect 3081 -596 3167 -540
rect 3223 -596 3309 -540
rect 3365 -596 3451 -540
rect 3507 -596 3593 -540
rect 3649 -596 3735 -540
rect 3791 -596 3877 -540
rect 3933 -596 4019 -540
rect 4075 -596 4161 -540
rect 4217 -596 4303 -540
rect 4359 -596 4445 -540
rect 4501 -596 4587 -540
rect 4643 -596 4729 -540
rect 4785 -596 4871 -540
rect 4927 -596 5013 -540
rect 5069 -596 5155 -540
rect 5211 -596 5297 -540
rect 5353 -596 5439 -540
rect 5495 -596 5581 -540
rect 5637 -596 5723 -540
rect 5779 -596 5865 -540
rect 5921 -596 6007 -540
rect 6063 -596 6149 -540
rect 6205 -596 6291 -540
rect 6347 -596 6433 -540
rect 6489 -596 6575 -540
rect 6631 -596 6717 -540
rect 6773 -596 6859 -540
rect 6915 -596 7001 -540
rect 7057 -596 7143 -540
rect 7199 -596 7285 -540
rect 7341 -596 7351 -540
rect -7351 -606 7351 -596
<< via3 >>
rect -7341 540 -7285 596
rect -7199 540 -7143 596
rect -7057 540 -7001 596
rect -6915 540 -6859 596
rect -6773 540 -6717 596
rect -6631 540 -6575 596
rect -6489 540 -6433 596
rect -6347 540 -6291 596
rect -6205 540 -6149 596
rect -6063 540 -6007 596
rect -5921 540 -5865 596
rect -5779 540 -5723 596
rect -5637 540 -5581 596
rect -5495 540 -5439 596
rect -5353 540 -5297 596
rect -5211 540 -5155 596
rect -5069 540 -5013 596
rect -4927 540 -4871 596
rect -4785 540 -4729 596
rect -4643 540 -4587 596
rect -4501 540 -4445 596
rect -4359 540 -4303 596
rect -4217 540 -4161 596
rect -4075 540 -4019 596
rect -3933 540 -3877 596
rect -3791 540 -3735 596
rect -3649 540 -3593 596
rect -3507 540 -3451 596
rect -3365 540 -3309 596
rect -3223 540 -3167 596
rect -3081 540 -3025 596
rect -2939 540 -2883 596
rect -2797 540 -2741 596
rect -2655 540 -2599 596
rect -2513 540 -2457 596
rect -2371 540 -2315 596
rect -2229 540 -2173 596
rect -2087 540 -2031 596
rect -1945 540 -1889 596
rect -1803 540 -1747 596
rect -1661 540 -1605 596
rect -1519 540 -1463 596
rect -1377 540 -1321 596
rect -1235 540 -1179 596
rect -1093 540 -1037 596
rect -951 540 -895 596
rect -809 540 -753 596
rect -667 540 -611 596
rect -525 540 -469 596
rect -383 540 -327 596
rect -241 540 -185 596
rect -99 540 -43 596
rect 43 540 99 596
rect 185 540 241 596
rect 327 540 383 596
rect 469 540 525 596
rect 611 540 667 596
rect 753 540 809 596
rect 895 540 951 596
rect 1037 540 1093 596
rect 1179 540 1235 596
rect 1321 540 1377 596
rect 1463 540 1519 596
rect 1605 540 1661 596
rect 1747 540 1803 596
rect 1889 540 1945 596
rect 2031 540 2087 596
rect 2173 540 2229 596
rect 2315 540 2371 596
rect 2457 540 2513 596
rect 2599 540 2655 596
rect 2741 540 2797 596
rect 2883 540 2939 596
rect 3025 540 3081 596
rect 3167 540 3223 596
rect 3309 540 3365 596
rect 3451 540 3507 596
rect 3593 540 3649 596
rect 3735 540 3791 596
rect 3877 540 3933 596
rect 4019 540 4075 596
rect 4161 540 4217 596
rect 4303 540 4359 596
rect 4445 540 4501 596
rect 4587 540 4643 596
rect 4729 540 4785 596
rect 4871 540 4927 596
rect 5013 540 5069 596
rect 5155 540 5211 596
rect 5297 540 5353 596
rect 5439 540 5495 596
rect 5581 540 5637 596
rect 5723 540 5779 596
rect 5865 540 5921 596
rect 6007 540 6063 596
rect 6149 540 6205 596
rect 6291 540 6347 596
rect 6433 540 6489 596
rect 6575 540 6631 596
rect 6717 540 6773 596
rect 6859 540 6915 596
rect 7001 540 7057 596
rect 7143 540 7199 596
rect 7285 540 7341 596
rect -7341 398 -7285 454
rect -7199 398 -7143 454
rect -7057 398 -7001 454
rect -6915 398 -6859 454
rect -6773 398 -6717 454
rect -6631 398 -6575 454
rect -6489 398 -6433 454
rect -6347 398 -6291 454
rect -6205 398 -6149 454
rect -6063 398 -6007 454
rect -5921 398 -5865 454
rect -5779 398 -5723 454
rect -5637 398 -5581 454
rect -5495 398 -5439 454
rect -5353 398 -5297 454
rect -5211 398 -5155 454
rect -5069 398 -5013 454
rect -4927 398 -4871 454
rect -4785 398 -4729 454
rect -4643 398 -4587 454
rect -4501 398 -4445 454
rect -4359 398 -4303 454
rect -4217 398 -4161 454
rect -4075 398 -4019 454
rect -3933 398 -3877 454
rect -3791 398 -3735 454
rect -3649 398 -3593 454
rect -3507 398 -3451 454
rect -3365 398 -3309 454
rect -3223 398 -3167 454
rect -3081 398 -3025 454
rect -2939 398 -2883 454
rect -2797 398 -2741 454
rect -2655 398 -2599 454
rect -2513 398 -2457 454
rect -2371 398 -2315 454
rect -2229 398 -2173 454
rect -2087 398 -2031 454
rect -1945 398 -1889 454
rect -1803 398 -1747 454
rect -1661 398 -1605 454
rect -1519 398 -1463 454
rect -1377 398 -1321 454
rect -1235 398 -1179 454
rect -1093 398 -1037 454
rect -951 398 -895 454
rect -809 398 -753 454
rect -667 398 -611 454
rect -525 398 -469 454
rect -383 398 -327 454
rect -241 398 -185 454
rect -99 398 -43 454
rect 43 398 99 454
rect 185 398 241 454
rect 327 398 383 454
rect 469 398 525 454
rect 611 398 667 454
rect 753 398 809 454
rect 895 398 951 454
rect 1037 398 1093 454
rect 1179 398 1235 454
rect 1321 398 1377 454
rect 1463 398 1519 454
rect 1605 398 1661 454
rect 1747 398 1803 454
rect 1889 398 1945 454
rect 2031 398 2087 454
rect 2173 398 2229 454
rect 2315 398 2371 454
rect 2457 398 2513 454
rect 2599 398 2655 454
rect 2741 398 2797 454
rect 2883 398 2939 454
rect 3025 398 3081 454
rect 3167 398 3223 454
rect 3309 398 3365 454
rect 3451 398 3507 454
rect 3593 398 3649 454
rect 3735 398 3791 454
rect 3877 398 3933 454
rect 4019 398 4075 454
rect 4161 398 4217 454
rect 4303 398 4359 454
rect 4445 398 4501 454
rect 4587 398 4643 454
rect 4729 398 4785 454
rect 4871 398 4927 454
rect 5013 398 5069 454
rect 5155 398 5211 454
rect 5297 398 5353 454
rect 5439 398 5495 454
rect 5581 398 5637 454
rect 5723 398 5779 454
rect 5865 398 5921 454
rect 6007 398 6063 454
rect 6149 398 6205 454
rect 6291 398 6347 454
rect 6433 398 6489 454
rect 6575 398 6631 454
rect 6717 398 6773 454
rect 6859 398 6915 454
rect 7001 398 7057 454
rect 7143 398 7199 454
rect 7285 398 7341 454
rect -7341 256 -7285 312
rect -7199 256 -7143 312
rect -7057 256 -7001 312
rect -6915 256 -6859 312
rect -6773 256 -6717 312
rect -6631 256 -6575 312
rect -6489 256 -6433 312
rect -6347 256 -6291 312
rect -6205 256 -6149 312
rect -6063 256 -6007 312
rect -5921 256 -5865 312
rect -5779 256 -5723 312
rect -5637 256 -5581 312
rect -5495 256 -5439 312
rect -5353 256 -5297 312
rect -5211 256 -5155 312
rect -5069 256 -5013 312
rect -4927 256 -4871 312
rect -4785 256 -4729 312
rect -4643 256 -4587 312
rect -4501 256 -4445 312
rect -4359 256 -4303 312
rect -4217 256 -4161 312
rect -4075 256 -4019 312
rect -3933 256 -3877 312
rect -3791 256 -3735 312
rect -3649 256 -3593 312
rect -3507 256 -3451 312
rect -3365 256 -3309 312
rect -3223 256 -3167 312
rect -3081 256 -3025 312
rect -2939 256 -2883 312
rect -2797 256 -2741 312
rect -2655 256 -2599 312
rect -2513 256 -2457 312
rect -2371 256 -2315 312
rect -2229 256 -2173 312
rect -2087 256 -2031 312
rect -1945 256 -1889 312
rect -1803 256 -1747 312
rect -1661 256 -1605 312
rect -1519 256 -1463 312
rect -1377 256 -1321 312
rect -1235 256 -1179 312
rect -1093 256 -1037 312
rect -951 256 -895 312
rect -809 256 -753 312
rect -667 256 -611 312
rect -525 256 -469 312
rect -383 256 -327 312
rect -241 256 -185 312
rect -99 256 -43 312
rect 43 256 99 312
rect 185 256 241 312
rect 327 256 383 312
rect 469 256 525 312
rect 611 256 667 312
rect 753 256 809 312
rect 895 256 951 312
rect 1037 256 1093 312
rect 1179 256 1235 312
rect 1321 256 1377 312
rect 1463 256 1519 312
rect 1605 256 1661 312
rect 1747 256 1803 312
rect 1889 256 1945 312
rect 2031 256 2087 312
rect 2173 256 2229 312
rect 2315 256 2371 312
rect 2457 256 2513 312
rect 2599 256 2655 312
rect 2741 256 2797 312
rect 2883 256 2939 312
rect 3025 256 3081 312
rect 3167 256 3223 312
rect 3309 256 3365 312
rect 3451 256 3507 312
rect 3593 256 3649 312
rect 3735 256 3791 312
rect 3877 256 3933 312
rect 4019 256 4075 312
rect 4161 256 4217 312
rect 4303 256 4359 312
rect 4445 256 4501 312
rect 4587 256 4643 312
rect 4729 256 4785 312
rect 4871 256 4927 312
rect 5013 256 5069 312
rect 5155 256 5211 312
rect 5297 256 5353 312
rect 5439 256 5495 312
rect 5581 256 5637 312
rect 5723 256 5779 312
rect 5865 256 5921 312
rect 6007 256 6063 312
rect 6149 256 6205 312
rect 6291 256 6347 312
rect 6433 256 6489 312
rect 6575 256 6631 312
rect 6717 256 6773 312
rect 6859 256 6915 312
rect 7001 256 7057 312
rect 7143 256 7199 312
rect 7285 256 7341 312
rect -7341 114 -7285 170
rect -7199 114 -7143 170
rect -7057 114 -7001 170
rect -6915 114 -6859 170
rect -6773 114 -6717 170
rect -6631 114 -6575 170
rect -6489 114 -6433 170
rect -6347 114 -6291 170
rect -6205 114 -6149 170
rect -6063 114 -6007 170
rect -5921 114 -5865 170
rect -5779 114 -5723 170
rect -5637 114 -5581 170
rect -5495 114 -5439 170
rect -5353 114 -5297 170
rect -5211 114 -5155 170
rect -5069 114 -5013 170
rect -4927 114 -4871 170
rect -4785 114 -4729 170
rect -4643 114 -4587 170
rect -4501 114 -4445 170
rect -4359 114 -4303 170
rect -4217 114 -4161 170
rect -4075 114 -4019 170
rect -3933 114 -3877 170
rect -3791 114 -3735 170
rect -3649 114 -3593 170
rect -3507 114 -3451 170
rect -3365 114 -3309 170
rect -3223 114 -3167 170
rect -3081 114 -3025 170
rect -2939 114 -2883 170
rect -2797 114 -2741 170
rect -2655 114 -2599 170
rect -2513 114 -2457 170
rect -2371 114 -2315 170
rect -2229 114 -2173 170
rect -2087 114 -2031 170
rect -1945 114 -1889 170
rect -1803 114 -1747 170
rect -1661 114 -1605 170
rect -1519 114 -1463 170
rect -1377 114 -1321 170
rect -1235 114 -1179 170
rect -1093 114 -1037 170
rect -951 114 -895 170
rect -809 114 -753 170
rect -667 114 -611 170
rect -525 114 -469 170
rect -383 114 -327 170
rect -241 114 -185 170
rect -99 114 -43 170
rect 43 114 99 170
rect 185 114 241 170
rect 327 114 383 170
rect 469 114 525 170
rect 611 114 667 170
rect 753 114 809 170
rect 895 114 951 170
rect 1037 114 1093 170
rect 1179 114 1235 170
rect 1321 114 1377 170
rect 1463 114 1519 170
rect 1605 114 1661 170
rect 1747 114 1803 170
rect 1889 114 1945 170
rect 2031 114 2087 170
rect 2173 114 2229 170
rect 2315 114 2371 170
rect 2457 114 2513 170
rect 2599 114 2655 170
rect 2741 114 2797 170
rect 2883 114 2939 170
rect 3025 114 3081 170
rect 3167 114 3223 170
rect 3309 114 3365 170
rect 3451 114 3507 170
rect 3593 114 3649 170
rect 3735 114 3791 170
rect 3877 114 3933 170
rect 4019 114 4075 170
rect 4161 114 4217 170
rect 4303 114 4359 170
rect 4445 114 4501 170
rect 4587 114 4643 170
rect 4729 114 4785 170
rect 4871 114 4927 170
rect 5013 114 5069 170
rect 5155 114 5211 170
rect 5297 114 5353 170
rect 5439 114 5495 170
rect 5581 114 5637 170
rect 5723 114 5779 170
rect 5865 114 5921 170
rect 6007 114 6063 170
rect 6149 114 6205 170
rect 6291 114 6347 170
rect 6433 114 6489 170
rect 6575 114 6631 170
rect 6717 114 6773 170
rect 6859 114 6915 170
rect 7001 114 7057 170
rect 7143 114 7199 170
rect 7285 114 7341 170
rect -7341 -28 -7285 28
rect -7199 -28 -7143 28
rect -7057 -28 -7001 28
rect -6915 -28 -6859 28
rect -6773 -28 -6717 28
rect -6631 -28 -6575 28
rect -6489 -28 -6433 28
rect -6347 -28 -6291 28
rect -6205 -28 -6149 28
rect -6063 -28 -6007 28
rect -5921 -28 -5865 28
rect -5779 -28 -5723 28
rect -5637 -28 -5581 28
rect -5495 -28 -5439 28
rect -5353 -28 -5297 28
rect -5211 -28 -5155 28
rect -5069 -28 -5013 28
rect -4927 -28 -4871 28
rect -4785 -28 -4729 28
rect -4643 -28 -4587 28
rect -4501 -28 -4445 28
rect -4359 -28 -4303 28
rect -4217 -28 -4161 28
rect -4075 -28 -4019 28
rect -3933 -28 -3877 28
rect -3791 -28 -3735 28
rect -3649 -28 -3593 28
rect -3507 -28 -3451 28
rect -3365 -28 -3309 28
rect -3223 -28 -3167 28
rect -3081 -28 -3025 28
rect -2939 -28 -2883 28
rect -2797 -28 -2741 28
rect -2655 -28 -2599 28
rect -2513 -28 -2457 28
rect -2371 -28 -2315 28
rect -2229 -28 -2173 28
rect -2087 -28 -2031 28
rect -1945 -28 -1889 28
rect -1803 -28 -1747 28
rect -1661 -28 -1605 28
rect -1519 -28 -1463 28
rect -1377 -28 -1321 28
rect -1235 -28 -1179 28
rect -1093 -28 -1037 28
rect -951 -28 -895 28
rect -809 -28 -753 28
rect -667 -28 -611 28
rect -525 -28 -469 28
rect -383 -28 -327 28
rect -241 -28 -185 28
rect -99 -28 -43 28
rect 43 -28 99 28
rect 185 -28 241 28
rect 327 -28 383 28
rect 469 -28 525 28
rect 611 -28 667 28
rect 753 -28 809 28
rect 895 -28 951 28
rect 1037 -28 1093 28
rect 1179 -28 1235 28
rect 1321 -28 1377 28
rect 1463 -28 1519 28
rect 1605 -28 1661 28
rect 1747 -28 1803 28
rect 1889 -28 1945 28
rect 2031 -28 2087 28
rect 2173 -28 2229 28
rect 2315 -28 2371 28
rect 2457 -28 2513 28
rect 2599 -28 2655 28
rect 2741 -28 2797 28
rect 2883 -28 2939 28
rect 3025 -28 3081 28
rect 3167 -28 3223 28
rect 3309 -28 3365 28
rect 3451 -28 3507 28
rect 3593 -28 3649 28
rect 3735 -28 3791 28
rect 3877 -28 3933 28
rect 4019 -28 4075 28
rect 4161 -28 4217 28
rect 4303 -28 4359 28
rect 4445 -28 4501 28
rect 4587 -28 4643 28
rect 4729 -28 4785 28
rect 4871 -28 4927 28
rect 5013 -28 5069 28
rect 5155 -28 5211 28
rect 5297 -28 5353 28
rect 5439 -28 5495 28
rect 5581 -28 5637 28
rect 5723 -28 5779 28
rect 5865 -28 5921 28
rect 6007 -28 6063 28
rect 6149 -28 6205 28
rect 6291 -28 6347 28
rect 6433 -28 6489 28
rect 6575 -28 6631 28
rect 6717 -28 6773 28
rect 6859 -28 6915 28
rect 7001 -28 7057 28
rect 7143 -28 7199 28
rect 7285 -28 7341 28
rect -7341 -170 -7285 -114
rect -7199 -170 -7143 -114
rect -7057 -170 -7001 -114
rect -6915 -170 -6859 -114
rect -6773 -170 -6717 -114
rect -6631 -170 -6575 -114
rect -6489 -170 -6433 -114
rect -6347 -170 -6291 -114
rect -6205 -170 -6149 -114
rect -6063 -170 -6007 -114
rect -5921 -170 -5865 -114
rect -5779 -170 -5723 -114
rect -5637 -170 -5581 -114
rect -5495 -170 -5439 -114
rect -5353 -170 -5297 -114
rect -5211 -170 -5155 -114
rect -5069 -170 -5013 -114
rect -4927 -170 -4871 -114
rect -4785 -170 -4729 -114
rect -4643 -170 -4587 -114
rect -4501 -170 -4445 -114
rect -4359 -170 -4303 -114
rect -4217 -170 -4161 -114
rect -4075 -170 -4019 -114
rect -3933 -170 -3877 -114
rect -3791 -170 -3735 -114
rect -3649 -170 -3593 -114
rect -3507 -170 -3451 -114
rect -3365 -170 -3309 -114
rect -3223 -170 -3167 -114
rect -3081 -170 -3025 -114
rect -2939 -170 -2883 -114
rect -2797 -170 -2741 -114
rect -2655 -170 -2599 -114
rect -2513 -170 -2457 -114
rect -2371 -170 -2315 -114
rect -2229 -170 -2173 -114
rect -2087 -170 -2031 -114
rect -1945 -170 -1889 -114
rect -1803 -170 -1747 -114
rect -1661 -170 -1605 -114
rect -1519 -170 -1463 -114
rect -1377 -170 -1321 -114
rect -1235 -170 -1179 -114
rect -1093 -170 -1037 -114
rect -951 -170 -895 -114
rect -809 -170 -753 -114
rect -667 -170 -611 -114
rect -525 -170 -469 -114
rect -383 -170 -327 -114
rect -241 -170 -185 -114
rect -99 -170 -43 -114
rect 43 -170 99 -114
rect 185 -170 241 -114
rect 327 -170 383 -114
rect 469 -170 525 -114
rect 611 -170 667 -114
rect 753 -170 809 -114
rect 895 -170 951 -114
rect 1037 -170 1093 -114
rect 1179 -170 1235 -114
rect 1321 -170 1377 -114
rect 1463 -170 1519 -114
rect 1605 -170 1661 -114
rect 1747 -170 1803 -114
rect 1889 -170 1945 -114
rect 2031 -170 2087 -114
rect 2173 -170 2229 -114
rect 2315 -170 2371 -114
rect 2457 -170 2513 -114
rect 2599 -170 2655 -114
rect 2741 -170 2797 -114
rect 2883 -170 2939 -114
rect 3025 -170 3081 -114
rect 3167 -170 3223 -114
rect 3309 -170 3365 -114
rect 3451 -170 3507 -114
rect 3593 -170 3649 -114
rect 3735 -170 3791 -114
rect 3877 -170 3933 -114
rect 4019 -170 4075 -114
rect 4161 -170 4217 -114
rect 4303 -170 4359 -114
rect 4445 -170 4501 -114
rect 4587 -170 4643 -114
rect 4729 -170 4785 -114
rect 4871 -170 4927 -114
rect 5013 -170 5069 -114
rect 5155 -170 5211 -114
rect 5297 -170 5353 -114
rect 5439 -170 5495 -114
rect 5581 -170 5637 -114
rect 5723 -170 5779 -114
rect 5865 -170 5921 -114
rect 6007 -170 6063 -114
rect 6149 -170 6205 -114
rect 6291 -170 6347 -114
rect 6433 -170 6489 -114
rect 6575 -170 6631 -114
rect 6717 -170 6773 -114
rect 6859 -170 6915 -114
rect 7001 -170 7057 -114
rect 7143 -170 7199 -114
rect 7285 -170 7341 -114
rect -7341 -312 -7285 -256
rect -7199 -312 -7143 -256
rect -7057 -312 -7001 -256
rect -6915 -312 -6859 -256
rect -6773 -312 -6717 -256
rect -6631 -312 -6575 -256
rect -6489 -312 -6433 -256
rect -6347 -312 -6291 -256
rect -6205 -312 -6149 -256
rect -6063 -312 -6007 -256
rect -5921 -312 -5865 -256
rect -5779 -312 -5723 -256
rect -5637 -312 -5581 -256
rect -5495 -312 -5439 -256
rect -5353 -312 -5297 -256
rect -5211 -312 -5155 -256
rect -5069 -312 -5013 -256
rect -4927 -312 -4871 -256
rect -4785 -312 -4729 -256
rect -4643 -312 -4587 -256
rect -4501 -312 -4445 -256
rect -4359 -312 -4303 -256
rect -4217 -312 -4161 -256
rect -4075 -312 -4019 -256
rect -3933 -312 -3877 -256
rect -3791 -312 -3735 -256
rect -3649 -312 -3593 -256
rect -3507 -312 -3451 -256
rect -3365 -312 -3309 -256
rect -3223 -312 -3167 -256
rect -3081 -312 -3025 -256
rect -2939 -312 -2883 -256
rect -2797 -312 -2741 -256
rect -2655 -312 -2599 -256
rect -2513 -312 -2457 -256
rect -2371 -312 -2315 -256
rect -2229 -312 -2173 -256
rect -2087 -312 -2031 -256
rect -1945 -312 -1889 -256
rect -1803 -312 -1747 -256
rect -1661 -312 -1605 -256
rect -1519 -312 -1463 -256
rect -1377 -312 -1321 -256
rect -1235 -312 -1179 -256
rect -1093 -312 -1037 -256
rect -951 -312 -895 -256
rect -809 -312 -753 -256
rect -667 -312 -611 -256
rect -525 -312 -469 -256
rect -383 -312 -327 -256
rect -241 -312 -185 -256
rect -99 -312 -43 -256
rect 43 -312 99 -256
rect 185 -312 241 -256
rect 327 -312 383 -256
rect 469 -312 525 -256
rect 611 -312 667 -256
rect 753 -312 809 -256
rect 895 -312 951 -256
rect 1037 -312 1093 -256
rect 1179 -312 1235 -256
rect 1321 -312 1377 -256
rect 1463 -312 1519 -256
rect 1605 -312 1661 -256
rect 1747 -312 1803 -256
rect 1889 -312 1945 -256
rect 2031 -312 2087 -256
rect 2173 -312 2229 -256
rect 2315 -312 2371 -256
rect 2457 -312 2513 -256
rect 2599 -312 2655 -256
rect 2741 -312 2797 -256
rect 2883 -312 2939 -256
rect 3025 -312 3081 -256
rect 3167 -312 3223 -256
rect 3309 -312 3365 -256
rect 3451 -312 3507 -256
rect 3593 -312 3649 -256
rect 3735 -312 3791 -256
rect 3877 -312 3933 -256
rect 4019 -312 4075 -256
rect 4161 -312 4217 -256
rect 4303 -312 4359 -256
rect 4445 -312 4501 -256
rect 4587 -312 4643 -256
rect 4729 -312 4785 -256
rect 4871 -312 4927 -256
rect 5013 -312 5069 -256
rect 5155 -312 5211 -256
rect 5297 -312 5353 -256
rect 5439 -312 5495 -256
rect 5581 -312 5637 -256
rect 5723 -312 5779 -256
rect 5865 -312 5921 -256
rect 6007 -312 6063 -256
rect 6149 -312 6205 -256
rect 6291 -312 6347 -256
rect 6433 -312 6489 -256
rect 6575 -312 6631 -256
rect 6717 -312 6773 -256
rect 6859 -312 6915 -256
rect 7001 -312 7057 -256
rect 7143 -312 7199 -256
rect 7285 -312 7341 -256
rect -7341 -454 -7285 -398
rect -7199 -454 -7143 -398
rect -7057 -454 -7001 -398
rect -6915 -454 -6859 -398
rect -6773 -454 -6717 -398
rect -6631 -454 -6575 -398
rect -6489 -454 -6433 -398
rect -6347 -454 -6291 -398
rect -6205 -454 -6149 -398
rect -6063 -454 -6007 -398
rect -5921 -454 -5865 -398
rect -5779 -454 -5723 -398
rect -5637 -454 -5581 -398
rect -5495 -454 -5439 -398
rect -5353 -454 -5297 -398
rect -5211 -454 -5155 -398
rect -5069 -454 -5013 -398
rect -4927 -454 -4871 -398
rect -4785 -454 -4729 -398
rect -4643 -454 -4587 -398
rect -4501 -454 -4445 -398
rect -4359 -454 -4303 -398
rect -4217 -454 -4161 -398
rect -4075 -454 -4019 -398
rect -3933 -454 -3877 -398
rect -3791 -454 -3735 -398
rect -3649 -454 -3593 -398
rect -3507 -454 -3451 -398
rect -3365 -454 -3309 -398
rect -3223 -454 -3167 -398
rect -3081 -454 -3025 -398
rect -2939 -454 -2883 -398
rect -2797 -454 -2741 -398
rect -2655 -454 -2599 -398
rect -2513 -454 -2457 -398
rect -2371 -454 -2315 -398
rect -2229 -454 -2173 -398
rect -2087 -454 -2031 -398
rect -1945 -454 -1889 -398
rect -1803 -454 -1747 -398
rect -1661 -454 -1605 -398
rect -1519 -454 -1463 -398
rect -1377 -454 -1321 -398
rect -1235 -454 -1179 -398
rect -1093 -454 -1037 -398
rect -951 -454 -895 -398
rect -809 -454 -753 -398
rect -667 -454 -611 -398
rect -525 -454 -469 -398
rect -383 -454 -327 -398
rect -241 -454 -185 -398
rect -99 -454 -43 -398
rect 43 -454 99 -398
rect 185 -454 241 -398
rect 327 -454 383 -398
rect 469 -454 525 -398
rect 611 -454 667 -398
rect 753 -454 809 -398
rect 895 -454 951 -398
rect 1037 -454 1093 -398
rect 1179 -454 1235 -398
rect 1321 -454 1377 -398
rect 1463 -454 1519 -398
rect 1605 -454 1661 -398
rect 1747 -454 1803 -398
rect 1889 -454 1945 -398
rect 2031 -454 2087 -398
rect 2173 -454 2229 -398
rect 2315 -454 2371 -398
rect 2457 -454 2513 -398
rect 2599 -454 2655 -398
rect 2741 -454 2797 -398
rect 2883 -454 2939 -398
rect 3025 -454 3081 -398
rect 3167 -454 3223 -398
rect 3309 -454 3365 -398
rect 3451 -454 3507 -398
rect 3593 -454 3649 -398
rect 3735 -454 3791 -398
rect 3877 -454 3933 -398
rect 4019 -454 4075 -398
rect 4161 -454 4217 -398
rect 4303 -454 4359 -398
rect 4445 -454 4501 -398
rect 4587 -454 4643 -398
rect 4729 -454 4785 -398
rect 4871 -454 4927 -398
rect 5013 -454 5069 -398
rect 5155 -454 5211 -398
rect 5297 -454 5353 -398
rect 5439 -454 5495 -398
rect 5581 -454 5637 -398
rect 5723 -454 5779 -398
rect 5865 -454 5921 -398
rect 6007 -454 6063 -398
rect 6149 -454 6205 -398
rect 6291 -454 6347 -398
rect 6433 -454 6489 -398
rect 6575 -454 6631 -398
rect 6717 -454 6773 -398
rect 6859 -454 6915 -398
rect 7001 -454 7057 -398
rect 7143 -454 7199 -398
rect 7285 -454 7341 -398
rect -7341 -596 -7285 -540
rect -7199 -596 -7143 -540
rect -7057 -596 -7001 -540
rect -6915 -596 -6859 -540
rect -6773 -596 -6717 -540
rect -6631 -596 -6575 -540
rect -6489 -596 -6433 -540
rect -6347 -596 -6291 -540
rect -6205 -596 -6149 -540
rect -6063 -596 -6007 -540
rect -5921 -596 -5865 -540
rect -5779 -596 -5723 -540
rect -5637 -596 -5581 -540
rect -5495 -596 -5439 -540
rect -5353 -596 -5297 -540
rect -5211 -596 -5155 -540
rect -5069 -596 -5013 -540
rect -4927 -596 -4871 -540
rect -4785 -596 -4729 -540
rect -4643 -596 -4587 -540
rect -4501 -596 -4445 -540
rect -4359 -596 -4303 -540
rect -4217 -596 -4161 -540
rect -4075 -596 -4019 -540
rect -3933 -596 -3877 -540
rect -3791 -596 -3735 -540
rect -3649 -596 -3593 -540
rect -3507 -596 -3451 -540
rect -3365 -596 -3309 -540
rect -3223 -596 -3167 -540
rect -3081 -596 -3025 -540
rect -2939 -596 -2883 -540
rect -2797 -596 -2741 -540
rect -2655 -596 -2599 -540
rect -2513 -596 -2457 -540
rect -2371 -596 -2315 -540
rect -2229 -596 -2173 -540
rect -2087 -596 -2031 -540
rect -1945 -596 -1889 -540
rect -1803 -596 -1747 -540
rect -1661 -596 -1605 -540
rect -1519 -596 -1463 -540
rect -1377 -596 -1321 -540
rect -1235 -596 -1179 -540
rect -1093 -596 -1037 -540
rect -951 -596 -895 -540
rect -809 -596 -753 -540
rect -667 -596 -611 -540
rect -525 -596 -469 -540
rect -383 -596 -327 -540
rect -241 -596 -185 -540
rect -99 -596 -43 -540
rect 43 -596 99 -540
rect 185 -596 241 -540
rect 327 -596 383 -540
rect 469 -596 525 -540
rect 611 -596 667 -540
rect 753 -596 809 -540
rect 895 -596 951 -540
rect 1037 -596 1093 -540
rect 1179 -596 1235 -540
rect 1321 -596 1377 -540
rect 1463 -596 1519 -540
rect 1605 -596 1661 -540
rect 1747 -596 1803 -540
rect 1889 -596 1945 -540
rect 2031 -596 2087 -540
rect 2173 -596 2229 -540
rect 2315 -596 2371 -540
rect 2457 -596 2513 -540
rect 2599 -596 2655 -540
rect 2741 -596 2797 -540
rect 2883 -596 2939 -540
rect 3025 -596 3081 -540
rect 3167 -596 3223 -540
rect 3309 -596 3365 -540
rect 3451 -596 3507 -540
rect 3593 -596 3649 -540
rect 3735 -596 3791 -540
rect 3877 -596 3933 -540
rect 4019 -596 4075 -540
rect 4161 -596 4217 -540
rect 4303 -596 4359 -540
rect 4445 -596 4501 -540
rect 4587 -596 4643 -540
rect 4729 -596 4785 -540
rect 4871 -596 4927 -540
rect 5013 -596 5069 -540
rect 5155 -596 5211 -540
rect 5297 -596 5353 -540
rect 5439 -596 5495 -540
rect 5581 -596 5637 -540
rect 5723 -596 5779 -540
rect 5865 -596 5921 -540
rect 6007 -596 6063 -540
rect 6149 -596 6205 -540
rect 6291 -596 6347 -540
rect 6433 -596 6489 -540
rect 6575 -596 6631 -540
rect 6717 -596 6773 -540
rect 6859 -596 6915 -540
rect 7001 -596 7057 -540
rect 7143 -596 7199 -540
rect 7285 -596 7341 -540
<< metal4 >>
rect -7351 596 7351 606
rect -7351 540 -7341 596
rect -7285 540 -7199 596
rect -7143 540 -7057 596
rect -7001 540 -6915 596
rect -6859 540 -6773 596
rect -6717 540 -6631 596
rect -6575 540 -6489 596
rect -6433 540 -6347 596
rect -6291 540 -6205 596
rect -6149 540 -6063 596
rect -6007 540 -5921 596
rect -5865 540 -5779 596
rect -5723 540 -5637 596
rect -5581 540 -5495 596
rect -5439 540 -5353 596
rect -5297 540 -5211 596
rect -5155 540 -5069 596
rect -5013 540 -4927 596
rect -4871 540 -4785 596
rect -4729 540 -4643 596
rect -4587 540 -4501 596
rect -4445 540 -4359 596
rect -4303 540 -4217 596
rect -4161 540 -4075 596
rect -4019 540 -3933 596
rect -3877 540 -3791 596
rect -3735 540 -3649 596
rect -3593 540 -3507 596
rect -3451 540 -3365 596
rect -3309 540 -3223 596
rect -3167 540 -3081 596
rect -3025 540 -2939 596
rect -2883 540 -2797 596
rect -2741 540 -2655 596
rect -2599 540 -2513 596
rect -2457 540 -2371 596
rect -2315 540 -2229 596
rect -2173 540 -2087 596
rect -2031 540 -1945 596
rect -1889 540 -1803 596
rect -1747 540 -1661 596
rect -1605 540 -1519 596
rect -1463 540 -1377 596
rect -1321 540 -1235 596
rect -1179 540 -1093 596
rect -1037 540 -951 596
rect -895 540 -809 596
rect -753 540 -667 596
rect -611 540 -525 596
rect -469 540 -383 596
rect -327 540 -241 596
rect -185 540 -99 596
rect -43 540 43 596
rect 99 540 185 596
rect 241 540 327 596
rect 383 540 469 596
rect 525 540 611 596
rect 667 540 753 596
rect 809 540 895 596
rect 951 540 1037 596
rect 1093 540 1179 596
rect 1235 540 1321 596
rect 1377 540 1463 596
rect 1519 540 1605 596
rect 1661 540 1747 596
rect 1803 540 1889 596
rect 1945 540 2031 596
rect 2087 540 2173 596
rect 2229 540 2315 596
rect 2371 540 2457 596
rect 2513 540 2599 596
rect 2655 540 2741 596
rect 2797 540 2883 596
rect 2939 540 3025 596
rect 3081 540 3167 596
rect 3223 540 3309 596
rect 3365 540 3451 596
rect 3507 540 3593 596
rect 3649 540 3735 596
rect 3791 540 3877 596
rect 3933 540 4019 596
rect 4075 540 4161 596
rect 4217 540 4303 596
rect 4359 540 4445 596
rect 4501 540 4587 596
rect 4643 540 4729 596
rect 4785 540 4871 596
rect 4927 540 5013 596
rect 5069 540 5155 596
rect 5211 540 5297 596
rect 5353 540 5439 596
rect 5495 540 5581 596
rect 5637 540 5723 596
rect 5779 540 5865 596
rect 5921 540 6007 596
rect 6063 540 6149 596
rect 6205 540 6291 596
rect 6347 540 6433 596
rect 6489 540 6575 596
rect 6631 540 6717 596
rect 6773 540 6859 596
rect 6915 540 7001 596
rect 7057 540 7143 596
rect 7199 540 7285 596
rect 7341 540 7351 596
rect -7351 454 7351 540
rect -7351 398 -7341 454
rect -7285 398 -7199 454
rect -7143 398 -7057 454
rect -7001 398 -6915 454
rect -6859 398 -6773 454
rect -6717 398 -6631 454
rect -6575 398 -6489 454
rect -6433 398 -6347 454
rect -6291 398 -6205 454
rect -6149 398 -6063 454
rect -6007 398 -5921 454
rect -5865 398 -5779 454
rect -5723 398 -5637 454
rect -5581 398 -5495 454
rect -5439 398 -5353 454
rect -5297 398 -5211 454
rect -5155 398 -5069 454
rect -5013 398 -4927 454
rect -4871 398 -4785 454
rect -4729 398 -4643 454
rect -4587 398 -4501 454
rect -4445 398 -4359 454
rect -4303 398 -4217 454
rect -4161 398 -4075 454
rect -4019 398 -3933 454
rect -3877 398 -3791 454
rect -3735 398 -3649 454
rect -3593 398 -3507 454
rect -3451 398 -3365 454
rect -3309 398 -3223 454
rect -3167 398 -3081 454
rect -3025 398 -2939 454
rect -2883 398 -2797 454
rect -2741 398 -2655 454
rect -2599 398 -2513 454
rect -2457 398 -2371 454
rect -2315 398 -2229 454
rect -2173 398 -2087 454
rect -2031 398 -1945 454
rect -1889 398 -1803 454
rect -1747 398 -1661 454
rect -1605 398 -1519 454
rect -1463 398 -1377 454
rect -1321 398 -1235 454
rect -1179 398 -1093 454
rect -1037 398 -951 454
rect -895 398 -809 454
rect -753 398 -667 454
rect -611 398 -525 454
rect -469 398 -383 454
rect -327 398 -241 454
rect -185 398 -99 454
rect -43 398 43 454
rect 99 398 185 454
rect 241 398 327 454
rect 383 398 469 454
rect 525 398 611 454
rect 667 398 753 454
rect 809 398 895 454
rect 951 398 1037 454
rect 1093 398 1179 454
rect 1235 398 1321 454
rect 1377 398 1463 454
rect 1519 398 1605 454
rect 1661 398 1747 454
rect 1803 398 1889 454
rect 1945 398 2031 454
rect 2087 398 2173 454
rect 2229 398 2315 454
rect 2371 398 2457 454
rect 2513 398 2599 454
rect 2655 398 2741 454
rect 2797 398 2883 454
rect 2939 398 3025 454
rect 3081 398 3167 454
rect 3223 398 3309 454
rect 3365 398 3451 454
rect 3507 398 3593 454
rect 3649 398 3735 454
rect 3791 398 3877 454
rect 3933 398 4019 454
rect 4075 398 4161 454
rect 4217 398 4303 454
rect 4359 398 4445 454
rect 4501 398 4587 454
rect 4643 398 4729 454
rect 4785 398 4871 454
rect 4927 398 5013 454
rect 5069 398 5155 454
rect 5211 398 5297 454
rect 5353 398 5439 454
rect 5495 398 5581 454
rect 5637 398 5723 454
rect 5779 398 5865 454
rect 5921 398 6007 454
rect 6063 398 6149 454
rect 6205 398 6291 454
rect 6347 398 6433 454
rect 6489 398 6575 454
rect 6631 398 6717 454
rect 6773 398 6859 454
rect 6915 398 7001 454
rect 7057 398 7143 454
rect 7199 398 7285 454
rect 7341 398 7351 454
rect -7351 312 7351 398
rect -7351 256 -7341 312
rect -7285 256 -7199 312
rect -7143 256 -7057 312
rect -7001 256 -6915 312
rect -6859 256 -6773 312
rect -6717 256 -6631 312
rect -6575 256 -6489 312
rect -6433 256 -6347 312
rect -6291 256 -6205 312
rect -6149 256 -6063 312
rect -6007 256 -5921 312
rect -5865 256 -5779 312
rect -5723 256 -5637 312
rect -5581 256 -5495 312
rect -5439 256 -5353 312
rect -5297 256 -5211 312
rect -5155 256 -5069 312
rect -5013 256 -4927 312
rect -4871 256 -4785 312
rect -4729 256 -4643 312
rect -4587 256 -4501 312
rect -4445 256 -4359 312
rect -4303 256 -4217 312
rect -4161 256 -4075 312
rect -4019 256 -3933 312
rect -3877 256 -3791 312
rect -3735 256 -3649 312
rect -3593 256 -3507 312
rect -3451 256 -3365 312
rect -3309 256 -3223 312
rect -3167 256 -3081 312
rect -3025 256 -2939 312
rect -2883 256 -2797 312
rect -2741 256 -2655 312
rect -2599 256 -2513 312
rect -2457 256 -2371 312
rect -2315 256 -2229 312
rect -2173 256 -2087 312
rect -2031 256 -1945 312
rect -1889 256 -1803 312
rect -1747 256 -1661 312
rect -1605 256 -1519 312
rect -1463 256 -1377 312
rect -1321 256 -1235 312
rect -1179 256 -1093 312
rect -1037 256 -951 312
rect -895 256 -809 312
rect -753 256 -667 312
rect -611 256 -525 312
rect -469 256 -383 312
rect -327 256 -241 312
rect -185 256 -99 312
rect -43 256 43 312
rect 99 256 185 312
rect 241 256 327 312
rect 383 256 469 312
rect 525 256 611 312
rect 667 256 753 312
rect 809 256 895 312
rect 951 256 1037 312
rect 1093 256 1179 312
rect 1235 256 1321 312
rect 1377 256 1463 312
rect 1519 256 1605 312
rect 1661 256 1747 312
rect 1803 256 1889 312
rect 1945 256 2031 312
rect 2087 256 2173 312
rect 2229 256 2315 312
rect 2371 256 2457 312
rect 2513 256 2599 312
rect 2655 256 2741 312
rect 2797 256 2883 312
rect 2939 256 3025 312
rect 3081 256 3167 312
rect 3223 256 3309 312
rect 3365 256 3451 312
rect 3507 256 3593 312
rect 3649 256 3735 312
rect 3791 256 3877 312
rect 3933 256 4019 312
rect 4075 256 4161 312
rect 4217 256 4303 312
rect 4359 256 4445 312
rect 4501 256 4587 312
rect 4643 256 4729 312
rect 4785 256 4871 312
rect 4927 256 5013 312
rect 5069 256 5155 312
rect 5211 256 5297 312
rect 5353 256 5439 312
rect 5495 256 5581 312
rect 5637 256 5723 312
rect 5779 256 5865 312
rect 5921 256 6007 312
rect 6063 256 6149 312
rect 6205 256 6291 312
rect 6347 256 6433 312
rect 6489 256 6575 312
rect 6631 256 6717 312
rect 6773 256 6859 312
rect 6915 256 7001 312
rect 7057 256 7143 312
rect 7199 256 7285 312
rect 7341 256 7351 312
rect -7351 170 7351 256
rect -7351 114 -7341 170
rect -7285 114 -7199 170
rect -7143 114 -7057 170
rect -7001 114 -6915 170
rect -6859 114 -6773 170
rect -6717 114 -6631 170
rect -6575 114 -6489 170
rect -6433 114 -6347 170
rect -6291 114 -6205 170
rect -6149 114 -6063 170
rect -6007 114 -5921 170
rect -5865 114 -5779 170
rect -5723 114 -5637 170
rect -5581 114 -5495 170
rect -5439 114 -5353 170
rect -5297 114 -5211 170
rect -5155 114 -5069 170
rect -5013 114 -4927 170
rect -4871 114 -4785 170
rect -4729 114 -4643 170
rect -4587 114 -4501 170
rect -4445 114 -4359 170
rect -4303 114 -4217 170
rect -4161 114 -4075 170
rect -4019 114 -3933 170
rect -3877 114 -3791 170
rect -3735 114 -3649 170
rect -3593 114 -3507 170
rect -3451 114 -3365 170
rect -3309 114 -3223 170
rect -3167 114 -3081 170
rect -3025 114 -2939 170
rect -2883 114 -2797 170
rect -2741 114 -2655 170
rect -2599 114 -2513 170
rect -2457 114 -2371 170
rect -2315 114 -2229 170
rect -2173 114 -2087 170
rect -2031 114 -1945 170
rect -1889 114 -1803 170
rect -1747 114 -1661 170
rect -1605 114 -1519 170
rect -1463 114 -1377 170
rect -1321 114 -1235 170
rect -1179 114 -1093 170
rect -1037 114 -951 170
rect -895 114 -809 170
rect -753 114 -667 170
rect -611 114 -525 170
rect -469 114 -383 170
rect -327 114 -241 170
rect -185 114 -99 170
rect -43 114 43 170
rect 99 114 185 170
rect 241 114 327 170
rect 383 114 469 170
rect 525 114 611 170
rect 667 114 753 170
rect 809 114 895 170
rect 951 114 1037 170
rect 1093 114 1179 170
rect 1235 114 1321 170
rect 1377 114 1463 170
rect 1519 114 1605 170
rect 1661 114 1747 170
rect 1803 114 1889 170
rect 1945 114 2031 170
rect 2087 114 2173 170
rect 2229 114 2315 170
rect 2371 114 2457 170
rect 2513 114 2599 170
rect 2655 114 2741 170
rect 2797 114 2883 170
rect 2939 114 3025 170
rect 3081 114 3167 170
rect 3223 114 3309 170
rect 3365 114 3451 170
rect 3507 114 3593 170
rect 3649 114 3735 170
rect 3791 114 3877 170
rect 3933 114 4019 170
rect 4075 114 4161 170
rect 4217 114 4303 170
rect 4359 114 4445 170
rect 4501 114 4587 170
rect 4643 114 4729 170
rect 4785 114 4871 170
rect 4927 114 5013 170
rect 5069 114 5155 170
rect 5211 114 5297 170
rect 5353 114 5439 170
rect 5495 114 5581 170
rect 5637 114 5723 170
rect 5779 114 5865 170
rect 5921 114 6007 170
rect 6063 114 6149 170
rect 6205 114 6291 170
rect 6347 114 6433 170
rect 6489 114 6575 170
rect 6631 114 6717 170
rect 6773 114 6859 170
rect 6915 114 7001 170
rect 7057 114 7143 170
rect 7199 114 7285 170
rect 7341 114 7351 170
rect -7351 28 7351 114
rect -7351 -28 -7341 28
rect -7285 -28 -7199 28
rect -7143 -28 -7057 28
rect -7001 -28 -6915 28
rect -6859 -28 -6773 28
rect -6717 -28 -6631 28
rect -6575 -28 -6489 28
rect -6433 -28 -6347 28
rect -6291 -28 -6205 28
rect -6149 -28 -6063 28
rect -6007 -28 -5921 28
rect -5865 -28 -5779 28
rect -5723 -28 -5637 28
rect -5581 -28 -5495 28
rect -5439 -28 -5353 28
rect -5297 -28 -5211 28
rect -5155 -28 -5069 28
rect -5013 -28 -4927 28
rect -4871 -28 -4785 28
rect -4729 -28 -4643 28
rect -4587 -28 -4501 28
rect -4445 -28 -4359 28
rect -4303 -28 -4217 28
rect -4161 -28 -4075 28
rect -4019 -28 -3933 28
rect -3877 -28 -3791 28
rect -3735 -28 -3649 28
rect -3593 -28 -3507 28
rect -3451 -28 -3365 28
rect -3309 -28 -3223 28
rect -3167 -28 -3081 28
rect -3025 -28 -2939 28
rect -2883 -28 -2797 28
rect -2741 -28 -2655 28
rect -2599 -28 -2513 28
rect -2457 -28 -2371 28
rect -2315 -28 -2229 28
rect -2173 -28 -2087 28
rect -2031 -28 -1945 28
rect -1889 -28 -1803 28
rect -1747 -28 -1661 28
rect -1605 -28 -1519 28
rect -1463 -28 -1377 28
rect -1321 -28 -1235 28
rect -1179 -28 -1093 28
rect -1037 -28 -951 28
rect -895 -28 -809 28
rect -753 -28 -667 28
rect -611 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 611 28
rect 667 -28 753 28
rect 809 -28 895 28
rect 951 -28 1037 28
rect 1093 -28 1179 28
rect 1235 -28 1321 28
rect 1377 -28 1463 28
rect 1519 -28 1605 28
rect 1661 -28 1747 28
rect 1803 -28 1889 28
rect 1945 -28 2031 28
rect 2087 -28 2173 28
rect 2229 -28 2315 28
rect 2371 -28 2457 28
rect 2513 -28 2599 28
rect 2655 -28 2741 28
rect 2797 -28 2883 28
rect 2939 -28 3025 28
rect 3081 -28 3167 28
rect 3223 -28 3309 28
rect 3365 -28 3451 28
rect 3507 -28 3593 28
rect 3649 -28 3735 28
rect 3791 -28 3877 28
rect 3933 -28 4019 28
rect 4075 -28 4161 28
rect 4217 -28 4303 28
rect 4359 -28 4445 28
rect 4501 -28 4587 28
rect 4643 -28 4729 28
rect 4785 -28 4871 28
rect 4927 -28 5013 28
rect 5069 -28 5155 28
rect 5211 -28 5297 28
rect 5353 -28 5439 28
rect 5495 -28 5581 28
rect 5637 -28 5723 28
rect 5779 -28 5865 28
rect 5921 -28 6007 28
rect 6063 -28 6149 28
rect 6205 -28 6291 28
rect 6347 -28 6433 28
rect 6489 -28 6575 28
rect 6631 -28 6717 28
rect 6773 -28 6859 28
rect 6915 -28 7001 28
rect 7057 -28 7143 28
rect 7199 -28 7285 28
rect 7341 -28 7351 28
rect -7351 -114 7351 -28
rect -7351 -170 -7341 -114
rect -7285 -170 -7199 -114
rect -7143 -170 -7057 -114
rect -7001 -170 -6915 -114
rect -6859 -170 -6773 -114
rect -6717 -170 -6631 -114
rect -6575 -170 -6489 -114
rect -6433 -170 -6347 -114
rect -6291 -170 -6205 -114
rect -6149 -170 -6063 -114
rect -6007 -170 -5921 -114
rect -5865 -170 -5779 -114
rect -5723 -170 -5637 -114
rect -5581 -170 -5495 -114
rect -5439 -170 -5353 -114
rect -5297 -170 -5211 -114
rect -5155 -170 -5069 -114
rect -5013 -170 -4927 -114
rect -4871 -170 -4785 -114
rect -4729 -170 -4643 -114
rect -4587 -170 -4501 -114
rect -4445 -170 -4359 -114
rect -4303 -170 -4217 -114
rect -4161 -170 -4075 -114
rect -4019 -170 -3933 -114
rect -3877 -170 -3791 -114
rect -3735 -170 -3649 -114
rect -3593 -170 -3507 -114
rect -3451 -170 -3365 -114
rect -3309 -170 -3223 -114
rect -3167 -170 -3081 -114
rect -3025 -170 -2939 -114
rect -2883 -170 -2797 -114
rect -2741 -170 -2655 -114
rect -2599 -170 -2513 -114
rect -2457 -170 -2371 -114
rect -2315 -170 -2229 -114
rect -2173 -170 -2087 -114
rect -2031 -170 -1945 -114
rect -1889 -170 -1803 -114
rect -1747 -170 -1661 -114
rect -1605 -170 -1519 -114
rect -1463 -170 -1377 -114
rect -1321 -170 -1235 -114
rect -1179 -170 -1093 -114
rect -1037 -170 -951 -114
rect -895 -170 -809 -114
rect -753 -170 -667 -114
rect -611 -170 -525 -114
rect -469 -170 -383 -114
rect -327 -170 -241 -114
rect -185 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 185 -114
rect 241 -170 327 -114
rect 383 -170 469 -114
rect 525 -170 611 -114
rect 667 -170 753 -114
rect 809 -170 895 -114
rect 951 -170 1037 -114
rect 1093 -170 1179 -114
rect 1235 -170 1321 -114
rect 1377 -170 1463 -114
rect 1519 -170 1605 -114
rect 1661 -170 1747 -114
rect 1803 -170 1889 -114
rect 1945 -170 2031 -114
rect 2087 -170 2173 -114
rect 2229 -170 2315 -114
rect 2371 -170 2457 -114
rect 2513 -170 2599 -114
rect 2655 -170 2741 -114
rect 2797 -170 2883 -114
rect 2939 -170 3025 -114
rect 3081 -170 3167 -114
rect 3223 -170 3309 -114
rect 3365 -170 3451 -114
rect 3507 -170 3593 -114
rect 3649 -170 3735 -114
rect 3791 -170 3877 -114
rect 3933 -170 4019 -114
rect 4075 -170 4161 -114
rect 4217 -170 4303 -114
rect 4359 -170 4445 -114
rect 4501 -170 4587 -114
rect 4643 -170 4729 -114
rect 4785 -170 4871 -114
rect 4927 -170 5013 -114
rect 5069 -170 5155 -114
rect 5211 -170 5297 -114
rect 5353 -170 5439 -114
rect 5495 -170 5581 -114
rect 5637 -170 5723 -114
rect 5779 -170 5865 -114
rect 5921 -170 6007 -114
rect 6063 -170 6149 -114
rect 6205 -170 6291 -114
rect 6347 -170 6433 -114
rect 6489 -170 6575 -114
rect 6631 -170 6717 -114
rect 6773 -170 6859 -114
rect 6915 -170 7001 -114
rect 7057 -170 7143 -114
rect 7199 -170 7285 -114
rect 7341 -170 7351 -114
rect -7351 -256 7351 -170
rect -7351 -312 -7341 -256
rect -7285 -312 -7199 -256
rect -7143 -312 -7057 -256
rect -7001 -312 -6915 -256
rect -6859 -312 -6773 -256
rect -6717 -312 -6631 -256
rect -6575 -312 -6489 -256
rect -6433 -312 -6347 -256
rect -6291 -312 -6205 -256
rect -6149 -312 -6063 -256
rect -6007 -312 -5921 -256
rect -5865 -312 -5779 -256
rect -5723 -312 -5637 -256
rect -5581 -312 -5495 -256
rect -5439 -312 -5353 -256
rect -5297 -312 -5211 -256
rect -5155 -312 -5069 -256
rect -5013 -312 -4927 -256
rect -4871 -312 -4785 -256
rect -4729 -312 -4643 -256
rect -4587 -312 -4501 -256
rect -4445 -312 -4359 -256
rect -4303 -312 -4217 -256
rect -4161 -312 -4075 -256
rect -4019 -312 -3933 -256
rect -3877 -312 -3791 -256
rect -3735 -312 -3649 -256
rect -3593 -312 -3507 -256
rect -3451 -312 -3365 -256
rect -3309 -312 -3223 -256
rect -3167 -312 -3081 -256
rect -3025 -312 -2939 -256
rect -2883 -312 -2797 -256
rect -2741 -312 -2655 -256
rect -2599 -312 -2513 -256
rect -2457 -312 -2371 -256
rect -2315 -312 -2229 -256
rect -2173 -312 -2087 -256
rect -2031 -312 -1945 -256
rect -1889 -312 -1803 -256
rect -1747 -312 -1661 -256
rect -1605 -312 -1519 -256
rect -1463 -312 -1377 -256
rect -1321 -312 -1235 -256
rect -1179 -312 -1093 -256
rect -1037 -312 -951 -256
rect -895 -312 -809 -256
rect -753 -312 -667 -256
rect -611 -312 -525 -256
rect -469 -312 -383 -256
rect -327 -312 -241 -256
rect -185 -312 -99 -256
rect -43 -312 43 -256
rect 99 -312 185 -256
rect 241 -312 327 -256
rect 383 -312 469 -256
rect 525 -312 611 -256
rect 667 -312 753 -256
rect 809 -312 895 -256
rect 951 -312 1037 -256
rect 1093 -312 1179 -256
rect 1235 -312 1321 -256
rect 1377 -312 1463 -256
rect 1519 -312 1605 -256
rect 1661 -312 1747 -256
rect 1803 -312 1889 -256
rect 1945 -312 2031 -256
rect 2087 -312 2173 -256
rect 2229 -312 2315 -256
rect 2371 -312 2457 -256
rect 2513 -312 2599 -256
rect 2655 -312 2741 -256
rect 2797 -312 2883 -256
rect 2939 -312 3025 -256
rect 3081 -312 3167 -256
rect 3223 -312 3309 -256
rect 3365 -312 3451 -256
rect 3507 -312 3593 -256
rect 3649 -312 3735 -256
rect 3791 -312 3877 -256
rect 3933 -312 4019 -256
rect 4075 -312 4161 -256
rect 4217 -312 4303 -256
rect 4359 -312 4445 -256
rect 4501 -312 4587 -256
rect 4643 -312 4729 -256
rect 4785 -312 4871 -256
rect 4927 -312 5013 -256
rect 5069 -312 5155 -256
rect 5211 -312 5297 -256
rect 5353 -312 5439 -256
rect 5495 -312 5581 -256
rect 5637 -312 5723 -256
rect 5779 -312 5865 -256
rect 5921 -312 6007 -256
rect 6063 -312 6149 -256
rect 6205 -312 6291 -256
rect 6347 -312 6433 -256
rect 6489 -312 6575 -256
rect 6631 -312 6717 -256
rect 6773 -312 6859 -256
rect 6915 -312 7001 -256
rect 7057 -312 7143 -256
rect 7199 -312 7285 -256
rect 7341 -312 7351 -256
rect -7351 -398 7351 -312
rect -7351 -454 -7341 -398
rect -7285 -454 -7199 -398
rect -7143 -454 -7057 -398
rect -7001 -454 -6915 -398
rect -6859 -454 -6773 -398
rect -6717 -454 -6631 -398
rect -6575 -454 -6489 -398
rect -6433 -454 -6347 -398
rect -6291 -454 -6205 -398
rect -6149 -454 -6063 -398
rect -6007 -454 -5921 -398
rect -5865 -454 -5779 -398
rect -5723 -454 -5637 -398
rect -5581 -454 -5495 -398
rect -5439 -454 -5353 -398
rect -5297 -454 -5211 -398
rect -5155 -454 -5069 -398
rect -5013 -454 -4927 -398
rect -4871 -454 -4785 -398
rect -4729 -454 -4643 -398
rect -4587 -454 -4501 -398
rect -4445 -454 -4359 -398
rect -4303 -454 -4217 -398
rect -4161 -454 -4075 -398
rect -4019 -454 -3933 -398
rect -3877 -454 -3791 -398
rect -3735 -454 -3649 -398
rect -3593 -454 -3507 -398
rect -3451 -454 -3365 -398
rect -3309 -454 -3223 -398
rect -3167 -454 -3081 -398
rect -3025 -454 -2939 -398
rect -2883 -454 -2797 -398
rect -2741 -454 -2655 -398
rect -2599 -454 -2513 -398
rect -2457 -454 -2371 -398
rect -2315 -454 -2229 -398
rect -2173 -454 -2087 -398
rect -2031 -454 -1945 -398
rect -1889 -454 -1803 -398
rect -1747 -454 -1661 -398
rect -1605 -454 -1519 -398
rect -1463 -454 -1377 -398
rect -1321 -454 -1235 -398
rect -1179 -454 -1093 -398
rect -1037 -454 -951 -398
rect -895 -454 -809 -398
rect -753 -454 -667 -398
rect -611 -454 -525 -398
rect -469 -454 -383 -398
rect -327 -454 -241 -398
rect -185 -454 -99 -398
rect -43 -454 43 -398
rect 99 -454 185 -398
rect 241 -454 327 -398
rect 383 -454 469 -398
rect 525 -454 611 -398
rect 667 -454 753 -398
rect 809 -454 895 -398
rect 951 -454 1037 -398
rect 1093 -454 1179 -398
rect 1235 -454 1321 -398
rect 1377 -454 1463 -398
rect 1519 -454 1605 -398
rect 1661 -454 1747 -398
rect 1803 -454 1889 -398
rect 1945 -454 2031 -398
rect 2087 -454 2173 -398
rect 2229 -454 2315 -398
rect 2371 -454 2457 -398
rect 2513 -454 2599 -398
rect 2655 -454 2741 -398
rect 2797 -454 2883 -398
rect 2939 -454 3025 -398
rect 3081 -454 3167 -398
rect 3223 -454 3309 -398
rect 3365 -454 3451 -398
rect 3507 -454 3593 -398
rect 3649 -454 3735 -398
rect 3791 -454 3877 -398
rect 3933 -454 4019 -398
rect 4075 -454 4161 -398
rect 4217 -454 4303 -398
rect 4359 -454 4445 -398
rect 4501 -454 4587 -398
rect 4643 -454 4729 -398
rect 4785 -454 4871 -398
rect 4927 -454 5013 -398
rect 5069 -454 5155 -398
rect 5211 -454 5297 -398
rect 5353 -454 5439 -398
rect 5495 -454 5581 -398
rect 5637 -454 5723 -398
rect 5779 -454 5865 -398
rect 5921 -454 6007 -398
rect 6063 -454 6149 -398
rect 6205 -454 6291 -398
rect 6347 -454 6433 -398
rect 6489 -454 6575 -398
rect 6631 -454 6717 -398
rect 6773 -454 6859 -398
rect 6915 -454 7001 -398
rect 7057 -454 7143 -398
rect 7199 -454 7285 -398
rect 7341 -454 7351 -398
rect -7351 -540 7351 -454
rect -7351 -596 -7341 -540
rect -7285 -596 -7199 -540
rect -7143 -596 -7057 -540
rect -7001 -596 -6915 -540
rect -6859 -596 -6773 -540
rect -6717 -596 -6631 -540
rect -6575 -596 -6489 -540
rect -6433 -596 -6347 -540
rect -6291 -596 -6205 -540
rect -6149 -596 -6063 -540
rect -6007 -596 -5921 -540
rect -5865 -596 -5779 -540
rect -5723 -596 -5637 -540
rect -5581 -596 -5495 -540
rect -5439 -596 -5353 -540
rect -5297 -596 -5211 -540
rect -5155 -596 -5069 -540
rect -5013 -596 -4927 -540
rect -4871 -596 -4785 -540
rect -4729 -596 -4643 -540
rect -4587 -596 -4501 -540
rect -4445 -596 -4359 -540
rect -4303 -596 -4217 -540
rect -4161 -596 -4075 -540
rect -4019 -596 -3933 -540
rect -3877 -596 -3791 -540
rect -3735 -596 -3649 -540
rect -3593 -596 -3507 -540
rect -3451 -596 -3365 -540
rect -3309 -596 -3223 -540
rect -3167 -596 -3081 -540
rect -3025 -596 -2939 -540
rect -2883 -596 -2797 -540
rect -2741 -596 -2655 -540
rect -2599 -596 -2513 -540
rect -2457 -596 -2371 -540
rect -2315 -596 -2229 -540
rect -2173 -596 -2087 -540
rect -2031 -596 -1945 -540
rect -1889 -596 -1803 -540
rect -1747 -596 -1661 -540
rect -1605 -596 -1519 -540
rect -1463 -596 -1377 -540
rect -1321 -596 -1235 -540
rect -1179 -596 -1093 -540
rect -1037 -596 -951 -540
rect -895 -596 -809 -540
rect -753 -596 -667 -540
rect -611 -596 -525 -540
rect -469 -596 -383 -540
rect -327 -596 -241 -540
rect -185 -596 -99 -540
rect -43 -596 43 -540
rect 99 -596 185 -540
rect 241 -596 327 -540
rect 383 -596 469 -540
rect 525 -596 611 -540
rect 667 -596 753 -540
rect 809 -596 895 -540
rect 951 -596 1037 -540
rect 1093 -596 1179 -540
rect 1235 -596 1321 -540
rect 1377 -596 1463 -540
rect 1519 -596 1605 -540
rect 1661 -596 1747 -540
rect 1803 -596 1889 -540
rect 1945 -596 2031 -540
rect 2087 -596 2173 -540
rect 2229 -596 2315 -540
rect 2371 -596 2457 -540
rect 2513 -596 2599 -540
rect 2655 -596 2741 -540
rect 2797 -596 2883 -540
rect 2939 -596 3025 -540
rect 3081 -596 3167 -540
rect 3223 -596 3309 -540
rect 3365 -596 3451 -540
rect 3507 -596 3593 -540
rect 3649 -596 3735 -540
rect 3791 -596 3877 -540
rect 3933 -596 4019 -540
rect 4075 -596 4161 -540
rect 4217 -596 4303 -540
rect 4359 -596 4445 -540
rect 4501 -596 4587 -540
rect 4643 -596 4729 -540
rect 4785 -596 4871 -540
rect 4927 -596 5013 -540
rect 5069 -596 5155 -540
rect 5211 -596 5297 -540
rect 5353 -596 5439 -540
rect 5495 -596 5581 -540
rect 5637 -596 5723 -540
rect 5779 -596 5865 -540
rect 5921 -596 6007 -540
rect 6063 -596 6149 -540
rect 6205 -596 6291 -540
rect 6347 -596 6433 -540
rect 6489 -596 6575 -540
rect 6631 -596 6717 -540
rect 6773 -596 6859 -540
rect 6915 -596 7001 -540
rect 7057 -596 7143 -540
rect 7199 -596 7285 -540
rect 7341 -596 7351 -540
rect -7351 -606 7351 -596
<< end >>
