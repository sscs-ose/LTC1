* NGSPICE file created from gf_inv_mag_flat.ext - technology: gf180mcuC

.subckt gf_inv_mag_flat VSS OUT IN VDD
X0 VDD IN.t0 gf_inv_mag_1.IN VDD.t7 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X1 OUT gf_inv_mag_1.IN VDD.t19 VDD.t18 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X2 gf_inv_mag_1.IN IN.t1 VSS.t9 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X3 VSS IN.t2 gf_inv_mag_1.IN VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X4 VSS gf_inv_mag_1.IN OUT.t5 VSS.t17 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X5 gf_inv_mag_1.IN IN.t3 VSS.t4 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X6 gf_inv_mag_1.IN IN.t4 VDD.t6 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X7 VDD gf_inv_mag_1.IN OUT.t2 VDD.t15 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X8 OUT gf_inv_mag_1.IN VSS.t16 VSS.t15 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X9 VDD IN.t5 gf_inv_mag_1.IN VDD.t2 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X10 VSS gf_inv_mag_1.IN OUT.t4 VSS.t12 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X11 gf_inv_mag_1.IN IN.t6 VDD.t1 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X12 OUT gf_inv_mag_1.IN VSS.t11 VSS.t10 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X13 OUT gf_inv_mag_1.IN VDD.t14 VDD.t13 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X14 VDD gf_inv_mag_1.IN OUT.t0 VDD.t10 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X15 VSS IN.t7 gf_inv_mag_1.IN VSS.t0 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
R0 IN.n2 IN.t2 25.8422
R1 IN.n0 IN.t7 25.8105
R2 IN.n1 IN.t1 25.809
R3 IN.n0 IN.t0 25.6004
R4 IN.n1 IN.t4 25.6004
R5 IN.n2 IN.t5 25.5672
R6 IN.n3 IN.t3 24.6435
R7 IN.n4 IN.t6 23.8188
R8 IN.n3 IN.n2 11.9051
R9 IN.n1 IN.n0 11.7928
R10 IN.n2 IN.n1 11.6805
R11 IN IN.n4 4.186
R12 IN.n4 IN.n3 0.338463
R13 VDD.t7 VDD.t18 609.678
R14 VDD.t13 VDD.t15 280.646
R15 VDD.t18 VDD.t10 280.646
R16 VDD.t5 VDD.t7 280.646
R17 VDD.t2 VDD.t0 280.646
R18 VDD.n8 VDD.t13 158.065
R19 VDD.n9 VDD.t5 158.065
R20 VDD.t10 VDD.n8 122.582
R21 VDD.n9 VDD.t2 122.582
R22 VDD.n3 VDD.n2 6.57811
R23 VDD VDD.t1 6.57171
R24 VDD.n12 VDD.n5 6.4598
R25 VDD.n13 VDD.t19 6.4598
R26 VDD.n10 VDD.n9 6.3005
R27 VDD.n8 VDD.n4 6.3005
R28 VDD.n7 VDD.t6 3.6405
R29 VDD.n7 VDD.n6 3.6405
R30 VDD.n1 VDD.t14 3.6405
R31 VDD.n1 VDD.n0 3.6405
R32 VDD.n11 VDD.n7 2.8198
R33 VDD.n3 VDD.n1 2.8198
R34 VDD VDD.n13 0.112058
R35 VDD VDD.n11 0.104691
R36 VDD.n13 VDD.n12 0.0688333
R37 VDD.n12 VDD 0.0138333
R38 VDD.n11 VDD.n10 0.00353371
R39 VDD.n4 VDD.n3 0.00353371
R40 VDD.n10 VDD 0.00151124
R41 VDD VDD.n4 0.00151124
R42 OUT.n1 OUT.t0 3.6405
R43 OUT.n1 OUT.n0 3.6405
R44 OUT.n6 OUT.t2 3.6405
R45 OUT.n6 OUT.n5 3.6405
R46 OUT.n9 OUT.n8 3.48732
R47 OUT.n4 OUT.n3 3.47267
R48 OUT.n9 OUT.n6 2.9305
R49 OUT.n4 OUT.n1 2.91615
R50 OUT.n3 OUT.t4 1.6385
R51 OUT.n3 OUT.n2 1.6385
R52 OUT.n8 OUT.t5 1.6385
R53 OUT.n8 OUT.n7 1.6385
R54 OUT.n9 OUT.n4 0.384406
R55 OUT OUT.n9 0.294406
R56 VSS.t0 VSS.t10 1814.62
R57 VSS.t15 VSS.t17 835.303
R58 VSS.t10 VSS.t12 835.303
R59 VSS.t8 VSS.t0 835.303
R60 VSS.t5 VSS.t3 835.303
R61 VSS.n8 VSS.t15 686.485
R62 VSS.n9 VSS.t8 686.485
R63 VSS.t12 VSS.n8 148.819
R64 VSS.n9 VSS.t5 148.819
R65 VSS.n3 VSS.n2 5.20098
R66 VSS.n10 VSS.n9 5.2005
R67 VSS.n8 VSS.n4 5.2005
R68 VSS VSS.t4 5.15186
R69 VSS.n12 VSS.n5 5.04745
R70 VSS.n13 VSS.t11 5.02656
R71 VSS.n3 VSS.n1 3.37758
R72 VSS.n11 VSS.n7 3.37758
R73 VSS.n1 VSS.t16 1.6385
R74 VSS.n1 VSS.n0 1.6385
R75 VSS.n7 VSS.t9 1.6385
R76 VSS.n7 VSS.n6 1.6385
R77 VSS.n12 VSS.n11 0.154029
R78 VSS VSS.n13 0.125794
R79 VSS.n13 VSS 0.0702059
R80 VSS.n4 VSS.n3 0.0243235
R81 VSS.n11 VSS.n10 0.0243235
R82 VSS VSS.n12 0.0207941
R83 VSS VSS.n4 0.00491176
R84 VSS.n10 VSS 0.00491176
C0 gf_inv_mag_1.IN IN 0.376f
C1 OUT IN 0.0023f
C2 OUT gf_inv_mag_1.IN 0.381f
C3 VDD IN 0.604f
C4 gf_inv_mag_1.IN VDD 0.991f
C5 OUT VDD 0.397f
C6 OUT VSS 0.693f
C7 gf_inv_mag_1.IN VSS 1.84f
C8 IN VSS 1.27f
C9 VDD VSS 3.89f
.ends

