magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2144 -2083 15504 16940
<< metal1 >>
rect 12354 10602 13432 10703
rect 10095 7691 10347 7871
rect 9570 6237 10171 6313
rect 12737 6306 13403 6393
rect 9726 6101 10351 6177
rect 8310 5571 8815 5639
rect 13168 4882 13378 5374
rect 7991 4446 9118 4522
rect 12910 4326 13432 4439
rect 6733 4202 7000 4270
rect 7841 3169 9118 3245
rect 377 2969 12754 3045
rect 3329 2832 6238 2908
rect 8162 2833 10072 2909
rect 1784 2697 9490 2773
rect 9726 2697 10142 2773
rect 11457 2718 12859 2794
rect -144 2561 7619 2637
rect 9570 2561 11482 2637
rect 73 1592 1858 1956
rect 73 683 2698 1056
<< metal2 >>
rect 9906 9171 10977 9247
rect 9906 7712 9982 9171
rect 9414 7636 9982 7712
rect 6579 5511 6779 6291
rect 6579 5351 7000 5511
rect 2295 3129 2371 4152
rect 3045 3344 3640 3348
rect 2969 3272 3640 3344
rect 2295 3053 3237 3129
rect -144 1415 -68 2637
rect -144 1235 317 1415
rect -144 422 -68 1235
rect 377 422 453 3045
rect 3161 2832 3237 3053
rect 1784 2262 1860 2773
rect 1499 2186 1860 2262
rect 3564 1571 3640 3272
rect 6162 1958 6238 2891
rect 4334 1571 4410 1958
rect 3564 1495 4410 1571
rect 2953 1362 3029 1485
rect 1499 1286 3029 1362
rect 7543 1305 7619 2637
rect 8162 1305 8238 2909
rect 9414 2697 9490 7636
rect 9570 2561 9646 6313
rect 10095 6237 10171 7871
rect 9726 2697 9802 6177
rect 10275 6101 10351 7381
rect 11245 5705 11321 10865
rect 12164 7970 12240 9649
rect 9892 5629 11321 5705
rect 11457 7894 12240 7970
rect 9892 2833 9948 5629
rect 10066 1958 10142 2773
rect 11457 2718 11513 7894
rect 12136 3237 12316 6526
rect 13356 6384 13432 10673
rect 12736 3045 12812 6306
rect 12694 2969 12812 3045
rect 11406 1958 11482 2637
rect 12783 1305 12859 2794
use comp018green_in_cms_smt  comp018green_in_cms_smt_0
timestamp 1713338890
transform 1 0 1532 0 1 3158
box -1470 -83 6872 2575
use comp018green_in_drv  comp018green_in_drv_0
timestamp 1713338890
transform 1 0 8900 0 1 3158
box -496 -83 4434 2575
use comp018green_in_logic_pupd  comp018green_in_logic_pupd_0
timestamp 1713338890
transform -1 0 13932 0 1 9724
box 428 -3277 3307 2142
use comp018green_in_pupd  comp018green_in_pupd_0
timestamp 1713338890
transform 0 -1 2979 -1 0 14857
box -83 -7815 8992 3035
use comp018green_sigbuf  comp018green_sigbuf_0
timestamp 1713338890
transform 1 0 2619 0 -1 2492
box -83 -83 2795 2575
use comp018green_sigbuf  comp018green_sigbuf_1
timestamp 1713338890
transform -1 0 7953 0 -1 2492
box -83 -83 2795 2575
use comp018green_sigbuf  comp018green_sigbuf_2
timestamp 1713338890
transform 1 0 7863 0 -1 2492
box -83 -83 2795 2575
use comp018green_sigbuf  comp018green_sigbuf_3
timestamp 1713338890
transform -1 0 13197 0 -1 2492
box -83 -83 2795 2575
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_0
timestamp 1713338890
transform 1 0 1589 0 1 1324
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_1
timestamp 1713338890
transform 0 1 279 -1 0 1325
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_2
timestamp 1713338890
transform 1 0 1874 0 1 2735
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_3
timestamp 1713338890
transform 1 0 340 0 1 2224
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_4
timestamp 1713338890
transform 1 0 -54 0 1 2599
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_5
timestamp 1713338890
transform 1 0 1589 0 1 2224
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_6
timestamp 1713338890
transform 0 -1 415 1 0 3059
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_7
timestamp 1713338890
transform 1 0 3059 0 1 3321
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_8
timestamp 1713338890
transform 1 0 3261 0 1 2870
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_9
timestamp 1713338890
transform 1 0 6197 0 1 2870
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_10
timestamp 1713338890
transform 1 0 9982 0 1 2871
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_11
timestamp 1713338890
transform 1 0 10052 0 1 2735
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_12
timestamp 1713338890
transform 1 0 8148 0 1 2871
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_13
timestamp 1713338890
transform 1 0 7529 0 1 2599
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_14
timestamp 1713338890
transform 0 1 9452 -1 0 2683
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_15
timestamp 1713338890
transform 1 0 12627 0 1 3007
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_16
timestamp 1713338890
transform 1 0 11547 0 1 2756
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_17
timestamp 1713338890
transform 1 0 11392 0 1 2599
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_18
timestamp 1713338890
transform 1 0 12769 0 1 2756
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_19
timestamp 1713338890
transform 1 0 12226 0 1 3199
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_20
timestamp 1713338890
transform 1 0 6910 0 1 4240
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_21
timestamp 1713338890
transform 1 0 10081 0 1 6275
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_22
timestamp 1713338890
transform 1 0 9660 0 1 6275
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_23
timestamp 1713338890
transform 1 0 9816 0 1 6139
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_24
timestamp 1713338890
transform 1 0 10261 0 1 6139
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_25
timestamp 1713338890
transform 1 0 12226 0 1 6488
box -90 -38 90 38
use M2_M1_CDNS_69033583165523  M2_M1_CDNS_69033583165523_26
timestamp 1713338890
transform 1 0 11184 0 1 10827
box -90 -38 90 38
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_0
timestamp 1713338890
transform 1 0 2991 0 1 1395
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_1
timestamp 1713338890
transform 1 0 4372 0 1 2048
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_2
timestamp 1713338890
transform 1 0 6200 0 1 2048
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_3
timestamp 1713338890
transform 1 0 8200 0 1 1395
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_4
timestamp 1713338890
transform 1 0 7581 0 1 1395
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_5
timestamp 1713338890
transform 1 0 9608 0 1 2651
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_6
timestamp 1713338890
transform 1 0 10104 0 1 2048
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_7
timestamp 1713338890
transform 0 -1 9816 1 0 2735
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_8
timestamp 1713338890
transform 1 0 11444 0 1 2048
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_9
timestamp 1713338890
transform 1 0 12821 0 1 1395
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_10
timestamp 1713338890
transform 1 0 13394 0 1 4380
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_11
timestamp 1713338890
transform 1 0 10313 0 1 7291
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_12
timestamp 1713338890
transform 1 0 13394 0 1 6303
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_13
timestamp 1713338890
transform 1 0 12774 0 1 6303
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_14
timestamp 1713338890
transform 1 0 12202 0 1 9734
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_15
timestamp 1713338890
transform 1 0 13394 0 1 10613
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_16
timestamp 1713338890
transform 1 0 10133 0 1 7781
box -38 -90 38 90
use M2_M1_CDNS_69033583165614  M2_M1_CDNS_69033583165614_0
timestamp 1713338890
transform 1 0 10065 0 1 3942
box -38 -246 38 246
use M2_M1_CDNS_69033583165614  M2_M1_CDNS_69033583165614_1
timestamp 1713338890
transform 1 0 10065 0 1 5128
box -38 -246 38 246
use M2_M1_CDNS_69033583165614  M2_M1_CDNS_69033583165614_2
timestamp 1713338890
transform 1 0 13414 0 1 5128
box -38 -246 38 246
use M3_M2_CDNS_69033583165577  M3_M2_CDNS_69033583165577_0
timestamp 1713338890
transform 1 0 12226 0 1 3320
box -90 -38 90 38
use M3_M2_CDNS_69033583165615  M3_M2_CDNS_69033583165615_0
timestamp 1713338890
transform 1 0 10065 0 1 5128
box -38 -246 38 246
use M3_M2_CDNS_69033583165615  M3_M2_CDNS_69033583165615_1
timestamp 1713338890
transform 1 0 10065 0 1 3942
box -38 -246 38 246
use M3_M2_CDNS_69033583165615  M3_M2_CDNS_69033583165615_2
timestamp 1713338890
transform 1 0 13414 0 1 5128
box -38 -246 38 246
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_0
timestamp 1713338890
transform 1 0 1490 0 1 1224
box -216 -216 416 416
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_1
timestamp 1713338890
transform 1 0 241 0 1 1224
box -216 -216 416 416
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_2
timestamp 1713338890
transform 1 0 241 0 1 2124
box -216 -216 416 416
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_3
timestamp 1713338890
transform 1 0 1490 0 1 2124
box -216 -216 416 416
<< labels >>
rlabel metal1 s 11686 5601 11686 5601 4 VDD
port 1 nsew
rlabel metal2 s 414 522 414 522 4 PU
port 2 nsew
rlabel metal2 s 1822 2409 1822 2409 4 PD
port 3 nsew
rlabel metal2 s -107 526 -107 526 4 CS
port 4 nsew
rlabel metal2 s 2128 1324 2128 1324 4 IE
port 5 nsew
rlabel metal2 s 6679 6191 6679 6191 4 PAD
port 6 nsew
<< end >>
