magic
tech gf180mcuC
magscale 1 10
timestamp 1693073856
<< nwell >>
rect -264 -11682 264 11682
<< nsubdiff >>
rect -240 11586 240 11658
rect -240 -11586 -168 11586
rect 168 -11586 240 11586
rect -240 -11658 240 -11586
<< polysilicon >>
rect -80 11485 80 11498
rect -80 11439 -67 11485
rect 67 11439 80 11485
rect -80 11396 80 11439
rect -80 9351 80 9394
rect -80 9305 -67 9351
rect 67 9305 80 9351
rect -80 9292 80 9305
rect -80 9175 80 9188
rect -80 9129 -67 9175
rect 67 9129 80 9175
rect -80 9086 80 9129
rect -80 7041 80 7084
rect -80 6995 -67 7041
rect 67 6995 80 7041
rect -80 6982 80 6995
rect -80 6865 80 6878
rect -80 6819 -67 6865
rect 67 6819 80 6865
rect -80 6776 80 6819
rect -80 4731 80 4774
rect -80 4685 -67 4731
rect 67 4685 80 4731
rect -80 4672 80 4685
rect -80 4555 80 4568
rect -80 4509 -67 4555
rect 67 4509 80 4555
rect -80 4466 80 4509
rect -80 2421 80 2464
rect -80 2375 -67 2421
rect 67 2375 80 2421
rect -80 2362 80 2375
rect -80 2245 80 2258
rect -80 2199 -67 2245
rect 67 2199 80 2245
rect -80 2156 80 2199
rect -80 111 80 154
rect -80 65 -67 111
rect 67 65 80 111
rect -80 52 80 65
rect -80 -65 80 -52
rect -80 -111 -67 -65
rect 67 -111 80 -65
rect -80 -154 80 -111
rect -80 -2199 80 -2156
rect -80 -2245 -67 -2199
rect 67 -2245 80 -2199
rect -80 -2258 80 -2245
rect -80 -2375 80 -2362
rect -80 -2421 -67 -2375
rect 67 -2421 80 -2375
rect -80 -2464 80 -2421
rect -80 -4509 80 -4466
rect -80 -4555 -67 -4509
rect 67 -4555 80 -4509
rect -80 -4568 80 -4555
rect -80 -4685 80 -4672
rect -80 -4731 -67 -4685
rect 67 -4731 80 -4685
rect -80 -4774 80 -4731
rect -80 -6819 80 -6776
rect -80 -6865 -67 -6819
rect 67 -6865 80 -6819
rect -80 -6878 80 -6865
rect -80 -6995 80 -6982
rect -80 -7041 -67 -6995
rect 67 -7041 80 -6995
rect -80 -7084 80 -7041
rect -80 -9129 80 -9086
rect -80 -9175 -67 -9129
rect 67 -9175 80 -9129
rect -80 -9188 80 -9175
rect -80 -9305 80 -9292
rect -80 -9351 -67 -9305
rect 67 -9351 80 -9305
rect -80 -9394 80 -9351
rect -80 -11439 80 -11396
rect -80 -11485 -67 -11439
rect 67 -11485 80 -11439
rect -80 -11498 80 -11485
<< polycontact >>
rect -67 11439 67 11485
rect -67 9305 67 9351
rect -67 9129 67 9175
rect -67 6995 67 7041
rect -67 6819 67 6865
rect -67 4685 67 4731
rect -67 4509 67 4555
rect -67 2375 67 2421
rect -67 2199 67 2245
rect -67 65 67 111
rect -67 -111 67 -65
rect -67 -2245 67 -2199
rect -67 -2421 67 -2375
rect -67 -4555 67 -4509
rect -67 -4731 67 -4685
rect -67 -6865 67 -6819
rect -67 -7041 67 -6995
rect -67 -9175 67 -9129
rect -67 -9351 67 -9305
rect -67 -11485 67 -11439
<< ppolyres >>
rect -80 9394 80 11396
rect -80 7084 80 9086
rect -80 4774 80 6776
rect -80 2464 80 4466
rect -80 154 80 2156
rect -80 -2156 80 -154
rect -80 -4466 80 -2464
rect -80 -6776 80 -4774
rect -80 -9086 80 -7084
rect -80 -11396 80 -9394
<< metal1 >>
rect -78 11439 -67 11485
rect 67 11439 78 11485
rect -78 9305 -67 9351
rect 67 9305 78 9351
rect -78 9129 -67 9175
rect 67 9129 78 9175
rect -78 6995 -67 7041
rect 67 6995 78 7041
rect -78 6819 -67 6865
rect 67 6819 78 6865
rect -78 4685 -67 4731
rect 67 4685 78 4731
rect -78 4509 -67 4555
rect 67 4509 78 4555
rect -78 2375 -67 2421
rect 67 2375 78 2421
rect -78 2199 -67 2245
rect 67 2199 78 2245
rect -78 65 -67 111
rect 67 65 78 111
rect -78 -111 -67 -65
rect 67 -111 78 -65
rect -78 -2245 -67 -2199
rect 67 -2245 78 -2199
rect -78 -2421 -67 -2375
rect 67 -2421 78 -2375
rect -78 -4555 -67 -4509
rect 67 -4555 78 -4509
rect -78 -4731 -67 -4685
rect 67 -4731 78 -4685
rect -78 -6865 -67 -6819
rect 67 -6865 78 -6819
rect -78 -7041 -67 -6995
rect 67 -7041 78 -6995
rect -78 -9175 -67 -9129
rect 67 -9175 78 -9129
rect -78 -9351 -67 -9305
rect 67 -9351 78 -9305
rect -78 -11485 -67 -11439
rect 67 -11485 78 -11439
<< properties >>
string FIXED_BBOX -204 -11622 204 11622
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 10.01 m 10 nx 1 wmin 0.80 lmin 1.00 rho 315 val 4.319k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
