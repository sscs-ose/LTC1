magic
tech gf180mcuC
magscale 1 10
timestamp 1692615943
<< nwell >>
rect -554 -1534 554 1534
<< pmos >>
rect -380 804 -268 1404
rect -164 804 -52 1404
rect 52 804 164 1404
rect 268 804 380 1404
rect -380 68 -268 668
rect -164 68 -52 668
rect 52 68 164 668
rect 268 68 380 668
rect -380 -668 -268 -68
rect -164 -668 -52 -68
rect 52 -668 164 -68
rect 268 -668 380 -68
rect -380 -1404 -268 -804
rect -164 -1404 -52 -804
rect 52 -1404 164 -804
rect 268 -1404 380 -804
<< pdiff >>
rect -468 1391 -380 1404
rect -468 817 -455 1391
rect -409 817 -380 1391
rect -468 804 -380 817
rect -268 1391 -164 1404
rect -268 817 -239 1391
rect -193 817 -164 1391
rect -268 804 -164 817
rect -52 1391 52 1404
rect -52 817 -23 1391
rect 23 817 52 1391
rect -52 804 52 817
rect 164 1391 268 1404
rect 164 817 193 1391
rect 239 817 268 1391
rect 164 804 268 817
rect 380 1391 468 1404
rect 380 817 409 1391
rect 455 817 468 1391
rect 380 804 468 817
rect -468 655 -380 668
rect -468 81 -455 655
rect -409 81 -380 655
rect -468 68 -380 81
rect -268 655 -164 668
rect -268 81 -239 655
rect -193 81 -164 655
rect -268 68 -164 81
rect -52 655 52 668
rect -52 81 -23 655
rect 23 81 52 655
rect -52 68 52 81
rect 164 655 268 668
rect 164 81 193 655
rect 239 81 268 655
rect 164 68 268 81
rect 380 655 468 668
rect 380 81 409 655
rect 455 81 468 655
rect 380 68 468 81
rect -468 -81 -380 -68
rect -468 -655 -455 -81
rect -409 -655 -380 -81
rect -468 -668 -380 -655
rect -268 -81 -164 -68
rect -268 -655 -239 -81
rect -193 -655 -164 -81
rect -268 -668 -164 -655
rect -52 -81 52 -68
rect -52 -655 -23 -81
rect 23 -655 52 -81
rect -52 -668 52 -655
rect 164 -81 268 -68
rect 164 -655 193 -81
rect 239 -655 268 -81
rect 164 -668 268 -655
rect 380 -81 468 -68
rect 380 -655 409 -81
rect 455 -655 468 -81
rect 380 -668 468 -655
rect -468 -817 -380 -804
rect -468 -1391 -455 -817
rect -409 -1391 -380 -817
rect -468 -1404 -380 -1391
rect -268 -817 -164 -804
rect -268 -1391 -239 -817
rect -193 -1391 -164 -817
rect -268 -1404 -164 -1391
rect -52 -817 52 -804
rect -52 -1391 -23 -817
rect 23 -1391 52 -817
rect -52 -1404 52 -1391
rect 164 -817 268 -804
rect 164 -1391 193 -817
rect 239 -1391 268 -817
rect 164 -1404 268 -1391
rect 380 -817 468 -804
rect 380 -1391 409 -817
rect 455 -1391 468 -817
rect 380 -1404 468 -1391
<< pdiffc >>
rect -455 817 -409 1391
rect -239 817 -193 1391
rect -23 817 23 1391
rect 193 817 239 1391
rect 409 817 455 1391
rect -455 81 -409 655
rect -239 81 -193 655
rect -23 81 23 655
rect 193 81 239 655
rect 409 81 455 655
rect -455 -655 -409 -81
rect -239 -655 -193 -81
rect -23 -655 23 -81
rect 193 -655 239 -81
rect 409 -655 455 -81
rect -455 -1391 -409 -817
rect -239 -1391 -193 -817
rect -23 -1391 23 -817
rect 193 -1391 239 -817
rect 409 -1391 455 -817
<< polysilicon >>
rect -380 1404 -268 1448
rect -164 1404 -52 1448
rect 52 1404 164 1448
rect 268 1404 380 1448
rect -380 760 -268 804
rect -164 760 -52 804
rect 52 760 164 804
rect 268 760 380 804
rect -380 668 -268 712
rect -164 668 -52 712
rect 52 668 164 712
rect 268 668 380 712
rect -380 24 -268 68
rect -164 24 -52 68
rect 52 24 164 68
rect 268 24 380 68
rect -380 -68 -268 -24
rect -164 -68 -52 -24
rect 52 -68 164 -24
rect 268 -68 380 -24
rect -380 -712 -268 -668
rect -164 -712 -52 -668
rect 52 -712 164 -668
rect 268 -712 380 -668
rect -380 -804 -268 -760
rect -164 -804 -52 -760
rect 52 -804 164 -760
rect 268 -804 380 -760
rect -380 -1448 -268 -1404
rect -164 -1448 -52 -1404
rect 52 -1448 164 -1404
rect 268 -1448 380 -1404
<< metal1 >>
rect -455 1391 -409 1402
rect -455 806 -409 817
rect -239 1391 -193 1402
rect -239 806 -193 817
rect -23 1391 23 1402
rect -23 806 23 817
rect 193 1391 239 1402
rect 193 806 239 817
rect 409 1391 455 1402
rect 409 806 455 817
rect -455 655 -409 666
rect -455 70 -409 81
rect -239 655 -193 666
rect -239 70 -193 81
rect -23 655 23 666
rect -23 70 23 81
rect 193 655 239 666
rect 193 70 239 81
rect 409 655 455 666
rect 409 70 455 81
rect -455 -81 -409 -70
rect -455 -666 -409 -655
rect -239 -81 -193 -70
rect -239 -666 -193 -655
rect -23 -81 23 -70
rect -23 -666 23 -655
rect 193 -81 239 -70
rect 193 -666 239 -655
rect 409 -81 455 -70
rect 409 -666 455 -655
rect -455 -817 -409 -806
rect -455 -1402 -409 -1391
rect -239 -817 -193 -806
rect -239 -1402 -193 -1391
rect -23 -817 23 -806
rect -23 -1402 23 -1391
rect 193 -817 239 -806
rect 193 -1402 239 -1391
rect 409 -817 455 -806
rect 409 -1402 455 -1391
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 3 l 0.56 m 4 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
