** sch_path: /home/shahid/GF180Projects/CP_PFD_dff_inv_nand_/Xschem/a_mux/pex_analog_mux_test.sch
**.subckt pex_analog_mux_test
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V4 SEL VSS pulse(0 3.3 0 100p 100p 400n 800n)
.save i(v4)
V6 IN2 VSS 1.12
.save i(v6)
V3 IN1 VSS 2.0
.save i(v3)
x1 IN1 VDD VOUT SEL VSS IN2 pex_a2x1mux_mag
**** begin user architecture code


.include pex_a2x1mux_mag.spice
.control
save all
tran 50p 800n
plot v(S)  v(I0)+5 v(I1)+10 v(OUT)+15


**write analog_mux_TB.raw
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
