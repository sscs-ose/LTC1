magic
tech gf180mcuC
magscale 1 10
timestamp 1692187240
<< nwell >>
rect -1344 -1487 1344 1487
<< nsubdiff >>
rect -1320 1391 1320 1463
rect -1320 -1391 -1248 1391
rect 1248 -1391 1320 1391
rect -1320 -1463 1320 -1391
<< polysilicon >>
rect -1160 1290 -1000 1303
rect -1160 1244 -1147 1290
rect -1013 1244 -1000 1290
rect -1160 1200 -1000 1244
rect -1160 -1244 -1000 -1200
rect -1160 -1290 -1147 -1244
rect -1013 -1290 -1000 -1244
rect -1160 -1303 -1000 -1290
rect -920 1290 -760 1303
rect -920 1244 -907 1290
rect -773 1244 -760 1290
rect -920 1200 -760 1244
rect -920 -1244 -760 -1200
rect -920 -1290 -907 -1244
rect -773 -1290 -760 -1244
rect -920 -1303 -760 -1290
rect -680 1290 -520 1303
rect -680 1244 -667 1290
rect -533 1244 -520 1290
rect -680 1200 -520 1244
rect -680 -1244 -520 -1200
rect -680 -1290 -667 -1244
rect -533 -1290 -520 -1244
rect -680 -1303 -520 -1290
rect -440 1290 -280 1303
rect -440 1244 -427 1290
rect -293 1244 -280 1290
rect -440 1200 -280 1244
rect -440 -1244 -280 -1200
rect -440 -1290 -427 -1244
rect -293 -1290 -280 -1244
rect -440 -1303 -280 -1290
rect -200 1290 -40 1303
rect -200 1244 -187 1290
rect -53 1244 -40 1290
rect -200 1200 -40 1244
rect -200 -1244 -40 -1200
rect -200 -1290 -187 -1244
rect -53 -1290 -40 -1244
rect -200 -1303 -40 -1290
rect 40 1290 200 1303
rect 40 1244 53 1290
rect 187 1244 200 1290
rect 40 1200 200 1244
rect 40 -1244 200 -1200
rect 40 -1290 53 -1244
rect 187 -1290 200 -1244
rect 40 -1303 200 -1290
rect 280 1290 440 1303
rect 280 1244 293 1290
rect 427 1244 440 1290
rect 280 1200 440 1244
rect 280 -1244 440 -1200
rect 280 -1290 293 -1244
rect 427 -1290 440 -1244
rect 280 -1303 440 -1290
rect 520 1290 680 1303
rect 520 1244 533 1290
rect 667 1244 680 1290
rect 520 1200 680 1244
rect 520 -1244 680 -1200
rect 520 -1290 533 -1244
rect 667 -1290 680 -1244
rect 520 -1303 680 -1290
rect 760 1290 920 1303
rect 760 1244 773 1290
rect 907 1244 920 1290
rect 760 1200 920 1244
rect 760 -1244 920 -1200
rect 760 -1290 773 -1244
rect 907 -1290 920 -1244
rect 760 -1303 920 -1290
rect 1000 1290 1160 1303
rect 1000 1244 1013 1290
rect 1147 1244 1160 1290
rect 1000 1200 1160 1244
rect 1000 -1244 1160 -1200
rect 1000 -1290 1013 -1244
rect 1147 -1290 1160 -1244
rect 1000 -1303 1160 -1290
<< polycontact >>
rect -1147 1244 -1013 1290
rect -1147 -1290 -1013 -1244
rect -907 1244 -773 1290
rect -907 -1290 -773 -1244
rect -667 1244 -533 1290
rect -667 -1290 -533 -1244
rect -427 1244 -293 1290
rect -427 -1290 -293 -1244
rect -187 1244 -53 1290
rect -187 -1290 -53 -1244
rect 53 1244 187 1290
rect 53 -1290 187 -1244
rect 293 1244 427 1290
rect 293 -1290 427 -1244
rect 533 1244 667 1290
rect 533 -1290 667 -1244
rect 773 1244 907 1290
rect 773 -1290 907 -1244
rect 1013 1244 1147 1290
rect 1013 -1290 1147 -1244
<< ppolyres >>
rect -1160 -1200 -1000 1200
rect -920 -1200 -760 1200
rect -680 -1200 -520 1200
rect -440 -1200 -280 1200
rect -200 -1200 -40 1200
rect 40 -1200 200 1200
rect 280 -1200 440 1200
rect 520 -1200 680 1200
rect 760 -1200 920 1200
rect 1000 -1200 1160 1200
<< metal1 >>
rect -1158 1244 -1147 1290
rect -1013 1244 -1002 1290
rect -918 1244 -907 1290
rect -773 1244 -762 1290
rect -678 1244 -667 1290
rect -533 1244 -522 1290
rect -438 1244 -427 1290
rect -293 1244 -282 1290
rect -198 1244 -187 1290
rect -53 1244 -42 1290
rect 42 1244 53 1290
rect 187 1244 198 1290
rect 282 1244 293 1290
rect 427 1244 438 1290
rect 522 1244 533 1290
rect 667 1244 678 1290
rect 762 1244 773 1290
rect 907 1244 918 1290
rect 1002 1244 1013 1290
rect 1147 1244 1158 1290
rect -1158 -1290 -1147 -1244
rect -1013 -1290 -1002 -1244
rect -918 -1290 -907 -1244
rect -773 -1290 -762 -1244
rect -678 -1290 -667 -1244
rect -533 -1290 -522 -1244
rect -438 -1290 -427 -1244
rect -293 -1290 -282 -1244
rect -198 -1290 -187 -1244
rect -53 -1290 -42 -1244
rect 42 -1290 53 -1244
rect 187 -1290 198 -1244
rect 282 -1290 293 -1244
rect 427 -1290 438 -1244
rect 522 -1290 533 -1244
rect 667 -1290 678 -1244
rect 762 -1290 773 -1244
rect 907 -1290 918 -1244
rect 1002 -1290 1013 -1244
rect 1147 -1290 1158 -1244
<< properties >>
string FIXED_BBOX -1284 -1427 1284 1427
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 12.0 m 1 nx 10 wmin 0.80 lmin 1.00 rho 315 val 5.178k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
