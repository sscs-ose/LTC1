magic
tech gf180mcuC
magscale 1 10
timestamp 1694518401
<< nwell >>
rect 5446 15160 14427 15705
rect 5446 15038 13793 15160
rect 13845 15038 14427 15160
rect 5446 14888 14427 15038
rect 5446 14855 13586 14888
rect 13706 14855 14427 14888
rect 5446 14825 13574 14855
rect 13708 14825 14427 14855
rect 5446 14587 14427 14825
rect 5446 14585 14114 14587
rect 5446 14529 13884 14585
rect 14030 14550 14114 14585
rect 14237 14550 14427 14587
rect 5446 14514 13784 14529
rect 14030 14514 14427 14550
rect 5446 14501 13897 14514
rect 5446 14383 13369 14501
rect 13428 14500 13897 14501
rect 13460 14384 13897 14500
rect 13997 14384 14003 14514
rect 5446 14375 13411 14383
rect 13460 14382 14003 14384
rect 14073 14382 14427 14514
rect 13460 14375 14427 14382
rect 5446 12554 14427 14375
<< nsubdiff >>
rect 5488 15658 14402 15673
rect 5488 15612 5504 15658
rect 5550 15612 5598 15658
rect 5644 15612 5692 15658
rect 5738 15612 5786 15658
rect 5832 15612 5880 15658
rect 5926 15612 5974 15658
rect 6020 15612 6068 15658
rect 6114 15612 6162 15658
rect 6208 15612 6256 15658
rect 6302 15612 6350 15658
rect 6396 15612 6444 15658
rect 6490 15612 6538 15658
rect 6584 15612 6632 15658
rect 6678 15612 6726 15658
rect 6772 15612 6820 15658
rect 6866 15612 6914 15658
rect 6960 15612 7008 15658
rect 7054 15612 7102 15658
rect 7148 15612 7196 15658
rect 7242 15612 7290 15658
rect 7336 15612 7384 15658
rect 7430 15612 7478 15658
rect 7524 15612 7572 15658
rect 7618 15612 7666 15658
rect 7712 15612 7760 15658
rect 7806 15612 7854 15658
rect 7900 15612 7948 15658
rect 7994 15612 8042 15658
rect 8088 15612 8136 15658
rect 8182 15612 8230 15658
rect 8276 15612 8324 15658
rect 8370 15612 8418 15658
rect 8464 15612 8512 15658
rect 8558 15612 8606 15658
rect 8652 15612 8700 15658
rect 8746 15612 8794 15658
rect 8840 15612 8888 15658
rect 8934 15612 8982 15658
rect 9028 15612 9076 15658
rect 9122 15612 9170 15658
rect 9216 15612 9264 15658
rect 9310 15612 9358 15658
rect 9404 15612 9452 15658
rect 9498 15612 9546 15658
rect 9592 15612 9640 15658
rect 9686 15612 9734 15658
rect 9780 15612 9828 15658
rect 9874 15612 9922 15658
rect 9968 15612 10016 15658
rect 10062 15612 10110 15658
rect 10156 15612 10204 15658
rect 10250 15612 10298 15658
rect 10344 15612 10392 15658
rect 10438 15612 10486 15658
rect 10532 15612 10580 15658
rect 10626 15612 10674 15658
rect 10720 15612 10768 15658
rect 10814 15612 10862 15658
rect 10908 15612 10956 15658
rect 11002 15612 11050 15658
rect 11096 15612 11144 15658
rect 11190 15612 11238 15658
rect 11284 15612 11332 15658
rect 11378 15612 11426 15658
rect 11472 15612 11520 15658
rect 11566 15612 11614 15658
rect 11660 15612 11708 15658
rect 11754 15612 11802 15658
rect 11848 15612 11896 15658
rect 11942 15612 11990 15658
rect 12036 15612 12084 15658
rect 12130 15612 12178 15658
rect 12224 15612 12272 15658
rect 12318 15612 12366 15658
rect 12412 15612 12460 15658
rect 12506 15612 12554 15658
rect 12600 15612 12648 15658
rect 12694 15612 12742 15658
rect 12788 15612 12836 15658
rect 12882 15612 12930 15658
rect 12976 15612 13024 15658
rect 13070 15612 13118 15658
rect 13164 15612 13212 15658
rect 13258 15612 13306 15658
rect 13352 15612 13400 15658
rect 13446 15612 13494 15658
rect 13540 15612 13588 15658
rect 13634 15612 13682 15658
rect 13728 15612 13776 15658
rect 13822 15612 13870 15658
rect 13916 15612 13964 15658
rect 14010 15612 14058 15658
rect 14104 15612 14152 15658
rect 14198 15612 14246 15658
rect 14292 15612 14340 15658
rect 14386 15612 14402 15658
rect 5488 15597 14402 15612
rect 5488 15564 5564 15597
rect 5488 15518 5503 15564
rect 5549 15518 5564 15564
rect 5488 15470 5564 15518
rect 5488 15424 5503 15470
rect 5549 15424 5564 15470
rect 5488 15376 5564 15424
rect 5488 15330 5503 15376
rect 5549 15330 5564 15376
rect 5488 15282 5564 15330
rect 5488 15236 5503 15282
rect 5549 15236 5564 15282
rect 5488 15188 5564 15236
rect 5488 15142 5503 15188
rect 5549 15142 5564 15188
rect 5488 15094 5564 15142
rect 5488 15048 5503 15094
rect 5549 15048 5564 15094
rect 5488 15000 5564 15048
rect 5488 14954 5503 15000
rect 5549 14954 5564 15000
rect 5488 14906 5564 14954
rect 5488 14860 5503 14906
rect 5549 14860 5564 14906
rect 5488 14812 5564 14860
rect 5488 14766 5503 14812
rect 5549 14766 5564 14812
rect 5488 14718 5564 14766
rect 5488 14672 5503 14718
rect 5549 14672 5564 14718
rect 5488 14624 5564 14672
rect 5488 14578 5503 14624
rect 5549 14578 5564 14624
rect 5488 14530 5564 14578
rect 5488 14484 5503 14530
rect 5549 14484 5564 14530
rect 5488 14436 5564 14484
rect 5488 14390 5503 14436
rect 5549 14390 5564 14436
rect 5488 14342 5564 14390
rect 5488 14296 5503 14342
rect 5549 14296 5564 14342
rect 5488 14248 5564 14296
rect 5488 14202 5503 14248
rect 5549 14202 5564 14248
rect 5488 14154 5564 14202
rect 5488 14108 5503 14154
rect 5549 14108 5564 14154
rect 5488 14060 5564 14108
rect 5488 14014 5503 14060
rect 5549 14014 5564 14060
rect 5488 13966 5564 14014
rect 5488 13920 5503 13966
rect 5549 13920 5564 13966
rect 5488 13872 5564 13920
rect 5488 13826 5503 13872
rect 5549 13826 5564 13872
rect 5488 13778 5564 13826
rect 5488 13732 5503 13778
rect 5549 13732 5564 13778
rect 5488 13684 5564 13732
rect 5488 13638 5503 13684
rect 5549 13638 5564 13684
rect 5488 13590 5564 13638
rect 5488 13544 5503 13590
rect 5549 13544 5564 13590
rect 5488 13496 5564 13544
rect 5488 13450 5503 13496
rect 5549 13450 5564 13496
rect 5488 13402 5564 13450
rect 5488 13356 5503 13402
rect 5549 13356 5564 13402
rect 5488 13308 5564 13356
rect 5488 13262 5503 13308
rect 5549 13262 5564 13308
rect 5488 13214 5564 13262
rect 5488 13168 5503 13214
rect 5549 13168 5564 13214
rect 5488 13120 5564 13168
rect 5488 13074 5503 13120
rect 5549 13074 5564 13120
rect 5488 13026 5564 13074
rect 5488 12980 5503 13026
rect 5549 12980 5564 13026
rect 5488 12932 5564 12980
rect 5488 12886 5503 12932
rect 5549 12886 5564 12932
rect 5488 12838 5564 12886
rect 5488 12792 5503 12838
rect 5549 12792 5564 12838
rect 5488 12744 5564 12792
rect 5488 12698 5503 12744
rect 5549 12698 5564 12744
rect 5488 12665 5564 12698
rect 14326 15564 14402 15597
rect 14326 15518 14341 15564
rect 14387 15518 14402 15564
rect 14326 15470 14402 15518
rect 14326 15424 14341 15470
rect 14387 15424 14402 15470
rect 14326 15376 14402 15424
rect 14326 15330 14341 15376
rect 14387 15330 14402 15376
rect 14326 15282 14402 15330
rect 14326 15236 14341 15282
rect 14387 15236 14402 15282
rect 14326 15188 14402 15236
rect 14326 15142 14341 15188
rect 14387 15142 14402 15188
rect 14326 15094 14402 15142
rect 14326 15048 14341 15094
rect 14387 15048 14402 15094
rect 14326 15000 14402 15048
rect 14326 14954 14341 15000
rect 14387 14954 14402 15000
rect 14326 14906 14402 14954
rect 14326 14860 14341 14906
rect 14387 14860 14402 14906
rect 14326 14812 14402 14860
rect 14326 14766 14341 14812
rect 14387 14766 14402 14812
rect 14326 14718 14402 14766
rect 14326 14672 14341 14718
rect 14387 14672 14402 14718
rect 14326 14624 14402 14672
rect 14326 14578 14341 14624
rect 14387 14578 14402 14624
rect 14326 14530 14402 14578
rect 14326 14484 14341 14530
rect 14387 14484 14402 14530
rect 14326 14436 14402 14484
rect 14326 14390 14341 14436
rect 14387 14390 14402 14436
rect 14326 14342 14402 14390
rect 14326 14296 14341 14342
rect 14387 14296 14402 14342
rect 14326 14248 14402 14296
rect 14326 14202 14341 14248
rect 14387 14202 14402 14248
rect 14326 14154 14402 14202
rect 14326 14108 14341 14154
rect 14387 14108 14402 14154
rect 14326 14060 14402 14108
rect 14326 14014 14341 14060
rect 14387 14014 14402 14060
rect 14326 13966 14402 14014
rect 14326 13920 14341 13966
rect 14387 13920 14402 13966
rect 14326 13872 14402 13920
rect 14326 13826 14341 13872
rect 14387 13826 14402 13872
rect 14326 13778 14402 13826
rect 14326 13732 14341 13778
rect 14387 13732 14402 13778
rect 14326 13684 14402 13732
rect 14326 13638 14341 13684
rect 14387 13638 14402 13684
rect 14326 13590 14402 13638
rect 14326 13544 14341 13590
rect 14387 13544 14402 13590
rect 14326 13496 14402 13544
rect 14326 13450 14341 13496
rect 14387 13450 14402 13496
rect 14326 13402 14402 13450
rect 14326 13356 14341 13402
rect 14387 13356 14402 13402
rect 14326 13308 14402 13356
rect 14326 13262 14341 13308
rect 14387 13262 14402 13308
rect 14326 13214 14402 13262
rect 14326 13168 14341 13214
rect 14387 13168 14402 13214
rect 14326 13120 14402 13168
rect 14326 13074 14341 13120
rect 14387 13074 14402 13120
rect 14326 13026 14402 13074
rect 14326 12980 14341 13026
rect 14387 12980 14402 13026
rect 14326 12932 14402 12980
rect 14326 12886 14341 12932
rect 14387 12886 14402 12932
rect 14326 12838 14402 12886
rect 14326 12792 14341 12838
rect 14387 12792 14402 12838
rect 14326 12744 14402 12792
rect 14326 12698 14341 12744
rect 14387 12698 14402 12744
rect 14326 12665 14402 12698
rect 5488 12650 14402 12665
rect 5488 12604 5504 12650
rect 5550 12604 5598 12650
rect 5644 12604 5692 12650
rect 5738 12604 5786 12650
rect 5832 12604 5880 12650
rect 5926 12604 5974 12650
rect 6020 12604 6068 12650
rect 6114 12604 6162 12650
rect 6208 12604 6256 12650
rect 6302 12604 6350 12650
rect 6396 12604 6444 12650
rect 6490 12604 6538 12650
rect 6584 12604 6632 12650
rect 6678 12604 6726 12650
rect 6772 12604 6820 12650
rect 6866 12604 6914 12650
rect 6960 12604 7008 12650
rect 7054 12604 7102 12650
rect 7148 12604 7196 12650
rect 7242 12604 7290 12650
rect 7336 12604 7384 12650
rect 7430 12604 7478 12650
rect 7524 12604 7572 12650
rect 7618 12604 7666 12650
rect 7712 12604 7760 12650
rect 7806 12604 7854 12650
rect 7900 12604 7948 12650
rect 7994 12604 8042 12650
rect 8088 12604 8136 12650
rect 8182 12604 8230 12650
rect 8276 12604 8324 12650
rect 8370 12604 8418 12650
rect 8464 12604 8512 12650
rect 8558 12604 8606 12650
rect 8652 12604 8700 12650
rect 8746 12604 8794 12650
rect 8840 12604 8888 12650
rect 8934 12604 8982 12650
rect 9028 12604 9076 12650
rect 9122 12604 9170 12650
rect 9216 12604 9264 12650
rect 9310 12604 9358 12650
rect 9404 12604 9452 12650
rect 9498 12604 9546 12650
rect 9592 12604 9640 12650
rect 9686 12604 9734 12650
rect 9780 12604 9828 12650
rect 9874 12604 9922 12650
rect 9968 12604 10016 12650
rect 10062 12604 10110 12650
rect 10156 12604 10204 12650
rect 10250 12604 10298 12650
rect 10344 12604 10392 12650
rect 10438 12604 10486 12650
rect 10532 12604 10580 12650
rect 10626 12604 10674 12650
rect 10720 12604 10768 12650
rect 10814 12604 10862 12650
rect 10908 12604 10956 12650
rect 11002 12604 11050 12650
rect 11096 12604 11144 12650
rect 11190 12604 11238 12650
rect 11284 12604 11332 12650
rect 11378 12604 11426 12650
rect 11472 12604 11520 12650
rect 11566 12604 11614 12650
rect 11660 12604 11708 12650
rect 11754 12604 11802 12650
rect 11848 12604 11896 12650
rect 11942 12604 11990 12650
rect 12036 12604 12084 12650
rect 12130 12604 12178 12650
rect 12224 12604 12272 12650
rect 12318 12604 12366 12650
rect 12412 12604 12460 12650
rect 12506 12604 12554 12650
rect 12600 12604 12648 12650
rect 12694 12604 12742 12650
rect 12788 12604 12836 12650
rect 12882 12604 12930 12650
rect 12976 12604 13024 12650
rect 13070 12604 13118 12650
rect 13164 12604 13212 12650
rect 13258 12604 13306 12650
rect 13352 12604 13400 12650
rect 13446 12604 13494 12650
rect 13540 12604 13588 12650
rect 13634 12604 13682 12650
rect 13728 12604 13776 12650
rect 13822 12604 13870 12650
rect 13916 12604 13964 12650
rect 14010 12604 14058 12650
rect 14104 12604 14152 12650
rect 14198 12604 14246 12650
rect 14292 12604 14340 12650
rect 14386 12604 14402 12650
rect 5488 12589 14402 12604
<< nsubdiffcont >>
rect 5504 15612 5550 15658
rect 5598 15612 5644 15658
rect 5692 15612 5738 15658
rect 5786 15612 5832 15658
rect 5880 15612 5926 15658
rect 5974 15612 6020 15658
rect 6068 15612 6114 15658
rect 6162 15612 6208 15658
rect 6256 15612 6302 15658
rect 6350 15612 6396 15658
rect 6444 15612 6490 15658
rect 6538 15612 6584 15658
rect 6632 15612 6678 15658
rect 6726 15612 6772 15658
rect 6820 15612 6866 15658
rect 6914 15612 6960 15658
rect 7008 15612 7054 15658
rect 7102 15612 7148 15658
rect 7196 15612 7242 15658
rect 7290 15612 7336 15658
rect 7384 15612 7430 15658
rect 7478 15612 7524 15658
rect 7572 15612 7618 15658
rect 7666 15612 7712 15658
rect 7760 15612 7806 15658
rect 7854 15612 7900 15658
rect 7948 15612 7994 15658
rect 8042 15612 8088 15658
rect 8136 15612 8182 15658
rect 8230 15612 8276 15658
rect 8324 15612 8370 15658
rect 8418 15612 8464 15658
rect 8512 15612 8558 15658
rect 8606 15612 8652 15658
rect 8700 15612 8746 15658
rect 8794 15612 8840 15658
rect 8888 15612 8934 15658
rect 8982 15612 9028 15658
rect 9076 15612 9122 15658
rect 9170 15612 9216 15658
rect 9264 15612 9310 15658
rect 9358 15612 9404 15658
rect 9452 15612 9498 15658
rect 9546 15612 9592 15658
rect 9640 15612 9686 15658
rect 9734 15612 9780 15658
rect 9828 15612 9874 15658
rect 9922 15612 9968 15658
rect 10016 15612 10062 15658
rect 10110 15612 10156 15658
rect 10204 15612 10250 15658
rect 10298 15612 10344 15658
rect 10392 15612 10438 15658
rect 10486 15612 10532 15658
rect 10580 15612 10626 15658
rect 10674 15612 10720 15658
rect 10768 15612 10814 15658
rect 10862 15612 10908 15658
rect 10956 15612 11002 15658
rect 11050 15612 11096 15658
rect 11144 15612 11190 15658
rect 11238 15612 11284 15658
rect 11332 15612 11378 15658
rect 11426 15612 11472 15658
rect 11520 15612 11566 15658
rect 11614 15612 11660 15658
rect 11708 15612 11754 15658
rect 11802 15612 11848 15658
rect 11896 15612 11942 15658
rect 11990 15612 12036 15658
rect 12084 15612 12130 15658
rect 12178 15612 12224 15658
rect 12272 15612 12318 15658
rect 12366 15612 12412 15658
rect 12460 15612 12506 15658
rect 12554 15612 12600 15658
rect 12648 15612 12694 15658
rect 12742 15612 12788 15658
rect 12836 15612 12882 15658
rect 12930 15612 12976 15658
rect 13024 15612 13070 15658
rect 13118 15612 13164 15658
rect 13212 15612 13258 15658
rect 13306 15612 13352 15658
rect 13400 15612 13446 15658
rect 13494 15612 13540 15658
rect 13588 15612 13634 15658
rect 13682 15612 13728 15658
rect 13776 15612 13822 15658
rect 13870 15612 13916 15658
rect 13964 15612 14010 15658
rect 14058 15612 14104 15658
rect 14152 15612 14198 15658
rect 14246 15612 14292 15658
rect 14340 15612 14386 15658
rect 5503 15518 5549 15564
rect 5503 15424 5549 15470
rect 5503 15330 5549 15376
rect 5503 15236 5549 15282
rect 5503 15142 5549 15188
rect 5503 15048 5549 15094
rect 5503 14954 5549 15000
rect 5503 14860 5549 14906
rect 5503 14766 5549 14812
rect 5503 14672 5549 14718
rect 5503 14578 5549 14624
rect 5503 14484 5549 14530
rect 5503 14390 5549 14436
rect 5503 14296 5549 14342
rect 5503 14202 5549 14248
rect 5503 14108 5549 14154
rect 5503 14014 5549 14060
rect 5503 13920 5549 13966
rect 5503 13826 5549 13872
rect 5503 13732 5549 13778
rect 5503 13638 5549 13684
rect 5503 13544 5549 13590
rect 5503 13450 5549 13496
rect 5503 13356 5549 13402
rect 5503 13262 5549 13308
rect 5503 13168 5549 13214
rect 5503 13074 5549 13120
rect 5503 12980 5549 13026
rect 5503 12886 5549 12932
rect 5503 12792 5549 12838
rect 5503 12698 5549 12744
rect 14341 15518 14387 15564
rect 14341 15424 14387 15470
rect 14341 15330 14387 15376
rect 14341 15236 14387 15282
rect 14341 15142 14387 15188
rect 14341 15048 14387 15094
rect 14341 14954 14387 15000
rect 14341 14860 14387 14906
rect 14341 14766 14387 14812
rect 14341 14672 14387 14718
rect 14341 14578 14387 14624
rect 14341 14484 14387 14530
rect 14341 14390 14387 14436
rect 14341 14296 14387 14342
rect 14341 14202 14387 14248
rect 14341 14108 14387 14154
rect 14341 14014 14387 14060
rect 14341 13920 14387 13966
rect 14341 13826 14387 13872
rect 14341 13732 14387 13778
rect 14341 13638 14387 13684
rect 14341 13544 14387 13590
rect 14341 13450 14387 13496
rect 14341 13356 14387 13402
rect 14341 13262 14387 13308
rect 14341 13168 14387 13214
rect 14341 13074 14387 13120
rect 14341 12980 14387 13026
rect 14341 12886 14387 12932
rect 14341 12792 14387 12838
rect 14341 12698 14387 12744
rect 5504 12604 5550 12650
rect 5598 12604 5644 12650
rect 5692 12604 5738 12650
rect 5786 12604 5832 12650
rect 5880 12604 5926 12650
rect 5974 12604 6020 12650
rect 6068 12604 6114 12650
rect 6162 12604 6208 12650
rect 6256 12604 6302 12650
rect 6350 12604 6396 12650
rect 6444 12604 6490 12650
rect 6538 12604 6584 12650
rect 6632 12604 6678 12650
rect 6726 12604 6772 12650
rect 6820 12604 6866 12650
rect 6914 12604 6960 12650
rect 7008 12604 7054 12650
rect 7102 12604 7148 12650
rect 7196 12604 7242 12650
rect 7290 12604 7336 12650
rect 7384 12604 7430 12650
rect 7478 12604 7524 12650
rect 7572 12604 7618 12650
rect 7666 12604 7712 12650
rect 7760 12604 7806 12650
rect 7854 12604 7900 12650
rect 7948 12604 7994 12650
rect 8042 12604 8088 12650
rect 8136 12604 8182 12650
rect 8230 12604 8276 12650
rect 8324 12604 8370 12650
rect 8418 12604 8464 12650
rect 8512 12604 8558 12650
rect 8606 12604 8652 12650
rect 8700 12604 8746 12650
rect 8794 12604 8840 12650
rect 8888 12604 8934 12650
rect 8982 12604 9028 12650
rect 9076 12604 9122 12650
rect 9170 12604 9216 12650
rect 9264 12604 9310 12650
rect 9358 12604 9404 12650
rect 9452 12604 9498 12650
rect 9546 12604 9592 12650
rect 9640 12604 9686 12650
rect 9734 12604 9780 12650
rect 9828 12604 9874 12650
rect 9922 12604 9968 12650
rect 10016 12604 10062 12650
rect 10110 12604 10156 12650
rect 10204 12604 10250 12650
rect 10298 12604 10344 12650
rect 10392 12604 10438 12650
rect 10486 12604 10532 12650
rect 10580 12604 10626 12650
rect 10674 12604 10720 12650
rect 10768 12604 10814 12650
rect 10862 12604 10908 12650
rect 10956 12604 11002 12650
rect 11050 12604 11096 12650
rect 11144 12604 11190 12650
rect 11238 12604 11284 12650
rect 11332 12604 11378 12650
rect 11426 12604 11472 12650
rect 11520 12604 11566 12650
rect 11614 12604 11660 12650
rect 11708 12604 11754 12650
rect 11802 12604 11848 12650
rect 11896 12604 11942 12650
rect 11990 12604 12036 12650
rect 12084 12604 12130 12650
rect 12178 12604 12224 12650
rect 12272 12604 12318 12650
rect 12366 12604 12412 12650
rect 12460 12604 12506 12650
rect 12554 12604 12600 12650
rect 12648 12604 12694 12650
rect 12742 12604 12788 12650
rect 12836 12604 12882 12650
rect 12930 12604 12976 12650
rect 13024 12604 13070 12650
rect 13118 12604 13164 12650
rect 13212 12604 13258 12650
rect 13306 12604 13352 12650
rect 13400 12604 13446 12650
rect 13494 12604 13540 12650
rect 13588 12604 13634 12650
rect 13682 12604 13728 12650
rect 13776 12604 13822 12650
rect 13870 12604 13916 12650
rect 13964 12604 14010 12650
rect 14058 12604 14104 12650
rect 14152 12604 14198 12650
rect 14246 12604 14292 12650
rect 14340 12604 14386 12650
<< metal1 >>
rect 5477 15658 14413 15684
rect 5477 15612 5504 15658
rect 5550 15612 5598 15658
rect 5644 15612 5692 15658
rect 5738 15612 5786 15658
rect 5832 15612 5880 15658
rect 5926 15612 5974 15658
rect 6020 15612 6068 15658
rect 6114 15612 6162 15658
rect 6208 15612 6256 15658
rect 6302 15612 6350 15658
rect 6396 15612 6444 15658
rect 6490 15612 6538 15658
rect 6584 15612 6632 15658
rect 6678 15612 6726 15658
rect 6772 15612 6820 15658
rect 6866 15612 6914 15658
rect 6960 15612 7008 15658
rect 7054 15612 7102 15658
rect 7148 15612 7196 15658
rect 7242 15612 7290 15658
rect 7336 15612 7384 15658
rect 7430 15612 7478 15658
rect 7524 15612 7572 15658
rect 7618 15612 7666 15658
rect 7712 15612 7760 15658
rect 7806 15612 7854 15658
rect 7900 15612 7948 15658
rect 7994 15612 8042 15658
rect 8088 15612 8136 15658
rect 8182 15612 8230 15658
rect 8276 15612 8324 15658
rect 8370 15612 8418 15658
rect 8464 15612 8512 15658
rect 8558 15612 8606 15658
rect 8652 15612 8700 15658
rect 8746 15612 8794 15658
rect 8840 15612 8888 15658
rect 8934 15612 8982 15658
rect 9028 15612 9076 15658
rect 9122 15612 9170 15658
rect 9216 15612 9264 15658
rect 9310 15612 9358 15658
rect 9404 15612 9452 15658
rect 9498 15612 9546 15658
rect 9592 15612 9640 15658
rect 9686 15612 9734 15658
rect 9780 15612 9828 15658
rect 9874 15612 9922 15658
rect 9968 15612 10016 15658
rect 10062 15612 10110 15658
rect 10156 15612 10204 15658
rect 10250 15612 10298 15658
rect 10344 15612 10392 15658
rect 10438 15612 10486 15658
rect 10532 15612 10580 15658
rect 10626 15612 10674 15658
rect 10720 15612 10768 15658
rect 10814 15612 10862 15658
rect 10908 15612 10956 15658
rect 11002 15612 11050 15658
rect 11096 15612 11144 15658
rect 11190 15612 11238 15658
rect 11284 15612 11332 15658
rect 11378 15612 11426 15658
rect 11472 15612 11520 15658
rect 11566 15612 11614 15658
rect 11660 15612 11708 15658
rect 11754 15612 11802 15658
rect 11848 15612 11896 15658
rect 11942 15612 11990 15658
rect 12036 15612 12084 15658
rect 12130 15612 12178 15658
rect 12224 15612 12272 15658
rect 12318 15612 12366 15658
rect 12412 15612 12460 15658
rect 12506 15612 12554 15658
rect 12600 15612 12648 15658
rect 12694 15612 12742 15658
rect 12788 15612 12836 15658
rect 12882 15612 12930 15658
rect 12976 15612 13024 15658
rect 13070 15612 13118 15658
rect 13164 15612 13212 15658
rect 13258 15612 13306 15658
rect 13352 15612 13400 15658
rect 13446 15612 13494 15658
rect 13540 15612 13588 15658
rect 13634 15612 13682 15658
rect 13728 15612 13776 15658
rect 13822 15612 13870 15658
rect 13916 15612 13964 15658
rect 14010 15612 14058 15658
rect 14104 15612 14152 15658
rect 14198 15612 14246 15658
rect 14292 15612 14340 15658
rect 14386 15612 14413 15658
rect 5477 15586 14413 15612
rect 5477 15564 5575 15586
rect 5477 15518 5503 15564
rect 5549 15518 5575 15564
rect 5477 15470 5575 15518
rect 5477 15424 5503 15470
rect 5549 15424 5575 15470
rect 5477 15376 5575 15424
rect 5477 15330 5503 15376
rect 5549 15330 5575 15376
rect 5477 15282 5575 15330
rect 5477 15236 5503 15282
rect 5549 15236 5575 15282
rect 5477 15188 5575 15236
rect 5477 15142 5503 15188
rect 5549 15142 5575 15188
rect 5477 15094 5575 15142
rect 5477 15048 5503 15094
rect 5549 15048 5575 15094
rect 5477 15000 5575 15048
rect 5477 14954 5503 15000
rect 5549 14954 5575 15000
rect 5477 14906 5575 14954
rect 5477 14860 5503 14906
rect 5549 14860 5575 14906
rect 5477 14812 5575 14860
rect 5477 14766 5503 14812
rect 5549 14766 5575 14812
rect 5477 14718 5575 14766
rect 5477 14672 5503 14718
rect 5549 14672 5575 14718
rect 5667 14920 5755 14932
rect 5667 14856 5679 14920
rect 5743 14856 5755 14920
rect 5904 14919 5983 15586
rect 6149 15237 6160 15283
rect 6218 14976 6318 15386
rect 6374 15237 6385 15283
rect 6535 15141 6635 15416
rect 9419 15380 10475 15480
rect 6789 15237 6800 15283
rect 6851 15221 7294 15309
rect 7438 15301 7657 15313
rect 7438 15283 7451 15301
rect 7334 15237 7345 15283
rect 7429 15237 7451 15283
rect 7515 15237 7581 15301
rect 7645 15283 7657 15301
rect 7645 15237 7665 15283
rect 7749 15237 7760 15283
rect 7438 15225 7657 15237
rect 7831 15219 8223 15307
rect 8397 15301 8616 15313
rect 8397 15283 8409 15301
rect 8294 15237 8305 15283
rect 8389 15237 8409 15283
rect 8473 15237 8539 15301
rect 8603 15283 8616 15301
rect 8603 15237 8625 15283
rect 8709 15237 8720 15283
rect 8397 15225 8616 15237
rect 8760 15221 9203 15309
rect 9254 15237 9265 15283
rect 9349 15237 9360 15283
rect 9419 15241 9519 15380
rect 9574 15237 9585 15283
rect 9669 15237 9680 15283
rect 9749 15222 10147 15310
rect 10214 15237 10225 15283
rect 10309 15237 10320 15283
rect 10375 15241 10475 15380
rect 10534 15237 10545 15283
rect 10629 15237 10640 15283
rect 10691 15221 11134 15309
rect 11278 15301 11497 15313
rect 11278 15283 11291 15301
rect 11174 15237 11185 15283
rect 11269 15237 11291 15283
rect 11355 15237 11421 15301
rect 11485 15283 11497 15301
rect 11485 15237 11505 15283
rect 11589 15237 11600 15283
rect 11278 15225 11497 15237
rect 11671 15219 12063 15307
rect 12237 15301 12456 15313
rect 12237 15283 12249 15301
rect 12134 15237 12145 15283
rect 12229 15237 12249 15283
rect 12313 15237 12379 15301
rect 12443 15283 12456 15301
rect 12443 15237 12465 15283
rect 12549 15237 12560 15283
rect 12237 15225 12456 15237
rect 12600 15221 13043 15309
rect 13414 15304 13504 15453
rect 13094 15237 13105 15283
rect 13189 15237 13200 15283
rect 13264 15214 13676 15304
rect 13734 15237 13745 15283
rect 13916 15259 14001 15586
rect 14315 15564 14413 15586
rect 14315 15518 14341 15564
rect 14387 15518 14413 15564
rect 14315 15470 14413 15518
rect 14315 15424 14341 15470
rect 14387 15424 14413 15470
rect 14315 15376 14413 15424
rect 14315 15330 14341 15376
rect 14387 15330 14413 15376
rect 14315 15282 14413 15330
rect 6535 15041 6950 15141
rect 6158 14964 6377 14976
rect 6158 14951 6171 14964
rect 6149 14905 6171 14951
rect 6158 14900 6171 14905
rect 6235 14900 6301 14964
rect 6365 14951 6377 14964
rect 6475 14962 6694 14974
rect 6475 14951 6488 14962
rect 6365 14905 6385 14951
rect 6469 14905 6488 14951
rect 6365 14900 6377 14905
rect 6158 14888 6377 14900
rect 6475 14898 6488 14905
rect 6552 14898 6618 14962
rect 6682 14951 6694 14962
rect 6682 14905 6705 14951
rect 6850 14917 6950 15041
rect 7109 14905 7120 14951
rect 6682 14898 6694 14905
rect 6475 14886 6694 14898
rect 5667 14813 5755 14856
rect 7177 14824 7277 14949
rect 7334 14905 7345 14951
rect 7429 14905 7440 14951
rect 7486 14886 7929 14974
rect 8125 14886 8568 14974
rect 9037 14965 9256 14977
rect 9037 14951 9049 14965
rect 8614 14905 8625 14951
rect 8709 14905 8720 14951
rect 8777 14824 8877 14949
rect 8934 14905 8945 14951
rect 9029 14905 9049 14951
rect 9037 14901 9049 14905
rect 9113 14901 9179 14965
rect 9243 14951 9256 14965
rect 9360 14962 9579 14974
rect 9360 14951 9372 14962
rect 9243 14905 9265 14951
rect 9349 14905 9372 14951
rect 9243 14901 9256 14905
rect 9037 14889 9256 14901
rect 9360 14898 9372 14905
rect 9436 14898 9502 14962
rect 9566 14951 9579 14962
rect 9677 14964 9896 14976
rect 9677 14951 9689 14964
rect 9566 14905 9585 14951
rect 9669 14905 9689 14951
rect 9566 14898 9579 14905
rect 9360 14886 9579 14898
rect 9677 14900 9689 14905
rect 9753 14900 9819 14964
rect 9883 14951 9896 14964
rect 9998 14964 10217 14976
rect 9998 14951 10011 14964
rect 9883 14905 9905 14951
rect 9989 14905 10011 14951
rect 9883 14900 9896 14905
rect 9677 14888 9896 14900
rect 9998 14900 10011 14905
rect 10075 14900 10141 14964
rect 10205 14951 10217 14964
rect 10315 14962 10534 14974
rect 10315 14951 10328 14962
rect 10205 14905 10225 14951
rect 10309 14905 10328 14951
rect 10205 14900 10217 14905
rect 9998 14888 10217 14900
rect 10315 14898 10328 14905
rect 10392 14898 10458 14962
rect 10522 14951 10534 14962
rect 10638 14965 10857 14977
rect 10638 14951 10651 14965
rect 10522 14905 10545 14951
rect 10629 14905 10651 14951
rect 10522 14898 10534 14905
rect 10315 14886 10534 14898
rect 10638 14901 10651 14905
rect 10715 14901 10781 14965
rect 10845 14951 10857 14965
rect 10845 14905 10865 14951
rect 10949 14905 10960 14951
rect 10845 14901 10857 14905
rect 10638 14889 10857 14901
rect 5667 14790 6638 14813
rect 5667 14726 5679 14790
rect 5743 14726 6638 14790
rect 5667 14713 6638 14726
rect 7177 14724 7600 14824
rect 5477 14631 5575 14672
rect 5477 14624 5970 14631
rect 5477 14578 5503 14624
rect 5549 14583 5970 14624
rect 6171 14615 6306 14650
rect 5549 14578 5575 14583
rect 5477 14530 5575 14578
rect 6171 14562 6313 14615
rect 6374 14585 6385 14631
rect 6469 14585 6480 14631
rect 6538 14593 6638 14713
rect 6694 14585 6705 14631
rect 6789 14585 6800 14631
rect 6847 14566 7290 14654
rect 7334 14585 7345 14631
rect 7429 14585 7440 14631
rect 7500 14591 7600 14724
rect 8454 14724 8877 14824
rect 11017 14824 11117 14949
rect 11174 14905 11185 14951
rect 11269 14905 11280 14951
rect 11326 14886 11769 14974
rect 11965 14886 12408 14974
rect 12877 14965 13096 14977
rect 13576 14976 13676 15214
rect 14315 15236 14341 15282
rect 14387 15236 14413 15282
rect 14315 15188 14413 15236
rect 14315 15142 14341 15188
rect 14387 15142 14413 15188
rect 14315 15094 14413 15142
rect 14315 15048 14341 15094
rect 14387 15048 14413 15094
rect 14315 15000 14413 15048
rect 12877 14951 12889 14965
rect 12454 14905 12465 14951
rect 12549 14905 12560 14951
rect 12617 14824 12717 14949
rect 12774 14905 12785 14951
rect 12869 14905 12889 14951
rect 12877 14901 12889 14905
rect 12953 14901 13019 14965
rect 13083 14951 13096 14965
rect 13200 14962 13419 14974
rect 13200 14951 13212 14962
rect 13083 14905 13105 14951
rect 13189 14905 13212 14951
rect 13083 14901 13096 14905
rect 12877 14889 13096 14901
rect 13200 14898 13212 14905
rect 13276 14898 13342 14962
rect 13406 14951 13419 14962
rect 13517 14964 13736 14976
rect 13517 14951 13529 14964
rect 13406 14905 13425 14951
rect 13509 14905 13529 14951
rect 13406 14898 13419 14905
rect 13200 14886 13419 14898
rect 13517 14900 13529 14905
rect 13593 14900 13659 14964
rect 13723 14951 13736 14964
rect 14315 14954 14341 15000
rect 14387 14954 14413 15000
rect 14315 14953 14413 14954
rect 13723 14905 13745 14951
rect 13917 14906 14413 14953
rect 13723 14900 13736 14905
rect 13917 14903 14341 14906
rect 13517 14888 13736 14900
rect 7654 14585 7665 14631
rect 7749 14585 7760 14631
rect 7800 14578 8240 14666
rect 8294 14585 8305 14631
rect 8389 14585 8400 14631
rect 8454 14591 8554 14724
rect 9416 14713 10478 14813
rect 11017 14724 11440 14824
rect 8614 14585 8625 14631
rect 8709 14585 8720 14631
rect 8764 14566 9207 14654
rect 9254 14585 9265 14631
rect 9349 14585 9360 14631
rect 9416 14593 9516 14713
rect 9574 14585 9585 14631
rect 9669 14585 9680 14631
rect 9748 14562 10146 14650
rect 10214 14585 10225 14631
rect 10309 14585 10320 14631
rect 10378 14593 10478 14713
rect 10534 14585 10545 14631
rect 10629 14585 10640 14631
rect 10687 14566 11130 14654
rect 11174 14585 11185 14631
rect 11269 14585 11280 14631
rect 11340 14591 11440 14724
rect 12294 14724 12717 14824
rect 14315 14860 14341 14903
rect 14387 14860 14413 14906
rect 13256 14794 14227 14813
rect 13256 14730 14146 14794
rect 14210 14730 14227 14794
rect 11494 14585 11505 14631
rect 11589 14585 11600 14631
rect 11643 14576 12083 14664
rect 12134 14585 12145 14631
rect 12229 14585 12240 14631
rect 12294 14591 12394 14724
rect 13256 14713 14227 14730
rect 12454 14585 12465 14631
rect 12549 14585 12560 14631
rect 12604 14566 13047 14654
rect 13094 14585 13105 14631
rect 13189 14585 13200 14631
rect 13256 14593 13356 14713
rect 14127 14664 14227 14713
rect 13414 14585 13425 14631
rect 5477 14484 5503 14530
rect 5549 14484 5575 14530
rect 6213 14497 6313 14562
rect 5477 14436 5575 14484
rect 5477 14390 5503 14436
rect 5549 14390 5575 14436
rect 5477 14342 5575 14390
rect 5477 14296 5503 14342
rect 5549 14296 5575 14342
rect 5477 14248 5575 14296
rect 5477 14202 5503 14248
rect 5549 14202 5575 14248
rect 5477 14154 5575 14202
rect 5477 14108 5503 14154
rect 5549 14108 5575 14154
rect 5477 14060 5575 14108
rect 5477 14014 5503 14060
rect 5549 14014 5575 14060
rect 5477 13966 5575 14014
rect 5477 13920 5503 13966
rect 5549 13920 5575 13966
rect 5477 13872 5575 13920
rect 5477 13826 5503 13872
rect 5549 13826 5575 13872
rect 5477 13778 5575 13826
rect 5477 13732 5503 13778
rect 5549 13732 5575 13778
rect 5667 14397 6313 14497
rect 13574 14495 13674 14617
rect 5667 13847 5767 14397
rect 6213 14321 6313 14397
rect 7496 14395 8558 14495
rect 6155 14309 6374 14321
rect 6155 14299 6168 14309
rect 5900 14152 5983 14290
rect 6149 14253 6168 14299
rect 6155 14245 6168 14253
rect 6232 14245 6298 14309
rect 6362 14299 6374 14309
rect 6477 14308 6696 14320
rect 6477 14299 6490 14308
rect 6362 14253 6385 14299
rect 6469 14253 6490 14299
rect 6362 14245 6374 14253
rect 6155 14233 6374 14245
rect 6477 14244 6490 14253
rect 6554 14244 6620 14308
rect 6684 14299 6696 14308
rect 7119 14304 7338 14316
rect 7119 14299 7132 14304
rect 6684 14253 6705 14299
rect 6789 14253 6800 14299
rect 6684 14244 6696 14253
rect 6477 14232 6696 14244
rect 5869 14140 6088 14152
rect 6831 14150 6931 14290
rect 7014 14253 7025 14299
rect 7109 14253 7132 14299
rect 7119 14240 7132 14253
rect 7196 14240 7262 14304
rect 7326 14299 7338 14304
rect 7326 14253 7345 14299
rect 7429 14253 7440 14299
rect 7496 14258 7596 14395
rect 7759 14312 7978 14324
rect 7759 14299 7772 14312
rect 7654 14253 7665 14299
rect 7749 14253 7772 14299
rect 7326 14240 7338 14253
rect 7119 14228 7338 14240
rect 7759 14248 7772 14253
rect 7836 14248 7902 14312
rect 7966 14299 7978 14312
rect 8076 14312 8295 14324
rect 8076 14299 8088 14312
rect 7966 14253 7985 14299
rect 8069 14253 8088 14299
rect 7966 14248 7978 14253
rect 7759 14236 7978 14248
rect 8076 14248 8088 14253
rect 8152 14248 8218 14312
rect 8282 14299 8295 14312
rect 8282 14253 8305 14299
rect 8389 14253 8400 14299
rect 8458 14258 8558 14395
rect 11336 14395 12398 14495
rect 13574 14475 13890 14495
rect 13574 14411 13683 14475
rect 13747 14411 13813 14475
rect 13877 14411 13890 14475
rect 13574 14395 13890 14411
rect 8716 14304 8935 14316
rect 8716 14299 8728 14304
rect 8614 14253 8625 14299
rect 8709 14253 8728 14299
rect 8282 14248 8295 14253
rect 8076 14236 8295 14248
rect 8716 14240 8728 14253
rect 8792 14240 8858 14304
rect 8922 14299 8935 14304
rect 9358 14308 9577 14320
rect 9358 14299 9370 14308
rect 8922 14253 8945 14299
rect 9029 14253 9040 14299
rect 8922 14240 8935 14253
rect 8716 14228 8935 14240
rect 5869 14076 5881 14140
rect 5945 14076 6011 14140
rect 6075 14076 6088 14140
rect 5869 14064 6088 14076
rect 5900 13949 5983 14064
rect 6216 14050 6931 14150
rect 7502 14052 8552 14151
rect 6149 13933 6160 13979
rect 6216 13967 6316 14050
rect 7502 14041 7601 14052
rect 6475 13989 6694 14001
rect 7118 13991 7337 14003
rect 6475 13979 6488 13989
rect 6216 13939 6317 13967
rect 6217 13847 6317 13939
rect 6374 13933 6385 13979
rect 6469 13933 6488 13979
rect 6475 13925 6488 13933
rect 6552 13925 6618 13989
rect 6682 13979 6694 13989
rect 6796 13979 7015 13990
rect 7118 13979 7131 13991
rect 6682 13933 6705 13979
rect 6789 13978 7025 13979
rect 6789 13933 6809 13978
rect 6682 13925 6694 13933
rect 6475 13913 6694 13925
rect 6796 13914 6809 13933
rect 6873 13914 6939 13978
rect 7003 13933 7025 13978
rect 7109 13933 7131 13979
rect 7003 13914 7015 13933
rect 7118 13927 7131 13933
rect 7195 13927 7261 13991
rect 7325 13979 7337 13991
rect 7325 13933 7345 13979
rect 7429 13933 7440 13979
rect 7501 13944 7601 14041
rect 8453 14041 8552 14052
rect 9123 14150 9223 14290
rect 9254 14253 9265 14299
rect 9349 14253 9370 14299
rect 9358 14244 9370 14253
rect 9434 14244 9500 14308
rect 9564 14299 9577 14308
rect 9680 14309 9899 14321
rect 9680 14299 9692 14309
rect 9564 14253 9585 14299
rect 9669 14253 9692 14299
rect 9564 14244 9577 14253
rect 9358 14232 9577 14244
rect 9680 14245 9692 14253
rect 9756 14245 9822 14309
rect 9886 14299 9899 14309
rect 9995 14309 10214 14321
rect 9995 14299 10008 14309
rect 9886 14253 9905 14299
rect 9989 14253 10008 14299
rect 9886 14245 9899 14253
rect 9680 14233 9899 14245
rect 9995 14245 10008 14253
rect 10072 14245 10138 14309
rect 10202 14299 10214 14309
rect 10317 14308 10536 14320
rect 10317 14299 10330 14308
rect 10202 14253 10225 14299
rect 10309 14253 10330 14299
rect 10202 14245 10214 14253
rect 9995 14233 10214 14245
rect 10317 14244 10330 14253
rect 10394 14244 10460 14308
rect 10524 14299 10536 14308
rect 10959 14304 11178 14316
rect 10959 14299 10972 14304
rect 10524 14253 10545 14299
rect 10629 14253 10640 14299
rect 10524 14244 10536 14253
rect 10317 14232 10536 14244
rect 10671 14150 10771 14290
rect 10854 14253 10865 14299
rect 10949 14253 10972 14299
rect 10959 14240 10972 14253
rect 11036 14240 11102 14304
rect 11166 14299 11178 14304
rect 11166 14253 11185 14299
rect 11269 14253 11280 14299
rect 11336 14258 11436 14395
rect 11599 14312 11818 14324
rect 11599 14299 11612 14312
rect 11494 14253 11505 14299
rect 11589 14253 11612 14299
rect 11166 14240 11178 14253
rect 10959 14228 11178 14240
rect 11599 14248 11612 14253
rect 11676 14248 11742 14312
rect 11806 14299 11818 14312
rect 11916 14312 12135 14324
rect 11916 14299 11928 14312
rect 11806 14253 11825 14299
rect 11909 14253 11928 14299
rect 11806 14248 11818 14253
rect 11599 14236 11818 14248
rect 11916 14248 11928 14253
rect 11992 14248 12058 14312
rect 12122 14299 12135 14312
rect 12122 14253 12145 14299
rect 12229 14253 12240 14299
rect 12298 14258 12398 14395
rect 12556 14304 12775 14316
rect 12556 14299 12568 14304
rect 12454 14253 12465 14299
rect 12549 14253 12568 14299
rect 12122 14248 12135 14253
rect 11916 14236 12135 14248
rect 12556 14240 12568 14253
rect 12632 14240 12698 14304
rect 12762 14299 12775 14304
rect 13198 14308 13417 14320
rect 13198 14299 13210 14308
rect 12762 14253 12785 14299
rect 12869 14253 12880 14299
rect 12762 14240 12775 14253
rect 12556 14228 12775 14240
rect 9123 14050 9838 14150
rect 7758 13987 7977 13999
rect 7758 13979 7771 13987
rect 7654 13933 7665 13979
rect 7749 13933 7771 13979
rect 7325 13927 7337 13933
rect 7118 13915 7337 13927
rect 7758 13923 7771 13933
rect 7835 13923 7901 13987
rect 7965 13979 7977 13987
rect 8077 13987 8296 13999
rect 8077 13979 8089 13987
rect 7965 13933 7985 13979
rect 8069 13933 8089 13979
rect 7965 13923 7977 13933
rect 6796 13902 7015 13914
rect 7758 13911 7977 13923
rect 8077 13923 8089 13933
rect 8153 13923 8219 13987
rect 8283 13979 8296 13987
rect 8283 13933 8305 13979
rect 8389 13933 8400 13979
rect 8453 13944 8553 14041
rect 8717 13991 8936 14003
rect 8717 13979 8729 13991
rect 8614 13933 8625 13979
rect 8709 13933 8729 13979
rect 8283 13923 8296 13933
rect 8077 13911 8296 13923
rect 8717 13927 8729 13933
rect 8793 13927 8859 13991
rect 8923 13979 8936 13991
rect 9039 13979 9258 13990
rect 9360 13989 9579 14001
rect 9360 13979 9372 13989
rect 8923 13933 8945 13979
rect 9029 13978 9265 13979
rect 9029 13933 9051 13978
rect 8923 13927 8936 13933
rect 8717 13915 8936 13927
rect 9039 13914 9051 13933
rect 9115 13914 9181 13978
rect 9245 13933 9265 13978
rect 9349 13933 9372 13979
rect 9245 13914 9258 13933
rect 9039 13902 9258 13914
rect 9360 13925 9372 13933
rect 9436 13925 9502 13989
rect 9566 13979 9579 13989
rect 9566 13933 9585 13979
rect 9669 13933 9680 13979
rect 9738 13939 9838 14050
rect 10056 14050 10771 14150
rect 11342 14052 12392 14151
rect 10056 13939 10156 14050
rect 11342 14041 11441 14052
rect 10315 13989 10534 14001
rect 10958 13991 11177 14003
rect 10315 13979 10328 13989
rect 10214 13933 10225 13979
rect 10309 13933 10328 13979
rect 9566 13925 9579 13933
rect 9360 13913 9579 13925
rect 10315 13925 10328 13933
rect 10392 13925 10458 13989
rect 10522 13979 10534 13989
rect 10636 13979 10855 13990
rect 10958 13979 10971 13991
rect 10522 13933 10545 13979
rect 10629 13978 10865 13979
rect 10629 13933 10649 13978
rect 10522 13925 10534 13933
rect 10315 13913 10534 13925
rect 10636 13914 10649 13933
rect 10713 13914 10779 13978
rect 10843 13933 10865 13978
rect 10949 13933 10971 13979
rect 10843 13914 10855 13933
rect 10958 13927 10971 13933
rect 11035 13927 11101 13991
rect 11165 13979 11177 13991
rect 11165 13933 11185 13979
rect 11269 13933 11280 13979
rect 11341 13944 11441 14041
rect 12293 14041 12392 14052
rect 12963 14150 13063 14290
rect 13094 14253 13105 14299
rect 13189 14253 13210 14299
rect 13198 14244 13210 14253
rect 13274 14244 13340 14308
rect 13404 14299 13417 14308
rect 13520 14309 13739 14321
rect 13520 14299 13532 14309
rect 13404 14253 13425 14299
rect 13509 14253 13532 14299
rect 13404 14244 13417 14253
rect 13198 14232 13417 14244
rect 13520 14245 13532 14253
rect 13596 14245 13662 14309
rect 13726 14299 13739 14309
rect 13995 14308 14062 14619
rect 14127 14600 14146 14664
rect 14210 14600 14227 14664
rect 14127 14587 14227 14600
rect 14315 14812 14413 14860
rect 14315 14766 14341 14812
rect 14387 14766 14413 14812
rect 14315 14718 14413 14766
rect 14315 14672 14341 14718
rect 14387 14672 14413 14718
rect 14315 14624 14413 14672
rect 14315 14578 14341 14624
rect 14387 14578 14413 14624
rect 14315 14530 14413 14578
rect 14315 14484 14341 14530
rect 14387 14484 14413 14530
rect 14315 14436 14413 14484
rect 14315 14390 14341 14436
rect 14387 14390 14413 14436
rect 14315 14342 14413 14390
rect 14315 14308 14341 14342
rect 13726 14253 13745 14299
rect 13986 14296 14341 14308
rect 14387 14296 14413 14342
rect 13726 14245 13739 14253
rect 13986 14248 14413 14296
rect 13986 14245 14341 14248
rect 13520 14233 13739 14245
rect 14315 14202 14341 14245
rect 14387 14202 14413 14248
rect 14315 14154 14413 14202
rect 12963 14050 13678 14150
rect 11598 13987 11817 13999
rect 11598 13979 11611 13987
rect 11494 13933 11505 13979
rect 11589 13933 11611 13979
rect 11165 13927 11177 13933
rect 10958 13915 11177 13927
rect 11598 13923 11611 13933
rect 11675 13923 11741 13987
rect 11805 13979 11817 13987
rect 11917 13987 12136 13999
rect 11917 13979 11929 13987
rect 11805 13933 11825 13979
rect 11909 13933 11929 13979
rect 11805 13923 11817 13933
rect 10636 13902 10855 13914
rect 11598 13911 11817 13923
rect 11917 13923 11929 13933
rect 11993 13923 12059 13987
rect 12123 13979 12136 13987
rect 12123 13933 12145 13979
rect 12229 13933 12240 13979
rect 12293 13944 12393 14041
rect 12557 13991 12776 14003
rect 12557 13979 12569 13991
rect 12454 13933 12465 13979
rect 12549 13933 12569 13979
rect 12123 13923 12136 13933
rect 11917 13911 12136 13923
rect 12557 13927 12569 13933
rect 12633 13927 12699 13991
rect 12763 13979 12776 13991
rect 12879 13979 13098 13990
rect 13200 13989 13419 14001
rect 13200 13979 13212 13989
rect 12763 13933 12785 13979
rect 12869 13978 13105 13979
rect 12869 13933 12891 13978
rect 12763 13927 12776 13933
rect 12557 13915 12776 13927
rect 12879 13914 12891 13933
rect 12955 13914 13021 13978
rect 13085 13933 13105 13978
rect 13189 13933 13212 13979
rect 13085 13914 13098 13933
rect 12879 13902 13098 13914
rect 13200 13925 13212 13933
rect 13276 13925 13342 13989
rect 13406 13979 13419 13989
rect 13406 13933 13425 13979
rect 13509 13933 13520 13979
rect 13578 13939 13678 14050
rect 14315 14108 14341 14154
rect 14387 14108 14413 14154
rect 14315 14060 14413 14108
rect 14315 14014 14341 14060
rect 14387 14014 14413 14060
rect 14315 13988 14413 14014
rect 13734 13933 13745 13979
rect 13976 13966 14413 13988
rect 13406 13925 13419 13933
rect 13976 13925 14341 13966
rect 13200 13913 13419 13925
rect 14315 13920 14341 13925
rect 14387 13920 14413 13966
rect 5667 13747 6317 13847
rect 14315 13872 14413 13920
rect 5477 13684 5575 13732
rect 5477 13638 5503 13684
rect 5549 13657 5575 13684
rect 5549 13649 5917 13657
rect 5549 13638 5952 13649
rect 5477 13636 5952 13638
rect 5477 13594 5991 13636
rect 5477 13590 5575 13594
rect 5477 13544 5503 13590
rect 5549 13544 5575 13590
rect 5477 13496 5575 13544
rect 5908 13497 5991 13594
rect 6217 13579 6317 13747
rect 6534 13732 7599 13832
rect 6374 13601 6385 13647
rect 6469 13601 6480 13647
rect 6534 13606 6634 13732
rect 6694 13601 6705 13647
rect 6789 13601 6800 13647
rect 6854 13576 7297 13664
rect 7334 13601 7345 13647
rect 7429 13601 7440 13647
rect 7499 13602 7599 13732
rect 8455 13732 9520 13832
rect 7654 13601 7665 13647
rect 7749 13601 7760 13647
rect 7807 13578 8247 13666
rect 8294 13601 8305 13647
rect 8389 13601 8400 13647
rect 8455 13602 8555 13732
rect 8614 13601 8625 13647
rect 8709 13601 8720 13647
rect 8757 13576 9200 13664
rect 9254 13601 9265 13647
rect 9349 13601 9360 13647
rect 9420 13606 9520 13732
rect 10374 13732 11439 13832
rect 9574 13601 9585 13647
rect 9669 13601 9680 13647
rect 9770 13579 10124 13667
rect 10214 13601 10225 13647
rect 10309 13601 10320 13647
rect 10374 13606 10474 13732
rect 10534 13601 10545 13647
rect 10629 13601 10640 13647
rect 10694 13576 11137 13664
rect 11174 13601 11185 13647
rect 11269 13601 11280 13647
rect 11339 13602 11439 13732
rect 12295 13732 13360 13832
rect 11494 13601 11505 13647
rect 11589 13601 11600 13647
rect 11647 13578 12087 13666
rect 12134 13601 12145 13647
rect 12229 13601 12240 13647
rect 12295 13602 12395 13732
rect 12454 13601 12465 13647
rect 12549 13601 12560 13647
rect 12597 13576 13040 13664
rect 13094 13601 13105 13647
rect 13189 13601 13200 13647
rect 13260 13606 13360 13732
rect 13575 13812 14227 13830
rect 13575 13748 14014 13812
rect 14078 13748 14144 13812
rect 14208 13748 14227 13812
rect 13575 13730 14227 13748
rect 14315 13826 14341 13872
rect 14387 13826 14413 13872
rect 14315 13778 14413 13826
rect 14315 13732 14341 13778
rect 14387 13732 14413 13778
rect 13414 13601 13425 13647
rect 13575 13604 13675 13730
rect 14315 13684 14413 13732
rect 14315 13655 14341 13684
rect 13983 13638 14341 13655
rect 14387 13638 14413 13684
rect 13983 13592 14413 13638
rect 14315 13590 14413 13592
rect 14315 13544 14341 13590
rect 14387 13544 14413 13590
rect 5477 13450 5503 13496
rect 5549 13450 5575 13496
rect 5477 13402 5575 13450
rect 5869 13485 6088 13497
rect 5869 13421 5881 13485
rect 5945 13421 6011 13485
rect 6075 13421 6088 13485
rect 5869 13409 6088 13421
rect 5477 13356 5503 13402
rect 5549 13356 5575 13402
rect 5477 13308 5575 13356
rect 5477 13262 5503 13308
rect 5549 13262 5575 13308
rect 5477 13214 5575 13262
rect 5477 13168 5503 13214
rect 5549 13168 5575 13214
rect 5477 13120 5575 13168
rect 5477 13074 5503 13120
rect 5549 13074 5575 13120
rect 5667 13293 5755 13305
rect 5908 13295 5991 13409
rect 7179 13403 8875 13503
rect 5667 13229 5679 13293
rect 5743 13229 5755 13293
rect 6149 13281 6160 13327
rect 6211 13269 6654 13357
rect 6797 13339 7016 13351
rect 6797 13327 6810 13339
rect 6694 13281 6705 13327
rect 6789 13281 6810 13327
rect 6797 13275 6810 13281
rect 6874 13275 6940 13339
rect 7004 13327 7016 13339
rect 7004 13281 7025 13327
rect 7109 13281 7120 13327
rect 7179 13291 7279 13403
rect 7438 13332 7657 13344
rect 7438 13327 7451 13332
rect 7334 13281 7345 13327
rect 7429 13281 7451 13327
rect 7004 13275 7016 13281
rect 5667 13181 5755 13229
rect 6222 13181 6317 13269
rect 6797 13263 7016 13275
rect 7438 13268 7451 13281
rect 7515 13268 7581 13332
rect 7645 13327 7657 13332
rect 7758 13343 7977 13355
rect 7758 13327 7771 13343
rect 7645 13281 7665 13327
rect 7749 13281 7771 13327
rect 7645 13268 7657 13281
rect 7438 13256 7657 13268
rect 7758 13279 7771 13281
rect 7835 13279 7901 13343
rect 7965 13327 7977 13343
rect 8077 13343 8296 13355
rect 8077 13327 8089 13343
rect 7965 13281 7985 13327
rect 8069 13281 8089 13327
rect 7965 13279 7977 13281
rect 7758 13267 7977 13279
rect 8077 13279 8089 13281
rect 8153 13279 8219 13343
rect 8283 13327 8296 13343
rect 8397 13332 8616 13344
rect 8397 13327 8409 13332
rect 8283 13281 8305 13327
rect 8389 13281 8409 13327
rect 8283 13279 8296 13281
rect 8077 13267 8296 13279
rect 8397 13268 8409 13281
rect 8473 13268 8539 13332
rect 8603 13327 8616 13332
rect 8603 13281 8625 13327
rect 8709 13281 8720 13327
rect 8775 13291 8875 13403
rect 11019 13403 12715 13503
rect 9038 13339 9257 13351
rect 9038 13327 9050 13339
rect 8934 13281 8945 13327
rect 9029 13281 9050 13327
rect 8603 13268 8616 13281
rect 8397 13256 8616 13268
rect 9038 13275 9050 13281
rect 9114 13275 9180 13339
rect 9244 13327 9257 13339
rect 9244 13281 9265 13327
rect 9349 13281 9360 13327
rect 9244 13275 9257 13281
rect 9038 13263 9257 13275
rect 9400 13269 9843 13357
rect 10051 13269 10494 13357
rect 10637 13339 10856 13351
rect 10637 13327 10650 13339
rect 10534 13281 10545 13327
rect 10629 13281 10650 13327
rect 10637 13275 10650 13281
rect 10714 13275 10780 13339
rect 10844 13327 10856 13339
rect 10844 13281 10865 13327
rect 10949 13281 10960 13327
rect 11019 13291 11119 13403
rect 11278 13332 11497 13344
rect 11278 13327 11291 13332
rect 11174 13281 11185 13327
rect 11269 13281 11291 13327
rect 10844 13275 10856 13281
rect 10637 13263 10856 13275
rect 11278 13268 11291 13281
rect 11355 13268 11421 13332
rect 11485 13327 11497 13332
rect 11598 13343 11817 13355
rect 11598 13327 11611 13343
rect 11485 13281 11505 13327
rect 11589 13281 11611 13327
rect 11485 13268 11497 13281
rect 11278 13256 11497 13268
rect 11598 13279 11611 13281
rect 11675 13279 11741 13343
rect 11805 13327 11817 13343
rect 11917 13343 12136 13355
rect 11917 13327 11929 13343
rect 11805 13281 11825 13327
rect 11909 13281 11929 13327
rect 11805 13279 11817 13281
rect 11598 13267 11817 13279
rect 11917 13279 11929 13281
rect 11993 13279 12059 13343
rect 12123 13327 12136 13343
rect 12237 13332 12456 13344
rect 12237 13327 12249 13332
rect 12123 13281 12145 13327
rect 12229 13281 12249 13327
rect 12123 13279 12136 13281
rect 11917 13267 12136 13279
rect 12237 13268 12249 13281
rect 12313 13268 12379 13332
rect 12443 13327 12456 13332
rect 12443 13281 12465 13327
rect 12549 13281 12560 13327
rect 12615 13291 12715 13403
rect 14315 13496 14413 13544
rect 14315 13450 14341 13496
rect 14387 13450 14413 13496
rect 14315 13402 14413 13450
rect 12878 13339 13097 13351
rect 12878 13327 12890 13339
rect 12774 13281 12785 13327
rect 12869 13281 12890 13327
rect 12443 13268 12456 13281
rect 12237 13256 12456 13268
rect 12878 13275 12890 13281
rect 12954 13275 13020 13339
rect 13084 13327 13097 13339
rect 13084 13281 13105 13327
rect 13189 13281 13200 13327
rect 13084 13275 13097 13281
rect 12878 13263 13097 13275
rect 13240 13269 13683 13357
rect 14315 13356 14341 13402
rect 14387 13356 14413 13402
rect 14315 13334 14413 13356
rect 13734 13281 13745 13327
rect 13946 13308 14413 13334
rect 13946 13271 14341 13308
rect 5667 13163 6317 13181
rect 5667 13099 5679 13163
rect 5743 13099 6317 13163
rect 5667 13086 6317 13099
rect 5477 13026 5575 13074
rect 5477 12980 5503 13026
rect 5549 12980 5575 13026
rect 5477 12932 5575 12980
rect 5477 12886 5503 12932
rect 5549 12886 5575 12932
rect 5477 12838 5575 12886
rect 5898 12843 5981 12980
rect 6222 12925 6317 13086
rect 13581 13182 13676 13269
rect 14315 13262 14341 13271
rect 14387 13262 14413 13308
rect 14315 13214 14413 13262
rect 13581 13087 14227 13182
rect 14315 13168 14341 13214
rect 14387 13168 14413 13214
rect 14315 13120 14413 13168
rect 6374 12949 6385 12995
rect 6469 12949 6480 12995
rect 6538 12872 6638 12994
rect 6694 12949 6705 12995
rect 6789 12949 6800 12995
rect 6855 12928 7298 13016
rect 7334 12949 7345 12995
rect 7429 12949 7440 12995
rect 7491 12872 7591 12987
rect 7654 12949 7665 12995
rect 7749 12949 7760 12995
rect 7811 12924 8243 13012
rect 8294 12949 8305 12995
rect 8389 12949 8400 12995
rect 5477 12792 5503 12838
rect 5549 12792 5575 12838
rect 5477 12744 5575 12792
rect 5860 12831 6079 12843
rect 5860 12767 5872 12831
rect 5936 12767 6002 12831
rect 6066 12767 6079 12831
rect 6538 12772 7591 12872
rect 8463 12872 8563 12987
rect 8614 12949 8625 12995
rect 8709 12949 8720 12995
rect 8756 12928 9199 13016
rect 9254 12949 9265 12995
rect 9349 12949 9360 12995
rect 9416 12872 9516 12994
rect 9574 12949 9585 12995
rect 9669 12949 9680 12995
rect 9731 12925 10134 13013
rect 10214 12949 10225 12995
rect 10309 12949 10320 12995
rect 8463 12772 9516 12872
rect 10378 12872 10478 12994
rect 10534 12949 10545 12995
rect 10629 12949 10640 12995
rect 10695 12928 11138 13016
rect 11174 12949 11185 12995
rect 11269 12949 11280 12995
rect 11331 12872 11431 12987
rect 11494 12949 11505 12995
rect 11589 12949 11600 12995
rect 11651 12924 12083 13012
rect 12134 12949 12145 12995
rect 12229 12949 12240 12995
rect 10378 12772 11431 12872
rect 12303 12872 12403 12987
rect 12454 12949 12465 12995
rect 12549 12949 12560 12995
rect 12596 12928 13039 13016
rect 13581 13013 13676 13087
rect 13094 12949 13105 12995
rect 13189 12949 13200 12995
rect 13256 12872 13356 12994
rect 13414 12949 13425 12995
rect 13509 12949 13520 12995
rect 13572 12925 13676 13013
rect 14315 13074 14341 13120
rect 14387 13074 14413 13120
rect 14315 13026 14413 13074
rect 14315 13003 14341 13026
rect 13965 12980 14341 13003
rect 14387 12980 14413 13026
rect 13965 12940 14413 12980
rect 14315 12932 14413 12940
rect 12303 12772 13356 12872
rect 14315 12886 14341 12932
rect 14387 12886 14413 12932
rect 14315 12838 14413 12886
rect 14315 12792 14341 12838
rect 14387 12792 14413 12838
rect 5860 12755 6079 12767
rect 5477 12698 5503 12744
rect 5549 12698 5575 12744
rect 5477 12676 5575 12698
rect 5898 12676 5981 12755
rect 14315 12744 14413 12792
rect 14315 12698 14341 12744
rect 14387 12698 14413 12744
rect 14315 12676 14413 12698
rect 5477 12650 14413 12676
rect 5477 12604 5504 12650
rect 5550 12604 5598 12650
rect 5644 12604 5692 12650
rect 5738 12604 5786 12650
rect 5832 12604 5880 12650
rect 5926 12604 5974 12650
rect 6020 12604 6068 12650
rect 6114 12604 6162 12650
rect 6208 12604 6256 12650
rect 6302 12604 6350 12650
rect 6396 12604 6444 12650
rect 6490 12604 6538 12650
rect 6584 12604 6632 12650
rect 6678 12604 6726 12650
rect 6772 12604 6820 12650
rect 6866 12604 6914 12650
rect 6960 12604 7008 12650
rect 7054 12604 7102 12650
rect 7148 12604 7196 12650
rect 7242 12604 7290 12650
rect 7336 12604 7384 12650
rect 7430 12604 7478 12650
rect 7524 12604 7572 12650
rect 7618 12604 7666 12650
rect 7712 12604 7760 12650
rect 7806 12604 7854 12650
rect 7900 12604 7948 12650
rect 7994 12604 8042 12650
rect 8088 12604 8136 12650
rect 8182 12604 8230 12650
rect 8276 12604 8324 12650
rect 8370 12604 8418 12650
rect 8464 12604 8512 12650
rect 8558 12604 8606 12650
rect 8652 12604 8700 12650
rect 8746 12604 8794 12650
rect 8840 12604 8888 12650
rect 8934 12604 8982 12650
rect 9028 12604 9076 12650
rect 9122 12604 9170 12650
rect 9216 12604 9264 12650
rect 9310 12604 9358 12650
rect 9404 12604 9452 12650
rect 9498 12604 9546 12650
rect 9592 12604 9640 12650
rect 9686 12604 9734 12650
rect 9780 12604 9828 12650
rect 9874 12604 9922 12650
rect 9968 12604 10016 12650
rect 10062 12604 10110 12650
rect 10156 12604 10204 12650
rect 10250 12604 10298 12650
rect 10344 12604 10392 12650
rect 10438 12604 10486 12650
rect 10532 12604 10580 12650
rect 10626 12604 10674 12650
rect 10720 12604 10768 12650
rect 10814 12604 10862 12650
rect 10908 12604 10956 12650
rect 11002 12604 11050 12650
rect 11096 12604 11144 12650
rect 11190 12604 11238 12650
rect 11284 12604 11332 12650
rect 11378 12604 11426 12650
rect 11472 12604 11520 12650
rect 11566 12604 11614 12650
rect 11660 12604 11708 12650
rect 11754 12604 11802 12650
rect 11848 12604 11896 12650
rect 11942 12604 11990 12650
rect 12036 12604 12084 12650
rect 12130 12604 12178 12650
rect 12224 12604 12272 12650
rect 12318 12604 12366 12650
rect 12412 12604 12460 12650
rect 12506 12604 12554 12650
rect 12600 12604 12648 12650
rect 12694 12604 12742 12650
rect 12788 12604 12836 12650
rect 12882 12604 12930 12650
rect 12976 12604 13024 12650
rect 13070 12604 13118 12650
rect 13164 12604 13212 12650
rect 13258 12604 13306 12650
rect 13352 12604 13400 12650
rect 13446 12604 13494 12650
rect 13540 12604 13588 12650
rect 13634 12604 13682 12650
rect 13728 12604 13776 12650
rect 13822 12604 13870 12650
rect 13916 12604 13964 12650
rect 14010 12604 14058 12650
rect 14104 12604 14152 12650
rect 14198 12604 14246 12650
rect 14292 12604 14340 12650
rect 14386 12604 14413 12650
rect 5477 12578 14413 12604
<< via1 >>
rect 5679 14856 5743 14920
rect 7451 15237 7515 15301
rect 7581 15237 7645 15301
rect 8409 15237 8473 15301
rect 8539 15237 8603 15301
rect 11291 15237 11355 15301
rect 11421 15237 11485 15301
rect 12249 15237 12313 15301
rect 12379 15237 12443 15301
rect 6171 14900 6235 14964
rect 6301 14900 6365 14964
rect 6488 14898 6552 14962
rect 6618 14898 6682 14962
rect 9049 14901 9113 14965
rect 9179 14901 9243 14965
rect 9372 14898 9436 14962
rect 9502 14898 9566 14962
rect 9689 14900 9753 14964
rect 9819 14900 9883 14964
rect 10011 14900 10075 14964
rect 10141 14900 10205 14964
rect 10328 14898 10392 14962
rect 10458 14898 10522 14962
rect 10651 14901 10715 14965
rect 10781 14901 10845 14965
rect 5679 14726 5743 14790
rect 12889 14901 12953 14965
rect 13019 14901 13083 14965
rect 13212 14898 13276 14962
rect 13342 14898 13406 14962
rect 13529 14900 13593 14964
rect 13659 14900 13723 14964
rect 14146 14730 14210 14794
rect 6168 14245 6232 14309
rect 6298 14245 6362 14309
rect 6490 14244 6554 14308
rect 6620 14244 6684 14308
rect 7132 14240 7196 14304
rect 7262 14240 7326 14304
rect 7772 14248 7836 14312
rect 7902 14248 7966 14312
rect 8088 14248 8152 14312
rect 8218 14248 8282 14312
rect 13683 14411 13747 14475
rect 13813 14411 13877 14475
rect 8728 14240 8792 14304
rect 8858 14240 8922 14304
rect 5881 14076 5945 14140
rect 6011 14076 6075 14140
rect 6488 13925 6552 13989
rect 6618 13925 6682 13989
rect 6809 13914 6873 13978
rect 6939 13914 7003 13978
rect 7131 13927 7195 13991
rect 7261 13927 7325 13991
rect 9370 14244 9434 14308
rect 9500 14244 9564 14308
rect 9692 14245 9756 14309
rect 9822 14245 9886 14309
rect 10008 14245 10072 14309
rect 10138 14245 10202 14309
rect 10330 14244 10394 14308
rect 10460 14244 10524 14308
rect 10972 14240 11036 14304
rect 11102 14240 11166 14304
rect 11612 14248 11676 14312
rect 11742 14248 11806 14312
rect 11928 14248 11992 14312
rect 12058 14248 12122 14312
rect 12568 14240 12632 14304
rect 12698 14240 12762 14304
rect 7771 13923 7835 13987
rect 7901 13923 7965 13987
rect 8089 13923 8153 13987
rect 8219 13923 8283 13987
rect 8729 13927 8793 13991
rect 8859 13927 8923 13991
rect 9051 13914 9115 13978
rect 9181 13914 9245 13978
rect 9372 13925 9436 13989
rect 9502 13925 9566 13989
rect 10328 13925 10392 13989
rect 10458 13925 10522 13989
rect 10649 13914 10713 13978
rect 10779 13914 10843 13978
rect 10971 13927 11035 13991
rect 11101 13927 11165 13991
rect 13210 14244 13274 14308
rect 13340 14244 13404 14308
rect 13532 14245 13596 14309
rect 13662 14245 13726 14309
rect 14146 14600 14210 14664
rect 11611 13923 11675 13987
rect 11741 13923 11805 13987
rect 11929 13923 11993 13987
rect 12059 13923 12123 13987
rect 12569 13927 12633 13991
rect 12699 13927 12763 13991
rect 12891 13914 12955 13978
rect 13021 13914 13085 13978
rect 13212 13925 13276 13989
rect 13342 13925 13406 13989
rect 14014 13748 14078 13812
rect 14144 13748 14208 13812
rect 5881 13421 5945 13485
rect 6011 13421 6075 13485
rect 5679 13229 5743 13293
rect 6810 13275 6874 13339
rect 6940 13275 7004 13339
rect 7451 13268 7515 13332
rect 7581 13268 7645 13332
rect 7771 13279 7835 13343
rect 7901 13279 7965 13343
rect 8089 13279 8153 13343
rect 8219 13279 8283 13343
rect 8409 13268 8473 13332
rect 8539 13268 8603 13332
rect 9050 13275 9114 13339
rect 9180 13275 9244 13339
rect 10650 13275 10714 13339
rect 10780 13275 10844 13339
rect 11291 13268 11355 13332
rect 11421 13268 11485 13332
rect 11611 13279 11675 13343
rect 11741 13279 11805 13343
rect 11929 13279 11993 13343
rect 12059 13279 12123 13343
rect 12249 13268 12313 13332
rect 12379 13268 12443 13332
rect 12890 13275 12954 13339
rect 13020 13275 13084 13339
rect 5679 13099 5743 13163
rect 5872 12767 5936 12831
rect 6002 12767 6066 12831
<< metal2 >>
rect 9098 15380 10796 15480
rect 7438 15301 7657 15313
rect 7438 15237 7451 15301
rect 7515 15237 7581 15301
rect 7645 15237 7657 15301
rect 7438 15225 7657 15237
rect 8397 15301 8616 15313
rect 8397 15237 8409 15301
rect 8473 15237 8539 15301
rect 8603 15237 8616 15301
rect 8397 15225 8616 15237
rect 9098 14977 9198 15380
rect 10696 14977 10796 15380
rect 11278 15301 11497 15313
rect 11278 15237 11291 15301
rect 11355 15237 11421 15301
rect 11485 15237 11497 15301
rect 11278 15225 11497 15237
rect 12237 15301 12456 15313
rect 12237 15237 12249 15301
rect 12313 15237 12379 15301
rect 12443 15237 12456 15301
rect 12237 15225 12456 15237
rect 12938 15148 13038 15480
rect 12938 15048 13939 15148
rect 12938 14977 13038 15048
rect 6158 14964 6377 14976
rect 5667 14920 5755 14932
rect 5667 14856 5679 14920
rect 5743 14856 5755 14920
rect 6158 14900 6171 14964
rect 6235 14900 6301 14964
rect 6365 14900 6377 14964
rect 6158 14888 6377 14900
rect 6475 14962 6694 14974
rect 6475 14898 6488 14962
rect 6552 14898 6618 14962
rect 6682 14898 6694 14962
rect 5667 14790 5755 14856
rect 5667 14726 5679 14790
rect 5743 14726 5755 14790
rect 5667 13293 5755 14726
rect 6202 14490 6302 14888
rect 6475 14886 6694 14898
rect 9037 14965 9256 14977
rect 9037 14901 9049 14965
rect 9113 14901 9179 14965
rect 9243 14901 9256 14965
rect 9037 14889 9256 14901
rect 9360 14962 9579 14974
rect 9360 14898 9372 14962
rect 9436 14898 9502 14962
rect 9566 14898 9579 14962
rect 9360 14886 9579 14898
rect 9677 14964 9896 14976
rect 9677 14900 9689 14964
rect 9753 14900 9819 14964
rect 9883 14900 9896 14964
rect 9677 14888 9896 14900
rect 9998 14964 10217 14976
rect 9998 14900 10011 14964
rect 10075 14900 10141 14964
rect 10205 14900 10217 14964
rect 9998 14888 10217 14900
rect 10315 14962 10534 14974
rect 10315 14898 10328 14962
rect 10392 14898 10458 14962
rect 10522 14898 10534 14962
rect 6202 14390 6934 14490
rect 6155 14309 6374 14321
rect 6155 14245 6168 14309
rect 6232 14245 6298 14309
rect 6362 14245 6374 14309
rect 6155 14233 6374 14245
rect 6477 14308 6696 14320
rect 6477 14244 6490 14308
rect 6554 14244 6620 14308
rect 6684 14244 6696 14308
rect 5869 14140 6088 14152
rect 5869 14076 5881 14140
rect 5945 14076 6011 14140
rect 6075 14076 6088 14140
rect 5869 14064 6088 14076
rect 5914 13497 6031 14064
rect 6216 13839 6316 14233
rect 6477 14232 6696 14244
rect 6834 14150 6934 14390
rect 7173 14395 7586 14495
rect 7173 14316 7273 14395
rect 7119 14304 7338 14316
rect 7119 14240 7132 14304
rect 7196 14240 7262 14304
rect 7326 14240 7338 14304
rect 7119 14228 7338 14240
rect 6533 14050 6934 14150
rect 7486 14154 7586 14395
rect 8468 14395 8881 14495
rect 9752 14490 9852 14888
rect 7759 14312 7978 14324
rect 7759 14248 7772 14312
rect 7836 14248 7902 14312
rect 7966 14248 7978 14312
rect 7759 14236 7978 14248
rect 8076 14312 8295 14324
rect 8076 14248 8088 14312
rect 8152 14248 8218 14312
rect 8282 14248 8295 14312
rect 8076 14236 8295 14248
rect 8468 14154 8568 14395
rect 8781 14316 8881 14395
rect 9120 14390 9852 14490
rect 10042 14490 10142 14888
rect 10315 14886 10534 14898
rect 10638 14965 10857 14977
rect 10638 14901 10651 14965
rect 10715 14901 10781 14965
rect 10845 14901 10857 14965
rect 10638 14889 10857 14901
rect 12877 14965 13096 14977
rect 12877 14901 12889 14965
rect 12953 14901 13019 14965
rect 13083 14901 13096 14965
rect 12877 14889 13096 14901
rect 13200 14962 13419 14974
rect 13200 14898 13212 14962
rect 13276 14898 13342 14962
rect 13406 14898 13419 14962
rect 13200 14886 13419 14898
rect 13517 14964 13736 14976
rect 13517 14900 13529 14964
rect 13593 14900 13659 14964
rect 13723 14900 13736 14964
rect 13517 14888 13736 14900
rect 13571 14813 13671 14888
rect 13269 14713 13671 14813
rect 10042 14390 10774 14490
rect 8716 14304 8935 14316
rect 8716 14240 8728 14304
rect 8792 14240 8858 14304
rect 8922 14240 8935 14304
rect 8716 14228 8935 14240
rect 7486 14054 7913 14154
rect 6533 14001 6694 14050
rect 6475 13989 6694 14001
rect 7118 13991 7337 14003
rect 6475 13925 6488 13989
rect 6552 13925 6618 13989
rect 6682 13925 6694 13989
rect 6475 13913 6694 13925
rect 6796 13978 7015 13990
rect 6796 13914 6809 13978
rect 6873 13914 6939 13978
rect 7003 13914 7015 13978
rect 7118 13927 7131 13991
rect 7195 13927 7261 13991
rect 7325 13927 7337 13991
rect 7118 13915 7337 13927
rect 7758 13999 7913 14054
rect 8141 14054 8568 14154
rect 9120 14150 9220 14390
rect 9358 14308 9577 14320
rect 9358 14244 9370 14308
rect 9434 14244 9500 14308
rect 9564 14244 9577 14308
rect 9358 14232 9577 14244
rect 9680 14309 9899 14321
rect 9680 14245 9692 14309
rect 9756 14245 9822 14309
rect 9886 14245 9899 14309
rect 9680 14233 9899 14245
rect 9995 14309 10214 14321
rect 9995 14245 10008 14309
rect 10072 14245 10138 14309
rect 10202 14245 10214 14309
rect 9995 14233 10214 14245
rect 10317 14308 10536 14320
rect 10317 14244 10330 14308
rect 10394 14244 10460 14308
rect 10524 14244 10536 14308
rect 8141 13999 8296 14054
rect 9120 14050 9521 14150
rect 7758 13987 7977 13999
rect 7758 13923 7771 13987
rect 7835 13923 7901 13987
rect 7965 13923 7977 13987
rect 6796 13902 7015 13914
rect 6858 13839 6958 13902
rect 6216 13739 6958 13839
rect 7173 13836 7273 13915
rect 7758 13911 7977 13923
rect 8077 13987 8296 13999
rect 8077 13923 8089 13987
rect 8153 13923 8219 13987
rect 8283 13923 8296 13987
rect 8077 13911 8296 13923
rect 8717 13991 8936 14003
rect 8717 13927 8729 13991
rect 8793 13927 8859 13991
rect 8923 13927 8936 13991
rect 9360 14001 9521 14050
rect 8717 13915 8936 13927
rect 9039 13978 9258 13990
rect 8781 13836 8881 13915
rect 9039 13914 9051 13978
rect 9115 13914 9181 13978
rect 9245 13914 9258 13978
rect 9039 13902 9258 13914
rect 9360 13989 9579 14001
rect 9360 13925 9372 13989
rect 9436 13925 9502 13989
rect 9566 13925 9579 13989
rect 9360 13913 9579 13925
rect 7173 13818 7958 13836
rect 7173 13754 7762 13818
rect 7826 13754 7882 13818
rect 7946 13754 7958 13818
rect 7173 13736 7958 13754
rect 8096 13818 8881 13836
rect 8096 13754 8108 13818
rect 8172 13754 8228 13818
rect 8292 13754 8881 13818
rect 8096 13736 8881 13754
rect 9096 13839 9196 13902
rect 9738 13839 9838 14233
rect 9096 13739 9838 13839
rect 10056 13839 10156 14233
rect 10317 14232 10536 14244
rect 10674 14150 10774 14390
rect 11013 14395 11426 14495
rect 11013 14316 11113 14395
rect 10959 14304 11178 14316
rect 10959 14240 10972 14304
rect 11036 14240 11102 14304
rect 11166 14240 11178 14304
rect 10959 14228 11178 14240
rect 10373 14050 10774 14150
rect 11326 14154 11426 14395
rect 12308 14395 12721 14495
rect 13269 14490 13369 14713
rect 13839 14493 13939 15048
rect 11599 14312 11818 14324
rect 11599 14248 11612 14312
rect 11676 14248 11742 14312
rect 11806 14248 11818 14312
rect 11599 14236 11818 14248
rect 11916 14312 12135 14324
rect 11916 14248 11928 14312
rect 11992 14248 12058 14312
rect 12122 14248 12135 14312
rect 11916 14236 12135 14248
rect 12308 14154 12408 14395
rect 12621 14316 12721 14395
rect 12960 14390 13369 14490
rect 13663 14475 13939 14493
rect 13663 14411 13683 14475
rect 13747 14411 13813 14475
rect 13877 14411 13939 14475
rect 13663 14393 13939 14411
rect 14119 14806 14220 14807
rect 14119 14794 14222 14806
rect 14119 14730 14146 14794
rect 14210 14730 14222 14794
rect 14119 14664 14222 14730
rect 14119 14600 14146 14664
rect 14210 14600 14222 14664
rect 14119 14587 14222 14600
rect 12556 14304 12775 14316
rect 12556 14240 12568 14304
rect 12632 14240 12698 14304
rect 12762 14240 12775 14304
rect 12556 14228 12775 14240
rect 11326 14054 11753 14154
rect 10373 14001 10534 14050
rect 10315 13989 10534 14001
rect 10958 13991 11177 14003
rect 10315 13925 10328 13989
rect 10392 13925 10458 13989
rect 10522 13925 10534 13989
rect 10315 13913 10534 13925
rect 10636 13978 10855 13990
rect 10636 13914 10649 13978
rect 10713 13914 10779 13978
rect 10843 13914 10855 13978
rect 10958 13927 10971 13991
rect 11035 13927 11101 13991
rect 11165 13927 11177 13991
rect 10958 13915 11177 13927
rect 11598 13999 11753 14054
rect 11981 14054 12408 14154
rect 12960 14150 13060 14390
rect 13198 14308 13417 14320
rect 13198 14244 13210 14308
rect 13274 14244 13340 14308
rect 13404 14244 13417 14308
rect 13198 14232 13417 14244
rect 13520 14309 13739 14321
rect 13520 14245 13532 14309
rect 13596 14245 13662 14309
rect 13726 14245 13739 14309
rect 13520 14233 13739 14245
rect 11981 13999 12136 14054
rect 12960 14050 13361 14150
rect 11598 13987 11817 13999
rect 11598 13923 11611 13987
rect 11675 13923 11741 13987
rect 11805 13923 11817 13987
rect 10636 13902 10855 13914
rect 10698 13839 10798 13902
rect 10056 13739 10798 13839
rect 11013 13836 11113 13915
rect 11598 13911 11817 13923
rect 11917 13987 12136 13999
rect 11917 13923 11929 13987
rect 11993 13923 12059 13987
rect 12123 13923 12136 13987
rect 11917 13911 12136 13923
rect 12557 13991 12776 14003
rect 12557 13927 12569 13991
rect 12633 13927 12699 13991
rect 12763 13927 12776 13991
rect 13200 14001 13361 14050
rect 12557 13915 12776 13927
rect 12879 13978 13098 13990
rect 12621 13836 12721 13915
rect 12879 13914 12891 13978
rect 12955 13914 13021 13978
rect 13085 13914 13098 13978
rect 12879 13902 13098 13914
rect 13200 13989 13419 14001
rect 13200 13925 13212 13989
rect 13276 13925 13342 13989
rect 13406 13925 13419 13989
rect 13200 13913 13419 13925
rect 11013 13818 11798 13836
rect 11013 13754 11602 13818
rect 11666 13754 11722 13818
rect 11786 13754 11798 13818
rect 11013 13736 11798 13754
rect 11936 13818 12721 13836
rect 11936 13754 11948 13818
rect 12012 13754 12068 13818
rect 12132 13754 12721 13818
rect 11936 13736 12721 13754
rect 12936 13839 13036 13902
rect 13578 13839 13678 14233
rect 12936 13739 13678 13839
rect 14119 13824 14220 14587
rect 14001 13812 14220 13824
rect 14001 13748 14014 13812
rect 14078 13748 14144 13812
rect 14208 13748 14220 13812
rect 14001 13736 14220 13748
rect 5869 13485 6088 13497
rect 5869 13421 5881 13485
rect 5945 13421 6011 13485
rect 6075 13421 6088 13485
rect 5869 13409 6088 13421
rect 5667 13229 5679 13293
rect 5743 13229 5755 13293
rect 5667 13163 5755 13229
rect 5667 13099 5679 13163
rect 5743 13099 5755 13163
rect 5667 13086 5755 13099
rect 5914 12843 6031 13409
rect 6797 13339 7016 13351
rect 6797 13275 6810 13339
rect 6874 13275 6940 13339
rect 7004 13275 7016 13339
rect 6797 13263 7016 13275
rect 7438 13332 7657 13344
rect 7438 13268 7451 13332
rect 7515 13268 7581 13332
rect 7645 13268 7657 13332
rect 7438 13256 7657 13268
rect 7758 13343 7977 13355
rect 7758 13279 7771 13343
rect 7835 13279 7901 13343
rect 7965 13279 7977 13343
rect 7758 13267 7977 13279
rect 8077 13343 8296 13355
rect 8077 13279 8089 13343
rect 8153 13279 8219 13343
rect 8283 13279 8296 13343
rect 8077 13267 8296 13279
rect 8397 13332 8616 13344
rect 8397 13268 8409 13332
rect 8473 13268 8539 13332
rect 8603 13268 8616 13332
rect 8397 13256 8616 13268
rect 9038 13339 9257 13351
rect 9038 13275 9050 13339
rect 9114 13275 9180 13339
rect 9244 13275 9257 13339
rect 9038 13263 9257 13275
rect 10637 13339 10856 13351
rect 10637 13275 10650 13339
rect 10714 13275 10780 13339
rect 10844 13275 10856 13339
rect 10637 13263 10856 13275
rect 11278 13332 11497 13344
rect 11278 13268 11291 13332
rect 11355 13268 11421 13332
rect 11485 13268 11497 13332
rect 11278 13256 11497 13268
rect 11598 13343 11817 13355
rect 11598 13279 11611 13343
rect 11675 13279 11741 13343
rect 11805 13279 11817 13343
rect 11598 13267 11817 13279
rect 11917 13343 12136 13355
rect 11917 13279 11929 13343
rect 11993 13279 12059 13343
rect 12123 13279 12136 13343
rect 11917 13267 12136 13279
rect 12237 13332 12456 13344
rect 12237 13268 12249 13332
rect 12313 13268 12379 13332
rect 12443 13268 12456 13332
rect 12237 13256 12456 13268
rect 12878 13339 13097 13351
rect 12878 13275 12890 13339
rect 12954 13275 13020 13339
rect 13084 13275 13097 13339
rect 12878 13263 13097 13275
rect 5860 12831 6079 12843
rect 5860 12767 5872 12831
rect 5936 12767 6002 12831
rect 6066 12767 6079 12831
rect 5860 12755 6079 12767
<< via2 >>
rect 7451 15237 7515 15301
rect 7581 15237 7645 15301
rect 8409 15237 8473 15301
rect 8539 15237 8603 15301
rect 11291 15237 11355 15301
rect 11421 15237 11485 15301
rect 12249 15237 12313 15301
rect 12379 15237 12443 15301
rect 6488 14898 6552 14962
rect 6618 14898 6682 14962
rect 9372 14898 9436 14962
rect 9502 14898 9566 14962
rect 10328 14898 10392 14962
rect 10458 14898 10522 14962
rect 6490 14244 6554 14308
rect 6620 14244 6684 14308
rect 7772 14248 7836 14312
rect 7902 14248 7966 14312
rect 8088 14248 8152 14312
rect 8218 14248 8282 14312
rect 13212 14898 13276 14962
rect 13342 14898 13406 14962
rect 9370 14244 9434 14308
rect 9500 14244 9564 14308
rect 10330 14244 10394 14308
rect 10460 14244 10524 14308
rect 7762 13754 7826 13818
rect 7882 13754 7946 13818
rect 8108 13754 8172 13818
rect 8228 13754 8292 13818
rect 11612 14248 11676 14312
rect 11742 14248 11806 14312
rect 11928 14248 11992 14312
rect 12058 14248 12122 14312
rect 13210 14244 13274 14308
rect 13340 14244 13404 14308
rect 11602 13754 11666 13818
rect 11722 13754 11786 13818
rect 11948 13754 12012 13818
rect 12068 13754 12132 13818
rect 6810 13275 6874 13339
rect 6940 13275 7004 13339
rect 7451 13268 7515 13332
rect 7581 13268 7645 13332
rect 7771 13279 7835 13343
rect 7901 13279 7965 13343
rect 8089 13279 8153 13343
rect 8219 13279 8283 13343
rect 8409 13268 8473 13332
rect 8539 13268 8603 13332
rect 9050 13275 9114 13339
rect 9180 13275 9244 13339
rect 10650 13275 10714 13339
rect 10780 13275 10844 13339
rect 11291 13268 11355 13332
rect 11421 13268 11485 13332
rect 11611 13279 11675 13343
rect 11741 13279 11805 13343
rect 11929 13279 11993 13343
rect 12059 13279 12123 13343
rect 12249 13268 12313 13332
rect 12379 13268 12443 13332
rect 12890 13275 12954 13339
rect 13020 13275 13084 13339
<< metal3 >>
rect 7438 15301 7657 15313
rect 7438 15237 7451 15301
rect 7515 15237 7581 15301
rect 7645 15237 7657 15301
rect 7438 15225 7657 15237
rect 8397 15301 8616 15313
rect 8397 15237 8409 15301
rect 8473 15237 8539 15301
rect 8603 15237 8616 15301
rect 8397 15225 8616 15237
rect 11278 15301 11497 15313
rect 11278 15237 11291 15301
rect 11355 15237 11421 15301
rect 11485 15237 11497 15301
rect 11278 15225 11497 15237
rect 12237 15301 12456 15313
rect 12237 15237 12249 15301
rect 12313 15237 12379 15301
rect 12443 15237 12456 15301
rect 12237 15225 12456 15237
rect 6475 14962 6694 14974
rect 6475 14898 6488 14962
rect 6552 14898 6618 14962
rect 6682 14898 6694 14962
rect 6475 14886 6694 14898
rect 6515 14806 6615 14886
rect 6515 14706 7275 14806
rect 6477 14308 6696 14320
rect 6477 14244 6490 14308
rect 6554 14244 6620 14308
rect 6684 14244 6696 14308
rect 6477 14232 6696 14244
rect 6533 14171 6633 14232
rect 6533 14071 6956 14171
rect 6856 13351 6956 14071
rect 6797 13339 7016 13351
rect 6797 13275 6810 13339
rect 6874 13275 6940 13339
rect 7004 13275 7016 13339
rect 6797 13263 7016 13275
rect 7175 13199 7275 14706
rect 7494 13344 7594 15225
rect 7759 14312 7978 14324
rect 7759 14248 7772 14312
rect 7836 14248 7902 14312
rect 7966 14248 7978 14312
rect 7759 14236 7978 14248
rect 8076 14312 8295 14324
rect 8076 14248 8088 14312
rect 8152 14248 8218 14312
rect 8282 14248 8295 14312
rect 8076 14236 8295 14248
rect 7808 13836 7908 14236
rect 8146 13836 8246 14236
rect 7749 13818 7958 13836
rect 7749 13754 7762 13818
rect 7826 13754 7882 13818
rect 7946 13754 7958 13818
rect 7749 13736 7958 13754
rect 8096 13818 8305 13836
rect 8096 13754 8108 13818
rect 8172 13754 8228 13818
rect 8292 13754 8305 13818
rect 8096 13736 8305 13754
rect 7438 13332 7657 13344
rect 7438 13268 7451 13332
rect 7515 13268 7581 13332
rect 7645 13268 7657 13332
rect 7438 13256 7657 13268
rect 7758 13343 7977 13355
rect 7758 13279 7771 13343
rect 7835 13279 7901 13343
rect 7965 13279 7977 13343
rect 7758 13267 7977 13279
rect 8077 13343 8296 13355
rect 8460 13344 8560 15225
rect 9360 14962 9579 14974
rect 9360 14898 9372 14962
rect 9436 14898 9502 14962
rect 9566 14898 9579 14962
rect 9360 14886 9579 14898
rect 10315 14962 10534 14974
rect 10315 14898 10328 14962
rect 10392 14898 10458 14962
rect 10522 14898 10534 14962
rect 10315 14886 10534 14898
rect 9439 14806 9539 14886
rect 8779 14706 9539 14806
rect 10355 14806 10455 14886
rect 10355 14706 11115 14806
rect 8077 13279 8089 13343
rect 8153 13279 8219 13343
rect 8283 13279 8296 13343
rect 8077 13267 8296 13279
rect 8397 13332 8616 13344
rect 8397 13268 8409 13332
rect 8473 13268 8539 13332
rect 8603 13268 8616 13332
rect 7806 13199 7906 13267
rect 7175 13099 7906 13199
rect 8148 13199 8248 13267
rect 8397 13256 8616 13268
rect 8779 13199 8879 14706
rect 9358 14308 9577 14320
rect 9358 14244 9370 14308
rect 9434 14244 9500 14308
rect 9564 14244 9577 14308
rect 9358 14232 9577 14244
rect 10317 14308 10536 14320
rect 10317 14244 10330 14308
rect 10394 14244 10460 14308
rect 10524 14244 10536 14308
rect 10317 14232 10536 14244
rect 9421 14171 9521 14232
rect 9098 14071 9521 14171
rect 10373 14171 10473 14232
rect 10373 14071 10796 14171
rect 9098 13351 9198 14071
rect 10696 13351 10796 14071
rect 9038 13339 9257 13351
rect 9038 13275 9050 13339
rect 9114 13275 9180 13339
rect 9244 13275 9257 13339
rect 9038 13263 9257 13275
rect 10637 13339 10856 13351
rect 10637 13275 10650 13339
rect 10714 13275 10780 13339
rect 10844 13275 10856 13339
rect 10637 13263 10856 13275
rect 8148 13099 8879 13199
rect 11015 13199 11115 14706
rect 11334 13344 11434 15225
rect 11599 14312 11818 14324
rect 11599 14248 11612 14312
rect 11676 14248 11742 14312
rect 11806 14248 11818 14312
rect 11599 14236 11818 14248
rect 11916 14312 12135 14324
rect 11916 14248 11928 14312
rect 11992 14248 12058 14312
rect 12122 14248 12135 14312
rect 11916 14236 12135 14248
rect 11648 13836 11748 14236
rect 11986 13836 12086 14236
rect 11589 13818 11798 13836
rect 11589 13754 11602 13818
rect 11666 13754 11722 13818
rect 11786 13754 11798 13818
rect 11589 13736 11798 13754
rect 11936 13818 12145 13836
rect 11936 13754 11948 13818
rect 12012 13754 12068 13818
rect 12132 13754 12145 13818
rect 11936 13736 12145 13754
rect 11278 13332 11497 13344
rect 11278 13268 11291 13332
rect 11355 13268 11421 13332
rect 11485 13268 11497 13332
rect 11278 13256 11497 13268
rect 11598 13343 11817 13355
rect 11598 13279 11611 13343
rect 11675 13279 11741 13343
rect 11805 13279 11817 13343
rect 11598 13267 11817 13279
rect 11917 13343 12136 13355
rect 12300 13344 12400 15225
rect 13200 14962 13419 14974
rect 13200 14898 13212 14962
rect 13276 14898 13342 14962
rect 13406 14898 13419 14962
rect 13200 14886 13419 14898
rect 13279 14806 13379 14886
rect 12619 14706 13379 14806
rect 11917 13279 11929 13343
rect 11993 13279 12059 13343
rect 12123 13279 12136 13343
rect 11917 13267 12136 13279
rect 12237 13332 12456 13344
rect 12237 13268 12249 13332
rect 12313 13268 12379 13332
rect 12443 13268 12456 13332
rect 11646 13199 11746 13267
rect 11015 13099 11746 13199
rect 11988 13199 12088 13267
rect 12237 13256 12456 13268
rect 12619 13199 12719 14706
rect 13198 14308 13417 14320
rect 13198 14244 13210 14308
rect 13274 14244 13340 14308
rect 13404 14244 13417 14308
rect 13198 14232 13417 14244
rect 13261 14171 13361 14232
rect 12938 14071 13361 14171
rect 12938 13351 13038 14071
rect 12878 13339 13097 13351
rect 12878 13275 12890 13339
rect 12954 13275 13020 13339
rect 13084 13275 13097 13339
rect 12878 13263 13097 13275
rect 11988 13099 12719 13199
use ppolyf_u_W5AMT6  ppolyf_u_W5AMT6_0
timestamp 1694513024
transform 1 0 9947 0 1 13138
box -4304 -386 4304 386
use ppolyf_u_W5AMT6  ppolyf_u_W5AMT6_1
timestamp 1694513024
transform 1 0 9947 0 1 15094
box -4304 -386 4304 386
use ppolyf_u_W5AMT6  ppolyf_u_W5AMT6_2
timestamp 1694513024
transform 1 0 9947 0 1 14442
box -4304 -386 4304 386
use ppolyf_u_W5AMT6  ppolyf_u_W5AMT6_3
timestamp 1694513024
transform 1 0 9947 0 1 13790
box -4304 -386 4304 386
<< labels >>
flabel metal1 6263 15330 6263 15330 0 FreeSans 1600 0 0 0 A
port 1 nsew
flabel metal1 13459 15339 13459 15339 0 FreeSans 1600 0 0 0 B
port 3 nsew
flabel metal1 6588 15339 6588 15339 0 FreeSans 1600 0 0 0 C
port 5 nsew
flabel metal2 12986 15349 12986 15349 0 FreeSans 1600 0 0 0 D
port 7 nsew
flabel metal1 5746 14447 5746 14447 0 FreeSans 1600 0 0 0 E
port 9 nsew
flabel metal1 14122 14758 14122 14758 0 FreeSans 1600 0 0 0 F
port 10 nsew
flabel metal1 5794 14766 5794 14766 0 FreeSans 1600 0 0 0 G
port 14 nsew
flabel metal1 14151 13143 14151 13143 0 FreeSans 1600 0 0 0 H
port 15 nsew
flabel metal1 5938 15580 5938 15580 0 FreeSans 1600 0 0 0 VDD
port 16 nsew
<< end >>
