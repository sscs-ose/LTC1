magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1046 -2396 1046 2396
<< metal1 >>
rect -46 1390 46 1396
rect -46 1364 -40 1390
rect -14 1364 14 1390
rect 40 1364 46 1390
rect -46 1336 46 1364
rect -46 1310 -40 1336
rect -14 1310 14 1336
rect 40 1310 46 1336
rect -46 1282 46 1310
rect -46 1256 -40 1282
rect -14 1256 14 1282
rect 40 1256 46 1282
rect -46 1228 46 1256
rect -46 1202 -40 1228
rect -14 1202 14 1228
rect 40 1202 46 1228
rect -46 1174 46 1202
rect -46 1148 -40 1174
rect -14 1148 14 1174
rect 40 1148 46 1174
rect -46 1120 46 1148
rect -46 1094 -40 1120
rect -14 1094 14 1120
rect 40 1094 46 1120
rect -46 1066 46 1094
rect -46 1040 -40 1066
rect -14 1040 14 1066
rect 40 1040 46 1066
rect -46 1012 46 1040
rect -46 986 -40 1012
rect -14 986 14 1012
rect 40 986 46 1012
rect -46 958 46 986
rect -46 932 -40 958
rect -14 932 14 958
rect 40 932 46 958
rect -46 904 46 932
rect -46 878 -40 904
rect -14 878 14 904
rect 40 878 46 904
rect -46 850 46 878
rect -46 824 -40 850
rect -14 824 14 850
rect 40 824 46 850
rect -46 796 46 824
rect -46 770 -40 796
rect -14 770 14 796
rect 40 770 46 796
rect -46 742 46 770
rect -46 716 -40 742
rect -14 716 14 742
rect 40 716 46 742
rect -46 688 46 716
rect -46 662 -40 688
rect -14 662 14 688
rect 40 662 46 688
rect -46 634 46 662
rect -46 608 -40 634
rect -14 608 14 634
rect 40 608 46 634
rect -46 580 46 608
rect -46 554 -40 580
rect -14 554 14 580
rect 40 554 46 580
rect -46 526 46 554
rect -46 500 -40 526
rect -14 500 14 526
rect 40 500 46 526
rect -46 472 46 500
rect -46 446 -40 472
rect -14 446 14 472
rect 40 446 46 472
rect -46 418 46 446
rect -46 392 -40 418
rect -14 392 14 418
rect 40 392 46 418
rect -46 364 46 392
rect -46 338 -40 364
rect -14 338 14 364
rect 40 338 46 364
rect -46 310 46 338
rect -46 284 -40 310
rect -14 284 14 310
rect 40 284 46 310
rect -46 256 46 284
rect -46 230 -40 256
rect -14 230 14 256
rect 40 230 46 256
rect -46 202 46 230
rect -46 176 -40 202
rect -14 176 14 202
rect 40 176 46 202
rect -46 148 46 176
rect -46 122 -40 148
rect -14 122 14 148
rect 40 122 46 148
rect -46 94 46 122
rect -46 68 -40 94
rect -14 68 14 94
rect 40 68 46 94
rect -46 40 46 68
rect -46 14 -40 40
rect -14 14 14 40
rect 40 14 46 40
rect -46 -14 46 14
rect -46 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 46 -14
rect -46 -68 46 -40
rect -46 -94 -40 -68
rect -14 -94 14 -68
rect 40 -94 46 -68
rect -46 -122 46 -94
rect -46 -148 -40 -122
rect -14 -148 14 -122
rect 40 -148 46 -122
rect -46 -176 46 -148
rect -46 -202 -40 -176
rect -14 -202 14 -176
rect 40 -202 46 -176
rect -46 -230 46 -202
rect -46 -256 -40 -230
rect -14 -256 14 -230
rect 40 -256 46 -230
rect -46 -284 46 -256
rect -46 -310 -40 -284
rect -14 -310 14 -284
rect 40 -310 46 -284
rect -46 -338 46 -310
rect -46 -364 -40 -338
rect -14 -364 14 -338
rect 40 -364 46 -338
rect -46 -392 46 -364
rect -46 -418 -40 -392
rect -14 -418 14 -392
rect 40 -418 46 -392
rect -46 -446 46 -418
rect -46 -472 -40 -446
rect -14 -472 14 -446
rect 40 -472 46 -446
rect -46 -500 46 -472
rect -46 -526 -40 -500
rect -14 -526 14 -500
rect 40 -526 46 -500
rect -46 -554 46 -526
rect -46 -580 -40 -554
rect -14 -580 14 -554
rect 40 -580 46 -554
rect -46 -608 46 -580
rect -46 -634 -40 -608
rect -14 -634 14 -608
rect 40 -634 46 -608
rect -46 -662 46 -634
rect -46 -688 -40 -662
rect -14 -688 14 -662
rect 40 -688 46 -662
rect -46 -716 46 -688
rect -46 -742 -40 -716
rect -14 -742 14 -716
rect 40 -742 46 -716
rect -46 -770 46 -742
rect -46 -796 -40 -770
rect -14 -796 14 -770
rect 40 -796 46 -770
rect -46 -824 46 -796
rect -46 -850 -40 -824
rect -14 -850 14 -824
rect 40 -850 46 -824
rect -46 -878 46 -850
rect -46 -904 -40 -878
rect -14 -904 14 -878
rect 40 -904 46 -878
rect -46 -932 46 -904
rect -46 -958 -40 -932
rect -14 -958 14 -932
rect 40 -958 46 -932
rect -46 -986 46 -958
rect -46 -1012 -40 -986
rect -14 -1012 14 -986
rect 40 -1012 46 -986
rect -46 -1040 46 -1012
rect -46 -1066 -40 -1040
rect -14 -1066 14 -1040
rect 40 -1066 46 -1040
rect -46 -1094 46 -1066
rect -46 -1120 -40 -1094
rect -14 -1120 14 -1094
rect 40 -1120 46 -1094
rect -46 -1148 46 -1120
rect -46 -1174 -40 -1148
rect -14 -1174 14 -1148
rect 40 -1174 46 -1148
rect -46 -1202 46 -1174
rect -46 -1228 -40 -1202
rect -14 -1228 14 -1202
rect 40 -1228 46 -1202
rect -46 -1256 46 -1228
rect -46 -1282 -40 -1256
rect -14 -1282 14 -1256
rect 40 -1282 46 -1256
rect -46 -1310 46 -1282
rect -46 -1336 -40 -1310
rect -14 -1336 14 -1310
rect 40 -1336 46 -1310
rect -46 -1364 46 -1336
rect -46 -1390 -40 -1364
rect -14 -1390 14 -1364
rect 40 -1390 46 -1364
rect -46 -1396 46 -1390
<< via1 >>
rect -40 1364 -14 1390
rect 14 1364 40 1390
rect -40 1310 -14 1336
rect 14 1310 40 1336
rect -40 1256 -14 1282
rect 14 1256 40 1282
rect -40 1202 -14 1228
rect 14 1202 40 1228
rect -40 1148 -14 1174
rect 14 1148 40 1174
rect -40 1094 -14 1120
rect 14 1094 40 1120
rect -40 1040 -14 1066
rect 14 1040 40 1066
rect -40 986 -14 1012
rect 14 986 40 1012
rect -40 932 -14 958
rect 14 932 40 958
rect -40 878 -14 904
rect 14 878 40 904
rect -40 824 -14 850
rect 14 824 40 850
rect -40 770 -14 796
rect 14 770 40 796
rect -40 716 -14 742
rect 14 716 40 742
rect -40 662 -14 688
rect 14 662 40 688
rect -40 608 -14 634
rect 14 608 40 634
rect -40 554 -14 580
rect 14 554 40 580
rect -40 500 -14 526
rect 14 500 40 526
rect -40 446 -14 472
rect 14 446 40 472
rect -40 392 -14 418
rect 14 392 40 418
rect -40 338 -14 364
rect 14 338 40 364
rect -40 284 -14 310
rect 14 284 40 310
rect -40 230 -14 256
rect 14 230 40 256
rect -40 176 -14 202
rect 14 176 40 202
rect -40 122 -14 148
rect 14 122 40 148
rect -40 68 -14 94
rect 14 68 40 94
rect -40 14 -14 40
rect 14 14 40 40
rect -40 -40 -14 -14
rect 14 -40 40 -14
rect -40 -94 -14 -68
rect 14 -94 40 -68
rect -40 -148 -14 -122
rect 14 -148 40 -122
rect -40 -202 -14 -176
rect 14 -202 40 -176
rect -40 -256 -14 -230
rect 14 -256 40 -230
rect -40 -310 -14 -284
rect 14 -310 40 -284
rect -40 -364 -14 -338
rect 14 -364 40 -338
rect -40 -418 -14 -392
rect 14 -418 40 -392
rect -40 -472 -14 -446
rect 14 -472 40 -446
rect -40 -526 -14 -500
rect 14 -526 40 -500
rect -40 -580 -14 -554
rect 14 -580 40 -554
rect -40 -634 -14 -608
rect 14 -634 40 -608
rect -40 -688 -14 -662
rect 14 -688 40 -662
rect -40 -742 -14 -716
rect 14 -742 40 -716
rect -40 -796 -14 -770
rect 14 -796 40 -770
rect -40 -850 -14 -824
rect 14 -850 40 -824
rect -40 -904 -14 -878
rect 14 -904 40 -878
rect -40 -958 -14 -932
rect 14 -958 40 -932
rect -40 -1012 -14 -986
rect 14 -1012 40 -986
rect -40 -1066 -14 -1040
rect 14 -1066 40 -1040
rect -40 -1120 -14 -1094
rect 14 -1120 40 -1094
rect -40 -1174 -14 -1148
rect 14 -1174 40 -1148
rect -40 -1228 -14 -1202
rect 14 -1228 40 -1202
rect -40 -1282 -14 -1256
rect 14 -1282 40 -1256
rect -40 -1336 -14 -1310
rect 14 -1336 40 -1310
rect -40 -1390 -14 -1364
rect 14 -1390 40 -1364
<< metal2 >>
rect -46 1390 46 1396
rect -46 1364 -40 1390
rect -14 1364 14 1390
rect 40 1364 46 1390
rect -46 1336 46 1364
rect -46 1310 -40 1336
rect -14 1310 14 1336
rect 40 1310 46 1336
rect -46 1282 46 1310
rect -46 1256 -40 1282
rect -14 1256 14 1282
rect 40 1256 46 1282
rect -46 1228 46 1256
rect -46 1202 -40 1228
rect -14 1202 14 1228
rect 40 1202 46 1228
rect -46 1174 46 1202
rect -46 1148 -40 1174
rect -14 1148 14 1174
rect 40 1148 46 1174
rect -46 1120 46 1148
rect -46 1094 -40 1120
rect -14 1094 14 1120
rect 40 1094 46 1120
rect -46 1066 46 1094
rect -46 1040 -40 1066
rect -14 1040 14 1066
rect 40 1040 46 1066
rect -46 1012 46 1040
rect -46 986 -40 1012
rect -14 986 14 1012
rect 40 986 46 1012
rect -46 958 46 986
rect -46 932 -40 958
rect -14 932 14 958
rect 40 932 46 958
rect -46 904 46 932
rect -46 878 -40 904
rect -14 878 14 904
rect 40 878 46 904
rect -46 850 46 878
rect -46 824 -40 850
rect -14 824 14 850
rect 40 824 46 850
rect -46 796 46 824
rect -46 770 -40 796
rect -14 770 14 796
rect 40 770 46 796
rect -46 742 46 770
rect -46 716 -40 742
rect -14 716 14 742
rect 40 716 46 742
rect -46 688 46 716
rect -46 662 -40 688
rect -14 662 14 688
rect 40 662 46 688
rect -46 634 46 662
rect -46 608 -40 634
rect -14 608 14 634
rect 40 608 46 634
rect -46 580 46 608
rect -46 554 -40 580
rect -14 554 14 580
rect 40 554 46 580
rect -46 526 46 554
rect -46 500 -40 526
rect -14 500 14 526
rect 40 500 46 526
rect -46 472 46 500
rect -46 446 -40 472
rect -14 446 14 472
rect 40 446 46 472
rect -46 418 46 446
rect -46 392 -40 418
rect -14 392 14 418
rect 40 392 46 418
rect -46 364 46 392
rect -46 338 -40 364
rect -14 338 14 364
rect 40 338 46 364
rect -46 310 46 338
rect -46 284 -40 310
rect -14 284 14 310
rect 40 284 46 310
rect -46 256 46 284
rect -46 230 -40 256
rect -14 230 14 256
rect 40 230 46 256
rect -46 202 46 230
rect -46 176 -40 202
rect -14 176 14 202
rect 40 176 46 202
rect -46 148 46 176
rect -46 122 -40 148
rect -14 122 14 148
rect 40 122 46 148
rect -46 94 46 122
rect -46 68 -40 94
rect -14 68 14 94
rect 40 68 46 94
rect -46 40 46 68
rect -46 14 -40 40
rect -14 14 14 40
rect 40 14 46 40
rect -46 -14 46 14
rect -46 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 46 -14
rect -46 -68 46 -40
rect -46 -94 -40 -68
rect -14 -94 14 -68
rect 40 -94 46 -68
rect -46 -122 46 -94
rect -46 -148 -40 -122
rect -14 -148 14 -122
rect 40 -148 46 -122
rect -46 -176 46 -148
rect -46 -202 -40 -176
rect -14 -202 14 -176
rect 40 -202 46 -176
rect -46 -230 46 -202
rect -46 -256 -40 -230
rect -14 -256 14 -230
rect 40 -256 46 -230
rect -46 -284 46 -256
rect -46 -310 -40 -284
rect -14 -310 14 -284
rect 40 -310 46 -284
rect -46 -338 46 -310
rect -46 -364 -40 -338
rect -14 -364 14 -338
rect 40 -364 46 -338
rect -46 -392 46 -364
rect -46 -418 -40 -392
rect -14 -418 14 -392
rect 40 -418 46 -392
rect -46 -446 46 -418
rect -46 -472 -40 -446
rect -14 -472 14 -446
rect 40 -472 46 -446
rect -46 -500 46 -472
rect -46 -526 -40 -500
rect -14 -526 14 -500
rect 40 -526 46 -500
rect -46 -554 46 -526
rect -46 -580 -40 -554
rect -14 -580 14 -554
rect 40 -580 46 -554
rect -46 -608 46 -580
rect -46 -634 -40 -608
rect -14 -634 14 -608
rect 40 -634 46 -608
rect -46 -662 46 -634
rect -46 -688 -40 -662
rect -14 -688 14 -662
rect 40 -688 46 -662
rect -46 -716 46 -688
rect -46 -742 -40 -716
rect -14 -742 14 -716
rect 40 -742 46 -716
rect -46 -770 46 -742
rect -46 -796 -40 -770
rect -14 -796 14 -770
rect 40 -796 46 -770
rect -46 -824 46 -796
rect -46 -850 -40 -824
rect -14 -850 14 -824
rect 40 -850 46 -824
rect -46 -878 46 -850
rect -46 -904 -40 -878
rect -14 -904 14 -878
rect 40 -904 46 -878
rect -46 -932 46 -904
rect -46 -958 -40 -932
rect -14 -958 14 -932
rect 40 -958 46 -932
rect -46 -986 46 -958
rect -46 -1012 -40 -986
rect -14 -1012 14 -986
rect 40 -1012 46 -986
rect -46 -1040 46 -1012
rect -46 -1066 -40 -1040
rect -14 -1066 14 -1040
rect 40 -1066 46 -1040
rect -46 -1094 46 -1066
rect -46 -1120 -40 -1094
rect -14 -1120 14 -1094
rect 40 -1120 46 -1094
rect -46 -1148 46 -1120
rect -46 -1174 -40 -1148
rect -14 -1174 14 -1148
rect 40 -1174 46 -1148
rect -46 -1202 46 -1174
rect -46 -1228 -40 -1202
rect -14 -1228 14 -1202
rect 40 -1228 46 -1202
rect -46 -1256 46 -1228
rect -46 -1282 -40 -1256
rect -14 -1282 14 -1256
rect 40 -1282 46 -1256
rect -46 -1310 46 -1282
rect -46 -1336 -40 -1310
rect -14 -1336 14 -1310
rect 40 -1336 46 -1310
rect -46 -1364 46 -1336
rect -46 -1390 -40 -1364
rect -14 -1390 14 -1364
rect 40 -1390 46 -1364
rect -46 -1396 46 -1390
<< end >>
