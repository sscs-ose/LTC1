magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1143 -1267 1143 1267
<< metal1 >>
rect -143 261 143 267
rect -143 235 -137 261
rect -111 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 111 261
rect 137 235 143 261
rect -143 199 143 235
rect -143 173 -137 199
rect -111 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 111 199
rect 137 173 143 199
rect -143 137 143 173
rect -143 111 -137 137
rect -111 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 111 137
rect 137 111 143 137
rect -143 75 143 111
rect -143 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 143 75
rect -143 13 143 49
rect -143 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 143 13
rect -143 -49 143 -13
rect -143 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 143 -49
rect -143 -111 143 -75
rect -143 -137 -137 -111
rect -111 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 111 -111
rect 137 -137 143 -111
rect -143 -173 143 -137
rect -143 -199 -137 -173
rect -111 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 111 -173
rect 137 -199 143 -173
rect -143 -235 143 -199
rect -143 -261 -137 -235
rect -111 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 111 -235
rect 137 -261 143 -235
rect -143 -267 143 -261
<< via1 >>
rect -137 235 -111 261
rect -75 235 -49 261
rect -13 235 13 261
rect 49 235 75 261
rect 111 235 137 261
rect -137 173 -111 199
rect -75 173 -49 199
rect -13 173 13 199
rect 49 173 75 199
rect 111 173 137 199
rect -137 111 -111 137
rect -75 111 -49 137
rect -13 111 13 137
rect 49 111 75 137
rect 111 111 137 137
rect -137 49 -111 75
rect -75 49 -49 75
rect -13 49 13 75
rect 49 49 75 75
rect 111 49 137 75
rect -137 -13 -111 13
rect -75 -13 -49 13
rect -13 -13 13 13
rect 49 -13 75 13
rect 111 -13 137 13
rect -137 -75 -111 -49
rect -75 -75 -49 -49
rect -13 -75 13 -49
rect 49 -75 75 -49
rect 111 -75 137 -49
rect -137 -137 -111 -111
rect -75 -137 -49 -111
rect -13 -137 13 -111
rect 49 -137 75 -111
rect 111 -137 137 -111
rect -137 -199 -111 -173
rect -75 -199 -49 -173
rect -13 -199 13 -173
rect 49 -199 75 -173
rect 111 -199 137 -173
rect -137 -261 -111 -235
rect -75 -261 -49 -235
rect -13 -261 13 -235
rect 49 -261 75 -235
rect 111 -261 137 -235
<< metal2 >>
rect -143 261 143 267
rect -143 235 -137 261
rect -111 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 111 261
rect 137 235 143 261
rect -143 199 143 235
rect -143 173 -137 199
rect -111 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 111 199
rect 137 173 143 199
rect -143 137 143 173
rect -143 111 -137 137
rect -111 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 111 137
rect 137 111 143 137
rect -143 75 143 111
rect -143 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 143 75
rect -143 13 143 49
rect -143 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 143 13
rect -143 -49 143 -13
rect -143 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 143 -49
rect -143 -111 143 -75
rect -143 -137 -137 -111
rect -111 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 111 -111
rect 137 -137 143 -111
rect -143 -173 143 -137
rect -143 -199 -137 -173
rect -111 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 111 -173
rect 137 -199 143 -173
rect -143 -235 143 -199
rect -143 -261 -137 -235
rect -111 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 111 -235
rect 137 -261 143 -235
rect -143 -267 143 -261
<< end >>
