** sch_path: /home/shahid/GF180Projects/Top_test/Decoder_muxes/Xschem/8x1_mux_PEX_TB_ibr..sym
**.subckt 8x1_mux_PEX_TB_ibr.
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V4 S0 VSS pulse(3.3 0 0 100p 100p 100n 200n)
.save i(v4)
V5 S1 VSS pulse(3.3 0 0 100p 100p 200n 400n)
.save i(v5)
V6 I0 VSS 3.3
.save i(v6)
V7 I1 VSS 0
.save i(v7)
V8 I2 VSS 3.3
.save i(v8)
V9 I3 VSS 0
.save i(v9)
V10 I5 VSS 0
.save i(v10)
V11 I4 VSS 3.3
.save i(v11)
V12 I6 VSS 3.3
.save i(v12)
V13 I7 VSS 0
.save i(v13)
V14 S2 VSS pulse(3.3 0 0 100p 100p 400n 800n)
.save i(v14)
x1 VDD VSS S1 S0 OUT S2 I0 I7 I3 I2 I5 I1 I4 I6 pex_mux_8x1_ibr
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_mux_8x1_ibr.spice
.control
save all
tran 50p 800n
plot v(S0) v(S1)+3.5 v(S2)+7 v(I0)+10.5 v(I1)+14 v(I2)+17.5
plot v(I3) v(I4)+4.5 v(I5)+8 v(I6)+11.5 v(I7)+15
plot v(OUT)



*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
