magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -8008 -2115 8008 2115
<< metal4 >>
rect -6002 99 6002 109
rect -6002 43 -5992 99
rect -5936 43 -5850 99
rect -5794 43 -5708 99
rect -5652 43 -5566 99
rect -5510 43 -5424 99
rect -5368 43 -5282 99
rect -5226 43 -5140 99
rect -5084 43 -4998 99
rect -4942 43 -4856 99
rect -4800 43 -4714 99
rect -4658 43 -4572 99
rect -4516 43 -4430 99
rect -4374 43 -4288 99
rect -4232 43 -4146 99
rect -4090 43 -4004 99
rect -3948 43 -3862 99
rect -3806 43 -3720 99
rect -3664 43 -3578 99
rect -3522 43 -3436 99
rect -3380 43 -3294 99
rect -3238 43 -3152 99
rect -3096 43 -3010 99
rect -2954 43 -2868 99
rect -2812 43 -2726 99
rect -2670 43 -2584 99
rect -2528 43 -2442 99
rect -2386 43 -2300 99
rect -2244 43 -2158 99
rect -2102 43 -2016 99
rect -1960 43 -1874 99
rect -1818 43 -1732 99
rect -1676 43 -1590 99
rect -1534 43 -1448 99
rect -1392 43 -1306 99
rect -1250 43 -1164 99
rect -1108 43 -1022 99
rect -966 43 -880 99
rect -824 43 -738 99
rect -682 43 -596 99
rect -540 43 -454 99
rect -398 43 -312 99
rect -256 43 -170 99
rect -114 43 -28 99
rect 28 43 114 99
rect 170 43 256 99
rect 312 43 398 99
rect 454 43 540 99
rect 596 43 682 99
rect 738 43 824 99
rect 880 43 966 99
rect 1022 43 1108 99
rect 1164 43 1250 99
rect 1306 43 1392 99
rect 1448 43 1534 99
rect 1590 43 1676 99
rect 1732 43 1818 99
rect 1874 43 1960 99
rect 2016 43 2102 99
rect 2158 43 2244 99
rect 2300 43 2386 99
rect 2442 43 2528 99
rect 2584 43 2670 99
rect 2726 43 2812 99
rect 2868 43 2954 99
rect 3010 43 3096 99
rect 3152 43 3238 99
rect 3294 43 3380 99
rect 3436 43 3522 99
rect 3578 43 3664 99
rect 3720 43 3806 99
rect 3862 43 3948 99
rect 4004 43 4090 99
rect 4146 43 4232 99
rect 4288 43 4374 99
rect 4430 43 4516 99
rect 4572 43 4658 99
rect 4714 43 4800 99
rect 4856 43 4942 99
rect 4998 43 5084 99
rect 5140 43 5226 99
rect 5282 43 5368 99
rect 5424 43 5510 99
rect 5566 43 5652 99
rect 5708 43 5794 99
rect 5850 43 5936 99
rect 5992 43 6002 99
rect -6002 -43 6002 43
rect -6002 -99 -5992 -43
rect -5936 -99 -5850 -43
rect -5794 -99 -5708 -43
rect -5652 -99 -5566 -43
rect -5510 -99 -5424 -43
rect -5368 -99 -5282 -43
rect -5226 -99 -5140 -43
rect -5084 -99 -4998 -43
rect -4942 -99 -4856 -43
rect -4800 -99 -4714 -43
rect -4658 -99 -4572 -43
rect -4516 -99 -4430 -43
rect -4374 -99 -4288 -43
rect -4232 -99 -4146 -43
rect -4090 -99 -4004 -43
rect -3948 -99 -3862 -43
rect -3806 -99 -3720 -43
rect -3664 -99 -3578 -43
rect -3522 -99 -3436 -43
rect -3380 -99 -3294 -43
rect -3238 -99 -3152 -43
rect -3096 -99 -3010 -43
rect -2954 -99 -2868 -43
rect -2812 -99 -2726 -43
rect -2670 -99 -2584 -43
rect -2528 -99 -2442 -43
rect -2386 -99 -2300 -43
rect -2244 -99 -2158 -43
rect -2102 -99 -2016 -43
rect -1960 -99 -1874 -43
rect -1818 -99 -1732 -43
rect -1676 -99 -1590 -43
rect -1534 -99 -1448 -43
rect -1392 -99 -1306 -43
rect -1250 -99 -1164 -43
rect -1108 -99 -1022 -43
rect -966 -99 -880 -43
rect -824 -99 -738 -43
rect -682 -99 -596 -43
rect -540 -99 -454 -43
rect -398 -99 -312 -43
rect -256 -99 -170 -43
rect -114 -99 -28 -43
rect 28 -99 114 -43
rect 170 -99 256 -43
rect 312 -99 398 -43
rect 454 -99 540 -43
rect 596 -99 682 -43
rect 738 -99 824 -43
rect 880 -99 966 -43
rect 1022 -99 1108 -43
rect 1164 -99 1250 -43
rect 1306 -99 1392 -43
rect 1448 -99 1534 -43
rect 1590 -99 1676 -43
rect 1732 -99 1818 -43
rect 1874 -99 1960 -43
rect 2016 -99 2102 -43
rect 2158 -99 2244 -43
rect 2300 -99 2386 -43
rect 2442 -99 2528 -43
rect 2584 -99 2670 -43
rect 2726 -99 2812 -43
rect 2868 -99 2954 -43
rect 3010 -99 3096 -43
rect 3152 -99 3238 -43
rect 3294 -99 3380 -43
rect 3436 -99 3522 -43
rect 3578 -99 3664 -43
rect 3720 -99 3806 -43
rect 3862 -99 3948 -43
rect 4004 -99 4090 -43
rect 4146 -99 4232 -43
rect 4288 -99 4374 -43
rect 4430 -99 4516 -43
rect 4572 -99 4658 -43
rect 4714 -99 4800 -43
rect 4856 -99 4942 -43
rect 4998 -99 5084 -43
rect 5140 -99 5226 -43
rect 5282 -99 5368 -43
rect 5424 -99 5510 -43
rect 5566 -99 5652 -43
rect 5708 -99 5794 -43
rect 5850 -99 5936 -43
rect 5992 -99 6002 -43
rect -6002 -109 6002 -99
<< via4 >>
rect -5992 43 -5936 99
rect -5850 43 -5794 99
rect -5708 43 -5652 99
rect -5566 43 -5510 99
rect -5424 43 -5368 99
rect -5282 43 -5226 99
rect -5140 43 -5084 99
rect -4998 43 -4942 99
rect -4856 43 -4800 99
rect -4714 43 -4658 99
rect -4572 43 -4516 99
rect -4430 43 -4374 99
rect -4288 43 -4232 99
rect -4146 43 -4090 99
rect -4004 43 -3948 99
rect -3862 43 -3806 99
rect -3720 43 -3664 99
rect -3578 43 -3522 99
rect -3436 43 -3380 99
rect -3294 43 -3238 99
rect -3152 43 -3096 99
rect -3010 43 -2954 99
rect -2868 43 -2812 99
rect -2726 43 -2670 99
rect -2584 43 -2528 99
rect -2442 43 -2386 99
rect -2300 43 -2244 99
rect -2158 43 -2102 99
rect -2016 43 -1960 99
rect -1874 43 -1818 99
rect -1732 43 -1676 99
rect -1590 43 -1534 99
rect -1448 43 -1392 99
rect -1306 43 -1250 99
rect -1164 43 -1108 99
rect -1022 43 -966 99
rect -880 43 -824 99
rect -738 43 -682 99
rect -596 43 -540 99
rect -454 43 -398 99
rect -312 43 -256 99
rect -170 43 -114 99
rect -28 43 28 99
rect 114 43 170 99
rect 256 43 312 99
rect 398 43 454 99
rect 540 43 596 99
rect 682 43 738 99
rect 824 43 880 99
rect 966 43 1022 99
rect 1108 43 1164 99
rect 1250 43 1306 99
rect 1392 43 1448 99
rect 1534 43 1590 99
rect 1676 43 1732 99
rect 1818 43 1874 99
rect 1960 43 2016 99
rect 2102 43 2158 99
rect 2244 43 2300 99
rect 2386 43 2442 99
rect 2528 43 2584 99
rect 2670 43 2726 99
rect 2812 43 2868 99
rect 2954 43 3010 99
rect 3096 43 3152 99
rect 3238 43 3294 99
rect 3380 43 3436 99
rect 3522 43 3578 99
rect 3664 43 3720 99
rect 3806 43 3862 99
rect 3948 43 4004 99
rect 4090 43 4146 99
rect 4232 43 4288 99
rect 4374 43 4430 99
rect 4516 43 4572 99
rect 4658 43 4714 99
rect 4800 43 4856 99
rect 4942 43 4998 99
rect 5084 43 5140 99
rect 5226 43 5282 99
rect 5368 43 5424 99
rect 5510 43 5566 99
rect 5652 43 5708 99
rect 5794 43 5850 99
rect 5936 43 5992 99
rect -5992 -99 -5936 -43
rect -5850 -99 -5794 -43
rect -5708 -99 -5652 -43
rect -5566 -99 -5510 -43
rect -5424 -99 -5368 -43
rect -5282 -99 -5226 -43
rect -5140 -99 -5084 -43
rect -4998 -99 -4942 -43
rect -4856 -99 -4800 -43
rect -4714 -99 -4658 -43
rect -4572 -99 -4516 -43
rect -4430 -99 -4374 -43
rect -4288 -99 -4232 -43
rect -4146 -99 -4090 -43
rect -4004 -99 -3948 -43
rect -3862 -99 -3806 -43
rect -3720 -99 -3664 -43
rect -3578 -99 -3522 -43
rect -3436 -99 -3380 -43
rect -3294 -99 -3238 -43
rect -3152 -99 -3096 -43
rect -3010 -99 -2954 -43
rect -2868 -99 -2812 -43
rect -2726 -99 -2670 -43
rect -2584 -99 -2528 -43
rect -2442 -99 -2386 -43
rect -2300 -99 -2244 -43
rect -2158 -99 -2102 -43
rect -2016 -99 -1960 -43
rect -1874 -99 -1818 -43
rect -1732 -99 -1676 -43
rect -1590 -99 -1534 -43
rect -1448 -99 -1392 -43
rect -1306 -99 -1250 -43
rect -1164 -99 -1108 -43
rect -1022 -99 -966 -43
rect -880 -99 -824 -43
rect -738 -99 -682 -43
rect -596 -99 -540 -43
rect -454 -99 -398 -43
rect -312 -99 -256 -43
rect -170 -99 -114 -43
rect -28 -99 28 -43
rect 114 -99 170 -43
rect 256 -99 312 -43
rect 398 -99 454 -43
rect 540 -99 596 -43
rect 682 -99 738 -43
rect 824 -99 880 -43
rect 966 -99 1022 -43
rect 1108 -99 1164 -43
rect 1250 -99 1306 -43
rect 1392 -99 1448 -43
rect 1534 -99 1590 -43
rect 1676 -99 1732 -43
rect 1818 -99 1874 -43
rect 1960 -99 2016 -43
rect 2102 -99 2158 -43
rect 2244 -99 2300 -43
rect 2386 -99 2442 -43
rect 2528 -99 2584 -43
rect 2670 -99 2726 -43
rect 2812 -99 2868 -43
rect 2954 -99 3010 -43
rect 3096 -99 3152 -43
rect 3238 -99 3294 -43
rect 3380 -99 3436 -43
rect 3522 -99 3578 -43
rect 3664 -99 3720 -43
rect 3806 -99 3862 -43
rect 3948 -99 4004 -43
rect 4090 -99 4146 -43
rect 4232 -99 4288 -43
rect 4374 -99 4430 -43
rect 4516 -99 4572 -43
rect 4658 -99 4714 -43
rect 4800 -99 4856 -43
rect 4942 -99 4998 -43
rect 5084 -99 5140 -43
rect 5226 -99 5282 -43
rect 5368 -99 5424 -43
rect 5510 -99 5566 -43
rect 5652 -99 5708 -43
rect 5794 -99 5850 -43
rect 5936 -99 5992 -43
<< metal5 >>
rect -6008 99 6008 115
rect -6008 43 -5992 99
rect -5936 43 -5850 99
rect -5794 43 -5708 99
rect -5652 43 -5566 99
rect -5510 43 -5424 99
rect -5368 43 -5282 99
rect -5226 43 -5140 99
rect -5084 43 -4998 99
rect -4942 43 -4856 99
rect -4800 43 -4714 99
rect -4658 43 -4572 99
rect -4516 43 -4430 99
rect -4374 43 -4288 99
rect -4232 43 -4146 99
rect -4090 43 -4004 99
rect -3948 43 -3862 99
rect -3806 43 -3720 99
rect -3664 43 -3578 99
rect -3522 43 -3436 99
rect -3380 43 -3294 99
rect -3238 43 -3152 99
rect -3096 43 -3010 99
rect -2954 43 -2868 99
rect -2812 43 -2726 99
rect -2670 43 -2584 99
rect -2528 43 -2442 99
rect -2386 43 -2300 99
rect -2244 43 -2158 99
rect -2102 43 -2016 99
rect -1960 43 -1874 99
rect -1818 43 -1732 99
rect -1676 43 -1590 99
rect -1534 43 -1448 99
rect -1392 43 -1306 99
rect -1250 43 -1164 99
rect -1108 43 -1022 99
rect -966 43 -880 99
rect -824 43 -738 99
rect -682 43 -596 99
rect -540 43 -454 99
rect -398 43 -312 99
rect -256 43 -170 99
rect -114 43 -28 99
rect 28 43 114 99
rect 170 43 256 99
rect 312 43 398 99
rect 454 43 540 99
rect 596 43 682 99
rect 738 43 824 99
rect 880 43 966 99
rect 1022 43 1108 99
rect 1164 43 1250 99
rect 1306 43 1392 99
rect 1448 43 1534 99
rect 1590 43 1676 99
rect 1732 43 1818 99
rect 1874 43 1960 99
rect 2016 43 2102 99
rect 2158 43 2244 99
rect 2300 43 2386 99
rect 2442 43 2528 99
rect 2584 43 2670 99
rect 2726 43 2812 99
rect 2868 43 2954 99
rect 3010 43 3096 99
rect 3152 43 3238 99
rect 3294 43 3380 99
rect 3436 43 3522 99
rect 3578 43 3664 99
rect 3720 43 3806 99
rect 3862 43 3948 99
rect 4004 43 4090 99
rect 4146 43 4232 99
rect 4288 43 4374 99
rect 4430 43 4516 99
rect 4572 43 4658 99
rect 4714 43 4800 99
rect 4856 43 4942 99
rect 4998 43 5084 99
rect 5140 43 5226 99
rect 5282 43 5368 99
rect 5424 43 5510 99
rect 5566 43 5652 99
rect 5708 43 5794 99
rect 5850 43 5936 99
rect 5992 43 6008 99
rect -6008 -43 6008 43
rect -6008 -99 -5992 -43
rect -5936 -99 -5850 -43
rect -5794 -99 -5708 -43
rect -5652 -99 -5566 -43
rect -5510 -99 -5424 -43
rect -5368 -99 -5282 -43
rect -5226 -99 -5140 -43
rect -5084 -99 -4998 -43
rect -4942 -99 -4856 -43
rect -4800 -99 -4714 -43
rect -4658 -99 -4572 -43
rect -4516 -99 -4430 -43
rect -4374 -99 -4288 -43
rect -4232 -99 -4146 -43
rect -4090 -99 -4004 -43
rect -3948 -99 -3862 -43
rect -3806 -99 -3720 -43
rect -3664 -99 -3578 -43
rect -3522 -99 -3436 -43
rect -3380 -99 -3294 -43
rect -3238 -99 -3152 -43
rect -3096 -99 -3010 -43
rect -2954 -99 -2868 -43
rect -2812 -99 -2726 -43
rect -2670 -99 -2584 -43
rect -2528 -99 -2442 -43
rect -2386 -99 -2300 -43
rect -2244 -99 -2158 -43
rect -2102 -99 -2016 -43
rect -1960 -99 -1874 -43
rect -1818 -99 -1732 -43
rect -1676 -99 -1590 -43
rect -1534 -99 -1448 -43
rect -1392 -99 -1306 -43
rect -1250 -99 -1164 -43
rect -1108 -99 -1022 -43
rect -966 -99 -880 -43
rect -824 -99 -738 -43
rect -682 -99 -596 -43
rect -540 -99 -454 -43
rect -398 -99 -312 -43
rect -256 -99 -170 -43
rect -114 -99 -28 -43
rect 28 -99 114 -43
rect 170 -99 256 -43
rect 312 -99 398 -43
rect 454 -99 540 -43
rect 596 -99 682 -43
rect 738 -99 824 -43
rect 880 -99 966 -43
rect 1022 -99 1108 -43
rect 1164 -99 1250 -43
rect 1306 -99 1392 -43
rect 1448 -99 1534 -43
rect 1590 -99 1676 -43
rect 1732 -99 1818 -43
rect 1874 -99 1960 -43
rect 2016 -99 2102 -43
rect 2158 -99 2244 -43
rect 2300 -99 2386 -43
rect 2442 -99 2528 -43
rect 2584 -99 2670 -43
rect 2726 -99 2812 -43
rect 2868 -99 2954 -43
rect 3010 -99 3096 -43
rect 3152 -99 3238 -43
rect 3294 -99 3380 -43
rect 3436 -99 3522 -43
rect 3578 -99 3664 -43
rect 3720 -99 3806 -43
rect 3862 -99 3948 -43
rect 4004 -99 4090 -43
rect 4146 -99 4232 -43
rect 4288 -99 4374 -43
rect 4430 -99 4516 -43
rect 4572 -99 4658 -43
rect 4714 -99 4800 -43
rect 4856 -99 4942 -43
rect 4998 -99 5084 -43
rect 5140 -99 5226 -43
rect 5282 -99 5368 -43
rect 5424 -99 5510 -43
rect 5566 -99 5652 -43
rect 5708 -99 5794 -43
rect 5850 -99 5936 -43
rect 5992 -99 6008 -43
rect -6008 -115 6008 -99
<< end >>
