magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1329 -1019 1329 1019
<< metal2 >>
rect -329 14 329 19
rect -329 -14 -324 14
rect -296 -14 -262 14
rect -234 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 234 14
rect 262 -14 296 14
rect 324 -14 329 14
rect -329 -19 329 -14
<< via2 >>
rect -324 -14 -296 14
rect -262 -14 -234 14
rect -200 -14 -172 14
rect -138 -14 -110 14
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect 110 -14 138 14
rect 172 -14 200 14
rect 234 -14 262 14
rect 296 -14 324 14
<< metal3 >>
rect -329 14 329 19
rect -329 -14 -324 14
rect -296 -14 -262 14
rect -234 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 234 14
rect 262 -14 296 14
rect 324 -14 329 14
rect -329 -19 329 -14
<< end >>
