magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1349 -3230 1349 3230
<< metal3 >>
rect -349 2225 349 2230
rect -349 2197 -344 2225
rect -316 2197 -278 2225
rect -250 2197 -212 2225
rect -184 2197 -146 2225
rect -118 2197 -80 2225
rect -52 2197 -14 2225
rect 14 2197 52 2225
rect 80 2197 118 2225
rect 146 2197 184 2225
rect 212 2197 250 2225
rect 278 2197 316 2225
rect 344 2197 349 2225
rect -349 2159 349 2197
rect -349 2131 -344 2159
rect -316 2131 -278 2159
rect -250 2131 -212 2159
rect -184 2131 -146 2159
rect -118 2131 -80 2159
rect -52 2131 -14 2159
rect 14 2131 52 2159
rect 80 2131 118 2159
rect 146 2131 184 2159
rect 212 2131 250 2159
rect 278 2131 316 2159
rect 344 2131 349 2159
rect -349 2093 349 2131
rect -349 2065 -344 2093
rect -316 2065 -278 2093
rect -250 2065 -212 2093
rect -184 2065 -146 2093
rect -118 2065 -80 2093
rect -52 2065 -14 2093
rect 14 2065 52 2093
rect 80 2065 118 2093
rect 146 2065 184 2093
rect 212 2065 250 2093
rect 278 2065 316 2093
rect 344 2065 349 2093
rect -349 2027 349 2065
rect -349 1999 -344 2027
rect -316 1999 -278 2027
rect -250 1999 -212 2027
rect -184 1999 -146 2027
rect -118 1999 -80 2027
rect -52 1999 -14 2027
rect 14 1999 52 2027
rect 80 1999 118 2027
rect 146 1999 184 2027
rect 212 1999 250 2027
rect 278 1999 316 2027
rect 344 1999 349 2027
rect -349 1961 349 1999
rect -349 1933 -344 1961
rect -316 1933 -278 1961
rect -250 1933 -212 1961
rect -184 1933 -146 1961
rect -118 1933 -80 1961
rect -52 1933 -14 1961
rect 14 1933 52 1961
rect 80 1933 118 1961
rect 146 1933 184 1961
rect 212 1933 250 1961
rect 278 1933 316 1961
rect 344 1933 349 1961
rect -349 1895 349 1933
rect -349 1867 -344 1895
rect -316 1867 -278 1895
rect -250 1867 -212 1895
rect -184 1867 -146 1895
rect -118 1867 -80 1895
rect -52 1867 -14 1895
rect 14 1867 52 1895
rect 80 1867 118 1895
rect 146 1867 184 1895
rect 212 1867 250 1895
rect 278 1867 316 1895
rect 344 1867 349 1895
rect -349 1829 349 1867
rect -349 1801 -344 1829
rect -316 1801 -278 1829
rect -250 1801 -212 1829
rect -184 1801 -146 1829
rect -118 1801 -80 1829
rect -52 1801 -14 1829
rect 14 1801 52 1829
rect 80 1801 118 1829
rect 146 1801 184 1829
rect 212 1801 250 1829
rect 278 1801 316 1829
rect 344 1801 349 1829
rect -349 1763 349 1801
rect -349 1735 -344 1763
rect -316 1735 -278 1763
rect -250 1735 -212 1763
rect -184 1735 -146 1763
rect -118 1735 -80 1763
rect -52 1735 -14 1763
rect 14 1735 52 1763
rect 80 1735 118 1763
rect 146 1735 184 1763
rect 212 1735 250 1763
rect 278 1735 316 1763
rect 344 1735 349 1763
rect -349 1697 349 1735
rect -349 1669 -344 1697
rect -316 1669 -278 1697
rect -250 1669 -212 1697
rect -184 1669 -146 1697
rect -118 1669 -80 1697
rect -52 1669 -14 1697
rect 14 1669 52 1697
rect 80 1669 118 1697
rect 146 1669 184 1697
rect 212 1669 250 1697
rect 278 1669 316 1697
rect 344 1669 349 1697
rect -349 1631 349 1669
rect -349 1603 -344 1631
rect -316 1603 -278 1631
rect -250 1603 -212 1631
rect -184 1603 -146 1631
rect -118 1603 -80 1631
rect -52 1603 -14 1631
rect 14 1603 52 1631
rect 80 1603 118 1631
rect 146 1603 184 1631
rect 212 1603 250 1631
rect 278 1603 316 1631
rect 344 1603 349 1631
rect -349 1565 349 1603
rect -349 1537 -344 1565
rect -316 1537 -278 1565
rect -250 1537 -212 1565
rect -184 1537 -146 1565
rect -118 1537 -80 1565
rect -52 1537 -14 1565
rect 14 1537 52 1565
rect 80 1537 118 1565
rect 146 1537 184 1565
rect 212 1537 250 1565
rect 278 1537 316 1565
rect 344 1537 349 1565
rect -349 1499 349 1537
rect -349 1471 -344 1499
rect -316 1471 -278 1499
rect -250 1471 -212 1499
rect -184 1471 -146 1499
rect -118 1471 -80 1499
rect -52 1471 -14 1499
rect 14 1471 52 1499
rect 80 1471 118 1499
rect 146 1471 184 1499
rect 212 1471 250 1499
rect 278 1471 316 1499
rect 344 1471 349 1499
rect -349 1433 349 1471
rect -349 1405 -344 1433
rect -316 1405 -278 1433
rect -250 1405 -212 1433
rect -184 1405 -146 1433
rect -118 1405 -80 1433
rect -52 1405 -14 1433
rect 14 1405 52 1433
rect 80 1405 118 1433
rect 146 1405 184 1433
rect 212 1405 250 1433
rect 278 1405 316 1433
rect 344 1405 349 1433
rect -349 1367 349 1405
rect -349 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 349 1367
rect -349 1301 349 1339
rect -349 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 349 1301
rect -349 1235 349 1273
rect -349 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 349 1235
rect -349 1169 349 1207
rect -349 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 349 1169
rect -349 1103 349 1141
rect -349 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 349 1103
rect -349 1037 349 1075
rect -349 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 349 1037
rect -349 971 349 1009
rect -349 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 349 971
rect -349 905 349 943
rect -349 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 349 905
rect -349 839 349 877
rect -349 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 349 839
rect -349 773 349 811
rect -349 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 349 773
rect -349 707 349 745
rect -349 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 349 707
rect -349 641 349 679
rect -349 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 349 641
rect -349 575 349 613
rect -349 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 349 575
rect -349 509 349 547
rect -349 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 349 509
rect -349 443 349 481
rect -349 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 349 443
rect -349 377 349 415
rect -349 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 349 377
rect -349 311 349 349
rect -349 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 349 311
rect -349 245 349 283
rect -349 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 349 245
rect -349 179 349 217
rect -349 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 349 179
rect -349 113 349 151
rect -349 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 349 113
rect -349 47 349 85
rect -349 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 349 47
rect -349 -19 349 19
rect -349 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 349 -19
rect -349 -85 349 -47
rect -349 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 349 -85
rect -349 -151 349 -113
rect -349 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 349 -151
rect -349 -217 349 -179
rect -349 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 349 -217
rect -349 -283 349 -245
rect -349 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 349 -283
rect -349 -349 349 -311
rect -349 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 349 -349
rect -349 -415 349 -377
rect -349 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 349 -415
rect -349 -481 349 -443
rect -349 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 349 -481
rect -349 -547 349 -509
rect -349 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 349 -547
rect -349 -613 349 -575
rect -349 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 349 -613
rect -349 -679 349 -641
rect -349 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 349 -679
rect -349 -745 349 -707
rect -349 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 349 -745
rect -349 -811 349 -773
rect -349 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 349 -811
rect -349 -877 349 -839
rect -349 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 349 -877
rect -349 -943 349 -905
rect -349 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 349 -943
rect -349 -1009 349 -971
rect -349 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 349 -1009
rect -349 -1075 349 -1037
rect -349 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 349 -1075
rect -349 -1141 349 -1103
rect -349 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 349 -1141
rect -349 -1207 349 -1169
rect -349 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 349 -1207
rect -349 -1273 349 -1235
rect -349 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 349 -1273
rect -349 -1339 349 -1301
rect -349 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 349 -1339
rect -349 -1405 349 -1367
rect -349 -1433 -344 -1405
rect -316 -1433 -278 -1405
rect -250 -1433 -212 -1405
rect -184 -1433 -146 -1405
rect -118 -1433 -80 -1405
rect -52 -1433 -14 -1405
rect 14 -1433 52 -1405
rect 80 -1433 118 -1405
rect 146 -1433 184 -1405
rect 212 -1433 250 -1405
rect 278 -1433 316 -1405
rect 344 -1433 349 -1405
rect -349 -1471 349 -1433
rect -349 -1499 -344 -1471
rect -316 -1499 -278 -1471
rect -250 -1499 -212 -1471
rect -184 -1499 -146 -1471
rect -118 -1499 -80 -1471
rect -52 -1499 -14 -1471
rect 14 -1499 52 -1471
rect 80 -1499 118 -1471
rect 146 -1499 184 -1471
rect 212 -1499 250 -1471
rect 278 -1499 316 -1471
rect 344 -1499 349 -1471
rect -349 -1537 349 -1499
rect -349 -1565 -344 -1537
rect -316 -1565 -278 -1537
rect -250 -1565 -212 -1537
rect -184 -1565 -146 -1537
rect -118 -1565 -80 -1537
rect -52 -1565 -14 -1537
rect 14 -1565 52 -1537
rect 80 -1565 118 -1537
rect 146 -1565 184 -1537
rect 212 -1565 250 -1537
rect 278 -1565 316 -1537
rect 344 -1565 349 -1537
rect -349 -1603 349 -1565
rect -349 -1631 -344 -1603
rect -316 -1631 -278 -1603
rect -250 -1631 -212 -1603
rect -184 -1631 -146 -1603
rect -118 -1631 -80 -1603
rect -52 -1631 -14 -1603
rect 14 -1631 52 -1603
rect 80 -1631 118 -1603
rect 146 -1631 184 -1603
rect 212 -1631 250 -1603
rect 278 -1631 316 -1603
rect 344 -1631 349 -1603
rect -349 -1669 349 -1631
rect -349 -1697 -344 -1669
rect -316 -1697 -278 -1669
rect -250 -1697 -212 -1669
rect -184 -1697 -146 -1669
rect -118 -1697 -80 -1669
rect -52 -1697 -14 -1669
rect 14 -1697 52 -1669
rect 80 -1697 118 -1669
rect 146 -1697 184 -1669
rect 212 -1697 250 -1669
rect 278 -1697 316 -1669
rect 344 -1697 349 -1669
rect -349 -1735 349 -1697
rect -349 -1763 -344 -1735
rect -316 -1763 -278 -1735
rect -250 -1763 -212 -1735
rect -184 -1763 -146 -1735
rect -118 -1763 -80 -1735
rect -52 -1763 -14 -1735
rect 14 -1763 52 -1735
rect 80 -1763 118 -1735
rect 146 -1763 184 -1735
rect 212 -1763 250 -1735
rect 278 -1763 316 -1735
rect 344 -1763 349 -1735
rect -349 -1801 349 -1763
rect -349 -1829 -344 -1801
rect -316 -1829 -278 -1801
rect -250 -1829 -212 -1801
rect -184 -1829 -146 -1801
rect -118 -1829 -80 -1801
rect -52 -1829 -14 -1801
rect 14 -1829 52 -1801
rect 80 -1829 118 -1801
rect 146 -1829 184 -1801
rect 212 -1829 250 -1801
rect 278 -1829 316 -1801
rect 344 -1829 349 -1801
rect -349 -1867 349 -1829
rect -349 -1895 -344 -1867
rect -316 -1895 -278 -1867
rect -250 -1895 -212 -1867
rect -184 -1895 -146 -1867
rect -118 -1895 -80 -1867
rect -52 -1895 -14 -1867
rect 14 -1895 52 -1867
rect 80 -1895 118 -1867
rect 146 -1895 184 -1867
rect 212 -1895 250 -1867
rect 278 -1895 316 -1867
rect 344 -1895 349 -1867
rect -349 -1933 349 -1895
rect -349 -1961 -344 -1933
rect -316 -1961 -278 -1933
rect -250 -1961 -212 -1933
rect -184 -1961 -146 -1933
rect -118 -1961 -80 -1933
rect -52 -1961 -14 -1933
rect 14 -1961 52 -1933
rect 80 -1961 118 -1933
rect 146 -1961 184 -1933
rect 212 -1961 250 -1933
rect 278 -1961 316 -1933
rect 344 -1961 349 -1933
rect -349 -1999 349 -1961
rect -349 -2027 -344 -1999
rect -316 -2027 -278 -1999
rect -250 -2027 -212 -1999
rect -184 -2027 -146 -1999
rect -118 -2027 -80 -1999
rect -52 -2027 -14 -1999
rect 14 -2027 52 -1999
rect 80 -2027 118 -1999
rect 146 -2027 184 -1999
rect 212 -2027 250 -1999
rect 278 -2027 316 -1999
rect 344 -2027 349 -1999
rect -349 -2065 349 -2027
rect -349 -2093 -344 -2065
rect -316 -2093 -278 -2065
rect -250 -2093 -212 -2065
rect -184 -2093 -146 -2065
rect -118 -2093 -80 -2065
rect -52 -2093 -14 -2065
rect 14 -2093 52 -2065
rect 80 -2093 118 -2065
rect 146 -2093 184 -2065
rect 212 -2093 250 -2065
rect 278 -2093 316 -2065
rect 344 -2093 349 -2065
rect -349 -2131 349 -2093
rect -349 -2159 -344 -2131
rect -316 -2159 -278 -2131
rect -250 -2159 -212 -2131
rect -184 -2159 -146 -2131
rect -118 -2159 -80 -2131
rect -52 -2159 -14 -2131
rect 14 -2159 52 -2131
rect 80 -2159 118 -2131
rect 146 -2159 184 -2131
rect 212 -2159 250 -2131
rect 278 -2159 316 -2131
rect 344 -2159 349 -2131
rect -349 -2197 349 -2159
rect -349 -2225 -344 -2197
rect -316 -2225 -278 -2197
rect -250 -2225 -212 -2197
rect -184 -2225 -146 -2197
rect -118 -2225 -80 -2197
rect -52 -2225 -14 -2197
rect 14 -2225 52 -2197
rect 80 -2225 118 -2197
rect 146 -2225 184 -2197
rect 212 -2225 250 -2197
rect 278 -2225 316 -2197
rect 344 -2225 349 -2197
rect -349 -2230 349 -2225
<< via3 >>
rect -344 2197 -316 2225
rect -278 2197 -250 2225
rect -212 2197 -184 2225
rect -146 2197 -118 2225
rect -80 2197 -52 2225
rect -14 2197 14 2225
rect 52 2197 80 2225
rect 118 2197 146 2225
rect 184 2197 212 2225
rect 250 2197 278 2225
rect 316 2197 344 2225
rect -344 2131 -316 2159
rect -278 2131 -250 2159
rect -212 2131 -184 2159
rect -146 2131 -118 2159
rect -80 2131 -52 2159
rect -14 2131 14 2159
rect 52 2131 80 2159
rect 118 2131 146 2159
rect 184 2131 212 2159
rect 250 2131 278 2159
rect 316 2131 344 2159
rect -344 2065 -316 2093
rect -278 2065 -250 2093
rect -212 2065 -184 2093
rect -146 2065 -118 2093
rect -80 2065 -52 2093
rect -14 2065 14 2093
rect 52 2065 80 2093
rect 118 2065 146 2093
rect 184 2065 212 2093
rect 250 2065 278 2093
rect 316 2065 344 2093
rect -344 1999 -316 2027
rect -278 1999 -250 2027
rect -212 1999 -184 2027
rect -146 1999 -118 2027
rect -80 1999 -52 2027
rect -14 1999 14 2027
rect 52 1999 80 2027
rect 118 1999 146 2027
rect 184 1999 212 2027
rect 250 1999 278 2027
rect 316 1999 344 2027
rect -344 1933 -316 1961
rect -278 1933 -250 1961
rect -212 1933 -184 1961
rect -146 1933 -118 1961
rect -80 1933 -52 1961
rect -14 1933 14 1961
rect 52 1933 80 1961
rect 118 1933 146 1961
rect 184 1933 212 1961
rect 250 1933 278 1961
rect 316 1933 344 1961
rect -344 1867 -316 1895
rect -278 1867 -250 1895
rect -212 1867 -184 1895
rect -146 1867 -118 1895
rect -80 1867 -52 1895
rect -14 1867 14 1895
rect 52 1867 80 1895
rect 118 1867 146 1895
rect 184 1867 212 1895
rect 250 1867 278 1895
rect 316 1867 344 1895
rect -344 1801 -316 1829
rect -278 1801 -250 1829
rect -212 1801 -184 1829
rect -146 1801 -118 1829
rect -80 1801 -52 1829
rect -14 1801 14 1829
rect 52 1801 80 1829
rect 118 1801 146 1829
rect 184 1801 212 1829
rect 250 1801 278 1829
rect 316 1801 344 1829
rect -344 1735 -316 1763
rect -278 1735 -250 1763
rect -212 1735 -184 1763
rect -146 1735 -118 1763
rect -80 1735 -52 1763
rect -14 1735 14 1763
rect 52 1735 80 1763
rect 118 1735 146 1763
rect 184 1735 212 1763
rect 250 1735 278 1763
rect 316 1735 344 1763
rect -344 1669 -316 1697
rect -278 1669 -250 1697
rect -212 1669 -184 1697
rect -146 1669 -118 1697
rect -80 1669 -52 1697
rect -14 1669 14 1697
rect 52 1669 80 1697
rect 118 1669 146 1697
rect 184 1669 212 1697
rect 250 1669 278 1697
rect 316 1669 344 1697
rect -344 1603 -316 1631
rect -278 1603 -250 1631
rect -212 1603 -184 1631
rect -146 1603 -118 1631
rect -80 1603 -52 1631
rect -14 1603 14 1631
rect 52 1603 80 1631
rect 118 1603 146 1631
rect 184 1603 212 1631
rect 250 1603 278 1631
rect 316 1603 344 1631
rect -344 1537 -316 1565
rect -278 1537 -250 1565
rect -212 1537 -184 1565
rect -146 1537 -118 1565
rect -80 1537 -52 1565
rect -14 1537 14 1565
rect 52 1537 80 1565
rect 118 1537 146 1565
rect 184 1537 212 1565
rect 250 1537 278 1565
rect 316 1537 344 1565
rect -344 1471 -316 1499
rect -278 1471 -250 1499
rect -212 1471 -184 1499
rect -146 1471 -118 1499
rect -80 1471 -52 1499
rect -14 1471 14 1499
rect 52 1471 80 1499
rect 118 1471 146 1499
rect 184 1471 212 1499
rect 250 1471 278 1499
rect 316 1471 344 1499
rect -344 1405 -316 1433
rect -278 1405 -250 1433
rect -212 1405 -184 1433
rect -146 1405 -118 1433
rect -80 1405 -52 1433
rect -14 1405 14 1433
rect 52 1405 80 1433
rect 118 1405 146 1433
rect 184 1405 212 1433
rect 250 1405 278 1433
rect 316 1405 344 1433
rect -344 1339 -316 1367
rect -278 1339 -250 1367
rect -212 1339 -184 1367
rect -146 1339 -118 1367
rect -80 1339 -52 1367
rect -14 1339 14 1367
rect 52 1339 80 1367
rect 118 1339 146 1367
rect 184 1339 212 1367
rect 250 1339 278 1367
rect 316 1339 344 1367
rect -344 1273 -316 1301
rect -278 1273 -250 1301
rect -212 1273 -184 1301
rect -146 1273 -118 1301
rect -80 1273 -52 1301
rect -14 1273 14 1301
rect 52 1273 80 1301
rect 118 1273 146 1301
rect 184 1273 212 1301
rect 250 1273 278 1301
rect 316 1273 344 1301
rect -344 1207 -316 1235
rect -278 1207 -250 1235
rect -212 1207 -184 1235
rect -146 1207 -118 1235
rect -80 1207 -52 1235
rect -14 1207 14 1235
rect 52 1207 80 1235
rect 118 1207 146 1235
rect 184 1207 212 1235
rect 250 1207 278 1235
rect 316 1207 344 1235
rect -344 1141 -316 1169
rect -278 1141 -250 1169
rect -212 1141 -184 1169
rect -146 1141 -118 1169
rect -80 1141 -52 1169
rect -14 1141 14 1169
rect 52 1141 80 1169
rect 118 1141 146 1169
rect 184 1141 212 1169
rect 250 1141 278 1169
rect 316 1141 344 1169
rect -344 1075 -316 1103
rect -278 1075 -250 1103
rect -212 1075 -184 1103
rect -146 1075 -118 1103
rect -80 1075 -52 1103
rect -14 1075 14 1103
rect 52 1075 80 1103
rect 118 1075 146 1103
rect 184 1075 212 1103
rect 250 1075 278 1103
rect 316 1075 344 1103
rect -344 1009 -316 1037
rect -278 1009 -250 1037
rect -212 1009 -184 1037
rect -146 1009 -118 1037
rect -80 1009 -52 1037
rect -14 1009 14 1037
rect 52 1009 80 1037
rect 118 1009 146 1037
rect 184 1009 212 1037
rect 250 1009 278 1037
rect 316 1009 344 1037
rect -344 943 -316 971
rect -278 943 -250 971
rect -212 943 -184 971
rect -146 943 -118 971
rect -80 943 -52 971
rect -14 943 14 971
rect 52 943 80 971
rect 118 943 146 971
rect 184 943 212 971
rect 250 943 278 971
rect 316 943 344 971
rect -344 877 -316 905
rect -278 877 -250 905
rect -212 877 -184 905
rect -146 877 -118 905
rect -80 877 -52 905
rect -14 877 14 905
rect 52 877 80 905
rect 118 877 146 905
rect 184 877 212 905
rect 250 877 278 905
rect 316 877 344 905
rect -344 811 -316 839
rect -278 811 -250 839
rect -212 811 -184 839
rect -146 811 -118 839
rect -80 811 -52 839
rect -14 811 14 839
rect 52 811 80 839
rect 118 811 146 839
rect 184 811 212 839
rect 250 811 278 839
rect 316 811 344 839
rect -344 745 -316 773
rect -278 745 -250 773
rect -212 745 -184 773
rect -146 745 -118 773
rect -80 745 -52 773
rect -14 745 14 773
rect 52 745 80 773
rect 118 745 146 773
rect 184 745 212 773
rect 250 745 278 773
rect 316 745 344 773
rect -344 679 -316 707
rect -278 679 -250 707
rect -212 679 -184 707
rect -146 679 -118 707
rect -80 679 -52 707
rect -14 679 14 707
rect 52 679 80 707
rect 118 679 146 707
rect 184 679 212 707
rect 250 679 278 707
rect 316 679 344 707
rect -344 613 -316 641
rect -278 613 -250 641
rect -212 613 -184 641
rect -146 613 -118 641
rect -80 613 -52 641
rect -14 613 14 641
rect 52 613 80 641
rect 118 613 146 641
rect 184 613 212 641
rect 250 613 278 641
rect 316 613 344 641
rect -344 547 -316 575
rect -278 547 -250 575
rect -212 547 -184 575
rect -146 547 -118 575
rect -80 547 -52 575
rect -14 547 14 575
rect 52 547 80 575
rect 118 547 146 575
rect 184 547 212 575
rect 250 547 278 575
rect 316 547 344 575
rect -344 481 -316 509
rect -278 481 -250 509
rect -212 481 -184 509
rect -146 481 -118 509
rect -80 481 -52 509
rect -14 481 14 509
rect 52 481 80 509
rect 118 481 146 509
rect 184 481 212 509
rect 250 481 278 509
rect 316 481 344 509
rect -344 415 -316 443
rect -278 415 -250 443
rect -212 415 -184 443
rect -146 415 -118 443
rect -80 415 -52 443
rect -14 415 14 443
rect 52 415 80 443
rect 118 415 146 443
rect 184 415 212 443
rect 250 415 278 443
rect 316 415 344 443
rect -344 349 -316 377
rect -278 349 -250 377
rect -212 349 -184 377
rect -146 349 -118 377
rect -80 349 -52 377
rect -14 349 14 377
rect 52 349 80 377
rect 118 349 146 377
rect 184 349 212 377
rect 250 349 278 377
rect 316 349 344 377
rect -344 283 -316 311
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect 316 283 344 311
rect -344 217 -316 245
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect 316 217 344 245
rect -344 151 -316 179
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect 316 151 344 179
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect -344 -179 -316 -151
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect 316 -179 344 -151
rect -344 -245 -316 -217
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect 316 -245 344 -217
rect -344 -311 -316 -283
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
rect 316 -311 344 -283
rect -344 -377 -316 -349
rect -278 -377 -250 -349
rect -212 -377 -184 -349
rect -146 -377 -118 -349
rect -80 -377 -52 -349
rect -14 -377 14 -349
rect 52 -377 80 -349
rect 118 -377 146 -349
rect 184 -377 212 -349
rect 250 -377 278 -349
rect 316 -377 344 -349
rect -344 -443 -316 -415
rect -278 -443 -250 -415
rect -212 -443 -184 -415
rect -146 -443 -118 -415
rect -80 -443 -52 -415
rect -14 -443 14 -415
rect 52 -443 80 -415
rect 118 -443 146 -415
rect 184 -443 212 -415
rect 250 -443 278 -415
rect 316 -443 344 -415
rect -344 -509 -316 -481
rect -278 -509 -250 -481
rect -212 -509 -184 -481
rect -146 -509 -118 -481
rect -80 -509 -52 -481
rect -14 -509 14 -481
rect 52 -509 80 -481
rect 118 -509 146 -481
rect 184 -509 212 -481
rect 250 -509 278 -481
rect 316 -509 344 -481
rect -344 -575 -316 -547
rect -278 -575 -250 -547
rect -212 -575 -184 -547
rect -146 -575 -118 -547
rect -80 -575 -52 -547
rect -14 -575 14 -547
rect 52 -575 80 -547
rect 118 -575 146 -547
rect 184 -575 212 -547
rect 250 -575 278 -547
rect 316 -575 344 -547
rect -344 -641 -316 -613
rect -278 -641 -250 -613
rect -212 -641 -184 -613
rect -146 -641 -118 -613
rect -80 -641 -52 -613
rect -14 -641 14 -613
rect 52 -641 80 -613
rect 118 -641 146 -613
rect 184 -641 212 -613
rect 250 -641 278 -613
rect 316 -641 344 -613
rect -344 -707 -316 -679
rect -278 -707 -250 -679
rect -212 -707 -184 -679
rect -146 -707 -118 -679
rect -80 -707 -52 -679
rect -14 -707 14 -679
rect 52 -707 80 -679
rect 118 -707 146 -679
rect 184 -707 212 -679
rect 250 -707 278 -679
rect 316 -707 344 -679
rect -344 -773 -316 -745
rect -278 -773 -250 -745
rect -212 -773 -184 -745
rect -146 -773 -118 -745
rect -80 -773 -52 -745
rect -14 -773 14 -745
rect 52 -773 80 -745
rect 118 -773 146 -745
rect 184 -773 212 -745
rect 250 -773 278 -745
rect 316 -773 344 -745
rect -344 -839 -316 -811
rect -278 -839 -250 -811
rect -212 -839 -184 -811
rect -146 -839 -118 -811
rect -80 -839 -52 -811
rect -14 -839 14 -811
rect 52 -839 80 -811
rect 118 -839 146 -811
rect 184 -839 212 -811
rect 250 -839 278 -811
rect 316 -839 344 -811
rect -344 -905 -316 -877
rect -278 -905 -250 -877
rect -212 -905 -184 -877
rect -146 -905 -118 -877
rect -80 -905 -52 -877
rect -14 -905 14 -877
rect 52 -905 80 -877
rect 118 -905 146 -877
rect 184 -905 212 -877
rect 250 -905 278 -877
rect 316 -905 344 -877
rect -344 -971 -316 -943
rect -278 -971 -250 -943
rect -212 -971 -184 -943
rect -146 -971 -118 -943
rect -80 -971 -52 -943
rect -14 -971 14 -943
rect 52 -971 80 -943
rect 118 -971 146 -943
rect 184 -971 212 -943
rect 250 -971 278 -943
rect 316 -971 344 -943
rect -344 -1037 -316 -1009
rect -278 -1037 -250 -1009
rect -212 -1037 -184 -1009
rect -146 -1037 -118 -1009
rect -80 -1037 -52 -1009
rect -14 -1037 14 -1009
rect 52 -1037 80 -1009
rect 118 -1037 146 -1009
rect 184 -1037 212 -1009
rect 250 -1037 278 -1009
rect 316 -1037 344 -1009
rect -344 -1103 -316 -1075
rect -278 -1103 -250 -1075
rect -212 -1103 -184 -1075
rect -146 -1103 -118 -1075
rect -80 -1103 -52 -1075
rect -14 -1103 14 -1075
rect 52 -1103 80 -1075
rect 118 -1103 146 -1075
rect 184 -1103 212 -1075
rect 250 -1103 278 -1075
rect 316 -1103 344 -1075
rect -344 -1169 -316 -1141
rect -278 -1169 -250 -1141
rect -212 -1169 -184 -1141
rect -146 -1169 -118 -1141
rect -80 -1169 -52 -1141
rect -14 -1169 14 -1141
rect 52 -1169 80 -1141
rect 118 -1169 146 -1141
rect 184 -1169 212 -1141
rect 250 -1169 278 -1141
rect 316 -1169 344 -1141
rect -344 -1235 -316 -1207
rect -278 -1235 -250 -1207
rect -212 -1235 -184 -1207
rect -146 -1235 -118 -1207
rect -80 -1235 -52 -1207
rect -14 -1235 14 -1207
rect 52 -1235 80 -1207
rect 118 -1235 146 -1207
rect 184 -1235 212 -1207
rect 250 -1235 278 -1207
rect 316 -1235 344 -1207
rect -344 -1301 -316 -1273
rect -278 -1301 -250 -1273
rect -212 -1301 -184 -1273
rect -146 -1301 -118 -1273
rect -80 -1301 -52 -1273
rect -14 -1301 14 -1273
rect 52 -1301 80 -1273
rect 118 -1301 146 -1273
rect 184 -1301 212 -1273
rect 250 -1301 278 -1273
rect 316 -1301 344 -1273
rect -344 -1367 -316 -1339
rect -278 -1367 -250 -1339
rect -212 -1367 -184 -1339
rect -146 -1367 -118 -1339
rect -80 -1367 -52 -1339
rect -14 -1367 14 -1339
rect 52 -1367 80 -1339
rect 118 -1367 146 -1339
rect 184 -1367 212 -1339
rect 250 -1367 278 -1339
rect 316 -1367 344 -1339
rect -344 -1433 -316 -1405
rect -278 -1433 -250 -1405
rect -212 -1433 -184 -1405
rect -146 -1433 -118 -1405
rect -80 -1433 -52 -1405
rect -14 -1433 14 -1405
rect 52 -1433 80 -1405
rect 118 -1433 146 -1405
rect 184 -1433 212 -1405
rect 250 -1433 278 -1405
rect 316 -1433 344 -1405
rect -344 -1499 -316 -1471
rect -278 -1499 -250 -1471
rect -212 -1499 -184 -1471
rect -146 -1499 -118 -1471
rect -80 -1499 -52 -1471
rect -14 -1499 14 -1471
rect 52 -1499 80 -1471
rect 118 -1499 146 -1471
rect 184 -1499 212 -1471
rect 250 -1499 278 -1471
rect 316 -1499 344 -1471
rect -344 -1565 -316 -1537
rect -278 -1565 -250 -1537
rect -212 -1565 -184 -1537
rect -146 -1565 -118 -1537
rect -80 -1565 -52 -1537
rect -14 -1565 14 -1537
rect 52 -1565 80 -1537
rect 118 -1565 146 -1537
rect 184 -1565 212 -1537
rect 250 -1565 278 -1537
rect 316 -1565 344 -1537
rect -344 -1631 -316 -1603
rect -278 -1631 -250 -1603
rect -212 -1631 -184 -1603
rect -146 -1631 -118 -1603
rect -80 -1631 -52 -1603
rect -14 -1631 14 -1603
rect 52 -1631 80 -1603
rect 118 -1631 146 -1603
rect 184 -1631 212 -1603
rect 250 -1631 278 -1603
rect 316 -1631 344 -1603
rect -344 -1697 -316 -1669
rect -278 -1697 -250 -1669
rect -212 -1697 -184 -1669
rect -146 -1697 -118 -1669
rect -80 -1697 -52 -1669
rect -14 -1697 14 -1669
rect 52 -1697 80 -1669
rect 118 -1697 146 -1669
rect 184 -1697 212 -1669
rect 250 -1697 278 -1669
rect 316 -1697 344 -1669
rect -344 -1763 -316 -1735
rect -278 -1763 -250 -1735
rect -212 -1763 -184 -1735
rect -146 -1763 -118 -1735
rect -80 -1763 -52 -1735
rect -14 -1763 14 -1735
rect 52 -1763 80 -1735
rect 118 -1763 146 -1735
rect 184 -1763 212 -1735
rect 250 -1763 278 -1735
rect 316 -1763 344 -1735
rect -344 -1829 -316 -1801
rect -278 -1829 -250 -1801
rect -212 -1829 -184 -1801
rect -146 -1829 -118 -1801
rect -80 -1829 -52 -1801
rect -14 -1829 14 -1801
rect 52 -1829 80 -1801
rect 118 -1829 146 -1801
rect 184 -1829 212 -1801
rect 250 -1829 278 -1801
rect 316 -1829 344 -1801
rect -344 -1895 -316 -1867
rect -278 -1895 -250 -1867
rect -212 -1895 -184 -1867
rect -146 -1895 -118 -1867
rect -80 -1895 -52 -1867
rect -14 -1895 14 -1867
rect 52 -1895 80 -1867
rect 118 -1895 146 -1867
rect 184 -1895 212 -1867
rect 250 -1895 278 -1867
rect 316 -1895 344 -1867
rect -344 -1961 -316 -1933
rect -278 -1961 -250 -1933
rect -212 -1961 -184 -1933
rect -146 -1961 -118 -1933
rect -80 -1961 -52 -1933
rect -14 -1961 14 -1933
rect 52 -1961 80 -1933
rect 118 -1961 146 -1933
rect 184 -1961 212 -1933
rect 250 -1961 278 -1933
rect 316 -1961 344 -1933
rect -344 -2027 -316 -1999
rect -278 -2027 -250 -1999
rect -212 -2027 -184 -1999
rect -146 -2027 -118 -1999
rect -80 -2027 -52 -1999
rect -14 -2027 14 -1999
rect 52 -2027 80 -1999
rect 118 -2027 146 -1999
rect 184 -2027 212 -1999
rect 250 -2027 278 -1999
rect 316 -2027 344 -1999
rect -344 -2093 -316 -2065
rect -278 -2093 -250 -2065
rect -212 -2093 -184 -2065
rect -146 -2093 -118 -2065
rect -80 -2093 -52 -2065
rect -14 -2093 14 -2065
rect 52 -2093 80 -2065
rect 118 -2093 146 -2065
rect 184 -2093 212 -2065
rect 250 -2093 278 -2065
rect 316 -2093 344 -2065
rect -344 -2159 -316 -2131
rect -278 -2159 -250 -2131
rect -212 -2159 -184 -2131
rect -146 -2159 -118 -2131
rect -80 -2159 -52 -2131
rect -14 -2159 14 -2131
rect 52 -2159 80 -2131
rect 118 -2159 146 -2131
rect 184 -2159 212 -2131
rect 250 -2159 278 -2131
rect 316 -2159 344 -2131
rect -344 -2225 -316 -2197
rect -278 -2225 -250 -2197
rect -212 -2225 -184 -2197
rect -146 -2225 -118 -2197
rect -80 -2225 -52 -2197
rect -14 -2225 14 -2197
rect 52 -2225 80 -2197
rect 118 -2225 146 -2197
rect 184 -2225 212 -2197
rect 250 -2225 278 -2197
rect 316 -2225 344 -2197
<< metal4 >>
rect -349 2225 349 2230
rect -349 2197 -344 2225
rect -316 2197 -278 2225
rect -250 2197 -212 2225
rect -184 2197 -146 2225
rect -118 2197 -80 2225
rect -52 2197 -14 2225
rect 14 2197 52 2225
rect 80 2197 118 2225
rect 146 2197 184 2225
rect 212 2197 250 2225
rect 278 2197 316 2225
rect 344 2197 349 2225
rect -349 2159 349 2197
rect -349 2131 -344 2159
rect -316 2131 -278 2159
rect -250 2131 -212 2159
rect -184 2131 -146 2159
rect -118 2131 -80 2159
rect -52 2131 -14 2159
rect 14 2131 52 2159
rect 80 2131 118 2159
rect 146 2131 184 2159
rect 212 2131 250 2159
rect 278 2131 316 2159
rect 344 2131 349 2159
rect -349 2093 349 2131
rect -349 2065 -344 2093
rect -316 2065 -278 2093
rect -250 2065 -212 2093
rect -184 2065 -146 2093
rect -118 2065 -80 2093
rect -52 2065 -14 2093
rect 14 2065 52 2093
rect 80 2065 118 2093
rect 146 2065 184 2093
rect 212 2065 250 2093
rect 278 2065 316 2093
rect 344 2065 349 2093
rect -349 2027 349 2065
rect -349 1999 -344 2027
rect -316 1999 -278 2027
rect -250 1999 -212 2027
rect -184 1999 -146 2027
rect -118 1999 -80 2027
rect -52 1999 -14 2027
rect 14 1999 52 2027
rect 80 1999 118 2027
rect 146 1999 184 2027
rect 212 1999 250 2027
rect 278 1999 316 2027
rect 344 1999 349 2027
rect -349 1961 349 1999
rect -349 1933 -344 1961
rect -316 1933 -278 1961
rect -250 1933 -212 1961
rect -184 1933 -146 1961
rect -118 1933 -80 1961
rect -52 1933 -14 1961
rect 14 1933 52 1961
rect 80 1933 118 1961
rect 146 1933 184 1961
rect 212 1933 250 1961
rect 278 1933 316 1961
rect 344 1933 349 1961
rect -349 1895 349 1933
rect -349 1867 -344 1895
rect -316 1867 -278 1895
rect -250 1867 -212 1895
rect -184 1867 -146 1895
rect -118 1867 -80 1895
rect -52 1867 -14 1895
rect 14 1867 52 1895
rect 80 1867 118 1895
rect 146 1867 184 1895
rect 212 1867 250 1895
rect 278 1867 316 1895
rect 344 1867 349 1895
rect -349 1829 349 1867
rect -349 1801 -344 1829
rect -316 1801 -278 1829
rect -250 1801 -212 1829
rect -184 1801 -146 1829
rect -118 1801 -80 1829
rect -52 1801 -14 1829
rect 14 1801 52 1829
rect 80 1801 118 1829
rect 146 1801 184 1829
rect 212 1801 250 1829
rect 278 1801 316 1829
rect 344 1801 349 1829
rect -349 1763 349 1801
rect -349 1735 -344 1763
rect -316 1735 -278 1763
rect -250 1735 -212 1763
rect -184 1735 -146 1763
rect -118 1735 -80 1763
rect -52 1735 -14 1763
rect 14 1735 52 1763
rect 80 1735 118 1763
rect 146 1735 184 1763
rect 212 1735 250 1763
rect 278 1735 316 1763
rect 344 1735 349 1763
rect -349 1697 349 1735
rect -349 1669 -344 1697
rect -316 1669 -278 1697
rect -250 1669 -212 1697
rect -184 1669 -146 1697
rect -118 1669 -80 1697
rect -52 1669 -14 1697
rect 14 1669 52 1697
rect 80 1669 118 1697
rect 146 1669 184 1697
rect 212 1669 250 1697
rect 278 1669 316 1697
rect 344 1669 349 1697
rect -349 1631 349 1669
rect -349 1603 -344 1631
rect -316 1603 -278 1631
rect -250 1603 -212 1631
rect -184 1603 -146 1631
rect -118 1603 -80 1631
rect -52 1603 -14 1631
rect 14 1603 52 1631
rect 80 1603 118 1631
rect 146 1603 184 1631
rect 212 1603 250 1631
rect 278 1603 316 1631
rect 344 1603 349 1631
rect -349 1565 349 1603
rect -349 1537 -344 1565
rect -316 1537 -278 1565
rect -250 1537 -212 1565
rect -184 1537 -146 1565
rect -118 1537 -80 1565
rect -52 1537 -14 1565
rect 14 1537 52 1565
rect 80 1537 118 1565
rect 146 1537 184 1565
rect 212 1537 250 1565
rect 278 1537 316 1565
rect 344 1537 349 1565
rect -349 1499 349 1537
rect -349 1471 -344 1499
rect -316 1471 -278 1499
rect -250 1471 -212 1499
rect -184 1471 -146 1499
rect -118 1471 -80 1499
rect -52 1471 -14 1499
rect 14 1471 52 1499
rect 80 1471 118 1499
rect 146 1471 184 1499
rect 212 1471 250 1499
rect 278 1471 316 1499
rect 344 1471 349 1499
rect -349 1433 349 1471
rect -349 1405 -344 1433
rect -316 1405 -278 1433
rect -250 1405 -212 1433
rect -184 1405 -146 1433
rect -118 1405 -80 1433
rect -52 1405 -14 1433
rect 14 1405 52 1433
rect 80 1405 118 1433
rect 146 1405 184 1433
rect 212 1405 250 1433
rect 278 1405 316 1433
rect 344 1405 349 1433
rect -349 1367 349 1405
rect -349 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 349 1367
rect -349 1301 349 1339
rect -349 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 349 1301
rect -349 1235 349 1273
rect -349 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 349 1235
rect -349 1169 349 1207
rect -349 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 349 1169
rect -349 1103 349 1141
rect -349 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 349 1103
rect -349 1037 349 1075
rect -349 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 349 1037
rect -349 971 349 1009
rect -349 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 349 971
rect -349 905 349 943
rect -349 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 349 905
rect -349 839 349 877
rect -349 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 349 839
rect -349 773 349 811
rect -349 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 349 773
rect -349 707 349 745
rect -349 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 349 707
rect -349 641 349 679
rect -349 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 349 641
rect -349 575 349 613
rect -349 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 349 575
rect -349 509 349 547
rect -349 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 349 509
rect -349 443 349 481
rect -349 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 349 443
rect -349 377 349 415
rect -349 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 349 377
rect -349 311 349 349
rect -349 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 349 311
rect -349 245 349 283
rect -349 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 349 245
rect -349 179 349 217
rect -349 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 349 179
rect -349 113 349 151
rect -349 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 349 113
rect -349 47 349 85
rect -349 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 349 47
rect -349 -19 349 19
rect -349 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 349 -19
rect -349 -85 349 -47
rect -349 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 349 -85
rect -349 -151 349 -113
rect -349 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 349 -151
rect -349 -217 349 -179
rect -349 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 349 -217
rect -349 -283 349 -245
rect -349 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 349 -283
rect -349 -349 349 -311
rect -349 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 349 -349
rect -349 -415 349 -377
rect -349 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 349 -415
rect -349 -481 349 -443
rect -349 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 349 -481
rect -349 -547 349 -509
rect -349 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 349 -547
rect -349 -613 349 -575
rect -349 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 349 -613
rect -349 -679 349 -641
rect -349 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 349 -679
rect -349 -745 349 -707
rect -349 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 349 -745
rect -349 -811 349 -773
rect -349 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 349 -811
rect -349 -877 349 -839
rect -349 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 349 -877
rect -349 -943 349 -905
rect -349 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 349 -943
rect -349 -1009 349 -971
rect -349 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 349 -1009
rect -349 -1075 349 -1037
rect -349 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 349 -1075
rect -349 -1141 349 -1103
rect -349 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 349 -1141
rect -349 -1207 349 -1169
rect -349 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 349 -1207
rect -349 -1273 349 -1235
rect -349 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 349 -1273
rect -349 -1339 349 -1301
rect -349 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 349 -1339
rect -349 -1405 349 -1367
rect -349 -1433 -344 -1405
rect -316 -1433 -278 -1405
rect -250 -1433 -212 -1405
rect -184 -1433 -146 -1405
rect -118 -1433 -80 -1405
rect -52 -1433 -14 -1405
rect 14 -1433 52 -1405
rect 80 -1433 118 -1405
rect 146 -1433 184 -1405
rect 212 -1433 250 -1405
rect 278 -1433 316 -1405
rect 344 -1433 349 -1405
rect -349 -1471 349 -1433
rect -349 -1499 -344 -1471
rect -316 -1499 -278 -1471
rect -250 -1499 -212 -1471
rect -184 -1499 -146 -1471
rect -118 -1499 -80 -1471
rect -52 -1499 -14 -1471
rect 14 -1499 52 -1471
rect 80 -1499 118 -1471
rect 146 -1499 184 -1471
rect 212 -1499 250 -1471
rect 278 -1499 316 -1471
rect 344 -1499 349 -1471
rect -349 -1537 349 -1499
rect -349 -1565 -344 -1537
rect -316 -1565 -278 -1537
rect -250 -1565 -212 -1537
rect -184 -1565 -146 -1537
rect -118 -1565 -80 -1537
rect -52 -1565 -14 -1537
rect 14 -1565 52 -1537
rect 80 -1565 118 -1537
rect 146 -1565 184 -1537
rect 212 -1565 250 -1537
rect 278 -1565 316 -1537
rect 344 -1565 349 -1537
rect -349 -1603 349 -1565
rect -349 -1631 -344 -1603
rect -316 -1631 -278 -1603
rect -250 -1631 -212 -1603
rect -184 -1631 -146 -1603
rect -118 -1631 -80 -1603
rect -52 -1631 -14 -1603
rect 14 -1631 52 -1603
rect 80 -1631 118 -1603
rect 146 -1631 184 -1603
rect 212 -1631 250 -1603
rect 278 -1631 316 -1603
rect 344 -1631 349 -1603
rect -349 -1669 349 -1631
rect -349 -1697 -344 -1669
rect -316 -1697 -278 -1669
rect -250 -1697 -212 -1669
rect -184 -1697 -146 -1669
rect -118 -1697 -80 -1669
rect -52 -1697 -14 -1669
rect 14 -1697 52 -1669
rect 80 -1697 118 -1669
rect 146 -1697 184 -1669
rect 212 -1697 250 -1669
rect 278 -1697 316 -1669
rect 344 -1697 349 -1669
rect -349 -1735 349 -1697
rect -349 -1763 -344 -1735
rect -316 -1763 -278 -1735
rect -250 -1763 -212 -1735
rect -184 -1763 -146 -1735
rect -118 -1763 -80 -1735
rect -52 -1763 -14 -1735
rect 14 -1763 52 -1735
rect 80 -1763 118 -1735
rect 146 -1763 184 -1735
rect 212 -1763 250 -1735
rect 278 -1763 316 -1735
rect 344 -1763 349 -1735
rect -349 -1801 349 -1763
rect -349 -1829 -344 -1801
rect -316 -1829 -278 -1801
rect -250 -1829 -212 -1801
rect -184 -1829 -146 -1801
rect -118 -1829 -80 -1801
rect -52 -1829 -14 -1801
rect 14 -1829 52 -1801
rect 80 -1829 118 -1801
rect 146 -1829 184 -1801
rect 212 -1829 250 -1801
rect 278 -1829 316 -1801
rect 344 -1829 349 -1801
rect -349 -1867 349 -1829
rect -349 -1895 -344 -1867
rect -316 -1895 -278 -1867
rect -250 -1895 -212 -1867
rect -184 -1895 -146 -1867
rect -118 -1895 -80 -1867
rect -52 -1895 -14 -1867
rect 14 -1895 52 -1867
rect 80 -1895 118 -1867
rect 146 -1895 184 -1867
rect 212 -1895 250 -1867
rect 278 -1895 316 -1867
rect 344 -1895 349 -1867
rect -349 -1933 349 -1895
rect -349 -1961 -344 -1933
rect -316 -1961 -278 -1933
rect -250 -1961 -212 -1933
rect -184 -1961 -146 -1933
rect -118 -1961 -80 -1933
rect -52 -1961 -14 -1933
rect 14 -1961 52 -1933
rect 80 -1961 118 -1933
rect 146 -1961 184 -1933
rect 212 -1961 250 -1933
rect 278 -1961 316 -1933
rect 344 -1961 349 -1933
rect -349 -1999 349 -1961
rect -349 -2027 -344 -1999
rect -316 -2027 -278 -1999
rect -250 -2027 -212 -1999
rect -184 -2027 -146 -1999
rect -118 -2027 -80 -1999
rect -52 -2027 -14 -1999
rect 14 -2027 52 -1999
rect 80 -2027 118 -1999
rect 146 -2027 184 -1999
rect 212 -2027 250 -1999
rect 278 -2027 316 -1999
rect 344 -2027 349 -1999
rect -349 -2065 349 -2027
rect -349 -2093 -344 -2065
rect -316 -2093 -278 -2065
rect -250 -2093 -212 -2065
rect -184 -2093 -146 -2065
rect -118 -2093 -80 -2065
rect -52 -2093 -14 -2065
rect 14 -2093 52 -2065
rect 80 -2093 118 -2065
rect 146 -2093 184 -2065
rect 212 -2093 250 -2065
rect 278 -2093 316 -2065
rect 344 -2093 349 -2065
rect -349 -2131 349 -2093
rect -349 -2159 -344 -2131
rect -316 -2159 -278 -2131
rect -250 -2159 -212 -2131
rect -184 -2159 -146 -2131
rect -118 -2159 -80 -2131
rect -52 -2159 -14 -2131
rect 14 -2159 52 -2131
rect 80 -2159 118 -2131
rect 146 -2159 184 -2131
rect 212 -2159 250 -2131
rect 278 -2159 316 -2131
rect 344 -2159 349 -2131
rect -349 -2197 349 -2159
rect -349 -2225 -344 -2197
rect -316 -2225 -278 -2197
rect -250 -2225 -212 -2197
rect -184 -2225 -146 -2197
rect -118 -2225 -80 -2197
rect -52 -2225 -14 -2197
rect 14 -2225 52 -2197
rect 80 -2225 118 -2197
rect 146 -2225 184 -2197
rect 212 -2225 250 -2197
rect 278 -2225 316 -2197
rect 344 -2225 349 -2197
rect -349 -2230 349 -2225
<< end >>
