magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -3992 -2209 6486 9070
<< nwell >>
rect -1809 6365 86 7070
rect -1809 6364 360 6365
rect -1809 6065 3868 6364
rect -1809 5929 3861 6065
rect -1809 5685 740 5929
rect -1809 5664 360 5685
rect -62 4310 4299 4347
rect -62 4136 298 4310
rect 4262 4136 4299 4310
rect -62 3627 4299 4136
rect -62 3565 1081 3627
rect 1086 3565 4299 3627
rect -62 3490 661 3565
rect 4261 3490 4299 3565
rect -62 2767 4299 3490
rect 159 2695 619 2767
rect 4262 2695 4299 2767
rect -62 2403 4299 2695
<< pwell >>
rect 676 5063 757 5067
rect 773 5063 776 5067
rect 1956 5040 2387 5296
rect 1975 4687 2387 4943
<< psubdiff >>
rect -1778 5513 -1650 5562
rect -1778 5467 -1737 5513
rect -1691 5467 -1650 5513
rect -1778 5416 -1650 5467
rect -1511 5513 -1383 5562
rect -1511 5467 -1470 5513
rect -1424 5467 -1383 5513
rect -1511 5416 -1383 5467
rect -1301 5513 -1173 5562
rect -1301 5467 -1260 5513
rect -1214 5467 -1173 5513
rect -1301 5416 -1173 5467
rect -1091 5513 -963 5562
rect -1091 5467 -1050 5513
rect -1004 5467 -963 5513
rect -1091 5416 -963 5467
rect -881 5513 -753 5562
rect -881 5467 -840 5513
rect -794 5467 -753 5513
rect -881 5416 -753 5467
rect -671 5513 -543 5562
rect -671 5467 -630 5513
rect -584 5467 -543 5513
rect -671 5416 -543 5467
rect -461 5513 -333 5562
rect -461 5467 -420 5513
rect -374 5467 -333 5513
rect -461 5416 -333 5467
rect -251 5513 -123 5562
rect -251 5467 -210 5513
rect -164 5467 -123 5513
rect -251 5416 -123 5467
rect 360 5516 488 5565
rect 360 5470 401 5516
rect 447 5470 488 5516
rect 360 5419 488 5470
rect 570 5516 698 5565
rect 570 5470 611 5516
rect 657 5470 698 5516
rect 570 5419 698 5470
rect 780 5516 908 5565
rect 780 5470 821 5516
rect 867 5470 908 5516
rect 780 5419 908 5470
rect 990 5516 1118 5565
rect 990 5470 1031 5516
rect 1077 5470 1118 5516
rect 990 5419 1118 5470
rect 1200 5516 1328 5565
rect 1200 5470 1241 5516
rect 1287 5470 1328 5516
rect 1200 5419 1328 5470
rect 1410 5516 1538 5565
rect 1410 5470 1451 5516
rect 1497 5470 1538 5516
rect 1410 5419 1538 5470
rect 1620 5516 1748 5565
rect 1620 5470 1661 5516
rect 1707 5470 1748 5516
rect 1620 5419 1748 5470
rect 1830 5516 1958 5565
rect 1830 5470 1871 5516
rect 1917 5470 1958 5516
rect 1830 5419 1958 5470
rect 2040 5516 2168 5565
rect 2040 5470 2081 5516
rect 2127 5470 2168 5516
rect 2040 5419 2168 5470
rect 2250 5516 2378 5565
rect 2250 5470 2291 5516
rect 2337 5470 2378 5516
rect 2250 5419 2378 5470
rect 2460 5516 2588 5565
rect 2460 5470 2501 5516
rect 2547 5470 2588 5516
rect 2460 5419 2588 5470
rect 2670 5516 2798 5565
rect 2670 5470 2711 5516
rect 2757 5470 2798 5516
rect 2670 5419 2798 5470
rect 2880 5516 3008 5565
rect 2880 5470 2921 5516
rect 2967 5470 3008 5516
rect 2880 5419 3008 5470
rect 3090 5516 3218 5565
rect 3090 5470 3131 5516
rect 3177 5470 3218 5516
rect 3090 5419 3218 5470
rect 3300 5516 3428 5565
rect 3300 5470 3341 5516
rect 3387 5470 3428 5516
rect 3300 5419 3428 5470
rect 3510 5516 3638 5565
rect 3510 5470 3551 5516
rect 3597 5470 3638 5516
rect 3510 5419 3638 5470
rect 3720 5516 3848 5565
rect 3720 5470 3761 5516
rect 3807 5470 3848 5516
rect 3720 5419 3848 5470
rect -1637 4512 -1509 4561
rect -1637 4466 -1596 4512
rect -1550 4466 -1509 4512
rect -1637 4415 -1509 4466
rect -1427 4512 -1299 4561
rect -1427 4466 -1386 4512
rect -1340 4466 -1299 4512
rect -1427 4415 -1299 4466
rect -1217 4512 -1089 4561
rect -1217 4466 -1176 4512
rect -1130 4466 -1089 4512
rect -1217 4415 -1089 4466
rect -1007 4512 -879 4561
rect -1007 4466 -966 4512
rect -920 4466 -879 4512
rect -1007 4415 -879 4466
rect -797 4512 -669 4561
rect -797 4466 -756 4512
rect -710 4466 -669 4512
rect -797 4415 -669 4466
rect -587 4512 -459 4561
rect -587 4466 -546 4512
rect -500 4466 -459 4512
rect -587 4415 -459 4466
rect -377 4512 -249 4561
rect -377 4466 -336 4512
rect -290 4466 -249 4512
rect -377 4415 -249 4466
rect -167 4512 -39 4561
rect -167 4466 -126 4512
rect -80 4466 -39 4512
rect -167 4415 -39 4466
rect 360 4497 488 4546
rect 360 4451 401 4497
rect 447 4451 488 4497
rect 360 4400 488 4451
rect 570 4497 698 4546
rect 570 4451 611 4497
rect 657 4451 698 4497
rect 570 4400 698 4451
rect 780 4497 908 4546
rect 780 4451 821 4497
rect 867 4451 908 4497
rect 780 4400 908 4451
rect 990 4497 1118 4546
rect 990 4451 1031 4497
rect 1077 4451 1118 4497
rect 990 4400 1118 4451
rect 1200 4497 1328 4546
rect 1200 4451 1241 4497
rect 1287 4451 1328 4497
rect 1200 4400 1328 4451
rect 1410 4497 1538 4546
rect 1410 4451 1451 4497
rect 1497 4451 1538 4497
rect 1410 4400 1538 4451
rect 1620 4497 1748 4546
rect 1620 4451 1661 4497
rect 1707 4451 1748 4497
rect 1620 4400 1748 4451
rect 1830 4497 1958 4546
rect 1830 4451 1871 4497
rect 1917 4451 1958 4497
rect 1830 4400 1958 4451
rect 2040 4497 2168 4546
rect 2040 4451 2081 4497
rect 2127 4451 2168 4497
rect 2040 4400 2168 4451
rect 2250 4497 2378 4546
rect 2250 4451 2291 4497
rect 2337 4451 2378 4497
rect 2250 4400 2378 4451
rect 2460 4497 2588 4546
rect 2460 4451 2501 4497
rect 2547 4451 2588 4497
rect 2460 4400 2588 4451
rect 2670 4497 2798 4546
rect 2670 4451 2711 4497
rect 2757 4451 2798 4497
rect 2670 4400 2798 4451
rect 2880 4497 3008 4546
rect 2880 4451 2921 4497
rect 2967 4451 3008 4497
rect 2880 4400 3008 4451
rect 3090 4497 3218 4546
rect 3090 4451 3131 4497
rect 3177 4451 3218 4497
rect 3090 4400 3218 4451
rect 3300 4497 3428 4546
rect 3300 4451 3341 4497
rect 3387 4451 3428 4497
rect 3300 4400 3428 4451
rect 3510 4497 3638 4546
rect 3510 4451 3551 4497
rect 3597 4451 3638 4497
rect 3510 4400 3638 4451
rect 3720 4497 3848 4546
rect 3720 4451 3761 4497
rect 3807 4451 3848 4497
rect 3720 4400 3848 4451
rect 0 2308 128 2357
rect 0 2262 41 2308
rect 87 2262 128 2308
rect 0 2211 128 2262
rect 210 2308 338 2357
rect 210 2262 251 2308
rect 297 2262 338 2308
rect 210 2211 338 2262
rect 420 2308 548 2357
rect 420 2262 461 2308
rect 507 2262 548 2308
rect 420 2211 548 2262
rect 630 2308 758 2357
rect 630 2262 671 2308
rect 717 2262 758 2308
rect 630 2211 758 2262
rect 840 2308 968 2357
rect 840 2262 881 2308
rect 927 2262 968 2308
rect 840 2211 968 2262
rect 1050 2308 1178 2357
rect 1050 2262 1091 2308
rect 1137 2262 1178 2308
rect 1050 2211 1178 2262
rect 1260 2308 1388 2357
rect 1260 2262 1301 2308
rect 1347 2262 1388 2308
rect 1260 2211 1388 2262
rect 1470 2308 1598 2357
rect 1470 2262 1511 2308
rect 1557 2262 1598 2308
rect 1470 2211 1598 2262
rect 1680 2308 1808 2357
rect 1680 2262 1721 2308
rect 1767 2262 1808 2308
rect 1680 2211 1808 2262
rect 1890 2308 2018 2357
rect 1890 2262 1931 2308
rect 1977 2262 2018 2308
rect 1890 2211 2018 2262
rect 2100 2308 2228 2357
rect 2100 2262 2141 2308
rect 2187 2262 2228 2308
rect 2100 2211 2228 2262
rect 2310 2308 2438 2357
rect 2310 2262 2351 2308
rect 2397 2262 2438 2308
rect 2310 2211 2438 2262
rect 2520 2308 2648 2357
rect 2520 2262 2561 2308
rect 2607 2262 2648 2308
rect 2520 2211 2648 2262
rect 2730 2308 2858 2357
rect 2730 2262 2771 2308
rect 2817 2262 2858 2308
rect 2730 2211 2858 2262
rect 2940 2308 3068 2357
rect 2940 2262 2981 2308
rect 3027 2262 3068 2308
rect 2940 2211 3068 2262
rect 3150 2308 3278 2357
rect 3150 2262 3191 2308
rect 3237 2262 3278 2308
rect 3150 2211 3278 2262
rect 3360 2308 3488 2357
rect 3360 2262 3401 2308
rect 3447 2262 3488 2308
rect 3360 2211 3488 2262
rect 3570 2308 3698 2357
rect 3570 2262 3611 2308
rect 3657 2262 3698 2308
rect 3570 2211 3698 2262
rect 3780 2308 3908 2357
rect 3780 2262 3821 2308
rect 3867 2262 3908 2308
rect 3780 2211 3908 2262
rect 3990 2308 4118 2357
rect 3990 2262 4031 2308
rect 4077 2262 4118 2308
rect 3990 2211 4118 2262
rect 0 1093 128 1142
rect 0 1047 41 1093
rect 87 1047 128 1093
rect 0 996 128 1047
rect 210 1093 338 1142
rect 210 1047 251 1093
rect 297 1047 338 1093
rect 210 996 338 1047
rect 420 1093 548 1142
rect 420 1047 461 1093
rect 507 1047 548 1093
rect 420 996 548 1047
rect 630 1093 758 1142
rect 630 1047 671 1093
rect 717 1047 758 1093
rect 630 996 758 1047
rect 840 1093 968 1142
rect 840 1047 881 1093
rect 927 1047 968 1093
rect 840 996 968 1047
rect 1050 1093 1178 1142
rect 1050 1047 1091 1093
rect 1137 1047 1178 1093
rect 1050 996 1178 1047
rect 1260 1093 1388 1142
rect 1260 1047 1301 1093
rect 1347 1047 1388 1093
rect 1260 996 1388 1047
rect 1470 1093 1598 1142
rect 1470 1047 1511 1093
rect 1557 1047 1598 1093
rect 1470 996 1598 1047
rect 1680 1093 1808 1142
rect 1680 1047 1721 1093
rect 1767 1047 1808 1093
rect 1680 996 1808 1047
rect 1890 1093 2018 1142
rect 1890 1047 1931 1093
rect 1977 1047 2018 1093
rect 1890 996 2018 1047
rect 2100 1093 2228 1142
rect 2100 1047 2141 1093
rect 2187 1047 2228 1093
rect 2100 996 2228 1047
rect 2310 1093 2438 1142
rect 2310 1047 2351 1093
rect 2397 1047 2438 1093
rect 2310 996 2438 1047
rect 2520 1093 2648 1142
rect 2520 1047 2561 1093
rect 2607 1047 2648 1093
rect 2520 996 2648 1047
rect 2730 1093 2858 1142
rect 2730 1047 2771 1093
rect 2817 1047 2858 1093
rect 2730 996 2858 1047
rect 2940 1093 3068 1142
rect 2940 1047 2981 1093
rect 3027 1047 3068 1093
rect 2940 996 3068 1047
rect 3150 1093 3278 1142
rect 3150 1047 3191 1093
rect 3237 1047 3278 1093
rect 3150 996 3278 1047
rect 3360 1093 3488 1142
rect 3360 1047 3401 1093
rect 3447 1047 3488 1093
rect 3360 996 3488 1047
rect 3570 1093 3698 1142
rect 3570 1047 3611 1093
rect 3657 1047 3698 1093
rect 3570 996 3698 1047
rect 3780 1093 3908 1142
rect 3780 1047 3821 1093
rect 3867 1047 3908 1093
rect 3780 996 3908 1047
rect 3990 1093 4118 1142
rect 3990 1047 4031 1093
rect 4077 1047 4118 1093
rect 3990 996 4118 1047
rect 0 -112 128 -63
rect 0 -158 41 -112
rect 87 -158 128 -112
rect 0 -209 128 -158
rect 210 -112 338 -63
rect 210 -158 251 -112
rect 297 -158 338 -112
rect 210 -209 338 -158
rect 420 -112 548 -63
rect 420 -158 461 -112
rect 507 -158 548 -112
rect 420 -209 548 -158
rect 630 -112 758 -63
rect 630 -158 671 -112
rect 717 -158 758 -112
rect 630 -209 758 -158
rect 840 -112 968 -63
rect 840 -158 881 -112
rect 927 -158 968 -112
rect 840 -209 968 -158
rect 1050 -112 1178 -63
rect 1050 -158 1091 -112
rect 1137 -158 1178 -112
rect 1050 -209 1178 -158
rect 1260 -112 1388 -63
rect 1260 -158 1301 -112
rect 1347 -158 1388 -112
rect 1260 -209 1388 -158
rect 1470 -112 1598 -63
rect 1470 -158 1511 -112
rect 1557 -158 1598 -112
rect 1470 -209 1598 -158
rect 1680 -112 1808 -63
rect 1680 -158 1721 -112
rect 1767 -158 1808 -112
rect 1680 -209 1808 -158
rect 1890 -112 2018 -63
rect 1890 -158 1931 -112
rect 1977 -158 2018 -112
rect 1890 -209 2018 -158
rect 2100 -112 2228 -63
rect 2100 -158 2141 -112
rect 2187 -158 2228 -112
rect 2100 -209 2228 -158
rect 2310 -112 2438 -63
rect 2310 -158 2351 -112
rect 2397 -158 2438 -112
rect 2310 -209 2438 -158
rect 2520 -112 2648 -63
rect 2520 -158 2561 -112
rect 2607 -158 2648 -112
rect 2520 -209 2648 -158
rect 2730 -112 2858 -63
rect 2730 -158 2771 -112
rect 2817 -158 2858 -112
rect 2730 -209 2858 -158
rect 2940 -112 3068 -63
rect 2940 -158 2981 -112
rect 3027 -158 3068 -112
rect 2940 -209 3068 -158
rect 3150 -112 3278 -63
rect 3150 -158 3191 -112
rect 3237 -158 3278 -112
rect 3150 -209 3278 -158
rect 3360 -112 3488 -63
rect 3360 -158 3401 -112
rect 3447 -158 3488 -112
rect 3360 -209 3488 -158
rect 3570 -112 3698 -63
rect 3570 -158 3611 -112
rect 3657 -158 3698 -112
rect 3570 -209 3698 -158
rect 3780 -112 3908 -63
rect 3780 -158 3821 -112
rect 3867 -158 3908 -112
rect 3780 -209 3908 -158
rect 3990 -112 4118 -63
rect 3990 -158 4031 -112
rect 4077 -158 4118 -112
rect 3990 -209 4118 -158
<< nsubdiff >>
rect -1758 7032 -1588 7046
rect -1758 6892 -1745 7032
rect -1605 6892 -1588 7032
rect -1758 6878 -1588 6892
rect -1528 7032 -1358 7046
rect -1528 6892 -1515 7032
rect -1375 6892 -1358 7032
rect -1528 6878 -1358 6892
rect -1298 7032 -1128 7046
rect -1298 6892 -1285 7032
rect -1145 6892 -1128 7032
rect -1298 6878 -1128 6892
rect -1068 7032 -898 7046
rect -1068 6892 -1055 7032
rect -915 6892 -898 7032
rect -1068 6878 -898 6892
rect -838 7032 -668 7046
rect -838 6892 -825 7032
rect -685 6892 -668 7032
rect -838 6878 -668 6892
rect -608 7032 -438 7046
rect -608 6892 -595 7032
rect -455 6892 -438 7032
rect -608 6878 -438 6892
rect -378 7032 -208 7046
rect -378 6892 -365 7032
rect -225 6892 -208 7032
rect -378 6878 -208 6892
rect -133 7032 37 7046
rect -133 6892 -120 7032
rect 20 6892 37 7032
rect -133 6878 37 6892
rect 420 6326 590 6340
rect 420 6186 433 6326
rect 573 6186 590 6326
rect 420 6172 590 6186
rect 650 6326 820 6340
rect 650 6186 663 6326
rect 803 6186 820 6326
rect 650 6172 820 6186
rect 880 6326 1050 6340
rect 880 6186 893 6326
rect 1033 6186 1050 6326
rect 880 6172 1050 6186
rect 1110 6326 1280 6340
rect 1110 6186 1123 6326
rect 1263 6186 1280 6326
rect 1110 6172 1280 6186
rect 1340 6326 1510 6340
rect 1340 6186 1353 6326
rect 1493 6186 1510 6326
rect 1340 6172 1510 6186
rect 1570 6326 1740 6340
rect 1570 6186 1583 6326
rect 1723 6186 1740 6326
rect 1570 6172 1740 6186
rect 1800 6326 1970 6340
rect 1800 6186 1813 6326
rect 1953 6186 1970 6326
rect 1800 6172 1970 6186
rect 2030 6326 2200 6340
rect 2030 6186 2043 6326
rect 2183 6186 2200 6326
rect 2030 6172 2200 6186
rect 2260 6326 2430 6340
rect 2260 6186 2273 6326
rect 2413 6186 2430 6326
rect 2260 6172 2430 6186
rect 2490 6326 2660 6340
rect 2490 6186 2503 6326
rect 2643 6186 2660 6326
rect 2490 6172 2660 6186
rect 2720 6326 2890 6340
rect 2720 6186 2733 6326
rect 2873 6186 2890 6326
rect 2720 6172 2890 6186
rect 2950 6326 3120 6340
rect 2950 6186 2963 6326
rect 3103 6186 3120 6326
rect 2950 6172 3120 6186
rect 3180 6326 3350 6340
rect 3180 6186 3193 6326
rect 3333 6186 3350 6326
rect 3180 6172 3350 6186
rect 3410 6326 3580 6340
rect 3410 6186 3423 6326
rect 3563 6186 3580 6326
rect 3410 6172 3580 6186
rect 3640 6326 3810 6340
rect 3640 6186 3653 6326
rect 3793 6186 3810 6326
rect 3640 6172 3810 6186
rect -1758 5842 -1588 5856
rect -1758 5702 -1745 5842
rect -1605 5702 -1588 5842
rect -1758 5688 -1588 5702
rect -1528 5842 -1358 5856
rect -1528 5702 -1515 5842
rect -1375 5702 -1358 5842
rect -1528 5688 -1358 5702
rect -1298 5842 -1128 5856
rect -1298 5702 -1285 5842
rect -1145 5702 -1128 5842
rect -1298 5688 -1128 5702
rect -1068 5842 -898 5856
rect -1068 5702 -1055 5842
rect -915 5702 -898 5842
rect -1068 5688 -898 5702
rect -838 5842 -668 5856
rect -838 5702 -825 5842
rect -685 5702 -668 5842
rect -838 5688 -668 5702
rect -608 5842 -438 5856
rect -608 5702 -595 5842
rect -455 5702 -438 5842
rect -608 5688 -438 5702
rect -378 5842 -208 5856
rect -378 5702 -365 5842
rect -225 5702 -208 5842
rect -378 5688 -208 5702
rect -133 5842 37 5856
rect -133 5702 -120 5842
rect 20 5702 37 5842
rect -133 5688 37 5702
rect -35 3876 135 3890
rect -35 3736 -22 3876
rect 118 3736 135 3876
rect -35 3722 135 3736
rect 195 3876 365 3890
rect 195 3736 208 3876
rect 348 3736 365 3876
rect 195 3722 365 3736
rect 425 3876 595 3890
rect 425 3736 438 3876
rect 578 3736 595 3876
rect 425 3722 595 3736
rect 655 3876 825 3890
rect 655 3736 668 3876
rect 808 3736 825 3876
rect 655 3722 825 3736
rect 885 3876 1055 3890
rect 885 3736 898 3876
rect 1038 3736 1055 3876
rect 885 3722 1055 3736
rect 1115 3876 1285 3890
rect 1115 3736 1128 3876
rect 1268 3736 1285 3876
rect 1115 3722 1285 3736
rect 1345 3876 1515 3890
rect 1345 3736 1358 3876
rect 1498 3736 1515 3876
rect 1345 3722 1515 3736
rect 1575 3876 1745 3890
rect 1575 3736 1588 3876
rect 1728 3736 1745 3876
rect 1575 3722 1745 3736
rect 1805 3876 1975 3890
rect 1805 3736 1818 3876
rect 1958 3736 1975 3876
rect 1805 3722 1975 3736
rect 2035 3876 2205 3890
rect 2035 3736 2048 3876
rect 2188 3736 2205 3876
rect 2035 3722 2205 3736
rect 2265 3876 2435 3890
rect 2265 3736 2278 3876
rect 2418 3736 2435 3876
rect 2265 3722 2435 3736
rect 2495 3876 2665 3890
rect 2495 3736 2508 3876
rect 2648 3736 2665 3876
rect 2495 3722 2665 3736
rect 2725 3876 2895 3890
rect 2725 3736 2738 3876
rect 2878 3736 2895 3876
rect 2725 3722 2895 3736
rect 2955 3876 3125 3890
rect 2955 3736 2968 3876
rect 3108 3736 3125 3876
rect 2955 3722 3125 3736
rect 3185 3876 3355 3890
rect 3185 3736 3198 3876
rect 3338 3736 3355 3876
rect 3185 3722 3355 3736
rect 3415 3876 3585 3890
rect 3415 3736 3428 3876
rect 3568 3736 3585 3876
rect 3415 3722 3585 3736
rect 3645 3876 3815 3890
rect 3645 3736 3658 3876
rect 3798 3736 3815 3876
rect 3645 3722 3815 3736
rect 3875 3876 4045 3890
rect 3875 3736 3888 3876
rect 4028 3736 4045 3876
rect 3875 3722 4045 3736
rect 4105 3876 4275 3890
rect 4105 3736 4118 3876
rect 4258 3736 4275 3876
rect 4105 3722 4275 3736
rect -35 2581 135 2595
rect -35 2441 -22 2581
rect 118 2441 135 2581
rect -35 2427 135 2441
rect 195 2581 365 2595
rect 195 2441 208 2581
rect 348 2441 365 2581
rect 195 2427 365 2441
rect 425 2581 595 2595
rect 425 2441 438 2581
rect 578 2441 595 2581
rect 425 2427 595 2441
rect 655 2581 825 2595
rect 655 2441 668 2581
rect 808 2441 825 2581
rect 655 2427 825 2441
rect 885 2581 1055 2595
rect 885 2441 898 2581
rect 1038 2441 1055 2581
rect 885 2427 1055 2441
rect 1115 2581 1285 2595
rect 1115 2441 1128 2581
rect 1268 2441 1285 2581
rect 1115 2427 1285 2441
rect 1345 2581 1515 2595
rect 1345 2441 1358 2581
rect 1498 2441 1515 2581
rect 1345 2427 1515 2441
rect 1575 2581 1745 2595
rect 1575 2441 1588 2581
rect 1728 2441 1745 2581
rect 1575 2427 1745 2441
rect 1805 2581 1975 2595
rect 1805 2441 1818 2581
rect 1958 2441 1975 2581
rect 1805 2427 1975 2441
rect 2035 2581 2205 2595
rect 2035 2441 2048 2581
rect 2188 2441 2205 2581
rect 2035 2427 2205 2441
rect 2265 2581 2435 2595
rect 2265 2441 2278 2581
rect 2418 2441 2435 2581
rect 2265 2427 2435 2441
rect 2495 2581 2665 2595
rect 2495 2441 2508 2581
rect 2648 2441 2665 2581
rect 2495 2427 2665 2441
rect 2725 2581 2895 2595
rect 2725 2441 2738 2581
rect 2878 2441 2895 2581
rect 2725 2427 2895 2441
rect 2955 2581 3125 2595
rect 2955 2441 2968 2581
rect 3108 2441 3125 2581
rect 2955 2427 3125 2441
rect 3185 2581 3355 2595
rect 3185 2441 3198 2581
rect 3338 2441 3355 2581
rect 3185 2427 3355 2441
rect 3415 2581 3585 2595
rect 3415 2441 3428 2581
rect 3568 2441 3585 2581
rect 3415 2427 3585 2441
rect 3645 2581 3815 2595
rect 3645 2441 3658 2581
rect 3798 2441 3815 2581
rect 3645 2427 3815 2441
rect 3875 2581 4045 2595
rect 3875 2441 3888 2581
rect 4028 2441 4045 2581
rect 3875 2427 4045 2441
rect 4105 2581 4275 2595
rect 4105 2441 4118 2581
rect 4258 2441 4275 2581
rect 4105 2427 4275 2441
<< psubdiffcont >>
rect -1737 5467 -1691 5513
rect -1470 5467 -1424 5513
rect -1260 5467 -1214 5513
rect -1050 5467 -1004 5513
rect -840 5467 -794 5513
rect -630 5467 -584 5513
rect -420 5467 -374 5513
rect -210 5467 -164 5513
rect 401 5470 447 5516
rect 611 5470 657 5516
rect 821 5470 867 5516
rect 1031 5470 1077 5516
rect 1241 5470 1287 5516
rect 1451 5470 1497 5516
rect 1661 5470 1707 5516
rect 1871 5470 1917 5516
rect 2081 5470 2127 5516
rect 2291 5470 2337 5516
rect 2501 5470 2547 5516
rect 2711 5470 2757 5516
rect 2921 5470 2967 5516
rect 3131 5470 3177 5516
rect 3341 5470 3387 5516
rect 3551 5470 3597 5516
rect 3761 5470 3807 5516
rect -1596 4466 -1550 4512
rect -1386 4466 -1340 4512
rect -1176 4466 -1130 4512
rect -966 4466 -920 4512
rect -756 4466 -710 4512
rect -546 4466 -500 4512
rect -336 4466 -290 4512
rect -126 4466 -80 4512
rect 401 4451 447 4497
rect 611 4451 657 4497
rect 821 4451 867 4497
rect 1031 4451 1077 4497
rect 1241 4451 1287 4497
rect 1451 4451 1497 4497
rect 1661 4451 1707 4497
rect 1871 4451 1917 4497
rect 2081 4451 2127 4497
rect 2291 4451 2337 4497
rect 2501 4451 2547 4497
rect 2711 4451 2757 4497
rect 2921 4451 2967 4497
rect 3131 4451 3177 4497
rect 3341 4451 3387 4497
rect 3551 4451 3597 4497
rect 3761 4451 3807 4497
rect 41 2262 87 2308
rect 251 2262 297 2308
rect 461 2262 507 2308
rect 671 2262 717 2308
rect 881 2262 927 2308
rect 1091 2262 1137 2308
rect 1301 2262 1347 2308
rect 1511 2262 1557 2308
rect 1721 2262 1767 2308
rect 1931 2262 1977 2308
rect 2141 2262 2187 2308
rect 2351 2262 2397 2308
rect 2561 2262 2607 2308
rect 2771 2262 2817 2308
rect 2981 2262 3027 2308
rect 3191 2262 3237 2308
rect 3401 2262 3447 2308
rect 3611 2262 3657 2308
rect 3821 2262 3867 2308
rect 4031 2262 4077 2308
rect 41 1047 87 1093
rect 251 1047 297 1093
rect 461 1047 507 1093
rect 671 1047 717 1093
rect 881 1047 927 1093
rect 1091 1047 1137 1093
rect 1301 1047 1347 1093
rect 1511 1047 1557 1093
rect 1721 1047 1767 1093
rect 1931 1047 1977 1093
rect 2141 1047 2187 1093
rect 2351 1047 2397 1093
rect 2561 1047 2607 1093
rect 2771 1047 2817 1093
rect 2981 1047 3027 1093
rect 3191 1047 3237 1093
rect 3401 1047 3447 1093
rect 3611 1047 3657 1093
rect 3821 1047 3867 1093
rect 4031 1047 4077 1093
rect 41 -158 87 -112
rect 251 -158 297 -112
rect 461 -158 507 -112
rect 671 -158 717 -112
rect 881 -158 927 -112
rect 1091 -158 1137 -112
rect 1301 -158 1347 -112
rect 1511 -158 1557 -112
rect 1721 -158 1767 -112
rect 1931 -158 1977 -112
rect 2141 -158 2187 -112
rect 2351 -158 2397 -112
rect 2561 -158 2607 -112
rect 2771 -158 2817 -112
rect 2981 -158 3027 -112
rect 3191 -158 3237 -112
rect 3401 -158 3447 -112
rect 3611 -158 3657 -112
rect 3821 -158 3867 -112
rect 4031 -158 4077 -112
<< nsubdiffcont >>
rect -1745 6892 -1605 7032
rect -1515 6892 -1375 7032
rect -1285 6892 -1145 7032
rect -1055 6892 -915 7032
rect -825 6892 -685 7032
rect -595 6892 -455 7032
rect -365 6892 -225 7032
rect -120 6892 20 7032
rect 433 6186 573 6326
rect 663 6186 803 6326
rect 893 6186 1033 6326
rect 1123 6186 1263 6326
rect 1353 6186 1493 6326
rect 1583 6186 1723 6326
rect 1813 6186 1953 6326
rect 2043 6186 2183 6326
rect 2273 6186 2413 6326
rect 2503 6186 2643 6326
rect 2733 6186 2873 6326
rect 2963 6186 3103 6326
rect 3193 6186 3333 6326
rect 3423 6186 3563 6326
rect 3653 6186 3793 6326
rect -1745 5702 -1605 5842
rect -1515 5702 -1375 5842
rect -1285 5702 -1145 5842
rect -1055 5702 -915 5842
rect -825 5702 -685 5842
rect -595 5702 -455 5842
rect -365 5702 -225 5842
rect -120 5702 20 5842
rect -22 3736 118 3876
rect 208 3736 348 3876
rect 438 3736 578 3876
rect 668 3736 808 3876
rect 898 3736 1038 3876
rect 1128 3736 1268 3876
rect 1358 3736 1498 3876
rect 1588 3736 1728 3876
rect 1818 3736 1958 3876
rect 2048 3736 2188 3876
rect 2278 3736 2418 3876
rect 2508 3736 2648 3876
rect 2738 3736 2878 3876
rect 2968 3736 3108 3876
rect 3198 3736 3338 3876
rect 3428 3736 3568 3876
rect 3658 3736 3798 3876
rect 3888 3736 4028 3876
rect 4118 3736 4258 3876
rect -22 2441 118 2581
rect 208 2441 348 2581
rect 438 2441 578 2581
rect 668 2441 808 2581
rect 898 2441 1038 2581
rect 1128 2441 1268 2581
rect 1358 2441 1498 2581
rect 1588 2441 1728 2581
rect 1818 2441 1958 2581
rect 2048 2441 2188 2581
rect 2278 2441 2418 2581
rect 2508 2441 2648 2581
rect 2738 2441 2878 2581
rect 2968 2441 3108 2581
rect 3198 2441 3338 2581
rect 3428 2441 3568 2581
rect 3658 2441 3798 2581
rect 3888 2441 4028 2581
rect 4118 2441 4258 2581
<< polysilicon >>
rect -1635 6793 -107 6815
rect -1635 6762 -221 6793
rect -1635 6701 -1536 6762
rect -1635 6657 -1535 6701
rect -1023 6657 -923 6762
rect -819 6657 -719 6762
rect -240 6747 -221 6762
rect -175 6747 -107 6793
rect -240 6726 -107 6747
rect -207 6657 -107 6726
rect -1431 6310 -1331 6518
rect -1227 6310 -1127 6499
rect -615 6310 -515 6511
rect -411 6310 -311 6514
rect -1635 6270 -107 6310
rect -1635 6221 -1536 6270
rect -1635 6177 -1535 6221
rect -1023 6177 -923 6270
rect -819 6177 -719 6270
rect -1431 6007 -1331 6059
rect -1456 5982 -1331 6007
rect -1456 5936 -1428 5982
rect -1382 5958 -1331 5982
rect -1227 5958 -1127 6059
rect -615 5958 -515 6059
rect -411 5958 -311 6059
rect -1382 5936 -311 5958
rect -207 6012 -107 6270
rect -207 5966 -180 6012
rect -134 5966 -107 6012
rect -207 5940 -107 5966
rect 534 6061 3694 6097
rect 534 6015 603 6061
rect 649 6015 685 6061
rect 534 5979 685 6015
rect 1095 6015 1131 6061
rect 1177 6015 1246 6061
rect 1095 5979 1246 6015
rect -1456 5919 -311 5936
rect 534 5935 634 5979
rect 1146 5935 1246 5979
rect 1350 6015 1419 6061
rect 1465 6015 1501 6061
rect 1350 5979 1501 6015
rect 1911 6015 1947 6061
rect 1993 6015 2062 6061
rect 1911 5979 2062 6015
rect 1350 5935 1450 5979
rect 1962 5935 2062 5979
rect 2166 6015 2235 6061
rect 2281 6015 2317 6061
rect 2166 5979 2317 6015
rect 2727 6015 2763 6061
rect 2809 6015 2878 6061
rect 2727 5979 2878 6015
rect 2166 5935 2266 5979
rect 2778 5935 2878 5979
rect 2982 6015 3051 6061
rect 3097 6015 3133 6061
rect 2982 5979 3133 6015
rect 3545 6015 3581 6061
rect 3627 6015 3694 6061
rect 3545 5979 3694 6015
rect 2982 5935 3082 5979
rect 3594 5935 3694 5979
rect -1456 5918 -1374 5919
rect 738 5712 838 5815
rect 942 5749 1042 5815
rect 942 5712 969 5749
rect 738 5703 969 5712
rect 1015 5712 1042 5749
rect 1554 5749 1654 5815
rect 1554 5712 1581 5749
rect 1015 5703 1581 5712
rect 1627 5712 1654 5749
rect 1758 5749 1858 5815
rect 1758 5712 1785 5749
rect 1627 5703 1785 5712
rect 1831 5712 1858 5749
rect 2370 5749 2470 5815
rect 2370 5712 2397 5749
rect 1831 5703 2397 5712
rect 2443 5712 2470 5749
rect 2574 5749 2674 5815
rect 2574 5712 2601 5749
rect 2443 5703 2601 5712
rect 2647 5712 2674 5749
rect 3186 5749 3286 5815
rect 3186 5712 3213 5749
rect 2647 5703 3213 5712
rect 3259 5712 3286 5749
rect 3390 5749 3490 5815
rect 3390 5712 3417 5749
rect 3259 5703 3417 5712
rect 3463 5703 3490 5749
rect 738 5676 3490 5703
rect -1678 5360 508 5363
rect -1678 5338 3771 5360
rect -1678 5310 492 5338
rect -1678 5249 -1579 5310
rect -1066 5249 -966 5310
rect -862 5249 -762 5310
rect -250 5249 -150 5310
rect 472 5292 492 5310
rect 538 5333 3771 5338
rect 538 5324 1111 5333
rect 538 5292 572 5324
rect 472 5260 572 5292
rect 1084 5287 1111 5324
rect 1157 5324 1927 5333
rect 1157 5287 1184 5324
rect 1084 5260 1184 5287
rect 1288 5272 1388 5324
rect 1900 5287 1927 5324
rect 1973 5324 3771 5333
rect 1973 5287 2000 5324
rect 1900 5260 2000 5287
rect 2243 5228 2343 5324
rect 2855 5228 2955 5324
rect 3059 5228 3159 5324
rect 3671 5228 3771 5324
rect -1474 4992 -1374 5041
rect -1270 4992 -1170 5042
rect -658 4992 -558 5043
rect -454 4992 -354 5043
rect 676 5041 776 5071
rect 676 5007 696 5041
rect 472 4995 696 5007
rect 742 5007 776 5041
rect 880 5068 980 5071
rect 880 5064 894 5068
rect 880 5041 980 5064
rect 880 5007 908 5041
rect 742 4995 908 5007
rect 954 5007 980 5041
rect 1492 5044 1592 5071
rect 1492 5007 1519 5044
rect 954 4998 1519 5007
rect 1565 5007 1592 5044
rect 1696 5044 1796 5071
rect 1696 5007 1723 5044
rect 1565 4998 1723 5007
rect 1769 5007 1796 5044
rect 2447 5007 2547 5108
rect 2651 5007 2751 5108
rect 3263 5007 3363 5108
rect 3467 5007 3567 5108
rect 1769 4998 3771 5007
rect 954 4995 3771 4998
rect 472 4992 3771 4995
rect -1678 4971 3771 4992
rect -1678 4952 572 4971
rect -1678 4903 -1579 4952
rect -1678 4859 -1578 4903
rect -1066 4859 -966 4952
rect -862 4859 -762 4952
rect -250 4911 572 4952
rect -250 4859 -150 4911
rect 472 4875 572 4911
rect 1084 4875 1184 4971
rect 1288 4875 1388 4971
rect 1900 4875 2000 4971
rect 2243 4875 2343 4971
rect 2855 4875 2955 4971
rect 3059 4875 3159 4971
rect 3671 4875 3771 4971
rect 676 4721 776 4723
rect 676 4714 771 4721
rect 676 4696 776 4714
rect -1474 4638 -1374 4695
rect -1270 4638 -1170 4695
rect -658 4638 -558 4695
rect -454 4638 -354 4695
rect 676 4659 703 4696
rect -75 4650 703 4659
rect 749 4659 776 4696
rect 880 4659 980 4711
rect 1492 4659 1592 4711
rect 1696 4696 1796 4723
rect 1696 4659 1723 4696
rect 749 4650 1723 4659
rect 1769 4659 1796 4696
rect 2447 4659 2547 4755
rect 2651 4659 2751 4755
rect 3263 4659 3363 4755
rect 3467 4659 3567 4755
rect 1769 4650 3567 4659
rect -75 4638 3567 4650
rect -1474 4623 3567 4638
rect -1474 4599 784 4623
rect 112 4332 4088 4359
rect 112 4286 139 4332
rect 185 4323 4015 4332
rect 185 4286 212 4323
rect 112 4217 212 4286
rect 724 4217 824 4323
rect 928 4217 1028 4323
rect 1540 4217 1640 4323
rect 1744 4217 1844 4323
rect 2356 4217 2456 4323
rect 2560 4217 2660 4323
rect 3172 4217 3272 4323
rect 3376 4217 3476 4323
rect 3988 4286 4015 4323
rect 4061 4286 4088 4332
rect 3988 4217 4088 4286
rect 316 4014 416 4117
rect 520 4014 620 4117
rect 1132 4051 1232 4117
rect 1132 4014 1159 4051
rect 316 4005 1159 4014
rect 1205 4014 1232 4051
rect 1336 4014 1436 4117
rect 1948 4014 2048 4117
rect 2152 4014 2252 4117
rect 2764 4051 2864 4117
rect 2764 4014 2791 4051
rect 1205 4005 2791 4014
rect 2837 4014 2864 4051
rect 2968 4014 3068 4117
rect 3580 4014 3680 4117
rect 3784 4014 3884 4117
rect 2837 4005 3884 4014
rect 316 3978 3884 4005
rect 112 3637 4088 3663
rect 112 3591 192 3637
rect 238 3627 705 3637
rect 238 3591 264 3627
rect 112 3565 264 3591
rect 679 3591 705 3627
rect 751 3627 1009 3637
rect 751 3591 824 3627
rect 679 3565 824 3591
rect 112 3521 212 3565
rect 724 3521 824 3565
rect 928 3591 1009 3627
rect 1055 3627 1516 3637
rect 1055 3591 1081 3627
rect 928 3565 1081 3591
rect 1490 3591 1516 3627
rect 1562 3627 1825 3637
rect 1562 3591 1640 3627
rect 1490 3565 1640 3591
rect 928 3521 1028 3565
rect 1540 3521 1640 3565
rect 1744 3591 1825 3627
rect 1871 3627 2332 3637
rect 1871 3591 1897 3627
rect 1744 3565 1897 3591
rect 2306 3591 2332 3627
rect 2378 3627 2640 3637
rect 2378 3591 2456 3627
rect 2306 3565 2456 3591
rect 1744 3521 1844 3565
rect 2356 3521 2456 3565
rect 2560 3591 2640 3627
rect 2686 3627 3146 3637
rect 2686 3591 2712 3627
rect 2560 3565 2712 3591
rect 3120 3591 3146 3627
rect 3192 3627 3455 3637
rect 3192 3591 3272 3627
rect 3120 3565 3272 3591
rect 2560 3521 2660 3565
rect 3172 3521 3272 3565
rect 3376 3591 3455 3627
rect 3501 3627 3959 3637
rect 3501 3591 3527 3627
rect 3376 3565 3527 3591
rect 3933 3591 3959 3627
rect 4005 3591 4088 3637
rect 3933 3565 4088 3591
rect 3376 3521 3476 3565
rect 3988 3521 4088 3565
rect 316 3210 416 3321
rect 520 3210 620 3321
rect 316 3179 620 3210
rect 316 3173 429 3179
rect 112 3133 429 3173
rect 475 3173 620 3179
rect 1132 3215 1232 3321
rect 1336 3215 1436 3321
rect 1132 3181 1436 3215
rect 1132 3173 1262 3181
rect 475 3139 1262 3173
rect 475 3133 848 3139
rect 112 3102 848 3133
rect 112 2996 212 3102
rect 724 3093 848 3102
rect 894 3135 1262 3139
rect 1308 3173 1436 3181
rect 1948 3213 2048 3321
rect 2152 3213 2252 3321
rect 1948 3180 2252 3213
rect 1948 3173 2075 3180
rect 1308 3137 2075 3173
rect 1308 3135 1676 3137
rect 894 3102 1676 3135
rect 894 3093 1028 3102
rect 724 3060 1028 3093
rect 724 2996 824 3060
rect 928 2996 1028 3060
rect 1540 3091 1676 3102
rect 1722 3134 2075 3137
rect 2121 3173 2252 3180
rect 2764 3217 2864 3321
rect 2968 3217 3068 3321
rect 2764 3182 3068 3217
rect 2764 3173 2891 3182
rect 2121 3140 2891 3173
rect 2121 3134 2472 3140
rect 1722 3102 2472 3134
rect 1722 3091 1844 3102
rect 1540 3056 1844 3091
rect 1540 2996 1640 3056
rect 1744 2996 1844 3056
rect 2356 3094 2472 3102
rect 2518 3136 2891 3140
rect 2937 3173 3068 3182
rect 3580 3215 3680 3321
rect 3784 3215 3884 3321
rect 3580 3181 3884 3215
rect 3580 3173 3719 3181
rect 2937 3139 3719 3173
rect 2937 3136 3303 3139
rect 2518 3102 3303 3136
rect 2518 3094 2660 3102
rect 2356 3061 2660 3094
rect 2356 2996 2456 3061
rect 2560 2996 2660 3061
rect 3172 3093 3303 3102
rect 3349 3135 3719 3139
rect 3765 3173 3884 3181
rect 3765 3135 4088 3173
rect 3349 3102 4088 3135
rect 3349 3093 3476 3102
rect 3172 3059 3476 3093
rect 3172 2996 3272 3059
rect 3376 2996 3476 3059
rect 3988 2996 4088 3102
rect 316 2752 416 2796
rect 264 2727 416 2752
rect 264 2681 288 2727
rect 334 2693 416 2727
rect 520 2752 620 2796
rect 1132 2752 1232 2796
rect 520 2727 673 2752
rect 520 2693 602 2727
rect 334 2681 602 2693
rect 648 2693 673 2727
rect 1079 2727 1232 2752
rect 1079 2693 1103 2727
rect 648 2681 1103 2693
rect 1149 2693 1232 2727
rect 1336 2752 1436 2796
rect 1948 2752 2048 2796
rect 1336 2727 1486 2752
rect 1336 2693 1415 2727
rect 1149 2681 1415 2693
rect 1461 2693 1486 2727
rect 1900 2727 2048 2752
rect 1900 2693 1924 2727
rect 1461 2681 1924 2693
rect 1970 2693 2048 2727
rect 2152 2752 2252 2796
rect 2764 2752 2864 2796
rect 2152 2727 2305 2752
rect 2152 2693 2234 2727
rect 1970 2681 2234 2693
rect 2280 2693 2305 2727
rect 2714 2727 2864 2752
rect 2714 2693 2738 2727
rect 2280 2681 2738 2693
rect 2784 2693 2864 2727
rect 2968 2752 3068 2796
rect 2968 2727 3121 2752
rect 3580 2748 3680 2796
rect 2968 2693 3050 2727
rect 2784 2681 3050 2693
rect 3096 2693 3121 2727
rect 3527 2725 3680 2748
rect 3527 2693 3549 2725
rect 3096 2681 3549 2693
rect 264 2679 3549 2681
rect 3595 2693 3680 2725
rect 3784 2752 3884 2796
rect 3784 2727 3936 2752
rect 3784 2693 3865 2727
rect 3595 2681 3865 2693
rect 3911 2681 3936 2727
rect 3595 2679 3936 2681
rect 264 2657 3936 2679
rect 112 2117 4088 2144
rect 112 2108 1771 2117
rect 112 2046 212 2108
rect 724 2046 824 2108
rect 928 2046 1028 2108
rect 1540 2046 1640 2108
rect 1744 2071 1771 2108
rect 1817 2115 4088 2117
rect 1817 2108 2383 2115
rect 1817 2071 1844 2108
rect 1744 2044 1844 2071
rect 2356 2069 2383 2108
rect 2429 2108 4088 2115
rect 2429 2069 2456 2108
rect 2356 2042 2456 2069
rect 2560 2046 2660 2108
rect 3172 2046 3272 2108
rect 3376 2046 3476 2108
rect 3988 2046 4088 2108
rect 316 1693 416 1758
rect 520 1693 620 1758
rect 1132 1693 1232 1758
rect 1336 1693 1436 1758
rect 1948 1693 2048 1758
rect 2152 1693 2252 1758
rect 2764 1693 2864 1758
rect 2968 1693 3068 1758
rect 3580 1693 3680 1758
rect 3784 1693 3884 1758
rect -151 1657 4354 1693
rect -151 1579 -115 1657
rect -181 1561 -92 1579
rect -181 1515 -161 1561
rect -115 1515 -92 1561
rect 112 1551 212 1657
rect 724 1551 824 1657
rect 928 1551 1028 1657
rect 1540 1551 1640 1657
rect 1744 1551 1844 1657
rect 2356 1551 2456 1657
rect 2560 1551 2660 1657
rect 3172 1551 3272 1657
rect 3376 1551 3476 1657
rect 3988 1551 4088 1657
rect 4318 1598 4354 1657
rect 4296 1578 4385 1598
rect 4296 1532 4317 1578
rect 4363 1532 4385 1578
rect 4296 1515 4385 1532
rect -181 1498 -92 1515
rect 316 1248 416 1307
rect 520 1248 620 1307
rect 1132 1248 1232 1307
rect 1336 1285 1436 1312
rect 1336 1248 1363 1285
rect 316 1239 1363 1248
rect 1409 1248 1436 1285
rect 1948 1248 2048 1307
rect 2152 1285 2252 1312
rect 2152 1248 2179 1285
rect 1409 1239 2179 1248
rect 2225 1248 2252 1285
rect 2764 1285 2864 1312
rect 2764 1248 2791 1285
rect 2225 1239 2791 1248
rect 2837 1248 2864 1285
rect 2968 1248 3068 1307
rect 3580 1248 3680 1307
rect 3784 1248 3884 1307
rect 2837 1239 3884 1248
rect 316 1212 3884 1239
rect 112 902 4088 929
rect 112 856 139 902
rect 185 901 955 902
rect 185 893 751 901
rect 185 856 212 893
rect 112 829 212 856
rect 724 855 751 893
rect 797 893 955 901
rect 797 855 824 893
rect 724 828 824 855
rect 928 856 955 893
rect 1001 893 1567 902
rect 1001 856 1028 893
rect 928 829 1028 856
rect 1540 856 1567 893
rect 1613 893 1771 902
rect 1613 856 1640 893
rect 1540 829 1640 856
rect 1744 856 1771 893
rect 1817 893 2383 902
rect 1817 856 1844 893
rect 1744 829 1844 856
rect 2356 856 2383 893
rect 2429 893 2587 902
rect 2429 856 2456 893
rect 2356 829 2456 856
rect 2560 856 2587 893
rect 2633 893 3199 902
rect 2633 856 2660 893
rect 2560 829 2660 856
rect 3172 856 3199 893
rect 3245 893 3403 902
rect 3245 856 3272 893
rect 3172 829 3272 856
rect 3376 856 3403 893
rect 3449 893 4015 902
rect 3449 856 3476 893
rect 3376 829 3476 856
rect 3988 856 4015 893
rect 4061 856 4088 902
rect 3988 829 4088 856
rect 316 518 416 545
rect 316 481 343 518
rect 112 472 343 481
rect 389 481 416 518
rect 520 518 620 545
rect 520 481 547 518
rect 389 472 547 481
rect 593 481 620 518
rect 1132 518 1232 545
rect 1132 481 1159 518
rect 593 472 1159 481
rect 1205 481 1232 518
rect 1336 518 1436 545
rect 1336 481 1363 518
rect 1205 472 1363 481
rect 1409 481 1436 518
rect 1948 518 2048 545
rect 1948 481 1975 518
rect 1409 472 1975 481
rect 2021 481 2048 518
rect 2152 518 2252 545
rect 2152 481 2179 518
rect 2021 472 2179 481
rect 2225 481 2252 518
rect 2764 518 2864 545
rect 2764 481 2791 518
rect 2225 472 2791 481
rect 2837 481 2864 518
rect 2968 518 3068 545
rect 2968 481 2995 518
rect 2837 472 2995 481
rect 3041 481 3068 518
rect 3580 518 3680 545
rect 3580 481 3607 518
rect 3041 472 3607 481
rect 3653 481 3680 518
rect 3784 518 3884 545
rect 3784 481 3811 518
rect 3653 472 3811 481
rect 3857 481 3884 518
rect 3857 472 4088 481
rect 112 454 4088 472
rect 112 445 751 454
rect 112 339 212 445
rect 724 408 751 445
rect 797 445 955 454
rect 797 408 824 445
rect 724 339 824 408
rect 928 408 955 445
rect 1001 445 1567 454
rect 1001 408 1028 445
rect 928 339 1028 408
rect 1540 408 1567 445
rect 1613 445 1771 454
rect 1613 408 1640 445
rect 1540 339 1640 408
rect 1744 408 1771 445
rect 1817 445 2383 454
rect 1817 408 1844 445
rect 1744 339 1844 408
rect 2356 408 2383 445
rect 2429 445 2587 454
rect 2429 408 2456 445
rect 2356 339 2456 408
rect 2560 408 2587 445
rect 2633 445 3199 454
rect 2633 408 2660 445
rect 2560 339 2660 408
rect 3172 408 3199 445
rect 3245 445 3403 454
rect 3245 408 3272 445
rect 3172 339 3272 408
rect 3376 408 3403 445
rect 3449 445 4088 454
rect 3449 408 3476 445
rect 3376 339 3476 408
rect 3988 339 4088 445
rect 316 73 416 100
rect 316 27 343 73
rect 389 36 416 73
rect 520 73 620 100
rect 520 36 547 73
rect 389 27 547 36
rect 593 36 620 73
rect 1132 73 1232 100
rect 1132 36 1159 73
rect 593 27 1159 36
rect 1205 36 1232 73
rect 1336 73 1436 100
rect 1336 36 1363 73
rect 1205 27 1363 36
rect 1409 36 1436 73
rect 1948 73 2048 100
rect 1948 36 1975 73
rect 1409 27 1975 36
rect 2021 36 2048 73
rect 2152 73 2252 100
rect 2152 36 2179 73
rect 2021 27 2179 36
rect 2225 36 2252 73
rect 2764 73 2864 100
rect 2764 36 2791 73
rect 2225 27 2791 36
rect 2837 36 2864 73
rect 2968 73 3068 100
rect 2968 36 2995 73
rect 2837 27 2995 36
rect 3041 36 3068 73
rect 3580 73 3680 100
rect 3580 36 3607 73
rect 3041 27 3607 36
rect 3653 36 3680 73
rect 3784 73 3884 100
rect 3784 36 3811 73
rect 3653 27 3811 36
rect 3857 27 3884 73
rect 316 0 3884 27
<< polycontact >>
rect -221 6747 -175 6793
rect -1428 5936 -1382 5982
rect -180 5966 -134 6012
rect 603 6015 649 6061
rect 1131 6015 1177 6061
rect 1419 6015 1465 6061
rect 1947 6015 1993 6061
rect 2235 6015 2281 6061
rect 2763 6015 2809 6061
rect 3051 6015 3097 6061
rect 3581 6015 3627 6061
rect 969 5703 1015 5749
rect 1581 5703 1627 5749
rect 1785 5703 1831 5749
rect 2397 5703 2443 5749
rect 2601 5703 2647 5749
rect 3213 5703 3259 5749
rect 3417 5703 3463 5749
rect 492 5292 538 5338
rect 1111 5287 1157 5333
rect 1927 5287 1973 5333
rect 696 4995 742 5041
rect 908 4995 954 5041
rect 1519 4998 1565 5044
rect 1723 4998 1769 5044
rect 703 4650 749 4696
rect 1723 4650 1769 4696
rect 139 4286 185 4332
rect 4015 4286 4061 4332
rect 1159 4005 1205 4051
rect 2791 4005 2837 4051
rect 192 3591 238 3637
rect 705 3591 751 3637
rect 1009 3591 1055 3637
rect 1516 3591 1562 3637
rect 1825 3591 1871 3637
rect 2332 3591 2378 3637
rect 2640 3591 2686 3637
rect 3146 3591 3192 3637
rect 3455 3591 3501 3637
rect 3959 3591 4005 3637
rect 429 3133 475 3179
rect 848 3093 894 3139
rect 1262 3135 1308 3181
rect 1676 3091 1722 3137
rect 2075 3134 2121 3180
rect 2472 3094 2518 3140
rect 2891 3136 2937 3182
rect 3303 3093 3349 3139
rect 3719 3135 3765 3181
rect 288 2681 334 2727
rect 602 2681 648 2727
rect 1103 2681 1149 2727
rect 1415 2681 1461 2727
rect 1924 2681 1970 2727
rect 2234 2681 2280 2727
rect 2738 2681 2784 2727
rect 3050 2681 3096 2727
rect 3549 2679 3595 2725
rect 3865 2681 3911 2727
rect 1771 2071 1817 2117
rect 2383 2069 2429 2115
rect -161 1515 -115 1561
rect 4317 1532 4363 1578
rect 1363 1239 1409 1285
rect 2179 1239 2225 1285
rect 2791 1239 2837 1285
rect 139 856 185 902
rect 751 855 797 901
rect 955 856 1001 902
rect 1567 856 1613 902
rect 1771 856 1817 902
rect 2383 856 2429 902
rect 2587 856 2633 902
rect 3199 856 3245 902
rect 3403 856 3449 902
rect 4015 856 4061 902
rect 343 472 389 518
rect 547 472 593 518
rect 1159 472 1205 518
rect 1363 472 1409 518
rect 1975 472 2021 518
rect 2179 472 2225 518
rect 2791 472 2837 518
rect 2995 472 3041 518
rect 3607 472 3653 518
rect 3811 472 3857 518
rect 751 408 797 454
rect 955 408 1001 454
rect 1567 408 1613 454
rect 1771 408 1817 454
rect 2383 408 2429 454
rect 2587 408 2633 454
rect 3199 408 3245 454
rect 3403 408 3449 454
rect 343 27 389 73
rect 547 27 593 73
rect 1159 27 1205 73
rect 1363 27 1409 73
rect 1975 27 2021 73
rect 2179 27 2225 73
rect 2791 27 2837 73
rect 2995 27 3041 73
rect 3607 27 3653 73
rect 3811 27 3857 73
<< metal1 >>
rect -1809 7032 314 7070
rect -1809 6892 -1745 7032
rect -1605 6892 -1515 7032
rect -1375 6892 -1285 7032
rect -1145 6892 -1055 7032
rect -915 6892 -825 7032
rect -685 6892 -595 7032
rect -455 6892 -365 7032
rect -225 6892 -120 7032
rect 20 6892 314 7032
rect -1809 6878 314 6892
rect -1710 6655 -1664 6878
rect -894 6655 -848 6878
rect -238 6796 -164 6811
rect -238 6744 -224 6796
rect -172 6744 -164 6796
rect -238 6729 -164 6744
rect -78 6655 -32 6878
rect -1527 6626 -1450 6637
rect -1527 6574 -1513 6626
rect -1461 6574 -1450 6626
rect -1527 6560 -1450 6574
rect -1116 6625 -1039 6636
rect -1116 6573 -1102 6625
rect -1050 6573 -1039 6625
rect -1116 6559 -1039 6573
rect -708 6625 -631 6636
rect -708 6573 -694 6625
rect -642 6573 -631 6625
rect -708 6559 -631 6573
rect -302 6625 -225 6636
rect -302 6573 -288 6625
rect -236 6573 -225 6625
rect -302 6559 -225 6573
rect -1302 6413 -1256 6539
rect -487 6413 -441 6557
rect -1992 6316 -32 6413
rect -1710 6175 -1664 6316
rect -894 6175 -848 6316
rect -78 6175 -32 6316
rect 166 6364 314 6878
rect 166 6326 3868 6364
rect 166 6186 433 6326
rect 573 6186 663 6326
rect 803 6186 893 6326
rect 1033 6186 1123 6326
rect 1263 6186 1353 6326
rect 1493 6186 1583 6326
rect 1723 6186 1813 6326
rect 1953 6186 2043 6326
rect 2183 6186 2273 6326
rect 2413 6186 2503 6326
rect 2643 6186 2733 6326
rect 2873 6186 2963 6326
rect 3103 6186 3193 6326
rect 3333 6186 3423 6326
rect 3563 6186 3653 6326
rect 3793 6324 3868 6326
rect 3793 6226 4230 6324
rect 3793 6186 3868 6226
rect 166 6172 3868 6186
rect -1527 6158 -1450 6169
rect -1527 6106 -1513 6158
rect -1461 6106 -1450 6158
rect -1527 6092 -1450 6106
rect -1116 6144 -1039 6155
rect -1116 6092 -1102 6144
rect -1050 6092 -1039 6144
rect -1116 6078 -1039 6092
rect -711 6144 -634 6155
rect -711 6092 -697 6144
rect -645 6092 -634 6144
rect -711 6078 -634 6092
rect -302 6154 -225 6165
rect -302 6102 -288 6154
rect -236 6102 -225 6154
rect -302 6088 -225 6102
rect -1441 5985 -1368 6004
rect -1441 5933 -1428 5985
rect -1376 5933 -1368 5985
rect -1441 5914 -1368 5933
rect -1302 5856 -1256 6078
rect -486 5856 -440 6075
rect -193 6017 -116 6032
rect -193 6012 -177 6017
rect -193 5966 -180 6012
rect -193 5965 -177 5966
rect -125 5965 -116 6017
rect -193 5947 -116 5965
rect 166 5856 314 6172
rect 459 5933 505 6172
rect 572 6079 680 6092
rect 1100 6079 1208 6092
rect 572 6064 1208 6079
rect 572 6012 599 6064
rect 651 6061 1208 6064
rect 651 6033 1131 6061
rect 651 6012 709 6033
rect 572 5984 709 6012
rect -1809 5842 314 5856
rect -1809 5702 -1745 5842
rect -1605 5702 -1515 5842
rect -1375 5702 -1285 5842
rect -1145 5702 -1055 5842
rect -915 5702 -825 5842
rect -685 5702 -595 5842
rect -455 5702 -365 5842
rect -225 5702 -120 5842
rect 20 5708 314 5842
rect 663 5812 709 5984
rect 1071 6015 1131 6033
rect 1177 6015 1208 6061
rect 1071 5984 1208 6015
rect 1071 5933 1117 5984
rect 1275 5933 1321 6172
rect 1388 6073 1496 6092
rect 1916 6073 2024 6092
rect 1388 6061 2024 6073
rect 1388 6015 1419 6061
rect 1465 6027 1947 6061
rect 1465 6015 1525 6027
rect 1388 5984 1525 6015
rect 1479 5933 1525 5984
rect 1887 6015 1947 6027
rect 1993 6015 2024 6061
rect 1887 5984 2024 6015
rect 1887 5933 1933 5984
rect 2091 5933 2137 6172
rect 2204 6070 2312 6092
rect 2732 6070 2840 6092
rect 2204 6061 2840 6070
rect 2204 6015 2235 6061
rect 2281 6024 2763 6061
rect 2281 6015 2341 6024
rect 2204 5984 2341 6015
rect 2295 5933 2341 5984
rect 2703 6015 2763 6024
rect 2809 6015 2840 6061
rect 2703 5984 2840 6015
rect 2703 5933 2749 5984
rect 2907 5933 2953 6172
rect 3020 6076 3128 6092
rect 3550 6076 3658 6092
rect 3020 6061 3658 6076
rect 3020 6015 3051 6061
rect 3097 6030 3581 6061
rect 3097 6015 3157 6030
rect 3020 5984 3157 6015
rect 3111 5933 3157 5984
rect 3519 6015 3581 6030
rect 3627 6015 3658 6061
rect 3519 5984 3658 6015
rect 3519 5933 3565 5984
rect 3723 5933 3769 6172
rect 636 5724 709 5812
rect 867 5771 913 5817
rect 1683 5771 1729 5817
rect 2499 5771 2545 5817
rect 3315 5771 3361 5817
rect 867 5749 3485 5771
rect 867 5716 969 5749
rect 20 5702 86 5708
rect -1809 5664 86 5702
rect 835 5703 969 5716
rect 1015 5725 1581 5749
rect 1015 5703 1037 5725
rect 835 5681 1037 5703
rect 1559 5703 1581 5725
rect 1627 5725 1778 5749
rect 1627 5703 1649 5725
rect 1559 5681 1649 5703
rect 1763 5697 1778 5725
rect 1831 5725 2397 5749
rect 1831 5703 1853 5725
rect 1830 5697 1853 5703
rect 1763 5681 1853 5697
rect 2375 5697 2397 5725
rect 2449 5725 2601 5749
rect 2449 5697 2465 5725
rect 2375 5681 2465 5697
rect 2579 5703 2601 5725
rect 2647 5725 3213 5749
rect 2647 5703 2669 5725
rect 2579 5681 2669 5703
rect 3191 5703 3213 5725
rect 3259 5725 3417 5749
rect 3259 5703 3281 5725
rect 3191 5681 3281 5703
rect 3395 5703 3417 5725
rect 3463 5703 3485 5749
rect 3395 5681 3485 5703
rect 835 5632 913 5681
rect 360 5562 3883 5565
rect -1793 5528 3883 5562
rect -1793 5513 395 5528
rect 447 5516 3883 5528
rect -1793 5467 -1737 5513
rect -1691 5467 -1470 5513
rect -1424 5467 -1260 5513
rect -1214 5467 -1050 5513
rect -1004 5467 -840 5513
rect -794 5467 -630 5513
rect -584 5467 -420 5513
rect -374 5467 -210 5513
rect -164 5476 395 5513
rect -164 5470 401 5476
rect 447 5470 611 5516
rect 657 5470 821 5516
rect 867 5470 1031 5516
rect 1077 5470 1241 5516
rect 1287 5470 1451 5516
rect 1497 5470 1661 5516
rect 1707 5470 1871 5516
rect 1917 5470 2081 5516
rect 2127 5470 2291 5516
rect 2337 5470 2501 5516
rect 2547 5470 2711 5516
rect 2757 5470 2921 5516
rect 2967 5470 3131 5516
rect 3177 5470 3341 5516
rect 3387 5470 3551 5516
rect 3597 5510 3761 5516
rect 3597 5470 3754 5510
rect 3807 5470 3883 5516
rect -164 5467 3754 5470
rect -1793 5458 3754 5467
rect 3806 5458 3883 5470
rect -1793 5419 3883 5458
rect -1793 5416 448 5419
rect -1345 5203 -1299 5416
rect -529 5203 -483 5416
rect 477 5338 567 5355
rect 477 5311 492 5338
rect 291 5292 492 5311
rect 538 5292 567 5338
rect 291 5265 567 5292
rect 291 5258 513 5265
rect 397 5226 443 5258
rect 805 5226 851 5419
rect 1089 5334 1179 5355
rect 1089 5282 1105 5334
rect 1157 5315 1179 5334
rect 1157 5282 1259 5315
rect 1089 5265 1259 5282
rect 1213 5226 1259 5265
rect 1621 5226 1667 5419
rect 1905 5333 1995 5355
rect 1905 5287 1927 5333
rect 1973 5311 1995 5333
rect 1973 5287 2075 5311
rect 1905 5265 2075 5287
rect 2029 5226 2075 5265
rect 2576 5226 2622 5419
rect 3392 5226 3438 5419
rect 2355 5197 2430 5210
rect -1565 5176 -1488 5187
rect -1565 5124 -1551 5176
rect -1499 5124 -1488 5176
rect -1565 5110 -1488 5124
rect -1158 5175 -1081 5186
rect -1158 5123 -1144 5175
rect -1092 5123 -1081 5175
rect -1158 5109 -1081 5123
rect -751 5175 -674 5186
rect -751 5123 -737 5175
rect -685 5123 -674 5175
rect -751 5109 -674 5123
rect -343 5175 -266 5186
rect -343 5123 -329 5175
rect -277 5123 -266 5175
rect 2355 5145 2366 5197
rect 2418 5145 2430 5197
rect -343 5109 -266 5123
rect -1753 5016 -1707 5087
rect -937 5016 -891 5087
rect -121 5016 -75 5087
rect 601 5067 647 5132
rect 601 5046 757 5067
rect 1009 5064 1055 5117
rect -1905 4948 -75 5016
rect 289 5041 757 5046
rect 289 4995 696 5041
rect 742 4995 757 5041
rect 289 4990 757 4995
rect 601 4976 757 4990
rect 890 5041 1055 5064
rect 890 4995 908 5041
rect 954 4995 1055 5041
rect -1345 4857 -1299 4948
rect -529 4857 -483 4948
rect 601 4873 647 4976
rect 890 4971 1055 4995
rect 1009 4873 1055 4971
rect 1417 5066 1463 5121
rect 1825 5066 1871 5116
rect 1417 5044 1587 5066
rect 1417 4998 1519 5044
rect 1565 4998 1587 5044
rect 1417 4976 1587 4998
rect 1701 5044 1871 5066
rect 1701 4998 1723 5044
rect 1769 4998 1871 5044
rect 2168 5043 2214 5135
rect 2355 5131 2430 5145
rect 2763 5193 2838 5206
rect 2763 5141 2774 5193
rect 2826 5141 2838 5193
rect 2763 5127 2838 5141
rect 3170 5194 3245 5207
rect 3170 5142 3181 5194
rect 3233 5142 3245 5194
rect 1701 4976 1871 4998
rect 1417 4873 1463 4976
rect 1825 4873 1871 4976
rect 2146 5023 2236 5043
rect 2146 4971 2165 5023
rect 2217 5020 2236 5023
rect 2984 5020 3030 5137
rect 3170 5128 3245 5142
rect 3580 5194 3655 5207
rect 3580 5142 3591 5194
rect 3643 5142 3655 5194
rect 3580 5128 3655 5142
rect 3800 5020 3846 5143
rect 2217 4974 3846 5020
rect 2217 4971 2236 4974
rect 2146 4953 2236 4971
rect 2576 4873 2622 4974
rect 3392 4873 3438 4974
rect 2356 4848 2431 4861
rect -1566 4830 -1489 4841
rect -1566 4778 -1552 4830
rect -1500 4778 -1489 4830
rect -1566 4764 -1489 4778
rect -1158 4830 -1081 4841
rect -1158 4778 -1144 4830
rect -1092 4778 -1081 4830
rect -1158 4764 -1081 4778
rect -751 4830 -674 4841
rect -751 4778 -737 4830
rect -685 4778 -674 4830
rect -751 4764 -674 4778
rect -343 4830 -266 4841
rect -343 4778 -329 4830
rect -277 4778 -266 4830
rect -343 4764 -266 4778
rect -1753 4561 -1707 4741
rect -937 4561 -891 4742
rect -121 4561 -75 4743
rect -1753 4514 -39 4561
rect 397 4546 443 4757
rect 805 4714 851 4764
rect 678 4696 851 4714
rect 678 4644 697 4696
rect 749 4668 851 4696
rect 749 4644 771 4668
rect 678 4626 771 4644
rect 687 4625 771 4626
rect 1213 4546 1259 4760
rect 1621 4722 1667 4757
rect 1621 4718 1743 4722
rect 1621 4696 1791 4718
rect 1621 4676 1723 4696
rect 1701 4650 1723 4676
rect 1769 4650 1791 4696
rect 1701 4628 1791 4650
rect 2029 4546 2075 4757
rect 2168 4546 2214 4826
rect 2356 4796 2367 4848
rect 2419 4796 2431 4848
rect 2356 4782 2431 4796
rect 2761 4846 2836 4859
rect 2761 4794 2772 4846
rect 2824 4794 2836 4846
rect 2761 4780 2836 4794
rect 2984 4546 3030 4861
rect 3171 4846 3246 4859
rect 3171 4794 3182 4846
rect 3234 4794 3246 4846
rect 3171 4780 3246 4794
rect 3580 4848 3655 4861
rect 3580 4796 3591 4848
rect 3643 4796 3655 4848
rect 3580 4782 3655 4796
rect 3800 4546 3846 4852
rect -1753 4512 -127 4514
rect -1753 4466 -1596 4512
rect -1550 4466 -1386 4512
rect -1340 4466 -1176 4512
rect -1130 4466 -966 4512
rect -920 4466 -756 4512
rect -710 4466 -546 4512
rect -500 4466 -336 4512
rect -290 4466 -127 4512
rect -1753 4462 -127 4466
rect -75 4462 -39 4514
rect -1753 4415 -39 4462
rect 360 4499 3883 4546
rect 360 4447 395 4499
rect 447 4497 3883 4499
rect 447 4451 611 4497
rect 657 4451 821 4497
rect 867 4451 1031 4497
rect 1077 4451 1241 4497
rect 1287 4451 1451 4497
rect 1497 4451 1661 4497
rect 1707 4451 1871 4497
rect 1917 4451 2081 4497
rect 2127 4451 2291 4497
rect 2337 4451 2501 4497
rect 2547 4451 2711 4497
rect 2757 4451 2921 4497
rect 2967 4451 3131 4497
rect 3177 4451 3341 4497
rect 3387 4451 3551 4497
rect 3597 4451 3754 4497
rect 3807 4451 3883 4497
rect 447 4447 3754 4451
rect 360 4445 3754 4447
rect 3806 4445 3883 4451
rect 360 4400 3883 4445
rect 117 4333 207 4354
rect 3993 4335 4083 4354
rect 117 4281 133 4333
rect 185 4281 207 4333
rect 117 4264 207 4281
rect 431 4323 516 4333
rect 431 4318 3755 4323
rect 431 4266 450 4318
rect 502 4266 3755 4318
rect 431 4261 3755 4266
rect 3993 4283 4011 4335
rect 4063 4283 4083 4335
rect 3993 4264 4083 4283
rect 431 4249 516 4261
rect 228 4196 301 4209
rect 228 4144 238 4196
rect 290 4144 301 4196
rect 445 4163 491 4249
rect 636 4196 709 4209
rect 228 4130 301 4144
rect 636 4144 646 4196
rect 698 4144 709 4196
rect 636 4130 709 4144
rect 1043 4196 1116 4209
rect 1043 4144 1053 4196
rect 1105 4144 1116 4196
rect 1261 4173 1307 4261
rect 1453 4196 1526 4209
rect 1043 4130 1116 4144
rect 1453 4144 1463 4196
rect 1515 4144 1526 4196
rect 1453 4130 1526 4144
rect 1859 4196 1932 4209
rect 1859 4144 1869 4196
rect 1921 4144 1932 4196
rect 2077 4161 2123 4261
rect 2265 4196 2338 4209
rect 1859 4130 1932 4144
rect 2265 4144 2275 4196
rect 2327 4144 2338 4196
rect 2265 4130 2338 4144
rect 2675 4196 2748 4209
rect 2675 4144 2685 4196
rect 2737 4144 2748 4196
rect 2893 4169 2939 4261
rect 3080 4196 3153 4209
rect 2675 4130 2748 4144
rect 3080 4144 3090 4196
rect 3142 4144 3153 4196
rect 3080 4130 3153 4144
rect 3492 4196 3565 4209
rect 3492 4144 3502 4196
rect 3554 4144 3565 4196
rect 3709 4172 3755 4261
rect 3899 4196 3972 4209
rect 3492 4130 3565 4144
rect 3899 4144 3909 4196
rect 3961 4144 3972 4196
rect 3899 4130 3972 4144
rect 4132 4119 4230 6226
rect 37 3914 83 4119
rect 853 3914 899 4119
rect 1137 4054 1227 4073
rect 1137 4002 1154 4054
rect 1206 4002 1227 4054
rect 1137 3983 1227 4002
rect 1669 3914 1715 4119
rect 2485 3914 2531 4119
rect 2769 4053 2859 4073
rect 2769 4001 2786 4053
rect 2838 4001 2859 4053
rect 2769 3983 2859 4001
rect 3301 3914 3347 4119
rect 4117 3914 4230 4119
rect -62 3876 4299 3914
rect -62 3736 -22 3876
rect 118 3736 208 3876
rect 348 3736 438 3876
rect 578 3736 668 3876
rect 808 3736 898 3876
rect 1038 3736 1128 3876
rect 1268 3736 1358 3876
rect 1498 3736 1588 3876
rect 1728 3736 1818 3876
rect 1958 3736 2048 3876
rect 2188 3736 2278 3876
rect 2418 3736 2508 3876
rect 2648 3736 2738 3876
rect 2878 3736 2968 3876
rect 3108 3736 3198 3876
rect 3338 3736 3428 3876
rect 3568 3736 3658 3876
rect 3798 3736 3888 3876
rect 4028 3736 4118 3876
rect 4258 3736 4299 3876
rect -62 3722 4299 3736
rect 37 3519 83 3722
rect 171 3639 259 3658
rect 171 3587 187 3639
rect 239 3619 259 3639
rect 684 3637 772 3658
rect 684 3619 705 3637
rect 239 3587 287 3619
rect 171 3570 287 3587
rect 241 3519 287 3570
rect 649 3591 705 3619
rect 751 3591 772 3637
rect 649 3570 772 3591
rect 649 3519 695 3570
rect 853 3519 899 3722
rect 988 3637 1076 3658
rect 988 3591 1009 3637
rect 1055 3619 1076 3637
rect 1495 3637 1583 3658
rect 1495 3619 1516 3637
rect 1055 3591 1103 3619
rect 988 3570 1103 3591
rect 1057 3519 1103 3570
rect 1465 3591 1516 3619
rect 1562 3591 1583 3637
rect 1465 3570 1583 3591
rect 1465 3519 1511 3570
rect 1669 3519 1715 3722
rect 1804 3640 1892 3658
rect 1804 3588 1819 3640
rect 1871 3619 1892 3640
rect 2311 3641 2399 3658
rect 2311 3619 2331 3641
rect 1871 3588 1919 3619
rect 1804 3570 1919 3588
rect 1873 3519 1919 3570
rect 2281 3589 2331 3619
rect 2383 3589 2399 3641
rect 2281 3570 2399 3589
rect 2281 3519 2327 3570
rect 2485 3519 2531 3722
rect 2619 3637 2707 3658
rect 2619 3591 2640 3637
rect 2686 3619 2707 3637
rect 3125 3637 3213 3658
rect 3125 3619 3146 3637
rect 2686 3591 2735 3619
rect 2619 3570 2735 3591
rect 2689 3519 2735 3570
rect 3097 3591 3146 3619
rect 3192 3591 3213 3637
rect 3097 3570 3213 3591
rect 3097 3519 3143 3570
rect 3301 3519 3347 3722
rect 3434 3637 3522 3658
rect 3434 3591 3455 3637
rect 3501 3619 3522 3637
rect 3938 3639 4026 3658
rect 3938 3619 3955 3639
rect 3501 3591 3551 3619
rect 3434 3570 3551 3591
rect 3505 3519 3551 3570
rect 3913 3587 3955 3619
rect 4007 3587 4026 3639
rect 3913 3570 4026 3587
rect 3913 3519 3959 3570
rect 4117 3519 4163 3722
rect 445 3205 491 3323
rect 1261 3210 1307 3323
rect 403 3181 501 3205
rect 1232 3183 1338 3210
rect 2077 3208 2123 3323
rect 2893 3212 2939 3323
rect 1232 3181 1258 3183
rect 1310 3181 1338 3183
rect 2046 3181 2150 3208
rect 2860 3184 2968 3212
rect 3709 3210 3755 3323
rect 2860 3181 2886 3184
rect 37 3179 1258 3181
rect 37 3135 429 3179
rect 37 2994 83 3135
rect 403 3133 429 3135
rect 475 3139 1258 3179
rect 475 3135 848 3139
rect 475 3133 501 3135
rect 403 3107 501 3133
rect 818 3093 848 3135
rect 894 3135 1258 3139
rect 1310 3180 2886 3181
rect 1310 3137 2075 3180
rect 1310 3135 1676 3137
rect 894 3093 924 3135
rect 1232 3131 1258 3135
rect 1310 3131 1338 3135
rect 1232 3107 1338 3131
rect 818 3065 924 3093
rect 1644 3091 1676 3135
rect 1722 3135 2075 3137
rect 1722 3091 1754 3135
rect 2046 3134 2075 3135
rect 2121 3140 2886 3180
rect 2121 3135 2472 3140
rect 2121 3134 2150 3135
rect 2046 3107 2150 3134
rect 853 2994 899 3065
rect 1644 3061 1754 3091
rect 2444 3094 2472 3135
rect 2518 3135 2886 3140
rect 2938 3181 2968 3184
rect 3689 3181 3795 3210
rect 2938 3139 3719 3181
rect 2518 3094 2546 3135
rect 2860 3132 2886 3135
rect 2938 3135 3303 3139
rect 2938 3132 2968 3135
rect 2860 3107 2968 3132
rect 2444 3066 2546 3094
rect 3274 3093 3303 3135
rect 3349 3135 3719 3139
rect 3765 3135 4163 3181
rect 3349 3093 3378 3135
rect 3689 3107 3795 3135
rect 1669 2994 1715 3061
rect 2485 2994 2531 3066
rect 3274 3064 3378 3093
rect 3301 2994 3347 3064
rect 4117 2994 4163 3135
rect -182 2850 60 2915
rect 4131 2856 4486 2921
rect -182 1718 -117 2850
rect 241 2747 287 2798
rect 241 2727 354 2747
rect 241 2699 288 2727
rect 269 2681 288 2699
rect 334 2681 354 2727
rect 269 2662 354 2681
rect 445 2595 491 2798
rect 649 2747 695 2798
rect 583 2727 695 2747
rect 583 2681 602 2727
rect 648 2699 695 2727
rect 1057 2747 1103 2798
rect 1057 2734 1169 2747
rect 1057 2699 1090 2734
rect 1142 2727 1169 2734
rect 648 2681 668 2699
rect 583 2662 668 2681
rect 1080 2682 1090 2699
rect 1080 2681 1103 2682
rect 1149 2681 1169 2727
rect 1080 2668 1169 2681
rect 1084 2662 1169 2668
rect 1261 2595 1307 2798
rect 1465 2747 1511 2798
rect 1396 2727 1511 2747
rect 1396 2681 1415 2727
rect 1461 2699 1511 2727
rect 1873 2747 1919 2798
rect 1873 2730 1990 2747
rect 1873 2699 1917 2730
rect 1969 2727 1990 2730
rect 1461 2681 1481 2699
rect 1396 2662 1481 2681
rect 1905 2678 1917 2699
rect 1970 2681 1990 2727
rect 1969 2678 1990 2681
rect 1905 2662 1990 2678
rect 2077 2595 2123 2798
rect 2281 2747 2327 2798
rect 2215 2727 2327 2747
rect 2215 2681 2234 2727
rect 2280 2699 2327 2727
rect 2689 2748 2735 2798
rect 2689 2747 2801 2748
rect 2689 2735 2804 2747
rect 2689 2699 2738 2735
rect 2280 2681 2300 2699
rect 2215 2662 2300 2681
rect 2719 2681 2738 2699
rect 2790 2683 2804 2735
rect 2784 2681 2804 2683
rect 2719 2662 2804 2681
rect 2893 2595 2939 2798
rect 3097 2747 3143 2798
rect 3031 2727 3143 2747
rect 3031 2681 3050 2727
rect 3096 2699 3143 2727
rect 3505 2743 3551 2798
rect 3505 2725 3613 2743
rect 3505 2699 3549 2725
rect 3096 2681 3116 2699
rect 3031 2662 3116 2681
rect 3532 2679 3549 2699
rect 3595 2679 3613 2725
rect 3532 2662 3613 2679
rect 3709 2595 3755 2798
rect 3913 2747 3959 2798
rect 3846 2727 3959 2747
rect 3846 2681 3865 2727
rect 3911 2699 3959 2727
rect 3911 2681 3931 2699
rect 3846 2662 3931 2681
rect -62 2581 4299 2595
rect -62 2441 -22 2581
rect 118 2441 208 2581
rect 348 2441 438 2581
rect 578 2441 668 2581
rect 808 2441 898 2581
rect 1038 2441 1128 2581
rect 1268 2441 1358 2581
rect 1498 2441 1588 2581
rect 1728 2441 1818 2581
rect 1958 2441 2048 2581
rect 2188 2441 2278 2581
rect 2418 2441 2508 2581
rect 2648 2441 2738 2581
rect 2878 2441 2968 2581
rect 3108 2441 3198 2581
rect 3338 2441 3428 2581
rect 3568 2441 3658 2581
rect 3798 2441 3888 2581
rect 4028 2441 4118 2581
rect 4258 2441 4299 2581
rect -62 2403 4299 2441
rect 0 2320 4200 2357
rect 0 2268 35 2320
rect 87 2308 4200 2320
rect 0 2262 41 2268
rect 87 2262 251 2308
rect 297 2262 461 2308
rect 507 2262 671 2308
rect 717 2262 881 2308
rect 927 2262 1091 2308
rect 1137 2262 1301 2308
rect 1347 2262 1511 2308
rect 1557 2262 1721 2308
rect 1767 2262 1931 2308
rect 1977 2262 2141 2308
rect 2187 2262 2351 2308
rect 2397 2262 2561 2308
rect 2607 2262 2771 2308
rect 2817 2262 2981 2308
rect 3027 2262 3191 2308
rect 3237 2262 3401 2308
rect 3447 2262 3611 2308
rect 3657 2262 3821 2308
rect 3867 2262 4023 2308
rect 4077 2262 4200 2308
rect 0 2256 4023 2262
rect 4075 2256 4200 2262
rect 0 2211 4200 2256
rect 445 2000 491 2211
rect 1261 2000 1307 2211
rect 1749 2118 1839 2139
rect 1749 2066 1765 2118
rect 1817 2066 1839 2118
rect 1749 2049 1839 2066
rect 2077 2000 2123 2211
rect 2361 2119 2451 2137
rect 2361 2067 2380 2119
rect 2432 2067 2451 2119
rect 2361 2047 2451 2067
rect 2893 2000 2939 2211
rect 3709 2000 3755 2211
rect 220 1923 293 1936
rect 220 1871 230 1923
rect 282 1871 293 1923
rect 220 1857 293 1871
rect 631 1931 704 1944
rect 631 1879 641 1931
rect 693 1879 704 1931
rect 631 1865 704 1879
rect 1038 1930 1111 1943
rect 1038 1878 1048 1930
rect 1100 1878 1111 1930
rect 1038 1864 1111 1878
rect 1448 1930 1521 1943
rect 1448 1878 1458 1930
rect 1510 1878 1521 1930
rect 1448 1864 1521 1878
rect 1854 1930 1927 1943
rect 1854 1878 1864 1930
rect 1916 1878 1927 1930
rect 1854 1864 1927 1878
rect 2264 1930 2337 1943
rect 2264 1878 2274 1930
rect 2326 1878 2337 1930
rect 2264 1864 2337 1878
rect 2671 1930 2744 1943
rect 2671 1878 2681 1930
rect 2733 1878 2744 1930
rect 2671 1864 2744 1878
rect 3076 1930 3149 1943
rect 3076 1878 3086 1930
rect 3138 1878 3149 1930
rect 3076 1864 3149 1878
rect 3486 1930 3559 1943
rect 3486 1878 3496 1930
rect 3548 1878 3559 1930
rect 3486 1864 3559 1878
rect 3897 1934 3970 1947
rect 3897 1882 3907 1934
rect 3959 1882 3970 1934
rect 3897 1868 3970 1882
rect 37 1718 83 1804
rect 853 1718 899 1809
rect 1669 1718 1715 1808
rect 2485 1718 2531 1811
rect 3301 1718 3347 1810
rect 4117 1718 4163 1807
rect 4421 1718 4486 2856
rect -182 1653 4486 1718
rect -181 1561 -92 1579
rect -181 1515 -161 1561
rect -115 1515 -92 1561
rect 445 1549 491 1653
rect 1261 1549 1307 1653
rect 2077 1549 2123 1653
rect 2893 1549 2939 1653
rect 3709 1549 3755 1653
rect 4296 1578 4385 1598
rect -181 530 -92 1515
rect 4296 1532 4317 1578
rect 4363 1532 4385 1578
rect 224 1479 297 1492
rect 224 1427 234 1479
rect 286 1427 297 1479
rect 224 1413 297 1427
rect 634 1478 707 1491
rect 634 1426 644 1478
rect 696 1426 707 1478
rect 634 1412 707 1426
rect 1043 1477 1116 1490
rect 1043 1425 1053 1477
rect 1105 1425 1116 1477
rect 1043 1411 1116 1425
rect 1452 1476 1525 1489
rect 1452 1424 1462 1476
rect 1514 1424 1525 1476
rect 1452 1410 1525 1424
rect 1861 1476 1934 1489
rect 1861 1424 1871 1476
rect 1923 1424 1934 1476
rect 1861 1410 1934 1424
rect 2267 1476 2340 1489
rect 2267 1424 2277 1476
rect 2329 1424 2340 1476
rect 2267 1410 2340 1424
rect 2674 1476 2747 1489
rect 2674 1424 2684 1476
rect 2736 1424 2747 1476
rect 2674 1410 2747 1424
rect 3082 1475 3155 1488
rect 3082 1423 3092 1475
rect 3144 1423 3155 1475
rect 3082 1409 3155 1423
rect 3490 1477 3563 1490
rect 3490 1425 3500 1477
rect 3552 1425 3563 1477
rect 3490 1411 3563 1425
rect 3898 1476 3971 1489
rect 3898 1424 3908 1476
rect 3960 1424 3971 1476
rect 3898 1410 3971 1424
rect 37 1142 83 1353
rect 853 1142 899 1353
rect 1341 1287 1431 1307
rect 1341 1235 1359 1287
rect 1411 1235 1431 1287
rect 1341 1217 1431 1235
rect 1669 1142 1715 1353
rect 2157 1288 2247 1307
rect 2157 1236 2175 1288
rect 2227 1236 2247 1288
rect 2157 1217 2247 1236
rect 2485 1142 2531 1353
rect 2769 1287 2859 1307
rect 2769 1235 2786 1287
rect 2838 1235 2859 1287
rect 2769 1217 2859 1235
rect 3301 1142 3347 1353
rect 4117 1142 4163 1353
rect 0 1105 4200 1142
rect 0 1053 35 1105
rect 87 1093 4200 1105
rect 0 1047 41 1053
rect 87 1047 251 1093
rect 297 1047 461 1093
rect 507 1047 671 1093
rect 717 1047 881 1093
rect 927 1047 1091 1093
rect 1137 1047 1301 1093
rect 1347 1047 1511 1093
rect 1557 1047 1721 1093
rect 1767 1047 1931 1093
rect 1977 1047 2141 1093
rect 2187 1047 2351 1093
rect 2397 1047 2561 1093
rect 2607 1047 2771 1093
rect 2817 1047 2981 1093
rect 3027 1047 3191 1093
rect 3237 1047 3401 1093
rect 3447 1047 3611 1093
rect 3657 1047 3821 1093
rect 3867 1047 4023 1093
rect 4077 1047 4200 1093
rect 0 1041 4023 1047
rect 4075 1041 4200 1047
rect 0 996 4200 1041
rect 117 908 207 924
rect 117 880 137 908
rect 37 856 137 880
rect 189 856 207 908
rect 37 834 207 856
rect 37 785 83 834
rect 445 785 491 996
rect 729 901 819 923
rect 729 855 751 901
rect 797 880 819 901
rect 933 902 1023 924
rect 933 880 955 902
rect 797 856 955 880
rect 1001 856 1023 902
rect 797 855 1023 856
rect 729 834 1023 855
rect 729 833 933 834
rect 853 785 899 833
rect 1261 785 1307 996
rect 1545 904 1635 924
rect 1545 852 1562 904
rect 1614 881 1635 904
rect 1749 902 1839 924
rect 1749 881 1771 902
rect 1614 856 1771 881
rect 1817 856 1839 902
rect 1614 852 1839 856
rect 1545 834 1839 852
rect 1669 785 1715 834
rect 2077 785 2123 996
rect 2361 906 2451 924
rect 2361 854 2380 906
rect 2432 881 2451 906
rect 2565 902 2655 924
rect 2565 881 2587 902
rect 2432 856 2587 881
rect 2633 856 2655 902
rect 2432 854 2655 856
rect 2361 834 2655 854
rect 2485 785 2531 834
rect 2893 785 2939 996
rect 3177 902 3267 924
rect 3177 856 3199 902
rect 3245 881 3267 902
rect 3381 902 3471 924
rect 3381 881 3403 902
rect 3245 856 3403 881
rect 3449 856 3471 902
rect 3177 834 3471 856
rect 3301 785 3347 834
rect 3709 785 3755 996
rect 3993 902 4083 924
rect 3993 856 4015 902
rect 4061 880 4083 902
rect 4061 856 4163 880
rect 3993 834 4163 856
rect 4117 785 4163 834
rect 241 548 287 589
rect 241 540 359 548
rect 649 547 695 589
rect 601 540 695 547
rect 241 530 411 540
rect 525 530 695 540
rect 1057 543 1103 594
rect 1465 554 1511 597
rect 1057 540 1169 543
rect 1405 540 1511 554
rect 1057 530 1227 540
rect 1341 530 1511 540
rect 1873 543 1919 599
rect 2281 560 2327 596
rect 1873 540 1974 543
rect 2224 540 2327 560
rect 1873 530 2043 540
rect 2157 530 2327 540
rect 2689 556 2735 598
rect 3097 564 3143 596
rect 2689 540 2785 556
rect 3031 540 3143 564
rect 2689 530 2859 540
rect 2973 530 3143 540
rect 3505 567 3551 600
rect 3505 540 3625 567
rect 3913 566 3959 600
rect 3858 540 3959 566
rect 3505 530 3675 540
rect 3789 530 3959 540
rect 4296 530 4385 1532
rect -181 518 4385 530
rect -181 472 343 518
rect 389 472 547 518
rect 593 472 1159 518
rect 1205 472 1363 518
rect 1409 472 1975 518
rect 2021 472 2179 518
rect 2225 472 2791 518
rect 2837 472 2995 518
rect 3041 472 3607 518
rect 3653 472 3811 518
rect 3857 472 4385 518
rect -181 454 4385 472
rect -181 441 751 454
rect 241 430 358 441
rect 241 337 287 430
rect 649 408 751 441
rect 797 441 955 454
rect 797 408 819 441
rect 649 386 819 408
rect 933 408 955 441
rect 1001 441 1567 454
rect 1001 408 1103 441
rect 933 386 1103 408
rect 649 337 695 386
rect 987 379 1103 386
rect 1057 337 1103 379
rect 1465 408 1567 441
rect 1613 441 1771 454
rect 1613 408 1635 441
rect 1465 386 1635 408
rect 1749 408 1771 441
rect 1817 441 2383 454
rect 1817 408 1919 441
rect 1749 386 1919 408
rect 1465 383 1610 386
rect 1465 337 1511 383
rect 1781 377 1919 386
rect 1873 337 1919 377
rect 2281 408 2383 441
rect 2429 441 2587 454
rect 2429 408 2451 441
rect 2281 386 2451 408
rect 2565 408 2587 441
rect 2633 441 3199 454
rect 2633 408 2735 441
rect 2565 386 2735 408
rect 2281 367 2389 386
rect 2622 372 2735 386
rect 2281 337 2327 367
rect 2689 337 2735 372
rect 3097 408 3199 441
rect 3245 441 3403 454
rect 3245 408 3267 441
rect 3097 386 3267 408
rect 3381 408 3403 441
rect 3449 441 4385 454
rect 3449 408 3551 441
rect 3381 386 3551 408
rect 3097 378 3229 386
rect 3097 337 3143 378
rect 3439 368 3551 386
rect 3505 337 3551 368
rect 3913 337 3959 441
rect -186 165 -87 196
rect -186 113 -161 165
rect -109 113 -87 165
rect -186 76 -87 113
rect 37 -63 83 141
rect 445 95 491 141
rect 321 73 615 95
rect 321 27 343 73
rect 389 48 547 73
rect 389 27 411 48
rect 321 5 411 27
rect 525 27 547 48
rect 593 27 615 73
rect 525 5 615 27
rect 853 -63 899 141
rect 1261 95 1307 141
rect 1137 75 1431 95
rect 1137 23 1154 75
rect 1206 73 1431 75
rect 1206 48 1363 73
rect 1206 23 1227 48
rect 1137 5 1227 23
rect 1341 27 1363 48
rect 1409 27 1431 73
rect 1341 5 1431 27
rect 1669 -63 1715 141
rect 2077 95 2123 141
rect 1953 76 2247 95
rect 1953 24 1975 76
rect 2027 73 2247 76
rect 2027 48 2179 73
rect 2027 24 2043 48
rect 1953 5 2043 24
rect 2157 27 2179 48
rect 2225 27 2247 73
rect 2157 5 2247 27
rect 2485 -63 2531 141
rect 2893 95 2939 141
rect 2769 76 3063 95
rect 2769 24 2787 76
rect 2839 73 3063 76
rect 2839 48 2995 73
rect 2839 24 2859 48
rect 2769 5 2859 24
rect 2973 27 2995 48
rect 3041 27 3063 73
rect 2973 5 3063 27
rect 3301 -63 3347 141
rect 3709 95 3755 141
rect 3585 73 3879 95
rect 3585 27 3607 73
rect 3653 48 3811 73
rect 3653 27 3675 48
rect 3585 5 3675 27
rect 3789 27 3811 48
rect 3857 27 3879 73
rect 3789 5 3879 27
rect 4117 -63 4163 141
rect 0 -110 4200 -63
rect 0 -162 35 -110
rect 87 -112 4200 -110
rect 87 -158 251 -112
rect 297 -158 461 -112
rect 507 -158 671 -112
rect 717 -158 881 -112
rect 927 -158 1091 -112
rect 1137 -158 1301 -112
rect 1347 -158 1511 -112
rect 1557 -158 1721 -112
rect 1767 -158 1931 -112
rect 1977 -158 2141 -112
rect 2187 -158 2351 -112
rect 2397 -158 2561 -112
rect 2607 -158 2771 -112
rect 2817 -158 2981 -112
rect 3027 -158 3191 -112
rect 3237 -158 3401 -112
rect 3447 -158 3611 -112
rect 3657 -158 3821 -112
rect 3867 -113 4031 -112
rect 4077 -113 4200 -112
rect 3867 -158 4026 -113
rect 87 -162 4026 -158
rect 0 -165 4026 -162
rect 4078 -165 4200 -113
rect 0 -209 4200 -165
<< via1 >>
rect -224 6793 -172 6796
rect -224 6747 -221 6793
rect -221 6747 -175 6793
rect -175 6747 -172 6793
rect -224 6744 -172 6747
rect -1513 6574 -1461 6626
rect -1102 6573 -1050 6625
rect -694 6573 -642 6625
rect -288 6573 -236 6625
rect -1513 6106 -1461 6158
rect -1102 6092 -1050 6144
rect -697 6092 -645 6144
rect -288 6102 -236 6154
rect -1428 5982 -1376 5985
rect -1428 5936 -1382 5982
rect -1382 5936 -1376 5982
rect -1428 5933 -1376 5936
rect -177 6012 -125 6017
rect -177 5966 -134 6012
rect -134 5966 -125 6012
rect -177 5965 -125 5966
rect 599 6061 651 6064
rect 599 6015 603 6061
rect 603 6015 649 6061
rect 649 6015 651 6061
rect 599 6012 651 6015
rect 1778 5703 1785 5749
rect 1785 5703 1830 5749
rect 1778 5697 1830 5703
rect 2397 5703 2443 5749
rect 2443 5703 2449 5749
rect 2397 5697 2449 5703
rect 395 5516 447 5528
rect 395 5476 401 5516
rect 401 5476 447 5516
rect 3754 5470 3761 5510
rect 3761 5470 3806 5510
rect 3754 5458 3806 5470
rect 1105 5333 1157 5334
rect 1105 5287 1111 5333
rect 1111 5287 1157 5333
rect 1105 5282 1157 5287
rect -1551 5124 -1499 5176
rect -1144 5123 -1092 5175
rect -737 5123 -685 5175
rect -329 5123 -277 5175
rect 2366 5145 2418 5197
rect 2774 5141 2826 5193
rect 3181 5142 3233 5194
rect 2165 4971 2217 5023
rect 3591 5142 3643 5194
rect -1552 4778 -1500 4830
rect -1144 4778 -1092 4830
rect -737 4778 -685 4830
rect -329 4778 -277 4830
rect 697 4650 703 4696
rect 703 4650 749 4696
rect 697 4644 749 4650
rect 2367 4796 2419 4848
rect 2772 4794 2824 4846
rect 3182 4794 3234 4846
rect 3591 4796 3643 4848
rect -127 4512 -75 4514
rect -127 4466 -126 4512
rect -126 4466 -80 4512
rect -80 4466 -75 4512
rect -127 4462 -75 4466
rect 395 4497 447 4499
rect 395 4451 401 4497
rect 401 4451 447 4497
rect 3754 4451 3761 4497
rect 3761 4451 3806 4497
rect 395 4447 447 4451
rect 3754 4445 3806 4451
rect 133 4332 185 4333
rect 133 4286 139 4332
rect 139 4286 185 4332
rect 133 4281 185 4286
rect 450 4266 502 4318
rect 4011 4332 4063 4335
rect 4011 4286 4015 4332
rect 4015 4286 4061 4332
rect 4061 4286 4063 4332
rect 4011 4283 4063 4286
rect 238 4144 290 4196
rect 646 4144 698 4196
rect 1053 4144 1105 4196
rect 1463 4144 1515 4196
rect 1869 4144 1921 4196
rect 2275 4144 2327 4196
rect 2685 4144 2737 4196
rect 3090 4144 3142 4196
rect 3502 4144 3554 4196
rect 3909 4144 3961 4196
rect 1154 4051 1206 4054
rect 1154 4005 1159 4051
rect 1159 4005 1205 4051
rect 1205 4005 1206 4051
rect 1154 4002 1206 4005
rect 2786 4051 2838 4053
rect 2786 4005 2791 4051
rect 2791 4005 2837 4051
rect 2837 4005 2838 4051
rect 2786 4001 2838 4005
rect 6 3775 58 3827
rect 4151 3775 4203 3827
rect 187 3637 239 3639
rect 187 3591 192 3637
rect 192 3591 238 3637
rect 238 3591 239 3637
rect 187 3587 239 3591
rect 1819 3637 1871 3640
rect 1819 3591 1825 3637
rect 1825 3591 1871 3637
rect 2331 3637 2383 3641
rect 1819 3588 1871 3591
rect 2331 3591 2332 3637
rect 2332 3591 2378 3637
rect 2378 3591 2383 3637
rect 2331 3589 2383 3591
rect 3955 3637 4007 3639
rect 3955 3591 3959 3637
rect 3959 3591 4005 3637
rect 4005 3591 4007 3637
rect 3955 3587 4007 3591
rect 1258 3181 1310 3183
rect 2886 3182 2938 3184
rect 1258 3135 1262 3181
rect 1262 3135 1308 3181
rect 1308 3135 1310 3181
rect 1258 3131 1310 3135
rect 2886 3136 2891 3182
rect 2891 3136 2937 3182
rect 2937 3136 2938 3182
rect 2886 3132 2938 3136
rect 1090 2727 1142 2734
rect 1090 2682 1103 2727
rect 1103 2682 1142 2727
rect 1917 2727 1969 2730
rect 1917 2681 1924 2727
rect 1924 2681 1969 2727
rect 1917 2678 1969 2681
rect 2738 2727 2790 2735
rect 2738 2683 2784 2727
rect 2784 2683 2790 2727
rect 26 2505 78 2557
rect 4155 2484 4207 2536
rect 35 2308 87 2320
rect 35 2268 41 2308
rect 41 2268 87 2308
rect 4023 2262 4031 2308
rect 4031 2262 4075 2308
rect 4023 2256 4075 2262
rect 1765 2117 1817 2118
rect 1765 2071 1771 2117
rect 1771 2071 1817 2117
rect 1765 2066 1817 2071
rect 2380 2115 2432 2119
rect 2380 2069 2383 2115
rect 2383 2069 2429 2115
rect 2429 2069 2432 2115
rect 2380 2067 2432 2069
rect 230 1871 282 1923
rect 641 1879 693 1931
rect 1048 1878 1100 1930
rect 1458 1878 1510 1930
rect 1864 1878 1916 1930
rect 2274 1878 2326 1930
rect 2681 1878 2733 1930
rect 3086 1878 3138 1930
rect 3496 1878 3548 1930
rect 3907 1882 3959 1934
rect 234 1427 286 1479
rect 644 1426 696 1478
rect 1053 1425 1105 1477
rect 1462 1424 1514 1476
rect 1871 1424 1923 1476
rect 2277 1424 2329 1476
rect 2684 1424 2736 1476
rect 3092 1423 3144 1475
rect 3500 1425 3552 1477
rect 3908 1424 3960 1476
rect 1359 1285 1411 1287
rect 1359 1239 1363 1285
rect 1363 1239 1409 1285
rect 1409 1239 1411 1285
rect 1359 1235 1411 1239
rect 2175 1285 2227 1288
rect 2175 1239 2179 1285
rect 2179 1239 2225 1285
rect 2225 1239 2227 1285
rect 2175 1236 2227 1239
rect 2786 1285 2838 1287
rect 2786 1239 2791 1285
rect 2791 1239 2837 1285
rect 2837 1239 2838 1285
rect 2786 1235 2838 1239
rect 35 1093 87 1105
rect 35 1053 41 1093
rect 41 1053 87 1093
rect 4023 1047 4031 1093
rect 4031 1047 4075 1093
rect 4023 1041 4075 1047
rect 137 902 189 908
rect 137 856 139 902
rect 139 856 185 902
rect 185 856 189 902
rect 1562 902 1614 904
rect 1562 856 1567 902
rect 1567 856 1613 902
rect 1613 856 1614 902
rect 1562 852 1614 856
rect 2380 902 2432 906
rect 2380 856 2383 902
rect 2383 856 2429 902
rect 2429 856 2432 902
rect 2380 854 2432 856
rect -161 113 -109 165
rect 1154 73 1206 75
rect 1154 27 1159 73
rect 1159 27 1205 73
rect 1205 27 1206 73
rect 1154 23 1206 27
rect 1975 73 2027 76
rect 1975 27 2021 73
rect 2021 27 2027 73
rect 1975 24 2027 27
rect 2787 73 2839 76
rect 2787 27 2791 73
rect 2791 27 2837 73
rect 2837 27 2839 73
rect 2787 24 2839 27
rect 35 -112 87 -110
rect 35 -158 41 -112
rect 41 -158 87 -112
rect 4026 -158 4031 -113
rect 4031 -158 4077 -113
rect 4077 -158 4078 -113
rect 35 -162 87 -158
rect 4026 -165 4078 -158
<< metal2 >>
rect -1705 6796 657 6815
rect -1705 6748 -224 6796
rect -1705 5978 -1638 6748
rect -235 6744 -224 6748
rect -172 6748 657 6796
rect -172 6744 -167 6748
rect -235 6732 -167 6744
rect -1527 6626 -1450 6637
rect -1527 6574 -1513 6626
rect -1461 6616 -1450 6626
rect -1116 6625 -1039 6636
rect -1116 6616 -1102 6625
rect -1461 6574 -1102 6616
rect -1527 6573 -1102 6574
rect -1050 6616 -1039 6625
rect -708 6625 -631 6636
rect -708 6616 -694 6625
rect -1050 6573 -694 6616
rect -642 6616 -631 6625
rect -302 6625 -225 6636
rect -302 6616 -288 6625
rect -642 6573 -288 6616
rect -236 6573 -225 6625
rect -1527 6560 -225 6573
rect -1516 6559 -225 6560
rect -1516 6205 -1459 6559
rect -1099 6205 -1042 6559
rect -694 6205 -637 6559
rect -287 6205 -230 6559
rect -1516 6169 -230 6205
rect -1527 6165 -230 6169
rect -1527 6158 -225 6165
rect -1527 6106 -1513 6158
rect -1461 6154 -225 6158
rect -1461 6148 -288 6154
rect -1461 6106 -1450 6148
rect -1527 6092 -1450 6106
rect -1116 6144 -1039 6148
rect -1116 6092 -1102 6144
rect -1050 6092 -1039 6144
rect -1116 6078 -1039 6092
rect -711 6144 -634 6148
rect -711 6092 -697 6144
rect -645 6092 -634 6144
rect -711 6078 -634 6092
rect -302 6102 -288 6148
rect -236 6102 -225 6154
rect -302 6088 -225 6102
rect 590 6085 657 6748
rect 579 6064 674 6085
rect -130 6033 -74 6034
rect -188 6017 -74 6033
rect -1441 5985 -1368 6004
rect -1441 5978 -1428 5985
rect -1705 5933 -1428 5978
rect -1376 5933 -1368 5985
rect -188 5965 -177 6017
rect -125 5965 -74 6017
rect 579 6012 599 6064
rect 651 6012 674 6064
rect 579 5992 674 6012
rect -188 5938 -74 5965
rect -1705 5914 -1368 5933
rect -1705 5911 -1394 5914
rect -130 5751 -74 5938
rect 1763 5751 1853 5771
rect 2375 5751 2465 5771
rect -130 5749 2465 5751
rect -130 5697 1778 5749
rect 1830 5697 2397 5749
rect 2449 5697 2465 5749
rect -130 5695 2465 5697
rect 1763 5681 1853 5695
rect 384 5528 461 5540
rect 384 5476 395 5528
rect 447 5476 461 5528
rect 384 5464 461 5476
rect -1565 5178 -1488 5187
rect -1158 5178 -1081 5186
rect -751 5178 -674 5186
rect -343 5178 -266 5186
rect -1565 5176 -266 5178
rect -1565 5124 -1551 5176
rect -1499 5175 -266 5176
rect -1499 5124 -1144 5175
rect -1565 5123 -1144 5124
rect -1092 5123 -737 5175
rect -685 5123 -329 5175
rect -277 5123 -266 5175
rect -1565 5120 -266 5123
rect -1565 5110 -1488 5120
rect -1555 4841 -1497 5110
rect -1158 5109 -1081 5120
rect -751 5109 -674 5120
rect -343 5109 -266 5120
rect -1146 4841 -1088 5109
rect -736 4841 -678 5109
rect -333 4841 -275 5109
rect -1566 4830 -1489 4841
rect -1566 4778 -1552 4830
rect -1500 4825 -1489 4830
rect -1158 4830 -1081 4841
rect -1158 4825 -1144 4830
rect -1500 4778 -1144 4825
rect -1092 4825 -1081 4830
rect -751 4830 -674 4841
rect -751 4825 -737 4830
rect -1092 4778 -737 4825
rect -685 4825 -674 4830
rect -343 4830 -266 4841
rect -343 4825 -329 4830
rect -685 4778 -329 4825
rect -277 4778 -266 4830
rect -1566 4767 -266 4778
rect -1566 4764 -1489 4767
rect -1158 4764 -1081 4767
rect -751 4764 -674 4767
rect -343 4764 -266 4767
rect -128 4526 -72 4561
rect -140 4521 -63 4526
rect -140 4514 -39 4521
rect -140 4499 -127 4514
rect -182 4462 -127 4499
rect -75 4499 -39 4514
rect 393 4511 449 5464
rect 1089 5334 1179 5355
rect 1089 5332 1105 5334
rect 690 5282 1105 5332
rect 1157 5282 1179 5334
rect 690 5276 1179 5282
rect 690 4723 746 5276
rect 1089 5265 1179 5276
rect 2163 5043 2219 5695
rect 2375 5681 2465 5695
rect 3743 5510 3818 5523
rect 3743 5458 3754 5510
rect 3806 5458 3818 5510
rect 3743 5444 3818 5458
rect 2355 5198 2430 5210
rect 2763 5198 2838 5206
rect 3170 5198 3245 5207
rect 3580 5198 3655 5207
rect 2355 5197 3655 5198
rect 2355 5145 2366 5197
rect 2418 5194 3655 5197
rect 2418 5193 3181 5194
rect 2418 5145 2774 5193
rect 2355 5142 2774 5145
rect 2355 5131 2430 5142
rect 2763 5141 2774 5142
rect 2826 5142 3181 5193
rect 3233 5142 3591 5194
rect 3643 5142 3655 5194
rect 2826 5141 2838 5142
rect 2146 5023 2236 5043
rect 2146 4971 2165 5023
rect 2217 4971 2236 5023
rect 2146 4953 2236 4971
rect 2370 4861 2426 5131
rect 2763 5127 2838 5141
rect 3170 5128 3245 5142
rect 3580 5128 3655 5142
rect 2356 4848 2431 4861
rect 2772 4859 2828 5127
rect 3178 4859 3234 5128
rect 3585 4861 3641 5128
rect 2356 4796 2367 4848
rect 2419 4796 2431 4848
rect 2356 4782 2431 4796
rect 2761 4846 2836 4859
rect 2761 4794 2772 4846
rect 2824 4794 2836 4846
rect 2761 4780 2836 4794
rect 3171 4846 3246 4859
rect 3171 4794 3182 4846
rect 3234 4794 3246 4846
rect 3171 4780 3246 4794
rect 3580 4848 3655 4861
rect 3580 4796 3591 4848
rect 3643 4796 3655 4848
rect 3580 4782 3655 4796
rect 678 4722 746 4723
rect 678 4696 771 4722
rect 678 4644 697 4696
rect 749 4644 771 4696
rect 678 4626 771 4644
rect 687 4625 771 4626
rect 384 4506 461 4511
rect 256 4499 461 4506
rect -75 4462 395 4499
rect -182 4447 395 4462
rect 447 4447 461 4499
rect -182 4435 461 4447
rect -182 4434 446 4435
rect -182 4427 418 4434
rect -182 2329 -110 4427
rect 117 4348 206 4355
rect 92 4333 206 4348
rect 690 4333 746 4625
rect 3757 4510 3813 5444
rect 3743 4502 3818 4510
rect 3743 4497 4484 4502
rect 3743 4445 3754 4497
rect 3806 4445 4484 4497
rect 3743 4431 4484 4445
rect 3766 4430 4484 4431
rect 92 4281 133 4333
rect 185 4281 206 4333
rect 92 4264 206 4281
rect 431 4318 746 4333
rect 431 4266 450 4318
rect 502 4277 746 4318
rect 3993 4346 4083 4354
rect 3993 4335 4115 4346
rect 3993 4283 4011 4335
rect 4063 4283 4115 4335
rect 502 4266 516 4277
rect 92 4021 148 4264
rect 431 4249 516 4266
rect 3993 4264 4115 4283
rect 228 4196 301 4209
rect 228 4144 238 4196
rect 290 4193 301 4196
rect 636 4196 709 4209
rect 636 4193 646 4196
rect 290 4144 646 4193
rect 698 4193 709 4196
rect 1043 4196 1116 4209
rect 1043 4193 1053 4196
rect 698 4144 1053 4193
rect 1105 4193 1116 4196
rect 1453 4196 1526 4209
rect 1453 4193 1463 4196
rect 1105 4144 1463 4193
rect 1515 4193 1526 4196
rect 1859 4196 1932 4209
rect 1859 4193 1869 4196
rect 1515 4144 1869 4193
rect 1921 4193 1932 4196
rect 2265 4196 2338 4209
rect 2265 4193 2275 4196
rect 1921 4144 2275 4193
rect 2327 4193 2338 4196
rect 2675 4196 2748 4209
rect 2675 4193 2685 4196
rect 2327 4144 2685 4193
rect 2737 4193 2748 4196
rect 3080 4196 3153 4209
rect 3080 4193 3090 4196
rect 2737 4144 3090 4193
rect 3142 4193 3153 4196
rect 3492 4196 3565 4209
rect 3492 4193 3502 4196
rect 3142 4144 3502 4193
rect 3554 4193 3565 4196
rect 3899 4196 3972 4209
rect 3899 4193 3909 4196
rect 3554 4144 3909 4193
rect 3961 4144 3972 4196
rect 228 4137 3972 4144
rect 228 4130 301 4137
rect 636 4130 709 4137
rect 1043 4130 1116 4137
rect 1453 4130 1526 4137
rect 1859 4130 1932 4137
rect 2265 4130 2338 4137
rect 2675 4130 2748 4137
rect 3080 4130 3153 4137
rect 3492 4130 3565 4137
rect 3899 4130 3972 4137
rect 1137 4054 1227 4073
rect 92 3965 246 4021
rect 1137 4002 1154 4054
rect 1206 4033 1227 4054
rect 2769 4053 2859 4073
rect 1206 4002 1309 4033
rect 1137 3983 1309 4002
rect 2769 4001 2786 4053
rect 2838 4035 2859 4053
rect 2838 4001 2946 4035
rect 4059 4021 4115 4264
rect 2769 3983 2946 4001
rect 1153 3977 1309 3983
rect 2810 3979 2946 3983
rect -4 3832 69 3840
rect -4 3827 79 3832
rect -4 3775 6 3827
rect 58 3775 79 3827
rect -4 3761 79 3775
rect 23 2570 79 3761
rect 190 3658 246 3965
rect 171 3639 259 3658
rect 171 3587 187 3639
rect 239 3587 259 3639
rect 171 3570 259 3587
rect 1253 3210 1309 3977
rect 1809 3646 1882 3653
rect 2321 3646 2394 3654
rect 1809 3641 2394 3646
rect 1809 3640 2331 3641
rect 1809 3588 1819 3640
rect 1871 3590 2331 3640
rect 1871 3588 1882 3590
rect 1809 3574 1882 3588
rect 2310 3589 2331 3590
rect 2383 3589 2394 3641
rect 2310 3575 2394 3589
rect 1231 3183 1337 3210
rect 1231 3131 1258 3183
rect 1310 3131 1337 3183
rect 1231 3108 1337 3131
rect 1080 2734 1153 2747
rect 1080 2682 1090 2734
rect 1142 2723 1153 2734
rect 1814 2743 1870 3574
rect 1814 2730 1980 2743
rect 1814 2723 1917 2730
rect 1142 2682 1917 2723
rect 1080 2678 1917 2682
rect 1969 2723 1980 2730
rect 2310 2723 2366 3575
rect 2890 3208 2946 3979
rect 3956 3965 4115 4021
rect 3956 3658 4012 3965
rect 4141 3827 4214 3840
rect 4141 3775 4151 3827
rect 4203 3775 4214 3827
rect 4141 3761 4214 3775
rect 3938 3639 4026 3658
rect 3938 3587 3955 3639
rect 4007 3587 4026 3639
rect 3938 3570 4026 3587
rect 2863 3184 2964 3208
rect 2863 3132 2886 3184
rect 2938 3132 2964 3184
rect 2863 3111 2964 3132
rect 2728 2735 2801 2748
rect 2728 2723 2738 2735
rect 1969 2683 2738 2723
rect 2790 2683 2801 2735
rect 1969 2678 2801 2683
rect 1080 2669 2801 2678
rect 1080 2668 2772 2669
rect 1123 2667 2772 2668
rect 1907 2664 1980 2667
rect 16 2557 89 2570
rect 16 2505 26 2557
rect 78 2505 89 2557
rect 4151 2549 4207 3761
rect 16 2491 89 2505
rect 4145 2536 4218 2549
rect 4145 2484 4155 2536
rect 4207 2484 4218 2536
rect 4145 2470 4218 2484
rect 24 2329 101 2332
rect -182 2320 101 2329
rect -182 2268 35 2320
rect 87 2268 101 2320
rect -182 2257 101 2268
rect 24 2256 101 2257
rect 4012 2316 4089 2320
rect 4412 2316 4484 4430
rect 4012 2308 4484 2316
rect 4012 2256 4023 2308
rect 4075 2256 4484 2308
rect 33 1117 89 2256
rect 4012 2244 4484 2256
rect 1749 2122 1839 2139
rect 1749 2118 1766 2122
rect 1749 2066 1765 2118
rect 1822 2066 1839 2122
rect 1749 2049 1839 2066
rect 2361 2120 2451 2137
rect 2361 2064 2378 2120
rect 2434 2064 2451 2120
rect 2361 2047 2451 2064
rect 220 1923 293 1936
rect 220 1871 230 1923
rect 282 1919 293 1923
rect 631 1931 704 1944
rect 631 1919 641 1931
rect 282 1879 641 1919
rect 693 1919 704 1931
rect 1038 1930 1111 1943
rect 1038 1919 1048 1930
rect 693 1879 1048 1919
rect 282 1878 1048 1879
rect 1100 1919 1111 1930
rect 1448 1930 1521 1943
rect 1448 1919 1458 1930
rect 1100 1878 1458 1919
rect 1510 1919 1521 1930
rect 1854 1930 1927 1943
rect 1854 1919 1864 1930
rect 1510 1878 1864 1919
rect 1916 1919 1927 1930
rect 2264 1930 2337 1943
rect 2264 1919 2274 1930
rect 1916 1878 2274 1919
rect 2326 1919 2337 1930
rect 2671 1930 2744 1943
rect 2671 1919 2681 1930
rect 2326 1878 2681 1919
rect 2733 1919 2744 1930
rect 3076 1930 3149 1943
rect 3076 1919 3086 1930
rect 2733 1878 3086 1919
rect 3138 1919 3149 1930
rect 3486 1930 3559 1943
rect 3486 1919 3496 1930
rect 3138 1878 3496 1919
rect 3548 1919 3559 1930
rect 3897 1934 3970 1947
rect 3897 1919 3907 1934
rect 3548 1882 3907 1919
rect 3959 1882 3970 1934
rect 3548 1878 3970 1882
rect 282 1871 3970 1878
rect 220 1868 3970 1871
rect 220 1863 3966 1868
rect 220 1857 293 1863
rect 229 1492 285 1857
rect 224 1479 297 1492
rect 638 1491 694 1863
rect 224 1427 234 1479
rect 286 1427 297 1479
rect 224 1413 297 1427
rect 634 1478 707 1491
rect 1047 1490 1103 1863
rect 634 1426 644 1478
rect 696 1426 707 1478
rect 634 1412 707 1426
rect 1043 1477 1116 1490
rect 1458 1489 1514 1863
rect 1865 1489 1921 1863
rect 2280 1489 2336 1863
rect 2677 1489 2733 1863
rect 1043 1425 1053 1477
rect 1105 1425 1116 1477
rect 1043 1411 1116 1425
rect 1452 1476 1525 1489
rect 1452 1424 1462 1476
rect 1514 1424 1525 1476
rect 1452 1410 1525 1424
rect 1861 1476 1934 1489
rect 1861 1424 1871 1476
rect 1923 1424 1934 1476
rect 1861 1410 1934 1424
rect 2267 1476 2340 1489
rect 2267 1424 2277 1476
rect 2329 1424 2340 1476
rect 2267 1410 2340 1424
rect 2674 1476 2747 1489
rect 3088 1488 3144 1863
rect 3504 1490 3560 1863
rect 2674 1424 2684 1476
rect 2736 1424 2747 1476
rect 2674 1410 2747 1424
rect 3082 1475 3155 1488
rect 3082 1423 3092 1475
rect 3144 1423 3155 1475
rect 3082 1409 3155 1423
rect 3490 1477 3563 1490
rect 3910 1489 3966 1863
rect 3490 1425 3500 1477
rect 3552 1425 3563 1477
rect 3490 1411 3563 1425
rect 3898 1476 3971 1489
rect 3898 1424 3908 1476
rect 3960 1424 3971 1476
rect 3898 1410 3971 1424
rect 1341 1290 1431 1307
rect 2157 1290 2246 1307
rect 2769 1290 2859 1307
rect 1341 1289 2173 1290
rect 1341 1233 1357 1289
rect 1413 1234 2173 1289
rect 2229 1289 2859 1290
rect 2229 1234 2784 1289
rect 1413 1233 1431 1234
rect 1341 1217 1431 1233
rect 2157 1217 2263 1234
rect 2769 1233 2784 1234
rect 2840 1233 2859 1289
rect 2769 1217 2859 1233
rect 24 1105 101 1117
rect 24 1053 35 1105
rect 87 1084 101 1105
rect 87 1053 808 1084
rect 24 1041 808 1053
rect 27 1028 808 1041
rect 127 908 200 919
rect 127 856 137 908
rect 189 856 200 908
rect -186 176 -87 196
rect 127 176 200 856
rect -186 165 200 176
rect -186 113 -161 165
rect -109 113 200 165
rect -186 103 200 113
rect -186 76 -87 103
rect 24 -110 101 -98
rect 24 -162 35 -110
rect 87 -112 101 -110
rect 752 -112 808 1028
rect 1367 904 1423 1217
rect 1548 904 1630 921
rect 2207 904 2263 1217
rect 2366 906 2447 920
rect 2366 904 2380 906
rect 1367 852 1562 904
rect 1614 854 2380 904
rect 2432 904 2447 906
rect 2799 904 2855 1217
rect 4029 1105 4085 2244
rect 4012 1093 4089 1105
rect 4012 1041 4023 1093
rect 4075 1041 4089 1093
rect 4012 1029 4089 1041
rect 2432 854 2855 904
rect 1614 852 2855 854
rect 1367 848 2855 852
rect 1548 837 1630 848
rect 2363 840 2447 848
rect 1139 75 1222 91
rect 1554 75 1610 837
rect 1961 76 2044 91
rect 1961 75 1975 76
rect 1139 23 1154 75
rect 1206 24 1975 75
rect 2027 75 2044 76
rect 2363 75 2419 840
rect 2772 76 2855 92
rect 2772 75 2787 76
rect 2027 24 2787 75
rect 2839 24 2855 76
rect 1206 23 2855 24
rect 1139 19 2855 23
rect 1139 8 1222 19
rect 1961 8 2044 19
rect 2772 8 2855 19
rect 4029 -101 4085 1029
rect 87 -162 808 -112
rect 24 -168 808 -162
rect 4015 -113 4092 -101
rect 4015 -165 4026 -113
rect 4078 -165 4092 -113
rect 24 -174 101 -168
rect 4015 -177 4092 -165
<< via2 >>
rect 1766 2118 1822 2122
rect 1766 2066 1817 2118
rect 1817 2066 1822 2118
rect 2378 2119 2434 2120
rect 2378 2067 2380 2119
rect 2380 2067 2432 2119
rect 2432 2067 2434 2119
rect 2378 2064 2434 2067
rect 1357 1287 1413 1289
rect 1357 1235 1359 1287
rect 1359 1235 1411 1287
rect 1411 1235 1413 1287
rect 1357 1233 1413 1235
rect 2173 1288 2229 1290
rect 2173 1236 2175 1288
rect 2175 1236 2227 1288
rect 2227 1236 2229 1288
rect 2173 1234 2229 1236
rect 2784 1287 2840 1289
rect 2784 1235 2786 1287
rect 2786 1235 2838 1287
rect 2838 1235 2840 1287
rect 2784 1233 2840 1235
<< metal3 >>
rect 1749 2128 1839 2139
rect 2361 2128 2451 2137
rect 1749 2122 2451 2128
rect 1749 2066 1766 2122
rect 1822 2120 2451 2122
rect 1822 2067 2378 2120
rect 1822 2066 1839 2067
rect 1749 2049 1839 2066
rect 2361 2064 2378 2067
rect 2434 2064 2451 2120
rect 1341 1291 1431 1307
rect 1341 1290 1478 1291
rect 1769 1290 1830 2049
rect 2361 2047 2451 2064
rect 2157 1290 2247 1307
rect 2375 1290 2436 2047
rect 2769 1290 2859 1307
rect 1341 1289 2173 1290
rect 1341 1233 1357 1289
rect 1413 1234 2173 1289
rect 2229 1289 2859 1290
rect 2229 1234 2784 1289
rect 1413 1233 2784 1234
rect 2840 1233 2859 1289
rect 1341 1229 2859 1233
rect 1341 1217 1431 1229
rect 2157 1217 2247 1229
rect 2769 1217 2859 1229
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_0
timestamp 1713185578
transform 1 0 1236 0 1 5168
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_1
timestamp 1713185578
transform 1 0 3007 0 1 4815
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_2
timestamp 1713185578
transform 1 0 -914 0 1 5145
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_3
timestamp 1713185578
transform 1 0 3007 0 1 5168
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_4
timestamp 1713185578
transform 1 0 1236 0 1 4815
box -876 -128 876 128
use nmos_3p3_AJEA3B  nmos_3p3_AJEA3B_5
timestamp 1713185578
transform 1 0 -914 0 1 4799
box -876 -128 876 128
use nmos_3p3_Z2JHD6  nmos_3p3_Z2JHD6_0
timestamp 1713185578
transform 1 0 2100 0 1 1902
box -2100 -168 2100 168
use nmos_3p3_Z2JHD6  nmos_3p3_Z2JHD6_1
timestamp 1713185578
transform 1 0 2100 0 1 239
box -2100 -168 2100 168
use nmos_3p3_Z2JHD6  nmos_3p3_Z2JHD6_2
timestamp 1713185578
transform 1 0 2100 0 1 687
box -2100 -168 2100 168
use nmos_3p3_Z2JHD6  nmos_3p3_Z2JHD6_3
timestamp 1713185578
transform 1 0 2100 0 1 1451
box -2100 -168 2100 168
use pfet_03v3_TTE2U8  pfet_03v3_TTE2U8_0
timestamp 1713185578
transform 1 0 -871 0 1 6117
box -938 -190 938 190
use pfet_03v3_TTE2U8  pfet_03v3_TTE2U8_1
timestamp 1713185578
transform 1 0 -871 0 1 6597
box -938 -190 938 190
use pmos_3p3_5QR9E7  pmos_3p3_5QR9E7_0
timestamp 1713185578
transform 1 0 2100 0 1 4157
box -2162 -170 2162 170
use pmos_3p3_DVJ9E7  pmos_3p3_DVJ9E7_0
timestamp 1713185578
transform 1 0 2114 0 1 5875
box -1754 -190 1754 190
use pmos_3p3_ZBCND7  pmos_3p3_ZBCND7_0
timestamp 1713185578
transform 1 0 2100 0 1 3421
box -2162 -230 2162 230
use pmos_3p3_ZBCND7  pmos_3p3_ZBCND7_1
timestamp 1713185578
transform 1 0 2100 0 1 2896
box -2162 -230 2162 230
<< labels >>
flabel nsubdiffcont 505 6259 505 6259 0 FreeSans 750 0 0 0 VDD
flabel polycontact 160 4312 160 4312 0 FreeSans 750 0 0 0 G1_2
flabel polycontact 1175 4023 1175 4023 0 FreeSans 750 0 0 0 G1_1
flabel polycontact 361 499 361 499 0 FreeSans 750 0 0 0 G2_1
flabel metal1 s 651 5747 651 5747 0 FreeSans 750 0 0 0 G_source_up
port 1 nsew
flabel metal1 s 851 5654 851 5654 0 FreeSans 750 0 0 0 G_source_dn
port 2 nsew
flabel metal1 s 513 5478 513 5478 0 FreeSans 750 0 0 0 VSS
port 3 nsew
flabel metal1 s 314 5279 314 5279 0 FreeSans 750 0 0 0 G_sink_up
port 4 nsew
flabel metal1 s 307 5018 307 5018 0 FreeSans 750 0 0 0 G_sink_dn
port 5 nsew
flabel metal1 s 2395 5173 2395 5173 0 FreeSans 750 0 0 0 SD0_1
port 6 nsew
flabel metal1 s 263 4170 263 4170 0 FreeSans 750 0 0 0 SD1_1
port 7 nsew
flabel metal1 s 252 1901 252 1901 0 FreeSans 750 0 0 0 SD2_1
port 8 nsew
flabel metal1 s -143 138 -143 138 0 FreeSans 750 0 0 0 ITAIL
port 9 nsew
flabel metal1 s -1875 4982 -1875 4982 0 FreeSans 2500 0 0 0 ITAIL_SINK
port 10 nsew
flabel metal1 s -1963 6357 -1963 6357 0 FreeSans 2500 0 0 0 ITAIL_SRC
port 11 nsew
flabel metal1 s -260 6600 -260 6600 0 FreeSans 2500 0 0 0 A1
port 12 nsew
flabel metal1 s -303 5146 -303 5146 0 FreeSans 2500 0 0 0 A2
port 13 nsew
<< end >>
