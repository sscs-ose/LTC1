magic
tech gf180mcuC
magscale 1 10
timestamp 1695100097
<< nwell >>
rect -1544 -676 1544 676
<< nsubdiff >>
rect -1520 580 1520 652
rect -1520 -580 -1448 580
rect 1448 -580 1520 580
rect -1520 -652 1520 -580
<< polysilicon >>
rect -1360 479 -1160 492
rect -1360 433 -1347 479
rect -1173 433 -1160 479
rect -1360 390 -1160 433
rect -1360 -433 -1160 -390
rect -1360 -479 -1347 -433
rect -1173 -479 -1160 -433
rect -1360 -492 -1160 -479
rect -1080 479 -880 492
rect -1080 433 -1067 479
rect -893 433 -880 479
rect -1080 390 -880 433
rect -1080 -433 -880 -390
rect -1080 -479 -1067 -433
rect -893 -479 -880 -433
rect -1080 -492 -880 -479
rect -800 479 -600 492
rect -800 433 -787 479
rect -613 433 -600 479
rect -800 390 -600 433
rect -800 -433 -600 -390
rect -800 -479 -787 -433
rect -613 -479 -600 -433
rect -800 -492 -600 -479
rect -520 479 -320 492
rect -520 433 -507 479
rect -333 433 -320 479
rect -520 390 -320 433
rect -520 -433 -320 -390
rect -520 -479 -507 -433
rect -333 -479 -320 -433
rect -520 -492 -320 -479
rect -240 479 -40 492
rect -240 433 -227 479
rect -53 433 -40 479
rect -240 390 -40 433
rect -240 -433 -40 -390
rect -240 -479 -227 -433
rect -53 -479 -40 -433
rect -240 -492 -40 -479
rect 40 479 240 492
rect 40 433 53 479
rect 227 433 240 479
rect 40 390 240 433
rect 40 -433 240 -390
rect 40 -479 53 -433
rect 227 -479 240 -433
rect 40 -492 240 -479
rect 320 479 520 492
rect 320 433 333 479
rect 507 433 520 479
rect 320 390 520 433
rect 320 -433 520 -390
rect 320 -479 333 -433
rect 507 -479 520 -433
rect 320 -492 520 -479
rect 600 479 800 492
rect 600 433 613 479
rect 787 433 800 479
rect 600 390 800 433
rect 600 -433 800 -390
rect 600 -479 613 -433
rect 787 -479 800 -433
rect 600 -492 800 -479
rect 880 479 1080 492
rect 880 433 893 479
rect 1067 433 1080 479
rect 880 390 1080 433
rect 880 -433 1080 -390
rect 880 -479 893 -433
rect 1067 -479 1080 -433
rect 880 -492 1080 -479
rect 1160 479 1360 492
rect 1160 433 1173 479
rect 1347 433 1360 479
rect 1160 390 1360 433
rect 1160 -433 1360 -390
rect 1160 -479 1173 -433
rect 1347 -479 1360 -433
rect 1160 -492 1360 -479
<< polycontact >>
rect -1347 433 -1173 479
rect -1347 -479 -1173 -433
rect -1067 433 -893 479
rect -1067 -479 -893 -433
rect -787 433 -613 479
rect -787 -479 -613 -433
rect -507 433 -333 479
rect -507 -479 -333 -433
rect -227 433 -53 479
rect -227 -479 -53 -433
rect 53 433 227 479
rect 53 -479 227 -433
rect 333 433 507 479
rect 333 -479 507 -433
rect 613 433 787 479
rect 613 -479 787 -433
rect 893 433 1067 479
rect 893 -479 1067 -433
rect 1173 433 1347 479
rect 1173 -479 1347 -433
<< ppolyres >>
rect -1360 -390 -1160 390
rect -1080 -390 -880 390
rect -800 -390 -600 390
rect -520 -390 -320 390
rect -240 -390 -40 390
rect 40 -390 240 390
rect 320 -390 520 390
rect 600 -390 800 390
rect 880 -390 1080 390
rect 1160 -390 1360 390
<< metal1 >>
rect -1358 433 -1347 479
rect -1173 433 -1162 479
rect -1078 433 -1067 479
rect -893 433 -882 479
rect -798 433 -787 479
rect -613 433 -602 479
rect -518 433 -507 479
rect -333 433 -322 479
rect -238 433 -227 479
rect -53 433 -42 479
rect 42 433 53 479
rect 227 433 238 479
rect 322 433 333 479
rect 507 433 518 479
rect 602 433 613 479
rect 787 433 798 479
rect 882 433 893 479
rect 1067 433 1078 479
rect 1162 433 1173 479
rect 1347 433 1358 479
rect -1358 -479 -1347 -433
rect -1173 -479 -1162 -433
rect -1078 -479 -1067 -433
rect -893 -479 -882 -433
rect -798 -479 -787 -433
rect -613 -479 -602 -433
rect -518 -479 -507 -433
rect -333 -479 -322 -433
rect -238 -479 -227 -433
rect -53 -479 -42 -433
rect 42 -479 53 -433
rect 227 -479 238 -433
rect 322 -479 333 -433
rect 507 -479 518 -433
rect 602 -479 613 -433
rect 787 -479 798 -433
rect 882 -479 893 -433
rect 1067 -479 1078 -433
rect 1162 -479 1173 -433
rect 1347 -479 1358 -433
<< properties >>
string FIXED_BBOX -1484 -616 1484 616
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 3.9 m 1 nx 10 wmin 0.80 lmin 1.00 rho 315 val 1.32k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
