magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2172 -2196 2172 2196
<< pwell >>
rect -172 -196 172 196
<< nmos >>
rect -56 68 56 124
rect -56 -124 56 -68
<< ndiff >>
rect -148 124 -76 132
rect 76 124 148 132
rect -148 119 -56 124
rect -148 73 -135 119
rect -89 73 -56 119
rect -148 68 -56 73
rect 56 119 148 124
rect 56 73 89 119
rect 135 73 148 119
rect 56 68 148 73
rect -148 60 -76 68
rect 76 60 148 68
rect -148 -68 -76 -60
rect 76 -68 148 -60
rect -148 -73 -56 -68
rect -148 -119 -135 -73
rect -89 -119 -56 -73
rect -148 -124 -56 -119
rect 56 -73 148 -68
rect 56 -119 89 -73
rect 135 -119 148 -73
rect 56 -124 148 -119
rect -148 -132 -76 -124
rect 76 -132 148 -124
<< ndiffc >>
rect -135 73 -89 119
rect 89 73 135 119
rect -135 -119 -89 -73
rect 89 -119 135 -73
<< polysilicon >>
rect -56 124 56 168
rect -56 24 56 68
rect -56 -68 56 -24
rect -56 -168 56 -124
<< metal1 >>
rect -146 73 -135 119
rect -89 73 -78 119
rect 78 73 89 119
rect 135 73 146 119
rect -146 -119 -135 -73
rect -89 -119 -78 -73
rect 78 -119 89 -73
rect 135 -119 146 -73
<< end >>
