magic
tech gf180mcuC
magscale 1 10
timestamp 1694586619
<< nwell >>
rect -1264 -386 1264 386
<< nsubdiff >>
rect -1240 290 1240 362
rect -1240 -290 -1168 290
rect 1168 -290 1240 290
rect -1240 -362 1240 -290
<< polysilicon >>
rect -1080 189 -880 202
rect -1080 143 -1067 189
rect -893 143 -880 189
rect -1080 100 -880 143
rect -1080 -143 -880 -100
rect -1080 -189 -1067 -143
rect -893 -189 -880 -143
rect -1080 -202 -880 -189
rect -800 189 -600 202
rect -800 143 -787 189
rect -613 143 -600 189
rect -800 100 -600 143
rect -800 -143 -600 -100
rect -800 -189 -787 -143
rect -613 -189 -600 -143
rect -800 -202 -600 -189
rect -520 189 -320 202
rect -520 143 -507 189
rect -333 143 -320 189
rect -520 100 -320 143
rect -520 -143 -320 -100
rect -520 -189 -507 -143
rect -333 -189 -320 -143
rect -520 -202 -320 -189
rect -240 189 -40 202
rect -240 143 -227 189
rect -53 143 -40 189
rect -240 100 -40 143
rect -240 -143 -40 -100
rect -240 -189 -227 -143
rect -53 -189 -40 -143
rect -240 -202 -40 -189
rect 40 189 240 202
rect 40 143 53 189
rect 227 143 240 189
rect 40 100 240 143
rect 40 -143 240 -100
rect 40 -189 53 -143
rect 227 -189 240 -143
rect 40 -202 240 -189
rect 320 189 520 202
rect 320 143 333 189
rect 507 143 520 189
rect 320 100 520 143
rect 320 -143 520 -100
rect 320 -189 333 -143
rect 507 -189 520 -143
rect 320 -202 520 -189
rect 600 189 800 202
rect 600 143 613 189
rect 787 143 800 189
rect 600 100 800 143
rect 600 -143 800 -100
rect 600 -189 613 -143
rect 787 -189 800 -143
rect 600 -202 800 -189
rect 880 189 1080 202
rect 880 143 893 189
rect 1067 143 1080 189
rect 880 100 1080 143
rect 880 -143 1080 -100
rect 880 -189 893 -143
rect 1067 -189 1080 -143
rect 880 -202 1080 -189
<< polycontact >>
rect -1067 143 -893 189
rect -1067 -189 -893 -143
rect -787 143 -613 189
rect -787 -189 -613 -143
rect -507 143 -333 189
rect -507 -189 -333 -143
rect -227 143 -53 189
rect -227 -189 -53 -143
rect 53 143 227 189
rect 53 -189 227 -143
rect 333 143 507 189
rect 333 -189 507 -143
rect 613 143 787 189
rect 613 -189 787 -143
rect 893 143 1067 189
rect 893 -189 1067 -143
<< ppolyres >>
rect -1080 -100 -880 100
rect -800 -100 -600 100
rect -520 -100 -320 100
rect -240 -100 -40 100
rect 40 -100 240 100
rect 320 -100 520 100
rect 600 -100 800 100
rect 880 -100 1080 100
<< metal1 >>
rect -1078 143 -1067 189
rect -893 143 -882 189
rect -798 143 -787 189
rect -613 143 -602 189
rect -518 143 -507 189
rect -333 143 -322 189
rect -238 143 -227 189
rect -53 143 -42 189
rect 42 143 53 189
rect 227 143 238 189
rect 322 143 333 189
rect 507 143 518 189
rect 602 143 613 189
rect 787 143 798 189
rect 882 143 893 189
rect 1067 143 1078 189
rect -1078 -189 -1067 -143
rect -893 -189 -882 -143
rect -798 -189 -787 -143
rect -613 -189 -602 -143
rect -518 -189 -507 -143
rect -333 -189 -322 -143
rect -238 -189 -227 -143
rect -53 -189 -42 -143
rect 42 -189 53 -143
rect 227 -189 238 -143
rect 322 -189 333 -143
rect 507 -189 518 -143
rect 602 -189 613 -143
rect 787 -189 798 -143
rect 882 -189 893 -143
rect 1067 -189 1078 -143
<< properties >>
string FIXED_BBOX -1204 -326 1204 326
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nx 8 wmin 0.80 lmin 1.00 rho 315 val 338.709 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
