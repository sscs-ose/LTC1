magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2045 -3251 4616 2545
<< nwell >>
rect 0 365 2488 545
rect 280 300 358 363
rect 282 289 358 300
rect 507 233 553 365
rect 1849 355 1945 365
rect 303 80 349 170
rect 619 87 665 164
rect 619 83 681 87
rect 619 82 665 83
rect 253 2 349 80
rect 615 16 687 82
rect 2341 8 2418 10
rect 1852 -76 1926 -8
rect 2341 -66 2421 8
rect 1700 -314 2062 -268
<< polysilicon >>
rect 280 348 358 363
rect 280 314 296 348
rect 172 302 296 314
rect 342 314 358 348
rect 342 302 2314 314
rect 172 278 2314 302
rect 2341 8 2418 10
rect 2341 -6 2421 8
rect 1398 -26 1498 -7
rect 1398 -72 1425 -26
rect 1471 -72 1498 -26
rect 1852 -24 1926 -8
rect 1852 -45 1866 -24
rect 1398 -81 1498 -72
rect 1730 -70 1866 -45
rect 1912 -45 1926 -24
rect 2341 -45 2357 -6
rect 1912 -70 2034 -45
rect 1730 -81 2034 -70
rect 2137 -52 2357 -45
rect 2403 -45 2421 -6
rect 2403 -52 2441 -45
rect 2137 -81 2441 -52
rect 1829 -86 1935 -81
rect 174 -310 274 -266
rect 378 -310 478 -269
rect 582 -305 1498 -269
rect 174 -381 478 -310
rect 174 -409 274 -381
rect 378 -409 478 -381
rect 1130 -315 1498 -305
rect 1130 -409 1230 -315
rect 2168 -372 2250 -359
rect 1742 -373 2250 -372
rect 1742 -408 2184 -373
rect 2183 -419 2184 -408
rect 2230 -408 2250 -373
rect 2230 -419 2232 -408
rect 2183 -424 2232 -419
rect 582 -627 886 -594
rect 1130 -608 1230 -593
rect 1334 -608 1434 -593
rect 1538 -608 1638 -593
rect 582 -649 909 -627
rect 816 -659 909 -649
rect 816 -705 839 -659
rect 885 -705 909 -659
rect 1130 -654 1638 -608
rect 1130 -663 1230 -654
rect 1334 -663 1434 -654
rect 1538 -663 1638 -654
rect 816 -723 909 -705
rect 173 -859 273 -840
rect 377 -859 477 -840
rect 2150 -844 2250 -843
rect 173 -872 477 -859
rect 173 -895 404 -872
rect 173 -912 273 -895
rect 377 -918 404 -895
rect 450 -918 477 -872
rect 1946 -868 2250 -844
rect 1946 -896 2175 -868
rect 377 -954 477 -918
rect 2150 -914 2175 -896
rect 2221 -914 2250 -868
rect 2150 -931 2250 -914
<< polycontact >>
rect 296 302 342 348
rect 1425 -72 1471 -26
rect 1866 -70 1912 -24
rect 2357 -52 2403 -6
rect 2184 -419 2230 -373
rect 839 -705 885 -659
rect 404 -918 450 -872
rect 2175 -914 2221 -868
<< metal1 >>
rect -1 460 2488 545
rect 99 -223 145 460
rect 282 350 354 360
rect 282 348 455 350
rect 282 302 296 348
rect 342 302 455 348
rect 282 301 455 302
rect 282 289 354 301
rect 303 80 349 233
rect 253 66 349 80
rect 253 14 271 66
rect 323 14 349 66
rect 253 2 349 14
rect 297 -150 358 -127
rect 409 -150 455 301
rect 297 -153 455 -150
rect 297 -205 303 -153
rect 355 -198 455 -153
rect 507 -35 553 460
rect 711 210 757 233
rect 618 163 757 210
rect 609 138 757 163
rect 915 138 961 460
rect 1112 389 1192 404
rect 1112 337 1127 389
rect 1179 337 1192 389
rect 1112 322 1192 337
rect 609 87 712 138
rect 1119 87 1165 322
rect 1323 137 1369 460
rect 1521 393 1600 407
rect 1521 341 1535 393
rect 1587 341 1600 393
rect 1521 326 1600 341
rect 1527 137 1573 326
rect 1731 138 1777 460
rect 1926 397 2009 409
rect 1926 345 1941 397
rect 1993 345 2009 397
rect 1926 331 2009 345
rect 1935 90 1981 331
rect 2139 221 2185 460
rect 2115 201 2198 221
rect 2115 149 2131 201
rect 2183 149 2198 201
rect 2115 136 2198 149
rect 2343 91 2389 233
rect 2343 90 2400 91
rect 609 83 1165 87
rect 609 31 623 83
rect 675 33 1165 83
rect 1422 43 2400 90
rect 675 31 712 33
rect 609 14 712 31
rect 1422 -14 1485 43
rect 2354 8 2400 43
rect 2354 -6 2418 8
rect 1407 -26 1485 -14
rect 1851 -20 1928 -11
rect 1812 -21 1928 -20
rect 1812 -23 1864 -21
rect 507 -81 1277 -35
rect 355 -205 358 -198
rect 297 -225 358 -205
rect 507 -223 553 -81
rect 711 -269 757 -127
rect 915 -223 961 -81
rect 1119 -269 1165 -127
rect 1231 -162 1277 -81
rect 1407 -72 1425 -26
rect 1471 -72 1485 -26
rect 1407 -80 1485 -72
rect 1811 -73 1864 -23
rect 1916 -73 1928 -21
rect 1811 -74 1928 -73
rect 2354 -52 2357 -6
rect 2403 -52 2418 -6
rect 2354 -66 2418 -52
rect 1855 -78 1923 -74
rect 2354 -76 2410 -66
rect 1407 -83 1484 -80
rect 1323 -162 1369 -127
rect 1231 -211 1369 -162
rect 1323 -223 1369 -211
rect 711 -315 1305 -269
rect 262 -318 349 -315
rect 711 -317 1190 -315
rect 262 -370 278 -318
rect 330 -370 349 -318
rect 262 -374 349 -370
rect 99 -465 145 -452
rect 94 -479 171 -465
rect 94 -531 107 -479
rect 159 -531 171 -479
rect 94 -545 171 -531
rect 99 -548 145 -545
rect 303 -548 349 -374
rect 1259 -360 1305 -315
rect 1527 -360 1573 -127
rect 1654 -268 1701 -127
rect 1859 -138 1905 -127
rect 1859 -150 1929 -138
rect 2062 -140 2109 -127
rect 1859 -202 1865 -150
rect 1917 -202 1929 -150
rect 1859 -214 1929 -202
rect 1859 -221 1905 -214
rect 2056 -217 2110 -140
rect 2266 -146 2312 -127
rect 2362 -146 2410 -76
rect 2266 -192 2410 -146
rect 2062 -263 2109 -217
rect 2266 -221 2312 -192
rect 2061 -267 2109 -263
rect 2471 -267 2517 -127
rect 2061 -268 2517 -267
rect 1654 -313 2517 -268
rect 1654 -314 2111 -313
rect 1259 -406 2021 -360
rect 516 -474 573 -461
rect 516 -526 518 -474
rect 570 -526 573 -474
rect 516 -538 573 -526
rect 98 -651 552 -605
rect 98 -794 145 -651
rect 302 -708 348 -699
rect 302 -723 374 -708
rect 302 -775 310 -723
rect 362 -775 374 -723
rect 302 -789 374 -775
rect 505 -770 552 -651
rect 302 -793 348 -789
rect 505 -794 573 -770
rect 505 -807 599 -794
rect 505 -816 534 -807
rect 377 -855 452 -852
rect 377 -872 466 -855
rect 522 -859 534 -816
rect 586 -859 599 -807
rect 522 -865 599 -859
rect 377 -873 404 -872
rect 377 -925 395 -873
rect 450 -918 466 -872
rect 447 -925 466 -918
rect 377 -938 466 -925
rect 377 -944 452 -938
rect 711 -994 757 -455
rect 915 -469 961 -452
rect 895 -482 973 -469
rect 895 -534 907 -482
rect 959 -534 973 -482
rect 895 -547 973 -534
rect 915 -548 961 -547
rect 1055 -598 1101 -453
rect 1259 -548 1305 -406
rect 1463 -598 1509 -453
rect 1667 -548 1713 -406
rect 819 -659 898 -642
rect 819 -711 835 -659
rect 887 -711 898 -659
rect 819 -723 898 -711
rect 1055 -645 1509 -598
rect 832 -728 893 -723
rect 1055 -805 1101 -645
rect 1259 -721 1305 -709
rect 1258 -933 1305 -721
rect 1463 -805 1509 -645
rect 1871 -601 1917 -452
rect 1975 -463 2021 -406
rect 2181 -373 2486 -359
rect 2181 -419 2184 -373
rect 2230 -405 2486 -373
rect 2230 -419 2233 -405
rect 2181 -430 2233 -419
rect 2075 -463 2121 -452
rect 1975 -483 2124 -463
rect 1975 -532 2065 -483
rect 2047 -535 2065 -532
rect 2117 -535 2124 -483
rect 2047 -553 2124 -535
rect 2279 -601 2325 -451
rect 2439 -455 2486 -405
rect 2439 -463 2517 -455
rect 2439 -469 2518 -463
rect 2439 -521 2457 -469
rect 2509 -521 2518 -469
rect 2439 -534 2518 -521
rect 1871 -648 2325 -601
rect 1258 -994 1304 -933
rect 1667 -994 1713 -709
rect 1871 -788 1917 -648
rect 2052 -730 2121 -703
rect 2052 -782 2060 -730
rect 2112 -782 2121 -730
rect 2052 -789 2121 -782
rect 2052 -794 2117 -789
rect 2052 -797 2100 -794
rect 2162 -862 2232 -855
rect 2107 -868 2232 -862
rect 2107 -914 2175 -868
rect 2221 -914 2232 -868
rect 2107 -915 2232 -914
rect 2162 -925 2232 -915
rect 2279 -994 2325 -648
rect 29 -1186 2367 -994
<< via1 >>
rect 271 14 323 66
rect 303 -205 355 -153
rect 1127 337 1179 389
rect 1535 341 1587 393
rect 1941 345 1993 397
rect 2131 149 2183 201
rect 623 31 675 83
rect 1864 -24 1916 -21
rect 1864 -70 1866 -24
rect 1866 -70 1912 -24
rect 1912 -70 1916 -24
rect 1864 -73 1916 -70
rect 278 -370 330 -318
rect 107 -531 159 -479
rect 1865 -202 1917 -150
rect 518 -526 570 -474
rect 310 -775 362 -723
rect 534 -859 586 -807
rect 395 -918 404 -873
rect 404 -918 447 -873
rect 395 -925 447 -918
rect 907 -534 959 -482
rect 835 -705 839 -659
rect 839 -705 885 -659
rect 885 -705 887 -659
rect 835 -711 887 -705
rect 2065 -535 2117 -483
rect 2457 -521 2509 -469
rect 2060 -782 2112 -730
<< metal2 >>
rect 1112 395 1192 404
rect 1521 397 1600 407
rect 1926 397 2009 409
rect 1521 395 1941 397
rect 1112 393 1941 395
rect 1112 389 1535 393
rect 1112 337 1127 389
rect 1179 341 1535 389
rect 1587 345 1941 393
rect 1993 345 2009 397
rect 1587 341 2009 345
rect 1179 339 2009 341
rect 1179 337 1600 339
rect 1112 336 1600 337
rect 1112 322 1192 336
rect 1521 326 1600 336
rect 1926 331 2009 339
rect 2125 221 2190 226
rect 2115 201 2198 221
rect 609 83 712 163
rect 2115 149 2131 201
rect 2183 149 2198 201
rect 2115 132 2198 149
rect 257 70 339 77
rect 609 70 623 83
rect 257 66 623 70
rect 257 14 271 66
rect 323 31 623 66
rect 675 31 712 83
rect 323 14 712 31
rect 257 2 339 14
rect 297 -148 358 -127
rect -45 -153 358 -148
rect -45 -204 303 -153
rect -45 -717 11 -204
rect 297 -205 303 -204
rect 355 -205 358 -153
rect 297 -225 358 -205
rect 623 -314 679 14
rect 1851 -16 1929 -8
rect 1776 -21 1929 -16
rect 1776 -73 1864 -21
rect 1916 -73 1929 -21
rect 1776 -74 1929 -73
rect 1851 -78 1929 -74
rect 2125 -148 2190 132
rect 1853 -150 2190 -148
rect 1853 -202 1865 -150
rect 1917 -202 2190 -150
rect 1853 -214 2190 -202
rect 2246 19 2603 84
rect 262 -318 679 -314
rect 262 -370 278 -318
rect 330 -370 679 -318
rect 262 -374 679 -370
rect 276 -381 332 -374
rect 94 -476 171 -465
rect 507 -472 578 -452
rect 895 -472 973 -469
rect 507 -474 973 -472
rect 507 -476 518 -474
rect 94 -479 518 -476
rect 94 -531 107 -479
rect 159 -526 518 -479
rect 570 -482 973 -474
rect 570 -526 907 -482
rect 159 -528 907 -526
rect 159 -531 578 -528
rect 94 -532 578 -531
rect 94 -545 171 -532
rect 507 -548 578 -532
rect 895 -534 907 -528
rect 959 -534 973 -482
rect 895 -547 973 -534
rect 2050 -476 2125 -471
rect 2246 -476 2311 19
rect 2050 -483 2311 -476
rect 2050 -535 2065 -483
rect 2117 -535 2311 -483
rect 2443 -469 2524 -455
rect 2443 -491 2457 -469
rect 2050 -540 2311 -535
rect 2440 -521 2457 -491
rect 2509 -521 2524 -469
rect 2440 -533 2524 -521
rect 2050 -553 2125 -540
rect 310 -650 366 -646
rect 814 -650 901 -642
rect 310 -659 901 -650
rect 310 -708 835 -659
rect 307 -710 835 -708
rect 307 -717 374 -710
rect -45 -723 374 -717
rect 814 -711 835 -710
rect 887 -711 901 -659
rect 814 -722 901 -711
rect 814 -723 900 -722
rect -45 -773 310 -723
rect 307 -775 310 -773
rect 362 -775 374 -723
rect 2055 -726 2128 -717
rect 307 -789 374 -775
rect 1461 -730 2128 -726
rect 1461 -782 2060 -730
rect 2112 -782 2128 -730
rect 1461 -785 2128 -782
rect 522 -801 599 -794
rect 1461 -801 1520 -785
rect 2055 -797 2128 -785
rect 522 -807 1520 -801
rect 368 -873 462 -847
rect 522 -859 534 -807
rect 586 -859 1520 -807
rect 522 -860 1520 -859
rect 522 -865 599 -860
rect 368 -925 395 -873
rect 447 -925 462 -873
rect 368 -960 462 -925
rect 391 -1195 447 -960
rect 2440 -1195 2496 -533
rect 391 -1251 2496 -1195
use nmos_3p3_3JEA4B  nmos_3p3_3JEA4B_0
timestamp 1713185578
transform 1 0 1996 0 1 -502
box -366 -118 366 118
use nmos_3p3_3JEA4B  nmos_3p3_3JEA4B_1
timestamp 1713185578
transform 1 0 1384 0 1 -502
box -366 -118 366 118
use nmos_3p3_3JEA4B  nmos_3p3_3JEA4B_2
timestamp 1713185578
transform 1 0 1384 0 1 -757
box -366 -118 366 118
use nmos_3p3_8FEA4B  nmos_3p3_8FEA4B_0
timestamp 1713185578
transform 1 0 734 0 1 -503
box -264 -118 264 118
use nmos_3p3_8FEA4B  nmos_3p3_8FEA4B_1
timestamp 1713185578
transform 1 0 326 0 1 -503
box -264 -118 264 118
use nmos_3p3_8FEA4B  nmos_3p3_8FEA4B_2
timestamp 1713185578
transform 1 0 325 0 1 -746
box -264 -118 264 118
use nmos_3p3_8FEA4B  nmos_3p3_8FEA4B_3
timestamp 1713185578
transform 1 0 2098 0 1 -750
box -264 -118 264 118
use pmos_3p3_HMK9E7  pmos_3p3_HMK9E7_0
timestamp 1713185578
transform 1 0 1244 0 1 185
box -1244 -180 1244 180
use pmos_3p3_K82TLV  pmos_3p3_K82TLV_0
timestamp 1713185578
transform 1 0 1448 0 1 -175
box -224 -180 224 180
use pmos_3p3_KG2TLV  pmos_3p3_KG2TLV_0
timestamp 1713185578
transform 1 0 2290 0 1 -173
box -326 -180 326 180
use pmos_3p3_KG2TLV  pmos_3p3_KG2TLV_1
timestamp 1713185578
transform 1 0 326 0 1 -175
box -326 -180 326 180
use pmos_3p3_KG2TLV  pmos_3p3_KG2TLV_2
timestamp 1713185578
transform 1 0 1882 0 1 -173
box -326 -180 326 180
use pmos_3p3_KG2TLV  pmos_3p3_KG2TLV_3
timestamp 1713185578
transform 1 0 734 0 1 -175
box -326 -180 326 180
use pmos_3p3_KG2TLV  pmos_3p3_KG2TLV_4
timestamp 1713185578
transform 1 0 1142 0 1 -175
box -326 -180 326 180
<< end >>
