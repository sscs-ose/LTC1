magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1745 -6563 1745 6563
<< metal3 >>
rect -745 5558 745 5563
rect -745 5530 -740 5558
rect -712 5530 -674 5558
rect -646 5530 -608 5558
rect -580 5530 -542 5558
rect -514 5530 -476 5558
rect -448 5530 -410 5558
rect -382 5530 -344 5558
rect -316 5530 -278 5558
rect -250 5530 -212 5558
rect -184 5530 -146 5558
rect -118 5530 -80 5558
rect -52 5530 -14 5558
rect 14 5530 52 5558
rect 80 5530 118 5558
rect 146 5530 184 5558
rect 212 5530 250 5558
rect 278 5530 316 5558
rect 344 5530 382 5558
rect 410 5530 448 5558
rect 476 5530 514 5558
rect 542 5530 580 5558
rect 608 5530 646 5558
rect 674 5530 712 5558
rect 740 5530 745 5558
rect -745 5492 745 5530
rect -745 5464 -740 5492
rect -712 5464 -674 5492
rect -646 5464 -608 5492
rect -580 5464 -542 5492
rect -514 5464 -476 5492
rect -448 5464 -410 5492
rect -382 5464 -344 5492
rect -316 5464 -278 5492
rect -250 5464 -212 5492
rect -184 5464 -146 5492
rect -118 5464 -80 5492
rect -52 5464 -14 5492
rect 14 5464 52 5492
rect 80 5464 118 5492
rect 146 5464 184 5492
rect 212 5464 250 5492
rect 278 5464 316 5492
rect 344 5464 382 5492
rect 410 5464 448 5492
rect 476 5464 514 5492
rect 542 5464 580 5492
rect 608 5464 646 5492
rect 674 5464 712 5492
rect 740 5464 745 5492
rect -745 5426 745 5464
rect -745 5398 -740 5426
rect -712 5398 -674 5426
rect -646 5398 -608 5426
rect -580 5398 -542 5426
rect -514 5398 -476 5426
rect -448 5398 -410 5426
rect -382 5398 -344 5426
rect -316 5398 -278 5426
rect -250 5398 -212 5426
rect -184 5398 -146 5426
rect -118 5398 -80 5426
rect -52 5398 -14 5426
rect 14 5398 52 5426
rect 80 5398 118 5426
rect 146 5398 184 5426
rect 212 5398 250 5426
rect 278 5398 316 5426
rect 344 5398 382 5426
rect 410 5398 448 5426
rect 476 5398 514 5426
rect 542 5398 580 5426
rect 608 5398 646 5426
rect 674 5398 712 5426
rect 740 5398 745 5426
rect -745 5360 745 5398
rect -745 5332 -740 5360
rect -712 5332 -674 5360
rect -646 5332 -608 5360
rect -580 5332 -542 5360
rect -514 5332 -476 5360
rect -448 5332 -410 5360
rect -382 5332 -344 5360
rect -316 5332 -278 5360
rect -250 5332 -212 5360
rect -184 5332 -146 5360
rect -118 5332 -80 5360
rect -52 5332 -14 5360
rect 14 5332 52 5360
rect 80 5332 118 5360
rect 146 5332 184 5360
rect 212 5332 250 5360
rect 278 5332 316 5360
rect 344 5332 382 5360
rect 410 5332 448 5360
rect 476 5332 514 5360
rect 542 5332 580 5360
rect 608 5332 646 5360
rect 674 5332 712 5360
rect 740 5332 745 5360
rect -745 5294 745 5332
rect -745 5266 -740 5294
rect -712 5266 -674 5294
rect -646 5266 -608 5294
rect -580 5266 -542 5294
rect -514 5266 -476 5294
rect -448 5266 -410 5294
rect -382 5266 -344 5294
rect -316 5266 -278 5294
rect -250 5266 -212 5294
rect -184 5266 -146 5294
rect -118 5266 -80 5294
rect -52 5266 -14 5294
rect 14 5266 52 5294
rect 80 5266 118 5294
rect 146 5266 184 5294
rect 212 5266 250 5294
rect 278 5266 316 5294
rect 344 5266 382 5294
rect 410 5266 448 5294
rect 476 5266 514 5294
rect 542 5266 580 5294
rect 608 5266 646 5294
rect 674 5266 712 5294
rect 740 5266 745 5294
rect -745 5228 745 5266
rect -745 5200 -740 5228
rect -712 5200 -674 5228
rect -646 5200 -608 5228
rect -580 5200 -542 5228
rect -514 5200 -476 5228
rect -448 5200 -410 5228
rect -382 5200 -344 5228
rect -316 5200 -278 5228
rect -250 5200 -212 5228
rect -184 5200 -146 5228
rect -118 5200 -80 5228
rect -52 5200 -14 5228
rect 14 5200 52 5228
rect 80 5200 118 5228
rect 146 5200 184 5228
rect 212 5200 250 5228
rect 278 5200 316 5228
rect 344 5200 382 5228
rect 410 5200 448 5228
rect 476 5200 514 5228
rect 542 5200 580 5228
rect 608 5200 646 5228
rect 674 5200 712 5228
rect 740 5200 745 5228
rect -745 5162 745 5200
rect -745 5134 -740 5162
rect -712 5134 -674 5162
rect -646 5134 -608 5162
rect -580 5134 -542 5162
rect -514 5134 -476 5162
rect -448 5134 -410 5162
rect -382 5134 -344 5162
rect -316 5134 -278 5162
rect -250 5134 -212 5162
rect -184 5134 -146 5162
rect -118 5134 -80 5162
rect -52 5134 -14 5162
rect 14 5134 52 5162
rect 80 5134 118 5162
rect 146 5134 184 5162
rect 212 5134 250 5162
rect 278 5134 316 5162
rect 344 5134 382 5162
rect 410 5134 448 5162
rect 476 5134 514 5162
rect 542 5134 580 5162
rect 608 5134 646 5162
rect 674 5134 712 5162
rect 740 5134 745 5162
rect -745 5096 745 5134
rect -745 5068 -740 5096
rect -712 5068 -674 5096
rect -646 5068 -608 5096
rect -580 5068 -542 5096
rect -514 5068 -476 5096
rect -448 5068 -410 5096
rect -382 5068 -344 5096
rect -316 5068 -278 5096
rect -250 5068 -212 5096
rect -184 5068 -146 5096
rect -118 5068 -80 5096
rect -52 5068 -14 5096
rect 14 5068 52 5096
rect 80 5068 118 5096
rect 146 5068 184 5096
rect 212 5068 250 5096
rect 278 5068 316 5096
rect 344 5068 382 5096
rect 410 5068 448 5096
rect 476 5068 514 5096
rect 542 5068 580 5096
rect 608 5068 646 5096
rect 674 5068 712 5096
rect 740 5068 745 5096
rect -745 5030 745 5068
rect -745 5002 -740 5030
rect -712 5002 -674 5030
rect -646 5002 -608 5030
rect -580 5002 -542 5030
rect -514 5002 -476 5030
rect -448 5002 -410 5030
rect -382 5002 -344 5030
rect -316 5002 -278 5030
rect -250 5002 -212 5030
rect -184 5002 -146 5030
rect -118 5002 -80 5030
rect -52 5002 -14 5030
rect 14 5002 52 5030
rect 80 5002 118 5030
rect 146 5002 184 5030
rect 212 5002 250 5030
rect 278 5002 316 5030
rect 344 5002 382 5030
rect 410 5002 448 5030
rect 476 5002 514 5030
rect 542 5002 580 5030
rect 608 5002 646 5030
rect 674 5002 712 5030
rect 740 5002 745 5030
rect -745 4964 745 5002
rect -745 4936 -740 4964
rect -712 4936 -674 4964
rect -646 4936 -608 4964
rect -580 4936 -542 4964
rect -514 4936 -476 4964
rect -448 4936 -410 4964
rect -382 4936 -344 4964
rect -316 4936 -278 4964
rect -250 4936 -212 4964
rect -184 4936 -146 4964
rect -118 4936 -80 4964
rect -52 4936 -14 4964
rect 14 4936 52 4964
rect 80 4936 118 4964
rect 146 4936 184 4964
rect 212 4936 250 4964
rect 278 4936 316 4964
rect 344 4936 382 4964
rect 410 4936 448 4964
rect 476 4936 514 4964
rect 542 4936 580 4964
rect 608 4936 646 4964
rect 674 4936 712 4964
rect 740 4936 745 4964
rect -745 4898 745 4936
rect -745 4870 -740 4898
rect -712 4870 -674 4898
rect -646 4870 -608 4898
rect -580 4870 -542 4898
rect -514 4870 -476 4898
rect -448 4870 -410 4898
rect -382 4870 -344 4898
rect -316 4870 -278 4898
rect -250 4870 -212 4898
rect -184 4870 -146 4898
rect -118 4870 -80 4898
rect -52 4870 -14 4898
rect 14 4870 52 4898
rect 80 4870 118 4898
rect 146 4870 184 4898
rect 212 4870 250 4898
rect 278 4870 316 4898
rect 344 4870 382 4898
rect 410 4870 448 4898
rect 476 4870 514 4898
rect 542 4870 580 4898
rect 608 4870 646 4898
rect 674 4870 712 4898
rect 740 4870 745 4898
rect -745 4832 745 4870
rect -745 4804 -740 4832
rect -712 4804 -674 4832
rect -646 4804 -608 4832
rect -580 4804 -542 4832
rect -514 4804 -476 4832
rect -448 4804 -410 4832
rect -382 4804 -344 4832
rect -316 4804 -278 4832
rect -250 4804 -212 4832
rect -184 4804 -146 4832
rect -118 4804 -80 4832
rect -52 4804 -14 4832
rect 14 4804 52 4832
rect 80 4804 118 4832
rect 146 4804 184 4832
rect 212 4804 250 4832
rect 278 4804 316 4832
rect 344 4804 382 4832
rect 410 4804 448 4832
rect 476 4804 514 4832
rect 542 4804 580 4832
rect 608 4804 646 4832
rect 674 4804 712 4832
rect 740 4804 745 4832
rect -745 4766 745 4804
rect -745 4738 -740 4766
rect -712 4738 -674 4766
rect -646 4738 -608 4766
rect -580 4738 -542 4766
rect -514 4738 -476 4766
rect -448 4738 -410 4766
rect -382 4738 -344 4766
rect -316 4738 -278 4766
rect -250 4738 -212 4766
rect -184 4738 -146 4766
rect -118 4738 -80 4766
rect -52 4738 -14 4766
rect 14 4738 52 4766
rect 80 4738 118 4766
rect 146 4738 184 4766
rect 212 4738 250 4766
rect 278 4738 316 4766
rect 344 4738 382 4766
rect 410 4738 448 4766
rect 476 4738 514 4766
rect 542 4738 580 4766
rect 608 4738 646 4766
rect 674 4738 712 4766
rect 740 4738 745 4766
rect -745 4700 745 4738
rect -745 4672 -740 4700
rect -712 4672 -674 4700
rect -646 4672 -608 4700
rect -580 4672 -542 4700
rect -514 4672 -476 4700
rect -448 4672 -410 4700
rect -382 4672 -344 4700
rect -316 4672 -278 4700
rect -250 4672 -212 4700
rect -184 4672 -146 4700
rect -118 4672 -80 4700
rect -52 4672 -14 4700
rect 14 4672 52 4700
rect 80 4672 118 4700
rect 146 4672 184 4700
rect 212 4672 250 4700
rect 278 4672 316 4700
rect 344 4672 382 4700
rect 410 4672 448 4700
rect 476 4672 514 4700
rect 542 4672 580 4700
rect 608 4672 646 4700
rect 674 4672 712 4700
rect 740 4672 745 4700
rect -745 4634 745 4672
rect -745 4606 -740 4634
rect -712 4606 -674 4634
rect -646 4606 -608 4634
rect -580 4606 -542 4634
rect -514 4606 -476 4634
rect -448 4606 -410 4634
rect -382 4606 -344 4634
rect -316 4606 -278 4634
rect -250 4606 -212 4634
rect -184 4606 -146 4634
rect -118 4606 -80 4634
rect -52 4606 -14 4634
rect 14 4606 52 4634
rect 80 4606 118 4634
rect 146 4606 184 4634
rect 212 4606 250 4634
rect 278 4606 316 4634
rect 344 4606 382 4634
rect 410 4606 448 4634
rect 476 4606 514 4634
rect 542 4606 580 4634
rect 608 4606 646 4634
rect 674 4606 712 4634
rect 740 4606 745 4634
rect -745 4568 745 4606
rect -745 4540 -740 4568
rect -712 4540 -674 4568
rect -646 4540 -608 4568
rect -580 4540 -542 4568
rect -514 4540 -476 4568
rect -448 4540 -410 4568
rect -382 4540 -344 4568
rect -316 4540 -278 4568
rect -250 4540 -212 4568
rect -184 4540 -146 4568
rect -118 4540 -80 4568
rect -52 4540 -14 4568
rect 14 4540 52 4568
rect 80 4540 118 4568
rect 146 4540 184 4568
rect 212 4540 250 4568
rect 278 4540 316 4568
rect 344 4540 382 4568
rect 410 4540 448 4568
rect 476 4540 514 4568
rect 542 4540 580 4568
rect 608 4540 646 4568
rect 674 4540 712 4568
rect 740 4540 745 4568
rect -745 4502 745 4540
rect -745 4474 -740 4502
rect -712 4474 -674 4502
rect -646 4474 -608 4502
rect -580 4474 -542 4502
rect -514 4474 -476 4502
rect -448 4474 -410 4502
rect -382 4474 -344 4502
rect -316 4474 -278 4502
rect -250 4474 -212 4502
rect -184 4474 -146 4502
rect -118 4474 -80 4502
rect -52 4474 -14 4502
rect 14 4474 52 4502
rect 80 4474 118 4502
rect 146 4474 184 4502
rect 212 4474 250 4502
rect 278 4474 316 4502
rect 344 4474 382 4502
rect 410 4474 448 4502
rect 476 4474 514 4502
rect 542 4474 580 4502
rect 608 4474 646 4502
rect 674 4474 712 4502
rect 740 4474 745 4502
rect -745 4436 745 4474
rect -745 4408 -740 4436
rect -712 4408 -674 4436
rect -646 4408 -608 4436
rect -580 4408 -542 4436
rect -514 4408 -476 4436
rect -448 4408 -410 4436
rect -382 4408 -344 4436
rect -316 4408 -278 4436
rect -250 4408 -212 4436
rect -184 4408 -146 4436
rect -118 4408 -80 4436
rect -52 4408 -14 4436
rect 14 4408 52 4436
rect 80 4408 118 4436
rect 146 4408 184 4436
rect 212 4408 250 4436
rect 278 4408 316 4436
rect 344 4408 382 4436
rect 410 4408 448 4436
rect 476 4408 514 4436
rect 542 4408 580 4436
rect 608 4408 646 4436
rect 674 4408 712 4436
rect 740 4408 745 4436
rect -745 4370 745 4408
rect -745 4342 -740 4370
rect -712 4342 -674 4370
rect -646 4342 -608 4370
rect -580 4342 -542 4370
rect -514 4342 -476 4370
rect -448 4342 -410 4370
rect -382 4342 -344 4370
rect -316 4342 -278 4370
rect -250 4342 -212 4370
rect -184 4342 -146 4370
rect -118 4342 -80 4370
rect -52 4342 -14 4370
rect 14 4342 52 4370
rect 80 4342 118 4370
rect 146 4342 184 4370
rect 212 4342 250 4370
rect 278 4342 316 4370
rect 344 4342 382 4370
rect 410 4342 448 4370
rect 476 4342 514 4370
rect 542 4342 580 4370
rect 608 4342 646 4370
rect 674 4342 712 4370
rect 740 4342 745 4370
rect -745 4304 745 4342
rect -745 4276 -740 4304
rect -712 4276 -674 4304
rect -646 4276 -608 4304
rect -580 4276 -542 4304
rect -514 4276 -476 4304
rect -448 4276 -410 4304
rect -382 4276 -344 4304
rect -316 4276 -278 4304
rect -250 4276 -212 4304
rect -184 4276 -146 4304
rect -118 4276 -80 4304
rect -52 4276 -14 4304
rect 14 4276 52 4304
rect 80 4276 118 4304
rect 146 4276 184 4304
rect 212 4276 250 4304
rect 278 4276 316 4304
rect 344 4276 382 4304
rect 410 4276 448 4304
rect 476 4276 514 4304
rect 542 4276 580 4304
rect 608 4276 646 4304
rect 674 4276 712 4304
rect 740 4276 745 4304
rect -745 4238 745 4276
rect -745 4210 -740 4238
rect -712 4210 -674 4238
rect -646 4210 -608 4238
rect -580 4210 -542 4238
rect -514 4210 -476 4238
rect -448 4210 -410 4238
rect -382 4210 -344 4238
rect -316 4210 -278 4238
rect -250 4210 -212 4238
rect -184 4210 -146 4238
rect -118 4210 -80 4238
rect -52 4210 -14 4238
rect 14 4210 52 4238
rect 80 4210 118 4238
rect 146 4210 184 4238
rect 212 4210 250 4238
rect 278 4210 316 4238
rect 344 4210 382 4238
rect 410 4210 448 4238
rect 476 4210 514 4238
rect 542 4210 580 4238
rect 608 4210 646 4238
rect 674 4210 712 4238
rect 740 4210 745 4238
rect -745 4172 745 4210
rect -745 4144 -740 4172
rect -712 4144 -674 4172
rect -646 4144 -608 4172
rect -580 4144 -542 4172
rect -514 4144 -476 4172
rect -448 4144 -410 4172
rect -382 4144 -344 4172
rect -316 4144 -278 4172
rect -250 4144 -212 4172
rect -184 4144 -146 4172
rect -118 4144 -80 4172
rect -52 4144 -14 4172
rect 14 4144 52 4172
rect 80 4144 118 4172
rect 146 4144 184 4172
rect 212 4144 250 4172
rect 278 4144 316 4172
rect 344 4144 382 4172
rect 410 4144 448 4172
rect 476 4144 514 4172
rect 542 4144 580 4172
rect 608 4144 646 4172
rect 674 4144 712 4172
rect 740 4144 745 4172
rect -745 4106 745 4144
rect -745 4078 -740 4106
rect -712 4078 -674 4106
rect -646 4078 -608 4106
rect -580 4078 -542 4106
rect -514 4078 -476 4106
rect -448 4078 -410 4106
rect -382 4078 -344 4106
rect -316 4078 -278 4106
rect -250 4078 -212 4106
rect -184 4078 -146 4106
rect -118 4078 -80 4106
rect -52 4078 -14 4106
rect 14 4078 52 4106
rect 80 4078 118 4106
rect 146 4078 184 4106
rect 212 4078 250 4106
rect 278 4078 316 4106
rect 344 4078 382 4106
rect 410 4078 448 4106
rect 476 4078 514 4106
rect 542 4078 580 4106
rect 608 4078 646 4106
rect 674 4078 712 4106
rect 740 4078 745 4106
rect -745 4040 745 4078
rect -745 4012 -740 4040
rect -712 4012 -674 4040
rect -646 4012 -608 4040
rect -580 4012 -542 4040
rect -514 4012 -476 4040
rect -448 4012 -410 4040
rect -382 4012 -344 4040
rect -316 4012 -278 4040
rect -250 4012 -212 4040
rect -184 4012 -146 4040
rect -118 4012 -80 4040
rect -52 4012 -14 4040
rect 14 4012 52 4040
rect 80 4012 118 4040
rect 146 4012 184 4040
rect 212 4012 250 4040
rect 278 4012 316 4040
rect 344 4012 382 4040
rect 410 4012 448 4040
rect 476 4012 514 4040
rect 542 4012 580 4040
rect 608 4012 646 4040
rect 674 4012 712 4040
rect 740 4012 745 4040
rect -745 3974 745 4012
rect -745 3946 -740 3974
rect -712 3946 -674 3974
rect -646 3946 -608 3974
rect -580 3946 -542 3974
rect -514 3946 -476 3974
rect -448 3946 -410 3974
rect -382 3946 -344 3974
rect -316 3946 -278 3974
rect -250 3946 -212 3974
rect -184 3946 -146 3974
rect -118 3946 -80 3974
rect -52 3946 -14 3974
rect 14 3946 52 3974
rect 80 3946 118 3974
rect 146 3946 184 3974
rect 212 3946 250 3974
rect 278 3946 316 3974
rect 344 3946 382 3974
rect 410 3946 448 3974
rect 476 3946 514 3974
rect 542 3946 580 3974
rect 608 3946 646 3974
rect 674 3946 712 3974
rect 740 3946 745 3974
rect -745 3908 745 3946
rect -745 3880 -740 3908
rect -712 3880 -674 3908
rect -646 3880 -608 3908
rect -580 3880 -542 3908
rect -514 3880 -476 3908
rect -448 3880 -410 3908
rect -382 3880 -344 3908
rect -316 3880 -278 3908
rect -250 3880 -212 3908
rect -184 3880 -146 3908
rect -118 3880 -80 3908
rect -52 3880 -14 3908
rect 14 3880 52 3908
rect 80 3880 118 3908
rect 146 3880 184 3908
rect 212 3880 250 3908
rect 278 3880 316 3908
rect 344 3880 382 3908
rect 410 3880 448 3908
rect 476 3880 514 3908
rect 542 3880 580 3908
rect 608 3880 646 3908
rect 674 3880 712 3908
rect 740 3880 745 3908
rect -745 3842 745 3880
rect -745 3814 -740 3842
rect -712 3814 -674 3842
rect -646 3814 -608 3842
rect -580 3814 -542 3842
rect -514 3814 -476 3842
rect -448 3814 -410 3842
rect -382 3814 -344 3842
rect -316 3814 -278 3842
rect -250 3814 -212 3842
rect -184 3814 -146 3842
rect -118 3814 -80 3842
rect -52 3814 -14 3842
rect 14 3814 52 3842
rect 80 3814 118 3842
rect 146 3814 184 3842
rect 212 3814 250 3842
rect 278 3814 316 3842
rect 344 3814 382 3842
rect 410 3814 448 3842
rect 476 3814 514 3842
rect 542 3814 580 3842
rect 608 3814 646 3842
rect 674 3814 712 3842
rect 740 3814 745 3842
rect -745 3776 745 3814
rect -745 3748 -740 3776
rect -712 3748 -674 3776
rect -646 3748 -608 3776
rect -580 3748 -542 3776
rect -514 3748 -476 3776
rect -448 3748 -410 3776
rect -382 3748 -344 3776
rect -316 3748 -278 3776
rect -250 3748 -212 3776
rect -184 3748 -146 3776
rect -118 3748 -80 3776
rect -52 3748 -14 3776
rect 14 3748 52 3776
rect 80 3748 118 3776
rect 146 3748 184 3776
rect 212 3748 250 3776
rect 278 3748 316 3776
rect 344 3748 382 3776
rect 410 3748 448 3776
rect 476 3748 514 3776
rect 542 3748 580 3776
rect 608 3748 646 3776
rect 674 3748 712 3776
rect 740 3748 745 3776
rect -745 3710 745 3748
rect -745 3682 -740 3710
rect -712 3682 -674 3710
rect -646 3682 -608 3710
rect -580 3682 -542 3710
rect -514 3682 -476 3710
rect -448 3682 -410 3710
rect -382 3682 -344 3710
rect -316 3682 -278 3710
rect -250 3682 -212 3710
rect -184 3682 -146 3710
rect -118 3682 -80 3710
rect -52 3682 -14 3710
rect 14 3682 52 3710
rect 80 3682 118 3710
rect 146 3682 184 3710
rect 212 3682 250 3710
rect 278 3682 316 3710
rect 344 3682 382 3710
rect 410 3682 448 3710
rect 476 3682 514 3710
rect 542 3682 580 3710
rect 608 3682 646 3710
rect 674 3682 712 3710
rect 740 3682 745 3710
rect -745 3644 745 3682
rect -745 3616 -740 3644
rect -712 3616 -674 3644
rect -646 3616 -608 3644
rect -580 3616 -542 3644
rect -514 3616 -476 3644
rect -448 3616 -410 3644
rect -382 3616 -344 3644
rect -316 3616 -278 3644
rect -250 3616 -212 3644
rect -184 3616 -146 3644
rect -118 3616 -80 3644
rect -52 3616 -14 3644
rect 14 3616 52 3644
rect 80 3616 118 3644
rect 146 3616 184 3644
rect 212 3616 250 3644
rect 278 3616 316 3644
rect 344 3616 382 3644
rect 410 3616 448 3644
rect 476 3616 514 3644
rect 542 3616 580 3644
rect 608 3616 646 3644
rect 674 3616 712 3644
rect 740 3616 745 3644
rect -745 3578 745 3616
rect -745 3550 -740 3578
rect -712 3550 -674 3578
rect -646 3550 -608 3578
rect -580 3550 -542 3578
rect -514 3550 -476 3578
rect -448 3550 -410 3578
rect -382 3550 -344 3578
rect -316 3550 -278 3578
rect -250 3550 -212 3578
rect -184 3550 -146 3578
rect -118 3550 -80 3578
rect -52 3550 -14 3578
rect 14 3550 52 3578
rect 80 3550 118 3578
rect 146 3550 184 3578
rect 212 3550 250 3578
rect 278 3550 316 3578
rect 344 3550 382 3578
rect 410 3550 448 3578
rect 476 3550 514 3578
rect 542 3550 580 3578
rect 608 3550 646 3578
rect 674 3550 712 3578
rect 740 3550 745 3578
rect -745 3512 745 3550
rect -745 3484 -740 3512
rect -712 3484 -674 3512
rect -646 3484 -608 3512
rect -580 3484 -542 3512
rect -514 3484 -476 3512
rect -448 3484 -410 3512
rect -382 3484 -344 3512
rect -316 3484 -278 3512
rect -250 3484 -212 3512
rect -184 3484 -146 3512
rect -118 3484 -80 3512
rect -52 3484 -14 3512
rect 14 3484 52 3512
rect 80 3484 118 3512
rect 146 3484 184 3512
rect 212 3484 250 3512
rect 278 3484 316 3512
rect 344 3484 382 3512
rect 410 3484 448 3512
rect 476 3484 514 3512
rect 542 3484 580 3512
rect 608 3484 646 3512
rect 674 3484 712 3512
rect 740 3484 745 3512
rect -745 3446 745 3484
rect -745 3418 -740 3446
rect -712 3418 -674 3446
rect -646 3418 -608 3446
rect -580 3418 -542 3446
rect -514 3418 -476 3446
rect -448 3418 -410 3446
rect -382 3418 -344 3446
rect -316 3418 -278 3446
rect -250 3418 -212 3446
rect -184 3418 -146 3446
rect -118 3418 -80 3446
rect -52 3418 -14 3446
rect 14 3418 52 3446
rect 80 3418 118 3446
rect 146 3418 184 3446
rect 212 3418 250 3446
rect 278 3418 316 3446
rect 344 3418 382 3446
rect 410 3418 448 3446
rect 476 3418 514 3446
rect 542 3418 580 3446
rect 608 3418 646 3446
rect 674 3418 712 3446
rect 740 3418 745 3446
rect -745 3380 745 3418
rect -745 3352 -740 3380
rect -712 3352 -674 3380
rect -646 3352 -608 3380
rect -580 3352 -542 3380
rect -514 3352 -476 3380
rect -448 3352 -410 3380
rect -382 3352 -344 3380
rect -316 3352 -278 3380
rect -250 3352 -212 3380
rect -184 3352 -146 3380
rect -118 3352 -80 3380
rect -52 3352 -14 3380
rect 14 3352 52 3380
rect 80 3352 118 3380
rect 146 3352 184 3380
rect 212 3352 250 3380
rect 278 3352 316 3380
rect 344 3352 382 3380
rect 410 3352 448 3380
rect 476 3352 514 3380
rect 542 3352 580 3380
rect 608 3352 646 3380
rect 674 3352 712 3380
rect 740 3352 745 3380
rect -745 3314 745 3352
rect -745 3286 -740 3314
rect -712 3286 -674 3314
rect -646 3286 -608 3314
rect -580 3286 -542 3314
rect -514 3286 -476 3314
rect -448 3286 -410 3314
rect -382 3286 -344 3314
rect -316 3286 -278 3314
rect -250 3286 -212 3314
rect -184 3286 -146 3314
rect -118 3286 -80 3314
rect -52 3286 -14 3314
rect 14 3286 52 3314
rect 80 3286 118 3314
rect 146 3286 184 3314
rect 212 3286 250 3314
rect 278 3286 316 3314
rect 344 3286 382 3314
rect 410 3286 448 3314
rect 476 3286 514 3314
rect 542 3286 580 3314
rect 608 3286 646 3314
rect 674 3286 712 3314
rect 740 3286 745 3314
rect -745 3248 745 3286
rect -745 3220 -740 3248
rect -712 3220 -674 3248
rect -646 3220 -608 3248
rect -580 3220 -542 3248
rect -514 3220 -476 3248
rect -448 3220 -410 3248
rect -382 3220 -344 3248
rect -316 3220 -278 3248
rect -250 3220 -212 3248
rect -184 3220 -146 3248
rect -118 3220 -80 3248
rect -52 3220 -14 3248
rect 14 3220 52 3248
rect 80 3220 118 3248
rect 146 3220 184 3248
rect 212 3220 250 3248
rect 278 3220 316 3248
rect 344 3220 382 3248
rect 410 3220 448 3248
rect 476 3220 514 3248
rect 542 3220 580 3248
rect 608 3220 646 3248
rect 674 3220 712 3248
rect 740 3220 745 3248
rect -745 3182 745 3220
rect -745 3154 -740 3182
rect -712 3154 -674 3182
rect -646 3154 -608 3182
rect -580 3154 -542 3182
rect -514 3154 -476 3182
rect -448 3154 -410 3182
rect -382 3154 -344 3182
rect -316 3154 -278 3182
rect -250 3154 -212 3182
rect -184 3154 -146 3182
rect -118 3154 -80 3182
rect -52 3154 -14 3182
rect 14 3154 52 3182
rect 80 3154 118 3182
rect 146 3154 184 3182
rect 212 3154 250 3182
rect 278 3154 316 3182
rect 344 3154 382 3182
rect 410 3154 448 3182
rect 476 3154 514 3182
rect 542 3154 580 3182
rect 608 3154 646 3182
rect 674 3154 712 3182
rect 740 3154 745 3182
rect -745 3116 745 3154
rect -745 3088 -740 3116
rect -712 3088 -674 3116
rect -646 3088 -608 3116
rect -580 3088 -542 3116
rect -514 3088 -476 3116
rect -448 3088 -410 3116
rect -382 3088 -344 3116
rect -316 3088 -278 3116
rect -250 3088 -212 3116
rect -184 3088 -146 3116
rect -118 3088 -80 3116
rect -52 3088 -14 3116
rect 14 3088 52 3116
rect 80 3088 118 3116
rect 146 3088 184 3116
rect 212 3088 250 3116
rect 278 3088 316 3116
rect 344 3088 382 3116
rect 410 3088 448 3116
rect 476 3088 514 3116
rect 542 3088 580 3116
rect 608 3088 646 3116
rect 674 3088 712 3116
rect 740 3088 745 3116
rect -745 3050 745 3088
rect -745 3022 -740 3050
rect -712 3022 -674 3050
rect -646 3022 -608 3050
rect -580 3022 -542 3050
rect -514 3022 -476 3050
rect -448 3022 -410 3050
rect -382 3022 -344 3050
rect -316 3022 -278 3050
rect -250 3022 -212 3050
rect -184 3022 -146 3050
rect -118 3022 -80 3050
rect -52 3022 -14 3050
rect 14 3022 52 3050
rect 80 3022 118 3050
rect 146 3022 184 3050
rect 212 3022 250 3050
rect 278 3022 316 3050
rect 344 3022 382 3050
rect 410 3022 448 3050
rect 476 3022 514 3050
rect 542 3022 580 3050
rect 608 3022 646 3050
rect 674 3022 712 3050
rect 740 3022 745 3050
rect -745 2984 745 3022
rect -745 2956 -740 2984
rect -712 2956 -674 2984
rect -646 2956 -608 2984
rect -580 2956 -542 2984
rect -514 2956 -476 2984
rect -448 2956 -410 2984
rect -382 2956 -344 2984
rect -316 2956 -278 2984
rect -250 2956 -212 2984
rect -184 2956 -146 2984
rect -118 2956 -80 2984
rect -52 2956 -14 2984
rect 14 2956 52 2984
rect 80 2956 118 2984
rect 146 2956 184 2984
rect 212 2956 250 2984
rect 278 2956 316 2984
rect 344 2956 382 2984
rect 410 2956 448 2984
rect 476 2956 514 2984
rect 542 2956 580 2984
rect 608 2956 646 2984
rect 674 2956 712 2984
rect 740 2956 745 2984
rect -745 2918 745 2956
rect -745 2890 -740 2918
rect -712 2890 -674 2918
rect -646 2890 -608 2918
rect -580 2890 -542 2918
rect -514 2890 -476 2918
rect -448 2890 -410 2918
rect -382 2890 -344 2918
rect -316 2890 -278 2918
rect -250 2890 -212 2918
rect -184 2890 -146 2918
rect -118 2890 -80 2918
rect -52 2890 -14 2918
rect 14 2890 52 2918
rect 80 2890 118 2918
rect 146 2890 184 2918
rect 212 2890 250 2918
rect 278 2890 316 2918
rect 344 2890 382 2918
rect 410 2890 448 2918
rect 476 2890 514 2918
rect 542 2890 580 2918
rect 608 2890 646 2918
rect 674 2890 712 2918
rect 740 2890 745 2918
rect -745 2852 745 2890
rect -745 2824 -740 2852
rect -712 2824 -674 2852
rect -646 2824 -608 2852
rect -580 2824 -542 2852
rect -514 2824 -476 2852
rect -448 2824 -410 2852
rect -382 2824 -344 2852
rect -316 2824 -278 2852
rect -250 2824 -212 2852
rect -184 2824 -146 2852
rect -118 2824 -80 2852
rect -52 2824 -14 2852
rect 14 2824 52 2852
rect 80 2824 118 2852
rect 146 2824 184 2852
rect 212 2824 250 2852
rect 278 2824 316 2852
rect 344 2824 382 2852
rect 410 2824 448 2852
rect 476 2824 514 2852
rect 542 2824 580 2852
rect 608 2824 646 2852
rect 674 2824 712 2852
rect 740 2824 745 2852
rect -745 2786 745 2824
rect -745 2758 -740 2786
rect -712 2758 -674 2786
rect -646 2758 -608 2786
rect -580 2758 -542 2786
rect -514 2758 -476 2786
rect -448 2758 -410 2786
rect -382 2758 -344 2786
rect -316 2758 -278 2786
rect -250 2758 -212 2786
rect -184 2758 -146 2786
rect -118 2758 -80 2786
rect -52 2758 -14 2786
rect 14 2758 52 2786
rect 80 2758 118 2786
rect 146 2758 184 2786
rect 212 2758 250 2786
rect 278 2758 316 2786
rect 344 2758 382 2786
rect 410 2758 448 2786
rect 476 2758 514 2786
rect 542 2758 580 2786
rect 608 2758 646 2786
rect 674 2758 712 2786
rect 740 2758 745 2786
rect -745 2720 745 2758
rect -745 2692 -740 2720
rect -712 2692 -674 2720
rect -646 2692 -608 2720
rect -580 2692 -542 2720
rect -514 2692 -476 2720
rect -448 2692 -410 2720
rect -382 2692 -344 2720
rect -316 2692 -278 2720
rect -250 2692 -212 2720
rect -184 2692 -146 2720
rect -118 2692 -80 2720
rect -52 2692 -14 2720
rect 14 2692 52 2720
rect 80 2692 118 2720
rect 146 2692 184 2720
rect 212 2692 250 2720
rect 278 2692 316 2720
rect 344 2692 382 2720
rect 410 2692 448 2720
rect 476 2692 514 2720
rect 542 2692 580 2720
rect 608 2692 646 2720
rect 674 2692 712 2720
rect 740 2692 745 2720
rect -745 2654 745 2692
rect -745 2626 -740 2654
rect -712 2626 -674 2654
rect -646 2626 -608 2654
rect -580 2626 -542 2654
rect -514 2626 -476 2654
rect -448 2626 -410 2654
rect -382 2626 -344 2654
rect -316 2626 -278 2654
rect -250 2626 -212 2654
rect -184 2626 -146 2654
rect -118 2626 -80 2654
rect -52 2626 -14 2654
rect 14 2626 52 2654
rect 80 2626 118 2654
rect 146 2626 184 2654
rect 212 2626 250 2654
rect 278 2626 316 2654
rect 344 2626 382 2654
rect 410 2626 448 2654
rect 476 2626 514 2654
rect 542 2626 580 2654
rect 608 2626 646 2654
rect 674 2626 712 2654
rect 740 2626 745 2654
rect -745 2588 745 2626
rect -745 2560 -740 2588
rect -712 2560 -674 2588
rect -646 2560 -608 2588
rect -580 2560 -542 2588
rect -514 2560 -476 2588
rect -448 2560 -410 2588
rect -382 2560 -344 2588
rect -316 2560 -278 2588
rect -250 2560 -212 2588
rect -184 2560 -146 2588
rect -118 2560 -80 2588
rect -52 2560 -14 2588
rect 14 2560 52 2588
rect 80 2560 118 2588
rect 146 2560 184 2588
rect 212 2560 250 2588
rect 278 2560 316 2588
rect 344 2560 382 2588
rect 410 2560 448 2588
rect 476 2560 514 2588
rect 542 2560 580 2588
rect 608 2560 646 2588
rect 674 2560 712 2588
rect 740 2560 745 2588
rect -745 2522 745 2560
rect -745 2494 -740 2522
rect -712 2494 -674 2522
rect -646 2494 -608 2522
rect -580 2494 -542 2522
rect -514 2494 -476 2522
rect -448 2494 -410 2522
rect -382 2494 -344 2522
rect -316 2494 -278 2522
rect -250 2494 -212 2522
rect -184 2494 -146 2522
rect -118 2494 -80 2522
rect -52 2494 -14 2522
rect 14 2494 52 2522
rect 80 2494 118 2522
rect 146 2494 184 2522
rect 212 2494 250 2522
rect 278 2494 316 2522
rect 344 2494 382 2522
rect 410 2494 448 2522
rect 476 2494 514 2522
rect 542 2494 580 2522
rect 608 2494 646 2522
rect 674 2494 712 2522
rect 740 2494 745 2522
rect -745 2456 745 2494
rect -745 2428 -740 2456
rect -712 2428 -674 2456
rect -646 2428 -608 2456
rect -580 2428 -542 2456
rect -514 2428 -476 2456
rect -448 2428 -410 2456
rect -382 2428 -344 2456
rect -316 2428 -278 2456
rect -250 2428 -212 2456
rect -184 2428 -146 2456
rect -118 2428 -80 2456
rect -52 2428 -14 2456
rect 14 2428 52 2456
rect 80 2428 118 2456
rect 146 2428 184 2456
rect 212 2428 250 2456
rect 278 2428 316 2456
rect 344 2428 382 2456
rect 410 2428 448 2456
rect 476 2428 514 2456
rect 542 2428 580 2456
rect 608 2428 646 2456
rect 674 2428 712 2456
rect 740 2428 745 2456
rect -745 2390 745 2428
rect -745 2362 -740 2390
rect -712 2362 -674 2390
rect -646 2362 -608 2390
rect -580 2362 -542 2390
rect -514 2362 -476 2390
rect -448 2362 -410 2390
rect -382 2362 -344 2390
rect -316 2362 -278 2390
rect -250 2362 -212 2390
rect -184 2362 -146 2390
rect -118 2362 -80 2390
rect -52 2362 -14 2390
rect 14 2362 52 2390
rect 80 2362 118 2390
rect 146 2362 184 2390
rect 212 2362 250 2390
rect 278 2362 316 2390
rect 344 2362 382 2390
rect 410 2362 448 2390
rect 476 2362 514 2390
rect 542 2362 580 2390
rect 608 2362 646 2390
rect 674 2362 712 2390
rect 740 2362 745 2390
rect -745 2324 745 2362
rect -745 2296 -740 2324
rect -712 2296 -674 2324
rect -646 2296 -608 2324
rect -580 2296 -542 2324
rect -514 2296 -476 2324
rect -448 2296 -410 2324
rect -382 2296 -344 2324
rect -316 2296 -278 2324
rect -250 2296 -212 2324
rect -184 2296 -146 2324
rect -118 2296 -80 2324
rect -52 2296 -14 2324
rect 14 2296 52 2324
rect 80 2296 118 2324
rect 146 2296 184 2324
rect 212 2296 250 2324
rect 278 2296 316 2324
rect 344 2296 382 2324
rect 410 2296 448 2324
rect 476 2296 514 2324
rect 542 2296 580 2324
rect 608 2296 646 2324
rect 674 2296 712 2324
rect 740 2296 745 2324
rect -745 2258 745 2296
rect -745 2230 -740 2258
rect -712 2230 -674 2258
rect -646 2230 -608 2258
rect -580 2230 -542 2258
rect -514 2230 -476 2258
rect -448 2230 -410 2258
rect -382 2230 -344 2258
rect -316 2230 -278 2258
rect -250 2230 -212 2258
rect -184 2230 -146 2258
rect -118 2230 -80 2258
rect -52 2230 -14 2258
rect 14 2230 52 2258
rect 80 2230 118 2258
rect 146 2230 184 2258
rect 212 2230 250 2258
rect 278 2230 316 2258
rect 344 2230 382 2258
rect 410 2230 448 2258
rect 476 2230 514 2258
rect 542 2230 580 2258
rect 608 2230 646 2258
rect 674 2230 712 2258
rect 740 2230 745 2258
rect -745 2192 745 2230
rect -745 2164 -740 2192
rect -712 2164 -674 2192
rect -646 2164 -608 2192
rect -580 2164 -542 2192
rect -514 2164 -476 2192
rect -448 2164 -410 2192
rect -382 2164 -344 2192
rect -316 2164 -278 2192
rect -250 2164 -212 2192
rect -184 2164 -146 2192
rect -118 2164 -80 2192
rect -52 2164 -14 2192
rect 14 2164 52 2192
rect 80 2164 118 2192
rect 146 2164 184 2192
rect 212 2164 250 2192
rect 278 2164 316 2192
rect 344 2164 382 2192
rect 410 2164 448 2192
rect 476 2164 514 2192
rect 542 2164 580 2192
rect 608 2164 646 2192
rect 674 2164 712 2192
rect 740 2164 745 2192
rect -745 2126 745 2164
rect -745 2098 -740 2126
rect -712 2098 -674 2126
rect -646 2098 -608 2126
rect -580 2098 -542 2126
rect -514 2098 -476 2126
rect -448 2098 -410 2126
rect -382 2098 -344 2126
rect -316 2098 -278 2126
rect -250 2098 -212 2126
rect -184 2098 -146 2126
rect -118 2098 -80 2126
rect -52 2098 -14 2126
rect 14 2098 52 2126
rect 80 2098 118 2126
rect 146 2098 184 2126
rect 212 2098 250 2126
rect 278 2098 316 2126
rect 344 2098 382 2126
rect 410 2098 448 2126
rect 476 2098 514 2126
rect 542 2098 580 2126
rect 608 2098 646 2126
rect 674 2098 712 2126
rect 740 2098 745 2126
rect -745 2060 745 2098
rect -745 2032 -740 2060
rect -712 2032 -674 2060
rect -646 2032 -608 2060
rect -580 2032 -542 2060
rect -514 2032 -476 2060
rect -448 2032 -410 2060
rect -382 2032 -344 2060
rect -316 2032 -278 2060
rect -250 2032 -212 2060
rect -184 2032 -146 2060
rect -118 2032 -80 2060
rect -52 2032 -14 2060
rect 14 2032 52 2060
rect 80 2032 118 2060
rect 146 2032 184 2060
rect 212 2032 250 2060
rect 278 2032 316 2060
rect 344 2032 382 2060
rect 410 2032 448 2060
rect 476 2032 514 2060
rect 542 2032 580 2060
rect 608 2032 646 2060
rect 674 2032 712 2060
rect 740 2032 745 2060
rect -745 1994 745 2032
rect -745 1966 -740 1994
rect -712 1966 -674 1994
rect -646 1966 -608 1994
rect -580 1966 -542 1994
rect -514 1966 -476 1994
rect -448 1966 -410 1994
rect -382 1966 -344 1994
rect -316 1966 -278 1994
rect -250 1966 -212 1994
rect -184 1966 -146 1994
rect -118 1966 -80 1994
rect -52 1966 -14 1994
rect 14 1966 52 1994
rect 80 1966 118 1994
rect 146 1966 184 1994
rect 212 1966 250 1994
rect 278 1966 316 1994
rect 344 1966 382 1994
rect 410 1966 448 1994
rect 476 1966 514 1994
rect 542 1966 580 1994
rect 608 1966 646 1994
rect 674 1966 712 1994
rect 740 1966 745 1994
rect -745 1928 745 1966
rect -745 1900 -740 1928
rect -712 1900 -674 1928
rect -646 1900 -608 1928
rect -580 1900 -542 1928
rect -514 1900 -476 1928
rect -448 1900 -410 1928
rect -382 1900 -344 1928
rect -316 1900 -278 1928
rect -250 1900 -212 1928
rect -184 1900 -146 1928
rect -118 1900 -80 1928
rect -52 1900 -14 1928
rect 14 1900 52 1928
rect 80 1900 118 1928
rect 146 1900 184 1928
rect 212 1900 250 1928
rect 278 1900 316 1928
rect 344 1900 382 1928
rect 410 1900 448 1928
rect 476 1900 514 1928
rect 542 1900 580 1928
rect 608 1900 646 1928
rect 674 1900 712 1928
rect 740 1900 745 1928
rect -745 1862 745 1900
rect -745 1834 -740 1862
rect -712 1834 -674 1862
rect -646 1834 -608 1862
rect -580 1834 -542 1862
rect -514 1834 -476 1862
rect -448 1834 -410 1862
rect -382 1834 -344 1862
rect -316 1834 -278 1862
rect -250 1834 -212 1862
rect -184 1834 -146 1862
rect -118 1834 -80 1862
rect -52 1834 -14 1862
rect 14 1834 52 1862
rect 80 1834 118 1862
rect 146 1834 184 1862
rect 212 1834 250 1862
rect 278 1834 316 1862
rect 344 1834 382 1862
rect 410 1834 448 1862
rect 476 1834 514 1862
rect 542 1834 580 1862
rect 608 1834 646 1862
rect 674 1834 712 1862
rect 740 1834 745 1862
rect -745 1796 745 1834
rect -745 1768 -740 1796
rect -712 1768 -674 1796
rect -646 1768 -608 1796
rect -580 1768 -542 1796
rect -514 1768 -476 1796
rect -448 1768 -410 1796
rect -382 1768 -344 1796
rect -316 1768 -278 1796
rect -250 1768 -212 1796
rect -184 1768 -146 1796
rect -118 1768 -80 1796
rect -52 1768 -14 1796
rect 14 1768 52 1796
rect 80 1768 118 1796
rect 146 1768 184 1796
rect 212 1768 250 1796
rect 278 1768 316 1796
rect 344 1768 382 1796
rect 410 1768 448 1796
rect 476 1768 514 1796
rect 542 1768 580 1796
rect 608 1768 646 1796
rect 674 1768 712 1796
rect 740 1768 745 1796
rect -745 1730 745 1768
rect -745 1702 -740 1730
rect -712 1702 -674 1730
rect -646 1702 -608 1730
rect -580 1702 -542 1730
rect -514 1702 -476 1730
rect -448 1702 -410 1730
rect -382 1702 -344 1730
rect -316 1702 -278 1730
rect -250 1702 -212 1730
rect -184 1702 -146 1730
rect -118 1702 -80 1730
rect -52 1702 -14 1730
rect 14 1702 52 1730
rect 80 1702 118 1730
rect 146 1702 184 1730
rect 212 1702 250 1730
rect 278 1702 316 1730
rect 344 1702 382 1730
rect 410 1702 448 1730
rect 476 1702 514 1730
rect 542 1702 580 1730
rect 608 1702 646 1730
rect 674 1702 712 1730
rect 740 1702 745 1730
rect -745 1664 745 1702
rect -745 1636 -740 1664
rect -712 1636 -674 1664
rect -646 1636 -608 1664
rect -580 1636 -542 1664
rect -514 1636 -476 1664
rect -448 1636 -410 1664
rect -382 1636 -344 1664
rect -316 1636 -278 1664
rect -250 1636 -212 1664
rect -184 1636 -146 1664
rect -118 1636 -80 1664
rect -52 1636 -14 1664
rect 14 1636 52 1664
rect 80 1636 118 1664
rect 146 1636 184 1664
rect 212 1636 250 1664
rect 278 1636 316 1664
rect 344 1636 382 1664
rect 410 1636 448 1664
rect 476 1636 514 1664
rect 542 1636 580 1664
rect 608 1636 646 1664
rect 674 1636 712 1664
rect 740 1636 745 1664
rect -745 1598 745 1636
rect -745 1570 -740 1598
rect -712 1570 -674 1598
rect -646 1570 -608 1598
rect -580 1570 -542 1598
rect -514 1570 -476 1598
rect -448 1570 -410 1598
rect -382 1570 -344 1598
rect -316 1570 -278 1598
rect -250 1570 -212 1598
rect -184 1570 -146 1598
rect -118 1570 -80 1598
rect -52 1570 -14 1598
rect 14 1570 52 1598
rect 80 1570 118 1598
rect 146 1570 184 1598
rect 212 1570 250 1598
rect 278 1570 316 1598
rect 344 1570 382 1598
rect 410 1570 448 1598
rect 476 1570 514 1598
rect 542 1570 580 1598
rect 608 1570 646 1598
rect 674 1570 712 1598
rect 740 1570 745 1598
rect -745 1532 745 1570
rect -745 1504 -740 1532
rect -712 1504 -674 1532
rect -646 1504 -608 1532
rect -580 1504 -542 1532
rect -514 1504 -476 1532
rect -448 1504 -410 1532
rect -382 1504 -344 1532
rect -316 1504 -278 1532
rect -250 1504 -212 1532
rect -184 1504 -146 1532
rect -118 1504 -80 1532
rect -52 1504 -14 1532
rect 14 1504 52 1532
rect 80 1504 118 1532
rect 146 1504 184 1532
rect 212 1504 250 1532
rect 278 1504 316 1532
rect 344 1504 382 1532
rect 410 1504 448 1532
rect 476 1504 514 1532
rect 542 1504 580 1532
rect 608 1504 646 1532
rect 674 1504 712 1532
rect 740 1504 745 1532
rect -745 1466 745 1504
rect -745 1438 -740 1466
rect -712 1438 -674 1466
rect -646 1438 -608 1466
rect -580 1438 -542 1466
rect -514 1438 -476 1466
rect -448 1438 -410 1466
rect -382 1438 -344 1466
rect -316 1438 -278 1466
rect -250 1438 -212 1466
rect -184 1438 -146 1466
rect -118 1438 -80 1466
rect -52 1438 -14 1466
rect 14 1438 52 1466
rect 80 1438 118 1466
rect 146 1438 184 1466
rect 212 1438 250 1466
rect 278 1438 316 1466
rect 344 1438 382 1466
rect 410 1438 448 1466
rect 476 1438 514 1466
rect 542 1438 580 1466
rect 608 1438 646 1466
rect 674 1438 712 1466
rect 740 1438 745 1466
rect -745 1400 745 1438
rect -745 1372 -740 1400
rect -712 1372 -674 1400
rect -646 1372 -608 1400
rect -580 1372 -542 1400
rect -514 1372 -476 1400
rect -448 1372 -410 1400
rect -382 1372 -344 1400
rect -316 1372 -278 1400
rect -250 1372 -212 1400
rect -184 1372 -146 1400
rect -118 1372 -80 1400
rect -52 1372 -14 1400
rect 14 1372 52 1400
rect 80 1372 118 1400
rect 146 1372 184 1400
rect 212 1372 250 1400
rect 278 1372 316 1400
rect 344 1372 382 1400
rect 410 1372 448 1400
rect 476 1372 514 1400
rect 542 1372 580 1400
rect 608 1372 646 1400
rect 674 1372 712 1400
rect 740 1372 745 1400
rect -745 1334 745 1372
rect -745 1306 -740 1334
rect -712 1306 -674 1334
rect -646 1306 -608 1334
rect -580 1306 -542 1334
rect -514 1306 -476 1334
rect -448 1306 -410 1334
rect -382 1306 -344 1334
rect -316 1306 -278 1334
rect -250 1306 -212 1334
rect -184 1306 -146 1334
rect -118 1306 -80 1334
rect -52 1306 -14 1334
rect 14 1306 52 1334
rect 80 1306 118 1334
rect 146 1306 184 1334
rect 212 1306 250 1334
rect 278 1306 316 1334
rect 344 1306 382 1334
rect 410 1306 448 1334
rect 476 1306 514 1334
rect 542 1306 580 1334
rect 608 1306 646 1334
rect 674 1306 712 1334
rect 740 1306 745 1334
rect -745 1268 745 1306
rect -745 1240 -740 1268
rect -712 1240 -674 1268
rect -646 1240 -608 1268
rect -580 1240 -542 1268
rect -514 1240 -476 1268
rect -448 1240 -410 1268
rect -382 1240 -344 1268
rect -316 1240 -278 1268
rect -250 1240 -212 1268
rect -184 1240 -146 1268
rect -118 1240 -80 1268
rect -52 1240 -14 1268
rect 14 1240 52 1268
rect 80 1240 118 1268
rect 146 1240 184 1268
rect 212 1240 250 1268
rect 278 1240 316 1268
rect 344 1240 382 1268
rect 410 1240 448 1268
rect 476 1240 514 1268
rect 542 1240 580 1268
rect 608 1240 646 1268
rect 674 1240 712 1268
rect 740 1240 745 1268
rect -745 1202 745 1240
rect -745 1174 -740 1202
rect -712 1174 -674 1202
rect -646 1174 -608 1202
rect -580 1174 -542 1202
rect -514 1174 -476 1202
rect -448 1174 -410 1202
rect -382 1174 -344 1202
rect -316 1174 -278 1202
rect -250 1174 -212 1202
rect -184 1174 -146 1202
rect -118 1174 -80 1202
rect -52 1174 -14 1202
rect 14 1174 52 1202
rect 80 1174 118 1202
rect 146 1174 184 1202
rect 212 1174 250 1202
rect 278 1174 316 1202
rect 344 1174 382 1202
rect 410 1174 448 1202
rect 476 1174 514 1202
rect 542 1174 580 1202
rect 608 1174 646 1202
rect 674 1174 712 1202
rect 740 1174 745 1202
rect -745 1136 745 1174
rect -745 1108 -740 1136
rect -712 1108 -674 1136
rect -646 1108 -608 1136
rect -580 1108 -542 1136
rect -514 1108 -476 1136
rect -448 1108 -410 1136
rect -382 1108 -344 1136
rect -316 1108 -278 1136
rect -250 1108 -212 1136
rect -184 1108 -146 1136
rect -118 1108 -80 1136
rect -52 1108 -14 1136
rect 14 1108 52 1136
rect 80 1108 118 1136
rect 146 1108 184 1136
rect 212 1108 250 1136
rect 278 1108 316 1136
rect 344 1108 382 1136
rect 410 1108 448 1136
rect 476 1108 514 1136
rect 542 1108 580 1136
rect 608 1108 646 1136
rect 674 1108 712 1136
rect 740 1108 745 1136
rect -745 1070 745 1108
rect -745 1042 -740 1070
rect -712 1042 -674 1070
rect -646 1042 -608 1070
rect -580 1042 -542 1070
rect -514 1042 -476 1070
rect -448 1042 -410 1070
rect -382 1042 -344 1070
rect -316 1042 -278 1070
rect -250 1042 -212 1070
rect -184 1042 -146 1070
rect -118 1042 -80 1070
rect -52 1042 -14 1070
rect 14 1042 52 1070
rect 80 1042 118 1070
rect 146 1042 184 1070
rect 212 1042 250 1070
rect 278 1042 316 1070
rect 344 1042 382 1070
rect 410 1042 448 1070
rect 476 1042 514 1070
rect 542 1042 580 1070
rect 608 1042 646 1070
rect 674 1042 712 1070
rect 740 1042 745 1070
rect -745 1004 745 1042
rect -745 976 -740 1004
rect -712 976 -674 1004
rect -646 976 -608 1004
rect -580 976 -542 1004
rect -514 976 -476 1004
rect -448 976 -410 1004
rect -382 976 -344 1004
rect -316 976 -278 1004
rect -250 976 -212 1004
rect -184 976 -146 1004
rect -118 976 -80 1004
rect -52 976 -14 1004
rect 14 976 52 1004
rect 80 976 118 1004
rect 146 976 184 1004
rect 212 976 250 1004
rect 278 976 316 1004
rect 344 976 382 1004
rect 410 976 448 1004
rect 476 976 514 1004
rect 542 976 580 1004
rect 608 976 646 1004
rect 674 976 712 1004
rect 740 976 745 1004
rect -745 938 745 976
rect -745 910 -740 938
rect -712 910 -674 938
rect -646 910 -608 938
rect -580 910 -542 938
rect -514 910 -476 938
rect -448 910 -410 938
rect -382 910 -344 938
rect -316 910 -278 938
rect -250 910 -212 938
rect -184 910 -146 938
rect -118 910 -80 938
rect -52 910 -14 938
rect 14 910 52 938
rect 80 910 118 938
rect 146 910 184 938
rect 212 910 250 938
rect 278 910 316 938
rect 344 910 382 938
rect 410 910 448 938
rect 476 910 514 938
rect 542 910 580 938
rect 608 910 646 938
rect 674 910 712 938
rect 740 910 745 938
rect -745 872 745 910
rect -745 844 -740 872
rect -712 844 -674 872
rect -646 844 -608 872
rect -580 844 -542 872
rect -514 844 -476 872
rect -448 844 -410 872
rect -382 844 -344 872
rect -316 844 -278 872
rect -250 844 -212 872
rect -184 844 -146 872
rect -118 844 -80 872
rect -52 844 -14 872
rect 14 844 52 872
rect 80 844 118 872
rect 146 844 184 872
rect 212 844 250 872
rect 278 844 316 872
rect 344 844 382 872
rect 410 844 448 872
rect 476 844 514 872
rect 542 844 580 872
rect 608 844 646 872
rect 674 844 712 872
rect 740 844 745 872
rect -745 806 745 844
rect -745 778 -740 806
rect -712 778 -674 806
rect -646 778 -608 806
rect -580 778 -542 806
rect -514 778 -476 806
rect -448 778 -410 806
rect -382 778 -344 806
rect -316 778 -278 806
rect -250 778 -212 806
rect -184 778 -146 806
rect -118 778 -80 806
rect -52 778 -14 806
rect 14 778 52 806
rect 80 778 118 806
rect 146 778 184 806
rect 212 778 250 806
rect 278 778 316 806
rect 344 778 382 806
rect 410 778 448 806
rect 476 778 514 806
rect 542 778 580 806
rect 608 778 646 806
rect 674 778 712 806
rect 740 778 745 806
rect -745 740 745 778
rect -745 712 -740 740
rect -712 712 -674 740
rect -646 712 -608 740
rect -580 712 -542 740
rect -514 712 -476 740
rect -448 712 -410 740
rect -382 712 -344 740
rect -316 712 -278 740
rect -250 712 -212 740
rect -184 712 -146 740
rect -118 712 -80 740
rect -52 712 -14 740
rect 14 712 52 740
rect 80 712 118 740
rect 146 712 184 740
rect 212 712 250 740
rect 278 712 316 740
rect 344 712 382 740
rect 410 712 448 740
rect 476 712 514 740
rect 542 712 580 740
rect 608 712 646 740
rect 674 712 712 740
rect 740 712 745 740
rect -745 674 745 712
rect -745 646 -740 674
rect -712 646 -674 674
rect -646 646 -608 674
rect -580 646 -542 674
rect -514 646 -476 674
rect -448 646 -410 674
rect -382 646 -344 674
rect -316 646 -278 674
rect -250 646 -212 674
rect -184 646 -146 674
rect -118 646 -80 674
rect -52 646 -14 674
rect 14 646 52 674
rect 80 646 118 674
rect 146 646 184 674
rect 212 646 250 674
rect 278 646 316 674
rect 344 646 382 674
rect 410 646 448 674
rect 476 646 514 674
rect 542 646 580 674
rect 608 646 646 674
rect 674 646 712 674
rect 740 646 745 674
rect -745 608 745 646
rect -745 580 -740 608
rect -712 580 -674 608
rect -646 580 -608 608
rect -580 580 -542 608
rect -514 580 -476 608
rect -448 580 -410 608
rect -382 580 -344 608
rect -316 580 -278 608
rect -250 580 -212 608
rect -184 580 -146 608
rect -118 580 -80 608
rect -52 580 -14 608
rect 14 580 52 608
rect 80 580 118 608
rect 146 580 184 608
rect 212 580 250 608
rect 278 580 316 608
rect 344 580 382 608
rect 410 580 448 608
rect 476 580 514 608
rect 542 580 580 608
rect 608 580 646 608
rect 674 580 712 608
rect 740 580 745 608
rect -745 542 745 580
rect -745 514 -740 542
rect -712 514 -674 542
rect -646 514 -608 542
rect -580 514 -542 542
rect -514 514 -476 542
rect -448 514 -410 542
rect -382 514 -344 542
rect -316 514 -278 542
rect -250 514 -212 542
rect -184 514 -146 542
rect -118 514 -80 542
rect -52 514 -14 542
rect 14 514 52 542
rect 80 514 118 542
rect 146 514 184 542
rect 212 514 250 542
rect 278 514 316 542
rect 344 514 382 542
rect 410 514 448 542
rect 476 514 514 542
rect 542 514 580 542
rect 608 514 646 542
rect 674 514 712 542
rect 740 514 745 542
rect -745 476 745 514
rect -745 448 -740 476
rect -712 448 -674 476
rect -646 448 -608 476
rect -580 448 -542 476
rect -514 448 -476 476
rect -448 448 -410 476
rect -382 448 -344 476
rect -316 448 -278 476
rect -250 448 -212 476
rect -184 448 -146 476
rect -118 448 -80 476
rect -52 448 -14 476
rect 14 448 52 476
rect 80 448 118 476
rect 146 448 184 476
rect 212 448 250 476
rect 278 448 316 476
rect 344 448 382 476
rect 410 448 448 476
rect 476 448 514 476
rect 542 448 580 476
rect 608 448 646 476
rect 674 448 712 476
rect 740 448 745 476
rect -745 410 745 448
rect -745 382 -740 410
rect -712 382 -674 410
rect -646 382 -608 410
rect -580 382 -542 410
rect -514 382 -476 410
rect -448 382 -410 410
rect -382 382 -344 410
rect -316 382 -278 410
rect -250 382 -212 410
rect -184 382 -146 410
rect -118 382 -80 410
rect -52 382 -14 410
rect 14 382 52 410
rect 80 382 118 410
rect 146 382 184 410
rect 212 382 250 410
rect 278 382 316 410
rect 344 382 382 410
rect 410 382 448 410
rect 476 382 514 410
rect 542 382 580 410
rect 608 382 646 410
rect 674 382 712 410
rect 740 382 745 410
rect -745 344 745 382
rect -745 316 -740 344
rect -712 316 -674 344
rect -646 316 -608 344
rect -580 316 -542 344
rect -514 316 -476 344
rect -448 316 -410 344
rect -382 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 382 344
rect 410 316 448 344
rect 476 316 514 344
rect 542 316 580 344
rect 608 316 646 344
rect 674 316 712 344
rect 740 316 745 344
rect -745 278 745 316
rect -745 250 -740 278
rect -712 250 -674 278
rect -646 250 -608 278
rect -580 250 -542 278
rect -514 250 -476 278
rect -448 250 -410 278
rect -382 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 382 278
rect 410 250 448 278
rect 476 250 514 278
rect 542 250 580 278
rect 608 250 646 278
rect 674 250 712 278
rect 740 250 745 278
rect -745 212 745 250
rect -745 184 -740 212
rect -712 184 -674 212
rect -646 184 -608 212
rect -580 184 -542 212
rect -514 184 -476 212
rect -448 184 -410 212
rect -382 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 382 212
rect 410 184 448 212
rect 476 184 514 212
rect 542 184 580 212
rect 608 184 646 212
rect 674 184 712 212
rect 740 184 745 212
rect -745 146 745 184
rect -745 118 -740 146
rect -712 118 -674 146
rect -646 118 -608 146
rect -580 118 -542 146
rect -514 118 -476 146
rect -448 118 -410 146
rect -382 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 382 146
rect 410 118 448 146
rect 476 118 514 146
rect 542 118 580 146
rect 608 118 646 146
rect 674 118 712 146
rect 740 118 745 146
rect -745 80 745 118
rect -745 52 -740 80
rect -712 52 -674 80
rect -646 52 -608 80
rect -580 52 -542 80
rect -514 52 -476 80
rect -448 52 -410 80
rect -382 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 382 80
rect 410 52 448 80
rect 476 52 514 80
rect 542 52 580 80
rect 608 52 646 80
rect 674 52 712 80
rect 740 52 745 80
rect -745 14 745 52
rect -745 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 382 14
rect 410 -14 448 14
rect 476 -14 514 14
rect 542 -14 580 14
rect 608 -14 646 14
rect 674 -14 712 14
rect 740 -14 745 14
rect -745 -52 745 -14
rect -745 -80 -740 -52
rect -712 -80 -674 -52
rect -646 -80 -608 -52
rect -580 -80 -542 -52
rect -514 -80 -476 -52
rect -448 -80 -410 -52
rect -382 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 382 -52
rect 410 -80 448 -52
rect 476 -80 514 -52
rect 542 -80 580 -52
rect 608 -80 646 -52
rect 674 -80 712 -52
rect 740 -80 745 -52
rect -745 -118 745 -80
rect -745 -146 -740 -118
rect -712 -146 -674 -118
rect -646 -146 -608 -118
rect -580 -146 -542 -118
rect -514 -146 -476 -118
rect -448 -146 -410 -118
rect -382 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 382 -118
rect 410 -146 448 -118
rect 476 -146 514 -118
rect 542 -146 580 -118
rect 608 -146 646 -118
rect 674 -146 712 -118
rect 740 -146 745 -118
rect -745 -184 745 -146
rect -745 -212 -740 -184
rect -712 -212 -674 -184
rect -646 -212 -608 -184
rect -580 -212 -542 -184
rect -514 -212 -476 -184
rect -448 -212 -410 -184
rect -382 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 382 -184
rect 410 -212 448 -184
rect 476 -212 514 -184
rect 542 -212 580 -184
rect 608 -212 646 -184
rect 674 -212 712 -184
rect 740 -212 745 -184
rect -745 -250 745 -212
rect -745 -278 -740 -250
rect -712 -278 -674 -250
rect -646 -278 -608 -250
rect -580 -278 -542 -250
rect -514 -278 -476 -250
rect -448 -278 -410 -250
rect -382 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 382 -250
rect 410 -278 448 -250
rect 476 -278 514 -250
rect 542 -278 580 -250
rect 608 -278 646 -250
rect 674 -278 712 -250
rect 740 -278 745 -250
rect -745 -316 745 -278
rect -745 -344 -740 -316
rect -712 -344 -674 -316
rect -646 -344 -608 -316
rect -580 -344 -542 -316
rect -514 -344 -476 -316
rect -448 -344 -410 -316
rect -382 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 382 -316
rect 410 -344 448 -316
rect 476 -344 514 -316
rect 542 -344 580 -316
rect 608 -344 646 -316
rect 674 -344 712 -316
rect 740 -344 745 -316
rect -745 -382 745 -344
rect -745 -410 -740 -382
rect -712 -410 -674 -382
rect -646 -410 -608 -382
rect -580 -410 -542 -382
rect -514 -410 -476 -382
rect -448 -410 -410 -382
rect -382 -410 -344 -382
rect -316 -410 -278 -382
rect -250 -410 -212 -382
rect -184 -410 -146 -382
rect -118 -410 -80 -382
rect -52 -410 -14 -382
rect 14 -410 52 -382
rect 80 -410 118 -382
rect 146 -410 184 -382
rect 212 -410 250 -382
rect 278 -410 316 -382
rect 344 -410 382 -382
rect 410 -410 448 -382
rect 476 -410 514 -382
rect 542 -410 580 -382
rect 608 -410 646 -382
rect 674 -410 712 -382
rect 740 -410 745 -382
rect -745 -448 745 -410
rect -745 -476 -740 -448
rect -712 -476 -674 -448
rect -646 -476 -608 -448
rect -580 -476 -542 -448
rect -514 -476 -476 -448
rect -448 -476 -410 -448
rect -382 -476 -344 -448
rect -316 -476 -278 -448
rect -250 -476 -212 -448
rect -184 -476 -146 -448
rect -118 -476 -80 -448
rect -52 -476 -14 -448
rect 14 -476 52 -448
rect 80 -476 118 -448
rect 146 -476 184 -448
rect 212 -476 250 -448
rect 278 -476 316 -448
rect 344 -476 382 -448
rect 410 -476 448 -448
rect 476 -476 514 -448
rect 542 -476 580 -448
rect 608 -476 646 -448
rect 674 -476 712 -448
rect 740 -476 745 -448
rect -745 -514 745 -476
rect -745 -542 -740 -514
rect -712 -542 -674 -514
rect -646 -542 -608 -514
rect -580 -542 -542 -514
rect -514 -542 -476 -514
rect -448 -542 -410 -514
rect -382 -542 -344 -514
rect -316 -542 -278 -514
rect -250 -542 -212 -514
rect -184 -542 -146 -514
rect -118 -542 -80 -514
rect -52 -542 -14 -514
rect 14 -542 52 -514
rect 80 -542 118 -514
rect 146 -542 184 -514
rect 212 -542 250 -514
rect 278 -542 316 -514
rect 344 -542 382 -514
rect 410 -542 448 -514
rect 476 -542 514 -514
rect 542 -542 580 -514
rect 608 -542 646 -514
rect 674 -542 712 -514
rect 740 -542 745 -514
rect -745 -580 745 -542
rect -745 -608 -740 -580
rect -712 -608 -674 -580
rect -646 -608 -608 -580
rect -580 -608 -542 -580
rect -514 -608 -476 -580
rect -448 -608 -410 -580
rect -382 -608 -344 -580
rect -316 -608 -278 -580
rect -250 -608 -212 -580
rect -184 -608 -146 -580
rect -118 -608 -80 -580
rect -52 -608 -14 -580
rect 14 -608 52 -580
rect 80 -608 118 -580
rect 146 -608 184 -580
rect 212 -608 250 -580
rect 278 -608 316 -580
rect 344 -608 382 -580
rect 410 -608 448 -580
rect 476 -608 514 -580
rect 542 -608 580 -580
rect 608 -608 646 -580
rect 674 -608 712 -580
rect 740 -608 745 -580
rect -745 -646 745 -608
rect -745 -674 -740 -646
rect -712 -674 -674 -646
rect -646 -674 -608 -646
rect -580 -674 -542 -646
rect -514 -674 -476 -646
rect -448 -674 -410 -646
rect -382 -674 -344 -646
rect -316 -674 -278 -646
rect -250 -674 -212 -646
rect -184 -674 -146 -646
rect -118 -674 -80 -646
rect -52 -674 -14 -646
rect 14 -674 52 -646
rect 80 -674 118 -646
rect 146 -674 184 -646
rect 212 -674 250 -646
rect 278 -674 316 -646
rect 344 -674 382 -646
rect 410 -674 448 -646
rect 476 -674 514 -646
rect 542 -674 580 -646
rect 608 -674 646 -646
rect 674 -674 712 -646
rect 740 -674 745 -646
rect -745 -712 745 -674
rect -745 -740 -740 -712
rect -712 -740 -674 -712
rect -646 -740 -608 -712
rect -580 -740 -542 -712
rect -514 -740 -476 -712
rect -448 -740 -410 -712
rect -382 -740 -344 -712
rect -316 -740 -278 -712
rect -250 -740 -212 -712
rect -184 -740 -146 -712
rect -118 -740 -80 -712
rect -52 -740 -14 -712
rect 14 -740 52 -712
rect 80 -740 118 -712
rect 146 -740 184 -712
rect 212 -740 250 -712
rect 278 -740 316 -712
rect 344 -740 382 -712
rect 410 -740 448 -712
rect 476 -740 514 -712
rect 542 -740 580 -712
rect 608 -740 646 -712
rect 674 -740 712 -712
rect 740 -740 745 -712
rect -745 -778 745 -740
rect -745 -806 -740 -778
rect -712 -806 -674 -778
rect -646 -806 -608 -778
rect -580 -806 -542 -778
rect -514 -806 -476 -778
rect -448 -806 -410 -778
rect -382 -806 -344 -778
rect -316 -806 -278 -778
rect -250 -806 -212 -778
rect -184 -806 -146 -778
rect -118 -806 -80 -778
rect -52 -806 -14 -778
rect 14 -806 52 -778
rect 80 -806 118 -778
rect 146 -806 184 -778
rect 212 -806 250 -778
rect 278 -806 316 -778
rect 344 -806 382 -778
rect 410 -806 448 -778
rect 476 -806 514 -778
rect 542 -806 580 -778
rect 608 -806 646 -778
rect 674 -806 712 -778
rect 740 -806 745 -778
rect -745 -844 745 -806
rect -745 -872 -740 -844
rect -712 -872 -674 -844
rect -646 -872 -608 -844
rect -580 -872 -542 -844
rect -514 -872 -476 -844
rect -448 -872 -410 -844
rect -382 -872 -344 -844
rect -316 -872 -278 -844
rect -250 -872 -212 -844
rect -184 -872 -146 -844
rect -118 -872 -80 -844
rect -52 -872 -14 -844
rect 14 -872 52 -844
rect 80 -872 118 -844
rect 146 -872 184 -844
rect 212 -872 250 -844
rect 278 -872 316 -844
rect 344 -872 382 -844
rect 410 -872 448 -844
rect 476 -872 514 -844
rect 542 -872 580 -844
rect 608 -872 646 -844
rect 674 -872 712 -844
rect 740 -872 745 -844
rect -745 -910 745 -872
rect -745 -938 -740 -910
rect -712 -938 -674 -910
rect -646 -938 -608 -910
rect -580 -938 -542 -910
rect -514 -938 -476 -910
rect -448 -938 -410 -910
rect -382 -938 -344 -910
rect -316 -938 -278 -910
rect -250 -938 -212 -910
rect -184 -938 -146 -910
rect -118 -938 -80 -910
rect -52 -938 -14 -910
rect 14 -938 52 -910
rect 80 -938 118 -910
rect 146 -938 184 -910
rect 212 -938 250 -910
rect 278 -938 316 -910
rect 344 -938 382 -910
rect 410 -938 448 -910
rect 476 -938 514 -910
rect 542 -938 580 -910
rect 608 -938 646 -910
rect 674 -938 712 -910
rect 740 -938 745 -910
rect -745 -976 745 -938
rect -745 -1004 -740 -976
rect -712 -1004 -674 -976
rect -646 -1004 -608 -976
rect -580 -1004 -542 -976
rect -514 -1004 -476 -976
rect -448 -1004 -410 -976
rect -382 -1004 -344 -976
rect -316 -1004 -278 -976
rect -250 -1004 -212 -976
rect -184 -1004 -146 -976
rect -118 -1004 -80 -976
rect -52 -1004 -14 -976
rect 14 -1004 52 -976
rect 80 -1004 118 -976
rect 146 -1004 184 -976
rect 212 -1004 250 -976
rect 278 -1004 316 -976
rect 344 -1004 382 -976
rect 410 -1004 448 -976
rect 476 -1004 514 -976
rect 542 -1004 580 -976
rect 608 -1004 646 -976
rect 674 -1004 712 -976
rect 740 -1004 745 -976
rect -745 -1042 745 -1004
rect -745 -1070 -740 -1042
rect -712 -1070 -674 -1042
rect -646 -1070 -608 -1042
rect -580 -1070 -542 -1042
rect -514 -1070 -476 -1042
rect -448 -1070 -410 -1042
rect -382 -1070 -344 -1042
rect -316 -1070 -278 -1042
rect -250 -1070 -212 -1042
rect -184 -1070 -146 -1042
rect -118 -1070 -80 -1042
rect -52 -1070 -14 -1042
rect 14 -1070 52 -1042
rect 80 -1070 118 -1042
rect 146 -1070 184 -1042
rect 212 -1070 250 -1042
rect 278 -1070 316 -1042
rect 344 -1070 382 -1042
rect 410 -1070 448 -1042
rect 476 -1070 514 -1042
rect 542 -1070 580 -1042
rect 608 -1070 646 -1042
rect 674 -1070 712 -1042
rect 740 -1070 745 -1042
rect -745 -1108 745 -1070
rect -745 -1136 -740 -1108
rect -712 -1136 -674 -1108
rect -646 -1136 -608 -1108
rect -580 -1136 -542 -1108
rect -514 -1136 -476 -1108
rect -448 -1136 -410 -1108
rect -382 -1136 -344 -1108
rect -316 -1136 -278 -1108
rect -250 -1136 -212 -1108
rect -184 -1136 -146 -1108
rect -118 -1136 -80 -1108
rect -52 -1136 -14 -1108
rect 14 -1136 52 -1108
rect 80 -1136 118 -1108
rect 146 -1136 184 -1108
rect 212 -1136 250 -1108
rect 278 -1136 316 -1108
rect 344 -1136 382 -1108
rect 410 -1136 448 -1108
rect 476 -1136 514 -1108
rect 542 -1136 580 -1108
rect 608 -1136 646 -1108
rect 674 -1136 712 -1108
rect 740 -1136 745 -1108
rect -745 -1174 745 -1136
rect -745 -1202 -740 -1174
rect -712 -1202 -674 -1174
rect -646 -1202 -608 -1174
rect -580 -1202 -542 -1174
rect -514 -1202 -476 -1174
rect -448 -1202 -410 -1174
rect -382 -1202 -344 -1174
rect -316 -1202 -278 -1174
rect -250 -1202 -212 -1174
rect -184 -1202 -146 -1174
rect -118 -1202 -80 -1174
rect -52 -1202 -14 -1174
rect 14 -1202 52 -1174
rect 80 -1202 118 -1174
rect 146 -1202 184 -1174
rect 212 -1202 250 -1174
rect 278 -1202 316 -1174
rect 344 -1202 382 -1174
rect 410 -1202 448 -1174
rect 476 -1202 514 -1174
rect 542 -1202 580 -1174
rect 608 -1202 646 -1174
rect 674 -1202 712 -1174
rect 740 -1202 745 -1174
rect -745 -1240 745 -1202
rect -745 -1268 -740 -1240
rect -712 -1268 -674 -1240
rect -646 -1268 -608 -1240
rect -580 -1268 -542 -1240
rect -514 -1268 -476 -1240
rect -448 -1268 -410 -1240
rect -382 -1268 -344 -1240
rect -316 -1268 -278 -1240
rect -250 -1268 -212 -1240
rect -184 -1268 -146 -1240
rect -118 -1268 -80 -1240
rect -52 -1268 -14 -1240
rect 14 -1268 52 -1240
rect 80 -1268 118 -1240
rect 146 -1268 184 -1240
rect 212 -1268 250 -1240
rect 278 -1268 316 -1240
rect 344 -1268 382 -1240
rect 410 -1268 448 -1240
rect 476 -1268 514 -1240
rect 542 -1268 580 -1240
rect 608 -1268 646 -1240
rect 674 -1268 712 -1240
rect 740 -1268 745 -1240
rect -745 -1306 745 -1268
rect -745 -1334 -740 -1306
rect -712 -1334 -674 -1306
rect -646 -1334 -608 -1306
rect -580 -1334 -542 -1306
rect -514 -1334 -476 -1306
rect -448 -1334 -410 -1306
rect -382 -1334 -344 -1306
rect -316 -1334 -278 -1306
rect -250 -1334 -212 -1306
rect -184 -1334 -146 -1306
rect -118 -1334 -80 -1306
rect -52 -1334 -14 -1306
rect 14 -1334 52 -1306
rect 80 -1334 118 -1306
rect 146 -1334 184 -1306
rect 212 -1334 250 -1306
rect 278 -1334 316 -1306
rect 344 -1334 382 -1306
rect 410 -1334 448 -1306
rect 476 -1334 514 -1306
rect 542 -1334 580 -1306
rect 608 -1334 646 -1306
rect 674 -1334 712 -1306
rect 740 -1334 745 -1306
rect -745 -1372 745 -1334
rect -745 -1400 -740 -1372
rect -712 -1400 -674 -1372
rect -646 -1400 -608 -1372
rect -580 -1400 -542 -1372
rect -514 -1400 -476 -1372
rect -448 -1400 -410 -1372
rect -382 -1400 -344 -1372
rect -316 -1400 -278 -1372
rect -250 -1400 -212 -1372
rect -184 -1400 -146 -1372
rect -118 -1400 -80 -1372
rect -52 -1400 -14 -1372
rect 14 -1400 52 -1372
rect 80 -1400 118 -1372
rect 146 -1400 184 -1372
rect 212 -1400 250 -1372
rect 278 -1400 316 -1372
rect 344 -1400 382 -1372
rect 410 -1400 448 -1372
rect 476 -1400 514 -1372
rect 542 -1400 580 -1372
rect 608 -1400 646 -1372
rect 674 -1400 712 -1372
rect 740 -1400 745 -1372
rect -745 -1438 745 -1400
rect -745 -1466 -740 -1438
rect -712 -1466 -674 -1438
rect -646 -1466 -608 -1438
rect -580 -1466 -542 -1438
rect -514 -1466 -476 -1438
rect -448 -1466 -410 -1438
rect -382 -1466 -344 -1438
rect -316 -1466 -278 -1438
rect -250 -1466 -212 -1438
rect -184 -1466 -146 -1438
rect -118 -1466 -80 -1438
rect -52 -1466 -14 -1438
rect 14 -1466 52 -1438
rect 80 -1466 118 -1438
rect 146 -1466 184 -1438
rect 212 -1466 250 -1438
rect 278 -1466 316 -1438
rect 344 -1466 382 -1438
rect 410 -1466 448 -1438
rect 476 -1466 514 -1438
rect 542 -1466 580 -1438
rect 608 -1466 646 -1438
rect 674 -1466 712 -1438
rect 740 -1466 745 -1438
rect -745 -1504 745 -1466
rect -745 -1532 -740 -1504
rect -712 -1532 -674 -1504
rect -646 -1532 -608 -1504
rect -580 -1532 -542 -1504
rect -514 -1532 -476 -1504
rect -448 -1532 -410 -1504
rect -382 -1532 -344 -1504
rect -316 -1532 -278 -1504
rect -250 -1532 -212 -1504
rect -184 -1532 -146 -1504
rect -118 -1532 -80 -1504
rect -52 -1532 -14 -1504
rect 14 -1532 52 -1504
rect 80 -1532 118 -1504
rect 146 -1532 184 -1504
rect 212 -1532 250 -1504
rect 278 -1532 316 -1504
rect 344 -1532 382 -1504
rect 410 -1532 448 -1504
rect 476 -1532 514 -1504
rect 542 -1532 580 -1504
rect 608 -1532 646 -1504
rect 674 -1532 712 -1504
rect 740 -1532 745 -1504
rect -745 -1570 745 -1532
rect -745 -1598 -740 -1570
rect -712 -1598 -674 -1570
rect -646 -1598 -608 -1570
rect -580 -1598 -542 -1570
rect -514 -1598 -476 -1570
rect -448 -1598 -410 -1570
rect -382 -1598 -344 -1570
rect -316 -1598 -278 -1570
rect -250 -1598 -212 -1570
rect -184 -1598 -146 -1570
rect -118 -1598 -80 -1570
rect -52 -1598 -14 -1570
rect 14 -1598 52 -1570
rect 80 -1598 118 -1570
rect 146 -1598 184 -1570
rect 212 -1598 250 -1570
rect 278 -1598 316 -1570
rect 344 -1598 382 -1570
rect 410 -1598 448 -1570
rect 476 -1598 514 -1570
rect 542 -1598 580 -1570
rect 608 -1598 646 -1570
rect 674 -1598 712 -1570
rect 740 -1598 745 -1570
rect -745 -1636 745 -1598
rect -745 -1664 -740 -1636
rect -712 -1664 -674 -1636
rect -646 -1664 -608 -1636
rect -580 -1664 -542 -1636
rect -514 -1664 -476 -1636
rect -448 -1664 -410 -1636
rect -382 -1664 -344 -1636
rect -316 -1664 -278 -1636
rect -250 -1664 -212 -1636
rect -184 -1664 -146 -1636
rect -118 -1664 -80 -1636
rect -52 -1664 -14 -1636
rect 14 -1664 52 -1636
rect 80 -1664 118 -1636
rect 146 -1664 184 -1636
rect 212 -1664 250 -1636
rect 278 -1664 316 -1636
rect 344 -1664 382 -1636
rect 410 -1664 448 -1636
rect 476 -1664 514 -1636
rect 542 -1664 580 -1636
rect 608 -1664 646 -1636
rect 674 -1664 712 -1636
rect 740 -1664 745 -1636
rect -745 -1702 745 -1664
rect -745 -1730 -740 -1702
rect -712 -1730 -674 -1702
rect -646 -1730 -608 -1702
rect -580 -1730 -542 -1702
rect -514 -1730 -476 -1702
rect -448 -1730 -410 -1702
rect -382 -1730 -344 -1702
rect -316 -1730 -278 -1702
rect -250 -1730 -212 -1702
rect -184 -1730 -146 -1702
rect -118 -1730 -80 -1702
rect -52 -1730 -14 -1702
rect 14 -1730 52 -1702
rect 80 -1730 118 -1702
rect 146 -1730 184 -1702
rect 212 -1730 250 -1702
rect 278 -1730 316 -1702
rect 344 -1730 382 -1702
rect 410 -1730 448 -1702
rect 476 -1730 514 -1702
rect 542 -1730 580 -1702
rect 608 -1730 646 -1702
rect 674 -1730 712 -1702
rect 740 -1730 745 -1702
rect -745 -1768 745 -1730
rect -745 -1796 -740 -1768
rect -712 -1796 -674 -1768
rect -646 -1796 -608 -1768
rect -580 -1796 -542 -1768
rect -514 -1796 -476 -1768
rect -448 -1796 -410 -1768
rect -382 -1796 -344 -1768
rect -316 -1796 -278 -1768
rect -250 -1796 -212 -1768
rect -184 -1796 -146 -1768
rect -118 -1796 -80 -1768
rect -52 -1796 -14 -1768
rect 14 -1796 52 -1768
rect 80 -1796 118 -1768
rect 146 -1796 184 -1768
rect 212 -1796 250 -1768
rect 278 -1796 316 -1768
rect 344 -1796 382 -1768
rect 410 -1796 448 -1768
rect 476 -1796 514 -1768
rect 542 -1796 580 -1768
rect 608 -1796 646 -1768
rect 674 -1796 712 -1768
rect 740 -1796 745 -1768
rect -745 -1834 745 -1796
rect -745 -1862 -740 -1834
rect -712 -1862 -674 -1834
rect -646 -1862 -608 -1834
rect -580 -1862 -542 -1834
rect -514 -1862 -476 -1834
rect -448 -1862 -410 -1834
rect -382 -1862 -344 -1834
rect -316 -1862 -278 -1834
rect -250 -1862 -212 -1834
rect -184 -1862 -146 -1834
rect -118 -1862 -80 -1834
rect -52 -1862 -14 -1834
rect 14 -1862 52 -1834
rect 80 -1862 118 -1834
rect 146 -1862 184 -1834
rect 212 -1862 250 -1834
rect 278 -1862 316 -1834
rect 344 -1862 382 -1834
rect 410 -1862 448 -1834
rect 476 -1862 514 -1834
rect 542 -1862 580 -1834
rect 608 -1862 646 -1834
rect 674 -1862 712 -1834
rect 740 -1862 745 -1834
rect -745 -1900 745 -1862
rect -745 -1928 -740 -1900
rect -712 -1928 -674 -1900
rect -646 -1928 -608 -1900
rect -580 -1928 -542 -1900
rect -514 -1928 -476 -1900
rect -448 -1928 -410 -1900
rect -382 -1928 -344 -1900
rect -316 -1928 -278 -1900
rect -250 -1928 -212 -1900
rect -184 -1928 -146 -1900
rect -118 -1928 -80 -1900
rect -52 -1928 -14 -1900
rect 14 -1928 52 -1900
rect 80 -1928 118 -1900
rect 146 -1928 184 -1900
rect 212 -1928 250 -1900
rect 278 -1928 316 -1900
rect 344 -1928 382 -1900
rect 410 -1928 448 -1900
rect 476 -1928 514 -1900
rect 542 -1928 580 -1900
rect 608 -1928 646 -1900
rect 674 -1928 712 -1900
rect 740 -1928 745 -1900
rect -745 -1966 745 -1928
rect -745 -1994 -740 -1966
rect -712 -1994 -674 -1966
rect -646 -1994 -608 -1966
rect -580 -1994 -542 -1966
rect -514 -1994 -476 -1966
rect -448 -1994 -410 -1966
rect -382 -1994 -344 -1966
rect -316 -1994 -278 -1966
rect -250 -1994 -212 -1966
rect -184 -1994 -146 -1966
rect -118 -1994 -80 -1966
rect -52 -1994 -14 -1966
rect 14 -1994 52 -1966
rect 80 -1994 118 -1966
rect 146 -1994 184 -1966
rect 212 -1994 250 -1966
rect 278 -1994 316 -1966
rect 344 -1994 382 -1966
rect 410 -1994 448 -1966
rect 476 -1994 514 -1966
rect 542 -1994 580 -1966
rect 608 -1994 646 -1966
rect 674 -1994 712 -1966
rect 740 -1994 745 -1966
rect -745 -2032 745 -1994
rect -745 -2060 -740 -2032
rect -712 -2060 -674 -2032
rect -646 -2060 -608 -2032
rect -580 -2060 -542 -2032
rect -514 -2060 -476 -2032
rect -448 -2060 -410 -2032
rect -382 -2060 -344 -2032
rect -316 -2060 -278 -2032
rect -250 -2060 -212 -2032
rect -184 -2060 -146 -2032
rect -118 -2060 -80 -2032
rect -52 -2060 -14 -2032
rect 14 -2060 52 -2032
rect 80 -2060 118 -2032
rect 146 -2060 184 -2032
rect 212 -2060 250 -2032
rect 278 -2060 316 -2032
rect 344 -2060 382 -2032
rect 410 -2060 448 -2032
rect 476 -2060 514 -2032
rect 542 -2060 580 -2032
rect 608 -2060 646 -2032
rect 674 -2060 712 -2032
rect 740 -2060 745 -2032
rect -745 -2098 745 -2060
rect -745 -2126 -740 -2098
rect -712 -2126 -674 -2098
rect -646 -2126 -608 -2098
rect -580 -2126 -542 -2098
rect -514 -2126 -476 -2098
rect -448 -2126 -410 -2098
rect -382 -2126 -344 -2098
rect -316 -2126 -278 -2098
rect -250 -2126 -212 -2098
rect -184 -2126 -146 -2098
rect -118 -2126 -80 -2098
rect -52 -2126 -14 -2098
rect 14 -2126 52 -2098
rect 80 -2126 118 -2098
rect 146 -2126 184 -2098
rect 212 -2126 250 -2098
rect 278 -2126 316 -2098
rect 344 -2126 382 -2098
rect 410 -2126 448 -2098
rect 476 -2126 514 -2098
rect 542 -2126 580 -2098
rect 608 -2126 646 -2098
rect 674 -2126 712 -2098
rect 740 -2126 745 -2098
rect -745 -2164 745 -2126
rect -745 -2192 -740 -2164
rect -712 -2192 -674 -2164
rect -646 -2192 -608 -2164
rect -580 -2192 -542 -2164
rect -514 -2192 -476 -2164
rect -448 -2192 -410 -2164
rect -382 -2192 -344 -2164
rect -316 -2192 -278 -2164
rect -250 -2192 -212 -2164
rect -184 -2192 -146 -2164
rect -118 -2192 -80 -2164
rect -52 -2192 -14 -2164
rect 14 -2192 52 -2164
rect 80 -2192 118 -2164
rect 146 -2192 184 -2164
rect 212 -2192 250 -2164
rect 278 -2192 316 -2164
rect 344 -2192 382 -2164
rect 410 -2192 448 -2164
rect 476 -2192 514 -2164
rect 542 -2192 580 -2164
rect 608 -2192 646 -2164
rect 674 -2192 712 -2164
rect 740 -2192 745 -2164
rect -745 -2230 745 -2192
rect -745 -2258 -740 -2230
rect -712 -2258 -674 -2230
rect -646 -2258 -608 -2230
rect -580 -2258 -542 -2230
rect -514 -2258 -476 -2230
rect -448 -2258 -410 -2230
rect -382 -2258 -344 -2230
rect -316 -2258 -278 -2230
rect -250 -2258 -212 -2230
rect -184 -2258 -146 -2230
rect -118 -2258 -80 -2230
rect -52 -2258 -14 -2230
rect 14 -2258 52 -2230
rect 80 -2258 118 -2230
rect 146 -2258 184 -2230
rect 212 -2258 250 -2230
rect 278 -2258 316 -2230
rect 344 -2258 382 -2230
rect 410 -2258 448 -2230
rect 476 -2258 514 -2230
rect 542 -2258 580 -2230
rect 608 -2258 646 -2230
rect 674 -2258 712 -2230
rect 740 -2258 745 -2230
rect -745 -2296 745 -2258
rect -745 -2324 -740 -2296
rect -712 -2324 -674 -2296
rect -646 -2324 -608 -2296
rect -580 -2324 -542 -2296
rect -514 -2324 -476 -2296
rect -448 -2324 -410 -2296
rect -382 -2324 -344 -2296
rect -316 -2324 -278 -2296
rect -250 -2324 -212 -2296
rect -184 -2324 -146 -2296
rect -118 -2324 -80 -2296
rect -52 -2324 -14 -2296
rect 14 -2324 52 -2296
rect 80 -2324 118 -2296
rect 146 -2324 184 -2296
rect 212 -2324 250 -2296
rect 278 -2324 316 -2296
rect 344 -2324 382 -2296
rect 410 -2324 448 -2296
rect 476 -2324 514 -2296
rect 542 -2324 580 -2296
rect 608 -2324 646 -2296
rect 674 -2324 712 -2296
rect 740 -2324 745 -2296
rect -745 -2362 745 -2324
rect -745 -2390 -740 -2362
rect -712 -2390 -674 -2362
rect -646 -2390 -608 -2362
rect -580 -2390 -542 -2362
rect -514 -2390 -476 -2362
rect -448 -2390 -410 -2362
rect -382 -2390 -344 -2362
rect -316 -2390 -278 -2362
rect -250 -2390 -212 -2362
rect -184 -2390 -146 -2362
rect -118 -2390 -80 -2362
rect -52 -2390 -14 -2362
rect 14 -2390 52 -2362
rect 80 -2390 118 -2362
rect 146 -2390 184 -2362
rect 212 -2390 250 -2362
rect 278 -2390 316 -2362
rect 344 -2390 382 -2362
rect 410 -2390 448 -2362
rect 476 -2390 514 -2362
rect 542 -2390 580 -2362
rect 608 -2390 646 -2362
rect 674 -2390 712 -2362
rect 740 -2390 745 -2362
rect -745 -2428 745 -2390
rect -745 -2456 -740 -2428
rect -712 -2456 -674 -2428
rect -646 -2456 -608 -2428
rect -580 -2456 -542 -2428
rect -514 -2456 -476 -2428
rect -448 -2456 -410 -2428
rect -382 -2456 -344 -2428
rect -316 -2456 -278 -2428
rect -250 -2456 -212 -2428
rect -184 -2456 -146 -2428
rect -118 -2456 -80 -2428
rect -52 -2456 -14 -2428
rect 14 -2456 52 -2428
rect 80 -2456 118 -2428
rect 146 -2456 184 -2428
rect 212 -2456 250 -2428
rect 278 -2456 316 -2428
rect 344 -2456 382 -2428
rect 410 -2456 448 -2428
rect 476 -2456 514 -2428
rect 542 -2456 580 -2428
rect 608 -2456 646 -2428
rect 674 -2456 712 -2428
rect 740 -2456 745 -2428
rect -745 -2494 745 -2456
rect -745 -2522 -740 -2494
rect -712 -2522 -674 -2494
rect -646 -2522 -608 -2494
rect -580 -2522 -542 -2494
rect -514 -2522 -476 -2494
rect -448 -2522 -410 -2494
rect -382 -2522 -344 -2494
rect -316 -2522 -278 -2494
rect -250 -2522 -212 -2494
rect -184 -2522 -146 -2494
rect -118 -2522 -80 -2494
rect -52 -2522 -14 -2494
rect 14 -2522 52 -2494
rect 80 -2522 118 -2494
rect 146 -2522 184 -2494
rect 212 -2522 250 -2494
rect 278 -2522 316 -2494
rect 344 -2522 382 -2494
rect 410 -2522 448 -2494
rect 476 -2522 514 -2494
rect 542 -2522 580 -2494
rect 608 -2522 646 -2494
rect 674 -2522 712 -2494
rect 740 -2522 745 -2494
rect -745 -2560 745 -2522
rect -745 -2588 -740 -2560
rect -712 -2588 -674 -2560
rect -646 -2588 -608 -2560
rect -580 -2588 -542 -2560
rect -514 -2588 -476 -2560
rect -448 -2588 -410 -2560
rect -382 -2588 -344 -2560
rect -316 -2588 -278 -2560
rect -250 -2588 -212 -2560
rect -184 -2588 -146 -2560
rect -118 -2588 -80 -2560
rect -52 -2588 -14 -2560
rect 14 -2588 52 -2560
rect 80 -2588 118 -2560
rect 146 -2588 184 -2560
rect 212 -2588 250 -2560
rect 278 -2588 316 -2560
rect 344 -2588 382 -2560
rect 410 -2588 448 -2560
rect 476 -2588 514 -2560
rect 542 -2588 580 -2560
rect 608 -2588 646 -2560
rect 674 -2588 712 -2560
rect 740 -2588 745 -2560
rect -745 -2626 745 -2588
rect -745 -2654 -740 -2626
rect -712 -2654 -674 -2626
rect -646 -2654 -608 -2626
rect -580 -2654 -542 -2626
rect -514 -2654 -476 -2626
rect -448 -2654 -410 -2626
rect -382 -2654 -344 -2626
rect -316 -2654 -278 -2626
rect -250 -2654 -212 -2626
rect -184 -2654 -146 -2626
rect -118 -2654 -80 -2626
rect -52 -2654 -14 -2626
rect 14 -2654 52 -2626
rect 80 -2654 118 -2626
rect 146 -2654 184 -2626
rect 212 -2654 250 -2626
rect 278 -2654 316 -2626
rect 344 -2654 382 -2626
rect 410 -2654 448 -2626
rect 476 -2654 514 -2626
rect 542 -2654 580 -2626
rect 608 -2654 646 -2626
rect 674 -2654 712 -2626
rect 740 -2654 745 -2626
rect -745 -2692 745 -2654
rect -745 -2720 -740 -2692
rect -712 -2720 -674 -2692
rect -646 -2720 -608 -2692
rect -580 -2720 -542 -2692
rect -514 -2720 -476 -2692
rect -448 -2720 -410 -2692
rect -382 -2720 -344 -2692
rect -316 -2720 -278 -2692
rect -250 -2720 -212 -2692
rect -184 -2720 -146 -2692
rect -118 -2720 -80 -2692
rect -52 -2720 -14 -2692
rect 14 -2720 52 -2692
rect 80 -2720 118 -2692
rect 146 -2720 184 -2692
rect 212 -2720 250 -2692
rect 278 -2720 316 -2692
rect 344 -2720 382 -2692
rect 410 -2720 448 -2692
rect 476 -2720 514 -2692
rect 542 -2720 580 -2692
rect 608 -2720 646 -2692
rect 674 -2720 712 -2692
rect 740 -2720 745 -2692
rect -745 -2758 745 -2720
rect -745 -2786 -740 -2758
rect -712 -2786 -674 -2758
rect -646 -2786 -608 -2758
rect -580 -2786 -542 -2758
rect -514 -2786 -476 -2758
rect -448 -2786 -410 -2758
rect -382 -2786 -344 -2758
rect -316 -2786 -278 -2758
rect -250 -2786 -212 -2758
rect -184 -2786 -146 -2758
rect -118 -2786 -80 -2758
rect -52 -2786 -14 -2758
rect 14 -2786 52 -2758
rect 80 -2786 118 -2758
rect 146 -2786 184 -2758
rect 212 -2786 250 -2758
rect 278 -2786 316 -2758
rect 344 -2786 382 -2758
rect 410 -2786 448 -2758
rect 476 -2786 514 -2758
rect 542 -2786 580 -2758
rect 608 -2786 646 -2758
rect 674 -2786 712 -2758
rect 740 -2786 745 -2758
rect -745 -2824 745 -2786
rect -745 -2852 -740 -2824
rect -712 -2852 -674 -2824
rect -646 -2852 -608 -2824
rect -580 -2852 -542 -2824
rect -514 -2852 -476 -2824
rect -448 -2852 -410 -2824
rect -382 -2852 -344 -2824
rect -316 -2852 -278 -2824
rect -250 -2852 -212 -2824
rect -184 -2852 -146 -2824
rect -118 -2852 -80 -2824
rect -52 -2852 -14 -2824
rect 14 -2852 52 -2824
rect 80 -2852 118 -2824
rect 146 -2852 184 -2824
rect 212 -2852 250 -2824
rect 278 -2852 316 -2824
rect 344 -2852 382 -2824
rect 410 -2852 448 -2824
rect 476 -2852 514 -2824
rect 542 -2852 580 -2824
rect 608 -2852 646 -2824
rect 674 -2852 712 -2824
rect 740 -2852 745 -2824
rect -745 -2890 745 -2852
rect -745 -2918 -740 -2890
rect -712 -2918 -674 -2890
rect -646 -2918 -608 -2890
rect -580 -2918 -542 -2890
rect -514 -2918 -476 -2890
rect -448 -2918 -410 -2890
rect -382 -2918 -344 -2890
rect -316 -2918 -278 -2890
rect -250 -2918 -212 -2890
rect -184 -2918 -146 -2890
rect -118 -2918 -80 -2890
rect -52 -2918 -14 -2890
rect 14 -2918 52 -2890
rect 80 -2918 118 -2890
rect 146 -2918 184 -2890
rect 212 -2918 250 -2890
rect 278 -2918 316 -2890
rect 344 -2918 382 -2890
rect 410 -2918 448 -2890
rect 476 -2918 514 -2890
rect 542 -2918 580 -2890
rect 608 -2918 646 -2890
rect 674 -2918 712 -2890
rect 740 -2918 745 -2890
rect -745 -2956 745 -2918
rect -745 -2984 -740 -2956
rect -712 -2984 -674 -2956
rect -646 -2984 -608 -2956
rect -580 -2984 -542 -2956
rect -514 -2984 -476 -2956
rect -448 -2984 -410 -2956
rect -382 -2984 -344 -2956
rect -316 -2984 -278 -2956
rect -250 -2984 -212 -2956
rect -184 -2984 -146 -2956
rect -118 -2984 -80 -2956
rect -52 -2984 -14 -2956
rect 14 -2984 52 -2956
rect 80 -2984 118 -2956
rect 146 -2984 184 -2956
rect 212 -2984 250 -2956
rect 278 -2984 316 -2956
rect 344 -2984 382 -2956
rect 410 -2984 448 -2956
rect 476 -2984 514 -2956
rect 542 -2984 580 -2956
rect 608 -2984 646 -2956
rect 674 -2984 712 -2956
rect 740 -2984 745 -2956
rect -745 -3022 745 -2984
rect -745 -3050 -740 -3022
rect -712 -3050 -674 -3022
rect -646 -3050 -608 -3022
rect -580 -3050 -542 -3022
rect -514 -3050 -476 -3022
rect -448 -3050 -410 -3022
rect -382 -3050 -344 -3022
rect -316 -3050 -278 -3022
rect -250 -3050 -212 -3022
rect -184 -3050 -146 -3022
rect -118 -3050 -80 -3022
rect -52 -3050 -14 -3022
rect 14 -3050 52 -3022
rect 80 -3050 118 -3022
rect 146 -3050 184 -3022
rect 212 -3050 250 -3022
rect 278 -3050 316 -3022
rect 344 -3050 382 -3022
rect 410 -3050 448 -3022
rect 476 -3050 514 -3022
rect 542 -3050 580 -3022
rect 608 -3050 646 -3022
rect 674 -3050 712 -3022
rect 740 -3050 745 -3022
rect -745 -3088 745 -3050
rect -745 -3116 -740 -3088
rect -712 -3116 -674 -3088
rect -646 -3116 -608 -3088
rect -580 -3116 -542 -3088
rect -514 -3116 -476 -3088
rect -448 -3116 -410 -3088
rect -382 -3116 -344 -3088
rect -316 -3116 -278 -3088
rect -250 -3116 -212 -3088
rect -184 -3116 -146 -3088
rect -118 -3116 -80 -3088
rect -52 -3116 -14 -3088
rect 14 -3116 52 -3088
rect 80 -3116 118 -3088
rect 146 -3116 184 -3088
rect 212 -3116 250 -3088
rect 278 -3116 316 -3088
rect 344 -3116 382 -3088
rect 410 -3116 448 -3088
rect 476 -3116 514 -3088
rect 542 -3116 580 -3088
rect 608 -3116 646 -3088
rect 674 -3116 712 -3088
rect 740 -3116 745 -3088
rect -745 -3154 745 -3116
rect -745 -3182 -740 -3154
rect -712 -3182 -674 -3154
rect -646 -3182 -608 -3154
rect -580 -3182 -542 -3154
rect -514 -3182 -476 -3154
rect -448 -3182 -410 -3154
rect -382 -3182 -344 -3154
rect -316 -3182 -278 -3154
rect -250 -3182 -212 -3154
rect -184 -3182 -146 -3154
rect -118 -3182 -80 -3154
rect -52 -3182 -14 -3154
rect 14 -3182 52 -3154
rect 80 -3182 118 -3154
rect 146 -3182 184 -3154
rect 212 -3182 250 -3154
rect 278 -3182 316 -3154
rect 344 -3182 382 -3154
rect 410 -3182 448 -3154
rect 476 -3182 514 -3154
rect 542 -3182 580 -3154
rect 608 -3182 646 -3154
rect 674 -3182 712 -3154
rect 740 -3182 745 -3154
rect -745 -3220 745 -3182
rect -745 -3248 -740 -3220
rect -712 -3248 -674 -3220
rect -646 -3248 -608 -3220
rect -580 -3248 -542 -3220
rect -514 -3248 -476 -3220
rect -448 -3248 -410 -3220
rect -382 -3248 -344 -3220
rect -316 -3248 -278 -3220
rect -250 -3248 -212 -3220
rect -184 -3248 -146 -3220
rect -118 -3248 -80 -3220
rect -52 -3248 -14 -3220
rect 14 -3248 52 -3220
rect 80 -3248 118 -3220
rect 146 -3248 184 -3220
rect 212 -3248 250 -3220
rect 278 -3248 316 -3220
rect 344 -3248 382 -3220
rect 410 -3248 448 -3220
rect 476 -3248 514 -3220
rect 542 -3248 580 -3220
rect 608 -3248 646 -3220
rect 674 -3248 712 -3220
rect 740 -3248 745 -3220
rect -745 -3286 745 -3248
rect -745 -3314 -740 -3286
rect -712 -3314 -674 -3286
rect -646 -3314 -608 -3286
rect -580 -3314 -542 -3286
rect -514 -3314 -476 -3286
rect -448 -3314 -410 -3286
rect -382 -3314 -344 -3286
rect -316 -3314 -278 -3286
rect -250 -3314 -212 -3286
rect -184 -3314 -146 -3286
rect -118 -3314 -80 -3286
rect -52 -3314 -14 -3286
rect 14 -3314 52 -3286
rect 80 -3314 118 -3286
rect 146 -3314 184 -3286
rect 212 -3314 250 -3286
rect 278 -3314 316 -3286
rect 344 -3314 382 -3286
rect 410 -3314 448 -3286
rect 476 -3314 514 -3286
rect 542 -3314 580 -3286
rect 608 -3314 646 -3286
rect 674 -3314 712 -3286
rect 740 -3314 745 -3286
rect -745 -3352 745 -3314
rect -745 -3380 -740 -3352
rect -712 -3380 -674 -3352
rect -646 -3380 -608 -3352
rect -580 -3380 -542 -3352
rect -514 -3380 -476 -3352
rect -448 -3380 -410 -3352
rect -382 -3380 -344 -3352
rect -316 -3380 -278 -3352
rect -250 -3380 -212 -3352
rect -184 -3380 -146 -3352
rect -118 -3380 -80 -3352
rect -52 -3380 -14 -3352
rect 14 -3380 52 -3352
rect 80 -3380 118 -3352
rect 146 -3380 184 -3352
rect 212 -3380 250 -3352
rect 278 -3380 316 -3352
rect 344 -3380 382 -3352
rect 410 -3380 448 -3352
rect 476 -3380 514 -3352
rect 542 -3380 580 -3352
rect 608 -3380 646 -3352
rect 674 -3380 712 -3352
rect 740 -3380 745 -3352
rect -745 -3418 745 -3380
rect -745 -3446 -740 -3418
rect -712 -3446 -674 -3418
rect -646 -3446 -608 -3418
rect -580 -3446 -542 -3418
rect -514 -3446 -476 -3418
rect -448 -3446 -410 -3418
rect -382 -3446 -344 -3418
rect -316 -3446 -278 -3418
rect -250 -3446 -212 -3418
rect -184 -3446 -146 -3418
rect -118 -3446 -80 -3418
rect -52 -3446 -14 -3418
rect 14 -3446 52 -3418
rect 80 -3446 118 -3418
rect 146 -3446 184 -3418
rect 212 -3446 250 -3418
rect 278 -3446 316 -3418
rect 344 -3446 382 -3418
rect 410 -3446 448 -3418
rect 476 -3446 514 -3418
rect 542 -3446 580 -3418
rect 608 -3446 646 -3418
rect 674 -3446 712 -3418
rect 740 -3446 745 -3418
rect -745 -3484 745 -3446
rect -745 -3512 -740 -3484
rect -712 -3512 -674 -3484
rect -646 -3512 -608 -3484
rect -580 -3512 -542 -3484
rect -514 -3512 -476 -3484
rect -448 -3512 -410 -3484
rect -382 -3512 -344 -3484
rect -316 -3512 -278 -3484
rect -250 -3512 -212 -3484
rect -184 -3512 -146 -3484
rect -118 -3512 -80 -3484
rect -52 -3512 -14 -3484
rect 14 -3512 52 -3484
rect 80 -3512 118 -3484
rect 146 -3512 184 -3484
rect 212 -3512 250 -3484
rect 278 -3512 316 -3484
rect 344 -3512 382 -3484
rect 410 -3512 448 -3484
rect 476 -3512 514 -3484
rect 542 -3512 580 -3484
rect 608 -3512 646 -3484
rect 674 -3512 712 -3484
rect 740 -3512 745 -3484
rect -745 -3550 745 -3512
rect -745 -3578 -740 -3550
rect -712 -3578 -674 -3550
rect -646 -3578 -608 -3550
rect -580 -3578 -542 -3550
rect -514 -3578 -476 -3550
rect -448 -3578 -410 -3550
rect -382 -3578 -344 -3550
rect -316 -3578 -278 -3550
rect -250 -3578 -212 -3550
rect -184 -3578 -146 -3550
rect -118 -3578 -80 -3550
rect -52 -3578 -14 -3550
rect 14 -3578 52 -3550
rect 80 -3578 118 -3550
rect 146 -3578 184 -3550
rect 212 -3578 250 -3550
rect 278 -3578 316 -3550
rect 344 -3578 382 -3550
rect 410 -3578 448 -3550
rect 476 -3578 514 -3550
rect 542 -3578 580 -3550
rect 608 -3578 646 -3550
rect 674 -3578 712 -3550
rect 740 -3578 745 -3550
rect -745 -3616 745 -3578
rect -745 -3644 -740 -3616
rect -712 -3644 -674 -3616
rect -646 -3644 -608 -3616
rect -580 -3644 -542 -3616
rect -514 -3644 -476 -3616
rect -448 -3644 -410 -3616
rect -382 -3644 -344 -3616
rect -316 -3644 -278 -3616
rect -250 -3644 -212 -3616
rect -184 -3644 -146 -3616
rect -118 -3644 -80 -3616
rect -52 -3644 -14 -3616
rect 14 -3644 52 -3616
rect 80 -3644 118 -3616
rect 146 -3644 184 -3616
rect 212 -3644 250 -3616
rect 278 -3644 316 -3616
rect 344 -3644 382 -3616
rect 410 -3644 448 -3616
rect 476 -3644 514 -3616
rect 542 -3644 580 -3616
rect 608 -3644 646 -3616
rect 674 -3644 712 -3616
rect 740 -3644 745 -3616
rect -745 -3682 745 -3644
rect -745 -3710 -740 -3682
rect -712 -3710 -674 -3682
rect -646 -3710 -608 -3682
rect -580 -3710 -542 -3682
rect -514 -3710 -476 -3682
rect -448 -3710 -410 -3682
rect -382 -3710 -344 -3682
rect -316 -3710 -278 -3682
rect -250 -3710 -212 -3682
rect -184 -3710 -146 -3682
rect -118 -3710 -80 -3682
rect -52 -3710 -14 -3682
rect 14 -3710 52 -3682
rect 80 -3710 118 -3682
rect 146 -3710 184 -3682
rect 212 -3710 250 -3682
rect 278 -3710 316 -3682
rect 344 -3710 382 -3682
rect 410 -3710 448 -3682
rect 476 -3710 514 -3682
rect 542 -3710 580 -3682
rect 608 -3710 646 -3682
rect 674 -3710 712 -3682
rect 740 -3710 745 -3682
rect -745 -3748 745 -3710
rect -745 -3776 -740 -3748
rect -712 -3776 -674 -3748
rect -646 -3776 -608 -3748
rect -580 -3776 -542 -3748
rect -514 -3776 -476 -3748
rect -448 -3776 -410 -3748
rect -382 -3776 -344 -3748
rect -316 -3776 -278 -3748
rect -250 -3776 -212 -3748
rect -184 -3776 -146 -3748
rect -118 -3776 -80 -3748
rect -52 -3776 -14 -3748
rect 14 -3776 52 -3748
rect 80 -3776 118 -3748
rect 146 -3776 184 -3748
rect 212 -3776 250 -3748
rect 278 -3776 316 -3748
rect 344 -3776 382 -3748
rect 410 -3776 448 -3748
rect 476 -3776 514 -3748
rect 542 -3776 580 -3748
rect 608 -3776 646 -3748
rect 674 -3776 712 -3748
rect 740 -3776 745 -3748
rect -745 -3814 745 -3776
rect -745 -3842 -740 -3814
rect -712 -3842 -674 -3814
rect -646 -3842 -608 -3814
rect -580 -3842 -542 -3814
rect -514 -3842 -476 -3814
rect -448 -3842 -410 -3814
rect -382 -3842 -344 -3814
rect -316 -3842 -278 -3814
rect -250 -3842 -212 -3814
rect -184 -3842 -146 -3814
rect -118 -3842 -80 -3814
rect -52 -3842 -14 -3814
rect 14 -3842 52 -3814
rect 80 -3842 118 -3814
rect 146 -3842 184 -3814
rect 212 -3842 250 -3814
rect 278 -3842 316 -3814
rect 344 -3842 382 -3814
rect 410 -3842 448 -3814
rect 476 -3842 514 -3814
rect 542 -3842 580 -3814
rect 608 -3842 646 -3814
rect 674 -3842 712 -3814
rect 740 -3842 745 -3814
rect -745 -3880 745 -3842
rect -745 -3908 -740 -3880
rect -712 -3908 -674 -3880
rect -646 -3908 -608 -3880
rect -580 -3908 -542 -3880
rect -514 -3908 -476 -3880
rect -448 -3908 -410 -3880
rect -382 -3908 -344 -3880
rect -316 -3908 -278 -3880
rect -250 -3908 -212 -3880
rect -184 -3908 -146 -3880
rect -118 -3908 -80 -3880
rect -52 -3908 -14 -3880
rect 14 -3908 52 -3880
rect 80 -3908 118 -3880
rect 146 -3908 184 -3880
rect 212 -3908 250 -3880
rect 278 -3908 316 -3880
rect 344 -3908 382 -3880
rect 410 -3908 448 -3880
rect 476 -3908 514 -3880
rect 542 -3908 580 -3880
rect 608 -3908 646 -3880
rect 674 -3908 712 -3880
rect 740 -3908 745 -3880
rect -745 -3946 745 -3908
rect -745 -3974 -740 -3946
rect -712 -3974 -674 -3946
rect -646 -3974 -608 -3946
rect -580 -3974 -542 -3946
rect -514 -3974 -476 -3946
rect -448 -3974 -410 -3946
rect -382 -3974 -344 -3946
rect -316 -3974 -278 -3946
rect -250 -3974 -212 -3946
rect -184 -3974 -146 -3946
rect -118 -3974 -80 -3946
rect -52 -3974 -14 -3946
rect 14 -3974 52 -3946
rect 80 -3974 118 -3946
rect 146 -3974 184 -3946
rect 212 -3974 250 -3946
rect 278 -3974 316 -3946
rect 344 -3974 382 -3946
rect 410 -3974 448 -3946
rect 476 -3974 514 -3946
rect 542 -3974 580 -3946
rect 608 -3974 646 -3946
rect 674 -3974 712 -3946
rect 740 -3974 745 -3946
rect -745 -4012 745 -3974
rect -745 -4040 -740 -4012
rect -712 -4040 -674 -4012
rect -646 -4040 -608 -4012
rect -580 -4040 -542 -4012
rect -514 -4040 -476 -4012
rect -448 -4040 -410 -4012
rect -382 -4040 -344 -4012
rect -316 -4040 -278 -4012
rect -250 -4040 -212 -4012
rect -184 -4040 -146 -4012
rect -118 -4040 -80 -4012
rect -52 -4040 -14 -4012
rect 14 -4040 52 -4012
rect 80 -4040 118 -4012
rect 146 -4040 184 -4012
rect 212 -4040 250 -4012
rect 278 -4040 316 -4012
rect 344 -4040 382 -4012
rect 410 -4040 448 -4012
rect 476 -4040 514 -4012
rect 542 -4040 580 -4012
rect 608 -4040 646 -4012
rect 674 -4040 712 -4012
rect 740 -4040 745 -4012
rect -745 -4078 745 -4040
rect -745 -4106 -740 -4078
rect -712 -4106 -674 -4078
rect -646 -4106 -608 -4078
rect -580 -4106 -542 -4078
rect -514 -4106 -476 -4078
rect -448 -4106 -410 -4078
rect -382 -4106 -344 -4078
rect -316 -4106 -278 -4078
rect -250 -4106 -212 -4078
rect -184 -4106 -146 -4078
rect -118 -4106 -80 -4078
rect -52 -4106 -14 -4078
rect 14 -4106 52 -4078
rect 80 -4106 118 -4078
rect 146 -4106 184 -4078
rect 212 -4106 250 -4078
rect 278 -4106 316 -4078
rect 344 -4106 382 -4078
rect 410 -4106 448 -4078
rect 476 -4106 514 -4078
rect 542 -4106 580 -4078
rect 608 -4106 646 -4078
rect 674 -4106 712 -4078
rect 740 -4106 745 -4078
rect -745 -4144 745 -4106
rect -745 -4172 -740 -4144
rect -712 -4172 -674 -4144
rect -646 -4172 -608 -4144
rect -580 -4172 -542 -4144
rect -514 -4172 -476 -4144
rect -448 -4172 -410 -4144
rect -382 -4172 -344 -4144
rect -316 -4172 -278 -4144
rect -250 -4172 -212 -4144
rect -184 -4172 -146 -4144
rect -118 -4172 -80 -4144
rect -52 -4172 -14 -4144
rect 14 -4172 52 -4144
rect 80 -4172 118 -4144
rect 146 -4172 184 -4144
rect 212 -4172 250 -4144
rect 278 -4172 316 -4144
rect 344 -4172 382 -4144
rect 410 -4172 448 -4144
rect 476 -4172 514 -4144
rect 542 -4172 580 -4144
rect 608 -4172 646 -4144
rect 674 -4172 712 -4144
rect 740 -4172 745 -4144
rect -745 -4210 745 -4172
rect -745 -4238 -740 -4210
rect -712 -4238 -674 -4210
rect -646 -4238 -608 -4210
rect -580 -4238 -542 -4210
rect -514 -4238 -476 -4210
rect -448 -4238 -410 -4210
rect -382 -4238 -344 -4210
rect -316 -4238 -278 -4210
rect -250 -4238 -212 -4210
rect -184 -4238 -146 -4210
rect -118 -4238 -80 -4210
rect -52 -4238 -14 -4210
rect 14 -4238 52 -4210
rect 80 -4238 118 -4210
rect 146 -4238 184 -4210
rect 212 -4238 250 -4210
rect 278 -4238 316 -4210
rect 344 -4238 382 -4210
rect 410 -4238 448 -4210
rect 476 -4238 514 -4210
rect 542 -4238 580 -4210
rect 608 -4238 646 -4210
rect 674 -4238 712 -4210
rect 740 -4238 745 -4210
rect -745 -4276 745 -4238
rect -745 -4304 -740 -4276
rect -712 -4304 -674 -4276
rect -646 -4304 -608 -4276
rect -580 -4304 -542 -4276
rect -514 -4304 -476 -4276
rect -448 -4304 -410 -4276
rect -382 -4304 -344 -4276
rect -316 -4304 -278 -4276
rect -250 -4304 -212 -4276
rect -184 -4304 -146 -4276
rect -118 -4304 -80 -4276
rect -52 -4304 -14 -4276
rect 14 -4304 52 -4276
rect 80 -4304 118 -4276
rect 146 -4304 184 -4276
rect 212 -4304 250 -4276
rect 278 -4304 316 -4276
rect 344 -4304 382 -4276
rect 410 -4304 448 -4276
rect 476 -4304 514 -4276
rect 542 -4304 580 -4276
rect 608 -4304 646 -4276
rect 674 -4304 712 -4276
rect 740 -4304 745 -4276
rect -745 -4342 745 -4304
rect -745 -4370 -740 -4342
rect -712 -4370 -674 -4342
rect -646 -4370 -608 -4342
rect -580 -4370 -542 -4342
rect -514 -4370 -476 -4342
rect -448 -4370 -410 -4342
rect -382 -4370 -344 -4342
rect -316 -4370 -278 -4342
rect -250 -4370 -212 -4342
rect -184 -4370 -146 -4342
rect -118 -4370 -80 -4342
rect -52 -4370 -14 -4342
rect 14 -4370 52 -4342
rect 80 -4370 118 -4342
rect 146 -4370 184 -4342
rect 212 -4370 250 -4342
rect 278 -4370 316 -4342
rect 344 -4370 382 -4342
rect 410 -4370 448 -4342
rect 476 -4370 514 -4342
rect 542 -4370 580 -4342
rect 608 -4370 646 -4342
rect 674 -4370 712 -4342
rect 740 -4370 745 -4342
rect -745 -4408 745 -4370
rect -745 -4436 -740 -4408
rect -712 -4436 -674 -4408
rect -646 -4436 -608 -4408
rect -580 -4436 -542 -4408
rect -514 -4436 -476 -4408
rect -448 -4436 -410 -4408
rect -382 -4436 -344 -4408
rect -316 -4436 -278 -4408
rect -250 -4436 -212 -4408
rect -184 -4436 -146 -4408
rect -118 -4436 -80 -4408
rect -52 -4436 -14 -4408
rect 14 -4436 52 -4408
rect 80 -4436 118 -4408
rect 146 -4436 184 -4408
rect 212 -4436 250 -4408
rect 278 -4436 316 -4408
rect 344 -4436 382 -4408
rect 410 -4436 448 -4408
rect 476 -4436 514 -4408
rect 542 -4436 580 -4408
rect 608 -4436 646 -4408
rect 674 -4436 712 -4408
rect 740 -4436 745 -4408
rect -745 -4474 745 -4436
rect -745 -4502 -740 -4474
rect -712 -4502 -674 -4474
rect -646 -4502 -608 -4474
rect -580 -4502 -542 -4474
rect -514 -4502 -476 -4474
rect -448 -4502 -410 -4474
rect -382 -4502 -344 -4474
rect -316 -4502 -278 -4474
rect -250 -4502 -212 -4474
rect -184 -4502 -146 -4474
rect -118 -4502 -80 -4474
rect -52 -4502 -14 -4474
rect 14 -4502 52 -4474
rect 80 -4502 118 -4474
rect 146 -4502 184 -4474
rect 212 -4502 250 -4474
rect 278 -4502 316 -4474
rect 344 -4502 382 -4474
rect 410 -4502 448 -4474
rect 476 -4502 514 -4474
rect 542 -4502 580 -4474
rect 608 -4502 646 -4474
rect 674 -4502 712 -4474
rect 740 -4502 745 -4474
rect -745 -4540 745 -4502
rect -745 -4568 -740 -4540
rect -712 -4568 -674 -4540
rect -646 -4568 -608 -4540
rect -580 -4568 -542 -4540
rect -514 -4568 -476 -4540
rect -448 -4568 -410 -4540
rect -382 -4568 -344 -4540
rect -316 -4568 -278 -4540
rect -250 -4568 -212 -4540
rect -184 -4568 -146 -4540
rect -118 -4568 -80 -4540
rect -52 -4568 -14 -4540
rect 14 -4568 52 -4540
rect 80 -4568 118 -4540
rect 146 -4568 184 -4540
rect 212 -4568 250 -4540
rect 278 -4568 316 -4540
rect 344 -4568 382 -4540
rect 410 -4568 448 -4540
rect 476 -4568 514 -4540
rect 542 -4568 580 -4540
rect 608 -4568 646 -4540
rect 674 -4568 712 -4540
rect 740 -4568 745 -4540
rect -745 -4606 745 -4568
rect -745 -4634 -740 -4606
rect -712 -4634 -674 -4606
rect -646 -4634 -608 -4606
rect -580 -4634 -542 -4606
rect -514 -4634 -476 -4606
rect -448 -4634 -410 -4606
rect -382 -4634 -344 -4606
rect -316 -4634 -278 -4606
rect -250 -4634 -212 -4606
rect -184 -4634 -146 -4606
rect -118 -4634 -80 -4606
rect -52 -4634 -14 -4606
rect 14 -4634 52 -4606
rect 80 -4634 118 -4606
rect 146 -4634 184 -4606
rect 212 -4634 250 -4606
rect 278 -4634 316 -4606
rect 344 -4634 382 -4606
rect 410 -4634 448 -4606
rect 476 -4634 514 -4606
rect 542 -4634 580 -4606
rect 608 -4634 646 -4606
rect 674 -4634 712 -4606
rect 740 -4634 745 -4606
rect -745 -4672 745 -4634
rect -745 -4700 -740 -4672
rect -712 -4700 -674 -4672
rect -646 -4700 -608 -4672
rect -580 -4700 -542 -4672
rect -514 -4700 -476 -4672
rect -448 -4700 -410 -4672
rect -382 -4700 -344 -4672
rect -316 -4700 -278 -4672
rect -250 -4700 -212 -4672
rect -184 -4700 -146 -4672
rect -118 -4700 -80 -4672
rect -52 -4700 -14 -4672
rect 14 -4700 52 -4672
rect 80 -4700 118 -4672
rect 146 -4700 184 -4672
rect 212 -4700 250 -4672
rect 278 -4700 316 -4672
rect 344 -4700 382 -4672
rect 410 -4700 448 -4672
rect 476 -4700 514 -4672
rect 542 -4700 580 -4672
rect 608 -4700 646 -4672
rect 674 -4700 712 -4672
rect 740 -4700 745 -4672
rect -745 -4738 745 -4700
rect -745 -4766 -740 -4738
rect -712 -4766 -674 -4738
rect -646 -4766 -608 -4738
rect -580 -4766 -542 -4738
rect -514 -4766 -476 -4738
rect -448 -4766 -410 -4738
rect -382 -4766 -344 -4738
rect -316 -4766 -278 -4738
rect -250 -4766 -212 -4738
rect -184 -4766 -146 -4738
rect -118 -4766 -80 -4738
rect -52 -4766 -14 -4738
rect 14 -4766 52 -4738
rect 80 -4766 118 -4738
rect 146 -4766 184 -4738
rect 212 -4766 250 -4738
rect 278 -4766 316 -4738
rect 344 -4766 382 -4738
rect 410 -4766 448 -4738
rect 476 -4766 514 -4738
rect 542 -4766 580 -4738
rect 608 -4766 646 -4738
rect 674 -4766 712 -4738
rect 740 -4766 745 -4738
rect -745 -4804 745 -4766
rect -745 -4832 -740 -4804
rect -712 -4832 -674 -4804
rect -646 -4832 -608 -4804
rect -580 -4832 -542 -4804
rect -514 -4832 -476 -4804
rect -448 -4832 -410 -4804
rect -382 -4832 -344 -4804
rect -316 -4832 -278 -4804
rect -250 -4832 -212 -4804
rect -184 -4832 -146 -4804
rect -118 -4832 -80 -4804
rect -52 -4832 -14 -4804
rect 14 -4832 52 -4804
rect 80 -4832 118 -4804
rect 146 -4832 184 -4804
rect 212 -4832 250 -4804
rect 278 -4832 316 -4804
rect 344 -4832 382 -4804
rect 410 -4832 448 -4804
rect 476 -4832 514 -4804
rect 542 -4832 580 -4804
rect 608 -4832 646 -4804
rect 674 -4832 712 -4804
rect 740 -4832 745 -4804
rect -745 -4870 745 -4832
rect -745 -4898 -740 -4870
rect -712 -4898 -674 -4870
rect -646 -4898 -608 -4870
rect -580 -4898 -542 -4870
rect -514 -4898 -476 -4870
rect -448 -4898 -410 -4870
rect -382 -4898 -344 -4870
rect -316 -4898 -278 -4870
rect -250 -4898 -212 -4870
rect -184 -4898 -146 -4870
rect -118 -4898 -80 -4870
rect -52 -4898 -14 -4870
rect 14 -4898 52 -4870
rect 80 -4898 118 -4870
rect 146 -4898 184 -4870
rect 212 -4898 250 -4870
rect 278 -4898 316 -4870
rect 344 -4898 382 -4870
rect 410 -4898 448 -4870
rect 476 -4898 514 -4870
rect 542 -4898 580 -4870
rect 608 -4898 646 -4870
rect 674 -4898 712 -4870
rect 740 -4898 745 -4870
rect -745 -4936 745 -4898
rect -745 -4964 -740 -4936
rect -712 -4964 -674 -4936
rect -646 -4964 -608 -4936
rect -580 -4964 -542 -4936
rect -514 -4964 -476 -4936
rect -448 -4964 -410 -4936
rect -382 -4964 -344 -4936
rect -316 -4964 -278 -4936
rect -250 -4964 -212 -4936
rect -184 -4964 -146 -4936
rect -118 -4964 -80 -4936
rect -52 -4964 -14 -4936
rect 14 -4964 52 -4936
rect 80 -4964 118 -4936
rect 146 -4964 184 -4936
rect 212 -4964 250 -4936
rect 278 -4964 316 -4936
rect 344 -4964 382 -4936
rect 410 -4964 448 -4936
rect 476 -4964 514 -4936
rect 542 -4964 580 -4936
rect 608 -4964 646 -4936
rect 674 -4964 712 -4936
rect 740 -4964 745 -4936
rect -745 -5002 745 -4964
rect -745 -5030 -740 -5002
rect -712 -5030 -674 -5002
rect -646 -5030 -608 -5002
rect -580 -5030 -542 -5002
rect -514 -5030 -476 -5002
rect -448 -5030 -410 -5002
rect -382 -5030 -344 -5002
rect -316 -5030 -278 -5002
rect -250 -5030 -212 -5002
rect -184 -5030 -146 -5002
rect -118 -5030 -80 -5002
rect -52 -5030 -14 -5002
rect 14 -5030 52 -5002
rect 80 -5030 118 -5002
rect 146 -5030 184 -5002
rect 212 -5030 250 -5002
rect 278 -5030 316 -5002
rect 344 -5030 382 -5002
rect 410 -5030 448 -5002
rect 476 -5030 514 -5002
rect 542 -5030 580 -5002
rect 608 -5030 646 -5002
rect 674 -5030 712 -5002
rect 740 -5030 745 -5002
rect -745 -5068 745 -5030
rect -745 -5096 -740 -5068
rect -712 -5096 -674 -5068
rect -646 -5096 -608 -5068
rect -580 -5096 -542 -5068
rect -514 -5096 -476 -5068
rect -448 -5096 -410 -5068
rect -382 -5096 -344 -5068
rect -316 -5096 -278 -5068
rect -250 -5096 -212 -5068
rect -184 -5096 -146 -5068
rect -118 -5096 -80 -5068
rect -52 -5096 -14 -5068
rect 14 -5096 52 -5068
rect 80 -5096 118 -5068
rect 146 -5096 184 -5068
rect 212 -5096 250 -5068
rect 278 -5096 316 -5068
rect 344 -5096 382 -5068
rect 410 -5096 448 -5068
rect 476 -5096 514 -5068
rect 542 -5096 580 -5068
rect 608 -5096 646 -5068
rect 674 -5096 712 -5068
rect 740 -5096 745 -5068
rect -745 -5134 745 -5096
rect -745 -5162 -740 -5134
rect -712 -5162 -674 -5134
rect -646 -5162 -608 -5134
rect -580 -5162 -542 -5134
rect -514 -5162 -476 -5134
rect -448 -5162 -410 -5134
rect -382 -5162 -344 -5134
rect -316 -5162 -278 -5134
rect -250 -5162 -212 -5134
rect -184 -5162 -146 -5134
rect -118 -5162 -80 -5134
rect -52 -5162 -14 -5134
rect 14 -5162 52 -5134
rect 80 -5162 118 -5134
rect 146 -5162 184 -5134
rect 212 -5162 250 -5134
rect 278 -5162 316 -5134
rect 344 -5162 382 -5134
rect 410 -5162 448 -5134
rect 476 -5162 514 -5134
rect 542 -5162 580 -5134
rect 608 -5162 646 -5134
rect 674 -5162 712 -5134
rect 740 -5162 745 -5134
rect -745 -5200 745 -5162
rect -745 -5228 -740 -5200
rect -712 -5228 -674 -5200
rect -646 -5228 -608 -5200
rect -580 -5228 -542 -5200
rect -514 -5228 -476 -5200
rect -448 -5228 -410 -5200
rect -382 -5228 -344 -5200
rect -316 -5228 -278 -5200
rect -250 -5228 -212 -5200
rect -184 -5228 -146 -5200
rect -118 -5228 -80 -5200
rect -52 -5228 -14 -5200
rect 14 -5228 52 -5200
rect 80 -5228 118 -5200
rect 146 -5228 184 -5200
rect 212 -5228 250 -5200
rect 278 -5228 316 -5200
rect 344 -5228 382 -5200
rect 410 -5228 448 -5200
rect 476 -5228 514 -5200
rect 542 -5228 580 -5200
rect 608 -5228 646 -5200
rect 674 -5228 712 -5200
rect 740 -5228 745 -5200
rect -745 -5266 745 -5228
rect -745 -5294 -740 -5266
rect -712 -5294 -674 -5266
rect -646 -5294 -608 -5266
rect -580 -5294 -542 -5266
rect -514 -5294 -476 -5266
rect -448 -5294 -410 -5266
rect -382 -5294 -344 -5266
rect -316 -5294 -278 -5266
rect -250 -5294 -212 -5266
rect -184 -5294 -146 -5266
rect -118 -5294 -80 -5266
rect -52 -5294 -14 -5266
rect 14 -5294 52 -5266
rect 80 -5294 118 -5266
rect 146 -5294 184 -5266
rect 212 -5294 250 -5266
rect 278 -5294 316 -5266
rect 344 -5294 382 -5266
rect 410 -5294 448 -5266
rect 476 -5294 514 -5266
rect 542 -5294 580 -5266
rect 608 -5294 646 -5266
rect 674 -5294 712 -5266
rect 740 -5294 745 -5266
rect -745 -5332 745 -5294
rect -745 -5360 -740 -5332
rect -712 -5360 -674 -5332
rect -646 -5360 -608 -5332
rect -580 -5360 -542 -5332
rect -514 -5360 -476 -5332
rect -448 -5360 -410 -5332
rect -382 -5360 -344 -5332
rect -316 -5360 -278 -5332
rect -250 -5360 -212 -5332
rect -184 -5360 -146 -5332
rect -118 -5360 -80 -5332
rect -52 -5360 -14 -5332
rect 14 -5360 52 -5332
rect 80 -5360 118 -5332
rect 146 -5360 184 -5332
rect 212 -5360 250 -5332
rect 278 -5360 316 -5332
rect 344 -5360 382 -5332
rect 410 -5360 448 -5332
rect 476 -5360 514 -5332
rect 542 -5360 580 -5332
rect 608 -5360 646 -5332
rect 674 -5360 712 -5332
rect 740 -5360 745 -5332
rect -745 -5398 745 -5360
rect -745 -5426 -740 -5398
rect -712 -5426 -674 -5398
rect -646 -5426 -608 -5398
rect -580 -5426 -542 -5398
rect -514 -5426 -476 -5398
rect -448 -5426 -410 -5398
rect -382 -5426 -344 -5398
rect -316 -5426 -278 -5398
rect -250 -5426 -212 -5398
rect -184 -5426 -146 -5398
rect -118 -5426 -80 -5398
rect -52 -5426 -14 -5398
rect 14 -5426 52 -5398
rect 80 -5426 118 -5398
rect 146 -5426 184 -5398
rect 212 -5426 250 -5398
rect 278 -5426 316 -5398
rect 344 -5426 382 -5398
rect 410 -5426 448 -5398
rect 476 -5426 514 -5398
rect 542 -5426 580 -5398
rect 608 -5426 646 -5398
rect 674 -5426 712 -5398
rect 740 -5426 745 -5398
rect -745 -5464 745 -5426
rect -745 -5492 -740 -5464
rect -712 -5492 -674 -5464
rect -646 -5492 -608 -5464
rect -580 -5492 -542 -5464
rect -514 -5492 -476 -5464
rect -448 -5492 -410 -5464
rect -382 -5492 -344 -5464
rect -316 -5492 -278 -5464
rect -250 -5492 -212 -5464
rect -184 -5492 -146 -5464
rect -118 -5492 -80 -5464
rect -52 -5492 -14 -5464
rect 14 -5492 52 -5464
rect 80 -5492 118 -5464
rect 146 -5492 184 -5464
rect 212 -5492 250 -5464
rect 278 -5492 316 -5464
rect 344 -5492 382 -5464
rect 410 -5492 448 -5464
rect 476 -5492 514 -5464
rect 542 -5492 580 -5464
rect 608 -5492 646 -5464
rect 674 -5492 712 -5464
rect 740 -5492 745 -5464
rect -745 -5530 745 -5492
rect -745 -5558 -740 -5530
rect -712 -5558 -674 -5530
rect -646 -5558 -608 -5530
rect -580 -5558 -542 -5530
rect -514 -5558 -476 -5530
rect -448 -5558 -410 -5530
rect -382 -5558 -344 -5530
rect -316 -5558 -278 -5530
rect -250 -5558 -212 -5530
rect -184 -5558 -146 -5530
rect -118 -5558 -80 -5530
rect -52 -5558 -14 -5530
rect 14 -5558 52 -5530
rect 80 -5558 118 -5530
rect 146 -5558 184 -5530
rect 212 -5558 250 -5530
rect 278 -5558 316 -5530
rect 344 -5558 382 -5530
rect 410 -5558 448 -5530
rect 476 -5558 514 -5530
rect 542 -5558 580 -5530
rect 608 -5558 646 -5530
rect 674 -5558 712 -5530
rect 740 -5558 745 -5530
rect -745 -5563 745 -5558
<< via3 >>
rect -740 5530 -712 5558
rect -674 5530 -646 5558
rect -608 5530 -580 5558
rect -542 5530 -514 5558
rect -476 5530 -448 5558
rect -410 5530 -382 5558
rect -344 5530 -316 5558
rect -278 5530 -250 5558
rect -212 5530 -184 5558
rect -146 5530 -118 5558
rect -80 5530 -52 5558
rect -14 5530 14 5558
rect 52 5530 80 5558
rect 118 5530 146 5558
rect 184 5530 212 5558
rect 250 5530 278 5558
rect 316 5530 344 5558
rect 382 5530 410 5558
rect 448 5530 476 5558
rect 514 5530 542 5558
rect 580 5530 608 5558
rect 646 5530 674 5558
rect 712 5530 740 5558
rect -740 5464 -712 5492
rect -674 5464 -646 5492
rect -608 5464 -580 5492
rect -542 5464 -514 5492
rect -476 5464 -448 5492
rect -410 5464 -382 5492
rect -344 5464 -316 5492
rect -278 5464 -250 5492
rect -212 5464 -184 5492
rect -146 5464 -118 5492
rect -80 5464 -52 5492
rect -14 5464 14 5492
rect 52 5464 80 5492
rect 118 5464 146 5492
rect 184 5464 212 5492
rect 250 5464 278 5492
rect 316 5464 344 5492
rect 382 5464 410 5492
rect 448 5464 476 5492
rect 514 5464 542 5492
rect 580 5464 608 5492
rect 646 5464 674 5492
rect 712 5464 740 5492
rect -740 5398 -712 5426
rect -674 5398 -646 5426
rect -608 5398 -580 5426
rect -542 5398 -514 5426
rect -476 5398 -448 5426
rect -410 5398 -382 5426
rect -344 5398 -316 5426
rect -278 5398 -250 5426
rect -212 5398 -184 5426
rect -146 5398 -118 5426
rect -80 5398 -52 5426
rect -14 5398 14 5426
rect 52 5398 80 5426
rect 118 5398 146 5426
rect 184 5398 212 5426
rect 250 5398 278 5426
rect 316 5398 344 5426
rect 382 5398 410 5426
rect 448 5398 476 5426
rect 514 5398 542 5426
rect 580 5398 608 5426
rect 646 5398 674 5426
rect 712 5398 740 5426
rect -740 5332 -712 5360
rect -674 5332 -646 5360
rect -608 5332 -580 5360
rect -542 5332 -514 5360
rect -476 5332 -448 5360
rect -410 5332 -382 5360
rect -344 5332 -316 5360
rect -278 5332 -250 5360
rect -212 5332 -184 5360
rect -146 5332 -118 5360
rect -80 5332 -52 5360
rect -14 5332 14 5360
rect 52 5332 80 5360
rect 118 5332 146 5360
rect 184 5332 212 5360
rect 250 5332 278 5360
rect 316 5332 344 5360
rect 382 5332 410 5360
rect 448 5332 476 5360
rect 514 5332 542 5360
rect 580 5332 608 5360
rect 646 5332 674 5360
rect 712 5332 740 5360
rect -740 5266 -712 5294
rect -674 5266 -646 5294
rect -608 5266 -580 5294
rect -542 5266 -514 5294
rect -476 5266 -448 5294
rect -410 5266 -382 5294
rect -344 5266 -316 5294
rect -278 5266 -250 5294
rect -212 5266 -184 5294
rect -146 5266 -118 5294
rect -80 5266 -52 5294
rect -14 5266 14 5294
rect 52 5266 80 5294
rect 118 5266 146 5294
rect 184 5266 212 5294
rect 250 5266 278 5294
rect 316 5266 344 5294
rect 382 5266 410 5294
rect 448 5266 476 5294
rect 514 5266 542 5294
rect 580 5266 608 5294
rect 646 5266 674 5294
rect 712 5266 740 5294
rect -740 5200 -712 5228
rect -674 5200 -646 5228
rect -608 5200 -580 5228
rect -542 5200 -514 5228
rect -476 5200 -448 5228
rect -410 5200 -382 5228
rect -344 5200 -316 5228
rect -278 5200 -250 5228
rect -212 5200 -184 5228
rect -146 5200 -118 5228
rect -80 5200 -52 5228
rect -14 5200 14 5228
rect 52 5200 80 5228
rect 118 5200 146 5228
rect 184 5200 212 5228
rect 250 5200 278 5228
rect 316 5200 344 5228
rect 382 5200 410 5228
rect 448 5200 476 5228
rect 514 5200 542 5228
rect 580 5200 608 5228
rect 646 5200 674 5228
rect 712 5200 740 5228
rect -740 5134 -712 5162
rect -674 5134 -646 5162
rect -608 5134 -580 5162
rect -542 5134 -514 5162
rect -476 5134 -448 5162
rect -410 5134 -382 5162
rect -344 5134 -316 5162
rect -278 5134 -250 5162
rect -212 5134 -184 5162
rect -146 5134 -118 5162
rect -80 5134 -52 5162
rect -14 5134 14 5162
rect 52 5134 80 5162
rect 118 5134 146 5162
rect 184 5134 212 5162
rect 250 5134 278 5162
rect 316 5134 344 5162
rect 382 5134 410 5162
rect 448 5134 476 5162
rect 514 5134 542 5162
rect 580 5134 608 5162
rect 646 5134 674 5162
rect 712 5134 740 5162
rect -740 5068 -712 5096
rect -674 5068 -646 5096
rect -608 5068 -580 5096
rect -542 5068 -514 5096
rect -476 5068 -448 5096
rect -410 5068 -382 5096
rect -344 5068 -316 5096
rect -278 5068 -250 5096
rect -212 5068 -184 5096
rect -146 5068 -118 5096
rect -80 5068 -52 5096
rect -14 5068 14 5096
rect 52 5068 80 5096
rect 118 5068 146 5096
rect 184 5068 212 5096
rect 250 5068 278 5096
rect 316 5068 344 5096
rect 382 5068 410 5096
rect 448 5068 476 5096
rect 514 5068 542 5096
rect 580 5068 608 5096
rect 646 5068 674 5096
rect 712 5068 740 5096
rect -740 5002 -712 5030
rect -674 5002 -646 5030
rect -608 5002 -580 5030
rect -542 5002 -514 5030
rect -476 5002 -448 5030
rect -410 5002 -382 5030
rect -344 5002 -316 5030
rect -278 5002 -250 5030
rect -212 5002 -184 5030
rect -146 5002 -118 5030
rect -80 5002 -52 5030
rect -14 5002 14 5030
rect 52 5002 80 5030
rect 118 5002 146 5030
rect 184 5002 212 5030
rect 250 5002 278 5030
rect 316 5002 344 5030
rect 382 5002 410 5030
rect 448 5002 476 5030
rect 514 5002 542 5030
rect 580 5002 608 5030
rect 646 5002 674 5030
rect 712 5002 740 5030
rect -740 4936 -712 4964
rect -674 4936 -646 4964
rect -608 4936 -580 4964
rect -542 4936 -514 4964
rect -476 4936 -448 4964
rect -410 4936 -382 4964
rect -344 4936 -316 4964
rect -278 4936 -250 4964
rect -212 4936 -184 4964
rect -146 4936 -118 4964
rect -80 4936 -52 4964
rect -14 4936 14 4964
rect 52 4936 80 4964
rect 118 4936 146 4964
rect 184 4936 212 4964
rect 250 4936 278 4964
rect 316 4936 344 4964
rect 382 4936 410 4964
rect 448 4936 476 4964
rect 514 4936 542 4964
rect 580 4936 608 4964
rect 646 4936 674 4964
rect 712 4936 740 4964
rect -740 4870 -712 4898
rect -674 4870 -646 4898
rect -608 4870 -580 4898
rect -542 4870 -514 4898
rect -476 4870 -448 4898
rect -410 4870 -382 4898
rect -344 4870 -316 4898
rect -278 4870 -250 4898
rect -212 4870 -184 4898
rect -146 4870 -118 4898
rect -80 4870 -52 4898
rect -14 4870 14 4898
rect 52 4870 80 4898
rect 118 4870 146 4898
rect 184 4870 212 4898
rect 250 4870 278 4898
rect 316 4870 344 4898
rect 382 4870 410 4898
rect 448 4870 476 4898
rect 514 4870 542 4898
rect 580 4870 608 4898
rect 646 4870 674 4898
rect 712 4870 740 4898
rect -740 4804 -712 4832
rect -674 4804 -646 4832
rect -608 4804 -580 4832
rect -542 4804 -514 4832
rect -476 4804 -448 4832
rect -410 4804 -382 4832
rect -344 4804 -316 4832
rect -278 4804 -250 4832
rect -212 4804 -184 4832
rect -146 4804 -118 4832
rect -80 4804 -52 4832
rect -14 4804 14 4832
rect 52 4804 80 4832
rect 118 4804 146 4832
rect 184 4804 212 4832
rect 250 4804 278 4832
rect 316 4804 344 4832
rect 382 4804 410 4832
rect 448 4804 476 4832
rect 514 4804 542 4832
rect 580 4804 608 4832
rect 646 4804 674 4832
rect 712 4804 740 4832
rect -740 4738 -712 4766
rect -674 4738 -646 4766
rect -608 4738 -580 4766
rect -542 4738 -514 4766
rect -476 4738 -448 4766
rect -410 4738 -382 4766
rect -344 4738 -316 4766
rect -278 4738 -250 4766
rect -212 4738 -184 4766
rect -146 4738 -118 4766
rect -80 4738 -52 4766
rect -14 4738 14 4766
rect 52 4738 80 4766
rect 118 4738 146 4766
rect 184 4738 212 4766
rect 250 4738 278 4766
rect 316 4738 344 4766
rect 382 4738 410 4766
rect 448 4738 476 4766
rect 514 4738 542 4766
rect 580 4738 608 4766
rect 646 4738 674 4766
rect 712 4738 740 4766
rect -740 4672 -712 4700
rect -674 4672 -646 4700
rect -608 4672 -580 4700
rect -542 4672 -514 4700
rect -476 4672 -448 4700
rect -410 4672 -382 4700
rect -344 4672 -316 4700
rect -278 4672 -250 4700
rect -212 4672 -184 4700
rect -146 4672 -118 4700
rect -80 4672 -52 4700
rect -14 4672 14 4700
rect 52 4672 80 4700
rect 118 4672 146 4700
rect 184 4672 212 4700
rect 250 4672 278 4700
rect 316 4672 344 4700
rect 382 4672 410 4700
rect 448 4672 476 4700
rect 514 4672 542 4700
rect 580 4672 608 4700
rect 646 4672 674 4700
rect 712 4672 740 4700
rect -740 4606 -712 4634
rect -674 4606 -646 4634
rect -608 4606 -580 4634
rect -542 4606 -514 4634
rect -476 4606 -448 4634
rect -410 4606 -382 4634
rect -344 4606 -316 4634
rect -278 4606 -250 4634
rect -212 4606 -184 4634
rect -146 4606 -118 4634
rect -80 4606 -52 4634
rect -14 4606 14 4634
rect 52 4606 80 4634
rect 118 4606 146 4634
rect 184 4606 212 4634
rect 250 4606 278 4634
rect 316 4606 344 4634
rect 382 4606 410 4634
rect 448 4606 476 4634
rect 514 4606 542 4634
rect 580 4606 608 4634
rect 646 4606 674 4634
rect 712 4606 740 4634
rect -740 4540 -712 4568
rect -674 4540 -646 4568
rect -608 4540 -580 4568
rect -542 4540 -514 4568
rect -476 4540 -448 4568
rect -410 4540 -382 4568
rect -344 4540 -316 4568
rect -278 4540 -250 4568
rect -212 4540 -184 4568
rect -146 4540 -118 4568
rect -80 4540 -52 4568
rect -14 4540 14 4568
rect 52 4540 80 4568
rect 118 4540 146 4568
rect 184 4540 212 4568
rect 250 4540 278 4568
rect 316 4540 344 4568
rect 382 4540 410 4568
rect 448 4540 476 4568
rect 514 4540 542 4568
rect 580 4540 608 4568
rect 646 4540 674 4568
rect 712 4540 740 4568
rect -740 4474 -712 4502
rect -674 4474 -646 4502
rect -608 4474 -580 4502
rect -542 4474 -514 4502
rect -476 4474 -448 4502
rect -410 4474 -382 4502
rect -344 4474 -316 4502
rect -278 4474 -250 4502
rect -212 4474 -184 4502
rect -146 4474 -118 4502
rect -80 4474 -52 4502
rect -14 4474 14 4502
rect 52 4474 80 4502
rect 118 4474 146 4502
rect 184 4474 212 4502
rect 250 4474 278 4502
rect 316 4474 344 4502
rect 382 4474 410 4502
rect 448 4474 476 4502
rect 514 4474 542 4502
rect 580 4474 608 4502
rect 646 4474 674 4502
rect 712 4474 740 4502
rect -740 4408 -712 4436
rect -674 4408 -646 4436
rect -608 4408 -580 4436
rect -542 4408 -514 4436
rect -476 4408 -448 4436
rect -410 4408 -382 4436
rect -344 4408 -316 4436
rect -278 4408 -250 4436
rect -212 4408 -184 4436
rect -146 4408 -118 4436
rect -80 4408 -52 4436
rect -14 4408 14 4436
rect 52 4408 80 4436
rect 118 4408 146 4436
rect 184 4408 212 4436
rect 250 4408 278 4436
rect 316 4408 344 4436
rect 382 4408 410 4436
rect 448 4408 476 4436
rect 514 4408 542 4436
rect 580 4408 608 4436
rect 646 4408 674 4436
rect 712 4408 740 4436
rect -740 4342 -712 4370
rect -674 4342 -646 4370
rect -608 4342 -580 4370
rect -542 4342 -514 4370
rect -476 4342 -448 4370
rect -410 4342 -382 4370
rect -344 4342 -316 4370
rect -278 4342 -250 4370
rect -212 4342 -184 4370
rect -146 4342 -118 4370
rect -80 4342 -52 4370
rect -14 4342 14 4370
rect 52 4342 80 4370
rect 118 4342 146 4370
rect 184 4342 212 4370
rect 250 4342 278 4370
rect 316 4342 344 4370
rect 382 4342 410 4370
rect 448 4342 476 4370
rect 514 4342 542 4370
rect 580 4342 608 4370
rect 646 4342 674 4370
rect 712 4342 740 4370
rect -740 4276 -712 4304
rect -674 4276 -646 4304
rect -608 4276 -580 4304
rect -542 4276 -514 4304
rect -476 4276 -448 4304
rect -410 4276 -382 4304
rect -344 4276 -316 4304
rect -278 4276 -250 4304
rect -212 4276 -184 4304
rect -146 4276 -118 4304
rect -80 4276 -52 4304
rect -14 4276 14 4304
rect 52 4276 80 4304
rect 118 4276 146 4304
rect 184 4276 212 4304
rect 250 4276 278 4304
rect 316 4276 344 4304
rect 382 4276 410 4304
rect 448 4276 476 4304
rect 514 4276 542 4304
rect 580 4276 608 4304
rect 646 4276 674 4304
rect 712 4276 740 4304
rect -740 4210 -712 4238
rect -674 4210 -646 4238
rect -608 4210 -580 4238
rect -542 4210 -514 4238
rect -476 4210 -448 4238
rect -410 4210 -382 4238
rect -344 4210 -316 4238
rect -278 4210 -250 4238
rect -212 4210 -184 4238
rect -146 4210 -118 4238
rect -80 4210 -52 4238
rect -14 4210 14 4238
rect 52 4210 80 4238
rect 118 4210 146 4238
rect 184 4210 212 4238
rect 250 4210 278 4238
rect 316 4210 344 4238
rect 382 4210 410 4238
rect 448 4210 476 4238
rect 514 4210 542 4238
rect 580 4210 608 4238
rect 646 4210 674 4238
rect 712 4210 740 4238
rect -740 4144 -712 4172
rect -674 4144 -646 4172
rect -608 4144 -580 4172
rect -542 4144 -514 4172
rect -476 4144 -448 4172
rect -410 4144 -382 4172
rect -344 4144 -316 4172
rect -278 4144 -250 4172
rect -212 4144 -184 4172
rect -146 4144 -118 4172
rect -80 4144 -52 4172
rect -14 4144 14 4172
rect 52 4144 80 4172
rect 118 4144 146 4172
rect 184 4144 212 4172
rect 250 4144 278 4172
rect 316 4144 344 4172
rect 382 4144 410 4172
rect 448 4144 476 4172
rect 514 4144 542 4172
rect 580 4144 608 4172
rect 646 4144 674 4172
rect 712 4144 740 4172
rect -740 4078 -712 4106
rect -674 4078 -646 4106
rect -608 4078 -580 4106
rect -542 4078 -514 4106
rect -476 4078 -448 4106
rect -410 4078 -382 4106
rect -344 4078 -316 4106
rect -278 4078 -250 4106
rect -212 4078 -184 4106
rect -146 4078 -118 4106
rect -80 4078 -52 4106
rect -14 4078 14 4106
rect 52 4078 80 4106
rect 118 4078 146 4106
rect 184 4078 212 4106
rect 250 4078 278 4106
rect 316 4078 344 4106
rect 382 4078 410 4106
rect 448 4078 476 4106
rect 514 4078 542 4106
rect 580 4078 608 4106
rect 646 4078 674 4106
rect 712 4078 740 4106
rect -740 4012 -712 4040
rect -674 4012 -646 4040
rect -608 4012 -580 4040
rect -542 4012 -514 4040
rect -476 4012 -448 4040
rect -410 4012 -382 4040
rect -344 4012 -316 4040
rect -278 4012 -250 4040
rect -212 4012 -184 4040
rect -146 4012 -118 4040
rect -80 4012 -52 4040
rect -14 4012 14 4040
rect 52 4012 80 4040
rect 118 4012 146 4040
rect 184 4012 212 4040
rect 250 4012 278 4040
rect 316 4012 344 4040
rect 382 4012 410 4040
rect 448 4012 476 4040
rect 514 4012 542 4040
rect 580 4012 608 4040
rect 646 4012 674 4040
rect 712 4012 740 4040
rect -740 3946 -712 3974
rect -674 3946 -646 3974
rect -608 3946 -580 3974
rect -542 3946 -514 3974
rect -476 3946 -448 3974
rect -410 3946 -382 3974
rect -344 3946 -316 3974
rect -278 3946 -250 3974
rect -212 3946 -184 3974
rect -146 3946 -118 3974
rect -80 3946 -52 3974
rect -14 3946 14 3974
rect 52 3946 80 3974
rect 118 3946 146 3974
rect 184 3946 212 3974
rect 250 3946 278 3974
rect 316 3946 344 3974
rect 382 3946 410 3974
rect 448 3946 476 3974
rect 514 3946 542 3974
rect 580 3946 608 3974
rect 646 3946 674 3974
rect 712 3946 740 3974
rect -740 3880 -712 3908
rect -674 3880 -646 3908
rect -608 3880 -580 3908
rect -542 3880 -514 3908
rect -476 3880 -448 3908
rect -410 3880 -382 3908
rect -344 3880 -316 3908
rect -278 3880 -250 3908
rect -212 3880 -184 3908
rect -146 3880 -118 3908
rect -80 3880 -52 3908
rect -14 3880 14 3908
rect 52 3880 80 3908
rect 118 3880 146 3908
rect 184 3880 212 3908
rect 250 3880 278 3908
rect 316 3880 344 3908
rect 382 3880 410 3908
rect 448 3880 476 3908
rect 514 3880 542 3908
rect 580 3880 608 3908
rect 646 3880 674 3908
rect 712 3880 740 3908
rect -740 3814 -712 3842
rect -674 3814 -646 3842
rect -608 3814 -580 3842
rect -542 3814 -514 3842
rect -476 3814 -448 3842
rect -410 3814 -382 3842
rect -344 3814 -316 3842
rect -278 3814 -250 3842
rect -212 3814 -184 3842
rect -146 3814 -118 3842
rect -80 3814 -52 3842
rect -14 3814 14 3842
rect 52 3814 80 3842
rect 118 3814 146 3842
rect 184 3814 212 3842
rect 250 3814 278 3842
rect 316 3814 344 3842
rect 382 3814 410 3842
rect 448 3814 476 3842
rect 514 3814 542 3842
rect 580 3814 608 3842
rect 646 3814 674 3842
rect 712 3814 740 3842
rect -740 3748 -712 3776
rect -674 3748 -646 3776
rect -608 3748 -580 3776
rect -542 3748 -514 3776
rect -476 3748 -448 3776
rect -410 3748 -382 3776
rect -344 3748 -316 3776
rect -278 3748 -250 3776
rect -212 3748 -184 3776
rect -146 3748 -118 3776
rect -80 3748 -52 3776
rect -14 3748 14 3776
rect 52 3748 80 3776
rect 118 3748 146 3776
rect 184 3748 212 3776
rect 250 3748 278 3776
rect 316 3748 344 3776
rect 382 3748 410 3776
rect 448 3748 476 3776
rect 514 3748 542 3776
rect 580 3748 608 3776
rect 646 3748 674 3776
rect 712 3748 740 3776
rect -740 3682 -712 3710
rect -674 3682 -646 3710
rect -608 3682 -580 3710
rect -542 3682 -514 3710
rect -476 3682 -448 3710
rect -410 3682 -382 3710
rect -344 3682 -316 3710
rect -278 3682 -250 3710
rect -212 3682 -184 3710
rect -146 3682 -118 3710
rect -80 3682 -52 3710
rect -14 3682 14 3710
rect 52 3682 80 3710
rect 118 3682 146 3710
rect 184 3682 212 3710
rect 250 3682 278 3710
rect 316 3682 344 3710
rect 382 3682 410 3710
rect 448 3682 476 3710
rect 514 3682 542 3710
rect 580 3682 608 3710
rect 646 3682 674 3710
rect 712 3682 740 3710
rect -740 3616 -712 3644
rect -674 3616 -646 3644
rect -608 3616 -580 3644
rect -542 3616 -514 3644
rect -476 3616 -448 3644
rect -410 3616 -382 3644
rect -344 3616 -316 3644
rect -278 3616 -250 3644
rect -212 3616 -184 3644
rect -146 3616 -118 3644
rect -80 3616 -52 3644
rect -14 3616 14 3644
rect 52 3616 80 3644
rect 118 3616 146 3644
rect 184 3616 212 3644
rect 250 3616 278 3644
rect 316 3616 344 3644
rect 382 3616 410 3644
rect 448 3616 476 3644
rect 514 3616 542 3644
rect 580 3616 608 3644
rect 646 3616 674 3644
rect 712 3616 740 3644
rect -740 3550 -712 3578
rect -674 3550 -646 3578
rect -608 3550 -580 3578
rect -542 3550 -514 3578
rect -476 3550 -448 3578
rect -410 3550 -382 3578
rect -344 3550 -316 3578
rect -278 3550 -250 3578
rect -212 3550 -184 3578
rect -146 3550 -118 3578
rect -80 3550 -52 3578
rect -14 3550 14 3578
rect 52 3550 80 3578
rect 118 3550 146 3578
rect 184 3550 212 3578
rect 250 3550 278 3578
rect 316 3550 344 3578
rect 382 3550 410 3578
rect 448 3550 476 3578
rect 514 3550 542 3578
rect 580 3550 608 3578
rect 646 3550 674 3578
rect 712 3550 740 3578
rect -740 3484 -712 3512
rect -674 3484 -646 3512
rect -608 3484 -580 3512
rect -542 3484 -514 3512
rect -476 3484 -448 3512
rect -410 3484 -382 3512
rect -344 3484 -316 3512
rect -278 3484 -250 3512
rect -212 3484 -184 3512
rect -146 3484 -118 3512
rect -80 3484 -52 3512
rect -14 3484 14 3512
rect 52 3484 80 3512
rect 118 3484 146 3512
rect 184 3484 212 3512
rect 250 3484 278 3512
rect 316 3484 344 3512
rect 382 3484 410 3512
rect 448 3484 476 3512
rect 514 3484 542 3512
rect 580 3484 608 3512
rect 646 3484 674 3512
rect 712 3484 740 3512
rect -740 3418 -712 3446
rect -674 3418 -646 3446
rect -608 3418 -580 3446
rect -542 3418 -514 3446
rect -476 3418 -448 3446
rect -410 3418 -382 3446
rect -344 3418 -316 3446
rect -278 3418 -250 3446
rect -212 3418 -184 3446
rect -146 3418 -118 3446
rect -80 3418 -52 3446
rect -14 3418 14 3446
rect 52 3418 80 3446
rect 118 3418 146 3446
rect 184 3418 212 3446
rect 250 3418 278 3446
rect 316 3418 344 3446
rect 382 3418 410 3446
rect 448 3418 476 3446
rect 514 3418 542 3446
rect 580 3418 608 3446
rect 646 3418 674 3446
rect 712 3418 740 3446
rect -740 3352 -712 3380
rect -674 3352 -646 3380
rect -608 3352 -580 3380
rect -542 3352 -514 3380
rect -476 3352 -448 3380
rect -410 3352 -382 3380
rect -344 3352 -316 3380
rect -278 3352 -250 3380
rect -212 3352 -184 3380
rect -146 3352 -118 3380
rect -80 3352 -52 3380
rect -14 3352 14 3380
rect 52 3352 80 3380
rect 118 3352 146 3380
rect 184 3352 212 3380
rect 250 3352 278 3380
rect 316 3352 344 3380
rect 382 3352 410 3380
rect 448 3352 476 3380
rect 514 3352 542 3380
rect 580 3352 608 3380
rect 646 3352 674 3380
rect 712 3352 740 3380
rect -740 3286 -712 3314
rect -674 3286 -646 3314
rect -608 3286 -580 3314
rect -542 3286 -514 3314
rect -476 3286 -448 3314
rect -410 3286 -382 3314
rect -344 3286 -316 3314
rect -278 3286 -250 3314
rect -212 3286 -184 3314
rect -146 3286 -118 3314
rect -80 3286 -52 3314
rect -14 3286 14 3314
rect 52 3286 80 3314
rect 118 3286 146 3314
rect 184 3286 212 3314
rect 250 3286 278 3314
rect 316 3286 344 3314
rect 382 3286 410 3314
rect 448 3286 476 3314
rect 514 3286 542 3314
rect 580 3286 608 3314
rect 646 3286 674 3314
rect 712 3286 740 3314
rect -740 3220 -712 3248
rect -674 3220 -646 3248
rect -608 3220 -580 3248
rect -542 3220 -514 3248
rect -476 3220 -448 3248
rect -410 3220 -382 3248
rect -344 3220 -316 3248
rect -278 3220 -250 3248
rect -212 3220 -184 3248
rect -146 3220 -118 3248
rect -80 3220 -52 3248
rect -14 3220 14 3248
rect 52 3220 80 3248
rect 118 3220 146 3248
rect 184 3220 212 3248
rect 250 3220 278 3248
rect 316 3220 344 3248
rect 382 3220 410 3248
rect 448 3220 476 3248
rect 514 3220 542 3248
rect 580 3220 608 3248
rect 646 3220 674 3248
rect 712 3220 740 3248
rect -740 3154 -712 3182
rect -674 3154 -646 3182
rect -608 3154 -580 3182
rect -542 3154 -514 3182
rect -476 3154 -448 3182
rect -410 3154 -382 3182
rect -344 3154 -316 3182
rect -278 3154 -250 3182
rect -212 3154 -184 3182
rect -146 3154 -118 3182
rect -80 3154 -52 3182
rect -14 3154 14 3182
rect 52 3154 80 3182
rect 118 3154 146 3182
rect 184 3154 212 3182
rect 250 3154 278 3182
rect 316 3154 344 3182
rect 382 3154 410 3182
rect 448 3154 476 3182
rect 514 3154 542 3182
rect 580 3154 608 3182
rect 646 3154 674 3182
rect 712 3154 740 3182
rect -740 3088 -712 3116
rect -674 3088 -646 3116
rect -608 3088 -580 3116
rect -542 3088 -514 3116
rect -476 3088 -448 3116
rect -410 3088 -382 3116
rect -344 3088 -316 3116
rect -278 3088 -250 3116
rect -212 3088 -184 3116
rect -146 3088 -118 3116
rect -80 3088 -52 3116
rect -14 3088 14 3116
rect 52 3088 80 3116
rect 118 3088 146 3116
rect 184 3088 212 3116
rect 250 3088 278 3116
rect 316 3088 344 3116
rect 382 3088 410 3116
rect 448 3088 476 3116
rect 514 3088 542 3116
rect 580 3088 608 3116
rect 646 3088 674 3116
rect 712 3088 740 3116
rect -740 3022 -712 3050
rect -674 3022 -646 3050
rect -608 3022 -580 3050
rect -542 3022 -514 3050
rect -476 3022 -448 3050
rect -410 3022 -382 3050
rect -344 3022 -316 3050
rect -278 3022 -250 3050
rect -212 3022 -184 3050
rect -146 3022 -118 3050
rect -80 3022 -52 3050
rect -14 3022 14 3050
rect 52 3022 80 3050
rect 118 3022 146 3050
rect 184 3022 212 3050
rect 250 3022 278 3050
rect 316 3022 344 3050
rect 382 3022 410 3050
rect 448 3022 476 3050
rect 514 3022 542 3050
rect 580 3022 608 3050
rect 646 3022 674 3050
rect 712 3022 740 3050
rect -740 2956 -712 2984
rect -674 2956 -646 2984
rect -608 2956 -580 2984
rect -542 2956 -514 2984
rect -476 2956 -448 2984
rect -410 2956 -382 2984
rect -344 2956 -316 2984
rect -278 2956 -250 2984
rect -212 2956 -184 2984
rect -146 2956 -118 2984
rect -80 2956 -52 2984
rect -14 2956 14 2984
rect 52 2956 80 2984
rect 118 2956 146 2984
rect 184 2956 212 2984
rect 250 2956 278 2984
rect 316 2956 344 2984
rect 382 2956 410 2984
rect 448 2956 476 2984
rect 514 2956 542 2984
rect 580 2956 608 2984
rect 646 2956 674 2984
rect 712 2956 740 2984
rect -740 2890 -712 2918
rect -674 2890 -646 2918
rect -608 2890 -580 2918
rect -542 2890 -514 2918
rect -476 2890 -448 2918
rect -410 2890 -382 2918
rect -344 2890 -316 2918
rect -278 2890 -250 2918
rect -212 2890 -184 2918
rect -146 2890 -118 2918
rect -80 2890 -52 2918
rect -14 2890 14 2918
rect 52 2890 80 2918
rect 118 2890 146 2918
rect 184 2890 212 2918
rect 250 2890 278 2918
rect 316 2890 344 2918
rect 382 2890 410 2918
rect 448 2890 476 2918
rect 514 2890 542 2918
rect 580 2890 608 2918
rect 646 2890 674 2918
rect 712 2890 740 2918
rect -740 2824 -712 2852
rect -674 2824 -646 2852
rect -608 2824 -580 2852
rect -542 2824 -514 2852
rect -476 2824 -448 2852
rect -410 2824 -382 2852
rect -344 2824 -316 2852
rect -278 2824 -250 2852
rect -212 2824 -184 2852
rect -146 2824 -118 2852
rect -80 2824 -52 2852
rect -14 2824 14 2852
rect 52 2824 80 2852
rect 118 2824 146 2852
rect 184 2824 212 2852
rect 250 2824 278 2852
rect 316 2824 344 2852
rect 382 2824 410 2852
rect 448 2824 476 2852
rect 514 2824 542 2852
rect 580 2824 608 2852
rect 646 2824 674 2852
rect 712 2824 740 2852
rect -740 2758 -712 2786
rect -674 2758 -646 2786
rect -608 2758 -580 2786
rect -542 2758 -514 2786
rect -476 2758 -448 2786
rect -410 2758 -382 2786
rect -344 2758 -316 2786
rect -278 2758 -250 2786
rect -212 2758 -184 2786
rect -146 2758 -118 2786
rect -80 2758 -52 2786
rect -14 2758 14 2786
rect 52 2758 80 2786
rect 118 2758 146 2786
rect 184 2758 212 2786
rect 250 2758 278 2786
rect 316 2758 344 2786
rect 382 2758 410 2786
rect 448 2758 476 2786
rect 514 2758 542 2786
rect 580 2758 608 2786
rect 646 2758 674 2786
rect 712 2758 740 2786
rect -740 2692 -712 2720
rect -674 2692 -646 2720
rect -608 2692 -580 2720
rect -542 2692 -514 2720
rect -476 2692 -448 2720
rect -410 2692 -382 2720
rect -344 2692 -316 2720
rect -278 2692 -250 2720
rect -212 2692 -184 2720
rect -146 2692 -118 2720
rect -80 2692 -52 2720
rect -14 2692 14 2720
rect 52 2692 80 2720
rect 118 2692 146 2720
rect 184 2692 212 2720
rect 250 2692 278 2720
rect 316 2692 344 2720
rect 382 2692 410 2720
rect 448 2692 476 2720
rect 514 2692 542 2720
rect 580 2692 608 2720
rect 646 2692 674 2720
rect 712 2692 740 2720
rect -740 2626 -712 2654
rect -674 2626 -646 2654
rect -608 2626 -580 2654
rect -542 2626 -514 2654
rect -476 2626 -448 2654
rect -410 2626 -382 2654
rect -344 2626 -316 2654
rect -278 2626 -250 2654
rect -212 2626 -184 2654
rect -146 2626 -118 2654
rect -80 2626 -52 2654
rect -14 2626 14 2654
rect 52 2626 80 2654
rect 118 2626 146 2654
rect 184 2626 212 2654
rect 250 2626 278 2654
rect 316 2626 344 2654
rect 382 2626 410 2654
rect 448 2626 476 2654
rect 514 2626 542 2654
rect 580 2626 608 2654
rect 646 2626 674 2654
rect 712 2626 740 2654
rect -740 2560 -712 2588
rect -674 2560 -646 2588
rect -608 2560 -580 2588
rect -542 2560 -514 2588
rect -476 2560 -448 2588
rect -410 2560 -382 2588
rect -344 2560 -316 2588
rect -278 2560 -250 2588
rect -212 2560 -184 2588
rect -146 2560 -118 2588
rect -80 2560 -52 2588
rect -14 2560 14 2588
rect 52 2560 80 2588
rect 118 2560 146 2588
rect 184 2560 212 2588
rect 250 2560 278 2588
rect 316 2560 344 2588
rect 382 2560 410 2588
rect 448 2560 476 2588
rect 514 2560 542 2588
rect 580 2560 608 2588
rect 646 2560 674 2588
rect 712 2560 740 2588
rect -740 2494 -712 2522
rect -674 2494 -646 2522
rect -608 2494 -580 2522
rect -542 2494 -514 2522
rect -476 2494 -448 2522
rect -410 2494 -382 2522
rect -344 2494 -316 2522
rect -278 2494 -250 2522
rect -212 2494 -184 2522
rect -146 2494 -118 2522
rect -80 2494 -52 2522
rect -14 2494 14 2522
rect 52 2494 80 2522
rect 118 2494 146 2522
rect 184 2494 212 2522
rect 250 2494 278 2522
rect 316 2494 344 2522
rect 382 2494 410 2522
rect 448 2494 476 2522
rect 514 2494 542 2522
rect 580 2494 608 2522
rect 646 2494 674 2522
rect 712 2494 740 2522
rect -740 2428 -712 2456
rect -674 2428 -646 2456
rect -608 2428 -580 2456
rect -542 2428 -514 2456
rect -476 2428 -448 2456
rect -410 2428 -382 2456
rect -344 2428 -316 2456
rect -278 2428 -250 2456
rect -212 2428 -184 2456
rect -146 2428 -118 2456
rect -80 2428 -52 2456
rect -14 2428 14 2456
rect 52 2428 80 2456
rect 118 2428 146 2456
rect 184 2428 212 2456
rect 250 2428 278 2456
rect 316 2428 344 2456
rect 382 2428 410 2456
rect 448 2428 476 2456
rect 514 2428 542 2456
rect 580 2428 608 2456
rect 646 2428 674 2456
rect 712 2428 740 2456
rect -740 2362 -712 2390
rect -674 2362 -646 2390
rect -608 2362 -580 2390
rect -542 2362 -514 2390
rect -476 2362 -448 2390
rect -410 2362 -382 2390
rect -344 2362 -316 2390
rect -278 2362 -250 2390
rect -212 2362 -184 2390
rect -146 2362 -118 2390
rect -80 2362 -52 2390
rect -14 2362 14 2390
rect 52 2362 80 2390
rect 118 2362 146 2390
rect 184 2362 212 2390
rect 250 2362 278 2390
rect 316 2362 344 2390
rect 382 2362 410 2390
rect 448 2362 476 2390
rect 514 2362 542 2390
rect 580 2362 608 2390
rect 646 2362 674 2390
rect 712 2362 740 2390
rect -740 2296 -712 2324
rect -674 2296 -646 2324
rect -608 2296 -580 2324
rect -542 2296 -514 2324
rect -476 2296 -448 2324
rect -410 2296 -382 2324
rect -344 2296 -316 2324
rect -278 2296 -250 2324
rect -212 2296 -184 2324
rect -146 2296 -118 2324
rect -80 2296 -52 2324
rect -14 2296 14 2324
rect 52 2296 80 2324
rect 118 2296 146 2324
rect 184 2296 212 2324
rect 250 2296 278 2324
rect 316 2296 344 2324
rect 382 2296 410 2324
rect 448 2296 476 2324
rect 514 2296 542 2324
rect 580 2296 608 2324
rect 646 2296 674 2324
rect 712 2296 740 2324
rect -740 2230 -712 2258
rect -674 2230 -646 2258
rect -608 2230 -580 2258
rect -542 2230 -514 2258
rect -476 2230 -448 2258
rect -410 2230 -382 2258
rect -344 2230 -316 2258
rect -278 2230 -250 2258
rect -212 2230 -184 2258
rect -146 2230 -118 2258
rect -80 2230 -52 2258
rect -14 2230 14 2258
rect 52 2230 80 2258
rect 118 2230 146 2258
rect 184 2230 212 2258
rect 250 2230 278 2258
rect 316 2230 344 2258
rect 382 2230 410 2258
rect 448 2230 476 2258
rect 514 2230 542 2258
rect 580 2230 608 2258
rect 646 2230 674 2258
rect 712 2230 740 2258
rect -740 2164 -712 2192
rect -674 2164 -646 2192
rect -608 2164 -580 2192
rect -542 2164 -514 2192
rect -476 2164 -448 2192
rect -410 2164 -382 2192
rect -344 2164 -316 2192
rect -278 2164 -250 2192
rect -212 2164 -184 2192
rect -146 2164 -118 2192
rect -80 2164 -52 2192
rect -14 2164 14 2192
rect 52 2164 80 2192
rect 118 2164 146 2192
rect 184 2164 212 2192
rect 250 2164 278 2192
rect 316 2164 344 2192
rect 382 2164 410 2192
rect 448 2164 476 2192
rect 514 2164 542 2192
rect 580 2164 608 2192
rect 646 2164 674 2192
rect 712 2164 740 2192
rect -740 2098 -712 2126
rect -674 2098 -646 2126
rect -608 2098 -580 2126
rect -542 2098 -514 2126
rect -476 2098 -448 2126
rect -410 2098 -382 2126
rect -344 2098 -316 2126
rect -278 2098 -250 2126
rect -212 2098 -184 2126
rect -146 2098 -118 2126
rect -80 2098 -52 2126
rect -14 2098 14 2126
rect 52 2098 80 2126
rect 118 2098 146 2126
rect 184 2098 212 2126
rect 250 2098 278 2126
rect 316 2098 344 2126
rect 382 2098 410 2126
rect 448 2098 476 2126
rect 514 2098 542 2126
rect 580 2098 608 2126
rect 646 2098 674 2126
rect 712 2098 740 2126
rect -740 2032 -712 2060
rect -674 2032 -646 2060
rect -608 2032 -580 2060
rect -542 2032 -514 2060
rect -476 2032 -448 2060
rect -410 2032 -382 2060
rect -344 2032 -316 2060
rect -278 2032 -250 2060
rect -212 2032 -184 2060
rect -146 2032 -118 2060
rect -80 2032 -52 2060
rect -14 2032 14 2060
rect 52 2032 80 2060
rect 118 2032 146 2060
rect 184 2032 212 2060
rect 250 2032 278 2060
rect 316 2032 344 2060
rect 382 2032 410 2060
rect 448 2032 476 2060
rect 514 2032 542 2060
rect 580 2032 608 2060
rect 646 2032 674 2060
rect 712 2032 740 2060
rect -740 1966 -712 1994
rect -674 1966 -646 1994
rect -608 1966 -580 1994
rect -542 1966 -514 1994
rect -476 1966 -448 1994
rect -410 1966 -382 1994
rect -344 1966 -316 1994
rect -278 1966 -250 1994
rect -212 1966 -184 1994
rect -146 1966 -118 1994
rect -80 1966 -52 1994
rect -14 1966 14 1994
rect 52 1966 80 1994
rect 118 1966 146 1994
rect 184 1966 212 1994
rect 250 1966 278 1994
rect 316 1966 344 1994
rect 382 1966 410 1994
rect 448 1966 476 1994
rect 514 1966 542 1994
rect 580 1966 608 1994
rect 646 1966 674 1994
rect 712 1966 740 1994
rect -740 1900 -712 1928
rect -674 1900 -646 1928
rect -608 1900 -580 1928
rect -542 1900 -514 1928
rect -476 1900 -448 1928
rect -410 1900 -382 1928
rect -344 1900 -316 1928
rect -278 1900 -250 1928
rect -212 1900 -184 1928
rect -146 1900 -118 1928
rect -80 1900 -52 1928
rect -14 1900 14 1928
rect 52 1900 80 1928
rect 118 1900 146 1928
rect 184 1900 212 1928
rect 250 1900 278 1928
rect 316 1900 344 1928
rect 382 1900 410 1928
rect 448 1900 476 1928
rect 514 1900 542 1928
rect 580 1900 608 1928
rect 646 1900 674 1928
rect 712 1900 740 1928
rect -740 1834 -712 1862
rect -674 1834 -646 1862
rect -608 1834 -580 1862
rect -542 1834 -514 1862
rect -476 1834 -448 1862
rect -410 1834 -382 1862
rect -344 1834 -316 1862
rect -278 1834 -250 1862
rect -212 1834 -184 1862
rect -146 1834 -118 1862
rect -80 1834 -52 1862
rect -14 1834 14 1862
rect 52 1834 80 1862
rect 118 1834 146 1862
rect 184 1834 212 1862
rect 250 1834 278 1862
rect 316 1834 344 1862
rect 382 1834 410 1862
rect 448 1834 476 1862
rect 514 1834 542 1862
rect 580 1834 608 1862
rect 646 1834 674 1862
rect 712 1834 740 1862
rect -740 1768 -712 1796
rect -674 1768 -646 1796
rect -608 1768 -580 1796
rect -542 1768 -514 1796
rect -476 1768 -448 1796
rect -410 1768 -382 1796
rect -344 1768 -316 1796
rect -278 1768 -250 1796
rect -212 1768 -184 1796
rect -146 1768 -118 1796
rect -80 1768 -52 1796
rect -14 1768 14 1796
rect 52 1768 80 1796
rect 118 1768 146 1796
rect 184 1768 212 1796
rect 250 1768 278 1796
rect 316 1768 344 1796
rect 382 1768 410 1796
rect 448 1768 476 1796
rect 514 1768 542 1796
rect 580 1768 608 1796
rect 646 1768 674 1796
rect 712 1768 740 1796
rect -740 1702 -712 1730
rect -674 1702 -646 1730
rect -608 1702 -580 1730
rect -542 1702 -514 1730
rect -476 1702 -448 1730
rect -410 1702 -382 1730
rect -344 1702 -316 1730
rect -278 1702 -250 1730
rect -212 1702 -184 1730
rect -146 1702 -118 1730
rect -80 1702 -52 1730
rect -14 1702 14 1730
rect 52 1702 80 1730
rect 118 1702 146 1730
rect 184 1702 212 1730
rect 250 1702 278 1730
rect 316 1702 344 1730
rect 382 1702 410 1730
rect 448 1702 476 1730
rect 514 1702 542 1730
rect 580 1702 608 1730
rect 646 1702 674 1730
rect 712 1702 740 1730
rect -740 1636 -712 1664
rect -674 1636 -646 1664
rect -608 1636 -580 1664
rect -542 1636 -514 1664
rect -476 1636 -448 1664
rect -410 1636 -382 1664
rect -344 1636 -316 1664
rect -278 1636 -250 1664
rect -212 1636 -184 1664
rect -146 1636 -118 1664
rect -80 1636 -52 1664
rect -14 1636 14 1664
rect 52 1636 80 1664
rect 118 1636 146 1664
rect 184 1636 212 1664
rect 250 1636 278 1664
rect 316 1636 344 1664
rect 382 1636 410 1664
rect 448 1636 476 1664
rect 514 1636 542 1664
rect 580 1636 608 1664
rect 646 1636 674 1664
rect 712 1636 740 1664
rect -740 1570 -712 1598
rect -674 1570 -646 1598
rect -608 1570 -580 1598
rect -542 1570 -514 1598
rect -476 1570 -448 1598
rect -410 1570 -382 1598
rect -344 1570 -316 1598
rect -278 1570 -250 1598
rect -212 1570 -184 1598
rect -146 1570 -118 1598
rect -80 1570 -52 1598
rect -14 1570 14 1598
rect 52 1570 80 1598
rect 118 1570 146 1598
rect 184 1570 212 1598
rect 250 1570 278 1598
rect 316 1570 344 1598
rect 382 1570 410 1598
rect 448 1570 476 1598
rect 514 1570 542 1598
rect 580 1570 608 1598
rect 646 1570 674 1598
rect 712 1570 740 1598
rect -740 1504 -712 1532
rect -674 1504 -646 1532
rect -608 1504 -580 1532
rect -542 1504 -514 1532
rect -476 1504 -448 1532
rect -410 1504 -382 1532
rect -344 1504 -316 1532
rect -278 1504 -250 1532
rect -212 1504 -184 1532
rect -146 1504 -118 1532
rect -80 1504 -52 1532
rect -14 1504 14 1532
rect 52 1504 80 1532
rect 118 1504 146 1532
rect 184 1504 212 1532
rect 250 1504 278 1532
rect 316 1504 344 1532
rect 382 1504 410 1532
rect 448 1504 476 1532
rect 514 1504 542 1532
rect 580 1504 608 1532
rect 646 1504 674 1532
rect 712 1504 740 1532
rect -740 1438 -712 1466
rect -674 1438 -646 1466
rect -608 1438 -580 1466
rect -542 1438 -514 1466
rect -476 1438 -448 1466
rect -410 1438 -382 1466
rect -344 1438 -316 1466
rect -278 1438 -250 1466
rect -212 1438 -184 1466
rect -146 1438 -118 1466
rect -80 1438 -52 1466
rect -14 1438 14 1466
rect 52 1438 80 1466
rect 118 1438 146 1466
rect 184 1438 212 1466
rect 250 1438 278 1466
rect 316 1438 344 1466
rect 382 1438 410 1466
rect 448 1438 476 1466
rect 514 1438 542 1466
rect 580 1438 608 1466
rect 646 1438 674 1466
rect 712 1438 740 1466
rect -740 1372 -712 1400
rect -674 1372 -646 1400
rect -608 1372 -580 1400
rect -542 1372 -514 1400
rect -476 1372 -448 1400
rect -410 1372 -382 1400
rect -344 1372 -316 1400
rect -278 1372 -250 1400
rect -212 1372 -184 1400
rect -146 1372 -118 1400
rect -80 1372 -52 1400
rect -14 1372 14 1400
rect 52 1372 80 1400
rect 118 1372 146 1400
rect 184 1372 212 1400
rect 250 1372 278 1400
rect 316 1372 344 1400
rect 382 1372 410 1400
rect 448 1372 476 1400
rect 514 1372 542 1400
rect 580 1372 608 1400
rect 646 1372 674 1400
rect 712 1372 740 1400
rect -740 1306 -712 1334
rect -674 1306 -646 1334
rect -608 1306 -580 1334
rect -542 1306 -514 1334
rect -476 1306 -448 1334
rect -410 1306 -382 1334
rect -344 1306 -316 1334
rect -278 1306 -250 1334
rect -212 1306 -184 1334
rect -146 1306 -118 1334
rect -80 1306 -52 1334
rect -14 1306 14 1334
rect 52 1306 80 1334
rect 118 1306 146 1334
rect 184 1306 212 1334
rect 250 1306 278 1334
rect 316 1306 344 1334
rect 382 1306 410 1334
rect 448 1306 476 1334
rect 514 1306 542 1334
rect 580 1306 608 1334
rect 646 1306 674 1334
rect 712 1306 740 1334
rect -740 1240 -712 1268
rect -674 1240 -646 1268
rect -608 1240 -580 1268
rect -542 1240 -514 1268
rect -476 1240 -448 1268
rect -410 1240 -382 1268
rect -344 1240 -316 1268
rect -278 1240 -250 1268
rect -212 1240 -184 1268
rect -146 1240 -118 1268
rect -80 1240 -52 1268
rect -14 1240 14 1268
rect 52 1240 80 1268
rect 118 1240 146 1268
rect 184 1240 212 1268
rect 250 1240 278 1268
rect 316 1240 344 1268
rect 382 1240 410 1268
rect 448 1240 476 1268
rect 514 1240 542 1268
rect 580 1240 608 1268
rect 646 1240 674 1268
rect 712 1240 740 1268
rect -740 1174 -712 1202
rect -674 1174 -646 1202
rect -608 1174 -580 1202
rect -542 1174 -514 1202
rect -476 1174 -448 1202
rect -410 1174 -382 1202
rect -344 1174 -316 1202
rect -278 1174 -250 1202
rect -212 1174 -184 1202
rect -146 1174 -118 1202
rect -80 1174 -52 1202
rect -14 1174 14 1202
rect 52 1174 80 1202
rect 118 1174 146 1202
rect 184 1174 212 1202
rect 250 1174 278 1202
rect 316 1174 344 1202
rect 382 1174 410 1202
rect 448 1174 476 1202
rect 514 1174 542 1202
rect 580 1174 608 1202
rect 646 1174 674 1202
rect 712 1174 740 1202
rect -740 1108 -712 1136
rect -674 1108 -646 1136
rect -608 1108 -580 1136
rect -542 1108 -514 1136
rect -476 1108 -448 1136
rect -410 1108 -382 1136
rect -344 1108 -316 1136
rect -278 1108 -250 1136
rect -212 1108 -184 1136
rect -146 1108 -118 1136
rect -80 1108 -52 1136
rect -14 1108 14 1136
rect 52 1108 80 1136
rect 118 1108 146 1136
rect 184 1108 212 1136
rect 250 1108 278 1136
rect 316 1108 344 1136
rect 382 1108 410 1136
rect 448 1108 476 1136
rect 514 1108 542 1136
rect 580 1108 608 1136
rect 646 1108 674 1136
rect 712 1108 740 1136
rect -740 1042 -712 1070
rect -674 1042 -646 1070
rect -608 1042 -580 1070
rect -542 1042 -514 1070
rect -476 1042 -448 1070
rect -410 1042 -382 1070
rect -344 1042 -316 1070
rect -278 1042 -250 1070
rect -212 1042 -184 1070
rect -146 1042 -118 1070
rect -80 1042 -52 1070
rect -14 1042 14 1070
rect 52 1042 80 1070
rect 118 1042 146 1070
rect 184 1042 212 1070
rect 250 1042 278 1070
rect 316 1042 344 1070
rect 382 1042 410 1070
rect 448 1042 476 1070
rect 514 1042 542 1070
rect 580 1042 608 1070
rect 646 1042 674 1070
rect 712 1042 740 1070
rect -740 976 -712 1004
rect -674 976 -646 1004
rect -608 976 -580 1004
rect -542 976 -514 1004
rect -476 976 -448 1004
rect -410 976 -382 1004
rect -344 976 -316 1004
rect -278 976 -250 1004
rect -212 976 -184 1004
rect -146 976 -118 1004
rect -80 976 -52 1004
rect -14 976 14 1004
rect 52 976 80 1004
rect 118 976 146 1004
rect 184 976 212 1004
rect 250 976 278 1004
rect 316 976 344 1004
rect 382 976 410 1004
rect 448 976 476 1004
rect 514 976 542 1004
rect 580 976 608 1004
rect 646 976 674 1004
rect 712 976 740 1004
rect -740 910 -712 938
rect -674 910 -646 938
rect -608 910 -580 938
rect -542 910 -514 938
rect -476 910 -448 938
rect -410 910 -382 938
rect -344 910 -316 938
rect -278 910 -250 938
rect -212 910 -184 938
rect -146 910 -118 938
rect -80 910 -52 938
rect -14 910 14 938
rect 52 910 80 938
rect 118 910 146 938
rect 184 910 212 938
rect 250 910 278 938
rect 316 910 344 938
rect 382 910 410 938
rect 448 910 476 938
rect 514 910 542 938
rect 580 910 608 938
rect 646 910 674 938
rect 712 910 740 938
rect -740 844 -712 872
rect -674 844 -646 872
rect -608 844 -580 872
rect -542 844 -514 872
rect -476 844 -448 872
rect -410 844 -382 872
rect -344 844 -316 872
rect -278 844 -250 872
rect -212 844 -184 872
rect -146 844 -118 872
rect -80 844 -52 872
rect -14 844 14 872
rect 52 844 80 872
rect 118 844 146 872
rect 184 844 212 872
rect 250 844 278 872
rect 316 844 344 872
rect 382 844 410 872
rect 448 844 476 872
rect 514 844 542 872
rect 580 844 608 872
rect 646 844 674 872
rect 712 844 740 872
rect -740 778 -712 806
rect -674 778 -646 806
rect -608 778 -580 806
rect -542 778 -514 806
rect -476 778 -448 806
rect -410 778 -382 806
rect -344 778 -316 806
rect -278 778 -250 806
rect -212 778 -184 806
rect -146 778 -118 806
rect -80 778 -52 806
rect -14 778 14 806
rect 52 778 80 806
rect 118 778 146 806
rect 184 778 212 806
rect 250 778 278 806
rect 316 778 344 806
rect 382 778 410 806
rect 448 778 476 806
rect 514 778 542 806
rect 580 778 608 806
rect 646 778 674 806
rect 712 778 740 806
rect -740 712 -712 740
rect -674 712 -646 740
rect -608 712 -580 740
rect -542 712 -514 740
rect -476 712 -448 740
rect -410 712 -382 740
rect -344 712 -316 740
rect -278 712 -250 740
rect -212 712 -184 740
rect -146 712 -118 740
rect -80 712 -52 740
rect -14 712 14 740
rect 52 712 80 740
rect 118 712 146 740
rect 184 712 212 740
rect 250 712 278 740
rect 316 712 344 740
rect 382 712 410 740
rect 448 712 476 740
rect 514 712 542 740
rect 580 712 608 740
rect 646 712 674 740
rect 712 712 740 740
rect -740 646 -712 674
rect -674 646 -646 674
rect -608 646 -580 674
rect -542 646 -514 674
rect -476 646 -448 674
rect -410 646 -382 674
rect -344 646 -316 674
rect -278 646 -250 674
rect -212 646 -184 674
rect -146 646 -118 674
rect -80 646 -52 674
rect -14 646 14 674
rect 52 646 80 674
rect 118 646 146 674
rect 184 646 212 674
rect 250 646 278 674
rect 316 646 344 674
rect 382 646 410 674
rect 448 646 476 674
rect 514 646 542 674
rect 580 646 608 674
rect 646 646 674 674
rect 712 646 740 674
rect -740 580 -712 608
rect -674 580 -646 608
rect -608 580 -580 608
rect -542 580 -514 608
rect -476 580 -448 608
rect -410 580 -382 608
rect -344 580 -316 608
rect -278 580 -250 608
rect -212 580 -184 608
rect -146 580 -118 608
rect -80 580 -52 608
rect -14 580 14 608
rect 52 580 80 608
rect 118 580 146 608
rect 184 580 212 608
rect 250 580 278 608
rect 316 580 344 608
rect 382 580 410 608
rect 448 580 476 608
rect 514 580 542 608
rect 580 580 608 608
rect 646 580 674 608
rect 712 580 740 608
rect -740 514 -712 542
rect -674 514 -646 542
rect -608 514 -580 542
rect -542 514 -514 542
rect -476 514 -448 542
rect -410 514 -382 542
rect -344 514 -316 542
rect -278 514 -250 542
rect -212 514 -184 542
rect -146 514 -118 542
rect -80 514 -52 542
rect -14 514 14 542
rect 52 514 80 542
rect 118 514 146 542
rect 184 514 212 542
rect 250 514 278 542
rect 316 514 344 542
rect 382 514 410 542
rect 448 514 476 542
rect 514 514 542 542
rect 580 514 608 542
rect 646 514 674 542
rect 712 514 740 542
rect -740 448 -712 476
rect -674 448 -646 476
rect -608 448 -580 476
rect -542 448 -514 476
rect -476 448 -448 476
rect -410 448 -382 476
rect -344 448 -316 476
rect -278 448 -250 476
rect -212 448 -184 476
rect -146 448 -118 476
rect -80 448 -52 476
rect -14 448 14 476
rect 52 448 80 476
rect 118 448 146 476
rect 184 448 212 476
rect 250 448 278 476
rect 316 448 344 476
rect 382 448 410 476
rect 448 448 476 476
rect 514 448 542 476
rect 580 448 608 476
rect 646 448 674 476
rect 712 448 740 476
rect -740 382 -712 410
rect -674 382 -646 410
rect -608 382 -580 410
rect -542 382 -514 410
rect -476 382 -448 410
rect -410 382 -382 410
rect -344 382 -316 410
rect -278 382 -250 410
rect -212 382 -184 410
rect -146 382 -118 410
rect -80 382 -52 410
rect -14 382 14 410
rect 52 382 80 410
rect 118 382 146 410
rect 184 382 212 410
rect 250 382 278 410
rect 316 382 344 410
rect 382 382 410 410
rect 448 382 476 410
rect 514 382 542 410
rect 580 382 608 410
rect 646 382 674 410
rect 712 382 740 410
rect -740 316 -712 344
rect -674 316 -646 344
rect -608 316 -580 344
rect -542 316 -514 344
rect -476 316 -448 344
rect -410 316 -382 344
rect -344 316 -316 344
rect -278 316 -250 344
rect -212 316 -184 344
rect -146 316 -118 344
rect -80 316 -52 344
rect -14 316 14 344
rect 52 316 80 344
rect 118 316 146 344
rect 184 316 212 344
rect 250 316 278 344
rect 316 316 344 344
rect 382 316 410 344
rect 448 316 476 344
rect 514 316 542 344
rect 580 316 608 344
rect 646 316 674 344
rect 712 316 740 344
rect -740 250 -712 278
rect -674 250 -646 278
rect -608 250 -580 278
rect -542 250 -514 278
rect -476 250 -448 278
rect -410 250 -382 278
rect -344 250 -316 278
rect -278 250 -250 278
rect -212 250 -184 278
rect -146 250 -118 278
rect -80 250 -52 278
rect -14 250 14 278
rect 52 250 80 278
rect 118 250 146 278
rect 184 250 212 278
rect 250 250 278 278
rect 316 250 344 278
rect 382 250 410 278
rect 448 250 476 278
rect 514 250 542 278
rect 580 250 608 278
rect 646 250 674 278
rect 712 250 740 278
rect -740 184 -712 212
rect -674 184 -646 212
rect -608 184 -580 212
rect -542 184 -514 212
rect -476 184 -448 212
rect -410 184 -382 212
rect -344 184 -316 212
rect -278 184 -250 212
rect -212 184 -184 212
rect -146 184 -118 212
rect -80 184 -52 212
rect -14 184 14 212
rect 52 184 80 212
rect 118 184 146 212
rect 184 184 212 212
rect 250 184 278 212
rect 316 184 344 212
rect 382 184 410 212
rect 448 184 476 212
rect 514 184 542 212
rect 580 184 608 212
rect 646 184 674 212
rect 712 184 740 212
rect -740 118 -712 146
rect -674 118 -646 146
rect -608 118 -580 146
rect -542 118 -514 146
rect -476 118 -448 146
rect -410 118 -382 146
rect -344 118 -316 146
rect -278 118 -250 146
rect -212 118 -184 146
rect -146 118 -118 146
rect -80 118 -52 146
rect -14 118 14 146
rect 52 118 80 146
rect 118 118 146 146
rect 184 118 212 146
rect 250 118 278 146
rect 316 118 344 146
rect 382 118 410 146
rect 448 118 476 146
rect 514 118 542 146
rect 580 118 608 146
rect 646 118 674 146
rect 712 118 740 146
rect -740 52 -712 80
rect -674 52 -646 80
rect -608 52 -580 80
rect -542 52 -514 80
rect -476 52 -448 80
rect -410 52 -382 80
rect -344 52 -316 80
rect -278 52 -250 80
rect -212 52 -184 80
rect -146 52 -118 80
rect -80 52 -52 80
rect -14 52 14 80
rect 52 52 80 80
rect 118 52 146 80
rect 184 52 212 80
rect 250 52 278 80
rect 316 52 344 80
rect 382 52 410 80
rect 448 52 476 80
rect 514 52 542 80
rect 580 52 608 80
rect 646 52 674 80
rect 712 52 740 80
rect -740 -14 -712 14
rect -674 -14 -646 14
rect -608 -14 -580 14
rect -542 -14 -514 14
rect -476 -14 -448 14
rect -410 -14 -382 14
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
rect 52 -14 80 14
rect 118 -14 146 14
rect 184 -14 212 14
rect 250 -14 278 14
rect 316 -14 344 14
rect 382 -14 410 14
rect 448 -14 476 14
rect 514 -14 542 14
rect 580 -14 608 14
rect 646 -14 674 14
rect 712 -14 740 14
rect -740 -80 -712 -52
rect -674 -80 -646 -52
rect -608 -80 -580 -52
rect -542 -80 -514 -52
rect -476 -80 -448 -52
rect -410 -80 -382 -52
rect -344 -80 -316 -52
rect -278 -80 -250 -52
rect -212 -80 -184 -52
rect -146 -80 -118 -52
rect -80 -80 -52 -52
rect -14 -80 14 -52
rect 52 -80 80 -52
rect 118 -80 146 -52
rect 184 -80 212 -52
rect 250 -80 278 -52
rect 316 -80 344 -52
rect 382 -80 410 -52
rect 448 -80 476 -52
rect 514 -80 542 -52
rect 580 -80 608 -52
rect 646 -80 674 -52
rect 712 -80 740 -52
rect -740 -146 -712 -118
rect -674 -146 -646 -118
rect -608 -146 -580 -118
rect -542 -146 -514 -118
rect -476 -146 -448 -118
rect -410 -146 -382 -118
rect -344 -146 -316 -118
rect -278 -146 -250 -118
rect -212 -146 -184 -118
rect -146 -146 -118 -118
rect -80 -146 -52 -118
rect -14 -146 14 -118
rect 52 -146 80 -118
rect 118 -146 146 -118
rect 184 -146 212 -118
rect 250 -146 278 -118
rect 316 -146 344 -118
rect 382 -146 410 -118
rect 448 -146 476 -118
rect 514 -146 542 -118
rect 580 -146 608 -118
rect 646 -146 674 -118
rect 712 -146 740 -118
rect -740 -212 -712 -184
rect -674 -212 -646 -184
rect -608 -212 -580 -184
rect -542 -212 -514 -184
rect -476 -212 -448 -184
rect -410 -212 -382 -184
rect -344 -212 -316 -184
rect -278 -212 -250 -184
rect -212 -212 -184 -184
rect -146 -212 -118 -184
rect -80 -212 -52 -184
rect -14 -212 14 -184
rect 52 -212 80 -184
rect 118 -212 146 -184
rect 184 -212 212 -184
rect 250 -212 278 -184
rect 316 -212 344 -184
rect 382 -212 410 -184
rect 448 -212 476 -184
rect 514 -212 542 -184
rect 580 -212 608 -184
rect 646 -212 674 -184
rect 712 -212 740 -184
rect -740 -278 -712 -250
rect -674 -278 -646 -250
rect -608 -278 -580 -250
rect -542 -278 -514 -250
rect -476 -278 -448 -250
rect -410 -278 -382 -250
rect -344 -278 -316 -250
rect -278 -278 -250 -250
rect -212 -278 -184 -250
rect -146 -278 -118 -250
rect -80 -278 -52 -250
rect -14 -278 14 -250
rect 52 -278 80 -250
rect 118 -278 146 -250
rect 184 -278 212 -250
rect 250 -278 278 -250
rect 316 -278 344 -250
rect 382 -278 410 -250
rect 448 -278 476 -250
rect 514 -278 542 -250
rect 580 -278 608 -250
rect 646 -278 674 -250
rect 712 -278 740 -250
rect -740 -344 -712 -316
rect -674 -344 -646 -316
rect -608 -344 -580 -316
rect -542 -344 -514 -316
rect -476 -344 -448 -316
rect -410 -344 -382 -316
rect -344 -344 -316 -316
rect -278 -344 -250 -316
rect -212 -344 -184 -316
rect -146 -344 -118 -316
rect -80 -344 -52 -316
rect -14 -344 14 -316
rect 52 -344 80 -316
rect 118 -344 146 -316
rect 184 -344 212 -316
rect 250 -344 278 -316
rect 316 -344 344 -316
rect 382 -344 410 -316
rect 448 -344 476 -316
rect 514 -344 542 -316
rect 580 -344 608 -316
rect 646 -344 674 -316
rect 712 -344 740 -316
rect -740 -410 -712 -382
rect -674 -410 -646 -382
rect -608 -410 -580 -382
rect -542 -410 -514 -382
rect -476 -410 -448 -382
rect -410 -410 -382 -382
rect -344 -410 -316 -382
rect -278 -410 -250 -382
rect -212 -410 -184 -382
rect -146 -410 -118 -382
rect -80 -410 -52 -382
rect -14 -410 14 -382
rect 52 -410 80 -382
rect 118 -410 146 -382
rect 184 -410 212 -382
rect 250 -410 278 -382
rect 316 -410 344 -382
rect 382 -410 410 -382
rect 448 -410 476 -382
rect 514 -410 542 -382
rect 580 -410 608 -382
rect 646 -410 674 -382
rect 712 -410 740 -382
rect -740 -476 -712 -448
rect -674 -476 -646 -448
rect -608 -476 -580 -448
rect -542 -476 -514 -448
rect -476 -476 -448 -448
rect -410 -476 -382 -448
rect -344 -476 -316 -448
rect -278 -476 -250 -448
rect -212 -476 -184 -448
rect -146 -476 -118 -448
rect -80 -476 -52 -448
rect -14 -476 14 -448
rect 52 -476 80 -448
rect 118 -476 146 -448
rect 184 -476 212 -448
rect 250 -476 278 -448
rect 316 -476 344 -448
rect 382 -476 410 -448
rect 448 -476 476 -448
rect 514 -476 542 -448
rect 580 -476 608 -448
rect 646 -476 674 -448
rect 712 -476 740 -448
rect -740 -542 -712 -514
rect -674 -542 -646 -514
rect -608 -542 -580 -514
rect -542 -542 -514 -514
rect -476 -542 -448 -514
rect -410 -542 -382 -514
rect -344 -542 -316 -514
rect -278 -542 -250 -514
rect -212 -542 -184 -514
rect -146 -542 -118 -514
rect -80 -542 -52 -514
rect -14 -542 14 -514
rect 52 -542 80 -514
rect 118 -542 146 -514
rect 184 -542 212 -514
rect 250 -542 278 -514
rect 316 -542 344 -514
rect 382 -542 410 -514
rect 448 -542 476 -514
rect 514 -542 542 -514
rect 580 -542 608 -514
rect 646 -542 674 -514
rect 712 -542 740 -514
rect -740 -608 -712 -580
rect -674 -608 -646 -580
rect -608 -608 -580 -580
rect -542 -608 -514 -580
rect -476 -608 -448 -580
rect -410 -608 -382 -580
rect -344 -608 -316 -580
rect -278 -608 -250 -580
rect -212 -608 -184 -580
rect -146 -608 -118 -580
rect -80 -608 -52 -580
rect -14 -608 14 -580
rect 52 -608 80 -580
rect 118 -608 146 -580
rect 184 -608 212 -580
rect 250 -608 278 -580
rect 316 -608 344 -580
rect 382 -608 410 -580
rect 448 -608 476 -580
rect 514 -608 542 -580
rect 580 -608 608 -580
rect 646 -608 674 -580
rect 712 -608 740 -580
rect -740 -674 -712 -646
rect -674 -674 -646 -646
rect -608 -674 -580 -646
rect -542 -674 -514 -646
rect -476 -674 -448 -646
rect -410 -674 -382 -646
rect -344 -674 -316 -646
rect -278 -674 -250 -646
rect -212 -674 -184 -646
rect -146 -674 -118 -646
rect -80 -674 -52 -646
rect -14 -674 14 -646
rect 52 -674 80 -646
rect 118 -674 146 -646
rect 184 -674 212 -646
rect 250 -674 278 -646
rect 316 -674 344 -646
rect 382 -674 410 -646
rect 448 -674 476 -646
rect 514 -674 542 -646
rect 580 -674 608 -646
rect 646 -674 674 -646
rect 712 -674 740 -646
rect -740 -740 -712 -712
rect -674 -740 -646 -712
rect -608 -740 -580 -712
rect -542 -740 -514 -712
rect -476 -740 -448 -712
rect -410 -740 -382 -712
rect -344 -740 -316 -712
rect -278 -740 -250 -712
rect -212 -740 -184 -712
rect -146 -740 -118 -712
rect -80 -740 -52 -712
rect -14 -740 14 -712
rect 52 -740 80 -712
rect 118 -740 146 -712
rect 184 -740 212 -712
rect 250 -740 278 -712
rect 316 -740 344 -712
rect 382 -740 410 -712
rect 448 -740 476 -712
rect 514 -740 542 -712
rect 580 -740 608 -712
rect 646 -740 674 -712
rect 712 -740 740 -712
rect -740 -806 -712 -778
rect -674 -806 -646 -778
rect -608 -806 -580 -778
rect -542 -806 -514 -778
rect -476 -806 -448 -778
rect -410 -806 -382 -778
rect -344 -806 -316 -778
rect -278 -806 -250 -778
rect -212 -806 -184 -778
rect -146 -806 -118 -778
rect -80 -806 -52 -778
rect -14 -806 14 -778
rect 52 -806 80 -778
rect 118 -806 146 -778
rect 184 -806 212 -778
rect 250 -806 278 -778
rect 316 -806 344 -778
rect 382 -806 410 -778
rect 448 -806 476 -778
rect 514 -806 542 -778
rect 580 -806 608 -778
rect 646 -806 674 -778
rect 712 -806 740 -778
rect -740 -872 -712 -844
rect -674 -872 -646 -844
rect -608 -872 -580 -844
rect -542 -872 -514 -844
rect -476 -872 -448 -844
rect -410 -872 -382 -844
rect -344 -872 -316 -844
rect -278 -872 -250 -844
rect -212 -872 -184 -844
rect -146 -872 -118 -844
rect -80 -872 -52 -844
rect -14 -872 14 -844
rect 52 -872 80 -844
rect 118 -872 146 -844
rect 184 -872 212 -844
rect 250 -872 278 -844
rect 316 -872 344 -844
rect 382 -872 410 -844
rect 448 -872 476 -844
rect 514 -872 542 -844
rect 580 -872 608 -844
rect 646 -872 674 -844
rect 712 -872 740 -844
rect -740 -938 -712 -910
rect -674 -938 -646 -910
rect -608 -938 -580 -910
rect -542 -938 -514 -910
rect -476 -938 -448 -910
rect -410 -938 -382 -910
rect -344 -938 -316 -910
rect -278 -938 -250 -910
rect -212 -938 -184 -910
rect -146 -938 -118 -910
rect -80 -938 -52 -910
rect -14 -938 14 -910
rect 52 -938 80 -910
rect 118 -938 146 -910
rect 184 -938 212 -910
rect 250 -938 278 -910
rect 316 -938 344 -910
rect 382 -938 410 -910
rect 448 -938 476 -910
rect 514 -938 542 -910
rect 580 -938 608 -910
rect 646 -938 674 -910
rect 712 -938 740 -910
rect -740 -1004 -712 -976
rect -674 -1004 -646 -976
rect -608 -1004 -580 -976
rect -542 -1004 -514 -976
rect -476 -1004 -448 -976
rect -410 -1004 -382 -976
rect -344 -1004 -316 -976
rect -278 -1004 -250 -976
rect -212 -1004 -184 -976
rect -146 -1004 -118 -976
rect -80 -1004 -52 -976
rect -14 -1004 14 -976
rect 52 -1004 80 -976
rect 118 -1004 146 -976
rect 184 -1004 212 -976
rect 250 -1004 278 -976
rect 316 -1004 344 -976
rect 382 -1004 410 -976
rect 448 -1004 476 -976
rect 514 -1004 542 -976
rect 580 -1004 608 -976
rect 646 -1004 674 -976
rect 712 -1004 740 -976
rect -740 -1070 -712 -1042
rect -674 -1070 -646 -1042
rect -608 -1070 -580 -1042
rect -542 -1070 -514 -1042
rect -476 -1070 -448 -1042
rect -410 -1070 -382 -1042
rect -344 -1070 -316 -1042
rect -278 -1070 -250 -1042
rect -212 -1070 -184 -1042
rect -146 -1070 -118 -1042
rect -80 -1070 -52 -1042
rect -14 -1070 14 -1042
rect 52 -1070 80 -1042
rect 118 -1070 146 -1042
rect 184 -1070 212 -1042
rect 250 -1070 278 -1042
rect 316 -1070 344 -1042
rect 382 -1070 410 -1042
rect 448 -1070 476 -1042
rect 514 -1070 542 -1042
rect 580 -1070 608 -1042
rect 646 -1070 674 -1042
rect 712 -1070 740 -1042
rect -740 -1136 -712 -1108
rect -674 -1136 -646 -1108
rect -608 -1136 -580 -1108
rect -542 -1136 -514 -1108
rect -476 -1136 -448 -1108
rect -410 -1136 -382 -1108
rect -344 -1136 -316 -1108
rect -278 -1136 -250 -1108
rect -212 -1136 -184 -1108
rect -146 -1136 -118 -1108
rect -80 -1136 -52 -1108
rect -14 -1136 14 -1108
rect 52 -1136 80 -1108
rect 118 -1136 146 -1108
rect 184 -1136 212 -1108
rect 250 -1136 278 -1108
rect 316 -1136 344 -1108
rect 382 -1136 410 -1108
rect 448 -1136 476 -1108
rect 514 -1136 542 -1108
rect 580 -1136 608 -1108
rect 646 -1136 674 -1108
rect 712 -1136 740 -1108
rect -740 -1202 -712 -1174
rect -674 -1202 -646 -1174
rect -608 -1202 -580 -1174
rect -542 -1202 -514 -1174
rect -476 -1202 -448 -1174
rect -410 -1202 -382 -1174
rect -344 -1202 -316 -1174
rect -278 -1202 -250 -1174
rect -212 -1202 -184 -1174
rect -146 -1202 -118 -1174
rect -80 -1202 -52 -1174
rect -14 -1202 14 -1174
rect 52 -1202 80 -1174
rect 118 -1202 146 -1174
rect 184 -1202 212 -1174
rect 250 -1202 278 -1174
rect 316 -1202 344 -1174
rect 382 -1202 410 -1174
rect 448 -1202 476 -1174
rect 514 -1202 542 -1174
rect 580 -1202 608 -1174
rect 646 -1202 674 -1174
rect 712 -1202 740 -1174
rect -740 -1268 -712 -1240
rect -674 -1268 -646 -1240
rect -608 -1268 -580 -1240
rect -542 -1268 -514 -1240
rect -476 -1268 -448 -1240
rect -410 -1268 -382 -1240
rect -344 -1268 -316 -1240
rect -278 -1268 -250 -1240
rect -212 -1268 -184 -1240
rect -146 -1268 -118 -1240
rect -80 -1268 -52 -1240
rect -14 -1268 14 -1240
rect 52 -1268 80 -1240
rect 118 -1268 146 -1240
rect 184 -1268 212 -1240
rect 250 -1268 278 -1240
rect 316 -1268 344 -1240
rect 382 -1268 410 -1240
rect 448 -1268 476 -1240
rect 514 -1268 542 -1240
rect 580 -1268 608 -1240
rect 646 -1268 674 -1240
rect 712 -1268 740 -1240
rect -740 -1334 -712 -1306
rect -674 -1334 -646 -1306
rect -608 -1334 -580 -1306
rect -542 -1334 -514 -1306
rect -476 -1334 -448 -1306
rect -410 -1334 -382 -1306
rect -344 -1334 -316 -1306
rect -278 -1334 -250 -1306
rect -212 -1334 -184 -1306
rect -146 -1334 -118 -1306
rect -80 -1334 -52 -1306
rect -14 -1334 14 -1306
rect 52 -1334 80 -1306
rect 118 -1334 146 -1306
rect 184 -1334 212 -1306
rect 250 -1334 278 -1306
rect 316 -1334 344 -1306
rect 382 -1334 410 -1306
rect 448 -1334 476 -1306
rect 514 -1334 542 -1306
rect 580 -1334 608 -1306
rect 646 -1334 674 -1306
rect 712 -1334 740 -1306
rect -740 -1400 -712 -1372
rect -674 -1400 -646 -1372
rect -608 -1400 -580 -1372
rect -542 -1400 -514 -1372
rect -476 -1400 -448 -1372
rect -410 -1400 -382 -1372
rect -344 -1400 -316 -1372
rect -278 -1400 -250 -1372
rect -212 -1400 -184 -1372
rect -146 -1400 -118 -1372
rect -80 -1400 -52 -1372
rect -14 -1400 14 -1372
rect 52 -1400 80 -1372
rect 118 -1400 146 -1372
rect 184 -1400 212 -1372
rect 250 -1400 278 -1372
rect 316 -1400 344 -1372
rect 382 -1400 410 -1372
rect 448 -1400 476 -1372
rect 514 -1400 542 -1372
rect 580 -1400 608 -1372
rect 646 -1400 674 -1372
rect 712 -1400 740 -1372
rect -740 -1466 -712 -1438
rect -674 -1466 -646 -1438
rect -608 -1466 -580 -1438
rect -542 -1466 -514 -1438
rect -476 -1466 -448 -1438
rect -410 -1466 -382 -1438
rect -344 -1466 -316 -1438
rect -278 -1466 -250 -1438
rect -212 -1466 -184 -1438
rect -146 -1466 -118 -1438
rect -80 -1466 -52 -1438
rect -14 -1466 14 -1438
rect 52 -1466 80 -1438
rect 118 -1466 146 -1438
rect 184 -1466 212 -1438
rect 250 -1466 278 -1438
rect 316 -1466 344 -1438
rect 382 -1466 410 -1438
rect 448 -1466 476 -1438
rect 514 -1466 542 -1438
rect 580 -1466 608 -1438
rect 646 -1466 674 -1438
rect 712 -1466 740 -1438
rect -740 -1532 -712 -1504
rect -674 -1532 -646 -1504
rect -608 -1532 -580 -1504
rect -542 -1532 -514 -1504
rect -476 -1532 -448 -1504
rect -410 -1532 -382 -1504
rect -344 -1532 -316 -1504
rect -278 -1532 -250 -1504
rect -212 -1532 -184 -1504
rect -146 -1532 -118 -1504
rect -80 -1532 -52 -1504
rect -14 -1532 14 -1504
rect 52 -1532 80 -1504
rect 118 -1532 146 -1504
rect 184 -1532 212 -1504
rect 250 -1532 278 -1504
rect 316 -1532 344 -1504
rect 382 -1532 410 -1504
rect 448 -1532 476 -1504
rect 514 -1532 542 -1504
rect 580 -1532 608 -1504
rect 646 -1532 674 -1504
rect 712 -1532 740 -1504
rect -740 -1598 -712 -1570
rect -674 -1598 -646 -1570
rect -608 -1598 -580 -1570
rect -542 -1598 -514 -1570
rect -476 -1598 -448 -1570
rect -410 -1598 -382 -1570
rect -344 -1598 -316 -1570
rect -278 -1598 -250 -1570
rect -212 -1598 -184 -1570
rect -146 -1598 -118 -1570
rect -80 -1598 -52 -1570
rect -14 -1598 14 -1570
rect 52 -1598 80 -1570
rect 118 -1598 146 -1570
rect 184 -1598 212 -1570
rect 250 -1598 278 -1570
rect 316 -1598 344 -1570
rect 382 -1598 410 -1570
rect 448 -1598 476 -1570
rect 514 -1598 542 -1570
rect 580 -1598 608 -1570
rect 646 -1598 674 -1570
rect 712 -1598 740 -1570
rect -740 -1664 -712 -1636
rect -674 -1664 -646 -1636
rect -608 -1664 -580 -1636
rect -542 -1664 -514 -1636
rect -476 -1664 -448 -1636
rect -410 -1664 -382 -1636
rect -344 -1664 -316 -1636
rect -278 -1664 -250 -1636
rect -212 -1664 -184 -1636
rect -146 -1664 -118 -1636
rect -80 -1664 -52 -1636
rect -14 -1664 14 -1636
rect 52 -1664 80 -1636
rect 118 -1664 146 -1636
rect 184 -1664 212 -1636
rect 250 -1664 278 -1636
rect 316 -1664 344 -1636
rect 382 -1664 410 -1636
rect 448 -1664 476 -1636
rect 514 -1664 542 -1636
rect 580 -1664 608 -1636
rect 646 -1664 674 -1636
rect 712 -1664 740 -1636
rect -740 -1730 -712 -1702
rect -674 -1730 -646 -1702
rect -608 -1730 -580 -1702
rect -542 -1730 -514 -1702
rect -476 -1730 -448 -1702
rect -410 -1730 -382 -1702
rect -344 -1730 -316 -1702
rect -278 -1730 -250 -1702
rect -212 -1730 -184 -1702
rect -146 -1730 -118 -1702
rect -80 -1730 -52 -1702
rect -14 -1730 14 -1702
rect 52 -1730 80 -1702
rect 118 -1730 146 -1702
rect 184 -1730 212 -1702
rect 250 -1730 278 -1702
rect 316 -1730 344 -1702
rect 382 -1730 410 -1702
rect 448 -1730 476 -1702
rect 514 -1730 542 -1702
rect 580 -1730 608 -1702
rect 646 -1730 674 -1702
rect 712 -1730 740 -1702
rect -740 -1796 -712 -1768
rect -674 -1796 -646 -1768
rect -608 -1796 -580 -1768
rect -542 -1796 -514 -1768
rect -476 -1796 -448 -1768
rect -410 -1796 -382 -1768
rect -344 -1796 -316 -1768
rect -278 -1796 -250 -1768
rect -212 -1796 -184 -1768
rect -146 -1796 -118 -1768
rect -80 -1796 -52 -1768
rect -14 -1796 14 -1768
rect 52 -1796 80 -1768
rect 118 -1796 146 -1768
rect 184 -1796 212 -1768
rect 250 -1796 278 -1768
rect 316 -1796 344 -1768
rect 382 -1796 410 -1768
rect 448 -1796 476 -1768
rect 514 -1796 542 -1768
rect 580 -1796 608 -1768
rect 646 -1796 674 -1768
rect 712 -1796 740 -1768
rect -740 -1862 -712 -1834
rect -674 -1862 -646 -1834
rect -608 -1862 -580 -1834
rect -542 -1862 -514 -1834
rect -476 -1862 -448 -1834
rect -410 -1862 -382 -1834
rect -344 -1862 -316 -1834
rect -278 -1862 -250 -1834
rect -212 -1862 -184 -1834
rect -146 -1862 -118 -1834
rect -80 -1862 -52 -1834
rect -14 -1862 14 -1834
rect 52 -1862 80 -1834
rect 118 -1862 146 -1834
rect 184 -1862 212 -1834
rect 250 -1862 278 -1834
rect 316 -1862 344 -1834
rect 382 -1862 410 -1834
rect 448 -1862 476 -1834
rect 514 -1862 542 -1834
rect 580 -1862 608 -1834
rect 646 -1862 674 -1834
rect 712 -1862 740 -1834
rect -740 -1928 -712 -1900
rect -674 -1928 -646 -1900
rect -608 -1928 -580 -1900
rect -542 -1928 -514 -1900
rect -476 -1928 -448 -1900
rect -410 -1928 -382 -1900
rect -344 -1928 -316 -1900
rect -278 -1928 -250 -1900
rect -212 -1928 -184 -1900
rect -146 -1928 -118 -1900
rect -80 -1928 -52 -1900
rect -14 -1928 14 -1900
rect 52 -1928 80 -1900
rect 118 -1928 146 -1900
rect 184 -1928 212 -1900
rect 250 -1928 278 -1900
rect 316 -1928 344 -1900
rect 382 -1928 410 -1900
rect 448 -1928 476 -1900
rect 514 -1928 542 -1900
rect 580 -1928 608 -1900
rect 646 -1928 674 -1900
rect 712 -1928 740 -1900
rect -740 -1994 -712 -1966
rect -674 -1994 -646 -1966
rect -608 -1994 -580 -1966
rect -542 -1994 -514 -1966
rect -476 -1994 -448 -1966
rect -410 -1994 -382 -1966
rect -344 -1994 -316 -1966
rect -278 -1994 -250 -1966
rect -212 -1994 -184 -1966
rect -146 -1994 -118 -1966
rect -80 -1994 -52 -1966
rect -14 -1994 14 -1966
rect 52 -1994 80 -1966
rect 118 -1994 146 -1966
rect 184 -1994 212 -1966
rect 250 -1994 278 -1966
rect 316 -1994 344 -1966
rect 382 -1994 410 -1966
rect 448 -1994 476 -1966
rect 514 -1994 542 -1966
rect 580 -1994 608 -1966
rect 646 -1994 674 -1966
rect 712 -1994 740 -1966
rect -740 -2060 -712 -2032
rect -674 -2060 -646 -2032
rect -608 -2060 -580 -2032
rect -542 -2060 -514 -2032
rect -476 -2060 -448 -2032
rect -410 -2060 -382 -2032
rect -344 -2060 -316 -2032
rect -278 -2060 -250 -2032
rect -212 -2060 -184 -2032
rect -146 -2060 -118 -2032
rect -80 -2060 -52 -2032
rect -14 -2060 14 -2032
rect 52 -2060 80 -2032
rect 118 -2060 146 -2032
rect 184 -2060 212 -2032
rect 250 -2060 278 -2032
rect 316 -2060 344 -2032
rect 382 -2060 410 -2032
rect 448 -2060 476 -2032
rect 514 -2060 542 -2032
rect 580 -2060 608 -2032
rect 646 -2060 674 -2032
rect 712 -2060 740 -2032
rect -740 -2126 -712 -2098
rect -674 -2126 -646 -2098
rect -608 -2126 -580 -2098
rect -542 -2126 -514 -2098
rect -476 -2126 -448 -2098
rect -410 -2126 -382 -2098
rect -344 -2126 -316 -2098
rect -278 -2126 -250 -2098
rect -212 -2126 -184 -2098
rect -146 -2126 -118 -2098
rect -80 -2126 -52 -2098
rect -14 -2126 14 -2098
rect 52 -2126 80 -2098
rect 118 -2126 146 -2098
rect 184 -2126 212 -2098
rect 250 -2126 278 -2098
rect 316 -2126 344 -2098
rect 382 -2126 410 -2098
rect 448 -2126 476 -2098
rect 514 -2126 542 -2098
rect 580 -2126 608 -2098
rect 646 -2126 674 -2098
rect 712 -2126 740 -2098
rect -740 -2192 -712 -2164
rect -674 -2192 -646 -2164
rect -608 -2192 -580 -2164
rect -542 -2192 -514 -2164
rect -476 -2192 -448 -2164
rect -410 -2192 -382 -2164
rect -344 -2192 -316 -2164
rect -278 -2192 -250 -2164
rect -212 -2192 -184 -2164
rect -146 -2192 -118 -2164
rect -80 -2192 -52 -2164
rect -14 -2192 14 -2164
rect 52 -2192 80 -2164
rect 118 -2192 146 -2164
rect 184 -2192 212 -2164
rect 250 -2192 278 -2164
rect 316 -2192 344 -2164
rect 382 -2192 410 -2164
rect 448 -2192 476 -2164
rect 514 -2192 542 -2164
rect 580 -2192 608 -2164
rect 646 -2192 674 -2164
rect 712 -2192 740 -2164
rect -740 -2258 -712 -2230
rect -674 -2258 -646 -2230
rect -608 -2258 -580 -2230
rect -542 -2258 -514 -2230
rect -476 -2258 -448 -2230
rect -410 -2258 -382 -2230
rect -344 -2258 -316 -2230
rect -278 -2258 -250 -2230
rect -212 -2258 -184 -2230
rect -146 -2258 -118 -2230
rect -80 -2258 -52 -2230
rect -14 -2258 14 -2230
rect 52 -2258 80 -2230
rect 118 -2258 146 -2230
rect 184 -2258 212 -2230
rect 250 -2258 278 -2230
rect 316 -2258 344 -2230
rect 382 -2258 410 -2230
rect 448 -2258 476 -2230
rect 514 -2258 542 -2230
rect 580 -2258 608 -2230
rect 646 -2258 674 -2230
rect 712 -2258 740 -2230
rect -740 -2324 -712 -2296
rect -674 -2324 -646 -2296
rect -608 -2324 -580 -2296
rect -542 -2324 -514 -2296
rect -476 -2324 -448 -2296
rect -410 -2324 -382 -2296
rect -344 -2324 -316 -2296
rect -278 -2324 -250 -2296
rect -212 -2324 -184 -2296
rect -146 -2324 -118 -2296
rect -80 -2324 -52 -2296
rect -14 -2324 14 -2296
rect 52 -2324 80 -2296
rect 118 -2324 146 -2296
rect 184 -2324 212 -2296
rect 250 -2324 278 -2296
rect 316 -2324 344 -2296
rect 382 -2324 410 -2296
rect 448 -2324 476 -2296
rect 514 -2324 542 -2296
rect 580 -2324 608 -2296
rect 646 -2324 674 -2296
rect 712 -2324 740 -2296
rect -740 -2390 -712 -2362
rect -674 -2390 -646 -2362
rect -608 -2390 -580 -2362
rect -542 -2390 -514 -2362
rect -476 -2390 -448 -2362
rect -410 -2390 -382 -2362
rect -344 -2390 -316 -2362
rect -278 -2390 -250 -2362
rect -212 -2390 -184 -2362
rect -146 -2390 -118 -2362
rect -80 -2390 -52 -2362
rect -14 -2390 14 -2362
rect 52 -2390 80 -2362
rect 118 -2390 146 -2362
rect 184 -2390 212 -2362
rect 250 -2390 278 -2362
rect 316 -2390 344 -2362
rect 382 -2390 410 -2362
rect 448 -2390 476 -2362
rect 514 -2390 542 -2362
rect 580 -2390 608 -2362
rect 646 -2390 674 -2362
rect 712 -2390 740 -2362
rect -740 -2456 -712 -2428
rect -674 -2456 -646 -2428
rect -608 -2456 -580 -2428
rect -542 -2456 -514 -2428
rect -476 -2456 -448 -2428
rect -410 -2456 -382 -2428
rect -344 -2456 -316 -2428
rect -278 -2456 -250 -2428
rect -212 -2456 -184 -2428
rect -146 -2456 -118 -2428
rect -80 -2456 -52 -2428
rect -14 -2456 14 -2428
rect 52 -2456 80 -2428
rect 118 -2456 146 -2428
rect 184 -2456 212 -2428
rect 250 -2456 278 -2428
rect 316 -2456 344 -2428
rect 382 -2456 410 -2428
rect 448 -2456 476 -2428
rect 514 -2456 542 -2428
rect 580 -2456 608 -2428
rect 646 -2456 674 -2428
rect 712 -2456 740 -2428
rect -740 -2522 -712 -2494
rect -674 -2522 -646 -2494
rect -608 -2522 -580 -2494
rect -542 -2522 -514 -2494
rect -476 -2522 -448 -2494
rect -410 -2522 -382 -2494
rect -344 -2522 -316 -2494
rect -278 -2522 -250 -2494
rect -212 -2522 -184 -2494
rect -146 -2522 -118 -2494
rect -80 -2522 -52 -2494
rect -14 -2522 14 -2494
rect 52 -2522 80 -2494
rect 118 -2522 146 -2494
rect 184 -2522 212 -2494
rect 250 -2522 278 -2494
rect 316 -2522 344 -2494
rect 382 -2522 410 -2494
rect 448 -2522 476 -2494
rect 514 -2522 542 -2494
rect 580 -2522 608 -2494
rect 646 -2522 674 -2494
rect 712 -2522 740 -2494
rect -740 -2588 -712 -2560
rect -674 -2588 -646 -2560
rect -608 -2588 -580 -2560
rect -542 -2588 -514 -2560
rect -476 -2588 -448 -2560
rect -410 -2588 -382 -2560
rect -344 -2588 -316 -2560
rect -278 -2588 -250 -2560
rect -212 -2588 -184 -2560
rect -146 -2588 -118 -2560
rect -80 -2588 -52 -2560
rect -14 -2588 14 -2560
rect 52 -2588 80 -2560
rect 118 -2588 146 -2560
rect 184 -2588 212 -2560
rect 250 -2588 278 -2560
rect 316 -2588 344 -2560
rect 382 -2588 410 -2560
rect 448 -2588 476 -2560
rect 514 -2588 542 -2560
rect 580 -2588 608 -2560
rect 646 -2588 674 -2560
rect 712 -2588 740 -2560
rect -740 -2654 -712 -2626
rect -674 -2654 -646 -2626
rect -608 -2654 -580 -2626
rect -542 -2654 -514 -2626
rect -476 -2654 -448 -2626
rect -410 -2654 -382 -2626
rect -344 -2654 -316 -2626
rect -278 -2654 -250 -2626
rect -212 -2654 -184 -2626
rect -146 -2654 -118 -2626
rect -80 -2654 -52 -2626
rect -14 -2654 14 -2626
rect 52 -2654 80 -2626
rect 118 -2654 146 -2626
rect 184 -2654 212 -2626
rect 250 -2654 278 -2626
rect 316 -2654 344 -2626
rect 382 -2654 410 -2626
rect 448 -2654 476 -2626
rect 514 -2654 542 -2626
rect 580 -2654 608 -2626
rect 646 -2654 674 -2626
rect 712 -2654 740 -2626
rect -740 -2720 -712 -2692
rect -674 -2720 -646 -2692
rect -608 -2720 -580 -2692
rect -542 -2720 -514 -2692
rect -476 -2720 -448 -2692
rect -410 -2720 -382 -2692
rect -344 -2720 -316 -2692
rect -278 -2720 -250 -2692
rect -212 -2720 -184 -2692
rect -146 -2720 -118 -2692
rect -80 -2720 -52 -2692
rect -14 -2720 14 -2692
rect 52 -2720 80 -2692
rect 118 -2720 146 -2692
rect 184 -2720 212 -2692
rect 250 -2720 278 -2692
rect 316 -2720 344 -2692
rect 382 -2720 410 -2692
rect 448 -2720 476 -2692
rect 514 -2720 542 -2692
rect 580 -2720 608 -2692
rect 646 -2720 674 -2692
rect 712 -2720 740 -2692
rect -740 -2786 -712 -2758
rect -674 -2786 -646 -2758
rect -608 -2786 -580 -2758
rect -542 -2786 -514 -2758
rect -476 -2786 -448 -2758
rect -410 -2786 -382 -2758
rect -344 -2786 -316 -2758
rect -278 -2786 -250 -2758
rect -212 -2786 -184 -2758
rect -146 -2786 -118 -2758
rect -80 -2786 -52 -2758
rect -14 -2786 14 -2758
rect 52 -2786 80 -2758
rect 118 -2786 146 -2758
rect 184 -2786 212 -2758
rect 250 -2786 278 -2758
rect 316 -2786 344 -2758
rect 382 -2786 410 -2758
rect 448 -2786 476 -2758
rect 514 -2786 542 -2758
rect 580 -2786 608 -2758
rect 646 -2786 674 -2758
rect 712 -2786 740 -2758
rect -740 -2852 -712 -2824
rect -674 -2852 -646 -2824
rect -608 -2852 -580 -2824
rect -542 -2852 -514 -2824
rect -476 -2852 -448 -2824
rect -410 -2852 -382 -2824
rect -344 -2852 -316 -2824
rect -278 -2852 -250 -2824
rect -212 -2852 -184 -2824
rect -146 -2852 -118 -2824
rect -80 -2852 -52 -2824
rect -14 -2852 14 -2824
rect 52 -2852 80 -2824
rect 118 -2852 146 -2824
rect 184 -2852 212 -2824
rect 250 -2852 278 -2824
rect 316 -2852 344 -2824
rect 382 -2852 410 -2824
rect 448 -2852 476 -2824
rect 514 -2852 542 -2824
rect 580 -2852 608 -2824
rect 646 -2852 674 -2824
rect 712 -2852 740 -2824
rect -740 -2918 -712 -2890
rect -674 -2918 -646 -2890
rect -608 -2918 -580 -2890
rect -542 -2918 -514 -2890
rect -476 -2918 -448 -2890
rect -410 -2918 -382 -2890
rect -344 -2918 -316 -2890
rect -278 -2918 -250 -2890
rect -212 -2918 -184 -2890
rect -146 -2918 -118 -2890
rect -80 -2918 -52 -2890
rect -14 -2918 14 -2890
rect 52 -2918 80 -2890
rect 118 -2918 146 -2890
rect 184 -2918 212 -2890
rect 250 -2918 278 -2890
rect 316 -2918 344 -2890
rect 382 -2918 410 -2890
rect 448 -2918 476 -2890
rect 514 -2918 542 -2890
rect 580 -2918 608 -2890
rect 646 -2918 674 -2890
rect 712 -2918 740 -2890
rect -740 -2984 -712 -2956
rect -674 -2984 -646 -2956
rect -608 -2984 -580 -2956
rect -542 -2984 -514 -2956
rect -476 -2984 -448 -2956
rect -410 -2984 -382 -2956
rect -344 -2984 -316 -2956
rect -278 -2984 -250 -2956
rect -212 -2984 -184 -2956
rect -146 -2984 -118 -2956
rect -80 -2984 -52 -2956
rect -14 -2984 14 -2956
rect 52 -2984 80 -2956
rect 118 -2984 146 -2956
rect 184 -2984 212 -2956
rect 250 -2984 278 -2956
rect 316 -2984 344 -2956
rect 382 -2984 410 -2956
rect 448 -2984 476 -2956
rect 514 -2984 542 -2956
rect 580 -2984 608 -2956
rect 646 -2984 674 -2956
rect 712 -2984 740 -2956
rect -740 -3050 -712 -3022
rect -674 -3050 -646 -3022
rect -608 -3050 -580 -3022
rect -542 -3050 -514 -3022
rect -476 -3050 -448 -3022
rect -410 -3050 -382 -3022
rect -344 -3050 -316 -3022
rect -278 -3050 -250 -3022
rect -212 -3050 -184 -3022
rect -146 -3050 -118 -3022
rect -80 -3050 -52 -3022
rect -14 -3050 14 -3022
rect 52 -3050 80 -3022
rect 118 -3050 146 -3022
rect 184 -3050 212 -3022
rect 250 -3050 278 -3022
rect 316 -3050 344 -3022
rect 382 -3050 410 -3022
rect 448 -3050 476 -3022
rect 514 -3050 542 -3022
rect 580 -3050 608 -3022
rect 646 -3050 674 -3022
rect 712 -3050 740 -3022
rect -740 -3116 -712 -3088
rect -674 -3116 -646 -3088
rect -608 -3116 -580 -3088
rect -542 -3116 -514 -3088
rect -476 -3116 -448 -3088
rect -410 -3116 -382 -3088
rect -344 -3116 -316 -3088
rect -278 -3116 -250 -3088
rect -212 -3116 -184 -3088
rect -146 -3116 -118 -3088
rect -80 -3116 -52 -3088
rect -14 -3116 14 -3088
rect 52 -3116 80 -3088
rect 118 -3116 146 -3088
rect 184 -3116 212 -3088
rect 250 -3116 278 -3088
rect 316 -3116 344 -3088
rect 382 -3116 410 -3088
rect 448 -3116 476 -3088
rect 514 -3116 542 -3088
rect 580 -3116 608 -3088
rect 646 -3116 674 -3088
rect 712 -3116 740 -3088
rect -740 -3182 -712 -3154
rect -674 -3182 -646 -3154
rect -608 -3182 -580 -3154
rect -542 -3182 -514 -3154
rect -476 -3182 -448 -3154
rect -410 -3182 -382 -3154
rect -344 -3182 -316 -3154
rect -278 -3182 -250 -3154
rect -212 -3182 -184 -3154
rect -146 -3182 -118 -3154
rect -80 -3182 -52 -3154
rect -14 -3182 14 -3154
rect 52 -3182 80 -3154
rect 118 -3182 146 -3154
rect 184 -3182 212 -3154
rect 250 -3182 278 -3154
rect 316 -3182 344 -3154
rect 382 -3182 410 -3154
rect 448 -3182 476 -3154
rect 514 -3182 542 -3154
rect 580 -3182 608 -3154
rect 646 -3182 674 -3154
rect 712 -3182 740 -3154
rect -740 -3248 -712 -3220
rect -674 -3248 -646 -3220
rect -608 -3248 -580 -3220
rect -542 -3248 -514 -3220
rect -476 -3248 -448 -3220
rect -410 -3248 -382 -3220
rect -344 -3248 -316 -3220
rect -278 -3248 -250 -3220
rect -212 -3248 -184 -3220
rect -146 -3248 -118 -3220
rect -80 -3248 -52 -3220
rect -14 -3248 14 -3220
rect 52 -3248 80 -3220
rect 118 -3248 146 -3220
rect 184 -3248 212 -3220
rect 250 -3248 278 -3220
rect 316 -3248 344 -3220
rect 382 -3248 410 -3220
rect 448 -3248 476 -3220
rect 514 -3248 542 -3220
rect 580 -3248 608 -3220
rect 646 -3248 674 -3220
rect 712 -3248 740 -3220
rect -740 -3314 -712 -3286
rect -674 -3314 -646 -3286
rect -608 -3314 -580 -3286
rect -542 -3314 -514 -3286
rect -476 -3314 -448 -3286
rect -410 -3314 -382 -3286
rect -344 -3314 -316 -3286
rect -278 -3314 -250 -3286
rect -212 -3314 -184 -3286
rect -146 -3314 -118 -3286
rect -80 -3314 -52 -3286
rect -14 -3314 14 -3286
rect 52 -3314 80 -3286
rect 118 -3314 146 -3286
rect 184 -3314 212 -3286
rect 250 -3314 278 -3286
rect 316 -3314 344 -3286
rect 382 -3314 410 -3286
rect 448 -3314 476 -3286
rect 514 -3314 542 -3286
rect 580 -3314 608 -3286
rect 646 -3314 674 -3286
rect 712 -3314 740 -3286
rect -740 -3380 -712 -3352
rect -674 -3380 -646 -3352
rect -608 -3380 -580 -3352
rect -542 -3380 -514 -3352
rect -476 -3380 -448 -3352
rect -410 -3380 -382 -3352
rect -344 -3380 -316 -3352
rect -278 -3380 -250 -3352
rect -212 -3380 -184 -3352
rect -146 -3380 -118 -3352
rect -80 -3380 -52 -3352
rect -14 -3380 14 -3352
rect 52 -3380 80 -3352
rect 118 -3380 146 -3352
rect 184 -3380 212 -3352
rect 250 -3380 278 -3352
rect 316 -3380 344 -3352
rect 382 -3380 410 -3352
rect 448 -3380 476 -3352
rect 514 -3380 542 -3352
rect 580 -3380 608 -3352
rect 646 -3380 674 -3352
rect 712 -3380 740 -3352
rect -740 -3446 -712 -3418
rect -674 -3446 -646 -3418
rect -608 -3446 -580 -3418
rect -542 -3446 -514 -3418
rect -476 -3446 -448 -3418
rect -410 -3446 -382 -3418
rect -344 -3446 -316 -3418
rect -278 -3446 -250 -3418
rect -212 -3446 -184 -3418
rect -146 -3446 -118 -3418
rect -80 -3446 -52 -3418
rect -14 -3446 14 -3418
rect 52 -3446 80 -3418
rect 118 -3446 146 -3418
rect 184 -3446 212 -3418
rect 250 -3446 278 -3418
rect 316 -3446 344 -3418
rect 382 -3446 410 -3418
rect 448 -3446 476 -3418
rect 514 -3446 542 -3418
rect 580 -3446 608 -3418
rect 646 -3446 674 -3418
rect 712 -3446 740 -3418
rect -740 -3512 -712 -3484
rect -674 -3512 -646 -3484
rect -608 -3512 -580 -3484
rect -542 -3512 -514 -3484
rect -476 -3512 -448 -3484
rect -410 -3512 -382 -3484
rect -344 -3512 -316 -3484
rect -278 -3512 -250 -3484
rect -212 -3512 -184 -3484
rect -146 -3512 -118 -3484
rect -80 -3512 -52 -3484
rect -14 -3512 14 -3484
rect 52 -3512 80 -3484
rect 118 -3512 146 -3484
rect 184 -3512 212 -3484
rect 250 -3512 278 -3484
rect 316 -3512 344 -3484
rect 382 -3512 410 -3484
rect 448 -3512 476 -3484
rect 514 -3512 542 -3484
rect 580 -3512 608 -3484
rect 646 -3512 674 -3484
rect 712 -3512 740 -3484
rect -740 -3578 -712 -3550
rect -674 -3578 -646 -3550
rect -608 -3578 -580 -3550
rect -542 -3578 -514 -3550
rect -476 -3578 -448 -3550
rect -410 -3578 -382 -3550
rect -344 -3578 -316 -3550
rect -278 -3578 -250 -3550
rect -212 -3578 -184 -3550
rect -146 -3578 -118 -3550
rect -80 -3578 -52 -3550
rect -14 -3578 14 -3550
rect 52 -3578 80 -3550
rect 118 -3578 146 -3550
rect 184 -3578 212 -3550
rect 250 -3578 278 -3550
rect 316 -3578 344 -3550
rect 382 -3578 410 -3550
rect 448 -3578 476 -3550
rect 514 -3578 542 -3550
rect 580 -3578 608 -3550
rect 646 -3578 674 -3550
rect 712 -3578 740 -3550
rect -740 -3644 -712 -3616
rect -674 -3644 -646 -3616
rect -608 -3644 -580 -3616
rect -542 -3644 -514 -3616
rect -476 -3644 -448 -3616
rect -410 -3644 -382 -3616
rect -344 -3644 -316 -3616
rect -278 -3644 -250 -3616
rect -212 -3644 -184 -3616
rect -146 -3644 -118 -3616
rect -80 -3644 -52 -3616
rect -14 -3644 14 -3616
rect 52 -3644 80 -3616
rect 118 -3644 146 -3616
rect 184 -3644 212 -3616
rect 250 -3644 278 -3616
rect 316 -3644 344 -3616
rect 382 -3644 410 -3616
rect 448 -3644 476 -3616
rect 514 -3644 542 -3616
rect 580 -3644 608 -3616
rect 646 -3644 674 -3616
rect 712 -3644 740 -3616
rect -740 -3710 -712 -3682
rect -674 -3710 -646 -3682
rect -608 -3710 -580 -3682
rect -542 -3710 -514 -3682
rect -476 -3710 -448 -3682
rect -410 -3710 -382 -3682
rect -344 -3710 -316 -3682
rect -278 -3710 -250 -3682
rect -212 -3710 -184 -3682
rect -146 -3710 -118 -3682
rect -80 -3710 -52 -3682
rect -14 -3710 14 -3682
rect 52 -3710 80 -3682
rect 118 -3710 146 -3682
rect 184 -3710 212 -3682
rect 250 -3710 278 -3682
rect 316 -3710 344 -3682
rect 382 -3710 410 -3682
rect 448 -3710 476 -3682
rect 514 -3710 542 -3682
rect 580 -3710 608 -3682
rect 646 -3710 674 -3682
rect 712 -3710 740 -3682
rect -740 -3776 -712 -3748
rect -674 -3776 -646 -3748
rect -608 -3776 -580 -3748
rect -542 -3776 -514 -3748
rect -476 -3776 -448 -3748
rect -410 -3776 -382 -3748
rect -344 -3776 -316 -3748
rect -278 -3776 -250 -3748
rect -212 -3776 -184 -3748
rect -146 -3776 -118 -3748
rect -80 -3776 -52 -3748
rect -14 -3776 14 -3748
rect 52 -3776 80 -3748
rect 118 -3776 146 -3748
rect 184 -3776 212 -3748
rect 250 -3776 278 -3748
rect 316 -3776 344 -3748
rect 382 -3776 410 -3748
rect 448 -3776 476 -3748
rect 514 -3776 542 -3748
rect 580 -3776 608 -3748
rect 646 -3776 674 -3748
rect 712 -3776 740 -3748
rect -740 -3842 -712 -3814
rect -674 -3842 -646 -3814
rect -608 -3842 -580 -3814
rect -542 -3842 -514 -3814
rect -476 -3842 -448 -3814
rect -410 -3842 -382 -3814
rect -344 -3842 -316 -3814
rect -278 -3842 -250 -3814
rect -212 -3842 -184 -3814
rect -146 -3842 -118 -3814
rect -80 -3842 -52 -3814
rect -14 -3842 14 -3814
rect 52 -3842 80 -3814
rect 118 -3842 146 -3814
rect 184 -3842 212 -3814
rect 250 -3842 278 -3814
rect 316 -3842 344 -3814
rect 382 -3842 410 -3814
rect 448 -3842 476 -3814
rect 514 -3842 542 -3814
rect 580 -3842 608 -3814
rect 646 -3842 674 -3814
rect 712 -3842 740 -3814
rect -740 -3908 -712 -3880
rect -674 -3908 -646 -3880
rect -608 -3908 -580 -3880
rect -542 -3908 -514 -3880
rect -476 -3908 -448 -3880
rect -410 -3908 -382 -3880
rect -344 -3908 -316 -3880
rect -278 -3908 -250 -3880
rect -212 -3908 -184 -3880
rect -146 -3908 -118 -3880
rect -80 -3908 -52 -3880
rect -14 -3908 14 -3880
rect 52 -3908 80 -3880
rect 118 -3908 146 -3880
rect 184 -3908 212 -3880
rect 250 -3908 278 -3880
rect 316 -3908 344 -3880
rect 382 -3908 410 -3880
rect 448 -3908 476 -3880
rect 514 -3908 542 -3880
rect 580 -3908 608 -3880
rect 646 -3908 674 -3880
rect 712 -3908 740 -3880
rect -740 -3974 -712 -3946
rect -674 -3974 -646 -3946
rect -608 -3974 -580 -3946
rect -542 -3974 -514 -3946
rect -476 -3974 -448 -3946
rect -410 -3974 -382 -3946
rect -344 -3974 -316 -3946
rect -278 -3974 -250 -3946
rect -212 -3974 -184 -3946
rect -146 -3974 -118 -3946
rect -80 -3974 -52 -3946
rect -14 -3974 14 -3946
rect 52 -3974 80 -3946
rect 118 -3974 146 -3946
rect 184 -3974 212 -3946
rect 250 -3974 278 -3946
rect 316 -3974 344 -3946
rect 382 -3974 410 -3946
rect 448 -3974 476 -3946
rect 514 -3974 542 -3946
rect 580 -3974 608 -3946
rect 646 -3974 674 -3946
rect 712 -3974 740 -3946
rect -740 -4040 -712 -4012
rect -674 -4040 -646 -4012
rect -608 -4040 -580 -4012
rect -542 -4040 -514 -4012
rect -476 -4040 -448 -4012
rect -410 -4040 -382 -4012
rect -344 -4040 -316 -4012
rect -278 -4040 -250 -4012
rect -212 -4040 -184 -4012
rect -146 -4040 -118 -4012
rect -80 -4040 -52 -4012
rect -14 -4040 14 -4012
rect 52 -4040 80 -4012
rect 118 -4040 146 -4012
rect 184 -4040 212 -4012
rect 250 -4040 278 -4012
rect 316 -4040 344 -4012
rect 382 -4040 410 -4012
rect 448 -4040 476 -4012
rect 514 -4040 542 -4012
rect 580 -4040 608 -4012
rect 646 -4040 674 -4012
rect 712 -4040 740 -4012
rect -740 -4106 -712 -4078
rect -674 -4106 -646 -4078
rect -608 -4106 -580 -4078
rect -542 -4106 -514 -4078
rect -476 -4106 -448 -4078
rect -410 -4106 -382 -4078
rect -344 -4106 -316 -4078
rect -278 -4106 -250 -4078
rect -212 -4106 -184 -4078
rect -146 -4106 -118 -4078
rect -80 -4106 -52 -4078
rect -14 -4106 14 -4078
rect 52 -4106 80 -4078
rect 118 -4106 146 -4078
rect 184 -4106 212 -4078
rect 250 -4106 278 -4078
rect 316 -4106 344 -4078
rect 382 -4106 410 -4078
rect 448 -4106 476 -4078
rect 514 -4106 542 -4078
rect 580 -4106 608 -4078
rect 646 -4106 674 -4078
rect 712 -4106 740 -4078
rect -740 -4172 -712 -4144
rect -674 -4172 -646 -4144
rect -608 -4172 -580 -4144
rect -542 -4172 -514 -4144
rect -476 -4172 -448 -4144
rect -410 -4172 -382 -4144
rect -344 -4172 -316 -4144
rect -278 -4172 -250 -4144
rect -212 -4172 -184 -4144
rect -146 -4172 -118 -4144
rect -80 -4172 -52 -4144
rect -14 -4172 14 -4144
rect 52 -4172 80 -4144
rect 118 -4172 146 -4144
rect 184 -4172 212 -4144
rect 250 -4172 278 -4144
rect 316 -4172 344 -4144
rect 382 -4172 410 -4144
rect 448 -4172 476 -4144
rect 514 -4172 542 -4144
rect 580 -4172 608 -4144
rect 646 -4172 674 -4144
rect 712 -4172 740 -4144
rect -740 -4238 -712 -4210
rect -674 -4238 -646 -4210
rect -608 -4238 -580 -4210
rect -542 -4238 -514 -4210
rect -476 -4238 -448 -4210
rect -410 -4238 -382 -4210
rect -344 -4238 -316 -4210
rect -278 -4238 -250 -4210
rect -212 -4238 -184 -4210
rect -146 -4238 -118 -4210
rect -80 -4238 -52 -4210
rect -14 -4238 14 -4210
rect 52 -4238 80 -4210
rect 118 -4238 146 -4210
rect 184 -4238 212 -4210
rect 250 -4238 278 -4210
rect 316 -4238 344 -4210
rect 382 -4238 410 -4210
rect 448 -4238 476 -4210
rect 514 -4238 542 -4210
rect 580 -4238 608 -4210
rect 646 -4238 674 -4210
rect 712 -4238 740 -4210
rect -740 -4304 -712 -4276
rect -674 -4304 -646 -4276
rect -608 -4304 -580 -4276
rect -542 -4304 -514 -4276
rect -476 -4304 -448 -4276
rect -410 -4304 -382 -4276
rect -344 -4304 -316 -4276
rect -278 -4304 -250 -4276
rect -212 -4304 -184 -4276
rect -146 -4304 -118 -4276
rect -80 -4304 -52 -4276
rect -14 -4304 14 -4276
rect 52 -4304 80 -4276
rect 118 -4304 146 -4276
rect 184 -4304 212 -4276
rect 250 -4304 278 -4276
rect 316 -4304 344 -4276
rect 382 -4304 410 -4276
rect 448 -4304 476 -4276
rect 514 -4304 542 -4276
rect 580 -4304 608 -4276
rect 646 -4304 674 -4276
rect 712 -4304 740 -4276
rect -740 -4370 -712 -4342
rect -674 -4370 -646 -4342
rect -608 -4370 -580 -4342
rect -542 -4370 -514 -4342
rect -476 -4370 -448 -4342
rect -410 -4370 -382 -4342
rect -344 -4370 -316 -4342
rect -278 -4370 -250 -4342
rect -212 -4370 -184 -4342
rect -146 -4370 -118 -4342
rect -80 -4370 -52 -4342
rect -14 -4370 14 -4342
rect 52 -4370 80 -4342
rect 118 -4370 146 -4342
rect 184 -4370 212 -4342
rect 250 -4370 278 -4342
rect 316 -4370 344 -4342
rect 382 -4370 410 -4342
rect 448 -4370 476 -4342
rect 514 -4370 542 -4342
rect 580 -4370 608 -4342
rect 646 -4370 674 -4342
rect 712 -4370 740 -4342
rect -740 -4436 -712 -4408
rect -674 -4436 -646 -4408
rect -608 -4436 -580 -4408
rect -542 -4436 -514 -4408
rect -476 -4436 -448 -4408
rect -410 -4436 -382 -4408
rect -344 -4436 -316 -4408
rect -278 -4436 -250 -4408
rect -212 -4436 -184 -4408
rect -146 -4436 -118 -4408
rect -80 -4436 -52 -4408
rect -14 -4436 14 -4408
rect 52 -4436 80 -4408
rect 118 -4436 146 -4408
rect 184 -4436 212 -4408
rect 250 -4436 278 -4408
rect 316 -4436 344 -4408
rect 382 -4436 410 -4408
rect 448 -4436 476 -4408
rect 514 -4436 542 -4408
rect 580 -4436 608 -4408
rect 646 -4436 674 -4408
rect 712 -4436 740 -4408
rect -740 -4502 -712 -4474
rect -674 -4502 -646 -4474
rect -608 -4502 -580 -4474
rect -542 -4502 -514 -4474
rect -476 -4502 -448 -4474
rect -410 -4502 -382 -4474
rect -344 -4502 -316 -4474
rect -278 -4502 -250 -4474
rect -212 -4502 -184 -4474
rect -146 -4502 -118 -4474
rect -80 -4502 -52 -4474
rect -14 -4502 14 -4474
rect 52 -4502 80 -4474
rect 118 -4502 146 -4474
rect 184 -4502 212 -4474
rect 250 -4502 278 -4474
rect 316 -4502 344 -4474
rect 382 -4502 410 -4474
rect 448 -4502 476 -4474
rect 514 -4502 542 -4474
rect 580 -4502 608 -4474
rect 646 -4502 674 -4474
rect 712 -4502 740 -4474
rect -740 -4568 -712 -4540
rect -674 -4568 -646 -4540
rect -608 -4568 -580 -4540
rect -542 -4568 -514 -4540
rect -476 -4568 -448 -4540
rect -410 -4568 -382 -4540
rect -344 -4568 -316 -4540
rect -278 -4568 -250 -4540
rect -212 -4568 -184 -4540
rect -146 -4568 -118 -4540
rect -80 -4568 -52 -4540
rect -14 -4568 14 -4540
rect 52 -4568 80 -4540
rect 118 -4568 146 -4540
rect 184 -4568 212 -4540
rect 250 -4568 278 -4540
rect 316 -4568 344 -4540
rect 382 -4568 410 -4540
rect 448 -4568 476 -4540
rect 514 -4568 542 -4540
rect 580 -4568 608 -4540
rect 646 -4568 674 -4540
rect 712 -4568 740 -4540
rect -740 -4634 -712 -4606
rect -674 -4634 -646 -4606
rect -608 -4634 -580 -4606
rect -542 -4634 -514 -4606
rect -476 -4634 -448 -4606
rect -410 -4634 -382 -4606
rect -344 -4634 -316 -4606
rect -278 -4634 -250 -4606
rect -212 -4634 -184 -4606
rect -146 -4634 -118 -4606
rect -80 -4634 -52 -4606
rect -14 -4634 14 -4606
rect 52 -4634 80 -4606
rect 118 -4634 146 -4606
rect 184 -4634 212 -4606
rect 250 -4634 278 -4606
rect 316 -4634 344 -4606
rect 382 -4634 410 -4606
rect 448 -4634 476 -4606
rect 514 -4634 542 -4606
rect 580 -4634 608 -4606
rect 646 -4634 674 -4606
rect 712 -4634 740 -4606
rect -740 -4700 -712 -4672
rect -674 -4700 -646 -4672
rect -608 -4700 -580 -4672
rect -542 -4700 -514 -4672
rect -476 -4700 -448 -4672
rect -410 -4700 -382 -4672
rect -344 -4700 -316 -4672
rect -278 -4700 -250 -4672
rect -212 -4700 -184 -4672
rect -146 -4700 -118 -4672
rect -80 -4700 -52 -4672
rect -14 -4700 14 -4672
rect 52 -4700 80 -4672
rect 118 -4700 146 -4672
rect 184 -4700 212 -4672
rect 250 -4700 278 -4672
rect 316 -4700 344 -4672
rect 382 -4700 410 -4672
rect 448 -4700 476 -4672
rect 514 -4700 542 -4672
rect 580 -4700 608 -4672
rect 646 -4700 674 -4672
rect 712 -4700 740 -4672
rect -740 -4766 -712 -4738
rect -674 -4766 -646 -4738
rect -608 -4766 -580 -4738
rect -542 -4766 -514 -4738
rect -476 -4766 -448 -4738
rect -410 -4766 -382 -4738
rect -344 -4766 -316 -4738
rect -278 -4766 -250 -4738
rect -212 -4766 -184 -4738
rect -146 -4766 -118 -4738
rect -80 -4766 -52 -4738
rect -14 -4766 14 -4738
rect 52 -4766 80 -4738
rect 118 -4766 146 -4738
rect 184 -4766 212 -4738
rect 250 -4766 278 -4738
rect 316 -4766 344 -4738
rect 382 -4766 410 -4738
rect 448 -4766 476 -4738
rect 514 -4766 542 -4738
rect 580 -4766 608 -4738
rect 646 -4766 674 -4738
rect 712 -4766 740 -4738
rect -740 -4832 -712 -4804
rect -674 -4832 -646 -4804
rect -608 -4832 -580 -4804
rect -542 -4832 -514 -4804
rect -476 -4832 -448 -4804
rect -410 -4832 -382 -4804
rect -344 -4832 -316 -4804
rect -278 -4832 -250 -4804
rect -212 -4832 -184 -4804
rect -146 -4832 -118 -4804
rect -80 -4832 -52 -4804
rect -14 -4832 14 -4804
rect 52 -4832 80 -4804
rect 118 -4832 146 -4804
rect 184 -4832 212 -4804
rect 250 -4832 278 -4804
rect 316 -4832 344 -4804
rect 382 -4832 410 -4804
rect 448 -4832 476 -4804
rect 514 -4832 542 -4804
rect 580 -4832 608 -4804
rect 646 -4832 674 -4804
rect 712 -4832 740 -4804
rect -740 -4898 -712 -4870
rect -674 -4898 -646 -4870
rect -608 -4898 -580 -4870
rect -542 -4898 -514 -4870
rect -476 -4898 -448 -4870
rect -410 -4898 -382 -4870
rect -344 -4898 -316 -4870
rect -278 -4898 -250 -4870
rect -212 -4898 -184 -4870
rect -146 -4898 -118 -4870
rect -80 -4898 -52 -4870
rect -14 -4898 14 -4870
rect 52 -4898 80 -4870
rect 118 -4898 146 -4870
rect 184 -4898 212 -4870
rect 250 -4898 278 -4870
rect 316 -4898 344 -4870
rect 382 -4898 410 -4870
rect 448 -4898 476 -4870
rect 514 -4898 542 -4870
rect 580 -4898 608 -4870
rect 646 -4898 674 -4870
rect 712 -4898 740 -4870
rect -740 -4964 -712 -4936
rect -674 -4964 -646 -4936
rect -608 -4964 -580 -4936
rect -542 -4964 -514 -4936
rect -476 -4964 -448 -4936
rect -410 -4964 -382 -4936
rect -344 -4964 -316 -4936
rect -278 -4964 -250 -4936
rect -212 -4964 -184 -4936
rect -146 -4964 -118 -4936
rect -80 -4964 -52 -4936
rect -14 -4964 14 -4936
rect 52 -4964 80 -4936
rect 118 -4964 146 -4936
rect 184 -4964 212 -4936
rect 250 -4964 278 -4936
rect 316 -4964 344 -4936
rect 382 -4964 410 -4936
rect 448 -4964 476 -4936
rect 514 -4964 542 -4936
rect 580 -4964 608 -4936
rect 646 -4964 674 -4936
rect 712 -4964 740 -4936
rect -740 -5030 -712 -5002
rect -674 -5030 -646 -5002
rect -608 -5030 -580 -5002
rect -542 -5030 -514 -5002
rect -476 -5030 -448 -5002
rect -410 -5030 -382 -5002
rect -344 -5030 -316 -5002
rect -278 -5030 -250 -5002
rect -212 -5030 -184 -5002
rect -146 -5030 -118 -5002
rect -80 -5030 -52 -5002
rect -14 -5030 14 -5002
rect 52 -5030 80 -5002
rect 118 -5030 146 -5002
rect 184 -5030 212 -5002
rect 250 -5030 278 -5002
rect 316 -5030 344 -5002
rect 382 -5030 410 -5002
rect 448 -5030 476 -5002
rect 514 -5030 542 -5002
rect 580 -5030 608 -5002
rect 646 -5030 674 -5002
rect 712 -5030 740 -5002
rect -740 -5096 -712 -5068
rect -674 -5096 -646 -5068
rect -608 -5096 -580 -5068
rect -542 -5096 -514 -5068
rect -476 -5096 -448 -5068
rect -410 -5096 -382 -5068
rect -344 -5096 -316 -5068
rect -278 -5096 -250 -5068
rect -212 -5096 -184 -5068
rect -146 -5096 -118 -5068
rect -80 -5096 -52 -5068
rect -14 -5096 14 -5068
rect 52 -5096 80 -5068
rect 118 -5096 146 -5068
rect 184 -5096 212 -5068
rect 250 -5096 278 -5068
rect 316 -5096 344 -5068
rect 382 -5096 410 -5068
rect 448 -5096 476 -5068
rect 514 -5096 542 -5068
rect 580 -5096 608 -5068
rect 646 -5096 674 -5068
rect 712 -5096 740 -5068
rect -740 -5162 -712 -5134
rect -674 -5162 -646 -5134
rect -608 -5162 -580 -5134
rect -542 -5162 -514 -5134
rect -476 -5162 -448 -5134
rect -410 -5162 -382 -5134
rect -344 -5162 -316 -5134
rect -278 -5162 -250 -5134
rect -212 -5162 -184 -5134
rect -146 -5162 -118 -5134
rect -80 -5162 -52 -5134
rect -14 -5162 14 -5134
rect 52 -5162 80 -5134
rect 118 -5162 146 -5134
rect 184 -5162 212 -5134
rect 250 -5162 278 -5134
rect 316 -5162 344 -5134
rect 382 -5162 410 -5134
rect 448 -5162 476 -5134
rect 514 -5162 542 -5134
rect 580 -5162 608 -5134
rect 646 -5162 674 -5134
rect 712 -5162 740 -5134
rect -740 -5228 -712 -5200
rect -674 -5228 -646 -5200
rect -608 -5228 -580 -5200
rect -542 -5228 -514 -5200
rect -476 -5228 -448 -5200
rect -410 -5228 -382 -5200
rect -344 -5228 -316 -5200
rect -278 -5228 -250 -5200
rect -212 -5228 -184 -5200
rect -146 -5228 -118 -5200
rect -80 -5228 -52 -5200
rect -14 -5228 14 -5200
rect 52 -5228 80 -5200
rect 118 -5228 146 -5200
rect 184 -5228 212 -5200
rect 250 -5228 278 -5200
rect 316 -5228 344 -5200
rect 382 -5228 410 -5200
rect 448 -5228 476 -5200
rect 514 -5228 542 -5200
rect 580 -5228 608 -5200
rect 646 -5228 674 -5200
rect 712 -5228 740 -5200
rect -740 -5294 -712 -5266
rect -674 -5294 -646 -5266
rect -608 -5294 -580 -5266
rect -542 -5294 -514 -5266
rect -476 -5294 -448 -5266
rect -410 -5294 -382 -5266
rect -344 -5294 -316 -5266
rect -278 -5294 -250 -5266
rect -212 -5294 -184 -5266
rect -146 -5294 -118 -5266
rect -80 -5294 -52 -5266
rect -14 -5294 14 -5266
rect 52 -5294 80 -5266
rect 118 -5294 146 -5266
rect 184 -5294 212 -5266
rect 250 -5294 278 -5266
rect 316 -5294 344 -5266
rect 382 -5294 410 -5266
rect 448 -5294 476 -5266
rect 514 -5294 542 -5266
rect 580 -5294 608 -5266
rect 646 -5294 674 -5266
rect 712 -5294 740 -5266
rect -740 -5360 -712 -5332
rect -674 -5360 -646 -5332
rect -608 -5360 -580 -5332
rect -542 -5360 -514 -5332
rect -476 -5360 -448 -5332
rect -410 -5360 -382 -5332
rect -344 -5360 -316 -5332
rect -278 -5360 -250 -5332
rect -212 -5360 -184 -5332
rect -146 -5360 -118 -5332
rect -80 -5360 -52 -5332
rect -14 -5360 14 -5332
rect 52 -5360 80 -5332
rect 118 -5360 146 -5332
rect 184 -5360 212 -5332
rect 250 -5360 278 -5332
rect 316 -5360 344 -5332
rect 382 -5360 410 -5332
rect 448 -5360 476 -5332
rect 514 -5360 542 -5332
rect 580 -5360 608 -5332
rect 646 -5360 674 -5332
rect 712 -5360 740 -5332
rect -740 -5426 -712 -5398
rect -674 -5426 -646 -5398
rect -608 -5426 -580 -5398
rect -542 -5426 -514 -5398
rect -476 -5426 -448 -5398
rect -410 -5426 -382 -5398
rect -344 -5426 -316 -5398
rect -278 -5426 -250 -5398
rect -212 -5426 -184 -5398
rect -146 -5426 -118 -5398
rect -80 -5426 -52 -5398
rect -14 -5426 14 -5398
rect 52 -5426 80 -5398
rect 118 -5426 146 -5398
rect 184 -5426 212 -5398
rect 250 -5426 278 -5398
rect 316 -5426 344 -5398
rect 382 -5426 410 -5398
rect 448 -5426 476 -5398
rect 514 -5426 542 -5398
rect 580 -5426 608 -5398
rect 646 -5426 674 -5398
rect 712 -5426 740 -5398
rect -740 -5492 -712 -5464
rect -674 -5492 -646 -5464
rect -608 -5492 -580 -5464
rect -542 -5492 -514 -5464
rect -476 -5492 -448 -5464
rect -410 -5492 -382 -5464
rect -344 -5492 -316 -5464
rect -278 -5492 -250 -5464
rect -212 -5492 -184 -5464
rect -146 -5492 -118 -5464
rect -80 -5492 -52 -5464
rect -14 -5492 14 -5464
rect 52 -5492 80 -5464
rect 118 -5492 146 -5464
rect 184 -5492 212 -5464
rect 250 -5492 278 -5464
rect 316 -5492 344 -5464
rect 382 -5492 410 -5464
rect 448 -5492 476 -5464
rect 514 -5492 542 -5464
rect 580 -5492 608 -5464
rect 646 -5492 674 -5464
rect 712 -5492 740 -5464
rect -740 -5558 -712 -5530
rect -674 -5558 -646 -5530
rect -608 -5558 -580 -5530
rect -542 -5558 -514 -5530
rect -476 -5558 -448 -5530
rect -410 -5558 -382 -5530
rect -344 -5558 -316 -5530
rect -278 -5558 -250 -5530
rect -212 -5558 -184 -5530
rect -146 -5558 -118 -5530
rect -80 -5558 -52 -5530
rect -14 -5558 14 -5530
rect 52 -5558 80 -5530
rect 118 -5558 146 -5530
rect 184 -5558 212 -5530
rect 250 -5558 278 -5530
rect 316 -5558 344 -5530
rect 382 -5558 410 -5530
rect 448 -5558 476 -5530
rect 514 -5558 542 -5530
rect 580 -5558 608 -5530
rect 646 -5558 674 -5530
rect 712 -5558 740 -5530
<< metal4 >>
rect -745 5558 745 5563
rect -745 5530 -740 5558
rect -712 5530 -674 5558
rect -646 5530 -608 5558
rect -580 5530 -542 5558
rect -514 5530 -476 5558
rect -448 5530 -410 5558
rect -382 5530 -344 5558
rect -316 5530 -278 5558
rect -250 5530 -212 5558
rect -184 5530 -146 5558
rect -118 5530 -80 5558
rect -52 5530 -14 5558
rect 14 5530 52 5558
rect 80 5530 118 5558
rect 146 5530 184 5558
rect 212 5530 250 5558
rect 278 5530 316 5558
rect 344 5530 382 5558
rect 410 5530 448 5558
rect 476 5530 514 5558
rect 542 5530 580 5558
rect 608 5530 646 5558
rect 674 5530 712 5558
rect 740 5530 745 5558
rect -745 5492 745 5530
rect -745 5464 -740 5492
rect -712 5464 -674 5492
rect -646 5464 -608 5492
rect -580 5464 -542 5492
rect -514 5464 -476 5492
rect -448 5464 -410 5492
rect -382 5464 -344 5492
rect -316 5464 -278 5492
rect -250 5464 -212 5492
rect -184 5464 -146 5492
rect -118 5464 -80 5492
rect -52 5464 -14 5492
rect 14 5464 52 5492
rect 80 5464 118 5492
rect 146 5464 184 5492
rect 212 5464 250 5492
rect 278 5464 316 5492
rect 344 5464 382 5492
rect 410 5464 448 5492
rect 476 5464 514 5492
rect 542 5464 580 5492
rect 608 5464 646 5492
rect 674 5464 712 5492
rect 740 5464 745 5492
rect -745 5426 745 5464
rect -745 5398 -740 5426
rect -712 5398 -674 5426
rect -646 5398 -608 5426
rect -580 5398 -542 5426
rect -514 5398 -476 5426
rect -448 5398 -410 5426
rect -382 5398 -344 5426
rect -316 5398 -278 5426
rect -250 5398 -212 5426
rect -184 5398 -146 5426
rect -118 5398 -80 5426
rect -52 5398 -14 5426
rect 14 5398 52 5426
rect 80 5398 118 5426
rect 146 5398 184 5426
rect 212 5398 250 5426
rect 278 5398 316 5426
rect 344 5398 382 5426
rect 410 5398 448 5426
rect 476 5398 514 5426
rect 542 5398 580 5426
rect 608 5398 646 5426
rect 674 5398 712 5426
rect 740 5398 745 5426
rect -745 5360 745 5398
rect -745 5332 -740 5360
rect -712 5332 -674 5360
rect -646 5332 -608 5360
rect -580 5332 -542 5360
rect -514 5332 -476 5360
rect -448 5332 -410 5360
rect -382 5332 -344 5360
rect -316 5332 -278 5360
rect -250 5332 -212 5360
rect -184 5332 -146 5360
rect -118 5332 -80 5360
rect -52 5332 -14 5360
rect 14 5332 52 5360
rect 80 5332 118 5360
rect 146 5332 184 5360
rect 212 5332 250 5360
rect 278 5332 316 5360
rect 344 5332 382 5360
rect 410 5332 448 5360
rect 476 5332 514 5360
rect 542 5332 580 5360
rect 608 5332 646 5360
rect 674 5332 712 5360
rect 740 5332 745 5360
rect -745 5294 745 5332
rect -745 5266 -740 5294
rect -712 5266 -674 5294
rect -646 5266 -608 5294
rect -580 5266 -542 5294
rect -514 5266 -476 5294
rect -448 5266 -410 5294
rect -382 5266 -344 5294
rect -316 5266 -278 5294
rect -250 5266 -212 5294
rect -184 5266 -146 5294
rect -118 5266 -80 5294
rect -52 5266 -14 5294
rect 14 5266 52 5294
rect 80 5266 118 5294
rect 146 5266 184 5294
rect 212 5266 250 5294
rect 278 5266 316 5294
rect 344 5266 382 5294
rect 410 5266 448 5294
rect 476 5266 514 5294
rect 542 5266 580 5294
rect 608 5266 646 5294
rect 674 5266 712 5294
rect 740 5266 745 5294
rect -745 5228 745 5266
rect -745 5200 -740 5228
rect -712 5200 -674 5228
rect -646 5200 -608 5228
rect -580 5200 -542 5228
rect -514 5200 -476 5228
rect -448 5200 -410 5228
rect -382 5200 -344 5228
rect -316 5200 -278 5228
rect -250 5200 -212 5228
rect -184 5200 -146 5228
rect -118 5200 -80 5228
rect -52 5200 -14 5228
rect 14 5200 52 5228
rect 80 5200 118 5228
rect 146 5200 184 5228
rect 212 5200 250 5228
rect 278 5200 316 5228
rect 344 5200 382 5228
rect 410 5200 448 5228
rect 476 5200 514 5228
rect 542 5200 580 5228
rect 608 5200 646 5228
rect 674 5200 712 5228
rect 740 5200 745 5228
rect -745 5162 745 5200
rect -745 5134 -740 5162
rect -712 5134 -674 5162
rect -646 5134 -608 5162
rect -580 5134 -542 5162
rect -514 5134 -476 5162
rect -448 5134 -410 5162
rect -382 5134 -344 5162
rect -316 5134 -278 5162
rect -250 5134 -212 5162
rect -184 5134 -146 5162
rect -118 5134 -80 5162
rect -52 5134 -14 5162
rect 14 5134 52 5162
rect 80 5134 118 5162
rect 146 5134 184 5162
rect 212 5134 250 5162
rect 278 5134 316 5162
rect 344 5134 382 5162
rect 410 5134 448 5162
rect 476 5134 514 5162
rect 542 5134 580 5162
rect 608 5134 646 5162
rect 674 5134 712 5162
rect 740 5134 745 5162
rect -745 5096 745 5134
rect -745 5068 -740 5096
rect -712 5068 -674 5096
rect -646 5068 -608 5096
rect -580 5068 -542 5096
rect -514 5068 -476 5096
rect -448 5068 -410 5096
rect -382 5068 -344 5096
rect -316 5068 -278 5096
rect -250 5068 -212 5096
rect -184 5068 -146 5096
rect -118 5068 -80 5096
rect -52 5068 -14 5096
rect 14 5068 52 5096
rect 80 5068 118 5096
rect 146 5068 184 5096
rect 212 5068 250 5096
rect 278 5068 316 5096
rect 344 5068 382 5096
rect 410 5068 448 5096
rect 476 5068 514 5096
rect 542 5068 580 5096
rect 608 5068 646 5096
rect 674 5068 712 5096
rect 740 5068 745 5096
rect -745 5030 745 5068
rect -745 5002 -740 5030
rect -712 5002 -674 5030
rect -646 5002 -608 5030
rect -580 5002 -542 5030
rect -514 5002 -476 5030
rect -448 5002 -410 5030
rect -382 5002 -344 5030
rect -316 5002 -278 5030
rect -250 5002 -212 5030
rect -184 5002 -146 5030
rect -118 5002 -80 5030
rect -52 5002 -14 5030
rect 14 5002 52 5030
rect 80 5002 118 5030
rect 146 5002 184 5030
rect 212 5002 250 5030
rect 278 5002 316 5030
rect 344 5002 382 5030
rect 410 5002 448 5030
rect 476 5002 514 5030
rect 542 5002 580 5030
rect 608 5002 646 5030
rect 674 5002 712 5030
rect 740 5002 745 5030
rect -745 4964 745 5002
rect -745 4936 -740 4964
rect -712 4936 -674 4964
rect -646 4936 -608 4964
rect -580 4936 -542 4964
rect -514 4936 -476 4964
rect -448 4936 -410 4964
rect -382 4936 -344 4964
rect -316 4936 -278 4964
rect -250 4936 -212 4964
rect -184 4936 -146 4964
rect -118 4936 -80 4964
rect -52 4936 -14 4964
rect 14 4936 52 4964
rect 80 4936 118 4964
rect 146 4936 184 4964
rect 212 4936 250 4964
rect 278 4936 316 4964
rect 344 4936 382 4964
rect 410 4936 448 4964
rect 476 4936 514 4964
rect 542 4936 580 4964
rect 608 4936 646 4964
rect 674 4936 712 4964
rect 740 4936 745 4964
rect -745 4898 745 4936
rect -745 4870 -740 4898
rect -712 4870 -674 4898
rect -646 4870 -608 4898
rect -580 4870 -542 4898
rect -514 4870 -476 4898
rect -448 4870 -410 4898
rect -382 4870 -344 4898
rect -316 4870 -278 4898
rect -250 4870 -212 4898
rect -184 4870 -146 4898
rect -118 4870 -80 4898
rect -52 4870 -14 4898
rect 14 4870 52 4898
rect 80 4870 118 4898
rect 146 4870 184 4898
rect 212 4870 250 4898
rect 278 4870 316 4898
rect 344 4870 382 4898
rect 410 4870 448 4898
rect 476 4870 514 4898
rect 542 4870 580 4898
rect 608 4870 646 4898
rect 674 4870 712 4898
rect 740 4870 745 4898
rect -745 4832 745 4870
rect -745 4804 -740 4832
rect -712 4804 -674 4832
rect -646 4804 -608 4832
rect -580 4804 -542 4832
rect -514 4804 -476 4832
rect -448 4804 -410 4832
rect -382 4804 -344 4832
rect -316 4804 -278 4832
rect -250 4804 -212 4832
rect -184 4804 -146 4832
rect -118 4804 -80 4832
rect -52 4804 -14 4832
rect 14 4804 52 4832
rect 80 4804 118 4832
rect 146 4804 184 4832
rect 212 4804 250 4832
rect 278 4804 316 4832
rect 344 4804 382 4832
rect 410 4804 448 4832
rect 476 4804 514 4832
rect 542 4804 580 4832
rect 608 4804 646 4832
rect 674 4804 712 4832
rect 740 4804 745 4832
rect -745 4766 745 4804
rect -745 4738 -740 4766
rect -712 4738 -674 4766
rect -646 4738 -608 4766
rect -580 4738 -542 4766
rect -514 4738 -476 4766
rect -448 4738 -410 4766
rect -382 4738 -344 4766
rect -316 4738 -278 4766
rect -250 4738 -212 4766
rect -184 4738 -146 4766
rect -118 4738 -80 4766
rect -52 4738 -14 4766
rect 14 4738 52 4766
rect 80 4738 118 4766
rect 146 4738 184 4766
rect 212 4738 250 4766
rect 278 4738 316 4766
rect 344 4738 382 4766
rect 410 4738 448 4766
rect 476 4738 514 4766
rect 542 4738 580 4766
rect 608 4738 646 4766
rect 674 4738 712 4766
rect 740 4738 745 4766
rect -745 4700 745 4738
rect -745 4672 -740 4700
rect -712 4672 -674 4700
rect -646 4672 -608 4700
rect -580 4672 -542 4700
rect -514 4672 -476 4700
rect -448 4672 -410 4700
rect -382 4672 -344 4700
rect -316 4672 -278 4700
rect -250 4672 -212 4700
rect -184 4672 -146 4700
rect -118 4672 -80 4700
rect -52 4672 -14 4700
rect 14 4672 52 4700
rect 80 4672 118 4700
rect 146 4672 184 4700
rect 212 4672 250 4700
rect 278 4672 316 4700
rect 344 4672 382 4700
rect 410 4672 448 4700
rect 476 4672 514 4700
rect 542 4672 580 4700
rect 608 4672 646 4700
rect 674 4672 712 4700
rect 740 4672 745 4700
rect -745 4634 745 4672
rect -745 4606 -740 4634
rect -712 4606 -674 4634
rect -646 4606 -608 4634
rect -580 4606 -542 4634
rect -514 4606 -476 4634
rect -448 4606 -410 4634
rect -382 4606 -344 4634
rect -316 4606 -278 4634
rect -250 4606 -212 4634
rect -184 4606 -146 4634
rect -118 4606 -80 4634
rect -52 4606 -14 4634
rect 14 4606 52 4634
rect 80 4606 118 4634
rect 146 4606 184 4634
rect 212 4606 250 4634
rect 278 4606 316 4634
rect 344 4606 382 4634
rect 410 4606 448 4634
rect 476 4606 514 4634
rect 542 4606 580 4634
rect 608 4606 646 4634
rect 674 4606 712 4634
rect 740 4606 745 4634
rect -745 4568 745 4606
rect -745 4540 -740 4568
rect -712 4540 -674 4568
rect -646 4540 -608 4568
rect -580 4540 -542 4568
rect -514 4540 -476 4568
rect -448 4540 -410 4568
rect -382 4540 -344 4568
rect -316 4540 -278 4568
rect -250 4540 -212 4568
rect -184 4540 -146 4568
rect -118 4540 -80 4568
rect -52 4540 -14 4568
rect 14 4540 52 4568
rect 80 4540 118 4568
rect 146 4540 184 4568
rect 212 4540 250 4568
rect 278 4540 316 4568
rect 344 4540 382 4568
rect 410 4540 448 4568
rect 476 4540 514 4568
rect 542 4540 580 4568
rect 608 4540 646 4568
rect 674 4540 712 4568
rect 740 4540 745 4568
rect -745 4502 745 4540
rect -745 4474 -740 4502
rect -712 4474 -674 4502
rect -646 4474 -608 4502
rect -580 4474 -542 4502
rect -514 4474 -476 4502
rect -448 4474 -410 4502
rect -382 4474 -344 4502
rect -316 4474 -278 4502
rect -250 4474 -212 4502
rect -184 4474 -146 4502
rect -118 4474 -80 4502
rect -52 4474 -14 4502
rect 14 4474 52 4502
rect 80 4474 118 4502
rect 146 4474 184 4502
rect 212 4474 250 4502
rect 278 4474 316 4502
rect 344 4474 382 4502
rect 410 4474 448 4502
rect 476 4474 514 4502
rect 542 4474 580 4502
rect 608 4474 646 4502
rect 674 4474 712 4502
rect 740 4474 745 4502
rect -745 4436 745 4474
rect -745 4408 -740 4436
rect -712 4408 -674 4436
rect -646 4408 -608 4436
rect -580 4408 -542 4436
rect -514 4408 -476 4436
rect -448 4408 -410 4436
rect -382 4408 -344 4436
rect -316 4408 -278 4436
rect -250 4408 -212 4436
rect -184 4408 -146 4436
rect -118 4408 -80 4436
rect -52 4408 -14 4436
rect 14 4408 52 4436
rect 80 4408 118 4436
rect 146 4408 184 4436
rect 212 4408 250 4436
rect 278 4408 316 4436
rect 344 4408 382 4436
rect 410 4408 448 4436
rect 476 4408 514 4436
rect 542 4408 580 4436
rect 608 4408 646 4436
rect 674 4408 712 4436
rect 740 4408 745 4436
rect -745 4370 745 4408
rect -745 4342 -740 4370
rect -712 4342 -674 4370
rect -646 4342 -608 4370
rect -580 4342 -542 4370
rect -514 4342 -476 4370
rect -448 4342 -410 4370
rect -382 4342 -344 4370
rect -316 4342 -278 4370
rect -250 4342 -212 4370
rect -184 4342 -146 4370
rect -118 4342 -80 4370
rect -52 4342 -14 4370
rect 14 4342 52 4370
rect 80 4342 118 4370
rect 146 4342 184 4370
rect 212 4342 250 4370
rect 278 4342 316 4370
rect 344 4342 382 4370
rect 410 4342 448 4370
rect 476 4342 514 4370
rect 542 4342 580 4370
rect 608 4342 646 4370
rect 674 4342 712 4370
rect 740 4342 745 4370
rect -745 4304 745 4342
rect -745 4276 -740 4304
rect -712 4276 -674 4304
rect -646 4276 -608 4304
rect -580 4276 -542 4304
rect -514 4276 -476 4304
rect -448 4276 -410 4304
rect -382 4276 -344 4304
rect -316 4276 -278 4304
rect -250 4276 -212 4304
rect -184 4276 -146 4304
rect -118 4276 -80 4304
rect -52 4276 -14 4304
rect 14 4276 52 4304
rect 80 4276 118 4304
rect 146 4276 184 4304
rect 212 4276 250 4304
rect 278 4276 316 4304
rect 344 4276 382 4304
rect 410 4276 448 4304
rect 476 4276 514 4304
rect 542 4276 580 4304
rect 608 4276 646 4304
rect 674 4276 712 4304
rect 740 4276 745 4304
rect -745 4238 745 4276
rect -745 4210 -740 4238
rect -712 4210 -674 4238
rect -646 4210 -608 4238
rect -580 4210 -542 4238
rect -514 4210 -476 4238
rect -448 4210 -410 4238
rect -382 4210 -344 4238
rect -316 4210 -278 4238
rect -250 4210 -212 4238
rect -184 4210 -146 4238
rect -118 4210 -80 4238
rect -52 4210 -14 4238
rect 14 4210 52 4238
rect 80 4210 118 4238
rect 146 4210 184 4238
rect 212 4210 250 4238
rect 278 4210 316 4238
rect 344 4210 382 4238
rect 410 4210 448 4238
rect 476 4210 514 4238
rect 542 4210 580 4238
rect 608 4210 646 4238
rect 674 4210 712 4238
rect 740 4210 745 4238
rect -745 4172 745 4210
rect -745 4144 -740 4172
rect -712 4144 -674 4172
rect -646 4144 -608 4172
rect -580 4144 -542 4172
rect -514 4144 -476 4172
rect -448 4144 -410 4172
rect -382 4144 -344 4172
rect -316 4144 -278 4172
rect -250 4144 -212 4172
rect -184 4144 -146 4172
rect -118 4144 -80 4172
rect -52 4144 -14 4172
rect 14 4144 52 4172
rect 80 4144 118 4172
rect 146 4144 184 4172
rect 212 4144 250 4172
rect 278 4144 316 4172
rect 344 4144 382 4172
rect 410 4144 448 4172
rect 476 4144 514 4172
rect 542 4144 580 4172
rect 608 4144 646 4172
rect 674 4144 712 4172
rect 740 4144 745 4172
rect -745 4106 745 4144
rect -745 4078 -740 4106
rect -712 4078 -674 4106
rect -646 4078 -608 4106
rect -580 4078 -542 4106
rect -514 4078 -476 4106
rect -448 4078 -410 4106
rect -382 4078 -344 4106
rect -316 4078 -278 4106
rect -250 4078 -212 4106
rect -184 4078 -146 4106
rect -118 4078 -80 4106
rect -52 4078 -14 4106
rect 14 4078 52 4106
rect 80 4078 118 4106
rect 146 4078 184 4106
rect 212 4078 250 4106
rect 278 4078 316 4106
rect 344 4078 382 4106
rect 410 4078 448 4106
rect 476 4078 514 4106
rect 542 4078 580 4106
rect 608 4078 646 4106
rect 674 4078 712 4106
rect 740 4078 745 4106
rect -745 4040 745 4078
rect -745 4012 -740 4040
rect -712 4012 -674 4040
rect -646 4012 -608 4040
rect -580 4012 -542 4040
rect -514 4012 -476 4040
rect -448 4012 -410 4040
rect -382 4012 -344 4040
rect -316 4012 -278 4040
rect -250 4012 -212 4040
rect -184 4012 -146 4040
rect -118 4012 -80 4040
rect -52 4012 -14 4040
rect 14 4012 52 4040
rect 80 4012 118 4040
rect 146 4012 184 4040
rect 212 4012 250 4040
rect 278 4012 316 4040
rect 344 4012 382 4040
rect 410 4012 448 4040
rect 476 4012 514 4040
rect 542 4012 580 4040
rect 608 4012 646 4040
rect 674 4012 712 4040
rect 740 4012 745 4040
rect -745 3974 745 4012
rect -745 3946 -740 3974
rect -712 3946 -674 3974
rect -646 3946 -608 3974
rect -580 3946 -542 3974
rect -514 3946 -476 3974
rect -448 3946 -410 3974
rect -382 3946 -344 3974
rect -316 3946 -278 3974
rect -250 3946 -212 3974
rect -184 3946 -146 3974
rect -118 3946 -80 3974
rect -52 3946 -14 3974
rect 14 3946 52 3974
rect 80 3946 118 3974
rect 146 3946 184 3974
rect 212 3946 250 3974
rect 278 3946 316 3974
rect 344 3946 382 3974
rect 410 3946 448 3974
rect 476 3946 514 3974
rect 542 3946 580 3974
rect 608 3946 646 3974
rect 674 3946 712 3974
rect 740 3946 745 3974
rect -745 3908 745 3946
rect -745 3880 -740 3908
rect -712 3880 -674 3908
rect -646 3880 -608 3908
rect -580 3880 -542 3908
rect -514 3880 -476 3908
rect -448 3880 -410 3908
rect -382 3880 -344 3908
rect -316 3880 -278 3908
rect -250 3880 -212 3908
rect -184 3880 -146 3908
rect -118 3880 -80 3908
rect -52 3880 -14 3908
rect 14 3880 52 3908
rect 80 3880 118 3908
rect 146 3880 184 3908
rect 212 3880 250 3908
rect 278 3880 316 3908
rect 344 3880 382 3908
rect 410 3880 448 3908
rect 476 3880 514 3908
rect 542 3880 580 3908
rect 608 3880 646 3908
rect 674 3880 712 3908
rect 740 3880 745 3908
rect -745 3842 745 3880
rect -745 3814 -740 3842
rect -712 3814 -674 3842
rect -646 3814 -608 3842
rect -580 3814 -542 3842
rect -514 3814 -476 3842
rect -448 3814 -410 3842
rect -382 3814 -344 3842
rect -316 3814 -278 3842
rect -250 3814 -212 3842
rect -184 3814 -146 3842
rect -118 3814 -80 3842
rect -52 3814 -14 3842
rect 14 3814 52 3842
rect 80 3814 118 3842
rect 146 3814 184 3842
rect 212 3814 250 3842
rect 278 3814 316 3842
rect 344 3814 382 3842
rect 410 3814 448 3842
rect 476 3814 514 3842
rect 542 3814 580 3842
rect 608 3814 646 3842
rect 674 3814 712 3842
rect 740 3814 745 3842
rect -745 3776 745 3814
rect -745 3748 -740 3776
rect -712 3748 -674 3776
rect -646 3748 -608 3776
rect -580 3748 -542 3776
rect -514 3748 -476 3776
rect -448 3748 -410 3776
rect -382 3748 -344 3776
rect -316 3748 -278 3776
rect -250 3748 -212 3776
rect -184 3748 -146 3776
rect -118 3748 -80 3776
rect -52 3748 -14 3776
rect 14 3748 52 3776
rect 80 3748 118 3776
rect 146 3748 184 3776
rect 212 3748 250 3776
rect 278 3748 316 3776
rect 344 3748 382 3776
rect 410 3748 448 3776
rect 476 3748 514 3776
rect 542 3748 580 3776
rect 608 3748 646 3776
rect 674 3748 712 3776
rect 740 3748 745 3776
rect -745 3710 745 3748
rect -745 3682 -740 3710
rect -712 3682 -674 3710
rect -646 3682 -608 3710
rect -580 3682 -542 3710
rect -514 3682 -476 3710
rect -448 3682 -410 3710
rect -382 3682 -344 3710
rect -316 3682 -278 3710
rect -250 3682 -212 3710
rect -184 3682 -146 3710
rect -118 3682 -80 3710
rect -52 3682 -14 3710
rect 14 3682 52 3710
rect 80 3682 118 3710
rect 146 3682 184 3710
rect 212 3682 250 3710
rect 278 3682 316 3710
rect 344 3682 382 3710
rect 410 3682 448 3710
rect 476 3682 514 3710
rect 542 3682 580 3710
rect 608 3682 646 3710
rect 674 3682 712 3710
rect 740 3682 745 3710
rect -745 3644 745 3682
rect -745 3616 -740 3644
rect -712 3616 -674 3644
rect -646 3616 -608 3644
rect -580 3616 -542 3644
rect -514 3616 -476 3644
rect -448 3616 -410 3644
rect -382 3616 -344 3644
rect -316 3616 -278 3644
rect -250 3616 -212 3644
rect -184 3616 -146 3644
rect -118 3616 -80 3644
rect -52 3616 -14 3644
rect 14 3616 52 3644
rect 80 3616 118 3644
rect 146 3616 184 3644
rect 212 3616 250 3644
rect 278 3616 316 3644
rect 344 3616 382 3644
rect 410 3616 448 3644
rect 476 3616 514 3644
rect 542 3616 580 3644
rect 608 3616 646 3644
rect 674 3616 712 3644
rect 740 3616 745 3644
rect -745 3578 745 3616
rect -745 3550 -740 3578
rect -712 3550 -674 3578
rect -646 3550 -608 3578
rect -580 3550 -542 3578
rect -514 3550 -476 3578
rect -448 3550 -410 3578
rect -382 3550 -344 3578
rect -316 3550 -278 3578
rect -250 3550 -212 3578
rect -184 3550 -146 3578
rect -118 3550 -80 3578
rect -52 3550 -14 3578
rect 14 3550 52 3578
rect 80 3550 118 3578
rect 146 3550 184 3578
rect 212 3550 250 3578
rect 278 3550 316 3578
rect 344 3550 382 3578
rect 410 3550 448 3578
rect 476 3550 514 3578
rect 542 3550 580 3578
rect 608 3550 646 3578
rect 674 3550 712 3578
rect 740 3550 745 3578
rect -745 3512 745 3550
rect -745 3484 -740 3512
rect -712 3484 -674 3512
rect -646 3484 -608 3512
rect -580 3484 -542 3512
rect -514 3484 -476 3512
rect -448 3484 -410 3512
rect -382 3484 -344 3512
rect -316 3484 -278 3512
rect -250 3484 -212 3512
rect -184 3484 -146 3512
rect -118 3484 -80 3512
rect -52 3484 -14 3512
rect 14 3484 52 3512
rect 80 3484 118 3512
rect 146 3484 184 3512
rect 212 3484 250 3512
rect 278 3484 316 3512
rect 344 3484 382 3512
rect 410 3484 448 3512
rect 476 3484 514 3512
rect 542 3484 580 3512
rect 608 3484 646 3512
rect 674 3484 712 3512
rect 740 3484 745 3512
rect -745 3446 745 3484
rect -745 3418 -740 3446
rect -712 3418 -674 3446
rect -646 3418 -608 3446
rect -580 3418 -542 3446
rect -514 3418 -476 3446
rect -448 3418 -410 3446
rect -382 3418 -344 3446
rect -316 3418 -278 3446
rect -250 3418 -212 3446
rect -184 3418 -146 3446
rect -118 3418 -80 3446
rect -52 3418 -14 3446
rect 14 3418 52 3446
rect 80 3418 118 3446
rect 146 3418 184 3446
rect 212 3418 250 3446
rect 278 3418 316 3446
rect 344 3418 382 3446
rect 410 3418 448 3446
rect 476 3418 514 3446
rect 542 3418 580 3446
rect 608 3418 646 3446
rect 674 3418 712 3446
rect 740 3418 745 3446
rect -745 3380 745 3418
rect -745 3352 -740 3380
rect -712 3352 -674 3380
rect -646 3352 -608 3380
rect -580 3352 -542 3380
rect -514 3352 -476 3380
rect -448 3352 -410 3380
rect -382 3352 -344 3380
rect -316 3352 -278 3380
rect -250 3352 -212 3380
rect -184 3352 -146 3380
rect -118 3352 -80 3380
rect -52 3352 -14 3380
rect 14 3352 52 3380
rect 80 3352 118 3380
rect 146 3352 184 3380
rect 212 3352 250 3380
rect 278 3352 316 3380
rect 344 3352 382 3380
rect 410 3352 448 3380
rect 476 3352 514 3380
rect 542 3352 580 3380
rect 608 3352 646 3380
rect 674 3352 712 3380
rect 740 3352 745 3380
rect -745 3314 745 3352
rect -745 3286 -740 3314
rect -712 3286 -674 3314
rect -646 3286 -608 3314
rect -580 3286 -542 3314
rect -514 3286 -476 3314
rect -448 3286 -410 3314
rect -382 3286 -344 3314
rect -316 3286 -278 3314
rect -250 3286 -212 3314
rect -184 3286 -146 3314
rect -118 3286 -80 3314
rect -52 3286 -14 3314
rect 14 3286 52 3314
rect 80 3286 118 3314
rect 146 3286 184 3314
rect 212 3286 250 3314
rect 278 3286 316 3314
rect 344 3286 382 3314
rect 410 3286 448 3314
rect 476 3286 514 3314
rect 542 3286 580 3314
rect 608 3286 646 3314
rect 674 3286 712 3314
rect 740 3286 745 3314
rect -745 3248 745 3286
rect -745 3220 -740 3248
rect -712 3220 -674 3248
rect -646 3220 -608 3248
rect -580 3220 -542 3248
rect -514 3220 -476 3248
rect -448 3220 -410 3248
rect -382 3220 -344 3248
rect -316 3220 -278 3248
rect -250 3220 -212 3248
rect -184 3220 -146 3248
rect -118 3220 -80 3248
rect -52 3220 -14 3248
rect 14 3220 52 3248
rect 80 3220 118 3248
rect 146 3220 184 3248
rect 212 3220 250 3248
rect 278 3220 316 3248
rect 344 3220 382 3248
rect 410 3220 448 3248
rect 476 3220 514 3248
rect 542 3220 580 3248
rect 608 3220 646 3248
rect 674 3220 712 3248
rect 740 3220 745 3248
rect -745 3182 745 3220
rect -745 3154 -740 3182
rect -712 3154 -674 3182
rect -646 3154 -608 3182
rect -580 3154 -542 3182
rect -514 3154 -476 3182
rect -448 3154 -410 3182
rect -382 3154 -344 3182
rect -316 3154 -278 3182
rect -250 3154 -212 3182
rect -184 3154 -146 3182
rect -118 3154 -80 3182
rect -52 3154 -14 3182
rect 14 3154 52 3182
rect 80 3154 118 3182
rect 146 3154 184 3182
rect 212 3154 250 3182
rect 278 3154 316 3182
rect 344 3154 382 3182
rect 410 3154 448 3182
rect 476 3154 514 3182
rect 542 3154 580 3182
rect 608 3154 646 3182
rect 674 3154 712 3182
rect 740 3154 745 3182
rect -745 3116 745 3154
rect -745 3088 -740 3116
rect -712 3088 -674 3116
rect -646 3088 -608 3116
rect -580 3088 -542 3116
rect -514 3088 -476 3116
rect -448 3088 -410 3116
rect -382 3088 -344 3116
rect -316 3088 -278 3116
rect -250 3088 -212 3116
rect -184 3088 -146 3116
rect -118 3088 -80 3116
rect -52 3088 -14 3116
rect 14 3088 52 3116
rect 80 3088 118 3116
rect 146 3088 184 3116
rect 212 3088 250 3116
rect 278 3088 316 3116
rect 344 3088 382 3116
rect 410 3088 448 3116
rect 476 3088 514 3116
rect 542 3088 580 3116
rect 608 3088 646 3116
rect 674 3088 712 3116
rect 740 3088 745 3116
rect -745 3050 745 3088
rect -745 3022 -740 3050
rect -712 3022 -674 3050
rect -646 3022 -608 3050
rect -580 3022 -542 3050
rect -514 3022 -476 3050
rect -448 3022 -410 3050
rect -382 3022 -344 3050
rect -316 3022 -278 3050
rect -250 3022 -212 3050
rect -184 3022 -146 3050
rect -118 3022 -80 3050
rect -52 3022 -14 3050
rect 14 3022 52 3050
rect 80 3022 118 3050
rect 146 3022 184 3050
rect 212 3022 250 3050
rect 278 3022 316 3050
rect 344 3022 382 3050
rect 410 3022 448 3050
rect 476 3022 514 3050
rect 542 3022 580 3050
rect 608 3022 646 3050
rect 674 3022 712 3050
rect 740 3022 745 3050
rect -745 2984 745 3022
rect -745 2956 -740 2984
rect -712 2956 -674 2984
rect -646 2956 -608 2984
rect -580 2956 -542 2984
rect -514 2956 -476 2984
rect -448 2956 -410 2984
rect -382 2956 -344 2984
rect -316 2956 -278 2984
rect -250 2956 -212 2984
rect -184 2956 -146 2984
rect -118 2956 -80 2984
rect -52 2956 -14 2984
rect 14 2956 52 2984
rect 80 2956 118 2984
rect 146 2956 184 2984
rect 212 2956 250 2984
rect 278 2956 316 2984
rect 344 2956 382 2984
rect 410 2956 448 2984
rect 476 2956 514 2984
rect 542 2956 580 2984
rect 608 2956 646 2984
rect 674 2956 712 2984
rect 740 2956 745 2984
rect -745 2918 745 2956
rect -745 2890 -740 2918
rect -712 2890 -674 2918
rect -646 2890 -608 2918
rect -580 2890 -542 2918
rect -514 2890 -476 2918
rect -448 2890 -410 2918
rect -382 2890 -344 2918
rect -316 2890 -278 2918
rect -250 2890 -212 2918
rect -184 2890 -146 2918
rect -118 2890 -80 2918
rect -52 2890 -14 2918
rect 14 2890 52 2918
rect 80 2890 118 2918
rect 146 2890 184 2918
rect 212 2890 250 2918
rect 278 2890 316 2918
rect 344 2890 382 2918
rect 410 2890 448 2918
rect 476 2890 514 2918
rect 542 2890 580 2918
rect 608 2890 646 2918
rect 674 2890 712 2918
rect 740 2890 745 2918
rect -745 2852 745 2890
rect -745 2824 -740 2852
rect -712 2824 -674 2852
rect -646 2824 -608 2852
rect -580 2824 -542 2852
rect -514 2824 -476 2852
rect -448 2824 -410 2852
rect -382 2824 -344 2852
rect -316 2824 -278 2852
rect -250 2824 -212 2852
rect -184 2824 -146 2852
rect -118 2824 -80 2852
rect -52 2824 -14 2852
rect 14 2824 52 2852
rect 80 2824 118 2852
rect 146 2824 184 2852
rect 212 2824 250 2852
rect 278 2824 316 2852
rect 344 2824 382 2852
rect 410 2824 448 2852
rect 476 2824 514 2852
rect 542 2824 580 2852
rect 608 2824 646 2852
rect 674 2824 712 2852
rect 740 2824 745 2852
rect -745 2786 745 2824
rect -745 2758 -740 2786
rect -712 2758 -674 2786
rect -646 2758 -608 2786
rect -580 2758 -542 2786
rect -514 2758 -476 2786
rect -448 2758 -410 2786
rect -382 2758 -344 2786
rect -316 2758 -278 2786
rect -250 2758 -212 2786
rect -184 2758 -146 2786
rect -118 2758 -80 2786
rect -52 2758 -14 2786
rect 14 2758 52 2786
rect 80 2758 118 2786
rect 146 2758 184 2786
rect 212 2758 250 2786
rect 278 2758 316 2786
rect 344 2758 382 2786
rect 410 2758 448 2786
rect 476 2758 514 2786
rect 542 2758 580 2786
rect 608 2758 646 2786
rect 674 2758 712 2786
rect 740 2758 745 2786
rect -745 2720 745 2758
rect -745 2692 -740 2720
rect -712 2692 -674 2720
rect -646 2692 -608 2720
rect -580 2692 -542 2720
rect -514 2692 -476 2720
rect -448 2692 -410 2720
rect -382 2692 -344 2720
rect -316 2692 -278 2720
rect -250 2692 -212 2720
rect -184 2692 -146 2720
rect -118 2692 -80 2720
rect -52 2692 -14 2720
rect 14 2692 52 2720
rect 80 2692 118 2720
rect 146 2692 184 2720
rect 212 2692 250 2720
rect 278 2692 316 2720
rect 344 2692 382 2720
rect 410 2692 448 2720
rect 476 2692 514 2720
rect 542 2692 580 2720
rect 608 2692 646 2720
rect 674 2692 712 2720
rect 740 2692 745 2720
rect -745 2654 745 2692
rect -745 2626 -740 2654
rect -712 2626 -674 2654
rect -646 2626 -608 2654
rect -580 2626 -542 2654
rect -514 2626 -476 2654
rect -448 2626 -410 2654
rect -382 2626 -344 2654
rect -316 2626 -278 2654
rect -250 2626 -212 2654
rect -184 2626 -146 2654
rect -118 2626 -80 2654
rect -52 2626 -14 2654
rect 14 2626 52 2654
rect 80 2626 118 2654
rect 146 2626 184 2654
rect 212 2626 250 2654
rect 278 2626 316 2654
rect 344 2626 382 2654
rect 410 2626 448 2654
rect 476 2626 514 2654
rect 542 2626 580 2654
rect 608 2626 646 2654
rect 674 2626 712 2654
rect 740 2626 745 2654
rect -745 2588 745 2626
rect -745 2560 -740 2588
rect -712 2560 -674 2588
rect -646 2560 -608 2588
rect -580 2560 -542 2588
rect -514 2560 -476 2588
rect -448 2560 -410 2588
rect -382 2560 -344 2588
rect -316 2560 -278 2588
rect -250 2560 -212 2588
rect -184 2560 -146 2588
rect -118 2560 -80 2588
rect -52 2560 -14 2588
rect 14 2560 52 2588
rect 80 2560 118 2588
rect 146 2560 184 2588
rect 212 2560 250 2588
rect 278 2560 316 2588
rect 344 2560 382 2588
rect 410 2560 448 2588
rect 476 2560 514 2588
rect 542 2560 580 2588
rect 608 2560 646 2588
rect 674 2560 712 2588
rect 740 2560 745 2588
rect -745 2522 745 2560
rect -745 2494 -740 2522
rect -712 2494 -674 2522
rect -646 2494 -608 2522
rect -580 2494 -542 2522
rect -514 2494 -476 2522
rect -448 2494 -410 2522
rect -382 2494 -344 2522
rect -316 2494 -278 2522
rect -250 2494 -212 2522
rect -184 2494 -146 2522
rect -118 2494 -80 2522
rect -52 2494 -14 2522
rect 14 2494 52 2522
rect 80 2494 118 2522
rect 146 2494 184 2522
rect 212 2494 250 2522
rect 278 2494 316 2522
rect 344 2494 382 2522
rect 410 2494 448 2522
rect 476 2494 514 2522
rect 542 2494 580 2522
rect 608 2494 646 2522
rect 674 2494 712 2522
rect 740 2494 745 2522
rect -745 2456 745 2494
rect -745 2428 -740 2456
rect -712 2428 -674 2456
rect -646 2428 -608 2456
rect -580 2428 -542 2456
rect -514 2428 -476 2456
rect -448 2428 -410 2456
rect -382 2428 -344 2456
rect -316 2428 -278 2456
rect -250 2428 -212 2456
rect -184 2428 -146 2456
rect -118 2428 -80 2456
rect -52 2428 -14 2456
rect 14 2428 52 2456
rect 80 2428 118 2456
rect 146 2428 184 2456
rect 212 2428 250 2456
rect 278 2428 316 2456
rect 344 2428 382 2456
rect 410 2428 448 2456
rect 476 2428 514 2456
rect 542 2428 580 2456
rect 608 2428 646 2456
rect 674 2428 712 2456
rect 740 2428 745 2456
rect -745 2390 745 2428
rect -745 2362 -740 2390
rect -712 2362 -674 2390
rect -646 2362 -608 2390
rect -580 2362 -542 2390
rect -514 2362 -476 2390
rect -448 2362 -410 2390
rect -382 2362 -344 2390
rect -316 2362 -278 2390
rect -250 2362 -212 2390
rect -184 2362 -146 2390
rect -118 2362 -80 2390
rect -52 2362 -14 2390
rect 14 2362 52 2390
rect 80 2362 118 2390
rect 146 2362 184 2390
rect 212 2362 250 2390
rect 278 2362 316 2390
rect 344 2362 382 2390
rect 410 2362 448 2390
rect 476 2362 514 2390
rect 542 2362 580 2390
rect 608 2362 646 2390
rect 674 2362 712 2390
rect 740 2362 745 2390
rect -745 2324 745 2362
rect -745 2296 -740 2324
rect -712 2296 -674 2324
rect -646 2296 -608 2324
rect -580 2296 -542 2324
rect -514 2296 -476 2324
rect -448 2296 -410 2324
rect -382 2296 -344 2324
rect -316 2296 -278 2324
rect -250 2296 -212 2324
rect -184 2296 -146 2324
rect -118 2296 -80 2324
rect -52 2296 -14 2324
rect 14 2296 52 2324
rect 80 2296 118 2324
rect 146 2296 184 2324
rect 212 2296 250 2324
rect 278 2296 316 2324
rect 344 2296 382 2324
rect 410 2296 448 2324
rect 476 2296 514 2324
rect 542 2296 580 2324
rect 608 2296 646 2324
rect 674 2296 712 2324
rect 740 2296 745 2324
rect -745 2258 745 2296
rect -745 2230 -740 2258
rect -712 2230 -674 2258
rect -646 2230 -608 2258
rect -580 2230 -542 2258
rect -514 2230 -476 2258
rect -448 2230 -410 2258
rect -382 2230 -344 2258
rect -316 2230 -278 2258
rect -250 2230 -212 2258
rect -184 2230 -146 2258
rect -118 2230 -80 2258
rect -52 2230 -14 2258
rect 14 2230 52 2258
rect 80 2230 118 2258
rect 146 2230 184 2258
rect 212 2230 250 2258
rect 278 2230 316 2258
rect 344 2230 382 2258
rect 410 2230 448 2258
rect 476 2230 514 2258
rect 542 2230 580 2258
rect 608 2230 646 2258
rect 674 2230 712 2258
rect 740 2230 745 2258
rect -745 2192 745 2230
rect -745 2164 -740 2192
rect -712 2164 -674 2192
rect -646 2164 -608 2192
rect -580 2164 -542 2192
rect -514 2164 -476 2192
rect -448 2164 -410 2192
rect -382 2164 -344 2192
rect -316 2164 -278 2192
rect -250 2164 -212 2192
rect -184 2164 -146 2192
rect -118 2164 -80 2192
rect -52 2164 -14 2192
rect 14 2164 52 2192
rect 80 2164 118 2192
rect 146 2164 184 2192
rect 212 2164 250 2192
rect 278 2164 316 2192
rect 344 2164 382 2192
rect 410 2164 448 2192
rect 476 2164 514 2192
rect 542 2164 580 2192
rect 608 2164 646 2192
rect 674 2164 712 2192
rect 740 2164 745 2192
rect -745 2126 745 2164
rect -745 2098 -740 2126
rect -712 2098 -674 2126
rect -646 2098 -608 2126
rect -580 2098 -542 2126
rect -514 2098 -476 2126
rect -448 2098 -410 2126
rect -382 2098 -344 2126
rect -316 2098 -278 2126
rect -250 2098 -212 2126
rect -184 2098 -146 2126
rect -118 2098 -80 2126
rect -52 2098 -14 2126
rect 14 2098 52 2126
rect 80 2098 118 2126
rect 146 2098 184 2126
rect 212 2098 250 2126
rect 278 2098 316 2126
rect 344 2098 382 2126
rect 410 2098 448 2126
rect 476 2098 514 2126
rect 542 2098 580 2126
rect 608 2098 646 2126
rect 674 2098 712 2126
rect 740 2098 745 2126
rect -745 2060 745 2098
rect -745 2032 -740 2060
rect -712 2032 -674 2060
rect -646 2032 -608 2060
rect -580 2032 -542 2060
rect -514 2032 -476 2060
rect -448 2032 -410 2060
rect -382 2032 -344 2060
rect -316 2032 -278 2060
rect -250 2032 -212 2060
rect -184 2032 -146 2060
rect -118 2032 -80 2060
rect -52 2032 -14 2060
rect 14 2032 52 2060
rect 80 2032 118 2060
rect 146 2032 184 2060
rect 212 2032 250 2060
rect 278 2032 316 2060
rect 344 2032 382 2060
rect 410 2032 448 2060
rect 476 2032 514 2060
rect 542 2032 580 2060
rect 608 2032 646 2060
rect 674 2032 712 2060
rect 740 2032 745 2060
rect -745 1994 745 2032
rect -745 1966 -740 1994
rect -712 1966 -674 1994
rect -646 1966 -608 1994
rect -580 1966 -542 1994
rect -514 1966 -476 1994
rect -448 1966 -410 1994
rect -382 1966 -344 1994
rect -316 1966 -278 1994
rect -250 1966 -212 1994
rect -184 1966 -146 1994
rect -118 1966 -80 1994
rect -52 1966 -14 1994
rect 14 1966 52 1994
rect 80 1966 118 1994
rect 146 1966 184 1994
rect 212 1966 250 1994
rect 278 1966 316 1994
rect 344 1966 382 1994
rect 410 1966 448 1994
rect 476 1966 514 1994
rect 542 1966 580 1994
rect 608 1966 646 1994
rect 674 1966 712 1994
rect 740 1966 745 1994
rect -745 1928 745 1966
rect -745 1900 -740 1928
rect -712 1900 -674 1928
rect -646 1900 -608 1928
rect -580 1900 -542 1928
rect -514 1900 -476 1928
rect -448 1900 -410 1928
rect -382 1900 -344 1928
rect -316 1900 -278 1928
rect -250 1900 -212 1928
rect -184 1900 -146 1928
rect -118 1900 -80 1928
rect -52 1900 -14 1928
rect 14 1900 52 1928
rect 80 1900 118 1928
rect 146 1900 184 1928
rect 212 1900 250 1928
rect 278 1900 316 1928
rect 344 1900 382 1928
rect 410 1900 448 1928
rect 476 1900 514 1928
rect 542 1900 580 1928
rect 608 1900 646 1928
rect 674 1900 712 1928
rect 740 1900 745 1928
rect -745 1862 745 1900
rect -745 1834 -740 1862
rect -712 1834 -674 1862
rect -646 1834 -608 1862
rect -580 1834 -542 1862
rect -514 1834 -476 1862
rect -448 1834 -410 1862
rect -382 1834 -344 1862
rect -316 1834 -278 1862
rect -250 1834 -212 1862
rect -184 1834 -146 1862
rect -118 1834 -80 1862
rect -52 1834 -14 1862
rect 14 1834 52 1862
rect 80 1834 118 1862
rect 146 1834 184 1862
rect 212 1834 250 1862
rect 278 1834 316 1862
rect 344 1834 382 1862
rect 410 1834 448 1862
rect 476 1834 514 1862
rect 542 1834 580 1862
rect 608 1834 646 1862
rect 674 1834 712 1862
rect 740 1834 745 1862
rect -745 1796 745 1834
rect -745 1768 -740 1796
rect -712 1768 -674 1796
rect -646 1768 -608 1796
rect -580 1768 -542 1796
rect -514 1768 -476 1796
rect -448 1768 -410 1796
rect -382 1768 -344 1796
rect -316 1768 -278 1796
rect -250 1768 -212 1796
rect -184 1768 -146 1796
rect -118 1768 -80 1796
rect -52 1768 -14 1796
rect 14 1768 52 1796
rect 80 1768 118 1796
rect 146 1768 184 1796
rect 212 1768 250 1796
rect 278 1768 316 1796
rect 344 1768 382 1796
rect 410 1768 448 1796
rect 476 1768 514 1796
rect 542 1768 580 1796
rect 608 1768 646 1796
rect 674 1768 712 1796
rect 740 1768 745 1796
rect -745 1730 745 1768
rect -745 1702 -740 1730
rect -712 1702 -674 1730
rect -646 1702 -608 1730
rect -580 1702 -542 1730
rect -514 1702 -476 1730
rect -448 1702 -410 1730
rect -382 1702 -344 1730
rect -316 1702 -278 1730
rect -250 1702 -212 1730
rect -184 1702 -146 1730
rect -118 1702 -80 1730
rect -52 1702 -14 1730
rect 14 1702 52 1730
rect 80 1702 118 1730
rect 146 1702 184 1730
rect 212 1702 250 1730
rect 278 1702 316 1730
rect 344 1702 382 1730
rect 410 1702 448 1730
rect 476 1702 514 1730
rect 542 1702 580 1730
rect 608 1702 646 1730
rect 674 1702 712 1730
rect 740 1702 745 1730
rect -745 1664 745 1702
rect -745 1636 -740 1664
rect -712 1636 -674 1664
rect -646 1636 -608 1664
rect -580 1636 -542 1664
rect -514 1636 -476 1664
rect -448 1636 -410 1664
rect -382 1636 -344 1664
rect -316 1636 -278 1664
rect -250 1636 -212 1664
rect -184 1636 -146 1664
rect -118 1636 -80 1664
rect -52 1636 -14 1664
rect 14 1636 52 1664
rect 80 1636 118 1664
rect 146 1636 184 1664
rect 212 1636 250 1664
rect 278 1636 316 1664
rect 344 1636 382 1664
rect 410 1636 448 1664
rect 476 1636 514 1664
rect 542 1636 580 1664
rect 608 1636 646 1664
rect 674 1636 712 1664
rect 740 1636 745 1664
rect -745 1598 745 1636
rect -745 1570 -740 1598
rect -712 1570 -674 1598
rect -646 1570 -608 1598
rect -580 1570 -542 1598
rect -514 1570 -476 1598
rect -448 1570 -410 1598
rect -382 1570 -344 1598
rect -316 1570 -278 1598
rect -250 1570 -212 1598
rect -184 1570 -146 1598
rect -118 1570 -80 1598
rect -52 1570 -14 1598
rect 14 1570 52 1598
rect 80 1570 118 1598
rect 146 1570 184 1598
rect 212 1570 250 1598
rect 278 1570 316 1598
rect 344 1570 382 1598
rect 410 1570 448 1598
rect 476 1570 514 1598
rect 542 1570 580 1598
rect 608 1570 646 1598
rect 674 1570 712 1598
rect 740 1570 745 1598
rect -745 1532 745 1570
rect -745 1504 -740 1532
rect -712 1504 -674 1532
rect -646 1504 -608 1532
rect -580 1504 -542 1532
rect -514 1504 -476 1532
rect -448 1504 -410 1532
rect -382 1504 -344 1532
rect -316 1504 -278 1532
rect -250 1504 -212 1532
rect -184 1504 -146 1532
rect -118 1504 -80 1532
rect -52 1504 -14 1532
rect 14 1504 52 1532
rect 80 1504 118 1532
rect 146 1504 184 1532
rect 212 1504 250 1532
rect 278 1504 316 1532
rect 344 1504 382 1532
rect 410 1504 448 1532
rect 476 1504 514 1532
rect 542 1504 580 1532
rect 608 1504 646 1532
rect 674 1504 712 1532
rect 740 1504 745 1532
rect -745 1466 745 1504
rect -745 1438 -740 1466
rect -712 1438 -674 1466
rect -646 1438 -608 1466
rect -580 1438 -542 1466
rect -514 1438 -476 1466
rect -448 1438 -410 1466
rect -382 1438 -344 1466
rect -316 1438 -278 1466
rect -250 1438 -212 1466
rect -184 1438 -146 1466
rect -118 1438 -80 1466
rect -52 1438 -14 1466
rect 14 1438 52 1466
rect 80 1438 118 1466
rect 146 1438 184 1466
rect 212 1438 250 1466
rect 278 1438 316 1466
rect 344 1438 382 1466
rect 410 1438 448 1466
rect 476 1438 514 1466
rect 542 1438 580 1466
rect 608 1438 646 1466
rect 674 1438 712 1466
rect 740 1438 745 1466
rect -745 1400 745 1438
rect -745 1372 -740 1400
rect -712 1372 -674 1400
rect -646 1372 -608 1400
rect -580 1372 -542 1400
rect -514 1372 -476 1400
rect -448 1372 -410 1400
rect -382 1372 -344 1400
rect -316 1372 -278 1400
rect -250 1372 -212 1400
rect -184 1372 -146 1400
rect -118 1372 -80 1400
rect -52 1372 -14 1400
rect 14 1372 52 1400
rect 80 1372 118 1400
rect 146 1372 184 1400
rect 212 1372 250 1400
rect 278 1372 316 1400
rect 344 1372 382 1400
rect 410 1372 448 1400
rect 476 1372 514 1400
rect 542 1372 580 1400
rect 608 1372 646 1400
rect 674 1372 712 1400
rect 740 1372 745 1400
rect -745 1334 745 1372
rect -745 1306 -740 1334
rect -712 1306 -674 1334
rect -646 1306 -608 1334
rect -580 1306 -542 1334
rect -514 1306 -476 1334
rect -448 1306 -410 1334
rect -382 1306 -344 1334
rect -316 1306 -278 1334
rect -250 1306 -212 1334
rect -184 1306 -146 1334
rect -118 1306 -80 1334
rect -52 1306 -14 1334
rect 14 1306 52 1334
rect 80 1306 118 1334
rect 146 1306 184 1334
rect 212 1306 250 1334
rect 278 1306 316 1334
rect 344 1306 382 1334
rect 410 1306 448 1334
rect 476 1306 514 1334
rect 542 1306 580 1334
rect 608 1306 646 1334
rect 674 1306 712 1334
rect 740 1306 745 1334
rect -745 1268 745 1306
rect -745 1240 -740 1268
rect -712 1240 -674 1268
rect -646 1240 -608 1268
rect -580 1240 -542 1268
rect -514 1240 -476 1268
rect -448 1240 -410 1268
rect -382 1240 -344 1268
rect -316 1240 -278 1268
rect -250 1240 -212 1268
rect -184 1240 -146 1268
rect -118 1240 -80 1268
rect -52 1240 -14 1268
rect 14 1240 52 1268
rect 80 1240 118 1268
rect 146 1240 184 1268
rect 212 1240 250 1268
rect 278 1240 316 1268
rect 344 1240 382 1268
rect 410 1240 448 1268
rect 476 1240 514 1268
rect 542 1240 580 1268
rect 608 1240 646 1268
rect 674 1240 712 1268
rect 740 1240 745 1268
rect -745 1202 745 1240
rect -745 1174 -740 1202
rect -712 1174 -674 1202
rect -646 1174 -608 1202
rect -580 1174 -542 1202
rect -514 1174 -476 1202
rect -448 1174 -410 1202
rect -382 1174 -344 1202
rect -316 1174 -278 1202
rect -250 1174 -212 1202
rect -184 1174 -146 1202
rect -118 1174 -80 1202
rect -52 1174 -14 1202
rect 14 1174 52 1202
rect 80 1174 118 1202
rect 146 1174 184 1202
rect 212 1174 250 1202
rect 278 1174 316 1202
rect 344 1174 382 1202
rect 410 1174 448 1202
rect 476 1174 514 1202
rect 542 1174 580 1202
rect 608 1174 646 1202
rect 674 1174 712 1202
rect 740 1174 745 1202
rect -745 1136 745 1174
rect -745 1108 -740 1136
rect -712 1108 -674 1136
rect -646 1108 -608 1136
rect -580 1108 -542 1136
rect -514 1108 -476 1136
rect -448 1108 -410 1136
rect -382 1108 -344 1136
rect -316 1108 -278 1136
rect -250 1108 -212 1136
rect -184 1108 -146 1136
rect -118 1108 -80 1136
rect -52 1108 -14 1136
rect 14 1108 52 1136
rect 80 1108 118 1136
rect 146 1108 184 1136
rect 212 1108 250 1136
rect 278 1108 316 1136
rect 344 1108 382 1136
rect 410 1108 448 1136
rect 476 1108 514 1136
rect 542 1108 580 1136
rect 608 1108 646 1136
rect 674 1108 712 1136
rect 740 1108 745 1136
rect -745 1070 745 1108
rect -745 1042 -740 1070
rect -712 1042 -674 1070
rect -646 1042 -608 1070
rect -580 1042 -542 1070
rect -514 1042 -476 1070
rect -448 1042 -410 1070
rect -382 1042 -344 1070
rect -316 1042 -278 1070
rect -250 1042 -212 1070
rect -184 1042 -146 1070
rect -118 1042 -80 1070
rect -52 1042 -14 1070
rect 14 1042 52 1070
rect 80 1042 118 1070
rect 146 1042 184 1070
rect 212 1042 250 1070
rect 278 1042 316 1070
rect 344 1042 382 1070
rect 410 1042 448 1070
rect 476 1042 514 1070
rect 542 1042 580 1070
rect 608 1042 646 1070
rect 674 1042 712 1070
rect 740 1042 745 1070
rect -745 1004 745 1042
rect -745 976 -740 1004
rect -712 976 -674 1004
rect -646 976 -608 1004
rect -580 976 -542 1004
rect -514 976 -476 1004
rect -448 976 -410 1004
rect -382 976 -344 1004
rect -316 976 -278 1004
rect -250 976 -212 1004
rect -184 976 -146 1004
rect -118 976 -80 1004
rect -52 976 -14 1004
rect 14 976 52 1004
rect 80 976 118 1004
rect 146 976 184 1004
rect 212 976 250 1004
rect 278 976 316 1004
rect 344 976 382 1004
rect 410 976 448 1004
rect 476 976 514 1004
rect 542 976 580 1004
rect 608 976 646 1004
rect 674 976 712 1004
rect 740 976 745 1004
rect -745 938 745 976
rect -745 910 -740 938
rect -712 910 -674 938
rect -646 910 -608 938
rect -580 910 -542 938
rect -514 910 -476 938
rect -448 910 -410 938
rect -382 910 -344 938
rect -316 910 -278 938
rect -250 910 -212 938
rect -184 910 -146 938
rect -118 910 -80 938
rect -52 910 -14 938
rect 14 910 52 938
rect 80 910 118 938
rect 146 910 184 938
rect 212 910 250 938
rect 278 910 316 938
rect 344 910 382 938
rect 410 910 448 938
rect 476 910 514 938
rect 542 910 580 938
rect 608 910 646 938
rect 674 910 712 938
rect 740 910 745 938
rect -745 872 745 910
rect -745 844 -740 872
rect -712 844 -674 872
rect -646 844 -608 872
rect -580 844 -542 872
rect -514 844 -476 872
rect -448 844 -410 872
rect -382 844 -344 872
rect -316 844 -278 872
rect -250 844 -212 872
rect -184 844 -146 872
rect -118 844 -80 872
rect -52 844 -14 872
rect 14 844 52 872
rect 80 844 118 872
rect 146 844 184 872
rect 212 844 250 872
rect 278 844 316 872
rect 344 844 382 872
rect 410 844 448 872
rect 476 844 514 872
rect 542 844 580 872
rect 608 844 646 872
rect 674 844 712 872
rect 740 844 745 872
rect -745 806 745 844
rect -745 778 -740 806
rect -712 778 -674 806
rect -646 778 -608 806
rect -580 778 -542 806
rect -514 778 -476 806
rect -448 778 -410 806
rect -382 778 -344 806
rect -316 778 -278 806
rect -250 778 -212 806
rect -184 778 -146 806
rect -118 778 -80 806
rect -52 778 -14 806
rect 14 778 52 806
rect 80 778 118 806
rect 146 778 184 806
rect 212 778 250 806
rect 278 778 316 806
rect 344 778 382 806
rect 410 778 448 806
rect 476 778 514 806
rect 542 778 580 806
rect 608 778 646 806
rect 674 778 712 806
rect 740 778 745 806
rect -745 740 745 778
rect -745 712 -740 740
rect -712 712 -674 740
rect -646 712 -608 740
rect -580 712 -542 740
rect -514 712 -476 740
rect -448 712 -410 740
rect -382 712 -344 740
rect -316 712 -278 740
rect -250 712 -212 740
rect -184 712 -146 740
rect -118 712 -80 740
rect -52 712 -14 740
rect 14 712 52 740
rect 80 712 118 740
rect 146 712 184 740
rect 212 712 250 740
rect 278 712 316 740
rect 344 712 382 740
rect 410 712 448 740
rect 476 712 514 740
rect 542 712 580 740
rect 608 712 646 740
rect 674 712 712 740
rect 740 712 745 740
rect -745 674 745 712
rect -745 646 -740 674
rect -712 646 -674 674
rect -646 646 -608 674
rect -580 646 -542 674
rect -514 646 -476 674
rect -448 646 -410 674
rect -382 646 -344 674
rect -316 646 -278 674
rect -250 646 -212 674
rect -184 646 -146 674
rect -118 646 -80 674
rect -52 646 -14 674
rect 14 646 52 674
rect 80 646 118 674
rect 146 646 184 674
rect 212 646 250 674
rect 278 646 316 674
rect 344 646 382 674
rect 410 646 448 674
rect 476 646 514 674
rect 542 646 580 674
rect 608 646 646 674
rect 674 646 712 674
rect 740 646 745 674
rect -745 608 745 646
rect -745 580 -740 608
rect -712 580 -674 608
rect -646 580 -608 608
rect -580 580 -542 608
rect -514 580 -476 608
rect -448 580 -410 608
rect -382 580 -344 608
rect -316 580 -278 608
rect -250 580 -212 608
rect -184 580 -146 608
rect -118 580 -80 608
rect -52 580 -14 608
rect 14 580 52 608
rect 80 580 118 608
rect 146 580 184 608
rect 212 580 250 608
rect 278 580 316 608
rect 344 580 382 608
rect 410 580 448 608
rect 476 580 514 608
rect 542 580 580 608
rect 608 580 646 608
rect 674 580 712 608
rect 740 580 745 608
rect -745 542 745 580
rect -745 514 -740 542
rect -712 514 -674 542
rect -646 514 -608 542
rect -580 514 -542 542
rect -514 514 -476 542
rect -448 514 -410 542
rect -382 514 -344 542
rect -316 514 -278 542
rect -250 514 -212 542
rect -184 514 -146 542
rect -118 514 -80 542
rect -52 514 -14 542
rect 14 514 52 542
rect 80 514 118 542
rect 146 514 184 542
rect 212 514 250 542
rect 278 514 316 542
rect 344 514 382 542
rect 410 514 448 542
rect 476 514 514 542
rect 542 514 580 542
rect 608 514 646 542
rect 674 514 712 542
rect 740 514 745 542
rect -745 476 745 514
rect -745 448 -740 476
rect -712 448 -674 476
rect -646 448 -608 476
rect -580 448 -542 476
rect -514 448 -476 476
rect -448 448 -410 476
rect -382 448 -344 476
rect -316 448 -278 476
rect -250 448 -212 476
rect -184 448 -146 476
rect -118 448 -80 476
rect -52 448 -14 476
rect 14 448 52 476
rect 80 448 118 476
rect 146 448 184 476
rect 212 448 250 476
rect 278 448 316 476
rect 344 448 382 476
rect 410 448 448 476
rect 476 448 514 476
rect 542 448 580 476
rect 608 448 646 476
rect 674 448 712 476
rect 740 448 745 476
rect -745 410 745 448
rect -745 382 -740 410
rect -712 382 -674 410
rect -646 382 -608 410
rect -580 382 -542 410
rect -514 382 -476 410
rect -448 382 -410 410
rect -382 382 -344 410
rect -316 382 -278 410
rect -250 382 -212 410
rect -184 382 -146 410
rect -118 382 -80 410
rect -52 382 -14 410
rect 14 382 52 410
rect 80 382 118 410
rect 146 382 184 410
rect 212 382 250 410
rect 278 382 316 410
rect 344 382 382 410
rect 410 382 448 410
rect 476 382 514 410
rect 542 382 580 410
rect 608 382 646 410
rect 674 382 712 410
rect 740 382 745 410
rect -745 344 745 382
rect -745 316 -740 344
rect -712 316 -674 344
rect -646 316 -608 344
rect -580 316 -542 344
rect -514 316 -476 344
rect -448 316 -410 344
rect -382 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 382 344
rect 410 316 448 344
rect 476 316 514 344
rect 542 316 580 344
rect 608 316 646 344
rect 674 316 712 344
rect 740 316 745 344
rect -745 278 745 316
rect -745 250 -740 278
rect -712 250 -674 278
rect -646 250 -608 278
rect -580 250 -542 278
rect -514 250 -476 278
rect -448 250 -410 278
rect -382 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 382 278
rect 410 250 448 278
rect 476 250 514 278
rect 542 250 580 278
rect 608 250 646 278
rect 674 250 712 278
rect 740 250 745 278
rect -745 212 745 250
rect -745 184 -740 212
rect -712 184 -674 212
rect -646 184 -608 212
rect -580 184 -542 212
rect -514 184 -476 212
rect -448 184 -410 212
rect -382 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 382 212
rect 410 184 448 212
rect 476 184 514 212
rect 542 184 580 212
rect 608 184 646 212
rect 674 184 712 212
rect 740 184 745 212
rect -745 146 745 184
rect -745 118 -740 146
rect -712 118 -674 146
rect -646 118 -608 146
rect -580 118 -542 146
rect -514 118 -476 146
rect -448 118 -410 146
rect -382 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 382 146
rect 410 118 448 146
rect 476 118 514 146
rect 542 118 580 146
rect 608 118 646 146
rect 674 118 712 146
rect 740 118 745 146
rect -745 80 745 118
rect -745 52 -740 80
rect -712 52 -674 80
rect -646 52 -608 80
rect -580 52 -542 80
rect -514 52 -476 80
rect -448 52 -410 80
rect -382 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 382 80
rect 410 52 448 80
rect 476 52 514 80
rect 542 52 580 80
rect 608 52 646 80
rect 674 52 712 80
rect 740 52 745 80
rect -745 14 745 52
rect -745 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 382 14
rect 410 -14 448 14
rect 476 -14 514 14
rect 542 -14 580 14
rect 608 -14 646 14
rect 674 -14 712 14
rect 740 -14 745 14
rect -745 -52 745 -14
rect -745 -80 -740 -52
rect -712 -80 -674 -52
rect -646 -80 -608 -52
rect -580 -80 -542 -52
rect -514 -80 -476 -52
rect -448 -80 -410 -52
rect -382 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 382 -52
rect 410 -80 448 -52
rect 476 -80 514 -52
rect 542 -80 580 -52
rect 608 -80 646 -52
rect 674 -80 712 -52
rect 740 -80 745 -52
rect -745 -118 745 -80
rect -745 -146 -740 -118
rect -712 -146 -674 -118
rect -646 -146 -608 -118
rect -580 -146 -542 -118
rect -514 -146 -476 -118
rect -448 -146 -410 -118
rect -382 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 382 -118
rect 410 -146 448 -118
rect 476 -146 514 -118
rect 542 -146 580 -118
rect 608 -146 646 -118
rect 674 -146 712 -118
rect 740 -146 745 -118
rect -745 -184 745 -146
rect -745 -212 -740 -184
rect -712 -212 -674 -184
rect -646 -212 -608 -184
rect -580 -212 -542 -184
rect -514 -212 -476 -184
rect -448 -212 -410 -184
rect -382 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 382 -184
rect 410 -212 448 -184
rect 476 -212 514 -184
rect 542 -212 580 -184
rect 608 -212 646 -184
rect 674 -212 712 -184
rect 740 -212 745 -184
rect -745 -250 745 -212
rect -745 -278 -740 -250
rect -712 -278 -674 -250
rect -646 -278 -608 -250
rect -580 -278 -542 -250
rect -514 -278 -476 -250
rect -448 -278 -410 -250
rect -382 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 382 -250
rect 410 -278 448 -250
rect 476 -278 514 -250
rect 542 -278 580 -250
rect 608 -278 646 -250
rect 674 -278 712 -250
rect 740 -278 745 -250
rect -745 -316 745 -278
rect -745 -344 -740 -316
rect -712 -344 -674 -316
rect -646 -344 -608 -316
rect -580 -344 -542 -316
rect -514 -344 -476 -316
rect -448 -344 -410 -316
rect -382 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 382 -316
rect 410 -344 448 -316
rect 476 -344 514 -316
rect 542 -344 580 -316
rect 608 -344 646 -316
rect 674 -344 712 -316
rect 740 -344 745 -316
rect -745 -382 745 -344
rect -745 -410 -740 -382
rect -712 -410 -674 -382
rect -646 -410 -608 -382
rect -580 -410 -542 -382
rect -514 -410 -476 -382
rect -448 -410 -410 -382
rect -382 -410 -344 -382
rect -316 -410 -278 -382
rect -250 -410 -212 -382
rect -184 -410 -146 -382
rect -118 -410 -80 -382
rect -52 -410 -14 -382
rect 14 -410 52 -382
rect 80 -410 118 -382
rect 146 -410 184 -382
rect 212 -410 250 -382
rect 278 -410 316 -382
rect 344 -410 382 -382
rect 410 -410 448 -382
rect 476 -410 514 -382
rect 542 -410 580 -382
rect 608 -410 646 -382
rect 674 -410 712 -382
rect 740 -410 745 -382
rect -745 -448 745 -410
rect -745 -476 -740 -448
rect -712 -476 -674 -448
rect -646 -476 -608 -448
rect -580 -476 -542 -448
rect -514 -476 -476 -448
rect -448 -476 -410 -448
rect -382 -476 -344 -448
rect -316 -476 -278 -448
rect -250 -476 -212 -448
rect -184 -476 -146 -448
rect -118 -476 -80 -448
rect -52 -476 -14 -448
rect 14 -476 52 -448
rect 80 -476 118 -448
rect 146 -476 184 -448
rect 212 -476 250 -448
rect 278 -476 316 -448
rect 344 -476 382 -448
rect 410 -476 448 -448
rect 476 -476 514 -448
rect 542 -476 580 -448
rect 608 -476 646 -448
rect 674 -476 712 -448
rect 740 -476 745 -448
rect -745 -514 745 -476
rect -745 -542 -740 -514
rect -712 -542 -674 -514
rect -646 -542 -608 -514
rect -580 -542 -542 -514
rect -514 -542 -476 -514
rect -448 -542 -410 -514
rect -382 -542 -344 -514
rect -316 -542 -278 -514
rect -250 -542 -212 -514
rect -184 -542 -146 -514
rect -118 -542 -80 -514
rect -52 -542 -14 -514
rect 14 -542 52 -514
rect 80 -542 118 -514
rect 146 -542 184 -514
rect 212 -542 250 -514
rect 278 -542 316 -514
rect 344 -542 382 -514
rect 410 -542 448 -514
rect 476 -542 514 -514
rect 542 -542 580 -514
rect 608 -542 646 -514
rect 674 -542 712 -514
rect 740 -542 745 -514
rect -745 -580 745 -542
rect -745 -608 -740 -580
rect -712 -608 -674 -580
rect -646 -608 -608 -580
rect -580 -608 -542 -580
rect -514 -608 -476 -580
rect -448 -608 -410 -580
rect -382 -608 -344 -580
rect -316 -608 -278 -580
rect -250 -608 -212 -580
rect -184 -608 -146 -580
rect -118 -608 -80 -580
rect -52 -608 -14 -580
rect 14 -608 52 -580
rect 80 -608 118 -580
rect 146 -608 184 -580
rect 212 -608 250 -580
rect 278 -608 316 -580
rect 344 -608 382 -580
rect 410 -608 448 -580
rect 476 -608 514 -580
rect 542 -608 580 -580
rect 608 -608 646 -580
rect 674 -608 712 -580
rect 740 -608 745 -580
rect -745 -646 745 -608
rect -745 -674 -740 -646
rect -712 -674 -674 -646
rect -646 -674 -608 -646
rect -580 -674 -542 -646
rect -514 -674 -476 -646
rect -448 -674 -410 -646
rect -382 -674 -344 -646
rect -316 -674 -278 -646
rect -250 -674 -212 -646
rect -184 -674 -146 -646
rect -118 -674 -80 -646
rect -52 -674 -14 -646
rect 14 -674 52 -646
rect 80 -674 118 -646
rect 146 -674 184 -646
rect 212 -674 250 -646
rect 278 -674 316 -646
rect 344 -674 382 -646
rect 410 -674 448 -646
rect 476 -674 514 -646
rect 542 -674 580 -646
rect 608 -674 646 -646
rect 674 -674 712 -646
rect 740 -674 745 -646
rect -745 -712 745 -674
rect -745 -740 -740 -712
rect -712 -740 -674 -712
rect -646 -740 -608 -712
rect -580 -740 -542 -712
rect -514 -740 -476 -712
rect -448 -740 -410 -712
rect -382 -740 -344 -712
rect -316 -740 -278 -712
rect -250 -740 -212 -712
rect -184 -740 -146 -712
rect -118 -740 -80 -712
rect -52 -740 -14 -712
rect 14 -740 52 -712
rect 80 -740 118 -712
rect 146 -740 184 -712
rect 212 -740 250 -712
rect 278 -740 316 -712
rect 344 -740 382 -712
rect 410 -740 448 -712
rect 476 -740 514 -712
rect 542 -740 580 -712
rect 608 -740 646 -712
rect 674 -740 712 -712
rect 740 -740 745 -712
rect -745 -778 745 -740
rect -745 -806 -740 -778
rect -712 -806 -674 -778
rect -646 -806 -608 -778
rect -580 -806 -542 -778
rect -514 -806 -476 -778
rect -448 -806 -410 -778
rect -382 -806 -344 -778
rect -316 -806 -278 -778
rect -250 -806 -212 -778
rect -184 -806 -146 -778
rect -118 -806 -80 -778
rect -52 -806 -14 -778
rect 14 -806 52 -778
rect 80 -806 118 -778
rect 146 -806 184 -778
rect 212 -806 250 -778
rect 278 -806 316 -778
rect 344 -806 382 -778
rect 410 -806 448 -778
rect 476 -806 514 -778
rect 542 -806 580 -778
rect 608 -806 646 -778
rect 674 -806 712 -778
rect 740 -806 745 -778
rect -745 -844 745 -806
rect -745 -872 -740 -844
rect -712 -872 -674 -844
rect -646 -872 -608 -844
rect -580 -872 -542 -844
rect -514 -872 -476 -844
rect -448 -872 -410 -844
rect -382 -872 -344 -844
rect -316 -872 -278 -844
rect -250 -872 -212 -844
rect -184 -872 -146 -844
rect -118 -872 -80 -844
rect -52 -872 -14 -844
rect 14 -872 52 -844
rect 80 -872 118 -844
rect 146 -872 184 -844
rect 212 -872 250 -844
rect 278 -872 316 -844
rect 344 -872 382 -844
rect 410 -872 448 -844
rect 476 -872 514 -844
rect 542 -872 580 -844
rect 608 -872 646 -844
rect 674 -872 712 -844
rect 740 -872 745 -844
rect -745 -910 745 -872
rect -745 -938 -740 -910
rect -712 -938 -674 -910
rect -646 -938 -608 -910
rect -580 -938 -542 -910
rect -514 -938 -476 -910
rect -448 -938 -410 -910
rect -382 -938 -344 -910
rect -316 -938 -278 -910
rect -250 -938 -212 -910
rect -184 -938 -146 -910
rect -118 -938 -80 -910
rect -52 -938 -14 -910
rect 14 -938 52 -910
rect 80 -938 118 -910
rect 146 -938 184 -910
rect 212 -938 250 -910
rect 278 -938 316 -910
rect 344 -938 382 -910
rect 410 -938 448 -910
rect 476 -938 514 -910
rect 542 -938 580 -910
rect 608 -938 646 -910
rect 674 -938 712 -910
rect 740 -938 745 -910
rect -745 -976 745 -938
rect -745 -1004 -740 -976
rect -712 -1004 -674 -976
rect -646 -1004 -608 -976
rect -580 -1004 -542 -976
rect -514 -1004 -476 -976
rect -448 -1004 -410 -976
rect -382 -1004 -344 -976
rect -316 -1004 -278 -976
rect -250 -1004 -212 -976
rect -184 -1004 -146 -976
rect -118 -1004 -80 -976
rect -52 -1004 -14 -976
rect 14 -1004 52 -976
rect 80 -1004 118 -976
rect 146 -1004 184 -976
rect 212 -1004 250 -976
rect 278 -1004 316 -976
rect 344 -1004 382 -976
rect 410 -1004 448 -976
rect 476 -1004 514 -976
rect 542 -1004 580 -976
rect 608 -1004 646 -976
rect 674 -1004 712 -976
rect 740 -1004 745 -976
rect -745 -1042 745 -1004
rect -745 -1070 -740 -1042
rect -712 -1070 -674 -1042
rect -646 -1070 -608 -1042
rect -580 -1070 -542 -1042
rect -514 -1070 -476 -1042
rect -448 -1070 -410 -1042
rect -382 -1070 -344 -1042
rect -316 -1070 -278 -1042
rect -250 -1070 -212 -1042
rect -184 -1070 -146 -1042
rect -118 -1070 -80 -1042
rect -52 -1070 -14 -1042
rect 14 -1070 52 -1042
rect 80 -1070 118 -1042
rect 146 -1070 184 -1042
rect 212 -1070 250 -1042
rect 278 -1070 316 -1042
rect 344 -1070 382 -1042
rect 410 -1070 448 -1042
rect 476 -1070 514 -1042
rect 542 -1070 580 -1042
rect 608 -1070 646 -1042
rect 674 -1070 712 -1042
rect 740 -1070 745 -1042
rect -745 -1108 745 -1070
rect -745 -1136 -740 -1108
rect -712 -1136 -674 -1108
rect -646 -1136 -608 -1108
rect -580 -1136 -542 -1108
rect -514 -1136 -476 -1108
rect -448 -1136 -410 -1108
rect -382 -1136 -344 -1108
rect -316 -1136 -278 -1108
rect -250 -1136 -212 -1108
rect -184 -1136 -146 -1108
rect -118 -1136 -80 -1108
rect -52 -1136 -14 -1108
rect 14 -1136 52 -1108
rect 80 -1136 118 -1108
rect 146 -1136 184 -1108
rect 212 -1136 250 -1108
rect 278 -1136 316 -1108
rect 344 -1136 382 -1108
rect 410 -1136 448 -1108
rect 476 -1136 514 -1108
rect 542 -1136 580 -1108
rect 608 -1136 646 -1108
rect 674 -1136 712 -1108
rect 740 -1136 745 -1108
rect -745 -1174 745 -1136
rect -745 -1202 -740 -1174
rect -712 -1202 -674 -1174
rect -646 -1202 -608 -1174
rect -580 -1202 -542 -1174
rect -514 -1202 -476 -1174
rect -448 -1202 -410 -1174
rect -382 -1202 -344 -1174
rect -316 -1202 -278 -1174
rect -250 -1202 -212 -1174
rect -184 -1202 -146 -1174
rect -118 -1202 -80 -1174
rect -52 -1202 -14 -1174
rect 14 -1202 52 -1174
rect 80 -1202 118 -1174
rect 146 -1202 184 -1174
rect 212 -1202 250 -1174
rect 278 -1202 316 -1174
rect 344 -1202 382 -1174
rect 410 -1202 448 -1174
rect 476 -1202 514 -1174
rect 542 -1202 580 -1174
rect 608 -1202 646 -1174
rect 674 -1202 712 -1174
rect 740 -1202 745 -1174
rect -745 -1240 745 -1202
rect -745 -1268 -740 -1240
rect -712 -1268 -674 -1240
rect -646 -1268 -608 -1240
rect -580 -1268 -542 -1240
rect -514 -1268 -476 -1240
rect -448 -1268 -410 -1240
rect -382 -1268 -344 -1240
rect -316 -1268 -278 -1240
rect -250 -1268 -212 -1240
rect -184 -1268 -146 -1240
rect -118 -1268 -80 -1240
rect -52 -1268 -14 -1240
rect 14 -1268 52 -1240
rect 80 -1268 118 -1240
rect 146 -1268 184 -1240
rect 212 -1268 250 -1240
rect 278 -1268 316 -1240
rect 344 -1268 382 -1240
rect 410 -1268 448 -1240
rect 476 -1268 514 -1240
rect 542 -1268 580 -1240
rect 608 -1268 646 -1240
rect 674 -1268 712 -1240
rect 740 -1268 745 -1240
rect -745 -1306 745 -1268
rect -745 -1334 -740 -1306
rect -712 -1334 -674 -1306
rect -646 -1334 -608 -1306
rect -580 -1334 -542 -1306
rect -514 -1334 -476 -1306
rect -448 -1334 -410 -1306
rect -382 -1334 -344 -1306
rect -316 -1334 -278 -1306
rect -250 -1334 -212 -1306
rect -184 -1334 -146 -1306
rect -118 -1334 -80 -1306
rect -52 -1334 -14 -1306
rect 14 -1334 52 -1306
rect 80 -1334 118 -1306
rect 146 -1334 184 -1306
rect 212 -1334 250 -1306
rect 278 -1334 316 -1306
rect 344 -1334 382 -1306
rect 410 -1334 448 -1306
rect 476 -1334 514 -1306
rect 542 -1334 580 -1306
rect 608 -1334 646 -1306
rect 674 -1334 712 -1306
rect 740 -1334 745 -1306
rect -745 -1372 745 -1334
rect -745 -1400 -740 -1372
rect -712 -1400 -674 -1372
rect -646 -1400 -608 -1372
rect -580 -1400 -542 -1372
rect -514 -1400 -476 -1372
rect -448 -1400 -410 -1372
rect -382 -1400 -344 -1372
rect -316 -1400 -278 -1372
rect -250 -1400 -212 -1372
rect -184 -1400 -146 -1372
rect -118 -1400 -80 -1372
rect -52 -1400 -14 -1372
rect 14 -1400 52 -1372
rect 80 -1400 118 -1372
rect 146 -1400 184 -1372
rect 212 -1400 250 -1372
rect 278 -1400 316 -1372
rect 344 -1400 382 -1372
rect 410 -1400 448 -1372
rect 476 -1400 514 -1372
rect 542 -1400 580 -1372
rect 608 -1400 646 -1372
rect 674 -1400 712 -1372
rect 740 -1400 745 -1372
rect -745 -1438 745 -1400
rect -745 -1466 -740 -1438
rect -712 -1466 -674 -1438
rect -646 -1466 -608 -1438
rect -580 -1466 -542 -1438
rect -514 -1466 -476 -1438
rect -448 -1466 -410 -1438
rect -382 -1466 -344 -1438
rect -316 -1466 -278 -1438
rect -250 -1466 -212 -1438
rect -184 -1466 -146 -1438
rect -118 -1466 -80 -1438
rect -52 -1466 -14 -1438
rect 14 -1466 52 -1438
rect 80 -1466 118 -1438
rect 146 -1466 184 -1438
rect 212 -1466 250 -1438
rect 278 -1466 316 -1438
rect 344 -1466 382 -1438
rect 410 -1466 448 -1438
rect 476 -1466 514 -1438
rect 542 -1466 580 -1438
rect 608 -1466 646 -1438
rect 674 -1466 712 -1438
rect 740 -1466 745 -1438
rect -745 -1504 745 -1466
rect -745 -1532 -740 -1504
rect -712 -1532 -674 -1504
rect -646 -1532 -608 -1504
rect -580 -1532 -542 -1504
rect -514 -1532 -476 -1504
rect -448 -1532 -410 -1504
rect -382 -1532 -344 -1504
rect -316 -1532 -278 -1504
rect -250 -1532 -212 -1504
rect -184 -1532 -146 -1504
rect -118 -1532 -80 -1504
rect -52 -1532 -14 -1504
rect 14 -1532 52 -1504
rect 80 -1532 118 -1504
rect 146 -1532 184 -1504
rect 212 -1532 250 -1504
rect 278 -1532 316 -1504
rect 344 -1532 382 -1504
rect 410 -1532 448 -1504
rect 476 -1532 514 -1504
rect 542 -1532 580 -1504
rect 608 -1532 646 -1504
rect 674 -1532 712 -1504
rect 740 -1532 745 -1504
rect -745 -1570 745 -1532
rect -745 -1598 -740 -1570
rect -712 -1598 -674 -1570
rect -646 -1598 -608 -1570
rect -580 -1598 -542 -1570
rect -514 -1598 -476 -1570
rect -448 -1598 -410 -1570
rect -382 -1598 -344 -1570
rect -316 -1598 -278 -1570
rect -250 -1598 -212 -1570
rect -184 -1598 -146 -1570
rect -118 -1598 -80 -1570
rect -52 -1598 -14 -1570
rect 14 -1598 52 -1570
rect 80 -1598 118 -1570
rect 146 -1598 184 -1570
rect 212 -1598 250 -1570
rect 278 -1598 316 -1570
rect 344 -1598 382 -1570
rect 410 -1598 448 -1570
rect 476 -1598 514 -1570
rect 542 -1598 580 -1570
rect 608 -1598 646 -1570
rect 674 -1598 712 -1570
rect 740 -1598 745 -1570
rect -745 -1636 745 -1598
rect -745 -1664 -740 -1636
rect -712 -1664 -674 -1636
rect -646 -1664 -608 -1636
rect -580 -1664 -542 -1636
rect -514 -1664 -476 -1636
rect -448 -1664 -410 -1636
rect -382 -1664 -344 -1636
rect -316 -1664 -278 -1636
rect -250 -1664 -212 -1636
rect -184 -1664 -146 -1636
rect -118 -1664 -80 -1636
rect -52 -1664 -14 -1636
rect 14 -1664 52 -1636
rect 80 -1664 118 -1636
rect 146 -1664 184 -1636
rect 212 -1664 250 -1636
rect 278 -1664 316 -1636
rect 344 -1664 382 -1636
rect 410 -1664 448 -1636
rect 476 -1664 514 -1636
rect 542 -1664 580 -1636
rect 608 -1664 646 -1636
rect 674 -1664 712 -1636
rect 740 -1664 745 -1636
rect -745 -1702 745 -1664
rect -745 -1730 -740 -1702
rect -712 -1730 -674 -1702
rect -646 -1730 -608 -1702
rect -580 -1730 -542 -1702
rect -514 -1730 -476 -1702
rect -448 -1730 -410 -1702
rect -382 -1730 -344 -1702
rect -316 -1730 -278 -1702
rect -250 -1730 -212 -1702
rect -184 -1730 -146 -1702
rect -118 -1730 -80 -1702
rect -52 -1730 -14 -1702
rect 14 -1730 52 -1702
rect 80 -1730 118 -1702
rect 146 -1730 184 -1702
rect 212 -1730 250 -1702
rect 278 -1730 316 -1702
rect 344 -1730 382 -1702
rect 410 -1730 448 -1702
rect 476 -1730 514 -1702
rect 542 -1730 580 -1702
rect 608 -1730 646 -1702
rect 674 -1730 712 -1702
rect 740 -1730 745 -1702
rect -745 -1768 745 -1730
rect -745 -1796 -740 -1768
rect -712 -1796 -674 -1768
rect -646 -1796 -608 -1768
rect -580 -1796 -542 -1768
rect -514 -1796 -476 -1768
rect -448 -1796 -410 -1768
rect -382 -1796 -344 -1768
rect -316 -1796 -278 -1768
rect -250 -1796 -212 -1768
rect -184 -1796 -146 -1768
rect -118 -1796 -80 -1768
rect -52 -1796 -14 -1768
rect 14 -1796 52 -1768
rect 80 -1796 118 -1768
rect 146 -1796 184 -1768
rect 212 -1796 250 -1768
rect 278 -1796 316 -1768
rect 344 -1796 382 -1768
rect 410 -1796 448 -1768
rect 476 -1796 514 -1768
rect 542 -1796 580 -1768
rect 608 -1796 646 -1768
rect 674 -1796 712 -1768
rect 740 -1796 745 -1768
rect -745 -1834 745 -1796
rect -745 -1862 -740 -1834
rect -712 -1862 -674 -1834
rect -646 -1862 -608 -1834
rect -580 -1862 -542 -1834
rect -514 -1862 -476 -1834
rect -448 -1862 -410 -1834
rect -382 -1862 -344 -1834
rect -316 -1862 -278 -1834
rect -250 -1862 -212 -1834
rect -184 -1862 -146 -1834
rect -118 -1862 -80 -1834
rect -52 -1862 -14 -1834
rect 14 -1862 52 -1834
rect 80 -1862 118 -1834
rect 146 -1862 184 -1834
rect 212 -1862 250 -1834
rect 278 -1862 316 -1834
rect 344 -1862 382 -1834
rect 410 -1862 448 -1834
rect 476 -1862 514 -1834
rect 542 -1862 580 -1834
rect 608 -1862 646 -1834
rect 674 -1862 712 -1834
rect 740 -1862 745 -1834
rect -745 -1900 745 -1862
rect -745 -1928 -740 -1900
rect -712 -1928 -674 -1900
rect -646 -1928 -608 -1900
rect -580 -1928 -542 -1900
rect -514 -1928 -476 -1900
rect -448 -1928 -410 -1900
rect -382 -1928 -344 -1900
rect -316 -1928 -278 -1900
rect -250 -1928 -212 -1900
rect -184 -1928 -146 -1900
rect -118 -1928 -80 -1900
rect -52 -1928 -14 -1900
rect 14 -1928 52 -1900
rect 80 -1928 118 -1900
rect 146 -1928 184 -1900
rect 212 -1928 250 -1900
rect 278 -1928 316 -1900
rect 344 -1928 382 -1900
rect 410 -1928 448 -1900
rect 476 -1928 514 -1900
rect 542 -1928 580 -1900
rect 608 -1928 646 -1900
rect 674 -1928 712 -1900
rect 740 -1928 745 -1900
rect -745 -1966 745 -1928
rect -745 -1994 -740 -1966
rect -712 -1994 -674 -1966
rect -646 -1994 -608 -1966
rect -580 -1994 -542 -1966
rect -514 -1994 -476 -1966
rect -448 -1994 -410 -1966
rect -382 -1994 -344 -1966
rect -316 -1994 -278 -1966
rect -250 -1994 -212 -1966
rect -184 -1994 -146 -1966
rect -118 -1994 -80 -1966
rect -52 -1994 -14 -1966
rect 14 -1994 52 -1966
rect 80 -1994 118 -1966
rect 146 -1994 184 -1966
rect 212 -1994 250 -1966
rect 278 -1994 316 -1966
rect 344 -1994 382 -1966
rect 410 -1994 448 -1966
rect 476 -1994 514 -1966
rect 542 -1994 580 -1966
rect 608 -1994 646 -1966
rect 674 -1994 712 -1966
rect 740 -1994 745 -1966
rect -745 -2032 745 -1994
rect -745 -2060 -740 -2032
rect -712 -2060 -674 -2032
rect -646 -2060 -608 -2032
rect -580 -2060 -542 -2032
rect -514 -2060 -476 -2032
rect -448 -2060 -410 -2032
rect -382 -2060 -344 -2032
rect -316 -2060 -278 -2032
rect -250 -2060 -212 -2032
rect -184 -2060 -146 -2032
rect -118 -2060 -80 -2032
rect -52 -2060 -14 -2032
rect 14 -2060 52 -2032
rect 80 -2060 118 -2032
rect 146 -2060 184 -2032
rect 212 -2060 250 -2032
rect 278 -2060 316 -2032
rect 344 -2060 382 -2032
rect 410 -2060 448 -2032
rect 476 -2060 514 -2032
rect 542 -2060 580 -2032
rect 608 -2060 646 -2032
rect 674 -2060 712 -2032
rect 740 -2060 745 -2032
rect -745 -2098 745 -2060
rect -745 -2126 -740 -2098
rect -712 -2126 -674 -2098
rect -646 -2126 -608 -2098
rect -580 -2126 -542 -2098
rect -514 -2126 -476 -2098
rect -448 -2126 -410 -2098
rect -382 -2126 -344 -2098
rect -316 -2126 -278 -2098
rect -250 -2126 -212 -2098
rect -184 -2126 -146 -2098
rect -118 -2126 -80 -2098
rect -52 -2126 -14 -2098
rect 14 -2126 52 -2098
rect 80 -2126 118 -2098
rect 146 -2126 184 -2098
rect 212 -2126 250 -2098
rect 278 -2126 316 -2098
rect 344 -2126 382 -2098
rect 410 -2126 448 -2098
rect 476 -2126 514 -2098
rect 542 -2126 580 -2098
rect 608 -2126 646 -2098
rect 674 -2126 712 -2098
rect 740 -2126 745 -2098
rect -745 -2164 745 -2126
rect -745 -2192 -740 -2164
rect -712 -2192 -674 -2164
rect -646 -2192 -608 -2164
rect -580 -2192 -542 -2164
rect -514 -2192 -476 -2164
rect -448 -2192 -410 -2164
rect -382 -2192 -344 -2164
rect -316 -2192 -278 -2164
rect -250 -2192 -212 -2164
rect -184 -2192 -146 -2164
rect -118 -2192 -80 -2164
rect -52 -2192 -14 -2164
rect 14 -2192 52 -2164
rect 80 -2192 118 -2164
rect 146 -2192 184 -2164
rect 212 -2192 250 -2164
rect 278 -2192 316 -2164
rect 344 -2192 382 -2164
rect 410 -2192 448 -2164
rect 476 -2192 514 -2164
rect 542 -2192 580 -2164
rect 608 -2192 646 -2164
rect 674 -2192 712 -2164
rect 740 -2192 745 -2164
rect -745 -2230 745 -2192
rect -745 -2258 -740 -2230
rect -712 -2258 -674 -2230
rect -646 -2258 -608 -2230
rect -580 -2258 -542 -2230
rect -514 -2258 -476 -2230
rect -448 -2258 -410 -2230
rect -382 -2258 -344 -2230
rect -316 -2258 -278 -2230
rect -250 -2258 -212 -2230
rect -184 -2258 -146 -2230
rect -118 -2258 -80 -2230
rect -52 -2258 -14 -2230
rect 14 -2258 52 -2230
rect 80 -2258 118 -2230
rect 146 -2258 184 -2230
rect 212 -2258 250 -2230
rect 278 -2258 316 -2230
rect 344 -2258 382 -2230
rect 410 -2258 448 -2230
rect 476 -2258 514 -2230
rect 542 -2258 580 -2230
rect 608 -2258 646 -2230
rect 674 -2258 712 -2230
rect 740 -2258 745 -2230
rect -745 -2296 745 -2258
rect -745 -2324 -740 -2296
rect -712 -2324 -674 -2296
rect -646 -2324 -608 -2296
rect -580 -2324 -542 -2296
rect -514 -2324 -476 -2296
rect -448 -2324 -410 -2296
rect -382 -2324 -344 -2296
rect -316 -2324 -278 -2296
rect -250 -2324 -212 -2296
rect -184 -2324 -146 -2296
rect -118 -2324 -80 -2296
rect -52 -2324 -14 -2296
rect 14 -2324 52 -2296
rect 80 -2324 118 -2296
rect 146 -2324 184 -2296
rect 212 -2324 250 -2296
rect 278 -2324 316 -2296
rect 344 -2324 382 -2296
rect 410 -2324 448 -2296
rect 476 -2324 514 -2296
rect 542 -2324 580 -2296
rect 608 -2324 646 -2296
rect 674 -2324 712 -2296
rect 740 -2324 745 -2296
rect -745 -2362 745 -2324
rect -745 -2390 -740 -2362
rect -712 -2390 -674 -2362
rect -646 -2390 -608 -2362
rect -580 -2390 -542 -2362
rect -514 -2390 -476 -2362
rect -448 -2390 -410 -2362
rect -382 -2390 -344 -2362
rect -316 -2390 -278 -2362
rect -250 -2390 -212 -2362
rect -184 -2390 -146 -2362
rect -118 -2390 -80 -2362
rect -52 -2390 -14 -2362
rect 14 -2390 52 -2362
rect 80 -2390 118 -2362
rect 146 -2390 184 -2362
rect 212 -2390 250 -2362
rect 278 -2390 316 -2362
rect 344 -2390 382 -2362
rect 410 -2390 448 -2362
rect 476 -2390 514 -2362
rect 542 -2390 580 -2362
rect 608 -2390 646 -2362
rect 674 -2390 712 -2362
rect 740 -2390 745 -2362
rect -745 -2428 745 -2390
rect -745 -2456 -740 -2428
rect -712 -2456 -674 -2428
rect -646 -2456 -608 -2428
rect -580 -2456 -542 -2428
rect -514 -2456 -476 -2428
rect -448 -2456 -410 -2428
rect -382 -2456 -344 -2428
rect -316 -2456 -278 -2428
rect -250 -2456 -212 -2428
rect -184 -2456 -146 -2428
rect -118 -2456 -80 -2428
rect -52 -2456 -14 -2428
rect 14 -2456 52 -2428
rect 80 -2456 118 -2428
rect 146 -2456 184 -2428
rect 212 -2456 250 -2428
rect 278 -2456 316 -2428
rect 344 -2456 382 -2428
rect 410 -2456 448 -2428
rect 476 -2456 514 -2428
rect 542 -2456 580 -2428
rect 608 -2456 646 -2428
rect 674 -2456 712 -2428
rect 740 -2456 745 -2428
rect -745 -2494 745 -2456
rect -745 -2522 -740 -2494
rect -712 -2522 -674 -2494
rect -646 -2522 -608 -2494
rect -580 -2522 -542 -2494
rect -514 -2522 -476 -2494
rect -448 -2522 -410 -2494
rect -382 -2522 -344 -2494
rect -316 -2522 -278 -2494
rect -250 -2522 -212 -2494
rect -184 -2522 -146 -2494
rect -118 -2522 -80 -2494
rect -52 -2522 -14 -2494
rect 14 -2522 52 -2494
rect 80 -2522 118 -2494
rect 146 -2522 184 -2494
rect 212 -2522 250 -2494
rect 278 -2522 316 -2494
rect 344 -2522 382 -2494
rect 410 -2522 448 -2494
rect 476 -2522 514 -2494
rect 542 -2522 580 -2494
rect 608 -2522 646 -2494
rect 674 -2522 712 -2494
rect 740 -2522 745 -2494
rect -745 -2560 745 -2522
rect -745 -2588 -740 -2560
rect -712 -2588 -674 -2560
rect -646 -2588 -608 -2560
rect -580 -2588 -542 -2560
rect -514 -2588 -476 -2560
rect -448 -2588 -410 -2560
rect -382 -2588 -344 -2560
rect -316 -2588 -278 -2560
rect -250 -2588 -212 -2560
rect -184 -2588 -146 -2560
rect -118 -2588 -80 -2560
rect -52 -2588 -14 -2560
rect 14 -2588 52 -2560
rect 80 -2588 118 -2560
rect 146 -2588 184 -2560
rect 212 -2588 250 -2560
rect 278 -2588 316 -2560
rect 344 -2588 382 -2560
rect 410 -2588 448 -2560
rect 476 -2588 514 -2560
rect 542 -2588 580 -2560
rect 608 -2588 646 -2560
rect 674 -2588 712 -2560
rect 740 -2588 745 -2560
rect -745 -2626 745 -2588
rect -745 -2654 -740 -2626
rect -712 -2654 -674 -2626
rect -646 -2654 -608 -2626
rect -580 -2654 -542 -2626
rect -514 -2654 -476 -2626
rect -448 -2654 -410 -2626
rect -382 -2654 -344 -2626
rect -316 -2654 -278 -2626
rect -250 -2654 -212 -2626
rect -184 -2654 -146 -2626
rect -118 -2654 -80 -2626
rect -52 -2654 -14 -2626
rect 14 -2654 52 -2626
rect 80 -2654 118 -2626
rect 146 -2654 184 -2626
rect 212 -2654 250 -2626
rect 278 -2654 316 -2626
rect 344 -2654 382 -2626
rect 410 -2654 448 -2626
rect 476 -2654 514 -2626
rect 542 -2654 580 -2626
rect 608 -2654 646 -2626
rect 674 -2654 712 -2626
rect 740 -2654 745 -2626
rect -745 -2692 745 -2654
rect -745 -2720 -740 -2692
rect -712 -2720 -674 -2692
rect -646 -2720 -608 -2692
rect -580 -2720 -542 -2692
rect -514 -2720 -476 -2692
rect -448 -2720 -410 -2692
rect -382 -2720 -344 -2692
rect -316 -2720 -278 -2692
rect -250 -2720 -212 -2692
rect -184 -2720 -146 -2692
rect -118 -2720 -80 -2692
rect -52 -2720 -14 -2692
rect 14 -2720 52 -2692
rect 80 -2720 118 -2692
rect 146 -2720 184 -2692
rect 212 -2720 250 -2692
rect 278 -2720 316 -2692
rect 344 -2720 382 -2692
rect 410 -2720 448 -2692
rect 476 -2720 514 -2692
rect 542 -2720 580 -2692
rect 608 -2720 646 -2692
rect 674 -2720 712 -2692
rect 740 -2720 745 -2692
rect -745 -2758 745 -2720
rect -745 -2786 -740 -2758
rect -712 -2786 -674 -2758
rect -646 -2786 -608 -2758
rect -580 -2786 -542 -2758
rect -514 -2786 -476 -2758
rect -448 -2786 -410 -2758
rect -382 -2786 -344 -2758
rect -316 -2786 -278 -2758
rect -250 -2786 -212 -2758
rect -184 -2786 -146 -2758
rect -118 -2786 -80 -2758
rect -52 -2786 -14 -2758
rect 14 -2786 52 -2758
rect 80 -2786 118 -2758
rect 146 -2786 184 -2758
rect 212 -2786 250 -2758
rect 278 -2786 316 -2758
rect 344 -2786 382 -2758
rect 410 -2786 448 -2758
rect 476 -2786 514 -2758
rect 542 -2786 580 -2758
rect 608 -2786 646 -2758
rect 674 -2786 712 -2758
rect 740 -2786 745 -2758
rect -745 -2824 745 -2786
rect -745 -2852 -740 -2824
rect -712 -2852 -674 -2824
rect -646 -2852 -608 -2824
rect -580 -2852 -542 -2824
rect -514 -2852 -476 -2824
rect -448 -2852 -410 -2824
rect -382 -2852 -344 -2824
rect -316 -2852 -278 -2824
rect -250 -2852 -212 -2824
rect -184 -2852 -146 -2824
rect -118 -2852 -80 -2824
rect -52 -2852 -14 -2824
rect 14 -2852 52 -2824
rect 80 -2852 118 -2824
rect 146 -2852 184 -2824
rect 212 -2852 250 -2824
rect 278 -2852 316 -2824
rect 344 -2852 382 -2824
rect 410 -2852 448 -2824
rect 476 -2852 514 -2824
rect 542 -2852 580 -2824
rect 608 -2852 646 -2824
rect 674 -2852 712 -2824
rect 740 -2852 745 -2824
rect -745 -2890 745 -2852
rect -745 -2918 -740 -2890
rect -712 -2918 -674 -2890
rect -646 -2918 -608 -2890
rect -580 -2918 -542 -2890
rect -514 -2918 -476 -2890
rect -448 -2918 -410 -2890
rect -382 -2918 -344 -2890
rect -316 -2918 -278 -2890
rect -250 -2918 -212 -2890
rect -184 -2918 -146 -2890
rect -118 -2918 -80 -2890
rect -52 -2918 -14 -2890
rect 14 -2918 52 -2890
rect 80 -2918 118 -2890
rect 146 -2918 184 -2890
rect 212 -2918 250 -2890
rect 278 -2918 316 -2890
rect 344 -2918 382 -2890
rect 410 -2918 448 -2890
rect 476 -2918 514 -2890
rect 542 -2918 580 -2890
rect 608 -2918 646 -2890
rect 674 -2918 712 -2890
rect 740 -2918 745 -2890
rect -745 -2956 745 -2918
rect -745 -2984 -740 -2956
rect -712 -2984 -674 -2956
rect -646 -2984 -608 -2956
rect -580 -2984 -542 -2956
rect -514 -2984 -476 -2956
rect -448 -2984 -410 -2956
rect -382 -2984 -344 -2956
rect -316 -2984 -278 -2956
rect -250 -2984 -212 -2956
rect -184 -2984 -146 -2956
rect -118 -2984 -80 -2956
rect -52 -2984 -14 -2956
rect 14 -2984 52 -2956
rect 80 -2984 118 -2956
rect 146 -2984 184 -2956
rect 212 -2984 250 -2956
rect 278 -2984 316 -2956
rect 344 -2984 382 -2956
rect 410 -2984 448 -2956
rect 476 -2984 514 -2956
rect 542 -2984 580 -2956
rect 608 -2984 646 -2956
rect 674 -2984 712 -2956
rect 740 -2984 745 -2956
rect -745 -3022 745 -2984
rect -745 -3050 -740 -3022
rect -712 -3050 -674 -3022
rect -646 -3050 -608 -3022
rect -580 -3050 -542 -3022
rect -514 -3050 -476 -3022
rect -448 -3050 -410 -3022
rect -382 -3050 -344 -3022
rect -316 -3050 -278 -3022
rect -250 -3050 -212 -3022
rect -184 -3050 -146 -3022
rect -118 -3050 -80 -3022
rect -52 -3050 -14 -3022
rect 14 -3050 52 -3022
rect 80 -3050 118 -3022
rect 146 -3050 184 -3022
rect 212 -3050 250 -3022
rect 278 -3050 316 -3022
rect 344 -3050 382 -3022
rect 410 -3050 448 -3022
rect 476 -3050 514 -3022
rect 542 -3050 580 -3022
rect 608 -3050 646 -3022
rect 674 -3050 712 -3022
rect 740 -3050 745 -3022
rect -745 -3088 745 -3050
rect -745 -3116 -740 -3088
rect -712 -3116 -674 -3088
rect -646 -3116 -608 -3088
rect -580 -3116 -542 -3088
rect -514 -3116 -476 -3088
rect -448 -3116 -410 -3088
rect -382 -3116 -344 -3088
rect -316 -3116 -278 -3088
rect -250 -3116 -212 -3088
rect -184 -3116 -146 -3088
rect -118 -3116 -80 -3088
rect -52 -3116 -14 -3088
rect 14 -3116 52 -3088
rect 80 -3116 118 -3088
rect 146 -3116 184 -3088
rect 212 -3116 250 -3088
rect 278 -3116 316 -3088
rect 344 -3116 382 -3088
rect 410 -3116 448 -3088
rect 476 -3116 514 -3088
rect 542 -3116 580 -3088
rect 608 -3116 646 -3088
rect 674 -3116 712 -3088
rect 740 -3116 745 -3088
rect -745 -3154 745 -3116
rect -745 -3182 -740 -3154
rect -712 -3182 -674 -3154
rect -646 -3182 -608 -3154
rect -580 -3182 -542 -3154
rect -514 -3182 -476 -3154
rect -448 -3182 -410 -3154
rect -382 -3182 -344 -3154
rect -316 -3182 -278 -3154
rect -250 -3182 -212 -3154
rect -184 -3182 -146 -3154
rect -118 -3182 -80 -3154
rect -52 -3182 -14 -3154
rect 14 -3182 52 -3154
rect 80 -3182 118 -3154
rect 146 -3182 184 -3154
rect 212 -3182 250 -3154
rect 278 -3182 316 -3154
rect 344 -3182 382 -3154
rect 410 -3182 448 -3154
rect 476 -3182 514 -3154
rect 542 -3182 580 -3154
rect 608 -3182 646 -3154
rect 674 -3182 712 -3154
rect 740 -3182 745 -3154
rect -745 -3220 745 -3182
rect -745 -3248 -740 -3220
rect -712 -3248 -674 -3220
rect -646 -3248 -608 -3220
rect -580 -3248 -542 -3220
rect -514 -3248 -476 -3220
rect -448 -3248 -410 -3220
rect -382 -3248 -344 -3220
rect -316 -3248 -278 -3220
rect -250 -3248 -212 -3220
rect -184 -3248 -146 -3220
rect -118 -3248 -80 -3220
rect -52 -3248 -14 -3220
rect 14 -3248 52 -3220
rect 80 -3248 118 -3220
rect 146 -3248 184 -3220
rect 212 -3248 250 -3220
rect 278 -3248 316 -3220
rect 344 -3248 382 -3220
rect 410 -3248 448 -3220
rect 476 -3248 514 -3220
rect 542 -3248 580 -3220
rect 608 -3248 646 -3220
rect 674 -3248 712 -3220
rect 740 -3248 745 -3220
rect -745 -3286 745 -3248
rect -745 -3314 -740 -3286
rect -712 -3314 -674 -3286
rect -646 -3314 -608 -3286
rect -580 -3314 -542 -3286
rect -514 -3314 -476 -3286
rect -448 -3314 -410 -3286
rect -382 -3314 -344 -3286
rect -316 -3314 -278 -3286
rect -250 -3314 -212 -3286
rect -184 -3314 -146 -3286
rect -118 -3314 -80 -3286
rect -52 -3314 -14 -3286
rect 14 -3314 52 -3286
rect 80 -3314 118 -3286
rect 146 -3314 184 -3286
rect 212 -3314 250 -3286
rect 278 -3314 316 -3286
rect 344 -3314 382 -3286
rect 410 -3314 448 -3286
rect 476 -3314 514 -3286
rect 542 -3314 580 -3286
rect 608 -3314 646 -3286
rect 674 -3314 712 -3286
rect 740 -3314 745 -3286
rect -745 -3352 745 -3314
rect -745 -3380 -740 -3352
rect -712 -3380 -674 -3352
rect -646 -3380 -608 -3352
rect -580 -3380 -542 -3352
rect -514 -3380 -476 -3352
rect -448 -3380 -410 -3352
rect -382 -3380 -344 -3352
rect -316 -3380 -278 -3352
rect -250 -3380 -212 -3352
rect -184 -3380 -146 -3352
rect -118 -3380 -80 -3352
rect -52 -3380 -14 -3352
rect 14 -3380 52 -3352
rect 80 -3380 118 -3352
rect 146 -3380 184 -3352
rect 212 -3380 250 -3352
rect 278 -3380 316 -3352
rect 344 -3380 382 -3352
rect 410 -3380 448 -3352
rect 476 -3380 514 -3352
rect 542 -3380 580 -3352
rect 608 -3380 646 -3352
rect 674 -3380 712 -3352
rect 740 -3380 745 -3352
rect -745 -3418 745 -3380
rect -745 -3446 -740 -3418
rect -712 -3446 -674 -3418
rect -646 -3446 -608 -3418
rect -580 -3446 -542 -3418
rect -514 -3446 -476 -3418
rect -448 -3446 -410 -3418
rect -382 -3446 -344 -3418
rect -316 -3446 -278 -3418
rect -250 -3446 -212 -3418
rect -184 -3446 -146 -3418
rect -118 -3446 -80 -3418
rect -52 -3446 -14 -3418
rect 14 -3446 52 -3418
rect 80 -3446 118 -3418
rect 146 -3446 184 -3418
rect 212 -3446 250 -3418
rect 278 -3446 316 -3418
rect 344 -3446 382 -3418
rect 410 -3446 448 -3418
rect 476 -3446 514 -3418
rect 542 -3446 580 -3418
rect 608 -3446 646 -3418
rect 674 -3446 712 -3418
rect 740 -3446 745 -3418
rect -745 -3484 745 -3446
rect -745 -3512 -740 -3484
rect -712 -3512 -674 -3484
rect -646 -3512 -608 -3484
rect -580 -3512 -542 -3484
rect -514 -3512 -476 -3484
rect -448 -3512 -410 -3484
rect -382 -3512 -344 -3484
rect -316 -3512 -278 -3484
rect -250 -3512 -212 -3484
rect -184 -3512 -146 -3484
rect -118 -3512 -80 -3484
rect -52 -3512 -14 -3484
rect 14 -3512 52 -3484
rect 80 -3512 118 -3484
rect 146 -3512 184 -3484
rect 212 -3512 250 -3484
rect 278 -3512 316 -3484
rect 344 -3512 382 -3484
rect 410 -3512 448 -3484
rect 476 -3512 514 -3484
rect 542 -3512 580 -3484
rect 608 -3512 646 -3484
rect 674 -3512 712 -3484
rect 740 -3512 745 -3484
rect -745 -3550 745 -3512
rect -745 -3578 -740 -3550
rect -712 -3578 -674 -3550
rect -646 -3578 -608 -3550
rect -580 -3578 -542 -3550
rect -514 -3578 -476 -3550
rect -448 -3578 -410 -3550
rect -382 -3578 -344 -3550
rect -316 -3578 -278 -3550
rect -250 -3578 -212 -3550
rect -184 -3578 -146 -3550
rect -118 -3578 -80 -3550
rect -52 -3578 -14 -3550
rect 14 -3578 52 -3550
rect 80 -3578 118 -3550
rect 146 -3578 184 -3550
rect 212 -3578 250 -3550
rect 278 -3578 316 -3550
rect 344 -3578 382 -3550
rect 410 -3578 448 -3550
rect 476 -3578 514 -3550
rect 542 -3578 580 -3550
rect 608 -3578 646 -3550
rect 674 -3578 712 -3550
rect 740 -3578 745 -3550
rect -745 -3616 745 -3578
rect -745 -3644 -740 -3616
rect -712 -3644 -674 -3616
rect -646 -3644 -608 -3616
rect -580 -3644 -542 -3616
rect -514 -3644 -476 -3616
rect -448 -3644 -410 -3616
rect -382 -3644 -344 -3616
rect -316 -3644 -278 -3616
rect -250 -3644 -212 -3616
rect -184 -3644 -146 -3616
rect -118 -3644 -80 -3616
rect -52 -3644 -14 -3616
rect 14 -3644 52 -3616
rect 80 -3644 118 -3616
rect 146 -3644 184 -3616
rect 212 -3644 250 -3616
rect 278 -3644 316 -3616
rect 344 -3644 382 -3616
rect 410 -3644 448 -3616
rect 476 -3644 514 -3616
rect 542 -3644 580 -3616
rect 608 -3644 646 -3616
rect 674 -3644 712 -3616
rect 740 -3644 745 -3616
rect -745 -3682 745 -3644
rect -745 -3710 -740 -3682
rect -712 -3710 -674 -3682
rect -646 -3710 -608 -3682
rect -580 -3710 -542 -3682
rect -514 -3710 -476 -3682
rect -448 -3710 -410 -3682
rect -382 -3710 -344 -3682
rect -316 -3710 -278 -3682
rect -250 -3710 -212 -3682
rect -184 -3710 -146 -3682
rect -118 -3710 -80 -3682
rect -52 -3710 -14 -3682
rect 14 -3710 52 -3682
rect 80 -3710 118 -3682
rect 146 -3710 184 -3682
rect 212 -3710 250 -3682
rect 278 -3710 316 -3682
rect 344 -3710 382 -3682
rect 410 -3710 448 -3682
rect 476 -3710 514 -3682
rect 542 -3710 580 -3682
rect 608 -3710 646 -3682
rect 674 -3710 712 -3682
rect 740 -3710 745 -3682
rect -745 -3748 745 -3710
rect -745 -3776 -740 -3748
rect -712 -3776 -674 -3748
rect -646 -3776 -608 -3748
rect -580 -3776 -542 -3748
rect -514 -3776 -476 -3748
rect -448 -3776 -410 -3748
rect -382 -3776 -344 -3748
rect -316 -3776 -278 -3748
rect -250 -3776 -212 -3748
rect -184 -3776 -146 -3748
rect -118 -3776 -80 -3748
rect -52 -3776 -14 -3748
rect 14 -3776 52 -3748
rect 80 -3776 118 -3748
rect 146 -3776 184 -3748
rect 212 -3776 250 -3748
rect 278 -3776 316 -3748
rect 344 -3776 382 -3748
rect 410 -3776 448 -3748
rect 476 -3776 514 -3748
rect 542 -3776 580 -3748
rect 608 -3776 646 -3748
rect 674 -3776 712 -3748
rect 740 -3776 745 -3748
rect -745 -3814 745 -3776
rect -745 -3842 -740 -3814
rect -712 -3842 -674 -3814
rect -646 -3842 -608 -3814
rect -580 -3842 -542 -3814
rect -514 -3842 -476 -3814
rect -448 -3842 -410 -3814
rect -382 -3842 -344 -3814
rect -316 -3842 -278 -3814
rect -250 -3842 -212 -3814
rect -184 -3842 -146 -3814
rect -118 -3842 -80 -3814
rect -52 -3842 -14 -3814
rect 14 -3842 52 -3814
rect 80 -3842 118 -3814
rect 146 -3842 184 -3814
rect 212 -3842 250 -3814
rect 278 -3842 316 -3814
rect 344 -3842 382 -3814
rect 410 -3842 448 -3814
rect 476 -3842 514 -3814
rect 542 -3842 580 -3814
rect 608 -3842 646 -3814
rect 674 -3842 712 -3814
rect 740 -3842 745 -3814
rect -745 -3880 745 -3842
rect -745 -3908 -740 -3880
rect -712 -3908 -674 -3880
rect -646 -3908 -608 -3880
rect -580 -3908 -542 -3880
rect -514 -3908 -476 -3880
rect -448 -3908 -410 -3880
rect -382 -3908 -344 -3880
rect -316 -3908 -278 -3880
rect -250 -3908 -212 -3880
rect -184 -3908 -146 -3880
rect -118 -3908 -80 -3880
rect -52 -3908 -14 -3880
rect 14 -3908 52 -3880
rect 80 -3908 118 -3880
rect 146 -3908 184 -3880
rect 212 -3908 250 -3880
rect 278 -3908 316 -3880
rect 344 -3908 382 -3880
rect 410 -3908 448 -3880
rect 476 -3908 514 -3880
rect 542 -3908 580 -3880
rect 608 -3908 646 -3880
rect 674 -3908 712 -3880
rect 740 -3908 745 -3880
rect -745 -3946 745 -3908
rect -745 -3974 -740 -3946
rect -712 -3974 -674 -3946
rect -646 -3974 -608 -3946
rect -580 -3974 -542 -3946
rect -514 -3974 -476 -3946
rect -448 -3974 -410 -3946
rect -382 -3974 -344 -3946
rect -316 -3974 -278 -3946
rect -250 -3974 -212 -3946
rect -184 -3974 -146 -3946
rect -118 -3974 -80 -3946
rect -52 -3974 -14 -3946
rect 14 -3974 52 -3946
rect 80 -3974 118 -3946
rect 146 -3974 184 -3946
rect 212 -3974 250 -3946
rect 278 -3974 316 -3946
rect 344 -3974 382 -3946
rect 410 -3974 448 -3946
rect 476 -3974 514 -3946
rect 542 -3974 580 -3946
rect 608 -3974 646 -3946
rect 674 -3974 712 -3946
rect 740 -3974 745 -3946
rect -745 -4012 745 -3974
rect -745 -4040 -740 -4012
rect -712 -4040 -674 -4012
rect -646 -4040 -608 -4012
rect -580 -4040 -542 -4012
rect -514 -4040 -476 -4012
rect -448 -4040 -410 -4012
rect -382 -4040 -344 -4012
rect -316 -4040 -278 -4012
rect -250 -4040 -212 -4012
rect -184 -4040 -146 -4012
rect -118 -4040 -80 -4012
rect -52 -4040 -14 -4012
rect 14 -4040 52 -4012
rect 80 -4040 118 -4012
rect 146 -4040 184 -4012
rect 212 -4040 250 -4012
rect 278 -4040 316 -4012
rect 344 -4040 382 -4012
rect 410 -4040 448 -4012
rect 476 -4040 514 -4012
rect 542 -4040 580 -4012
rect 608 -4040 646 -4012
rect 674 -4040 712 -4012
rect 740 -4040 745 -4012
rect -745 -4078 745 -4040
rect -745 -4106 -740 -4078
rect -712 -4106 -674 -4078
rect -646 -4106 -608 -4078
rect -580 -4106 -542 -4078
rect -514 -4106 -476 -4078
rect -448 -4106 -410 -4078
rect -382 -4106 -344 -4078
rect -316 -4106 -278 -4078
rect -250 -4106 -212 -4078
rect -184 -4106 -146 -4078
rect -118 -4106 -80 -4078
rect -52 -4106 -14 -4078
rect 14 -4106 52 -4078
rect 80 -4106 118 -4078
rect 146 -4106 184 -4078
rect 212 -4106 250 -4078
rect 278 -4106 316 -4078
rect 344 -4106 382 -4078
rect 410 -4106 448 -4078
rect 476 -4106 514 -4078
rect 542 -4106 580 -4078
rect 608 -4106 646 -4078
rect 674 -4106 712 -4078
rect 740 -4106 745 -4078
rect -745 -4144 745 -4106
rect -745 -4172 -740 -4144
rect -712 -4172 -674 -4144
rect -646 -4172 -608 -4144
rect -580 -4172 -542 -4144
rect -514 -4172 -476 -4144
rect -448 -4172 -410 -4144
rect -382 -4172 -344 -4144
rect -316 -4172 -278 -4144
rect -250 -4172 -212 -4144
rect -184 -4172 -146 -4144
rect -118 -4172 -80 -4144
rect -52 -4172 -14 -4144
rect 14 -4172 52 -4144
rect 80 -4172 118 -4144
rect 146 -4172 184 -4144
rect 212 -4172 250 -4144
rect 278 -4172 316 -4144
rect 344 -4172 382 -4144
rect 410 -4172 448 -4144
rect 476 -4172 514 -4144
rect 542 -4172 580 -4144
rect 608 -4172 646 -4144
rect 674 -4172 712 -4144
rect 740 -4172 745 -4144
rect -745 -4210 745 -4172
rect -745 -4238 -740 -4210
rect -712 -4238 -674 -4210
rect -646 -4238 -608 -4210
rect -580 -4238 -542 -4210
rect -514 -4238 -476 -4210
rect -448 -4238 -410 -4210
rect -382 -4238 -344 -4210
rect -316 -4238 -278 -4210
rect -250 -4238 -212 -4210
rect -184 -4238 -146 -4210
rect -118 -4238 -80 -4210
rect -52 -4238 -14 -4210
rect 14 -4238 52 -4210
rect 80 -4238 118 -4210
rect 146 -4238 184 -4210
rect 212 -4238 250 -4210
rect 278 -4238 316 -4210
rect 344 -4238 382 -4210
rect 410 -4238 448 -4210
rect 476 -4238 514 -4210
rect 542 -4238 580 -4210
rect 608 -4238 646 -4210
rect 674 -4238 712 -4210
rect 740 -4238 745 -4210
rect -745 -4276 745 -4238
rect -745 -4304 -740 -4276
rect -712 -4304 -674 -4276
rect -646 -4304 -608 -4276
rect -580 -4304 -542 -4276
rect -514 -4304 -476 -4276
rect -448 -4304 -410 -4276
rect -382 -4304 -344 -4276
rect -316 -4304 -278 -4276
rect -250 -4304 -212 -4276
rect -184 -4304 -146 -4276
rect -118 -4304 -80 -4276
rect -52 -4304 -14 -4276
rect 14 -4304 52 -4276
rect 80 -4304 118 -4276
rect 146 -4304 184 -4276
rect 212 -4304 250 -4276
rect 278 -4304 316 -4276
rect 344 -4304 382 -4276
rect 410 -4304 448 -4276
rect 476 -4304 514 -4276
rect 542 -4304 580 -4276
rect 608 -4304 646 -4276
rect 674 -4304 712 -4276
rect 740 -4304 745 -4276
rect -745 -4342 745 -4304
rect -745 -4370 -740 -4342
rect -712 -4370 -674 -4342
rect -646 -4370 -608 -4342
rect -580 -4370 -542 -4342
rect -514 -4370 -476 -4342
rect -448 -4370 -410 -4342
rect -382 -4370 -344 -4342
rect -316 -4370 -278 -4342
rect -250 -4370 -212 -4342
rect -184 -4370 -146 -4342
rect -118 -4370 -80 -4342
rect -52 -4370 -14 -4342
rect 14 -4370 52 -4342
rect 80 -4370 118 -4342
rect 146 -4370 184 -4342
rect 212 -4370 250 -4342
rect 278 -4370 316 -4342
rect 344 -4370 382 -4342
rect 410 -4370 448 -4342
rect 476 -4370 514 -4342
rect 542 -4370 580 -4342
rect 608 -4370 646 -4342
rect 674 -4370 712 -4342
rect 740 -4370 745 -4342
rect -745 -4408 745 -4370
rect -745 -4436 -740 -4408
rect -712 -4436 -674 -4408
rect -646 -4436 -608 -4408
rect -580 -4436 -542 -4408
rect -514 -4436 -476 -4408
rect -448 -4436 -410 -4408
rect -382 -4436 -344 -4408
rect -316 -4436 -278 -4408
rect -250 -4436 -212 -4408
rect -184 -4436 -146 -4408
rect -118 -4436 -80 -4408
rect -52 -4436 -14 -4408
rect 14 -4436 52 -4408
rect 80 -4436 118 -4408
rect 146 -4436 184 -4408
rect 212 -4436 250 -4408
rect 278 -4436 316 -4408
rect 344 -4436 382 -4408
rect 410 -4436 448 -4408
rect 476 -4436 514 -4408
rect 542 -4436 580 -4408
rect 608 -4436 646 -4408
rect 674 -4436 712 -4408
rect 740 -4436 745 -4408
rect -745 -4474 745 -4436
rect -745 -4502 -740 -4474
rect -712 -4502 -674 -4474
rect -646 -4502 -608 -4474
rect -580 -4502 -542 -4474
rect -514 -4502 -476 -4474
rect -448 -4502 -410 -4474
rect -382 -4502 -344 -4474
rect -316 -4502 -278 -4474
rect -250 -4502 -212 -4474
rect -184 -4502 -146 -4474
rect -118 -4502 -80 -4474
rect -52 -4502 -14 -4474
rect 14 -4502 52 -4474
rect 80 -4502 118 -4474
rect 146 -4502 184 -4474
rect 212 -4502 250 -4474
rect 278 -4502 316 -4474
rect 344 -4502 382 -4474
rect 410 -4502 448 -4474
rect 476 -4502 514 -4474
rect 542 -4502 580 -4474
rect 608 -4502 646 -4474
rect 674 -4502 712 -4474
rect 740 -4502 745 -4474
rect -745 -4540 745 -4502
rect -745 -4568 -740 -4540
rect -712 -4568 -674 -4540
rect -646 -4568 -608 -4540
rect -580 -4568 -542 -4540
rect -514 -4568 -476 -4540
rect -448 -4568 -410 -4540
rect -382 -4568 -344 -4540
rect -316 -4568 -278 -4540
rect -250 -4568 -212 -4540
rect -184 -4568 -146 -4540
rect -118 -4568 -80 -4540
rect -52 -4568 -14 -4540
rect 14 -4568 52 -4540
rect 80 -4568 118 -4540
rect 146 -4568 184 -4540
rect 212 -4568 250 -4540
rect 278 -4568 316 -4540
rect 344 -4568 382 -4540
rect 410 -4568 448 -4540
rect 476 -4568 514 -4540
rect 542 -4568 580 -4540
rect 608 -4568 646 -4540
rect 674 -4568 712 -4540
rect 740 -4568 745 -4540
rect -745 -4606 745 -4568
rect -745 -4634 -740 -4606
rect -712 -4634 -674 -4606
rect -646 -4634 -608 -4606
rect -580 -4634 -542 -4606
rect -514 -4634 -476 -4606
rect -448 -4634 -410 -4606
rect -382 -4634 -344 -4606
rect -316 -4634 -278 -4606
rect -250 -4634 -212 -4606
rect -184 -4634 -146 -4606
rect -118 -4634 -80 -4606
rect -52 -4634 -14 -4606
rect 14 -4634 52 -4606
rect 80 -4634 118 -4606
rect 146 -4634 184 -4606
rect 212 -4634 250 -4606
rect 278 -4634 316 -4606
rect 344 -4634 382 -4606
rect 410 -4634 448 -4606
rect 476 -4634 514 -4606
rect 542 -4634 580 -4606
rect 608 -4634 646 -4606
rect 674 -4634 712 -4606
rect 740 -4634 745 -4606
rect -745 -4672 745 -4634
rect -745 -4700 -740 -4672
rect -712 -4700 -674 -4672
rect -646 -4700 -608 -4672
rect -580 -4700 -542 -4672
rect -514 -4700 -476 -4672
rect -448 -4700 -410 -4672
rect -382 -4700 -344 -4672
rect -316 -4700 -278 -4672
rect -250 -4700 -212 -4672
rect -184 -4700 -146 -4672
rect -118 -4700 -80 -4672
rect -52 -4700 -14 -4672
rect 14 -4700 52 -4672
rect 80 -4700 118 -4672
rect 146 -4700 184 -4672
rect 212 -4700 250 -4672
rect 278 -4700 316 -4672
rect 344 -4700 382 -4672
rect 410 -4700 448 -4672
rect 476 -4700 514 -4672
rect 542 -4700 580 -4672
rect 608 -4700 646 -4672
rect 674 -4700 712 -4672
rect 740 -4700 745 -4672
rect -745 -4738 745 -4700
rect -745 -4766 -740 -4738
rect -712 -4766 -674 -4738
rect -646 -4766 -608 -4738
rect -580 -4766 -542 -4738
rect -514 -4766 -476 -4738
rect -448 -4766 -410 -4738
rect -382 -4766 -344 -4738
rect -316 -4766 -278 -4738
rect -250 -4766 -212 -4738
rect -184 -4766 -146 -4738
rect -118 -4766 -80 -4738
rect -52 -4766 -14 -4738
rect 14 -4766 52 -4738
rect 80 -4766 118 -4738
rect 146 -4766 184 -4738
rect 212 -4766 250 -4738
rect 278 -4766 316 -4738
rect 344 -4766 382 -4738
rect 410 -4766 448 -4738
rect 476 -4766 514 -4738
rect 542 -4766 580 -4738
rect 608 -4766 646 -4738
rect 674 -4766 712 -4738
rect 740 -4766 745 -4738
rect -745 -4804 745 -4766
rect -745 -4832 -740 -4804
rect -712 -4832 -674 -4804
rect -646 -4832 -608 -4804
rect -580 -4832 -542 -4804
rect -514 -4832 -476 -4804
rect -448 -4832 -410 -4804
rect -382 -4832 -344 -4804
rect -316 -4832 -278 -4804
rect -250 -4832 -212 -4804
rect -184 -4832 -146 -4804
rect -118 -4832 -80 -4804
rect -52 -4832 -14 -4804
rect 14 -4832 52 -4804
rect 80 -4832 118 -4804
rect 146 -4832 184 -4804
rect 212 -4832 250 -4804
rect 278 -4832 316 -4804
rect 344 -4832 382 -4804
rect 410 -4832 448 -4804
rect 476 -4832 514 -4804
rect 542 -4832 580 -4804
rect 608 -4832 646 -4804
rect 674 -4832 712 -4804
rect 740 -4832 745 -4804
rect -745 -4870 745 -4832
rect -745 -4898 -740 -4870
rect -712 -4898 -674 -4870
rect -646 -4898 -608 -4870
rect -580 -4898 -542 -4870
rect -514 -4898 -476 -4870
rect -448 -4898 -410 -4870
rect -382 -4898 -344 -4870
rect -316 -4898 -278 -4870
rect -250 -4898 -212 -4870
rect -184 -4898 -146 -4870
rect -118 -4898 -80 -4870
rect -52 -4898 -14 -4870
rect 14 -4898 52 -4870
rect 80 -4898 118 -4870
rect 146 -4898 184 -4870
rect 212 -4898 250 -4870
rect 278 -4898 316 -4870
rect 344 -4898 382 -4870
rect 410 -4898 448 -4870
rect 476 -4898 514 -4870
rect 542 -4898 580 -4870
rect 608 -4898 646 -4870
rect 674 -4898 712 -4870
rect 740 -4898 745 -4870
rect -745 -4936 745 -4898
rect -745 -4964 -740 -4936
rect -712 -4964 -674 -4936
rect -646 -4964 -608 -4936
rect -580 -4964 -542 -4936
rect -514 -4964 -476 -4936
rect -448 -4964 -410 -4936
rect -382 -4964 -344 -4936
rect -316 -4964 -278 -4936
rect -250 -4964 -212 -4936
rect -184 -4964 -146 -4936
rect -118 -4964 -80 -4936
rect -52 -4964 -14 -4936
rect 14 -4964 52 -4936
rect 80 -4964 118 -4936
rect 146 -4964 184 -4936
rect 212 -4964 250 -4936
rect 278 -4964 316 -4936
rect 344 -4964 382 -4936
rect 410 -4964 448 -4936
rect 476 -4964 514 -4936
rect 542 -4964 580 -4936
rect 608 -4964 646 -4936
rect 674 -4964 712 -4936
rect 740 -4964 745 -4936
rect -745 -5002 745 -4964
rect -745 -5030 -740 -5002
rect -712 -5030 -674 -5002
rect -646 -5030 -608 -5002
rect -580 -5030 -542 -5002
rect -514 -5030 -476 -5002
rect -448 -5030 -410 -5002
rect -382 -5030 -344 -5002
rect -316 -5030 -278 -5002
rect -250 -5030 -212 -5002
rect -184 -5030 -146 -5002
rect -118 -5030 -80 -5002
rect -52 -5030 -14 -5002
rect 14 -5030 52 -5002
rect 80 -5030 118 -5002
rect 146 -5030 184 -5002
rect 212 -5030 250 -5002
rect 278 -5030 316 -5002
rect 344 -5030 382 -5002
rect 410 -5030 448 -5002
rect 476 -5030 514 -5002
rect 542 -5030 580 -5002
rect 608 -5030 646 -5002
rect 674 -5030 712 -5002
rect 740 -5030 745 -5002
rect -745 -5068 745 -5030
rect -745 -5096 -740 -5068
rect -712 -5096 -674 -5068
rect -646 -5096 -608 -5068
rect -580 -5096 -542 -5068
rect -514 -5096 -476 -5068
rect -448 -5096 -410 -5068
rect -382 -5096 -344 -5068
rect -316 -5096 -278 -5068
rect -250 -5096 -212 -5068
rect -184 -5096 -146 -5068
rect -118 -5096 -80 -5068
rect -52 -5096 -14 -5068
rect 14 -5096 52 -5068
rect 80 -5096 118 -5068
rect 146 -5096 184 -5068
rect 212 -5096 250 -5068
rect 278 -5096 316 -5068
rect 344 -5096 382 -5068
rect 410 -5096 448 -5068
rect 476 -5096 514 -5068
rect 542 -5096 580 -5068
rect 608 -5096 646 -5068
rect 674 -5096 712 -5068
rect 740 -5096 745 -5068
rect -745 -5134 745 -5096
rect -745 -5162 -740 -5134
rect -712 -5162 -674 -5134
rect -646 -5162 -608 -5134
rect -580 -5162 -542 -5134
rect -514 -5162 -476 -5134
rect -448 -5162 -410 -5134
rect -382 -5162 -344 -5134
rect -316 -5162 -278 -5134
rect -250 -5162 -212 -5134
rect -184 -5162 -146 -5134
rect -118 -5162 -80 -5134
rect -52 -5162 -14 -5134
rect 14 -5162 52 -5134
rect 80 -5162 118 -5134
rect 146 -5162 184 -5134
rect 212 -5162 250 -5134
rect 278 -5162 316 -5134
rect 344 -5162 382 -5134
rect 410 -5162 448 -5134
rect 476 -5162 514 -5134
rect 542 -5162 580 -5134
rect 608 -5162 646 -5134
rect 674 -5162 712 -5134
rect 740 -5162 745 -5134
rect -745 -5200 745 -5162
rect -745 -5228 -740 -5200
rect -712 -5228 -674 -5200
rect -646 -5228 -608 -5200
rect -580 -5228 -542 -5200
rect -514 -5228 -476 -5200
rect -448 -5228 -410 -5200
rect -382 -5228 -344 -5200
rect -316 -5228 -278 -5200
rect -250 -5228 -212 -5200
rect -184 -5228 -146 -5200
rect -118 -5228 -80 -5200
rect -52 -5228 -14 -5200
rect 14 -5228 52 -5200
rect 80 -5228 118 -5200
rect 146 -5228 184 -5200
rect 212 -5228 250 -5200
rect 278 -5228 316 -5200
rect 344 -5228 382 -5200
rect 410 -5228 448 -5200
rect 476 -5228 514 -5200
rect 542 -5228 580 -5200
rect 608 -5228 646 -5200
rect 674 -5228 712 -5200
rect 740 -5228 745 -5200
rect -745 -5266 745 -5228
rect -745 -5294 -740 -5266
rect -712 -5294 -674 -5266
rect -646 -5294 -608 -5266
rect -580 -5294 -542 -5266
rect -514 -5294 -476 -5266
rect -448 -5294 -410 -5266
rect -382 -5294 -344 -5266
rect -316 -5294 -278 -5266
rect -250 -5294 -212 -5266
rect -184 -5294 -146 -5266
rect -118 -5294 -80 -5266
rect -52 -5294 -14 -5266
rect 14 -5294 52 -5266
rect 80 -5294 118 -5266
rect 146 -5294 184 -5266
rect 212 -5294 250 -5266
rect 278 -5294 316 -5266
rect 344 -5294 382 -5266
rect 410 -5294 448 -5266
rect 476 -5294 514 -5266
rect 542 -5294 580 -5266
rect 608 -5294 646 -5266
rect 674 -5294 712 -5266
rect 740 -5294 745 -5266
rect -745 -5332 745 -5294
rect -745 -5360 -740 -5332
rect -712 -5360 -674 -5332
rect -646 -5360 -608 -5332
rect -580 -5360 -542 -5332
rect -514 -5360 -476 -5332
rect -448 -5360 -410 -5332
rect -382 -5360 -344 -5332
rect -316 -5360 -278 -5332
rect -250 -5360 -212 -5332
rect -184 -5360 -146 -5332
rect -118 -5360 -80 -5332
rect -52 -5360 -14 -5332
rect 14 -5360 52 -5332
rect 80 -5360 118 -5332
rect 146 -5360 184 -5332
rect 212 -5360 250 -5332
rect 278 -5360 316 -5332
rect 344 -5360 382 -5332
rect 410 -5360 448 -5332
rect 476 -5360 514 -5332
rect 542 -5360 580 -5332
rect 608 -5360 646 -5332
rect 674 -5360 712 -5332
rect 740 -5360 745 -5332
rect -745 -5398 745 -5360
rect -745 -5426 -740 -5398
rect -712 -5426 -674 -5398
rect -646 -5426 -608 -5398
rect -580 -5426 -542 -5398
rect -514 -5426 -476 -5398
rect -448 -5426 -410 -5398
rect -382 -5426 -344 -5398
rect -316 -5426 -278 -5398
rect -250 -5426 -212 -5398
rect -184 -5426 -146 -5398
rect -118 -5426 -80 -5398
rect -52 -5426 -14 -5398
rect 14 -5426 52 -5398
rect 80 -5426 118 -5398
rect 146 -5426 184 -5398
rect 212 -5426 250 -5398
rect 278 -5426 316 -5398
rect 344 -5426 382 -5398
rect 410 -5426 448 -5398
rect 476 -5426 514 -5398
rect 542 -5426 580 -5398
rect 608 -5426 646 -5398
rect 674 -5426 712 -5398
rect 740 -5426 745 -5398
rect -745 -5464 745 -5426
rect -745 -5492 -740 -5464
rect -712 -5492 -674 -5464
rect -646 -5492 -608 -5464
rect -580 -5492 -542 -5464
rect -514 -5492 -476 -5464
rect -448 -5492 -410 -5464
rect -382 -5492 -344 -5464
rect -316 -5492 -278 -5464
rect -250 -5492 -212 -5464
rect -184 -5492 -146 -5464
rect -118 -5492 -80 -5464
rect -52 -5492 -14 -5464
rect 14 -5492 52 -5464
rect 80 -5492 118 -5464
rect 146 -5492 184 -5464
rect 212 -5492 250 -5464
rect 278 -5492 316 -5464
rect 344 -5492 382 -5464
rect 410 -5492 448 -5464
rect 476 -5492 514 -5464
rect 542 -5492 580 -5464
rect 608 -5492 646 -5464
rect 674 -5492 712 -5464
rect 740 -5492 745 -5464
rect -745 -5530 745 -5492
rect -745 -5558 -740 -5530
rect -712 -5558 -674 -5530
rect -646 -5558 -608 -5530
rect -580 -5558 -542 -5530
rect -514 -5558 -476 -5530
rect -448 -5558 -410 -5530
rect -382 -5558 -344 -5530
rect -316 -5558 -278 -5530
rect -250 -5558 -212 -5530
rect -184 -5558 -146 -5530
rect -118 -5558 -80 -5530
rect -52 -5558 -14 -5530
rect 14 -5558 52 -5530
rect 80 -5558 118 -5530
rect 146 -5558 184 -5530
rect 212 -5558 250 -5530
rect 278 -5558 316 -5530
rect 344 -5558 382 -5530
rect 410 -5558 448 -5530
rect 476 -5558 514 -5530
rect 542 -5558 580 -5530
rect 608 -5558 646 -5530
rect 674 -5558 712 -5530
rect 740 -5558 745 -5530
rect -745 -5563 745 -5558
<< end >>
