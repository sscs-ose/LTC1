magic
tech gf180mcuC
magscale 1 10
timestamp 1691593880
<< error_p >>
rect -295 133 -284 179
rect -121 133 -110 179
rect 53 133 64 179
rect 227 133 238 179
rect -295 -179 -284 -133
rect -121 -179 -110 -133
rect 53 -179 64 -133
rect 227 -179 238 -133
<< pwell >>
rect -546 -308 546 308
<< nmos >>
rect -296 -100 -226 100
rect -122 -100 -52 100
rect 52 -100 122 100
rect 226 -100 296 100
<< ndiff >>
rect -384 87 -296 100
rect -384 -87 -371 87
rect -325 -87 -296 87
rect -384 -100 -296 -87
rect -226 87 -122 100
rect -226 -87 -197 87
rect -151 -87 -122 87
rect -226 -100 -122 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 122 87 226 100
rect 122 -87 151 87
rect 197 -87 226 87
rect 122 -100 226 -87
rect 296 87 384 100
rect 296 -87 325 87
rect 371 -87 384 87
rect 296 -100 384 -87
<< ndiffc >>
rect -371 -87 -325 87
rect -197 -87 -151 87
rect -23 -87 23 87
rect 151 -87 197 87
rect 325 -87 371 87
<< psubdiff >>
rect -522 212 522 284
rect -522 168 -450 212
rect -522 -168 -509 168
rect -463 -168 -450 168
rect 450 168 522 212
rect -522 -212 -450 -168
rect 450 -168 463 168
rect 509 -168 522 168
rect 450 -212 522 -168
rect -522 -284 522 -212
<< psubdiffcont >>
rect -509 -168 -463 168
rect 463 -168 509 168
<< polysilicon >>
rect -297 179 -225 192
rect -297 133 -284 179
rect -238 133 -225 179
rect -297 120 -225 133
rect -123 179 -51 192
rect -123 133 -110 179
rect -64 133 -51 179
rect -123 120 -51 133
rect 51 179 123 192
rect 51 133 64 179
rect 110 133 123 179
rect 51 120 123 133
rect 225 179 297 192
rect 225 133 238 179
rect 284 133 297 179
rect 225 120 297 133
rect -296 100 -226 120
rect -122 100 -52 120
rect 52 100 122 120
rect 226 100 296 120
rect -296 -120 -226 -100
rect -122 -120 -52 -100
rect 52 -120 122 -100
rect 226 -120 296 -100
rect -297 -133 -225 -120
rect -297 -179 -284 -133
rect -238 -179 -225 -133
rect -297 -192 -225 -179
rect -123 -133 -51 -120
rect -123 -179 -110 -133
rect -64 -179 -51 -133
rect -123 -192 -51 -179
rect 51 -133 123 -120
rect 51 -179 64 -133
rect 110 -179 123 -133
rect 51 -192 123 -179
rect 225 -133 297 -120
rect 225 -179 238 -133
rect 284 -179 297 -133
rect 225 -192 297 -179
<< polycontact >>
rect -284 133 -238 179
rect -110 133 -64 179
rect 64 133 110 179
rect 238 133 284 179
rect -284 -179 -238 -133
rect -110 -179 -64 -133
rect 64 -179 110 -133
rect 238 -179 284 -133
<< metal1 >>
rect -509 225 509 271
rect -509 168 -463 225
rect -295 133 -284 179
rect -238 133 -227 179
rect -121 133 -110 179
rect -64 133 -53 179
rect 53 133 64 179
rect 110 133 121 179
rect 227 133 238 179
rect 284 133 295 179
rect 463 168 509 225
rect -371 87 -325 98
rect -371 -98 -325 -87
rect -197 87 -151 98
rect -197 -98 -151 -87
rect -23 87 23 98
rect -23 -98 23 -87
rect 151 87 197 98
rect 151 -98 197 -87
rect 325 87 371 98
rect 325 -98 371 -87
rect -509 -225 -463 -168
rect -295 -179 -284 -133
rect -238 -179 -227 -133
rect -121 -179 -110 -133
rect -64 -179 -53 -133
rect 53 -179 64 -133
rect 110 -179 121 -133
rect 227 -179 238 -133
rect 284 -179 295 -133
rect 463 -225 509 -168
rect -509 -271 509 -225
<< properties >>
string FIXED_BBOX -486 -248 486 248
string gencell nmos_3p3
string library gf180mcu
string parameters w 1 l 0.35 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 1 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
