* NGSPICE file created from PLL_TOP_MUX_flat.ext - technology: gf180mcuC

.subckt PLL_TOP_MUX_flat S3 S2 S6 UP_INPUT PRE_SCALAR ITAIL1 OUTB VCTRL_IN S4 ITAIL
+ DIV_OUT DN_INPUT UP DN S1 VCTRL2 F_IN OUT VSS VDD
X0 a_42928_8770# a_43228_8148# VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X1 RES_74k_1.M VSS.t415 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X2 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.IN VSS.t425 VSS.t424 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.5u
X3 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN VDD.t419 VDD.t264 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X4 a_24437_9224# PFD_T2_0.INV_mag_0.IN VDD.t444 VDD.t443 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X5 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VSS.t134 VSS.t133 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X6 a_25706_n567# VCTRL2.t0 VSS.t149 VSS.t148 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X7 a_27875_9714# DN_INPUT.t0 VDD.t256 VDD.t255 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X8 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t360 VDD.t320 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X9 RES_74k_1.M VSS.t414 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X10 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VSS.t622 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X11 VSS VCTRL2.t1 a_25706_n567# VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X12 VSS mux_magic_3.OR_magic_0.A a_21443_9476# VSS.t726 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X13 a_43528_12082# a_43828_11460# VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X14 a_19897_11741# mux_magic_2.AND2_magic_0.A a_20097_11741# VSS.t662 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X15 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t338 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X16 VSS PFD_T2_0.Buffer_V_2_0.IN a_25557_8739# VSS.t166 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X17 a_34443_2598# VCTRL2.t2 VSS.t154 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X18 VSS.t283 VSS.t281 VSS.t283 VSS.t282 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X19 RES_74k_1.M VSS.t413 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X20 RES_74k_1.M VSS.t412 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X21 RES_74k_1.P RES_74k_1.P VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X22 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK VCO_DFF_C_0.VCTRL VSS.t108 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X23 VDD a_22967_8787# PFD_T2_0.INV_mag_1.IN VDD.t288 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X24 RES_74k_1.P RES_74k_1.P VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X25 VSS VCTRL2.t3 a_34443_2598# VSS.t155 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X26 a_21443_8068# mux_magic_3.OR_magic_0.A VDD.t787 VDD.t783 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X27 RES_74k_1.M VSS.t411 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X28 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.OUTB VSS.t756 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X29 VSS S6.t0 mux_magic_3.AND2_magic_0.A VSS.t169 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X30 a_29415_8145# mux_magic_1.OR_magic_0.B a_29415_9553# VDD.t474 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X31 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t12 VSS.t765 VSS.t625 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X32 a_25706_n567# VCTRL2.t4 VSS.t159 VSS.t158 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X33 VDD a_22967_8787# PFD_T2_0.INV_mag_1.IN VDD.t285 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X34 a_43828_11254# a_43528_10632# VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X35 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUT.t11 VSS.t630 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X36 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL VDD.t180 VDD.t147 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X37 VSS PFD_T2_0.INV_mag_1.OUT a_22879_10704# VSS.t5 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X38 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.IN VDD.t418 VDD.t417 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X39 VDD.t244 VDD.t242 VDD.t244 VDD.t243 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X40 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t706 VDD.t575 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X41 VDD.t241 VDD.t240 VDD.t241 VDD.t182 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X42 RES_74k_1.M VSS.t410 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X43 a_27875_8520# mux_magic_1.AND2_magic_0.A VDD.t381 VDD.t380 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X44 VSS.t280 VSS.t279 VSS.t280 VSS.t218 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X45 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT a_34443_2598# VSS.t503 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X46 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t520 VDD.t320 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X47 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCTRL VDD.t179 VDD.t152 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X48 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t338 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X49 VDD.t239 VDD.t237 VDD.t239 VDD.t238 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X50 RES_74k_1.M VSS.t409 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X51 mux_magic_2.OR_magic_0.B a_19897_10547# VDD.t544 VDD.t543 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X52 RES_74k_1.M VSS.t408 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X53 a_22966_11778# PFD_T2_0.INV_mag_0.OUT a_22879_10704# VSS.t701 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X54 a_27875_9714# S3.t0 VDD.t796 VDD.t795 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X55 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT a_34443_2598# VSS.t93 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X56 a_34443_2598# VCTRL2.t5 VSS.t161 VSS.t160 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X57 RES_74k_1.M VSS.t407 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X58 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t347 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X59 VSS VCTRL2.t6 a_34443_2598# VSS.t162 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X60 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_44716_n517# VSS.t651 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X61 VSS.t278 VSS.t277 VSS.t278 VSS.t270 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X62 VDD mux_magic_1.AND2_magic_0.A a_27875_8520# VDD.t377 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X63 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VSS.t79 VSS.t78 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X64 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT VDD.t133 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X65 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VSS.t82 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X66 a_22967_8787# PFD_T2_0.INV_mag_0.OUT a_22880_9797# VSS.t137 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X67 VSS ITAIL1.t6 ITAIL1.t7 VSS.t46 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X68 RES_74k_1.P RES_74k_1.P VDD.t54 ppolyf_u r_width=1.1u r_length=2.6u
X69 RES_74k_1.M VSS.t406 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X70 VSS.t276 VSS.t274 VSS.t276 VSS.t275 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X71 mux_magic_3.AND2_magic_0.A S6.t1 VDD.t398 VDD.t397 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X72 a_31940_9626# UP.t3 VSS.t145 VSS.t120 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X73 a_31940_9626# UP.t4 VSS.t660 VSS.t659 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X74 VDD S3.t1 a_27875_9714# VDD.t797 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X75 VSS.t273 VSS.t272 VSS.t273 VSS.t229 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X76 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t606 VDD.t598 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X77 a_20103_8443# DIV_OUT.t0 VSS.t56 VSS.t55 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X78 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCTRL VDD.t178 VDD.t149 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X79 a_44728_10426# a_44428_9804# VDD.t54 ppolyf_u r_width=1.1u r_length=2.6u
X80 VDD S4.t0 A_MUX_0.Tr_Gate_1.CLK VDD.t85 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X81 RES_74k_1.M VSS.t405 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X82 a_42628_9598# a_42928_8976# VDD.t93 ppolyf_u r_width=1.1u r_length=2.6u
X83 VSS.t271 VSS.t269 VSS.t271 VSS.t270 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X84 a_44728_12082# a_44428_11460# VDD.t54 ppolyf_u r_width=1.1u r_length=2.6u
X85 a_20103_9637# VSS.t266 VSS.t268 VSS.t267 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X86 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VSS.t586 VSS.t131 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X87 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VSS.t496 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X88 PFD_T2_0.FIN a_21437_10708# VSS.t136 VSS.t135 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X89 a_41879_1284# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VSS.t656 VSS.t652 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X90 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.IN VDD.t442 VDD.t417 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X91 a_27722_10564# S2.t0 a_27922_10564# VSS.t764 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X92 a_41879_1284# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD.t650 VDD.t260 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X93 a_25706_n567# VCTRL2.t7 VSS.t165 VSS.t148 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X94 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT a_25706_n567# VSS.t81 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X95 VSS S1.t0 mux_magic_2.AND2_magic_0.A VSS.t590 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X96 a_44428_11254# a_44728_10632# VDD.t54 ppolyf_u r_width=1.1u r_length=2.6u
X97 a_19897_11741# PRE_SCALAR.t0 VDD.t726 VDD.t725 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X98 VSS OUT.t13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VSS.t630 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X99 VSS VCTRL2.t8 a_25706_n567# VSS.t451 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X100 a_27722_11758# mux_magic_0.AND2_magic_0.A a_27922_11758# VSS.t54 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X101 ITAIL ITAIL.t14 VDD.t558 VDD.t537 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X102 a_29262_12133# mux_magic_0.OR_magic_0.A VDD.t482 VDD.t1 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X103 VSS PFD_T2_0.INV_mag_0.IN a_23836_10693# VSS.t475 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X104 VSS S3.t2 mux_magic_1.AND2_magic_0.A VSS.t740 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X105 a_45928_10426# a_46228_9804# VDD.t56 ppolyf_u r_width=1.1u r_length=2.6u
X106 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t605 VDD.t570 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X107 a_44428_9598# a_44128_8976# VDD.t55 ppolyf_u r_width=1.1u r_length=2.6u
X108 VDD S4.t1 a_42763_5679# VDD.t78 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X109 RES_74k_1.M VSS.t404 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X110 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB VSS.t499 VSS.t498 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X111 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD.t826 VDD.t819 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X112 RES_74k_1.M VSS.t403 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X113 a_27922_10564# S2.t1 a_27722_10564# VSS.t732 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X114 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t355 VDD.t336 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X115 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VSS.t80 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X116 a_29262_12133# mux_magic_0.OR_magic_0.A VDD.t481 VDD.t477 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X117 a_45928_8770# a_45628_8148# VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X118 OUTB a_41879_1284# VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD.t261 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X119 a_42628_8770# a_42628_8148# VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X120 RES_74k_1.M VSS.t402 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X121 a_31732_10267# ITAIL.t17 RES_74k_1.P VDD.t534 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X122 a_29415_9553# mux_magic_1.OR_magic_0.B a_29415_8145# VDD.t306 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X123 a_27922_11758# mux_magic_0.AND2_magic_0.A a_27722_11758# VSS.t53 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X124 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT a_25706_n567# VSS.t83 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X125 VSS DIV_OUT.t1 a_20103_8443# VSS.t587 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X126 RES_74k_1.P RES_74k_1.P VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X127 VSS VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT VSS.t75 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X128 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t604 VDD.t575 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X129 VDD.t236 VDD.t235 VDD.t236 VDD.t206 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X130 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t722 VDD.t712 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X131 VSS VCTRL2.t9 a_25706_n567# VSS.t451 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X132 a_19897_11741# mux_magic_2.AND2_magic_0.A VDD.t655 VDD.t654 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X133 RES_74k_1.P RES_74k_1.P VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X134 VSS OUT.t14 OUTB.t11 VSS.t768 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X135 PFD_T2_0.FDIV a_21443_9476# VDD.t764 VDD.t20 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X136 RES_74k_1.P RES_74k_1.P VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X137 VDD.t234 VDD.t233 VDD.t234 VDD.t152 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X138 PFD_T2_0.INV_mag_1.IN a_22967_8787# VDD.t284 VDD.t283 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X139 a_25557_8739# PFD_T2_0.Buffer_V_2_0.IN VDD.t396 VDD.t395 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X140 VDD ITAIL.t12 ITAIL.t13 VDD.t538 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X141 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t603 VDD.t580 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X142 RES_74k_1.M VSS.t401 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X143 a_24436_11277# PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.IN VDD.t441 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X144 VSS VSS.t262 a_20103_9637# VSS.t263 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X145 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t602 VDD.t589 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X146 VDD A_MUX_0.Tr_Gate_1.CLK a_45158_5339# VDD.t298 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X147 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t324 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X148 mux_magic_0.OR_magic_0.B a_27722_10564# VSS.t147 VSS.t146 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X149 a_22880_9797# PFD_T2_0.INV_mag_0.OUT a_22967_8787# VSS.t138 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X150 a_45328_12082# a_45628_11460# VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X151 a_41879_1284# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD.t649 VDD.t263 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X152 a_44128_8770# a_43828_8148# VDD.t25 ppolyf_u r_width=1.1u r_length=2.6u
X153 mux_magic_1.AND2_magic_0.A S3.t3 VDD.t801 VDD.t800 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X154 VDD.t232 VDD.t230 VDD.t232 VDD.t231 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X155 VDD S2.t2 a_27722_10564# VDD.t420 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X156 RES_74k_1.P ITAIL.t18 a_31732_10267# VDD.t539 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X157 VSS VCTRL2.t10 a_25706_n567# VSS.t517 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X158 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VSS.t676 VSS.t675 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X159 RES_74k_1.M VSS.t400 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X160 mux_magic_0.OR_magic_0.A a_27722_11758# VSS.t95 VSS.t94 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X161 RES_74k_1.M VSS.t399 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X162 VDD a_31468_10271# a_31732_10267# VDD.t122 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X163 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VDD.t332 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X164 RES_74k_1.M VSS.t398 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X165 a_31468_10271# DN.t3 VDD.t666 VDD.t104 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X166 a_45628_11254# a_45328_10632# VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X167 VDD A_MUX_0.Tr_Gate_1.CLK a_45158_5339# VDD.t295 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X168 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT a_34443_2598# VSS.t91 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X169 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VSS.t478 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X170 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_41879_1284# VDD.t261 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X171 a_22880_9797# PFD_T2_0.INV_mag_1.OUT VSS.t15 VSS.t14 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X172 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t705 VDD.t683 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X173 VDD OUT.t15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD.t48 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X174 VDD.t229 VDD.t228 VDD.t229 VDD.t182 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X175 VDD a_22966_11778# PFD_T2_0.INV_mag_0.IN VDD.t752 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X176 RES_74k_1.P RES_74k_1.P VDD.t25 ppolyf_u r_width=1.1u r_length=2.6u
X177 a_34443_2598# VCTRL2.t11 VSS.t547 VSS.t533 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X178 VSS VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VSS.t672 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X179 a_20097_10547# F_IN.t0 VSS.t734 VSS.t733 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X180 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t352 VDD.t327 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X181 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t517 VDD.t483 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X182 RES_74k_1.M VSS.t397 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X183 a_22880_10947# a_22966_11778# VSS.t706 VSS.t705 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X184 VSS UP.t5 a_31940_9626# VSS.t122 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X185 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD.t562 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X186 mux_magic_3.OR_magic_0.A a_19903_8443# VDD.t759 VDD.t758 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X187 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t324 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X188 RES_74k_1.M VSS.t396 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X189 a_21443_9476# mux_magic_3.OR_magic_0.B a_21443_8068# VDD.t22 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X190 RES_74k_1.M VSS.t395 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X191 VDD VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD.t461 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X192 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VSS.t621 VSS.t620 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X193 VDD a_31468_10271# a_31732_10267# VDD.t122 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X194 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD.t714 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X195 a_22880_10947# PFD_T2_0.FIN PFD_T2_0.INV_mag_0.IN VSS.t138 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X196 a_22967_8787# PFD_T2_0.FDIV VDD.t376 VDD.t283 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X197 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VSS.t755 VSS.t754 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X198 RES_74k_1.M VSS.t394 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X199 VDD mux_magic_2.OR_magic_0.A a_21437_12116# VDD.t17 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X200 RES_74k_1.M VSS.t393 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X201 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUT.t7 VDD.t31 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X202 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB VDD.t470 VDD.t459 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X203 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.OUTB VDD.t816 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X204 RES_74k_1.M VSS.t392 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X205 a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD.t646 VDD.t372 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X206 VSS VCTRL2.t12 a_25706_n567# VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X207 VDD.t227 VDD.t225 VDD.t227 VDD.t226 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X208 RES_74k_1.P RES_74k_1.P VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X209 VSS VCTRL2.t13 a_25706_n567# VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X210 RES_74k_1.P RES_74k_1.P VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X211 a_45158_5339# A_MUX_0.Tr_Gate_1.CLK VSS.t111 VSS.t107 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X212 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t591 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X213 a_42763_5679# S4.t2 VDD.t90 VDD.t77 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X214 UP a_29262_10725# VDD.t24 VDD.t3 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X215 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t329 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X216 mux_magic_2.OR_magic_0.A a_19897_11741# VSS.t59 VSS.t58 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X217 VSS a_22967_8787# a_22881_9554# VSS.t103 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X218 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t599 VDD.t598 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X219 RES_74k_1.M VSS.t391 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X220 a_20097_10547# S1.t1 a_19897_10547# VSS.t593 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X221 VDD a_25557_8739# PFD_T2_0.DOWN VDD.t66 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X222 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t514 VDD.t508 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X223 RES_74k_1.M a_42628_11460# VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X224 VDD OUT.t16 OUTB.t7 VDD.t45 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X225 mux_magic_0.AND2_magic_0.A S2.t3 VDD.t121 VDD.t120 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X226 a_46528_12082# a_46228_11460# VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X227 VSS.t261 VSS.t260 VSS.t261 VSS.t181 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X228 a_19903_9637# S6.t2 VDD.t400 VDD.t399 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X229 PFD_T2_0.INV_mag_0.IN a_22966_11778# VDD.t751 VDD.t439 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X230 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VSS.t501 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X231 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD.t638 VDD.t445 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X232 a_45328_10426# a_45628_9804# VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X233 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD.t144 VDD.t131 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X234 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t702 VDD.t575 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X235 RES_74k_1.P RES_74k_1.P VDD.t69 ppolyf_u r_width=1.1u r_length=2.6u
X236 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN VDD.t440 VDD.t439 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X237 VDD a_22967_8787# PFD_T2_0.INV_mag_1.IN VDD.t280 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X238 DN a_29415_9553# VDD.t476 VDD.t474 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X239 a_43828_9598# a_43528_8976# VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X240 VCO_DFF_C_0.VCTRL S4.t3 VCTRL_IN.t7 VSS.t57 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X241 VCTRL_IN a_42763_5679# VCO_DFF_C_0.VCTRL VDD.t78 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X242 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VSS.t92 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X243 VSS VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VSS.t669 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X244 RES_74k_1.M VSS.t390 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X245 mux_magic_2.AND2_magic_0.A S1.t2 VDD.t524 VDD.t523 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X246 a_42628_11254# a_42628_10426# VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X247 a_46228_11254# a_46528_10632# VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X248 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t567 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X249 RES_74k_1.M VSS.t389 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X250 a_21437_10708# mux_magic_2.OR_magic_0.B a_21437_12116# VDD.t548 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X251 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT a_34443_2598# VSS.t91 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X252 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t699 VDD.t565 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X253 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VSS.t646 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X254 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_0.OUT VSS.t700 VSS.t14 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X255 VDD DIV_OUT.t2 a_19903_8443# VDD.t301 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X256 VDD mux_magic_1.OR_magic_0.A a_29415_8145# VDD.t308 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X257 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t347 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X258 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD.t143 VDD.t139 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X259 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VSS.t132 VSS.t131 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X260 RES_74k_1.M VSS.t388 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X261 RES_74k_1.M VSS.t387 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X262 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB a_25706_n567# VSS.t83 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X263 mux_magic_0.OR_magic_0.A a_27722_11758# VDD.t254 VDD.t253 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X264 a_23837_9553# PFD_T2_0.INV_mag_1.IN PFD_T2_0.Buffer_V_2_0.IN VSS.t420 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X265 a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD.t645 VDD.t371 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X266 a_25706_n567# VCTRL2.t14 VSS.t552 VSS.t504 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X267 RES_74k_1.P RES_74k_1.P VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X268 VSS.t259 VSS.t257 VSS.t259 VSS.t258 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X269 RES_74k_1.M VSS.t386 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X270 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD.t692 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X271 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD.t371 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X272 VSS ITAIL1.t4 ITAIL1.t5 VSS.t43 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X273 a_45028_9598# a_45328_8976# VDD.t57 ppolyf_u r_width=1.1u r_length=2.6u
X274 a_34443_2598# VCTRL2.t15 VSS.t553 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X275 VSS VCTRL2.t16 a_34443_2598# VSS.t434 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X276 a_28075_8520# PFD_T2_0.DOWN VSS.t29 VSS.t28 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X277 RES_74k_1.P RES_74k_1.P VDD.t63 ppolyf_u r_width=1.1u r_length=2.6u
X278 RES_74k_1.P a_45158_5339# VCO_DFF_C_0.VCTRL VDD.t298 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X279 a_25706_n567# VCTRL2.t17 VSS.t556 VSS.t442 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X280 a_24436_11277# PFD_T2_0.INV_mag_1.IN VDD.t416 VDD.t415 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X281 VSS VCTRL2.t18 a_34443_2598# VSS.t155 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X282 VDD F_IN.t1 a_19897_10547# VDD.t790 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X283 RES_74k_1.P ITAIL.t19 a_31732_10267# VDD.t537 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X284 VDD PFD_T2_0.FDIV a_22967_8787# VDD.t280 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X285 a_46528_8770# RES_74k_1.P VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X286 mux_magic_0.AND2_magic_0.A S2.t4 VDD.t760 VDD.t608 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X287 a_43528_8770# a_43228_8148# VDD.t63 ppolyf_u r_width=1.1u r_length=2.6u
X288 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t347 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X289 a_28075_9714# DN_INPUT.t1 VSS.t97 VSS.t96 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X290 VDD S4.t4 A_MUX_0.Tr_Gate_1.CLK VDD.t85 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X291 VDD VCO_DFF_C_0.VCO_C_0.OUTB a_44716_1837# VDD.t373 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X292 VDD.t224 VDD.t223 VDD.t224 VDD.t197 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X293 a_25706_n567# VCTRL2.t19 VSS.t559 VSS.t148 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X294 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.OUT VSS.t13 VSS.t11 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X295 a_29262_10725# mux_magic_0.OR_magic_0.B VSS.t1 VSS.t0 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X296 a_43528_12082# a_43228_11460# VDD.t63 ppolyf_u r_width=1.1u r_length=2.6u
X297 RES_74k_1.P a_45158_5339# VCO_DFF_C_0.VCTRL VDD.t295 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X298 VSS.t256 VSS.t254 VSS.t256 VSS.t255 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X299 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT a_34443_2598# VSS.t88 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X300 a_34443_2598# VCTRL2.t20 VSS.t560 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X301 RES_74k_1.P RES_74k_1.P VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X302 VSS VCTRL2.t21 a_34443_2598# VSS.t155 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X303 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t591 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X304 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN a_23836_10693# VSS.t468 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X305 ITAIL1 ITAIL1.t2 VSS.t42 VSS.t41 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X306 mux_magic_1.AND2_magic_0.A S3.t4 VDD.t803 VDD.t802 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X307 RES_74k_1.P RES_74k_1.P VDD.t63 ppolyf_u r_width=1.1u r_length=2.6u
X308 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_n196# VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD.t263 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X309 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t572 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X310 VDD mux_magic_3.OR_magic_0.A a_21443_8068# VDD.t783 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X311 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK VCO_DFF_C_0.VCTRL VSS.t106 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X312 RES_74k_1.M VSS.t385 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X313 VSS.t253 VSS.t252 VSS.t253 VSS.t175 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X314 VSS S4.t5 A_MUX_0.Tr_Gate_1.CLK VSS.t62 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X315 mux_magic_2.AND2_magic_0.A S1.t3 VDD.t526 VDD.t525 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X316 a_43228_11254# a_43528_10632# VDD.t63 ppolyf_u r_width=1.1u r_length=2.6u
X317 RES_74k_1.M VSS.t384 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X318 VSS PFD_T2_0.INV_mag_1.IN a_23837_9553# VSS.t416 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X319 a_44728_8770# a_45028_8148# VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X320 a_22879_10704# PFD_T2_0.INV_mag_0.OUT a_22966_11778# VSS.t699 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X321 a_28075_8520# mux_magic_1.AND2_magic_0.A a_27875_8520# VSS.t142 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X322 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_44716_n517# VDD.t370 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X323 a_27922_10564# UP_INPUT.t0 VSS.t666 VSS.t665 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X324 RES_74k_1.M VSS.t383 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X325 VSS.t251 VSS.t250 VSS.t251 VSS.t178 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X326 VDD S4.t6 A_MUX_0.Tr_Gate_1.CLK VDD.t106 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X327 RES_74k_1.M VSS.t382 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X328 VDD mux_magic_2.AND2_magic_0.A a_19897_11741# VDD.t651 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X329 a_28075_9714# S3.t5 a_27875_9714# VSS.t743 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X330 VCO_DFF_C_0.VCTRL a_42763_5679# VCTRL_IN.t2 VDD.t77 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X331 VDD.t222 VDD.t220 VDD.t222 VDD.t221 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X332 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t152 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X333 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t591 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X334 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VSS.t491 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X335 VDD mux_magic_0.OR_magic_0.A a_29262_12133# VDD.t477 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X336 a_27922_11758# PFD_T2_0.UP VSS.t763 VSS.t762 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X337 RES_74k_1.P RES_74k_1.P VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X338 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t696 VDD.t668 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X339 RES_74k_1.M VSS.t381 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X340 VSS PFD_T2_0.DOWN a_28075_8520# VSS.t25 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X341 a_29262_10725# mux_magic_0.OR_magic_0.B a_29262_12133# VDD.t1 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X342 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD.t370 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X343 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT a_34443_2598# VSS.t90 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X344 VSS VCTRL2.t22 a_25706_n567# VSS.t457 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X345 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t695 VDD.t580 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X346 a_31468_10271# DN.t4 VDD.t105 VDD.t104 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X347 VDD.t219 VDD.t217 VDD.t219 VDD.t218 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X348 RES_74k_1.M VSS.t380 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X349 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VSS.t488 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X350 a_31468_10271# DN.t5 VSS.t634 VSS.t633 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X351 RES_74k_1.P RES_74k_1.P VDD.t55 ppolyf_u r_width=1.1u r_length=2.6u
X352 VSS VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VSS.t128 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X353 mux_magic_3.AND2_magic_0.A S6.t3 VSS.t173 VSS.t172 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X354 RES_74k_1.M VSS.t379 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X355 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT a_25706_n567# VSS.t83 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X356 ITAIL ITAIL.t10 VDD.t555 VDD.t539 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X357 VSS DN_INPUT.t2 a_28075_9714# VSS.t98 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X358 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD.t692 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X359 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_41879_1284# VSS.t650 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X360 PFD_T2_0.INV_mag_0.IN a_22966_11778# VDD.t750 VDD.t437 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X361 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t511 VDD.t322 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X362 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t590 VDD.t589 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X363 a_29415_9553# mux_magic_1.OR_magic_0.B a_29415_8145# VDD.t306 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X364 a_34443_2598# VCTRL2.t23 VSS.t565 VSS.t446 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X365 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VSS.t668 VSS.t667 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X366 PFD_T2_0.INV_mag_0.IN a_22966_11778# VDD.t749 VDD.t435 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X367 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN VDD.t438 VDD.t437 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X368 RES_74k_1.M VSS.t378 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X369 RES_74k_1.M VSS.t377 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X370 RES_74k_1.M VSS.t376 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X371 ITAIL1 ITAIL1.t0 VSS.t40 VSS.t39 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X372 VSS VCTRL2.t24 a_34443_2598# VSS.t448 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X373 a_41879_n196# VCO_DFF_C_0.VCO_C_0.OUTB VSS.t497 VSS.t496 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X374 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD.t823 VDD.t811 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X375 a_44128_12082# a_44428_11460# VDD.t55 ppolyf_u r_width=1.1u r_length=2.6u
X376 RES_74k_1.P VSS.t712 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X377 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t147 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X378 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN VDD.t436 VDD.t435 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X379 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB a_25706_n567# VSS.t83 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X380 VSS.t249 VSS.t248 VSS.t249 VSS.t237 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X381 RES_74k_1.M VSS.t375 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X382 VSS VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VSS.t493 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X383 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t567 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X384 VSS S2.t5 mux_magic_0.AND2_magic_0.A VSS.t715 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X385 mux_magic_1.OR_magic_0.A a_27875_8520# VDD.t386 VDD.t385 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X386 a_34443_2598# VCTRL2.t25 VSS.t568 VSS.t533 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X387 RES_74k_1.M VSS.t374 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X388 RES_74k_1.M VSS.t373 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X389 a_25706_n567# VCTRL2.t26 VSS.t569 VSS.t158 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X390 VSS mux_magic_2.OR_magic_0.A a_21437_10708# VSS.t18 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X391 VSS.t247 VSS.t245 VSS.t247 VSS.t246 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X392 a_44716_1837# VCO_DFF_C_0.VCO_C_0.OUTB VDD.t467 VDD.t372 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X393 RES_74k_1.M VSS.t372 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X394 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_44716_n517# VDD.t373 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X395 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_1284# OUTB.t14 VDD.t260 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X396 PFD_T2_0.UP a_25556_11637# VDD.t249 VDD.t248 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X397 a_44428_11254# a_44128_10632# VDD.t55 ppolyf_u r_width=1.1u r_length=2.6u
X398 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL VDD.t173 VDD.t155 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X399 mux_magic_1.OR_magic_0.B a_27875_9714# VDD.t103 VDD.t102 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X400 a_46528_10426# a_46228_9804# VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X401 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t559 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X402 a_42928_10426# a_43228_9804# VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X403 VSS OUT.t17 OUTB.t10 VSS.t771 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X404 VDD.t216 VDD.t215 VDD.t216 VDD.t147 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X405 a_25556_11637# PFD_T2_0.Buffer_V_2_1.IN VDD.t769 VDD.t768 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X406 a_44428_9598# a_44728_8976# VDD.t54 ppolyf_u r_width=1.1u r_length=2.6u
X407 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT a_41879_n196# VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD.t262 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X408 PFD_T2_0.DOWN a_25557_8739# VDD.t65 VDD.t64 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X409 RES_74k_1.M VSS.t371 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X410 RES_74k_1.M VSS.t370 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X411 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD.t707 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X412 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t510 VDD.t336 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X413 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t584 VDD.t565 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X414 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VSS.t645 VSS.t644 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X415 VSS VCTRL2.t27 a_25706_n567# VSS.t517 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X416 a_42928_8770# a_42628_8148# VDD.t93 ppolyf_u r_width=1.1u r_length=2.6u
X417 RES_74k_1.M VSS.t369 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X418 VSS F_IN.t2 a_20097_10547# VSS.t735 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X419 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD.t577 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X420 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t149 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X421 VDD ITAIL.t8 ITAIL.t9 VDD.t538 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X422 a_34443_2598# VCTRL2.t28 VSS.t573 VSS.t572 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X423 a_25706_n567# VCTRL2.t29 VSS.t505 VSS.t504 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X424 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD.t677 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X425 RES_74k_1.P RES_74k_1.P VDD.t57 ppolyf_u r_width=1.1u r_length=2.6u
X426 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT a_34443_2598# VSS.t90 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X427 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VDD.t317 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X428 RES_74k_1.M VSS.t368 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X429 mux_magic_2.OR_magic_0.A a_19897_11741# VDD.t98 VDD.t97 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X430 RES_74k_1.M VSS.t367 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X431 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_44716_1837# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD.t373 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X432 VDD mux_magic_0.AND2_magic_0.A a_27722_11758# VDD.t82 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X433 a_22879_10704# PFD_T2_0.INV_mag_1.OUT VSS.t12 VSS.t11 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X434 RES_74k_1.P RES_74k_1.P VDD.t93 ppolyf_u r_width=1.1u r_length=2.6u
X435 a_42763_5679# S4.t7 VSS.t66 VSS.t65 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X436 RES_74k_1.P VSS.t711 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X437 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN a_23836_10693# VSS.t475 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X438 a_46228_9598# a_45928_8976# VDD.t56 ppolyf_u r_width=1.1u r_length=2.6u
X439 RES_74k_1.M VSS.t366 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X440 a_29262_12133# mux_magic_0.OR_magic_0.B a_29262_10725# VDD.t3 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X441 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t344 VDD.t315 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X442 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t509 VDD.t508 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X443 a_45158_5339# A_MUX_0.Tr_Gate_1.CLK VDD.t294 VDD.t293 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X444 VSS.t244 VSS.t243 VSS.t244 VSS.t181 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X445 VSS.t242 VSS.t241 VSS.t242 VSS.t175 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X446 RES_74k_1.M VSS.t365 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X447 VDD OUT.t18 OUTB.t6 VDD.t31 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X448 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.OUTB VDD.t813 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X449 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN a_23837_9553# VSS.t417 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X450 VSS.t240 VSS.t239 VSS.t240 VSS.t221 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X451 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t19 VDD.t35 VDD.t34 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X452 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t581 VDD.t580 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X453 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VSS.t82 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X454 VDD S1.t4 mux_magic_2.AND2_magic_0.A VDD.t527 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X455 a_45328_12082# a_45028_11460# VDD.t57 ppolyf_u r_width=1.1u r_length=2.6u
X456 a_44128_8770# a_44428_8148# VDD.t55 ppolyf_u r_width=1.1u r_length=2.6u
X457 mux_magic_1.AND2_magic_0.A S3.t6 VSS.t745 VSS.t744 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X458 RES_74k_1.M VSS.t364 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X459 VSS.t238 VSS.t236 VSS.t238 VSS.t237 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X460 RES_74k_1.M VSS.t363 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X461 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t20 VDD.t37 VDD.t36 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X462 VDD OUT.t21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD.t38 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X463 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUT.t6 VDD.t45 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X464 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VSS.t617 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X465 mux_magic_3.OR_magic_0.B a_19903_9637# VDD.t734 VDD.t733 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X466 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD.t620 VDD.t43 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X467 PFD_T2_0.FIN a_21437_10708# VDD.t364 VDD.t363 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X468 VDD.t214 VDD.t212 VDD.t214 VDD.t213 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X469 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t155 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X470 a_45028_11254# a_45328_10632# VDD.t57 ppolyf_u r_width=1.1u r_length=2.6u
X471 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t343 VDD.t313 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X472 VDD VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD.t449 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X473 RES_74k_1.M VSS.t362 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X474 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VSS.t82 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X475 VSS.t235 VSS.t233 VSS.t235 VSS.t234 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X476 a_31940_9626# ITAIL1.t10 RES_74k_1.P VSS.t46 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X477 RES_74k_1.P RES_74k_1.P VDD.t55 ppolyf_u r_width=1.1u r_length=2.6u
X478 a_34443_2598# VCTRL2.t30 VSS.t506 VSS.t466 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X479 a_29415_8145# mux_magic_1.OR_magic_0.A VDD.t310 VDD.t308 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X480 VSS.t232 VSS.t231 VSS.t232 VSS.t175 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X481 a_25706_n567# VCTRL2.t31 VSS.t507 VSS.t504 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X482 RES_74k_1.P VSS.t710 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X483 RES_74k_1.M VSS.t361 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X484 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK OUTB.t19 VSS.t653 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X485 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t559 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X486 VSS A_MUX_0.Tr_Gate_1.CLK a_45158_5339# VSS.t108 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X487 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT a_34443_2598# VSS.t503 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X488 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB VDD.t464 VDD.t445 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X489 VDD a_22967_8787# PFD_T2_0.INV_mag_1.IN VDD.t277 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X490 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t717 VDD.t710 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X491 DN a_29415_9553# VDD.t475 VDD.t474 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X492 RES_74k_1.M VSS.t360 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X493 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t567 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X494 VSS VCTRL2.t32 a_34443_2598# VSS.t434 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X495 VDD a_19903_8443# mux_magic_3.OR_magic_0.A VDD.t755 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X496 mux_magic_3.AND2_magic_0.A S6.t4 VDD.t771 VDD.t770 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X497 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VDD.t501 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X498 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD.t637 VDD.t459 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X499 VDD a_19897_10547# mux_magic_2.OR_magic_0.B VDD.t540 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X500 OUTB OUT.t22 VDD.t42 VDD.t41 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X501 VDD UP_INPUT.t1 a_27722_10564# VDD.t663 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X502 RES_74k_1.M VSS.t359 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X503 RES_74k_1.M VSS.t358 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X504 VDD a_22967_8787# PFD_T2_0.INV_mag_1.IN VDD.t274 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X505 PFD_T2_0.INV_mag_0.IN a_22966_11778# VDD.t748 VDD.t368 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X506 RES_74k_1.P RES_74k_1.P VDD.t69 ppolyf_u r_width=1.1u r_length=2.6u
X507 RES_74k_1.P RES_74k_1.P VDD.t56 ppolyf_u r_width=1.1u r_length=2.6u
X508 OUTB OUT.t23 VDD.t44 VDD.t43 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X509 a_20103_8443# mux_magic_3.AND2_magic_0.A a_19903_8443# VSS.t52 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X510 VSS.t230 VSS.t228 VSS.t230 VSS.t229 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X511 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t685 VDD.t565 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X512 VSS VCTRL2.t33 a_25706_n567# VSS.t457 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X513 a_22966_11778# PFD_T2_0.FIN VDD.t369 VDD.t368 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X514 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t329 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X515 VSS VCTRL2.t34 a_34443_2598# VSS.t428 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X516 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCTRL VDD.t168 VDD.t149 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X517 a_20097_11741# PRE_SCALAR.t1 VSS.t688 VSS.t687 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X518 VSS.t227 VSS.t225 VSS.t227 VSS.t226 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X519 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VSS.t682 VSS.t644 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X520 a_20103_9637# S6.t5 a_19903_9637# VSS.t722 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X521 RES_74k_1.P RES_74k_1.P VDD.t69 ppolyf_u r_width=1.1u r_length=2.6u
X522 VCTRL_IN S4.t8 VCO_DFF_C_0.VCTRL VSS.t67 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X523 VDD.t211 VDD.t210 VDD.t211 VDD.t206 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X524 VSS.t224 VSS.t223 VSS.t224 VSS.t178 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X525 VSS PFD_T2_0.INV_mag_0.OUT PFD_T2_0.Buffer_V_2_0.IN VSS.t696 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X526 a_45928_12082# a_46228_11460# VDD.t56 ppolyf_u r_width=1.1u r_length=2.6u
X527 VSS.t222 VSS.t220 VSS.t222 VSS.t221 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X528 VSS VCTRL2.t35 a_34443_2598# VSS.t514 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X529 a_27722_10564# S2.t6 VDD.t762 VDD.t761 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X530 VDD VSS.t775 a_19903_9637# VDD.t836 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X531 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VSS.t482 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X532 VSS VCTRL2.t36 a_25706_n567# VSS.t517 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X533 VDD PFD_T2_0.INV_mag_1.IN PFD_T2_0.Buffer_V_2_0.IN VDD.t277 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X534 a_45928_10426# a_45628_9804# VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X535 a_25706_n567# VCTRL2.t37 VSS.t520 VSS.t148 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X536 RES_74k_1.M VSS.t357 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X537 VSS.t219 VSS.t217 VSS.t219 VSS.t218 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X538 a_21437_10708# mux_magic_2.OR_magic_0.B a_21437_12116# VDD.t547 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X539 a_42628_10426# a_42628_9804# VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X540 VSS VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VSS.t128 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X541 RES_74k_1.M VSS.t356 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X542 RES_74k_1.M VSS.t355 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X543 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_1837# VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t372 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X544 mux_magic_0.AND2_magic_0.A S2.t7 VDD.t607 VDD.t120 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X545 a_21443_8068# mux_magic_3.OR_magic_0.A VDD.t784 VDD.t783 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X546 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VSS.t641 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X547 VSS mux_magic_0.OR_magic_0.A a_29262_10725# VSS.t578 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X548 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VSS.t629 VSS.t30 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X549 PFD_T2_0.DOWN a_25557_8739# VSS.t50 VSS.t49 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X550 RES_74k_1.P RES_74k_1.P VDD.t69 ppolyf_u r_width=1.1u r_length=2.6u
X551 a_46228_11254# a_45928_10632# VDD.t56 ppolyf_u r_width=1.1u r_length=2.6u
X552 RES_74k_1.M VSS.t354 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X553 RES_74k_1.M VSS.t353 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X554 VSS.t216 VSS.t215 VSS.t216 VSS.t178 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X555 VSS.t214 VSS.t213 VSS.t214 VSS.t209 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X556 a_21437_10708# mux_magic_2.OR_magic_0.B a_21437_12116# VDD.t546 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X557 VDD a_31468_10271# a_31732_10267# VDD.t122 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X558 VDD PFD_T2_0.INV_mag_1.IN PFD_T2_0.Buffer_V_2_0.IN VDD.t274 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X559 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VSS.t89 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X560 VSS.t212 VSS.t211 VSS.t212 VSS.t184 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X561 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB a_25706_n567# VSS.t81 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X562 VDD PFD_T2_0.INV_mag_0.IN a_24437_9224# VDD.t432 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X563 VSS.t210 VSS.t208 VSS.t210 VSS.t209 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X564 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t684 VDD.t683 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X565 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VSS.t80 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X566 VDD S4.t9 A_MUX_0.Tr_Gate_1.CLK VDD.t106 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X567 VDD S6.t6 mux_magic_3.AND2_magic_0.A VDD.t772 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X568 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t682 VDD.t598 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X569 a_20097_11741# mux_magic_2.AND2_magic_0.A a_19897_11741# VSS.t661 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X570 a_31732_10267# ITAIL.t21 RES_74k_1.P VDD.t534 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X571 VDD PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.OUT VDD.t408 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X572 RES_74k_1.M VSS.t352 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X573 RES_74k_1.M VSS.t351 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X574 mux_magic_1.AND2_magic_0.A S3.t7 VDD.t804 VDD.t802 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X575 RES_74k_1.M VSS.t350 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X576 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL VDD.t167 VDD.t155 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X577 VDD a_27722_10564# mux_magic_0.OR_magic_0.B VDD.t389 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X578 RES_74k_1.P ITAIL.t22 a_31732_10267# VDD.t537 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X579 RES_74k_1.M VSS.t349 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X580 PFD_T2_0.INV_mag_1.IN a_22967_8787# VDD.t273 VDD.t272 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X581 a_44128_10426# a_43828_9804# VDD.t25 ppolyf_u r_width=1.1u r_length=2.6u
X582 a_45628_9598# a_45328_8976# VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X583 RES_74k_1.P RES_74k_1.P VDD.t69 ppolyf_u r_width=1.1u r_length=2.6u
X584 RES_74k_1.M VSS.t348 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X585 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT a_25706_n567# VSS.t81 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X586 VCO_DFF_C_0.VCTRL a_45158_5339# RES_74k_1.P VDD.t293 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X587 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VSS.t86 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X588 RES_74k_1.M VSS.t347 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X589 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VSS.t80 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X590 PFD_T2_0.UP a_25556_11637# VSS.t85 VSS.t84 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X591 PFD_T2_0.INV_mag_1.IN a_22967_8787# VDD.t271 VDD.t270 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X592 RES_74k_1.P RES_74k_1.P VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X593 a_34443_2598# VCTRL2.t38 VSS.t521 VSS.t446 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X594 RES_74k_1.P RES_74k_1.P VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X595 VSS S4.t10 A_MUX_0.Tr_Gate_1.CLK VSS.t62 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X596 a_44716_1837# VCO_DFF_C_0.VCO_C_0.OUTB VSS.t492 VSS.t491 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X597 a_43528_8770# a_43828_8148# VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X598 VSS VCTRL2.t39 a_34443_2598# VSS.t448 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X599 RES_74k_1.M VSS.t346 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X600 VDD a_31468_10271# a_31732_10267# VDD.t122 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X601 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VSS.t502 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X602 a_29262_12133# mux_magic_0.OR_magic_0.A VDD.t478 VDD.t477 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X603 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t505 VDD.t320 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X604 PFD_T2_0.INV_mag_0.IN a_22966_11778# VDD.t747 VDD.t746 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X605 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t572 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X606 a_23837_9553# PFD_T2_0.INV_mag_1.IN VSS.t421 VSS.t420 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X607 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t338 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X608 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD.t636 VDD.t445 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X609 mux_magic_0.AND2_magic_0.A S2.t8 VDD.t609 VDD.t608 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X610 a_42928_12082# a_43228_11460# VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X611 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t152 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X612 RES_74k_1.M VSS.t345 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X613 VSS UP.t6 a_31940_9626# VSS.t122 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X614 RES_74k_1.P RES_74k_1.P VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X615 a_19903_8443# DIV_OUT.t3 VDD.t305 VDD.t304 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X616 RES_74k_1.P RES_74k_1.P VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X617 RES_74k_1.M VSS.t344 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X618 RES_74k_1.P RES_74k_1.P VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X619 A_MUX_0.Tr_Gate_1.CLK S4.t11 VDD.t112 VDD.t111 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X620 RES_74k_1.M VSS.t343 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X621 a_25706_n567# VCTRL2.t40 VSS.t524 VSS.t158 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X622 RES_74k_1.M VSS.t342 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X623 RES_74k_1.M VSS.t341 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X624 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t504 VDD.t336 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X625 VSS VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VSS.t125 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X626 a_34443_2598# VCTRL2.t41 VSS.t526 VSS.t525 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X627 a_25706_n567# VCTRL2.t42 VSS.t527 VSS.t504 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X628 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t24 VSS.t31 VSS.t30 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X629 a_43228_11254# a_42928_10632# VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X630 RES_74k_1.P RES_74k_1.P VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X631 a_45328_8770# a_45028_8148# VDD.t57 ppolyf_u r_width=1.1u r_length=2.6u
X632 VSS VCTRL2.t43 a_34443_2598# VSS.t528 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X633 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VSS.t640 VSS.t639 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X634 VSS VCTRL2.t44 a_25706_n567# VSS.t517 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X635 a_31732_10267# ITAIL.t23 RES_74k_1.P VDD.t538 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X636 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN VDD.t407 VDD.t270 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X637 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VSS.t89 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X638 a_24437_9224# PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.IN VDD.t406 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X639 A_MUX_0.Tr_Gate_1.CLK S4.t12 VDD.t114 VDD.t113 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X640 RES_74k_1.M VSS.t340 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X641 mux_magic_2.AND2_magic_0.A S1.t5 VDD.t531 VDD.t530 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X642 a_31468_10271# DN.t6 VDD.t625 VDD.t104 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X643 UP a_29262_10725# VSS.t24 VSS.t23 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X644 RES_74k_1.P RES_74k_1.P VDD.t57 ppolyf_u r_width=1.1u r_length=2.6u
X645 RES_74k_1.M VSS.t339 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X646 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD.t577 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X647 RES_74k_1.M VSS.t338 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X648 VSS VCO_DFF_C_0.VCO_C_0.OUTB a_41879_n196# VSS.t488 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X649 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VSS.t641 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X650 VSS VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VSS.t485 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X651 VDD S3.t8 mux_magic_1.AND2_magic_0.A VDD.t805 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X652 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t337 VDD.t336 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X653 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL VDD.t164 VDD.t155 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X654 RES_74k_1.P RES_74k_1.P VDD.t25 ppolyf_u r_width=1.1u r_length=2.6u
X655 VSS.t207 VSS.t206 VSS.t207 VSS.t181 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X656 VSS.t205 VSS.t204 VSS.t205 VSS.t175 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X657 a_34443_2598# VCTRL2.t45 VSS.t534 VSS.t533 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X658 RES_74k_1.M VSS.t337 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X659 a_23836_10693# PFD_T2_0.INV_mag_0.IN VSS.t474 VSS.t471 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X660 RES_74k_1.M VSS.t336 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X661 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VSS.t648 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X662 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t335 VDD.t322 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X663 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT a_41879_n196# VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD.t261 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X664 VDD mux_magic_3.AND2_magic_0.A a_19903_8443# VDD.t72 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X665 a_42763_5679# S4.t13 VDD.t115 VDD.t76 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X666 mux_magic_2.AND2_magic_0.A S1.t6 VSS.t595 VSS.t594 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X667 a_44128_12082# a_43828_11460# VDD.t25 ppolyf_u r_width=1.1u r_length=2.6u
X668 VSS VCTRL2.t46 a_25706_n567# VSS.t451 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X669 RES_74k_1.M VSS.t335 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X670 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD.t714 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X671 OUTB OUT.t25 VSS.t33 VSS.t32 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X672 VDD PRE_SCALAR.t2 a_19897_11741# VDD.t727 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X673 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VSS.t501 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X674 PFD_T2_0.INV_mag_1.IN PFD_T2_0.FDIV a_22881_9554# VSS.t140 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X675 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK OUTB.t18 VSS.t652 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X676 a_34443_2598# VCTRL2.t47 VSS.t537 VSS.t533 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X677 a_29262_10725# mux_magic_0.OR_magic_0.B a_29262_12133# VDD.t2 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X678 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCTRL VDD.t163 VDD.t152 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X679 a_34443_2598# VCTRL2.t48 VSS.t538 VSS.t466 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X680 UP a_29262_10725# VDD.t23 VDD.t3 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X681 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.IN a_24436_11277# VDD.t431 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X682 a_29415_9553# mux_magic_1.OR_magic_0.B VSS.t575 VSS.t574 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X683 RES_74k_1.M VSS.t334 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X684 OUTB OUT.t26 VSS.t35 VSS.t34 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X685 VDD a_27875_8520# mux_magic_1.OR_magic_0.A VDD.t382 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X686 RES_74k_1.M VSS.t333 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X687 VSS.t203 VSS.t201 VSS.t203 VSS.t202 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X688 RES_74k_1.M VSS.t332 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X689 VDD PFD_T2_0.INV_mag_1.IN a_24436_11277# VDD.t403 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X690 a_43828_11254# a_44128_10632# VDD.t25 ppolyf_u r_width=1.1u r_length=2.6u
X691 a_46528_10426# a_46828_9598# VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X692 PFD_T2_0.FDIV a_21443_9476# VSS.t719 VSS.t718 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X693 a_43528_10426# a_43228_9804# VDD.t63 ppolyf_u r_width=1.1u r_length=2.6u
X694 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VSS.t82 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X695 VDD a_27875_9714# mux_magic_1.OR_magic_0.B VDD.t99 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X696 a_45158_5339# A_MUX_0.Tr_Gate_1.CLK VDD.t292 VDD.t291 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X697 PFD_T2_0.FDIV a_21443_9476# VDD.t763 VDD.t20 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X698 VDD OUT.t27 OUTB.t3 VDD.t45 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X699 VSS PFD_T2_0.INV_mag_1.OUT a_22880_9797# VSS.t8 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X700 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VDD.t332 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X701 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VDD.t501 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X702 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t329 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X703 VDD.t209 VDD.t208 VDD.t209 VDD.t188 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X704 RES_74k_1.M VSS.t331 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X705 VSS VCTRL2.t49 a_25706_n567# VSS.t457 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X706 a_29415_8145# mux_magic_1.OR_magic_0.A VDD.t309 VDD.t308 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X707 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD.t820 VDD.t819 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X708 a_34443_2598# VCTRL2.t50 VSS.t427 VSS.t426 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X709 VDD OUT.t28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD.t48 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X710 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t449 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X711 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t328 VDD.t327 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X712 VSS VCTRL2.t51 a_34443_2598# VSS.t428 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X713 a_25706_n567# VCTRL2.t52 VSS.t431 VSS.t148 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X714 RES_74k_1.P ITAIL1.t11 a_31940_9626# VSS.t41 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X715 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t576 VDD.t575 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X716 RES_74k_1.P RES_74k_1.P VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X717 VDD.t207 VDD.t205 VDD.t207 VDD.t206 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X718 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VSS.t479 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X719 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD.t677 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X720 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VSS.t679 VSS.t639 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X721 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD.t619 VDD.t41 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X722 VDD VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD.t461 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X723 PFD_T2_0.INV_mag_0.IN a_22966_11778# VDD.t745 VDD.t744 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X724 a_44728_10426# a_45028_9804# VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X725 VSS VCTRL2.t53 a_25706_n567# VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X726 RES_74k_1.M VSS.t330 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X727 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT a_25706_n567# VSS.t81 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X728 VDD PFD_T2_0.DOWN a_27875_8520# VDD.t28 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X729 a_46228_9598# a_46528_8976# VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X730 RES_74k_1.M VSS.t329 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X731 a_31940_9626# UP.t7 VSS.t121 VSS.t120 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X732 a_43228_9598# a_42928_8976# VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X733 a_27722_10564# UP_INPUT.t2 VDD.t789 VDD.t788 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X734 VDD ITAIL.t6 ITAIL.t7 VDD.t534 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X735 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t324 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X736 RES_74k_1.M VSS.t328 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X737 VDD S2.t9 mux_magic_0.AND2_magic_0.A VDD.t610 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X738 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD.t618 VDD.t43 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X739 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB VDD.t460 VDD.t459 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X740 a_21443_9476# mux_magic_3.OR_magic_0.B VSS.t22 VSS.t21 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X741 mux_magic_3.AND2_magic_0.A S6.t7 VDD.t775 VDD.t770 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X742 VDD S4.t14 a_42763_5679# VDD.t75 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X743 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t713 VDD.t712 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X744 a_44728_12082# a_45028_11460# VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X745 VSS.t200 VSS.t198 VSS.t200 VSS.t199 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X746 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VSS.t636 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X747 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.OUTB VSS.t751 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X748 VDD DN_INPUT.t3 a_27875_9714# VDD.t257 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X749 a_44728_8770# a_44428_8148# VDD.t54 ppolyf_u r_width=1.1u r_length=2.6u
X750 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t329 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X751 RES_74k_1.M VSS.t327 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X752 RES_74k_1.M VSS.t326 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X753 a_21443_9476# mux_magic_3.OR_magic_0.B a_21443_8068# VDD.t22 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X754 VSS.t197 VSS.t195 VSS.t197 VSS.t196 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X755 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VDD.t487 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X756 a_19897_10547# S1.t7 a_20097_10547# VSS.t596 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X757 a_31468_10271# DN.t7 VSS.t635 VSS.t633 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X758 VSS VCTRL2.t54 a_34443_2598# VSS.t434 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X759 VDD S1.t8 mux_magic_2.AND2_magic_0.A VDD.t527 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X760 VSS PRE_SCALAR.t3 a_20097_11741# VSS.t689 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X761 PFD_T2_0.FIN a_21437_10708# VDD.t362 VDD.t361 pfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X762 ITAIL ITAIL.t4 VDD.t550 VDD.t537 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X763 VSS VCTRL2.t55 a_34443_2598# VSS.t437 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X764 VDD.t204 VDD.t202 VDD.t204 VDD.t203 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X765 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VSS.t80 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X766 a_21437_12116# mux_magic_2.OR_magic_0.A VDD.t16 VDD.t15 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X767 VDD a_19903_9637# mux_magic_3.OR_magic_0.B VDD.t730 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X768 RES_74k_1.M VSS.t325 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X769 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t449 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X770 a_45028_11254# a_44728_10632# VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X771 RES_74k_1.P RES_74k_1.P VDD.t54 ppolyf_u r_width=1.1u r_length=2.6u
X772 VDD.t201 VDD.t199 VDD.t201 VDD.t200 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X773 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t496 VDD.t313 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X774 RES_74k_1.M VSS.t324 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X775 VSS VCO_DFF_C_0.VCO_C_0.OUTB a_44716_1837# VSS.t482 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X776 VDD PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.OUT VDD.t408 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X777 VSS.t194 VSS.t192 VSS.t194 VSS.t193 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X778 VSS.t191 VSS.t189 VSS.t191 VSS.t190 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X779 a_21437_12116# mux_magic_2.OR_magic_0.A VDD.t14 VDD.t13 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X780 VDD PFD_T2_0.UP a_27722_11758# VDD.t829 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X781 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.IN VSS.t473 VSS.t472 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.5u
X782 a_22881_9554# PFD_T2_0.FDIV PFD_T2_0.INV_mag_1.IN VSS.t139 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X783 PFD_T2_0.INV_mag_1.IN a_22967_8787# VDD.t269 VDD.t268 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X784 VDD a_22966_11778# PFD_T2_0.INV_mag_0.IN VDD.t426 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X785 VSS VCTRL2.t56 a_34443_2598# VSS.t434 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X786 VDD PFD_T2_0.INV_mag_0.IN PFD_T2_0.Buffer_V_2_1.IN VDD.t426 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X787 VSS PFD_T2_0.INV_mag_1.IN a_23837_9553# VSS.t417 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X788 RES_74k_1.M VSS.t323 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X789 VDD a_22966_11778# PFD_T2_0.INV_mag_0.IN VDD.t365 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X790 a_45928_8770# a_46228_8148# VDD.t56 ppolyf_u r_width=1.1u r_length=2.6u
X791 RES_74k_1.M VSS.t322 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X792 VSS PFD_T2_0.INV_mag_0.OUT PFD_T2_0.Buffer_V_2_0.IN VSS.t8 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X793 a_25706_n567# VCTRL2.t57 VSS.t443 VSS.t442 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X794 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT VDD.t136 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X795 VDD PFD_T2_0.FIN a_22966_11778# VDD.t365 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X796 ITAIL ITAIL.t2 VDD.t549 VDD.t539 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X797 VSS VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VSS.t125 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X798 a_19897_10547# F_IN.t3 VDD.t794 VDD.t793 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X799 DN a_29415_9553# VSS.t577 VSS.t576 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X800 VCO_DFF_C_0.VCTRL a_42763_5679# VCTRL_IN.t1 VDD.t76 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X801 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t591 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X802 RES_74k_1.M VSS.t321 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X803 a_27722_11758# mux_magic_0.AND2_magic_0.A VDD.t81 VDD.t80 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X804 RES_74k_1.P RES_74k_1.P VDD.t56 ppolyf_u r_width=1.1u r_length=2.6u
X805 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD.t631 VDD.t459 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X806 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.OUTB VDD.t816 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X807 VDD PFD_T2_0.Buffer_V_2_1.IN a_25556_11637# VDD.t765 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X808 a_19903_8443# mux_magic_3.AND2_magic_0.A a_20103_8443# VSS.t51 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X809 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD.t373 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X810 VDD VCO_DFF_C_0.VCO_C_0.OUTB a_41879_n196# VDD.t262 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X811 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t572 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X812 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.IN a_24437_9224# VDD.t402 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X813 VDD S6.t8 mux_magic_3.AND2_magic_0.A VDD.t772 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X814 a_25706_n567# VCTRL2.t58 VSS.t444 VSS.t442 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X815 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD.t140 VDD.t139 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X816 RES_74k_1.M VSS.t320 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X817 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t149 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X818 RES_74k_1.M VSS.t319 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X819 RES_74k_1.M VSS.t318 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X820 a_25706_n567# VCTRL2.t59 VSS.t445 VSS.t158 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X821 a_19903_9637# S6.t9 a_20103_9637# VSS.t723 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X822 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN VDD.t401 VDD.t268 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X823 RES_74k_1.M VSS.t317 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X824 RES_74k_1.M VSS.t316 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X825 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUT.t2 VDD.t31 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X826 a_42928_10426# a_42628_9804# VDD.t93 ppolyf_u r_width=1.1u r_length=2.6u
X827 A_MUX_0.Tr_Gate_1.CLK S4.t15 VDD.t118 VDD.t111 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X828 VCO_DFF_C_0.VCTRL A_MUX_0.Tr_Gate_1.CLK RES_74k_1.P VSS.t107 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X829 a_31468_10271# DN.t8 VDD.t626 VDD.t104 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X830 VDD.t198 VDD.t196 VDD.t198 VDD.t197 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X831 VCO_DFF_C_0.VCTRL a_45158_5339# RES_74k_1.P VDD.t291 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X832 VDD a_27722_11758# mux_magic_0.OR_magic_0.A VDD.t250 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X833 a_19897_10547# S1.t9 VDD.t657 VDD.t656 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X834 VDD.t195 VDD.t193 VDD.t195 VDD.t194 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X835 VSS UP_INPUT.t3 a_27922_10564# VSS.t729 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X836 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t347 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X837 RES_74k_1.M VSS.t315 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X838 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VSS.t651 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X839 A_MUX_0.Tr_Gate_1.CLK S4.t16 VDD.t119 VDD.t113 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X840 a_34443_2598# VCTRL2.t60 VSS.t447 VSS.t446 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X841 a_44716_1837# VCO_DFF_C_0.VCO_C_0.OUTB VDD.t456 VDD.t371 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X842 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_1284# OUTB.t13 VDD.t263 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X843 A_MUX_0.Tr_Gate_1.CLK S4.t17 VSS.t115 VSS.t62 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X844 VSS VCTRL2.t61 a_34443_2598# VSS.t448 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X845 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VSS.t636 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X846 VSS PFD_T2_0.UP a_27922_11758# VSS.t759 nfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X847 mux_magic_1.AND2_magic_0.A S3.t9 VSS.t747 VSS.t746 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X848 VCO_DFF_C_0.VCTRL S4.t18 VCTRL_IN.t5 VSS.t116 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X849 RES_74k_1.M VSS.t314 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X850 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL VDD.t160 VDD.t147 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X851 a_44128_10426# a_44428_9804# VDD.t55 ppolyf_u r_width=1.1u r_length=2.6u
X852 VSS VCTRL2.t62 a_25706_n567# VSS.t451 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X853 RES_74k_1.M VSS.t313 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X854 a_45628_9598# a_45928_8976# VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X855 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t323 VDD.t322 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X856 VSS a_22966_11778# a_22880_10947# VSS.t702 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X857 a_42628_9598# a_42628_8770# VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X858 RES_74k_1.M VSS.t312 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X859 A_MUX_0.Tr_Gate_1.CLK S4.t19 VSS.t117 VSS.t62 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X860 a_34443_2598# VCTRL2.t63 VSS.t454 VSS.t446 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X861 VDD.t192 VDD.t190 VDD.t192 VDD.t191 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X862 VCTRL_IN a_42763_5679# VCO_DFF_C_0.VCTRL VDD.t75 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X863 a_19903_9637# VSS.t776 VDD.t840 VDD.t839 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X864 VSS VCTRL2.t64 a_34443_2598# VSS.t448 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X865 RES_74k_1.M VSS.t311 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X866 RES_74k_1.M VSS.t310 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X867 VSS VCTRL2.t65 a_25706_n567# VSS.t457 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X868 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t321 VDD.t320 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X869 VSS.t188 VSS.t186 VSS.t188 VSS.t187 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X870 VDD a_19897_11741# mux_magic_2.OR_magic_0.A VDD.t94 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X871 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VSS.t87 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X872 a_34443_2598# VCTRL2.t66 VSS.t460 VSS.t153 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X873 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t338 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X874 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VSS.t74 VSS.t73 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X875 VSS VCTRL2.t67 a_34443_2598# VSS.t155 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X876 mux_magic_3.AND2_magic_0.A S6.t10 VDD.t778 VDD.t397 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X877 RES_74k_1.M VSS.t309 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X878 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t491 VDD.t322 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X879 VDD S3.t10 mux_magic_1.AND2_magic_0.A VDD.t805 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X880 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB a_25706_n567# VSS.t83 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X881 a_43828_9598# a_44128_8976# VDD.t25 ppolyf_u r_width=1.1u r_length=2.6u
X882 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD.t372 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X883 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUT.t9 VSS.t36 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X884 VDD a_22966_11778# PFD_T2_0.INV_mag_0.IN VDD.t737 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X885 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VSS.t581 VSS.t133 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X886 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t572 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X887 RES_74k_1.M VSS.t308 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X888 VSS.t185 VSS.t183 VSS.t185 VSS.t184 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X889 a_45328_8770# a_45628_8148# VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X890 PFD_T2_0.INV_mag_1.IN a_22967_8787# VDD.t267 VDD.t266 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X891 RES_74k_1.P RES_74k_1.P VDD.t69 ppolyf_u r_width=1.1u r_length=2.6u
X892 a_25706_n567# VCTRL2.t68 VSS.t463 VSS.t158 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X893 VSS.t182 VSS.t180 VSS.t182 VSS.t181 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X894 RES_74k_1.M VSS.t307 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X895 a_29415_9553# mux_magic_1.OR_magic_0.B a_29415_8145# VDD.t473 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X896 RES_74k_1.P RES_74k_1.P VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X897 VSS VCTRL2.t69 a_25706_n567# VSS.t150 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X898 VDD VCO_DFF_C_0.VCO_C_0.OUTB a_44716_1837# VDD.t370 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X899 RES_74k_1.M VSS.t306 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X900 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK VCO_DFF_C_0.VCTRL VSS.t106 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X901 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t461 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X902 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.OUTB VDD.t813 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X903 RES_74k_1.M VSS.t305 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X904 RES_74k_1.P RES_74k_1.P VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X905 a_41879_n196# VCO_DFF_C_0.VCO_C_0.OUTB VDD.t453 VDD.t260 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X906 RES_74k_1.P RES_74k_1.P VDD.t69 ppolyf_u r_width=1.1u r_length=2.6u
X907 RES_74k_1.M VSS.t304 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X908 RES_74k_1.P VSS.t709 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X909 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT VDD.t136 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X910 RES_74k_1.M VSS.t303 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X911 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_n196# VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD.t260 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X912 VDD.t189 VDD.t187 VDD.t189 VDD.t188 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X913 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB VSS.t481 VSS.t480 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X914 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t147 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X915 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t672 VDD.t580 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X916 VDD S6.t11 a_19903_9637# VDD.t779 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X917 RES_74k_1.M VSS.t302 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X918 a_45928_12082# a_45628_11460# VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X919 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT a_34443_2598# VSS.t88 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X920 RES_74k_1.M VSS.t301 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X921 VDD a_25556_11637# PFD_T2_0.UP VDD.t245 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X922 a_31940_9626# ITAIL1.t12 RES_74k_1.P VSS.t43 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X923 OUTB a_41879_1284# VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD.t262 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X924 RES_74k_1.P RES_74k_1.P VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X925 RES_74k_1.M VSS.t300 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X926 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD.t615 VDD.t41 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X927 OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VSS.t650 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X928 a_34443_2598# VCTRL2.t70 VSS.t467 VSS.t466 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X929 RES_74k_1.M VSS.t299 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X930 RES_74k_1.M VSS.t298 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X931 a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VSS.t649 VSS.t648 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X932 RES_74k_1.P VSS.t708 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X933 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT a_34443_2598# VSS.t500 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X934 mux_magic_0.AND2_magic_0.A S2.t10 VSS.t684 VSS.t683 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X935 VDD PFD_T2_0.Buffer_V_2_0.IN a_25557_8739# VDD.t392 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X936 a_21437_10708# mux_magic_2.OR_magic_0.B VSS.t614 VSS.t613 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X937 a_45628_11254# a_45928_10632# VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X938 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t711 VDD.t710 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X939 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VSS.t479 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X940 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VSS.t87 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X941 a_29262_10725# mux_magic_0.OR_magic_0.B a_29262_12133# VDD.t1 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X942 mux_magic_2.OR_magic_0.B a_19897_10547# VSS.t612 VSS.t611 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X943 RES_74k_1.P RES_74k_1.P VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X944 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t490 VDD.t313 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X945 RES_74k_1.M VSS.t297 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X946 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VSS.t478 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X947 RES_74k_1.P ITAIL.t26 a_31732_10267# VDD.t539 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X948 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t571 VDD.t570 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X949 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t567 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X950 VSS PFD_T2_0.INV_mag_1.OUT PFD_T2_0.Buffer_V_2_1.IN VSS.t5 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X951 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VDD.t317 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X952 a_34443_2598# VCTRL2.t71 VSS.t597 VSS.t466 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X953 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VDD.t487 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X954 VSS.t179 VSS.t177 VSS.t179 VSS.t178 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X955 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t559 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X956 OUTB OUT.t29 VDD.t51 VDD.t41 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X957 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK OUTB.t16 VSS.t647 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X958 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD.t812 VDD.t811 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X959 VDD.t186 VDD.t184 VDD.t186 VDD.t185 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X960 a_25706_n567# VCTRL2.t72 VSS.t598 VSS.t504 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X961 VSS OUT.t30 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VSS.t36 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X962 VSS VCTRL2.t73 a_25706_n567# VSS.t451 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X963 a_21437_12116# mux_magic_2.OR_magic_0.B a_21437_10708# VDD.t545 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X964 VSS PFD_T2_0.INV_mag_1.OUT PFD_T2_0.Buffer_V_2_1.IN VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X965 mux_magic_1.OR_magic_0.A a_27875_8520# VSS.t144 VSS.t143 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X966 a_21443_9476# mux_magic_3.OR_magic_0.B a_21443_8068# VDD.t21 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X967 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t316 VDD.t315 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X968 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_1837# VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t371 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X969 VSS PFD_T2_0.Buffer_V_2_1.IN a_25556_11637# VSS.t84 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X970 RES_74k_1.M VSS.t296 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X971 OUTB OUT.t31 VDD.t52 VDD.t43 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X972 a_23836_10693# PFD_T2_0.INV_mag_0.IN PFD_T2_0.Buffer_V_2_1.IN VSS.t471 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X973 a_29415_8145# mux_magic_1.OR_magic_0.A VDD.t307 VDD.t306 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X974 a_43528_10426# a_43828_9804# VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X975 VSS S4.t20 a_42763_5679# VSS.t67 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X976 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t32 VDD.t53 VDD.t34 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X977 VSS VCTRL2.t74 a_34443_2598# VSS.t428 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X978 a_25706_n567# VCTRL2.t75 VSS.t603 VSS.t442 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X979 mux_magic_1.OR_magic_0.B a_27875_9714# VSS.t61 VSS.t60 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X980 mux_magic_1.AND2_magic_0.A S3.t11 VDD.t810 VDD.t800 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X981 RES_74k_1.P RES_74k_1.P VDD.t93 ppolyf_u r_width=1.1u r_length=2.6u
X982 PFD_T2_0.INV_mag_0.IN PFD_T2_0.FIN a_22880_10947# VSS.t137 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X983 RES_74k_1.P RES_74k_1.P VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X984 a_41879_n196# VCO_DFF_C_0.VCO_C_0.OUTB VDD.t452 VDD.t263 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X985 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD.t566 VDD.t565 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X986 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t669 VDD.t668 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X987 RES_74k_1.M VSS.t295 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X988 VDD OUT.t33 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD.t38 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X989 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT.t34 VDD.t60 VDD.t36 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X990 a_21443_8068# mux_magic_3.OR_magic_0.B a_21443_9476# VDD.t20 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X991 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t314 VDD.t313 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X992 a_25706_n567# VCTRL2.t76 VSS.t604 VSS.t442 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X993 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t155 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X994 RES_74k_1.M VSS.t294 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X995 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VSS.t616 VSS.t615 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X996 a_27722_11758# PFD_T2_0.UP VDD.t828 VDD.t827 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X997 VDD VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD.t449 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X998 VDD.t183 VDD.t181 VDD.t183 VDD.t182 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X999 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VSS.t86 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1000 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VSS.t82 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1001 VSS VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT VSS.t70 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1002 RES_74k_1.M VSS.t293 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1003 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD.t707 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1004 VDD VCO_DFF_C_0.VCO_C_0.OUTB a_41879_n196# VDD.t261 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1005 VDD ITAIL.t0 ITAIL.t1 VDD.t534 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X1006 a_42928_12082# a_42628_11460# VDD.t93 ppolyf_u r_width=1.1u r_length=2.6u
X1007 a_46528_12082# a_46828_11254# VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X1008 VSS VCTRL2.t77 a_34443_2598# VSS.t428 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X1009 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VSS.t750 VSS.t749 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1010 RES_74k_1.M VSS.t292 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1011 mux_magic_0.AND2_magic_0.A S2.t11 VSS.t686 VSS.t685 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1012 RES_74k_1.M VSS.t291 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1013 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB VDD.t446 VDD.t445 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1014 mux_magic_2.AND2_magic_0.A S1.t10 VDD.t659 VDD.t658 pfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1015 a_27875_8520# mux_magic_1.AND2_magic_0.A a_28075_8520# VSS.t141 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1016 a_45328_10426# a_45028_9804# VDD.t57 ppolyf_u r_width=1.1u r_length=2.6u
X1017 OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VSS.t626 VSS.t625 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1018 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD.t461 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1019 a_46828_9598# a_46528_8976# VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X1020 RES_74k_1.M VSS.t290 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1021 VSS mux_magic_1.OR_magic_0.A a_29415_9553# VSS.t112 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1022 a_43228_9598# a_43528_8976# VDD.t63 ppolyf_u r_width=1.1u r_length=2.6u
X1023 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUT.t0 VDD.t45 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1024 a_22881_9554# a_22967_8787# VSS.t102 VSS.t101 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1025 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t152 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1026 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD.t324 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1027 VDD S1.t11 a_19897_10547# VDD.t660 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1028 PFD_T2_0.INV_mag_1.IN a_22967_8787# VDD.t265 VDD.t264 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1029 a_42628_11254# a_42928_10632# VDD.t93 ppolyf_u r_width=1.1u r_length=2.6u
X1030 VSS.t176 VSS.t174 VSS.t176 VSS.t175 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X1031 VDD a_22966_11778# PFD_T2_0.INV_mag_0.IN VDD.t423 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1032 mux_magic_3.AND2_magic_0.A S6.t12 VSS.t725 VSS.t724 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1033 a_46828_11254# a_46528_10632# VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X1034 a_19903_8443# mux_magic_3.AND2_magic_0.A VDD.t71 VDD.t70 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1035 a_27875_9714# S3.t12 a_28075_9714# VSS.t748 nfet_03v3 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.56u
X1036 mux_magic_3.OR_magic_0.A a_19903_8443# VSS.t714 VSS.t713 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1037 RES_74k_1.M VSS.t289 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1038 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VSS.t646 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1039 RES_74k_1.P ITAIL1.t13 a_31940_9626# VSS.t39 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X1040 VDD PFD_T2_0.INV_mag_0.IN PFD_T2_0.Buffer_V_2_1.IN VDD.t423 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1041 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t484 VDD.t483 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1042 VDD S2.t12 mux_magic_0.AND2_magic_0.A VDD.t610 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1043 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT VDD.t133 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1044 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB a_25706_n567# VSS.t81 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1045 RES_74k_1.M VSS.t288 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1046 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD.t562 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1047 a_21443_8068# mux_magic_3.OR_magic_0.A VDD.t782 VDD.t22 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1048 VDD OUT.t35 OUTB.t0 VDD.t31 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1049 mux_magic_2.AND2_magic_0.A S1.t12 VSS.t664 VSS.t663 nfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1050 a_31732_10267# ITAIL.t27 RES_74k_1.P VDD.t538 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X1051 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_41879_1284# VDD.t262 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1052 mux_magic_3.OR_magic_0.B a_19903_9637# VSS.t693 VSS.t692 nfet_03v3 ad=0.493p pd=3.12u as=0.493p ps=3.12u w=1.12u l=0.56u
X1053 VCO_DFF_C_0.VCTRL S4.t21 VCTRL_IN.t4 VSS.t65 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1054 RES_74k_1.P VSS.t707 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X1055 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t667 VDD.t598 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1056 VSS VCTRL2.t78 a_25706_n567# VSS.t517 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X1057 a_21437_12116# mux_magic_2.OR_magic_0.A VDD.t12 VDD.t11 pfet_03v3 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.56u
X1058 VSS PFD_T2_0.INV_mag_0.IN a_23836_10693# VSS.t468 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1059 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD.t132 VDD.t131 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1060 RES_74k_1.M VSS.t287 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1061 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_44716_1837# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD.t370 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1062 a_45028_9598# a_44728_8976# VDD.t79 ppolyf_u r_width=1.1u r_length=2.6u
X1063 RES_74k_1.M VSS.t286 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1064 VDD VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD.t149 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X1065 RES_74k_1.P RES_74k_1.P VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X1066 RES_74k_1.M VSS.t285 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1067 mux_magic_0.OR_magic_0.B a_27722_10564# VDD.t388 VDD.t387 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1068 a_27875_8520# PFD_T2_0.DOWN VDD.t27 VDD.t26 pfet_03v3 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.56u
X1069 VSS VCTRL2.t79 a_25706_n567# VSS.t457 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1070 RES_74k_1.M VSS.t284 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1071 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD.t559 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1072 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VSS.t80 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X1073 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN a_23837_9553# VSS.t416 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1074 a_46528_8770# a_46228_8148# VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X1075 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL VDD.t148 VDD.t147 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
R0 VDD.n1767 VDD.n569 130000
R1 VDD.n1548 VDD.n718 129000
R2 VDD.n1768 VDD.n1767 65000
R3 VDD.n1503 VDD.n718 64500
R4 VDD.n1957 VDD.n1956 6501.29
R5 VDD.t540 VDD.t11 1194.81
R6 VDD.n1715 VDD.n1714 947.995
R7 VDD.n1769 VDD.n561 947.995
R8 VDD.n1520 VDD.n1496 947.995
R9 VDD.n1511 VDD.n1504 947.995
R10 VDD.n1714 VDD.n1705 944.883
R11 VDD.n1705 VDD.n568 944.883
R12 VDD.n1513 VDD.n1512 944.883
R13 VDD.n1512 VDD.n1511 944.883
R14 VDD.n1769 VDD.n1768 842.52
R15 VDD.n1503 VDD.n1496 842.52
R16 VDD.n172 VDD.t361 841.558
R17 VDD.n156 VDD.t17 714.287
R18 VDD.t527 VDD.t658 566.929
R19 VDD.t527 VDD.t525 566.929
R20 VDD.t11 VDD.t546 561.039
R21 VDD.n172 VDD.t363 500
R22 VDD.t654 VDD.n197 481.685
R23 VDD.t80 VDD.n2041 450.401
R24 VDD.t70 VDD.n324 450.401
R25 VDD.n410 VDD.t380 450.401
R26 VDD.n1957 VDD.n1896 447.029
R27 VDD.t406 VDD.t395 432.243
R28 VDD.t389 VDD.n99 421.245
R29 VDD.t730 VDD.n302 421.245
R30 VDD.t99 VDD.n401 421.245
R31 VDD.t387 VDD.t389 395.604
R32 VDD.t663 VDD.t387 395.604
R33 VDD.t788 VDD.t420 395.604
R34 VDD.t420 VDD.t761 395.604
R35 VDD.t547 VDD.t545 395.604
R36 VDD.t17 VDD.t13 395.604
R37 VDD.t97 VDD.t727 395.604
R38 VDD.t543 VDD.t540 395.604
R39 VDD.t790 VDD.t543 395.604
R40 VDD.t793 VDD.t660 395.604
R41 VDD.t660 VDD.t656 395.604
R42 VDD.t733 VDD.t730 395.604
R43 VDD.t836 VDD.t733 395.604
R44 VDD.t839 VDD.t779 395.604
R45 VDD.t779 VDD.t399 395.604
R46 VDD.t102 VDD.t99 395.604
R47 VDD.t257 VDD.t102 395.604
R48 VDD.t255 VDD.t797 395.604
R49 VDD.t797 VDD.t795 395.604
R50 VDD.t253 VDD.t829 391.305
R51 VDD.t758 VDD.t301 391.305
R52 VDD.t385 VDD.t28 391.305
R53 VDD.t530 VDD.n189 384.615
R54 VDD.n1766 VDD.n527 371.986
R55 VDD.n1536 VDD.n725 371.986
R56 VDD.n1754 VDD.n1753 353.928
R57 VDD.n1551 VDD.n715 353.928
R58 VDD.n1755 VDD.n1754 350.877
R59 VDD.n1759 VDD.n570 350.877
R60 VDD.n1547 VDD.n720 350.877
R61 VDD.n1551 VDD.n1550 350.877
R62 VDD.t768 VDD.t441 339.613
R63 VDD.t548 VDD.t15 333.334
R64 VDD.t64 VDD.t66 316.279
R65 VDD.t395 VDD.t392 316.279
R66 VDD.n1759 VDD.n569 312.866
R67 VDD.n1548 VDD.n1547 312.866
R68 VDD.n1921 VDD.n1920 310.428
R69 VDD.n1922 VDD.n1921 307.495
R70 VDD.n1922 VDD.n1905 307.495
R71 VDD.n1907 VDD.n1906 307.495
R72 VDD.n1931 VDD.n1907 307.495
R73 VDD.n1954 VDD.n1898 307.495
R74 VDD.n1947 VDD.n1898 307.495
R75 VDD.n1945 VDD.n1944 307.495
R76 VDD.n1944 VDD.n1932 307.495
R77 VDD.n1937 VDD.n1896 307.495
R78 VDD.n1955 VDD.n1897 304.911
R79 VDD.t527 VDD.n188 294.873
R80 VDD.n99 VDD.n74 289.856
R81 VDD.n302 VDD.n301 289.856
R82 VDD.n401 VDD.n400 289.856
R83 VDD.t221 VDD.n1766 283.627
R84 VDD.n1536 VDD.t226 283.627
R85 VDD.t248 VDD.t245 282.159
R86 VDD.t765 VDD.t768 282.159
R87 VDD.t546 VDD.n172 280.519
R88 VDD.n1757 VDD.t152 279.885
R89 VDD.t147 VDD.n1549 279.885
R90 VDD.t206 VDD.n1945 263.567
R91 VDD.t725 VDD.n204 260.074
R92 VDD.t827 VDD.n84 246.871
R93 VDD.n292 VDD.t304 246.871
R94 VDD.n384 VDD.t26 246.871
R95 VDD.t206 VDD.n1906 235.143
R96 VDD.n207 VDD.n206 230.769
R97 VDD.n197 VDD.n196 230.769
R98 VDD.n198 VDD.n178 230.769
R99 VDD.n91 VDD.n90 228.262
R100 VDD.n335 VDD.n334 228.262
R101 VDD.n394 VDD.n379 228.262
R102 VDD.n2043 VDD.n2042 227.028
R103 VDD.n326 VDD.n325 227.028
R104 VDD.n386 VDD.n385 227.028
R105 VDD.t608 VDD.n113 225.081
R106 VDD.t397 VDD.n316 225.081
R107 VDD.t800 VDD.n2020 225.081
R108 VDD.t206 VDD.n1931 209.303
R109 VDD.n100 VDD.t663 197.803
R110 VDD.n100 VDD.t788 197.803
R111 VDD.n172 VDD.t547 197.803
R112 VDD.t727 VDD.n205 197.803
R113 VDD.n205 VDD.t725 197.803
R114 VDD.n173 VDD.t790 197.803
R115 VDD.n173 VDD.t793 197.803
R116 VDD.n303 VDD.t836 197.803
R117 VDD.n303 VDD.t839 197.803
R118 VDD.n402 VDD.t257 197.803
R119 VDD.n402 VDD.t255 197.803
R120 VDD.t829 VDD.n89 195.653
R121 VDD.n89 VDD.t827 195.653
R122 VDD.t301 VDD.n333 195.653
R123 VDD.n333 VDD.t304 195.653
R124 VDD.t28 VDD.n393 195.653
R125 VDD.n393 VDD.t26 195.653
R126 VDD.t737 VDD.t439 188.018
R127 VDD.t439 VDD.t423 188.018
R128 VDD.t423 VDD.t437 188.018
R129 VDD.t437 VDD.t426 188.018
R130 VDD.t426 VDD.t435 188.018
R131 VDD.t435 VDD.t365 188.018
R132 VDD.t365 VDD.t368 188.018
R133 VDD.t392 VDD.n256 184.496
R134 VDD.n1932 VDD.t194 180.88
R135 VDD.t270 VDD.t285 180.213
R136 VDD.t277 VDD.t270 180.213
R137 VDD.t264 VDD.t274 180.213
R138 VDD.t274 VDD.t268 180.213
R139 VDD.t268 VDD.t280 180.213
R140 VDD.t280 VDD.t283 180.213
R141 VDD.t610 VDD.n112 172.562
R142 VDD.t772 VDD.n315 172.562
R143 VDD.n412 VDD.t805 172.562
R144 VDD.n172 VDD.t548 166.667
R145 VDD.n119 VDD.t765 164.593
R146 VDD.n257 VDD.t264 161.661
R147 VDD.n1584 VDD.t191 160.7
R148 VDD.n1743 VDD.t218 160.284
R149 VDD.n172 VDD.n147 155.679
R150 VDD.n99 VDD.t477 145.662
R151 VDD.n302 VDD.t783 145.662
R152 VDD.n401 VDD.t308 145.662
R153 VDD.t2 VDD.t3 136.796
R154 VDD.t477 VDD.t1 136.796
R155 VDD.t21 VDD.t20 136.796
R156 VDD.t783 VDD.t22 136.796
R157 VDD.t473 VDD.t474 136.796
R158 VDD.t306 VDD.t308 136.796
R159 VDD.n204 VDD.t651 135.531
R160 VDD.n2041 VDD.n2040 135.048
R161 VDD.n324 VDD.n323 135.048
R162 VDD.n411 VDD.n410 135.048
R163 VDD.n84 VDD.t82 133.333
R164 VDD.t72 VDD.n292 133.333
R165 VDD.t377 VDD.n384 133.333
R166 VDD.n1684 VDD.n1683 132.696
R167 VDD.n1675 VDD.n1674 132.696
R168 VDD.n1609 VDD.n1608 132.696
R169 VDD.n693 VDD.n650 132.696
R170 VDD.n675 VDD.n674 132.696
R171 VDD.n1114 VDD.n1113 132.696
R172 VDD.n1204 VDD.n1203 132.696
R173 VDD.n1623 VDD.n1620 132.696
R174 VDD.n256 VDD.t64 131.784
R175 VDD.n196 VDD.t523 130.037
R176 VDD.n1685 VDD.n1684 128.591
R177 VDD.t508 VDD.n594 128.591
R178 VDD.n1691 VDD.n594 128.591
R179 VDD.n1693 VDD.n1692 128.591
R180 VDD.n1674 VDD.n1647 128.591
R181 VDD.n1657 VDD.t315 128.591
R182 VDD.n1667 VDD.n1657 128.591
R183 VDD.n1666 VDD.n1665 128.591
R184 VDD.n1601 VDD.n621 128.591
R185 VDD.n1603 VDD.n1602 128.591
R186 VDD.n1603 VDD.t677 128.591
R187 VDD.n1608 VDD.n612 128.591
R188 VDD.n707 VDD.n641 128.591
R189 VDD.n701 VDD.n700 128.591
R190 VDD.n700 VDD.t577 128.591
R191 VDD.n699 VDD.n650 128.591
R192 VDD.n684 VDD.n683 128.591
R193 VDD.n682 VDD.n659 128.591
R194 VDD.t813 VDD.n659 128.591
R195 VDD.n675 VDD.n670 128.591
R196 VDD.n1105 VDD.n1104 128.591
R197 VDD.n1111 VDD.n1088 128.591
R198 VDD.t38 VDD.n1111 128.591
R199 VDD.n1114 VDD.n1112 128.591
R200 VDD.n1211 VDD.n1189 128.591
R201 VDD.t707 VDD.n1189 128.591
R202 VDD.n1204 VDD.n1197 128.591
R203 VDD.n1619 VDD.n1618 128.591
R204 VDD.n1632 VDD.n1631 128.591
R205 VDD.n1631 VDD.t136 128.591
R206 VDD.n1630 VDD.n1620 128.591
R207 VDD.t94 VDD.n156 128.206
R208 VDD.t250 VDD.n74 126.812
R209 VDD.n301 VDD.t755 126.812
R210 VDD.n400 VDD.t382 126.812
R211 VDD.n1937 VDD.t194 126.615
R212 VDD.n98 VDD.t2 122.23
R213 VDD.n275 VDD.t21 122.23
R214 VDD.n372 VDD.t473 122.23
R215 VDD.n2062 VDD.t78 122.1
R216 VDD.t291 VDD.n2124 121.091
R217 VDD.n2026 VDD.t408 120.213
R218 VDD.t441 VDD.t744 118.191
R219 VDD.t431 VDD.t752 118.191
R220 VDD.t415 VDD.t746 118.191
R221 VDD.n1638 VDD.t487 118.061
R222 VDD.n1676 VDD.t317 118.061
R223 VDD.n1610 VDD.t668 118.061
R224 VDD.t570 VDD.n692 118.061
R225 VDD.t819 VDD.n673 118.061
R226 VDD.t710 VDD.n1202 118.061
R227 VDD.n1624 VDD.t139 118.061
R228 VDD.n119 VDD.t248 117.567
R229 VDD.t77 VDD.n2060 116.044
R230 VDD.t266 VDD.t406 113.275
R231 VDD.t288 VDD.t402 113.275
R232 VDD.t272 VDD.t443 113.275
R233 VDD.n1692 VDD.t501 110.808
R234 VDD.t332 VDD.n1666 110.808
R235 VDD.t683 VDD.n1601 110.808
R236 VDD.t589 VDD.n641 110.808
R237 VDD.n683 VDD.t811 110.808
R238 VDD.n1105 VDD.t34 110.808
R239 VDD.t131 VDD.n1619 110.808
R240 VDD.n1212 VDD.t712 109.439
R241 VDD.t403 VDD.t737 108.948
R242 VDD.n2061 VDD.t77 105.954
R243 VDD.n2125 VDD.t295 104.945
R244 VDD.t285 VDD.t432 104.418
R245 VDD.n207 VDD.t94 102.564
R246 VDD.n1768 VDD.n568 102.362
R247 VDD.n1513 VDD.n1503 102.362
R248 VDD.n91 VDD.t250 101.45
R249 VDD.n335 VDD.t755 101.45
R250 VDD.n379 VDD.t382 101.45
R251 VDD.n2125 VDD.t291 100.909
R252 VDD.n188 VDD.t523 100.734
R253 VDD.t78 VDD.n2061 99.8996
R254 VDD.n1767 VDD.t152 99.5009
R255 VDD.t147 VDD.n718 99.0846
R256 VDD.n1120 VDD.t36 98.4957
R257 VDD.t206 VDD.n1897 98.1917
R258 VDD.n1695 VDD.t483 97.5562
R259 VDD.n2026 VDD.t417 96.809
R260 VDD.t48 VDD.n1103 95.9239
R261 VDD.n1660 VDD.t327 95.9239
R262 VDD.n1594 VDD.t692 95.9239
R263 VDD.n708 VDD.t562 95.9239
R264 VDD.n687 VDD.t816 95.9239
R265 VDD.n1615 VDD.t133 95.9239
R266 VDD.n178 VDD.t651 95.2386
R267 VDD.n2043 VDD.t82 93.6942
R268 VDD.n326 VDD.t72 93.6942
R269 VDD.n386 VDD.t377 93.6942
R270 VDD.t213 VDD.n529 92.4235
R271 VDD.t203 VDD.n1535 92.4235
R272 VDD.n2060 VDD.t75 89.8088
R273 VDD.n2127 VDD.t293 88.7997
R274 VDD.n811 VDD.n810 86.1787
R275 VDD.t714 VDD.n1178 84.8158
R276 VDD.n2124 VDD.t298 84.7634
R277 VDD.n2062 VDD.t76 83.7543
R278 VDD.n2040 VDD.t120 76.0991
R279 VDD.n323 VDD.t770 76.0991
R280 VDD.t802 VDD.n411 76.0991
R281 VDD.n1223 VDD.n1179 73.8719
R282 VDD.t206 VDD.n1905 72.3519
R283 VDD.t744 VDD.t431 70.1759
R284 VDD.t752 VDD.t415 70.1759
R285 VDD.t746 VDD.t403 70.1759
R286 VDD.n1755 VDD.t152 70.1759
R287 VDD.n1550 VDD.t147 70.1759
R288 VDD.n198 VDD.t654 69.5976
R289 VDD.n2042 VDD.t80 68.469
R290 VDD.n325 VDD.t70 68.469
R291 VDD.n385 VDD.t380 68.469
R292 VDD.t402 VDD.t266 67.2571
R293 VDD.t443 VDD.t288 67.2571
R294 VDD.t432 VDD.t272 67.2571
R295 VDD.t221 VDD.n570 67.252
R296 VDD.t226 VDD.n720 67.252
R297 VDD.n1042 VDD.n1026 66.348
R298 VDD.n1043 VDD.n1042 64.296
R299 VDD.t41 VDD.n1022 64.296
R300 VDD.n1059 VDD.n1022 64.296
R301 VDD.n1063 VDD.n1062 64.296
R302 VDD.n1069 VDD.n1068 64.296
R303 VDD.n206 VDD.t97 62.2716
R304 VDD.n930 VDD.t263 61.8854
R305 VDD.n90 VDD.t253 61.5947
R306 VDD.n334 VDD.t758 61.5947
R307 VDD.n394 VDD.t385 61.5947
R308 VDD.n1142 VDD.t370 60.8721
R309 VDD.n929 VDD.t262 60.7435
R310 VDD.t372 VDD.n1144 59.702
R311 VDD.t260 VDD.n926 59.0509
R312 VDD.n112 VDD.t120 58.9501
R313 VDD.n315 VDD.t770 58.9501
R314 VDD.n412 VDD.t802 58.9501
R315 VDD.t371 VDD.n1146 58.9084
R316 VDD.t373 VDD.n1147 57.7119
R317 VDD.n1036 VDD.t45 57.456
R318 VDD.n191 VDD.t530 56.849
R319 VDD.n849 VDD.n848 56.5021
R320 VDD.n911 VDD.n910 56.5021
R321 VDD.n1062 VDD.t31 55.4041
R322 VDD.n1964 VDD.n1890 54.5384
R323 VDD.n1281 VDD.n1280 54.5384
R324 VDD.n981 VDD.n840 53.3521
R325 VDD.n967 VDD.n888 53.3521
R326 VDD.n964 VDD.n963 53.3521
R327 VDD.n909 VDD.n905 53.3521
R328 VDD.n927 VDD.t260 52.7113
R329 VDD.n1820 VDD.n1819 52.4568
R330 VDD.n1435 VDD.n740 52.0405
R331 VDD.n1148 VDD.t373 51.7418
R332 VDD.n15 VDD.t537 51.2378
R333 VDD.t226 VDD.n718 50.3542
R334 VDD.n1767 VDD.t221 49.9381
R335 VDD.n1148 VDD.t372 49.7517
R336 VDD.n927 VDD.t262 49.6993
R337 VDD.t5 VDD.t10 49.5054
R338 VDD.t10 VDD.t6 49.5054
R339 VDD.t6 VDD.t56 49.5054
R340 VDD.t8 VDD.t7 49.5054
R341 VDD.t57 VDD.t8 49.5054
R342 VDD.t79 VDD.t57 49.5054
R343 VDD.t54 VDD.t79 49.5054
R344 VDD.t54 VDD.t55 49.5054
R345 VDD.t55 VDD.t25 49.5054
R346 VDD.t25 VDD.t4 49.5054
R347 VDD.t4 VDD.t63 49.5054
R348 VDD.t93 VDD.t9 49.5054
R349 VDD.t0 VDD.t93 49.5054
R350 VDD.t69 VDD.t0 49.5054
R351 VDD.n24 VDD.t534 47.9334
R352 VDD.t445 VDD.n955 46.5121
R353 VDD.n1068 VDD.t43 46.5121
R354 VDD.n1827 VDD.n517 45.7957
R355 VDD.n1826 VDD.n518 45.7957
R356 VDD.n1833 VDD.n513 45.7957
R357 VDD.t336 VDD.n1834 45.7957
R358 VDD.n1853 VDD.n489 45.7957
R359 VDD.n1844 VDD.n1841 45.7957
R360 VDD.n2009 VDD.n423 45.7957
R361 VDD.n431 VDD.n430 45.7957
R362 VDD.n2002 VDD.n2001 45.7957
R363 VDD.n438 VDD.n432 45.7957
R364 VDD.n1995 VDD.n439 45.7957
R365 VDD.n450 VDD.n449 45.7957
R366 VDD.n458 VDD.n451 45.7957
R367 VDD.n1979 VDD.n457 45.7957
R368 VDD.n1880 VDD.n1879 45.7957
R369 VDD.n1888 VDD.n1881 45.7957
R370 VDD.n1965 VDD.n1889 45.7957
R371 VDD.n1288 VDD.n801 45.7957
R372 VDD.n1287 VDD.n803 45.7957
R373 VDD.n1296 VDD.n1295 45.7957
R374 VDD.n1305 VDD.n789 45.7957
R375 VDD.n794 VDD.n793 45.7957
R376 VDD.n1369 VDD.n780 45.7957
R377 VDD.n1379 VDD.n1378 45.7957
R378 VDD.n1386 VDD.n768 45.7957
R379 VDD.n1385 VDD.n769 45.7957
R380 VDD.n1393 VDD.n764 45.7957
R381 VDD.n1403 VDD.n758 45.7957
R382 VDD.n1410 VDD.n754 45.7957
R383 VDD.n1420 VDD.n748 45.7957
R384 VDD.n1426 VDD.n744 45.7957
R385 VDD.n1428 VDD.n1427 45.7957
R386 VDD.n1436 VDD.n739 45.7957
R387 VDD.n1419 VDD.t572 45.3794
R388 VDD.n968 VDD.n887 45.1441
R389 VDD.n1947 VDD.t206 43.9281
R390 VDD.n1147 VDD.t371 43.7816
R391 VDD.t347 VDD.n1971 43.2978
R392 VDD.n802 VDD.t580 42.8814
R393 VDD.t575 VDD.n1394 42.8814
R394 VDD.n2008 VDD.t338 42.4651
R395 VDD.t13 VDD.n147 42.125
R396 VDD.n1144 VDD.t370 41.7915
R397 VDD.n0 VDD.t5 41.7644
R398 VDD.n2050 VDD.t69 41.7644
R399 VDD.t263 VDD.n929 41.6672
R400 VDD.n1693 VDD.t483 39.6722
R401 VDD.n1665 VDD.t327 39.6722
R402 VDD.t692 VDD.n621 39.6722
R403 VDD.t562 VDD.n707 39.6722
R404 VDD.n684 VDD.t816 39.6722
R405 VDD.n894 VDD.n893 39.6722
R406 VDD.n1104 VDD.t48 39.6722
R407 VDD.n1618 VDD.t133 39.6722
R408 VDD.n2086 VDD.t113 39.6722
R409 VDD.n1818 VDD.n522 39.5509
R410 VDD.n1526 VDD.n734 39.5509
R411 VDD.n1806 VDD.n529 38.3019
R412 VDD.n791 VDD.t567 38.3019
R413 VDD.n1535 VDD.n726 38.3019
R414 VDD.n1757 VDD.n569 37.9019
R415 VDD.n1549 VDD.n1548 37.9019
R416 VDD.n459 VDD.t313 37.8856
R417 VDD.n448 VDD.t322 36.2203
R418 VDD.n1745 VDD.n577 35.8675
R419 VDD.n1557 VDD.n1556 35.8675
R420 VDD.n779 VDD.t591 35.804
R421 VDD.n866 VDD.t461 35.5682
R422 VDD.n318 VDD.t397 35.5071
R423 VDD.n28 VDD.t538 33.5535
R424 VDD.n114 VDD.t608 32.8941
R425 VDD.n2021 VDD.t800 32.8941
R426 VDD.n1225 VDD.t714 32.8322
R427 VDD.n1717 VDD.n1716 32.7175
R428 VDD.n1586 VDD.n625 32.7175
R429 VDD.n1806 VDD.n530 32.0571
R430 VDD.n1527 VDD.n726 32.0571
R431 VDD.n809 VDD.t231 31.6415
R432 VDD.n1840 VDD.t329 31.6408
R433 VDD.n1412 VDD.t598 31.2245
R434 VDD.n5 VDD.t104 31.1569
R435 VDD.n530 VDD.n522 30.8082
R436 VDD.n1527 VDD.n1526 30.8082
R437 VDD.n1213 VDD.n1179 30.0963
R438 VDD.n1177 VDD.n1168 28.8809
R439 VDD.t559 VDD.n759 28.7266
R440 VDD.n1846 VDD.t320 28.3102
R441 VDD.n1776 VDD.n1775 28.1746
R442 VDD.n1521 VDD.n736 28.1746
R443 VDD.n227 VDD.n116 26.1348
R444 VDD.n926 VDD.t261 24.6667
R445 VDD.n1224 VDD.n1223 24.6243
R446 VDD.n1370 VDD.t565 24.147
R447 VDD.n1987 VDD.t324 23.7307
R448 VDD.n1701 VDD.n1700 23.2342
R449 VDD.n2089 VDD.n2084 23.2342
R450 VDD.t324 VDD.n1986 22.0654
R451 VDD.t501 VDD.n1691 21.8883
R452 VDD.n1667 VDD.t332 21.8883
R453 VDD.n1602 VDD.t683 21.8883
R454 VDD.n701 VDD.t589 21.8883
R455 VDD.t811 VDD.n682 21.8883
R456 VDD.t34 VDD.n1088 21.8883
R457 VDD.t712 VDD.n1211 21.8883
R458 VDD.n1632 VDD.t131 21.8883
R459 VDD.n2102 VDD.t85 21.8883
R460 VDD.n792 VDD.t565 21.6491
R461 VDD.n1279 VDD.t182 21.2328
R462 VDD.t206 VDD.n1946 20.8165
R463 VDD.n1702 VDD.n1701 20.395
R464 VDD.n2089 VDD.n2085 20.3898
R465 VDD.n1063 VDD.t43 19.8363
R466 VDD.n88 VDD.n64 19.7184
R467 VDD.n203 VDD.n157 19.7184
R468 VDD.n332 VDD.n284 19.7184
R469 VDD.n392 VDD.n380 19.7184
R470 VDD.t243 VDD.n1818 19.5675
R471 VDD.t185 VDD.n734 19.5675
R472 VDD.n1121 VDD.n1120 19.0194
R473 VDD.n257 VDD.t277 18.5517
R474 VDD.n1242 VDD.n806 17.5593
R475 VDD.t320 VDD.n1845 17.4859
R476 VDD.n1402 VDD.t559 17.0696
R477 VDD.n1920 VDD.n1913 16.2393
R478 VDD.t598 VDD.n1411 14.5717
R479 VDD.t1 VDD.n98 14.5667
R480 VDD.t22 VDD.n275 14.5667
R481 VDD.n372 VDD.t306 14.5667
R482 VDD.n1852 VDD.t329 14.1554
R483 VDD.n1683 VDD.t487 13.6804
R484 VDD.t317 VDD.n1675 13.6804
R485 VDD.t668 VDD.n1609 13.6804
R486 VDD.n693 VDD.t570 13.6804
R487 VDD.n674 VDD.t819 13.6804
R488 VDD.n893 VDD.n841 13.6804
R489 VDD.n1113 VDD.t36 13.6804
R490 VDD.n1203 VDD.t710 13.6804
R491 VDD.t139 VDD.n1623 13.6804
R492 VDD.n2113 VDD.t106 13.6804
R493 VDD.n1817 VDD.n516 13.33
R494 VDD.n1434 VDD.n733 13.2637
R495 VDD.n865 VDD.n840 12.9964
R496 VDD.n956 VDD.n909 12.9964
R497 VDD.n2022 VDD.n2021 12.0091
R498 VDD.n2033 VDD.n114 12.0091
R499 VDD.n1821 VDD.n521 11.6418
R500 VDD.n1525 VDD.n735 11.6418
R501 VDD.n1765 VDD.n572 11.2373
R502 VDD.n1817 VDD.n523 11.2079
R503 VDD.n1528 VDD.n733 11.2079
R504 VDD.n1537 VDD.n724 11.1709
R505 VDD.n1274 VDD.n807 11.094
R506 VDD.n189 VDD.t527 10.9895
R507 VDD.n866 VDD.n864 10.9444
R508 VDD.n968 VDD.n967 10.9444
R509 VDD.t449 VDD.n888 10.9444
R510 VDD.n963 VDD.n905 10.9444
R511 VDD.n955 VDD.n910 10.9444
R512 VDD.n1059 VDD.t31 10.9444
R513 VDD.n1103 VDD.n1102 10.723
R514 VDD.n1661 VDD.n1660 10.7223
R515 VDD.n1594 VDD.n1593 10.7223
R516 VDD.n709 VDD.n708 10.7223
R517 VDD.n688 VDD.n687 10.7223
R518 VDD.n1615 VDD.n1614 10.7223
R519 VDD.n1913 VDD.n1887 10.4784
R520 VDD.n1282 VDD.n806 10.4784
R521 VDD.n1963 VDD.n1892 10.3407
R522 VDD.n1278 VDD.n800 10.3407
R523 VDD.n1786 VDD.n1785 10.2548
R524 VDD.n1486 VDD.n1485 10.2548
R525 VDD.n1274 VDD.n811 10.2279
R526 VDD.n1936 VDD.n1895 10.1865
R527 VDD.n1274 VDD.n1273 10.1865
R528 VDD.n1820 VDD.t188 9.99217
R529 VDD.n1377 VDD.t591 9.99217
R530 VDD.n740 VDD.t197 9.99217
R531 VDD.n1959 VDD.n1892 9.86137
R532 VDD.n1278 VDD.n807 9.86137
R533 VDD.n1776 VDD.n521 9.78981
R534 VDD.n1525 VDD.n736 9.78981
R535 VDD.n93 VDD.n92 9.68099
R536 VDD.n92 VDD.n83 9.68099
R537 VDD.n2044 VDD.n65 9.68099
R538 VDD.n2039 VDD.n66 9.68099
R539 VDD.n2039 VDD.n67 9.68099
R540 VDD.n203 VDD.n158 9.68099
R541 VDD.n199 VDD.n158 9.68099
R542 VDD.n208 VDD.n153 9.68099
R543 VDD.n208 VDD.n155 9.68099
R544 VDD.n195 VDD.n179 9.68099
R545 VDD.n195 VDD.n180 9.68099
R546 VDD.n322 VDD.n293 9.68099
R547 VDD.n322 VDD.n294 9.68099
R548 VDD.n327 VDD.n284 9.68099
R549 VDD.n327 VDD.n291 9.68099
R550 VDD.n336 VDD.n281 9.68099
R551 VDD.n336 VDD.n283 9.68099
R552 VDD.n409 VDD.n357 9.68099
R553 VDD.n413 VDD.n357 9.68099
R554 VDD.n387 VDD.n380 9.68099
R555 VDD.n387 VDD.n383 9.68099
R556 VDD.n399 VDD.n365 9.68099
R557 VDD.n395 VDD.n365 9.68099
R558 VDD.n2052 VDD.n2051 9.6468
R559 VDD.n1994 VDD.t322 9.57585
R560 VDD.n825 VDD.t181 9.55982
R561 VDD.n821 VDD.t240 9.55982
R562 VDD.n817 VDD.t228 9.55982
R563 VDD.n813 VDD.t230 9.55982
R564 VDD.n1915 VDD.t235 9.51591
R565 VDD.n1909 VDD.t205 9.51591
R566 VDD.n1902 VDD.t210 9.51591
R567 VDD.n1934 VDD.t193 9.51591
R568 VDD.n43 VDD.n42 9.4133
R569 VDD.n1966 VDD.n1887 9.28471
R570 VDD.n1282 VDD.n804 9.28471
R571 VDD.n1821 VDD.n519 9.24507
R572 VDD.n1437 VDD.n735 9.17659
R573 VDD.n1171 VDD.n1168 9.16567
R574 VDD.n2 VDD.n1 9.09976
R575 VDD.n728 VDD.n727 9.08576
R576 VDD.n6 VDD.t626 9.02932
R577 VDD.n1811 VDD.n1810 9.01945
R578 VDD.n981 VDD.n980 8.89243
R579 VDD.n45 VDD.n44 8.82188
R580 VDD.n1719 VDD.n581 8.80618
R581 VDD.n43 VDD.t549 8.79795
R582 VDD.n1804 VDD.n537 8.78029
R583 VDD.n1799 VDD.n1798 8.78029
R584 VDD.n1473 VDD.n1472 8.78029
R585 VDD.n1470 VDD.n1459 8.78029
R586 VDD.n1794 VDD.n1793 8.71327
R587 VDD.n1781 VDD.n1780 8.71327
R588 VDD.n1491 VDD.n1490 8.71327
R589 VDD.n1478 VDD.n1477 8.71327
R590 VDD.n6 VDD.t625 8.6005
R591 VDD.n7 VDD.t666 8.6005
R592 VDD.n8 VDD.t105 8.6005
R593 VDD.n1752 VDD.n575 8.59141
R594 VDD.n1756 VDD.n575 8.59141
R595 VDD.n1758 VDD.n1756 8.59141
R596 VDD.n1760 VDD.n1758 8.59141
R597 VDD.n1760 VDD.n571 8.59141
R598 VDD.n1765 VDD.n571 8.59141
R599 VDD.n1713 VDD.n1704 8.59141
R600 VDD.n1713 VDD.n1706 8.59141
R601 VDD.n1706 VDD.n566 8.59141
R602 VDD.n1770 VDD.n566 8.59141
R603 VDD.n1771 VDD.n1770 8.59141
R604 VDD.n1519 VDD.n1497 8.59141
R605 VDD.n1514 VDD.n1497 8.59141
R606 VDD.n1514 VDD.n1502 8.59141
R607 VDD.n1510 VDD.n1502 8.59141
R608 VDD.n1510 VDD.n1505 8.59141
R609 VDD.n1537 VDD.n721 8.59141
R610 VDD.n1546 VDD.n721 8.59141
R611 VDD.n1546 VDD.n719 8.59141
R612 VDD.n719 VDD.n717 8.59141
R613 VDD.n1552 VDD.n717 8.59141
R614 VDD.n1553 VDD.n1552 8.59141
R615 VDD.n1682 VDD.n1637 8.488
R616 VDD.n1686 VDD.n595 8.488
R617 VDD.n1690 VDD.n593 8.488
R618 VDD.n1673 VDD.n1646 8.488
R619 VDD.n1649 VDD.n1648 8.488
R620 VDD.n1668 VDD.n1656 8.488
R621 VDD.n1664 VDD.n1658 8.488
R622 VDD.n1595 VDD.n622 8.488
R623 VDD.n1600 VDD.n620 8.488
R624 VDD.n1604 VDD.n613 8.488
R625 VDD.n1607 VDD.n611 8.488
R626 VDD.n706 VDD.n640 8.488
R627 VDD.n702 VDD.n642 8.488
R628 VDD.n698 VDD.n649 8.488
R629 VDD.n694 VDD.n651 8.488
R630 VDD.n686 VDD.n685 8.488
R631 VDD.n681 VDD.n657 8.488
R632 VDD.n667 VDD.n660 8.488
R633 VDD.n676 VDD.n669 8.488
R634 VDD.n966 VDD.n965 8.488
R635 VDD.n957 VDD.n903 8.488
R636 VDD.n982 VDD.n838 8.488
R637 VDD.n969 VDD.n839 8.488
R638 VDD.n962 VDD.n886 8.488
R639 VDD.n954 VDD.n906 8.488
R640 VDD.n1097 VDD.n1096 8.488
R641 VDD.n1106 VDD.n1089 8.488
R642 VDD.n1110 VDD.n1087 8.488
R643 VDD.n1115 VDD.n1085 8.488
R644 VDD.n1041 VDD.n1040 8.488
R645 VDD.n1057 VDD.n1023 8.488
R646 VDD.n1058 VDD.n1019 8.488
R647 VDD.n1064 VDD.n1016 8.488
R648 VDD.n1038 VDD.n1025 8.488
R649 VDD.n1044 VDD.n1020 8.488
R650 VDD.n1061 VDD.n1060 8.488
R651 VDD.n1067 VDD.n1017 8.488
R652 VDD.n1206 VDD.n1190 8.488
R653 VDD.n1205 VDD.n1198 8.488
R654 VDD.n1617 VDD.n1616 8.488
R655 VDD.n1629 VDD.n604 8.488
R656 VDD.n1628 VDD.n1621 8.488
R657 VDD.n1716 VDD.n1715 8.48682
R658 VDD.n1775 VDD.n561 8.48682
R659 VDD.n1521 VDD.n1520 8.48682
R660 VDD.n1504 VDD.n625 8.48682
R661 VDD.n1210 VDD.n1188 8.4005
R662 VDD.n1722 VDD.n581 8.37664
R663 VDD.n1946 VDD.n1890 8.32689
R664 VDD.n1281 VDD.n1279 8.32689
R665 VDD.n1753 VDD.n577 8.31689
R666 VDD.n1556 VDD.n715 8.31615
R667 VDD.n1682 VDD.n1638 8.2255
R668 VDD.n1686 VDD.n1637 8.2255
R669 VDD.n1690 VDD.n595 8.2255
R670 VDD.n1694 VDD.n593 8.2255
R671 VDD.n1676 VDD.n1646 8.2255
R672 VDD.n1673 VDD.n1648 8.2255
R673 VDD.n1668 VDD.n1649 8.2255
R674 VDD.n1664 VDD.n1656 8.2255
R675 VDD.n1600 VDD.n622 8.2255
R676 VDD.n1604 VDD.n620 8.2255
R677 VDD.n1607 VDD.n613 8.2255
R678 VDD.n1610 VDD.n611 8.2255
R679 VDD.n706 VDD.n642 8.2255
R680 VDD.n702 VDD.n649 8.2255
R681 VDD.n698 VDD.n651 8.2255
R682 VDD.n694 VDD.n692 8.2255
R683 VDD.n685 VDD.n657 8.2255
R684 VDD.n681 VDD.n660 8.2255
R685 VDD.n676 VDD.n667 8.2255
R686 VDD.n673 VDD.n669 8.2255
R687 VDD.n965 VDD.n903 8.2255
R688 VDD.n957 VDD.n908 8.2255
R689 VDD.n858 VDD.n838 8.2255
R690 VDD.n982 VDD.n839 8.2255
R691 VDD.n969 VDD.n886 8.2255
R692 VDD.n962 VDD.n906 8.2255
R693 VDD.n954 VDD.n911 8.2255
R694 VDD.n1106 VDD.n1096 8.2255
R695 VDD.n1110 VDD.n1089 8.2255
R696 VDD.n1115 VDD.n1087 8.2255
R697 VDD.n1040 VDD.n1027 8.2255
R698 VDD.n1041 VDD.n1023 8.2255
R699 VDD.n1058 VDD.n1057 8.2255
R700 VDD.n1064 VDD.n1019 8.2255
R701 VDD.n1070 VDD.n1016 8.2255
R702 VDD.n1038 VDD.n1037 8.2255
R703 VDD.n1044 VDD.n1025 8.2255
R704 VDD.n1060 VDD.n1020 8.2255
R705 VDD.n1061 VDD.n1017 8.2255
R706 VDD.n1067 VDD.n1015 8.2255
R707 VDD.n1210 VDD.n1190 8.2255
R708 VDD.n1206 VDD.n1205 8.2255
R709 VDD.n1202 VDD.n1198 8.2255
R710 VDD.n1617 VDD.n603 8.2255
R711 VDD.n1633 VDD.n604 8.2255
R712 VDD.n1629 VDD.n1628 8.2255
R713 VDD.n1624 VDD.n1621 8.2255
R714 VDD.n2105 VDD.n2103 8.2255
R715 VDD.n895 VDD.n887 8.20843
R716 VDD.n1178 VDD.n1177 8.20843
R717 VDD.n1825 VDD.n519 8.14941
R718 VDD.n1825 VDD.n512 8.14941
R719 VDD.n1835 VDD.n512 8.14941
R720 VDD.n1835 VDD.n490 8.14941
R721 VDD.n1851 VDD.n490 8.14941
R722 VDD.n1851 VDD.n491 8.14941
R723 VDD.n1847 VDD.n491 8.14941
R724 VDD.n1847 VDD.n424 8.14941
R725 VDD.n2007 VDD.n424 8.14941
R726 VDD.n2007 VDD.n425 8.14941
R727 VDD.n2003 VDD.n425 8.14941
R728 VDD.n2003 VDD.n428 8.14941
R729 VDD.n440 VDD.n428 8.14941
R730 VDD.n1993 VDD.n440 8.14941
R731 VDD.n1993 VDD.n441 8.14941
R732 VDD.n1988 VDD.n441 8.14941
R733 VDD.n1988 VDD.n447 8.14941
R734 VDD.n460 VDD.n447 8.14941
R735 VDD.n1978 VDD.n460 8.14941
R736 VDD.n1978 VDD.n461 8.14941
R737 VDD.n1973 VDD.n461 8.14941
R738 VDD.n1973 VDD.n1878 8.14941
R739 VDD.n1891 VDD.n1878 8.14941
R740 VDD.n1963 VDD.n1891 8.14941
R741 VDD.n1289 VDD.n800 8.14941
R742 VDD.n1289 VDD.n798 8.14941
R743 VDD.n1293 VDD.n798 8.14941
R744 VDD.n1293 VDD.n787 8.14941
R745 VDD.n1306 VDD.n787 8.14941
R746 VDD.n1306 VDD.n788 8.14941
R747 VDD.n788 VDD.n778 8.14941
R748 VDD.n1371 VDD.n778 8.14941
R749 VDD.n1371 VDD.n773 8.14941
R750 VDD.n1376 VDD.n773 8.14941
R751 VDD.n1376 VDD.n767 8.14941
R752 VDD.n1387 VDD.n767 8.14941
R753 VDD.n1387 VDD.n765 8.14941
R754 VDD.n1392 VDD.n765 8.14941
R755 VDD.n1392 VDD.n757 8.14941
R756 VDD.n1404 VDD.n757 8.14941
R757 VDD.n1404 VDD.n755 8.14941
R758 VDD.n1409 VDD.n755 8.14941
R759 VDD.n1409 VDD.n747 8.14941
R760 VDD.n1421 VDD.n747 8.14941
R761 VDD.n1421 VDD.n745 8.14941
R762 VDD.n1425 VDD.n745 8.14941
R763 VDD.n1425 VDD.n738 8.14941
R764 VDD.n1437 VDD.n738 8.14941
R765 VDD.n979 VDD.n868 7.963
R766 VDD.n1980 VDD.t313 7.91057
R767 VDD.n1828 VDD.n516 7.89208
R768 VDD.n1828 VDD.n514 7.89208
R769 VDD.n1832 VDD.n514 7.89208
R770 VDD.n1832 VDD.n487 7.89208
R771 VDD.n1854 VDD.n487 7.89208
R772 VDD.n1854 VDD.n488 7.89208
R773 VDD.n1843 VDD.n488 7.89208
R774 VDD.n1843 VDD.n421 7.89208
R775 VDD.n2010 VDD.n421 7.89208
R776 VDD.n2010 VDD.n422 7.89208
R777 VDD.n433 VDD.n422 7.89208
R778 VDD.n2000 VDD.n433 7.89208
R779 VDD.n2000 VDD.n434 7.89208
R780 VDD.n1996 VDD.n434 7.89208
R781 VDD.n1996 VDD.n437 7.89208
R782 VDD.n452 VDD.n437 7.89208
R783 VDD.n1985 VDD.n452 7.89208
R784 VDD.n1985 VDD.n453 7.89208
R785 VDD.n1981 VDD.n453 7.89208
R786 VDD.n1981 VDD.n456 7.89208
R787 VDD.n1882 VDD.n456 7.89208
R788 VDD.n1970 VDD.n1882 7.89208
R789 VDD.n1970 VDD.n1883 7.89208
R790 VDD.n1966 VDD.n1883 7.89208
R791 VDD.n1286 VDD.n804 7.89208
R792 VDD.n1286 VDD.n797 7.89208
R793 VDD.n1297 VDD.n797 7.89208
R794 VDD.n1297 VDD.n790 7.89208
R795 VDD.n1303 VDD.n790 7.89208
R796 VDD.n1303 VDD.n795 7.89208
R797 VDD.n795 VDD.n781 7.89208
R798 VDD.n1368 VDD.n781 7.89208
R799 VDD.n1368 VDD.n772 7.89208
R800 VDD.n1380 VDD.n772 7.89208
R801 VDD.n1380 VDD.n770 7.89208
R802 VDD.n1384 VDD.n770 7.89208
R803 VDD.n1384 VDD.n763 7.89208
R804 VDD.n1396 VDD.n763 7.89208
R805 VDD.n1396 VDD.n760 7.89208
R806 VDD.n1401 VDD.n760 7.89208
R807 VDD.n1401 VDD.n753 7.89208
R808 VDD.n1413 VDD.n753 7.89208
R809 VDD.n1413 VDD.n750 7.89208
R810 VDD.n1418 VDD.n750 7.89208
R811 VDD.n1418 VDD.n743 7.89208
R812 VDD.n1429 VDD.n743 7.89208
R813 VDD.n1429 VDD.n741 7.89208
R814 VDD.n1434 VDD.n741 7.89208
R815 VDD.n862 VDD.n849 7.613
R816 VDD.n55 VDD.t550 7.58462
R817 VDD.n56 VDD.t558 7.58462
R818 VDD.n37 VDD.n23 7.58109
R819 VDD.n1226 VDD.n1166 7.5255
R820 VDD.n896 VDD.n895 7.52444
R821 VDD.n1304 VDD.t567 7.49426
R822 VDD.n1790 VDD.n1789 7.30582
R823 VDD.n1482 VDD.n1481 7.30582
R824 VDD.n1530 VDD.n732 7.30582
R825 VDD.n26 VDD.t539 7.19043
R826 VDD.n3 VDD.t122 7.19043
R827 VDD.n966 VDD.n902 7.1755
R828 VDD.n1119 VDD.n1085 7.1755
R829 VDD.n868 VDD.n867 7.088
R830 VDD.n1919 VDD.n1911 7.00704
R831 VDD.n1923 VDD.n1911 7.00704
R832 VDD.n1924 VDD.n1923 7.00704
R833 VDD.n1925 VDD.n1924 7.00704
R834 VDD.n1925 VDD.n1908 7.00704
R835 VDD.n1930 VDD.n1908 7.00704
R836 VDD.n1930 VDD.n1899 7.00704
R837 VDD.n1953 VDD.n1899 7.00704
R838 VDD.n1953 VDD.n1900 7.00704
R839 VDD.n1948 VDD.n1900 7.00704
R840 VDD.n1948 VDD.n1904 7.00704
R841 VDD.n1943 VDD.n1904 7.00704
R842 VDD.n1943 VDD.n1933 7.00704
R843 VDD.n1938 VDD.n1933 7.00704
R844 VDD.n1938 VDD.n1936 7.00704
R845 VDD.n1271 VDD.n812 7.00704
R846 VDD.n1266 VDD.n1265 7.00704
R847 VDD.n1263 VDD.n816 7.00704
R848 VDD.n1258 VDD.n1257 7.00704
R849 VDD.n1255 VDD.n820 7.00704
R850 VDD.n1250 VDD.n1249 7.00704
R851 VDD.n1247 VDD.n824 7.00704
R852 VDD.n145 VDD.t369 6.94485
R853 VDD.n272 VDD.t376 6.94485
R854 VDD.n557 VDD.n555 6.94485
R855 VDD.n1443 VDD.t160 6.94485
R856 VDD.t461 VDD.n865 6.84045
R857 VDD.n956 VDD.t445 6.84045
R858 VDD.t45 VDD.n1026 6.84045
R859 VDD.n1225 VDD.n1224 6.84045
R860 VDD.n1644 VDD.n1643 6.70224
R861 VDD.n1641 VDD.n1639 6.70224
R862 VDD.n671 VDD.t826 6.70224
R863 VDD.n652 VDD.t605 6.70224
R864 VDD.n913 VDD.t446 6.70224
R865 VDD.n852 VDD.n851 6.70224
R866 VDD.n1082 VDD.t60 6.70224
R867 VDD.n1030 VDD.n1028 6.70224
R868 VDD.n1033 VDD.n1032 6.70224
R869 VDD.n1200 VDD.t711 6.70224
R870 VDD.n609 VDD.t696 6.70224
R871 VDD.n1622 VDD.t140 6.70224
R872 VDD.n2110 VDD.n2109 6.70224
R873 VDD.n591 VDD.t484 6.68489
R874 VDD.n712 VDD.n710 6.68371
R875 VDD.n225 VDD.t769 6.68267
R876 VDD.n1659 VDD.t352 6.65503
R877 VDD.n655 VDD.n653 6.65503
R878 VDD.n941 VDD.t636 6.65503
R879 VDD.n855 VDD.n853 6.65503
R880 VDD.n1100 VDD.n1098 6.65503
R881 VDD.n997 VDD.t44 6.65503
R882 VDD.n1174 VDD.n1172 6.65503
R883 VDD.n1592 VDD.n1591 6.65503
R884 VDD.n608 VDD.n607 6.65503
R885 VDD.n2085 VDD.t119 6.65503
R886 VDD.n1075 VDD.t620 6.64521
R887 VDD.n1809 VDD.n1808 6.63561
R888 VDD.n2029 VDD.n2028 6.61305
R889 VDD.n230 VDD.n229 6.58706
R890 VDD.n1530 VDD.n1529 6.56859
R891 VDD.n2027 VDD.t442 6.54616
R892 VDD.n2027 VDD.t418 6.54616
R893 VDD.n253 VDD.t396 6.52811
R894 VDD.n233 VDD.n232 6.52199
R895 VDD.n2030 VDD.n2025 6.51831
R896 VDD.t204 VDD.n1498 6.50716
R897 VDD.n563 VDD.t214 6.50716
R898 VDD.n51 VDD.n50 6.44895
R899 VDD.n1456 VDD.t184 6.43191
R900 VDD.n113 VDD.t610 6.43137
R901 VDD.n316 VDD.t772 6.43137
R902 VDD.n2020 VDD.t805 6.43137
R903 VDD.n1442 VDD.t223 6.43124
R904 VDD.n1465 VDD.t196 6.4298
R905 VDD.n538 VDD.t187 6.42961
R906 VDD.n546 VDD.t242 6.37351
R907 VDD.n1446 VDD.t237 6.37275
R908 VDD.n553 VDD.t199 6.37256
R909 VDD.n559 VDD.t208 6.37217
R910 VDD.n573 VDD.t220 6.36486
R911 VDD.n1748 VDD.t233 6.36262
R912 VDD.n1708 VDD.t217 6.36128
R913 VDD.n1541 VDD.t215 6.30795
R914 VDD.n722 VDD.t225 6.30193
R915 VDD.n101 VDD.n100 6.3005
R916 VDD.n174 VDD.n173 6.3005
R917 VDD VDD.n189 6.3005
R918 VDD.n213 VDD.n147 6.3005
R919 VDD.n120 VDD.n119 6.3005
R920 VDD.n304 VDD.n303 6.3005
R921 VDD.n256 VDD.n255 6.3005
R922 VDD VDD.n257 6.3005
R923 VDD.n341 VDD.n275 6.3005
R924 VDD VDD.n316 6.3005
R925 VDD.n403 VDD.n402 6.3005
R926 VDD.n892 VDD.n891 6.3005
R927 VDD.n893 VDD.n892 6.3005
R928 VDD.n898 VDD.n897 6.3005
R929 VDD.n897 VDD.n896 6.3005
R930 VDD.n862 VDD.n861 6.3005
R931 VDD.n863 VDD.n862 6.3005
R932 VDD.n1119 VDD.n1118 6.3005
R933 VDD.n1120 VDD.n1119 6.3005
R934 VDD.n1170 VDD.n1169 6.3005
R935 VDD.n1188 VDD.n1187 6.3005
R936 VDD.n1212 VDD.n1188 6.3005
R937 VDD.n1227 VDD.n1226 6.3005
R938 VDD.n1226 VDD.n1225 6.3005
R939 VDD.n1167 VDD.n1165 6.3005
R940 VDD.n1224 VDD.n1167 6.3005
R941 VDD.n1215 VDD.n1214 6.3005
R942 VDD.n1214 VDD.n1213 6.3005
R943 VDD.n373 VDD.n372 6.3005
R944 VDD.n2020 VDD 6.3005
R945 VDD VDD.n113 6.3005
R946 VDD.n98 VDD.n97 6.3005
R947 VDD.n10 VDD.n5 6.3005
R948 VDD.n11 VDD.n4 6.3005
R949 VDD.n12 VDD.n3 6.3005
R950 VDD.n14 VDD.n13 6.3005
R951 VDD.n30 VDD.n29 6.3005
R952 VDD.n31 VDD.n28 6.3005
R953 VDD.n32 VDD.n27 6.3005
R954 VDD.n33 VDD.n26 6.3005
R955 VDD.n34 VDD.n25 6.3005
R956 VDD.n35 VDD.n24 6.3005
R957 VDD.n2070 VDD.n2060 6.3005
R958 VDD VDD.n2061 6.3005
R959 VDD.n2069 VDD.n2062 6.3005
R960 VDD.n2124 VDD.n2123 6.3005
R961 VDD.n2126 VDD.n2125 6.3005
R962 VDD.n2128 VDD.n2127 6.3005
R963 VDD.n1506 VDD.t190 6.29942
R964 VDD.n563 VDD.t212 6.29685
R965 VDD.n46 VDD.t555 6.27989
R966 VDD.n1075 VDD.t618 6.26273
R967 VDD.n712 VDD.n711 6.24167
R968 VDD.n145 VDD.t748 6.2405
R969 VDD.n272 VDD.t284 6.2405
R970 VDD.n557 VDD.n556 6.2405
R971 VDD.n591 VDD.t517 6.2405
R972 VDD.n1659 VDD.t328 6.2405
R973 VDD.n1644 VDD.n1642 6.2405
R974 VDD.n1641 VDD.n1640 6.2405
R975 VDD.n1499 VDD.t204 6.2405
R976 VDD.n1443 VDD.t173 6.2405
R977 VDD.n671 VDD.t820 6.2405
R978 VDD.n655 VDD.n654 6.2405
R979 VDD.n652 VDD.t571 6.2405
R980 VDD.n913 VDD.t464 6.2405
R981 VDD.n941 VDD.t638 6.2405
R982 VDD.n855 VDD.n854 6.2405
R983 VDD.n852 VDD.n850 6.2405
R984 VDD.n1100 VDD.n1099 6.2405
R985 VDD.n1082 VDD.t37 6.2405
R986 VDD.n1033 VDD.n1031 6.2405
R987 VDD.n1030 VDD.n1029 6.2405
R988 VDD.n997 VDD.t52 6.2405
R989 VDD.n1200 VDD.t717 6.2405
R990 VDD.n1174 VDD.n1173 6.2405
R991 VDD.n1592 VDD.n1590 6.2405
R992 VDD.n609 VDD.t669 6.2405
R993 VDD.n608 VDD.n606 6.2405
R994 VDD.n1622 VDD.t143 6.2405
R995 VDD.t214 VDD.n562 6.2405
R996 VDD.n2085 VDD.t114 6.2405
R997 VDD.n2110 VDD.n2108 6.2405
R998 VDD.n1498 VDD.t202 6.23498
R999 VDD.n863 VDD.n848 6.15645
R1000 VDD.n1529 VDD.n727 6.03524
R1001 VDD.n1810 VDD.n1809 5.96892
R1002 VDD.n934 VDD.n933 5.77744
R1003 VDD.n923 VDD.n922 5.77744
R1004 VDD.n1139 VDD.t645 5.77744
R1005 VDD.n1134 VDD.t456 5.77744
R1006 VDD.n2066 VDD.n2065 5.77744
R1007 VDD.n2119 VDD.t294 5.77744
R1008 VDD.n897 VDD.n892 5.7755
R1009 VDD.n20 VDD.n19 5.7405
R1010 VDD.n104 VDD.n103 5.72051
R1011 VDD.n177 VDD.n176 5.72051
R1012 VDD.n307 VDD.n306 5.72032
R1013 VDD.n406 VDD.n405 5.72032
R1014 VDD.n1122 VDD.n1121 5.2962
R1015 VDD.n278 VDD.t784 5.20342
R1016 VDD.n369 VDD.t310 5.20342
R1017 VDD.n78 VDD.t481 5.20242
R1018 VDD.n150 VDD.t12 5.20242
R1019 VDD.n22 VDD.n16 5.2005
R1020 VDD.n21 VDD.n17 5.2005
R1021 VDD.n20 VDD.n18 5.2005
R1022 VDD.n75 VDD.t24 5.17246
R1023 VDD.n146 VDD.t362 5.17246
R1024 VDD.n274 VDD.t764 5.17246
R1025 VDD.n371 VDD.t476 5.17246
R1026 VDD.n73 VDD.n72 5.107
R1027 VDD.n171 VDD.n170 5.107
R1028 VDD.n300 VDD.n299 5.107
R1029 VDD.n364 VDD.n363 5.107
R1030 VDD.n1809 VDD.n523 5.10682
R1031 VDD.n1529 VDD.n1528 5.10682
R1032 VDD.n924 VDD.t452 5.07264
R1033 VDD.n1141 VDD.n1140 5.07264
R1034 VDD.n1136 VDD.n1135 5.07264
R1035 VDD.n2067 VDD.t115 5.07264
R1036 VDD.n2121 VDD.n2120 5.07264
R1037 VDD.n231 VDD.n116 5.0405
R1038 VDD.n1956 VDD.t194 4.99634
R1039 VDD.n190 VDD.t526 4.92985
R1040 VDD.n317 VDD.t398 4.92985
R1041 VDD.n348 VDD.t801 4.92985
R1042 VDD.n115 VDD.t760 4.92985
R1043 VDD.n938 VDD.t649 4.79075
R1044 VDD.n864 VDD.n863 4.78846
R1045 VDD.n1222 VDD.n1180 4.7255
R1046 VDD.n103 VDD.t762 4.64447
R1047 VDD.n176 VDD.t657 4.64447
R1048 VDD.n306 VDD.t400 4.64447
R1049 VDD.n405 VDD.t796 4.64447
R1050 VDD.n95 VDD.n80 4.60311
R1051 VDD.n181 VDD.t655 4.60311
R1052 VDD.n211 VDD.n152 4.60311
R1053 VDD.n339 VDD.n280 4.60311
R1054 VDD.n308 VDD.t71 4.60311
R1055 VDD.n375 VDD.n366 4.60311
R1056 VDD.n407 VDD.t381 4.60311
R1057 VDD.n105 VDD.t81 4.60311
R1058 VDD.n949 VDD.n916 4.52789
R1059 VDD.n1218 VDD.n1217 4.52785
R1060 VDD.n847 VDD.n832 4.51855
R1061 VDD.n1122 VDD.n1081 4.5152
R1062 VDD.n973 VDD.n972 4.5084
R1063 VDD.n1011 VDD.n1010 4.50489
R1064 VDD.n948 VDD.n947 4.5005
R1065 VDD.n946 VDD.n917 4.5005
R1066 VDD.n942 VDD.n915 4.5005
R1067 VDD.n916 VDD.n907 4.5005
R1068 VDD.n952 VDD.n912 4.5005
R1069 VDD.n901 VDD.n900 4.5005
R1070 VDD.n902 VDD.n901 4.5005
R1071 VDD.n902 VDD.n887 4.5005
R1072 VDD.n985 VDD.n984 4.5005
R1073 VDD.n978 VDD.n977 4.5005
R1074 VDD.n979 VDD.n978 4.5005
R1075 VDD.n980 VDD.n979 4.5005
R1076 VDD.n867 VDD.n847 4.5005
R1077 VDD.n867 VDD.n866 4.5005
R1078 VDD.n844 VDD.n834 4.5005
R1079 VDD.n988 VDD.n987 4.5005
R1080 VDD.n974 VDD.n871 4.5005
R1081 VDD.n976 VDD.n975 4.5005
R1082 VDD.n986 VDD.n833 4.5005
R1083 VDD.n1126 VDD.n1080 4.5005
R1084 VDD.n1127 VDD.n1079 4.5005
R1085 VDD.n1011 VDD.n1000 4.5005
R1086 VDD.n1014 VDD.n1001 4.5005
R1087 VDD.n1072 VDD.n1071 4.5005
R1088 VDD.n1073 VDD.n1072 4.5005
R1089 VDD.n1014 VDD.n1013 4.5005
R1090 VDD.n1007 VDD.n1002 4.5005
R1091 VDD.n1004 VDD.n1003 4.5005
R1092 VDD.n995 VDD.n994 4.5005
R1093 VDD.n1009 VDD.n1008 4.5005
R1094 VDD.n1159 VDD.n1158 4.5005
R1095 VDD.n1153 VDD.n1152 4.5005
R1096 VDD.n1154 VDD.n992 4.5005
R1097 VDD.n1157 VDD.n991 4.5005
R1098 VDD.n1217 VDD.n1216 4.5005
R1099 VDD.n1216 VDD.n1180 4.5005
R1100 VDD.n1180 VDD.n1179 4.5005
R1101 VDD.n1186 VDD.n1183 4.5005
R1102 VDD.n1221 VDD.n1220 4.5005
R1103 VDD.n1222 VDD.n1221 4.5005
R1104 VDD.n1223 VDD.n1222 4.5005
R1105 VDD.n1185 VDD.n1182 4.5005
R1106 VDD.n1184 VDD.n1163 4.5005
R1107 VDD.n1229 VDD.n1228 4.5005
R1108 VDD.n1233 VDD.n1232 4.5005
R1109 VDD.n1170 VDD.n830 4.5005
R1110 VDD.n1170 VDD.n1166 4.5005
R1111 VDD.n1178 VDD.n1166 4.5005
R1112 VDD.n831 VDD.n829 4.5005
R1113 VDD.n2017 VDD.n2016 4.5005
R1114 VDD.n54 VDD.n53 4.5005
R1115 VDD.n75 VDD.t23 4.2255
R1116 VDD.n190 VDD.t531 4.2255
R1117 VDD.n146 VDD.t364 4.2255
R1118 VDD.n274 VDD.t763 4.2255
R1119 VDD.n317 VDD.t778 4.2255
R1120 VDD.n371 VDD.t475 4.2255
R1121 VDD.n348 VDD.t810 4.2255
R1122 VDD.n115 VDD.t609 4.2255
R1123 VDD.n1685 VDD.t508 4.10447
R1124 VDD.t315 VDD.n1647 4.10447
R1125 VDD.t677 VDD.n612 4.10447
R1126 VDD.t577 VDD.n699 4.10447
R1127 VDD.n670 VDD.t813 4.10447
R1128 VDD.n1112 VDD.t38 4.10447
R1129 VDD.n1197 VDD.t707 4.10447
R1130 VDD.t136 VDD.n1630 4.10447
R1131 VDD.n2095 VDD.t111 4.10447
R1132 VDD.n242 VDD.n241 3.99669
R1133 VDD.n125 VDD.n124 3.99665
R1134 VDD.n241 VDD.t444 3.80383
R1135 VDD.n124 VDD.t416 3.80304
R1136 VDD.n1819 VDD.n517 3.74738
R1137 VDD.n1827 VDD.n1826 3.74738
R1138 VDD.n518 VDD.n513 3.74738
R1139 VDD.t336 VDD.n1833 3.74738
R1140 VDD.n1834 VDD.n489 3.74738
R1141 VDD.n1853 VDD.n1852 3.74738
R1142 VDD.n1841 VDD.n1840 3.74738
R1143 VDD.n1846 VDD.n1844 3.74738
R1144 VDD.n1845 VDD.n423 3.74738
R1145 VDD.n2009 VDD.n2008 3.74738
R1146 VDD.n430 VDD.n429 3.74738
R1147 VDD.n2002 VDD.n431 3.74738
R1148 VDD.n2001 VDD.n432 3.74738
R1149 VDD.n439 VDD.n438 3.74738
R1150 VDD.n1995 VDD.n1994 3.74738
R1151 VDD.n449 VDD.n448 3.74738
R1152 VDD.n1987 VDD.n450 3.74738
R1153 VDD.n1986 VDD.n451 3.74738
R1154 VDD.n459 VDD.n458 3.74738
R1155 VDD.n1980 VDD.n1979 3.74738
R1156 VDD.n1879 VDD.n457 3.74738
R1157 VDD.n1972 VDD.n1880 3.74738
R1158 VDD.n1971 VDD.n1881 3.74738
R1159 VDD.n1889 VDD.n1888 3.74738
R1160 VDD.n1965 VDD.n1964 3.74738
R1161 VDD.n1280 VDD.n801 3.74738
R1162 VDD.n1288 VDD.n1287 3.74738
R1163 VDD.n803 VDD.n802 3.74738
R1164 VDD.n1296 VDD.n1294 3.74738
R1165 VDD.n1295 VDD.n789 3.74738
R1166 VDD.n1305 VDD.n1304 3.74738
R1167 VDD.n794 VDD.n791 3.74738
R1168 VDD.n793 VDD.n792 3.74738
R1169 VDD.n1370 VDD.n1369 3.74738
R1170 VDD.n780 VDD.n779 3.74738
R1171 VDD.n1379 VDD.n1377 3.74738
R1172 VDD.n1378 VDD.n768 3.74738
R1173 VDD.n1386 VDD.n1385 3.74738
R1174 VDD.n769 VDD.n764 3.74738
R1175 VDD.n1395 VDD.n1393 3.74738
R1176 VDD.n1394 VDD.n758 3.74738
R1177 VDD.n1403 VDD.n1402 3.74738
R1178 VDD.n759 VDD.n754 3.74738
R1179 VDD.n1412 VDD.n1410 3.74738
R1180 VDD.n1411 VDD.n748 3.74738
R1181 VDD.n1420 VDD.n1419 3.74738
R1182 VDD.n749 VDD.n744 3.74738
R1183 VDD.n1428 VDD.n1426 3.74738
R1184 VDD.n1427 VDD.n739 3.74738
R1185 VDD.n1436 VDD.n1435 3.74738
R1186 VDD.n134 VDD.t749 3.6405
R1187 VDD.n134 VDD.n133 3.6405
R1188 VDD.n136 VDD.t436 3.6405
R1189 VDD.n136 VDD.n135 3.6405
R1190 VDD.n138 VDD.t438 3.6405
R1191 VDD.n138 VDD.n137 3.6405
R1192 VDD.n140 VDD.t440 3.6405
R1193 VDD.n140 VDD.n139 3.6405
R1194 VDD.n132 VDD.t750 3.6405
R1195 VDD.n132 VDD.n131 3.6405
R1196 VDD.n129 VDD.t751 3.6405
R1197 VDD.n129 VDD.n128 3.6405
R1198 VDD.n127 VDD.t747 3.6405
R1199 VDD.n127 VDD.n126 3.6405
R1200 VDD.n122 VDD.t745 3.6405
R1201 VDD.n122 VDD.n121 3.6405
R1202 VDD.n118 VDD.t249 3.6405
R1203 VDD.n118 VDD.n117 3.6405
R1204 VDD.n252 VDD.t65 3.6405
R1205 VDD.n252 VDD.n251 3.6405
R1206 VDD.n239 VDD.t267 3.6405
R1207 VDD.n239 VDD.n238 3.6405
R1208 VDD.n237 VDD.t273 3.6405
R1209 VDD.n237 VDD.n236 3.6405
R1210 VDD.n249 VDD.t271 3.6405
R1211 VDD.n249 VDD.n248 3.6405
R1212 VDD.n247 VDD.t265 3.6405
R1213 VDD.n247 VDD.n246 3.6405
R1214 VDD.n269 VDD.t269 3.6405
R1215 VDD.n269 VDD.n268 3.6405
R1216 VDD.n261 VDD.t401 3.6405
R1217 VDD.n261 VDD.n260 3.6405
R1218 VDD.n265 VDD.t407 3.6405
R1219 VDD.n265 VDD.n264 3.6405
R1220 VDD.n263 VDD.t419 3.6405
R1221 VDD.n263 VDD.n262 3.6405
R1222 VDD.n1859 VDD.t504 3.6405
R1223 VDD.n1859 VDD.n1858 3.6405
R1224 VDD.n496 VDD.t520 3.6405
R1225 VDD.n496 VDD.n495 3.6405
R1226 VDD.n480 VDD.t505 3.6405
R1227 VDD.n480 VDD.n479 3.6405
R1228 VDD.n477 VDD.t360 3.6405
R1229 VDD.n477 VDD.n476 3.6405
R1230 VDD.n474 VDD.t511 3.6405
R1231 VDD.n474 VDD.n473 3.6405
R1232 VDD.n502 VDD.t491 3.6405
R1233 VDD.n502 VDD.n501 3.6405
R1234 VDD.n1871 VDD.t314 3.6405
R1235 VDD.n1871 VDD.n1870 3.6405
R1236 VDD.n1868 VDD.t343 3.6405
R1237 VDD.n1868 VDD.n1867 3.6405
R1238 VDD.n465 VDD.t490 3.6405
R1239 VDD.n465 VDD.n464 3.6405
R1240 VDD.n544 VDD.t178 3.6405
R1241 VDD.n544 VDD.n543 3.6405
R1242 VDD.n542 VDD.t163 3.6405
R1243 VDD.n542 VDD.n541 3.6405
R1244 VDD.n550 VDD.t168 3.6405
R1245 VDD.n550 VDD.n549 3.6405
R1246 VDD.n548 VDD.t179 3.6405
R1247 VDD.n548 VDD.n547 3.6405
R1248 VDD.n1699 VDD.t509 3.6405
R1249 VDD.n1699 VDD.n1698 3.6405
R1250 VDD.n1697 VDD.t514 3.6405
R1251 VDD.n1697 VDD.n1696 3.6405
R1252 VDD.n1651 VDD.t316 3.6405
R1253 VDD.n1651 VDD.n1650 3.6405
R1254 VDD.n1653 VDD.t344 3.6405
R1255 VDD.n1653 VDD.n1652 3.6405
R1256 VDD.n1461 VDD.t167 3.6405
R1257 VDD.n1461 VDD.n1460 3.6405
R1258 VDD.n1463 VDD.t148 3.6405
R1259 VDD.n1463 VDD.n1462 3.6405
R1260 VDD.n1450 VDD.t164 3.6405
R1261 VDD.n1450 VDD.n1449 3.6405
R1262 VDD.n1452 VDD.t180 3.6405
R1263 VDD.n1452 VDD.n1451 3.6405
R1264 VDD.n1340 VDD.t606 3.6405
R1265 VDD.n1340 VDD.n1339 3.6405
R1266 VDD.n1326 VDD.t604 3.6405
R1267 VDD.n1326 VDD.n1325 3.6405
R1268 VDD.n1328 VDD.t576 3.6405
R1269 VDD.n1328 VDD.n1327 3.6405
R1270 VDD.n1334 VDD.t667 3.6405
R1271 VDD.n1334 VDD.n1333 3.6405
R1272 VDD.n1337 VDD.t682 3.6405
R1273 VDD.n1337 VDD.n1336 3.6405
R1274 VDD.n1322 VDD.t599 3.6405
R1275 VDD.n1322 VDD.n1321 3.6405
R1276 VDD.n665 VDD.t812 3.6405
R1277 VDD.n665 VDD.n664 3.6405
R1278 VDD.n663 VDD.t823 3.6405
R1279 VDD.n663 VDD.n662 3.6405
R1280 VDD.n646 VDD.t602 3.6405
R1281 VDD.n646 VDD.n645 3.6405
R1282 VDD.n644 VDD.t590 3.6405
R1283 VDD.n644 VDD.n643 3.6405
R1284 VDD.n1330 VDD.t702 3.6405
R1285 VDD.n1330 VDD.n1329 3.6405
R1286 VDD.n1363 VDD.t685 3.6405
R1287 VDD.n1363 VDD.n1362 3.6405
R1288 VDD.n1358 VDD.t581 3.6405
R1289 VDD.n1358 VDD.n1357 3.6405
R1290 VDD.n1352 VDD.t695 3.6405
R1291 VDD.n1352 VDD.n1351 3.6405
R1292 VDD.n1355 VDD.t672 3.6405
R1293 VDD.n1355 VDD.n1354 3.6405
R1294 VDD.n1310 VDD.t603 3.6405
R1295 VDD.n1310 VDD.n1309 3.6405
R1296 VDD.n1315 VDD.t566 3.6405
R1297 VDD.n1315 VDD.n1314 3.6405
R1298 VDD.n1313 VDD.t584 3.6405
R1299 VDD.n1313 VDD.n1312 3.6405
R1300 VDD.n1319 VDD.t706 3.6405
R1301 VDD.n1319 VDD.n1318 3.6405
R1302 VDD.n775 VDD.t699 3.6405
R1303 VDD.n775 VDD.n774 3.6405
R1304 VDD.n878 VDD.t460 3.6405
R1305 VDD.n878 VDD.n877 3.6405
R1306 VDD.n876 VDD.t470 3.6405
R1307 VDD.n876 VDD.n875 3.6405
R1308 VDD.n882 VDD.t637 3.6405
R1309 VDD.n882 VDD.n881 3.6405
R1310 VDD.n884 VDD.t631 3.6405
R1311 VDD.n884 VDD.n883 3.6405
R1312 VDD.n1093 VDD.t35 3.6405
R1313 VDD.n1093 VDD.n1092 3.6405
R1314 VDD.n1091 VDD.t53 3.6405
R1315 VDD.n1091 VDD.n1090 3.6405
R1316 VDD.n1052 VDD.t619 3.6405
R1317 VDD.n1052 VDD.n1051 3.6405
R1318 VDD.n1054 VDD.t615 3.6405
R1319 VDD.n1054 VDD.n1053 3.6405
R1320 VDD.n1049 VDD.t51 3.6405
R1321 VDD.n1049 VDD.n1048 3.6405
R1322 VDD.n1047 VDD.t42 3.6405
R1323 VDD.n1047 VDD.n1046 3.6405
R1324 VDD.n1194 VDD.t713 3.6405
R1325 VDD.n1194 VDD.n1193 3.6405
R1326 VDD.n1192 VDD.t722 3.6405
R1327 VDD.n1192 VDD.n1191 3.6405
R1328 VDD.n615 VDD.t705 3.6405
R1329 VDD.n615 VDD.n614 3.6405
R1330 VDD.n617 VDD.t684 3.6405
R1331 VDD.n617 VDD.n616 3.6405
R1332 VDD.n598 VDD.t144 3.6405
R1333 VDD.n598 VDD.n597 3.6405
R1334 VDD.n600 VDD.t132 3.6405
R1335 VDD.n600 VDD.n599 3.6405
R1336 VDD.n1875 VDD.t496 3.6405
R1337 VDD.n1875 VDD.n1874 3.6405
R1338 VDD.n444 VDD.t335 3.6405
R1339 VDD.n444 VDD.n443 3.6405
R1340 VDD.n499 VDD.t321 3.6405
R1341 VDD.n499 VDD.n498 3.6405
R1342 VDD.n509 VDD.t510 3.6405
R1343 VDD.n509 VDD.n508 3.6405
R1344 VDD.n483 VDD.t355 3.6405
R1345 VDD.n483 VDD.n482 3.6405
R1346 VDD.n493 VDD.t337 3.6405
R1347 VDD.n493 VDD.n492 3.6405
R1348 VDD.n471 VDD.t323 3.6405
R1349 VDD.n471 VDD.n470 3.6405
R1350 VDD.n2081 VDD.t112 3.6405
R1351 VDD.n2081 VDD.n2080 3.6405
R1352 VDD.n2083 VDD.t118 3.6405
R1353 VDD.n2083 VDD.n2082 3.6405
R1354 VDD.n279 VDD.n278 3.60762
R1355 VDD.n370 VDD.n369 3.60762
R1356 VDD.n79 VDD.n78 3.60724
R1357 VDD.n151 VDD.n150 3.60724
R1358 VDD.n141 VDD.n140 3.54622
R1359 VDD.n266 VDD.n265 3.54622
R1360 VDD.n896 VDD.t459 3.42047
R1361 VDD.n2035 VDD.n114 3.35291
R1362 VDD.n2021 VDD.n350 3.35291
R1363 VDD.n429 VDD.t338 3.33106
R1364 VDD.n1238 VDD.n1236 3.32815
R1365 VDD.n187 VDD.n186 3.30485
R1366 VDD.n314 VDD.n311 3.30485
R1367 VDD.n355 VDD.n352 3.30485
R1368 VDD.n545 VDD.n542 3.30485
R1369 VDD.n551 VDD.n548 3.30485
R1370 VDD.n1464 VDD.n1463 3.30485
R1371 VDD.n1453 VDD.n1452 3.30485
R1372 VDD.n111 VDD.n110 3.30485
R1373 VDD.n1493 VDD.n736 3.28454
R1374 VDD.n1758 VDD.n1757 3.2486
R1375 VDD.n1549 VDD.n719 3.2486
R1376 VDD.n1915 VDD.t236 3.22394
R1377 VDD.n1909 VDD.t207 3.22394
R1378 VDD.n1902 VDD.t211 3.22394
R1379 VDD.n1934 VDD.t195 3.22394
R1380 VDD.n825 VDD.t183 3.22347
R1381 VDD.n821 VDD.t241 3.22347
R1382 VDD.n817 VDD.t229 3.22347
R1383 VDD.n813 VDD.t232 3.22347
R1384 VDD.n1446 VDD.t239 3.21802
R1385 VDD.n553 VDD.t201 3.21788
R1386 VDD.n538 VDD.t189 3.21785
R1387 VDD.n1442 VDD.t224 3.21781
R1388 VDD.n559 VDD.t209 3.21767
R1389 VDD.n1465 VDD.t198 3.21766
R1390 VDD.n1777 VDD.n1776 3.21752
R1391 VDD.n1456 VDD.t186 3.21671
R1392 VDD.n546 VDD.t244 3.21657
R1393 VDD.n55 VDD.n54 3.21512
R1394 VDD.n241 VDD.n240 3.20353
R1395 VDD.n124 VDD.n123 3.20342
R1396 VDD.n1541 VDD.t216 3.19864
R1397 VDD.n1506 VDD.t192 3.19113
R1398 VDD.n1708 VDD.t219 3.19113
R1399 VDD.n1748 VDD.t234 3.18927
R1400 VDD.n573 VDD.t222 3.1878
R1401 VDD.n722 VDD.t227 3.1878
R1402 VDD.n1275 VDD.n1274 3.16769
R1403 VDD.n1895 VDD.n1894 3.16769
R1404 VDD.n57 VDD.n56 3.16326
R1405 VDD.n47 VDD.n46 3.15744
R1406 VDD.n929 VDD.n928 3.15287
R1407 VDD VDD.n927 3.15287
R1408 VDD.n1147 VDD.n1145 3.15287
R1409 VDD.n1149 VDD.n1148 3.15287
R1410 VDD.n1144 VDD.n1143 3.15287
R1411 VDD VDD.n2026 3.15269
R1412 VDD.n1813 VDD.n525 3.15151
R1413 VDD.n182 VDD.n179 3.1505
R1414 VDD.n197 VDD.n179 3.1505
R1415 VDD.n195 VDD.n194 3.1505
R1416 VDD.n196 VDD.n195 3.1505
R1417 VDD.n193 VDD.n180 3.1505
R1418 VDD.n188 VDD.n180 3.1505
R1419 VDD.n210 VDD.n153 3.1505
R1420 VDD.n156 VDD.n153 3.1505
R1421 VDD.n209 VDD.n208 3.1505
R1422 VDD.n208 VDD.n207 3.1505
R1423 VDD.n155 VDD.n154 3.1505
R1424 VDD.n206 VDD.n155 3.1505
R1425 VDD.n164 VDD.n157 3.1505
R1426 VDD.n205 VDD.n157 3.1505
R1427 VDD.n203 VDD.n202 3.1505
R1428 VDD.n204 VDD.n203 3.1505
R1429 VDD.n201 VDD.n158 3.1505
R1430 VDD.n178 VDD.n158 3.1505
R1431 VDD.n200 VDD.n199 3.1505
R1432 VDD.n199 VDD.n198 3.1505
R1433 VDD.n338 VDD.n281 3.1505
R1434 VDD.n301 VDD.n281 3.1505
R1435 VDD.n337 VDD.n336 3.1505
R1436 VDD.n336 VDD.n335 3.1505
R1437 VDD.n283 VDD.n282 3.1505
R1438 VDD.n334 VDD.n283 3.1505
R1439 VDD.n329 VDD.n284 3.1505
R1440 VDD.n292 VDD.n284 3.1505
R1441 VDD.n328 VDD.n327 3.1505
R1442 VDD.n327 VDD.n326 3.1505
R1443 VDD.n291 VDD.n290 3.1505
R1444 VDD.n325 VDD.n291 3.1505
R1445 VDD.n332 VDD.n331 3.1505
R1446 VDD.n333 VDD.n332 3.1505
R1447 VDD.n309 VDD.n293 3.1505
R1448 VDD.n324 VDD.n293 3.1505
R1449 VDD.n322 VDD.n321 3.1505
R1450 VDD.n323 VDD.n322 3.1505
R1451 VDD.n320 VDD.n294 3.1505
R1452 VDD.n315 VDD.n294 3.1505
R1453 VDD.n1747 VDD.n577 3.1505
R1454 VDD.n1752 VDD.n1751 3.1505
R1455 VDD.n1750 VDD.n575 3.1505
R1456 VDD.n1754 VDD.n575 3.1505
R1457 VDD.n1756 VDD.n576 3.1505
R1458 VDD.n1756 VDD.n1755 3.1505
R1459 VDD.n1758 VDD.n574 3.1505
R1460 VDD.n1761 VDD.n1760 3.1505
R1461 VDD.n1760 VDD.n1759 3.1505
R1462 VDD.n1763 VDD.n571 3.1505
R1463 VDD.n571 VDD.n570 3.1505
R1464 VDD.n1765 VDD.n1764 3.1505
R1465 VDD.n1766 VDD.n1765 3.1505
R1466 VDD.n572 VDD.n526 3.1505
R1467 VDD.n1812 VDD.n1811 3.1505
R1468 VDD.n529 VDD.n525 3.1505
R1469 VDD.n1815 VDD.n523 3.1505
R1470 VDD.n530 VDD.n523 3.1505
R1471 VDD.n1817 VDD.n1816 3.1505
R1472 VDD.n1818 VDD.n1817 3.1505
R1473 VDD.n516 VDD.n515 3.1505
R1474 VDD.n1819 VDD.n516 3.1505
R1475 VDD.n1829 VDD.n1828 3.1505
R1476 VDD.n1828 VDD.n1827 3.1505
R1477 VDD.n1830 VDD.n514 3.1505
R1478 VDD.n518 VDD.n514 3.1505
R1479 VDD.n1832 VDD.n1831 3.1505
R1480 VDD.n1833 VDD.n1832 3.1505
R1481 VDD.n487 VDD.n485 3.1505
R1482 VDD.n1834 VDD.n487 3.1505
R1483 VDD.n1855 VDD.n1854 3.1505
R1484 VDD.n1854 VDD.n1853 3.1505
R1485 VDD.n488 VDD.n486 3.1505
R1486 VDD.n1840 VDD.n488 3.1505
R1487 VDD.n1843 VDD.n1842 3.1505
R1488 VDD.n1844 VDD.n1843 3.1505
R1489 VDD.n421 VDD.n418 3.1505
R1490 VDD.n1845 VDD.n421 3.1505
R1491 VDD.n1808 VDD.n524 3.1505
R1492 VDD.n539 VDD.n528 3.1505
R1493 VDD.n1804 VDD.n1803 3.1505
R1494 VDD.n1801 VDD.n537 3.1505
R1495 VDD.n1800 VDD.n1799 3.1505
R1496 VDD.n1798 VDD.n1797 3.1505
R1497 VDD.n1795 VDD.n1794 3.1505
R1498 VDD.n1793 VDD.n1792 3.1505
R1499 VDD.n1791 VDD.n1790 3.1505
R1500 VDD.n1789 VDD.n1788 3.1505
R1501 VDD.n1787 VDD.n1786 3.1505
R1502 VDD.n1785 VDD.n1784 3.1505
R1503 VDD.n1782 VDD.n1781 3.1505
R1504 VDD.n1780 VDD.n1779 3.1505
R1505 VDD.n1778 VDD.n1777 3.1505
R1506 VDD.n1723 VDD.n1722 3.1505
R1507 VDD.n1725 VDD.n1724 3.1505
R1508 VDD.n1727 VDD.n1726 3.1505
R1509 VDD.n1729 VDD.n1728 3.1505
R1510 VDD.n1731 VDD.n1730 3.1505
R1511 VDD.n1733 VDD.n1732 3.1505
R1512 VDD.n1735 VDD.n1734 3.1505
R1513 VDD.n1737 VDD.n1736 3.1505
R1514 VDD.n1739 VDD.n1738 3.1505
R1515 VDD.n1741 VDD.n1740 3.1505
R1516 VDD.n579 VDD.n578 3.1505
R1517 VDD.n1746 VDD.n1745 3.1505
R1518 VDD VDD.n1649 3.1505
R1519 VDD.n1657 VDD.n1649 3.1505
R1520 VDD.n1669 VDD.n1668 3.1505
R1521 VDD.n1668 VDD.n1667 3.1505
R1522 VDD.n1656 VDD.n1655 3.1505
R1523 VDD.n1666 VDD.n1656 3.1505
R1524 VDD.n1664 VDD.n1663 3.1505
R1525 VDD.n1665 VDD.n1664 3.1505
R1526 VDD.n1662 VDD.n1658 3.1505
R1527 VDD.n1677 VDD.n1676 3.1505
R1528 VDD.n1646 VDD.n1645 3.1505
R1529 VDD.n1675 VDD.n1646 3.1505
R1530 VDD.n1673 VDD.n1672 3.1505
R1531 VDD.n1674 VDD.n1673 3.1505
R1532 VDD.n1671 VDD.n1648 3.1505
R1533 VDD.n1648 VDD.n1647 3.1505
R1534 VDD.n1637 VDD.n1636 3.1505
R1535 VDD.n1684 VDD.n1637 3.1505
R1536 VDD.n1682 VDD.n1681 3.1505
R1537 VDD.n1683 VDD.n1682 3.1505
R1538 VDD.n1680 VDD.n1638 3.1505
R1539 VDD.n678 VDD.n667 3.1505
R1540 VDD.n670 VDD.n667 3.1505
R1541 VDD.n677 VDD.n676 3.1505
R1542 VDD.n676 VDD.n675 3.1505
R1543 VDD.n669 VDD.n668 3.1505
R1544 VDD.n674 VDD.n669 3.1505
R1545 VDD.n673 VDD.n672 3.1505
R1546 VDD.n686 VDD.n656 3.1505
R1547 VDD.n685 VDD.n658 3.1505
R1548 VDD.n685 VDD.n684 3.1505
R1549 VDD.n661 VDD.n657 3.1505
R1550 VDD.n683 VDD.n657 3.1505
R1551 VDD.n681 VDD.n680 3.1505
R1552 VDD.n682 VDD.n681 3.1505
R1553 VDD VDD.n660 3.1505
R1554 VDD.n660 VDD.n659 3.1505
R1555 VDD.n692 VDD.n691 3.1505
R1556 VDD.n698 VDD.n697 3.1505
R1557 VDD.n699 VDD.n698 3.1505
R1558 VDD.n696 VDD.n651 3.1505
R1559 VDD.n651 VDD.n650 3.1505
R1560 VDD.n695 VDD.n694 3.1505
R1561 VDD.n694 VDD.n693 3.1505
R1562 VDD.n640 VDD.n639 3.1505
R1563 VDD.n706 VDD.n705 3.1505
R1564 VDD.n707 VDD.n706 3.1505
R1565 VDD.n704 VDD.n642 3.1505
R1566 VDD.n642 VDD.n641 3.1505
R1567 VDD.n703 VDD.n702 3.1505
R1568 VDD.n702 VDD.n701 3.1505
R1569 VDD VDD.n649 3.1505
R1570 VDD.n700 VDD.n649 3.1505
R1571 VDD.n1556 VDD.n1555 3.1505
R1572 VDD.n1539 VDD.n721 3.1505
R1573 VDD.n721 VDD.n720 3.1505
R1574 VDD.n1546 VDD.n1545 3.1505
R1575 VDD.n1547 VDD.n1546 3.1505
R1576 VDD.n1544 VDD.n719 3.1505
R1577 VDD.n1543 VDD.n717 3.1505
R1578 VDD.n1550 VDD.n717 3.1505
R1579 VDD.n1552 VDD.n716 3.1505
R1580 VDD.n1552 VDD.n1551 3.1505
R1581 VDD.n1554 VDD.n1553 3.1505
R1582 VDD.n1538 VDD.n1537 3.1505
R1583 VDD.n1537 VDD.n1536 3.1505
R1584 VDD.n729 VDD.n728 3.1505
R1585 VDD.n724 VDD.n723 3.1505
R1586 VDD.n1283 VDD.n1282 3.1505
R1587 VDD.n1282 VDD.n1281 3.1505
R1588 VDD.n1284 VDD.n804 3.1505
R1589 VDD.n804 VDD.n801 3.1505
R1590 VDD.n1286 VDD.n1285 3.1505
R1591 VDD.n1287 VDD.n1286 3.1505
R1592 VDD.n797 VDD.n796 3.1505
R1593 VDD.n802 VDD.n797 3.1505
R1594 VDD.n1298 VDD.n1297 3.1505
R1595 VDD.n1297 VDD.n1296 3.1505
R1596 VDD.n1299 VDD.n790 3.1505
R1597 VDD.n790 VDD.n789 3.1505
R1598 VDD.n1303 VDD.n1302 3.1505
R1599 VDD.n1304 VDD.n1303 3.1505
R1600 VDD.n1301 VDD.n795 3.1505
R1601 VDD.n795 VDD.n794 3.1505
R1602 VDD.n782 VDD.n781 3.1505
R1603 VDD.n792 VDD.n781 3.1505
R1604 VDD.n1368 VDD.n1367 3.1505
R1605 VDD.n1369 VDD.n1368 3.1505
R1606 VDD.n772 VDD.n771 3.1505
R1607 VDD.n779 VDD.n772 3.1505
R1608 VDD.n1381 VDD.n1380 3.1505
R1609 VDD.n1380 VDD.n1379 3.1505
R1610 VDD.n1382 VDD.n770 3.1505
R1611 VDD.n770 VDD.n768 3.1505
R1612 VDD.n1384 VDD.n1383 3.1505
R1613 VDD.n1385 VDD.n1384 3.1505
R1614 VDD.n763 VDD.n762 3.1505
R1615 VDD.n764 VDD.n763 3.1505
R1616 VDD.n1397 VDD.n1396 3.1505
R1617 VDD.n1396 VDD.n1395 3.1505
R1618 VDD.n1398 VDD.n760 3.1505
R1619 VDD.n760 VDD.n758 3.1505
R1620 VDD.n1401 VDD.n1400 3.1505
R1621 VDD.n1402 VDD.n1401 3.1505
R1622 VDD.n753 VDD.n752 3.1505
R1623 VDD.n754 VDD.n753 3.1505
R1624 VDD.n1414 VDD.n1413 3.1505
R1625 VDD.n1413 VDD.n1412 3.1505
R1626 VDD.n1415 VDD.n750 3.1505
R1627 VDD.n750 VDD.n748 3.1505
R1628 VDD.n806 VDD.n805 3.1505
R1629 VDD.n809 VDD.n806 3.1505
R1630 VDD.n943 VDD.n911 3.1505
R1631 VDD.n886 VDD.n880 3.1505
R1632 VDD.n888 VDD.n886 3.1505
R1633 VDD.n962 VDD.n961 3.1505
R1634 VDD.n963 VDD.n962 3.1505
R1635 VDD.n959 VDD.n906 3.1505
R1636 VDD.n909 VDD.n906 3.1505
R1637 VDD.n954 VDD.n953 3.1505
R1638 VDD.n955 VDD.n954 3.1505
R1639 VDD.n965 VDD.n904 3.1505
R1640 VDD.n965 VDD.n964 3.1505
R1641 VDD.n960 VDD.n903 3.1505
R1642 VDD.n905 VDD.n903 3.1505
R1643 VDD.n958 VDD.n957 3.1505
R1644 VDD.n957 VDD.n956 3.1505
R1645 VDD VDD.n969 3.1505
R1646 VDD.n969 VDD.n968 3.1505
R1647 VDD.n966 VDD 3.1505
R1648 VDD.n967 VDD.n966 3.1505
R1649 VDD.n843 VDD.n838 3.1505
R1650 VDD.n865 VDD.n838 3.1505
R1651 VDD.n983 VDD.n982 3.1505
R1652 VDD.n982 VDD.n981 3.1505
R1653 VDD.n890 VDD.n839 3.1505
R1654 VDD.n894 VDD.n839 3.1505
R1655 VDD.n859 VDD.n858 3.1505
R1656 VDD.n858 VDD.n848 3.1505
R1657 VDD.n869 VDD.n841 3.1505
R1658 VDD.n870 VDD.n869 3.1505
R1659 VDD.n899 VDD.n889 3.1505
R1660 VDD.n895 VDD.n889 3.1505
R1661 VDD.n864 VDD.n842 3.1505
R1662 VDD.n856 VDD.n849 3.1505
R1663 VDD.n860 VDD.n842 3.1505
R1664 VDD.n868 VDD.n836 3.1505
R1665 VDD.n868 VDD.n840 3.1505
R1666 VDD.n1101 VDD.n1097 3.1505
R1667 VDD.n1096 VDD.n1095 3.1505
R1668 VDD.n1104 VDD.n1096 3.1505
R1669 VDD.n1107 VDD.n1106 3.1505
R1670 VDD.n1106 VDD.n1105 3.1505
R1671 VDD.n1108 VDD.n1089 3.1505
R1672 VDD.n1089 VDD.n1088 3.1505
R1673 VDD.n1110 VDD 3.1505
R1674 VDD.n1111 VDD.n1110 3.1505
R1675 VDD.n1087 VDD.n1086 3.1505
R1676 VDD.n1112 VDD.n1087 3.1505
R1677 VDD.n1116 VDD.n1115 3.1505
R1678 VDD.n1115 VDD.n1114 3.1505
R1679 VDD.n1117 VDD.n1085 3.1505
R1680 VDD.n1113 VDD.n1085 3.1505
R1681 VDD.n1084 VDD.n1083 3.1505
R1682 VDD.n1037 VDD.n1035 3.1505
R1683 VDD.n1037 VDD.n1036 3.1505
R1684 VDD.n1039 VDD.n1038 3.1505
R1685 VDD.n1038 VDD.n1026 3.1505
R1686 VDD.n1025 VDD.n1024 3.1505
R1687 VDD.n1042 VDD.n1025 3.1505
R1688 VDD.n1045 VDD.n1044 3.1505
R1689 VDD.n1044 VDD.n1043 3.1505
R1690 VDD.n1035 VDD.n1027 3.1505
R1691 VDD.n1036 VDD.n1027 3.1505
R1692 VDD.n1040 VDD.n1039 3.1505
R1693 VDD.n1040 VDD.n1026 3.1505
R1694 VDD.n1041 VDD.n1024 3.1505
R1695 VDD.n1042 VDD.n1041 3.1505
R1696 VDD.n1045 VDD.n1023 3.1505
R1697 VDD.n1043 VDD.n1023 3.1505
R1698 VDD VDD.n1020 3.1505
R1699 VDD.n1022 VDD.n1020 3.1505
R1700 VDD.n1060 VDD.n1021 3.1505
R1701 VDD.n1060 VDD.n1059 3.1505
R1702 VDD.n1061 VDD.n1018 3.1505
R1703 VDD.n1062 VDD.n1061 3.1505
R1704 VDD.n1065 VDD.n1017 3.1505
R1705 VDD.n1063 VDD.n1017 3.1505
R1706 VDD.n1067 VDD.n1066 3.1505
R1707 VDD.n1068 VDD.n1067 3.1505
R1708 VDD.n1071 VDD.n1015 3.1505
R1709 VDD.n1069 VDD.n1015 3.1505
R1710 VDD.n1057 VDD 3.1505
R1711 VDD.n1057 VDD.n1022 3.1505
R1712 VDD.n1058 VDD.n1021 3.1505
R1713 VDD.n1059 VDD.n1058 3.1505
R1714 VDD.n1019 VDD.n1018 3.1505
R1715 VDD.n1062 VDD.n1019 3.1505
R1716 VDD.n1065 VDD.n1064 3.1505
R1717 VDD.n1064 VDD.n1063 3.1505
R1718 VDD.n1066 VDD.n1016 3.1505
R1719 VDD.n1068 VDD.n1016 3.1505
R1720 VDD.n1207 VDD.n1206 3.1505
R1721 VDD.n1206 VDD.n1197 3.1505
R1722 VDD.n1205 VDD.n1196 3.1505
R1723 VDD.n1205 VDD.n1204 3.1505
R1724 VDD.n1199 VDD.n1198 3.1505
R1725 VDD.n1203 VDD.n1198 3.1505
R1726 VDD.n1202 VDD.n1201 3.1505
R1727 VDD.n1177 VDD.n1176 3.1505
R1728 VDD.n1210 VDD.n1209 3.1505
R1729 VDD.n1211 VDD.n1210 3.1505
R1730 VDD VDD.n1190 3.1505
R1731 VDD.n1190 VDD.n1189 3.1505
R1732 VDD.n1273 VDD.n808 3.1505
R1733 VDD.n1271 VDD.n1270 3.1505
R1734 VDD.n1269 VDD.n812 3.1505
R1735 VDD.n1267 VDD.n1266 3.1505
R1736 VDD.n1265 VDD.n814 3.1505
R1737 VDD.n1263 VDD.n1262 3.1505
R1738 VDD.n1261 VDD.n816 3.1505
R1739 VDD.n1259 VDD.n1258 3.1505
R1740 VDD.n1257 VDD.n818 3.1505
R1741 VDD.n1255 VDD.n1254 3.1505
R1742 VDD.n1252 VDD.n820 3.1505
R1743 VDD.n1251 VDD.n1250 3.1505
R1744 VDD.n1249 VDD.n822 3.1505
R1745 VDD.n1247 VDD.n1246 3.1505
R1746 VDD.n1244 VDD.n824 3.1505
R1747 VDD.n1243 VDD.n1242 3.1505
R1748 VDD.n1276 VDD.n807 3.1505
R1749 VDD.n810 VDD.n807 3.1505
R1750 VDD.n1278 VDD.n1277 3.1505
R1751 VDD.n1279 VDD.n1278 3.1505
R1752 VDD.n800 VDD.n799 3.1505
R1753 VDD.n1280 VDD.n800 3.1505
R1754 VDD.n1290 VDD.n1289 3.1505
R1755 VDD.n1289 VDD.n1288 3.1505
R1756 VDD.n1291 VDD.n798 3.1505
R1757 VDD.n803 VDD.n798 3.1505
R1758 VDD.n1293 VDD.n1292 3.1505
R1759 VDD.n1294 VDD.n1293 3.1505
R1760 VDD.n787 VDD.n785 3.1505
R1761 VDD.n1295 VDD.n787 3.1505
R1762 VDD.n1307 VDD.n1306 3.1505
R1763 VDD.n1306 VDD.n1305 3.1505
R1764 VDD.n788 VDD.n786 3.1505
R1765 VDD.n791 VDD.n788 3.1505
R1766 VDD.n778 VDD.n777 3.1505
R1767 VDD.n793 VDD.n778 3.1505
R1768 VDD.n1372 VDD.n1371 3.1505
R1769 VDD.n1371 VDD.n1370 3.1505
R1770 VDD.n1374 VDD.n773 3.1505
R1771 VDD.n780 VDD.n773 3.1505
R1772 VDD.n1376 VDD.n1375 3.1505
R1773 VDD.n1377 VDD.n1376 3.1505
R1774 VDD.n767 VDD.n766 3.1505
R1775 VDD.n1378 VDD.n767 3.1505
R1776 VDD.n1388 VDD.n1387 3.1505
R1777 VDD.n1387 VDD.n1386 3.1505
R1778 VDD.n1389 VDD.n765 3.1505
R1779 VDD.n769 VDD.n765 3.1505
R1780 VDD.n1392 VDD.n1391 3.1505
R1781 VDD.n1393 VDD.n1392 3.1505
R1782 VDD.n1390 VDD.n757 3.1505
R1783 VDD.n1394 VDD.n757 3.1505
R1784 VDD.n1405 VDD.n1404 3.1505
R1785 VDD.n1404 VDD.n1403 3.1505
R1786 VDD.n1406 VDD.n755 3.1505
R1787 VDD.n759 VDD.n755 3.1505
R1788 VDD.n1409 VDD.n1408 3.1505
R1789 VDD.n1410 VDD.n1409 3.1505
R1790 VDD.n1407 VDD.n747 3.1505
R1791 VDD.n1411 VDD.n747 3.1505
R1792 VDD.n1422 VDD.n1421 3.1505
R1793 VDD.n1421 VDD.n1420 3.1505
R1794 VDD.n1423 VDD.n745 3.1505
R1795 VDD.n749 VDD.n745 3.1505
R1796 VDD.n1425 VDD.n1424 3.1505
R1797 VDD.n1426 VDD.n1425 3.1505
R1798 VDD.n738 VDD.n737 3.1505
R1799 VDD.n1427 VDD.n738 3.1505
R1800 VDD.n1438 VDD.n1437 3.1505
R1801 VDD.n1437 VDD.n1436 3.1505
R1802 VDD.n1439 VDD.n735 3.1505
R1803 VDD.n740 VDD.n735 3.1505
R1804 VDD.n1525 VDD.n1524 3.1505
R1805 VDD.n1526 VDD.n1525 3.1505
R1806 VDD.n1418 VDD.n1417 3.1505
R1807 VDD.n1419 VDD.n1418 3.1505
R1808 VDD.n743 VDD.n742 3.1505
R1809 VDD.n744 VDD.n743 3.1505
R1810 VDD.n1430 VDD.n1429 3.1505
R1811 VDD.n1429 VDD.n1428 3.1505
R1812 VDD.n1431 VDD.n741 3.1505
R1813 VDD.n741 VDD.n739 3.1505
R1814 VDD.n1434 VDD.n1433 3.1505
R1815 VDD.n1435 VDD.n1434 3.1505
R1816 VDD.n1432 VDD.n733 3.1505
R1817 VDD.n734 VDD.n733 3.1505
R1818 VDD.n1528 VDD.n730 3.1505
R1819 VDD.n1528 VDD.n1527 3.1505
R1820 VDD.n1534 VDD.n1533 3.1505
R1821 VDD.n1535 VDD.n1534 3.1505
R1822 VDD.n1491 VDD.n1440 3.1505
R1823 VDD.n1490 VDD.n1489 3.1505
R1824 VDD.n1487 VDD.n1486 3.1505
R1825 VDD.n1485 VDD.n1484 3.1505
R1826 VDD.n1483 VDD.n1482 3.1505
R1827 VDD.n1481 VDD.n1480 3.1505
R1828 VDD.n1479 VDD.n1478 3.1505
R1829 VDD.n1477 VDD.n1476 3.1505
R1830 VDD.n1474 VDD.n1473 3.1505
R1831 VDD.n1472 VDD.n1457 3.1505
R1832 VDD.n1470 VDD.n1469 3.1505
R1833 VDD.n1467 VDD.n1459 3.1505
R1834 VDD.n732 VDD.n731 3.1505
R1835 VDD.n1531 VDD.n1530 3.1505
R1836 VDD.n1530 VDD.n726 3.1505
R1837 VDD.n1494 VDD.n1493 3.1505
R1838 VDD.n1522 VDD.n1521 3.1505
R1839 VDD.n1519 VDD.n1518 3.1505
R1840 VDD.n1516 VDD.n1497 3.1505
R1841 VDD.n1497 VDD.n1496 3.1505
R1842 VDD.n1515 VDD.n1514 3.1505
R1843 VDD.n1514 VDD.n1513 3.1505
R1844 VDD.n1502 VDD.n1501 3.1505
R1845 VDD.n1512 VDD.n1502 3.1505
R1846 VDD.n1510 VDD.n1509 3.1505
R1847 VDD.n1511 VDD.n1510 3.1505
R1848 VDD.n1508 VDD.n1505 3.1505
R1849 VDD.n625 VDD.n623 3.1505
R1850 VDD.n1558 VDD.n1557 3.1505
R1851 VDD.n1560 VDD.n1559 3.1505
R1852 VDD.n1562 VDD.n1561 3.1505
R1853 VDD.n1564 VDD.n1563 3.1505
R1854 VDD.n1566 VDD.n1565 3.1505
R1855 VDD.n1568 VDD.n1567 3.1505
R1856 VDD.n1570 VDD.n1569 3.1505
R1857 VDD.n1572 VDD.n1571 3.1505
R1858 VDD.n1574 VDD.n1573 3.1505
R1859 VDD.n1576 VDD.n1575 3.1505
R1860 VDD.n1578 VDD.n1577 3.1505
R1861 VDD.n1580 VDD.n1579 3.1505
R1862 VDD.n1582 VDD.n1581 3.1505
R1863 VDD.n626 VDD.n624 3.1505
R1864 VDD.n1587 VDD.n1586 3.1505
R1865 VDD VDD.n1604 3.1505
R1866 VDD.n1604 VDD.n1603 3.1505
R1867 VDD.n1596 VDD.n1595 3.1505
R1868 VDD.n1597 VDD.n622 3.1505
R1869 VDD.n622 VDD.n621 3.1505
R1870 VDD.n1600 VDD.n1599 3.1505
R1871 VDD.n1601 VDD.n1600 3.1505
R1872 VDD.n1598 VDD.n620 3.1505
R1873 VDD.n1602 VDD.n620 3.1505
R1874 VDD.n1605 VDD.n613 3.1505
R1875 VDD.n613 VDD.n612 3.1505
R1876 VDD.n1607 VDD.n1606 3.1505
R1877 VDD.n1608 VDD.n1607 3.1505
R1878 VDD.n611 VDD.n610 3.1505
R1879 VDD.n1609 VDD.n611 3.1505
R1880 VDD.n1611 VDD.n1610 3.1505
R1881 VDD.n1625 VDD.n1624 3.1505
R1882 VDD.n1629 VDD.n596 3.1505
R1883 VDD.n1630 VDD.n1629 3.1505
R1884 VDD.n1628 VDD.n1627 3.1505
R1885 VDD.n1628 VDD.n1620 3.1505
R1886 VDD.n1626 VDD.n1621 3.1505
R1887 VDD.n1623 VDD.n1621 3.1505
R1888 VDD.n604 VDD 3.1505
R1889 VDD.n1631 VDD.n604 3.1505
R1890 VDD.n1616 VDD.n605 3.1505
R1891 VDD.n1617 VDD.n602 3.1505
R1892 VDD.n1618 VDD.n1617 3.1505
R1893 VDD.n1619 VDD.n603 3.1505
R1894 VDD.n1633 VDD.n1632 3.1505
R1895 VDD.n1687 VDD.n1686 3.1505
R1896 VDD.n1686 VDD.n1685 3.1505
R1897 VDD VDD.n595 3.1505
R1898 VDD.n595 VDD.n594 3.1505
R1899 VDD.n1690 VDD.n1689 3.1505
R1900 VDD.n1691 VDD.n1690 3.1505
R1901 VDD.n593 VDD.n592 3.1505
R1902 VDD.n1692 VDD.n593 3.1505
R1903 VDD.n1694 VDD.n1693 3.1505
R1904 VDD.n1721 VDD.n581 3.1505
R1905 VDD.n1743 VDD.n581 3.1505
R1906 VDD.n1720 VDD.n1719 3.1505
R1907 VDD.n1718 VDD.n1717 3.1505
R1908 VDD.n1707 VDD.n1704 3.1505
R1909 VDD.n1713 VDD.n1712 3.1505
R1910 VDD.n1714 VDD.n1713 3.1505
R1911 VDD.n1710 VDD.n1706 3.1505
R1912 VDD.n1706 VDD.n1705 3.1505
R1913 VDD.n1709 VDD.n566 3.1505
R1914 VDD.n568 VDD.n566 3.1505
R1915 VDD.n1770 VDD.n567 3.1505
R1916 VDD.n1770 VDD.n1769 3.1505
R1917 VDD.n1772 VDD.n1771 3.1505
R1918 VDD.n1775 VDD.n1774 3.1505
R1919 VDD.n1716 VDD.n1703 3.1505
R1920 VDD.n521 VDD.n520 3.1505
R1921 VDD.n522 VDD.n521 3.1505
R1922 VDD.n1822 VDD.n1821 3.1505
R1923 VDD.n1821 VDD.n1820 3.1505
R1924 VDD.n1823 VDD.n519 3.1505
R1925 VDD.n519 VDD.n517 3.1505
R1926 VDD.n1825 VDD.n1824 3.1505
R1927 VDD.n1826 VDD.n1825 3.1505
R1928 VDD.n512 VDD.n511 3.1505
R1929 VDD.n513 VDD.n512 3.1505
R1930 VDD.n1836 VDD.n1835 3.1505
R1931 VDD.n1835 VDD.t336 3.1505
R1932 VDD.n1837 VDD.n490 3.1505
R1933 VDD.n490 VDD.n489 3.1505
R1934 VDD.n1851 VDD.n1850 3.1505
R1935 VDD.n1852 VDD.n1851 3.1505
R1936 VDD.n1849 VDD.n491 3.1505
R1937 VDD.n1841 VDD.n491 3.1505
R1938 VDD.n1848 VDD.n1847 3.1505
R1939 VDD.n1847 VDD.n1846 3.1505
R1940 VDD.n1839 VDD.n424 3.1505
R1941 VDD.n424 VDD.n423 3.1505
R1942 VDD.n2007 VDD.n2006 3.1505
R1943 VDD.n2008 VDD.n2007 3.1505
R1944 VDD.n2005 VDD.n425 3.1505
R1945 VDD.n430 VDD.n425 3.1505
R1946 VDD.n2004 VDD.n2003 3.1505
R1947 VDD.n2003 VDD.n2002 3.1505
R1948 VDD.n428 VDD.n427 3.1505
R1949 VDD.n432 VDD.n428 3.1505
R1950 VDD.n442 VDD.n440 3.1505
R1951 VDD.n440 VDD.n439 3.1505
R1952 VDD.n1993 VDD.n1992 3.1505
R1953 VDD.n1994 VDD.n1993 3.1505
R1954 VDD.n1991 VDD.n441 3.1505
R1955 VDD.n449 VDD.n441 3.1505
R1956 VDD.n1989 VDD.n1988 3.1505
R1957 VDD.n1988 VDD.n1987 3.1505
R1958 VDD.n447 VDD.n446 3.1505
R1959 VDD.n451 VDD.n447 3.1505
R1960 VDD.n462 VDD.n460 3.1505
R1961 VDD.n460 VDD.n459 3.1505
R1962 VDD.n1978 VDD.n1977 3.1505
R1963 VDD.n1979 VDD.n1978 3.1505
R1964 VDD.n1975 VDD.n461 3.1505
R1965 VDD.n1879 VDD.n461 3.1505
R1966 VDD.n1974 VDD.n1973 3.1505
R1967 VDD.n1973 VDD.n1972 3.1505
R1968 VDD.n1878 VDD.n1877 3.1505
R1969 VDD.n1881 VDD.n1878 3.1505
R1970 VDD.n1893 VDD.n1891 3.1505
R1971 VDD.n1891 VDD.n1889 3.1505
R1972 VDD.n1963 VDD.n1962 3.1505
R1973 VDD.n1964 VDD.n1963 3.1505
R1974 VDD.n1961 VDD.n1892 3.1505
R1975 VDD.n1946 VDD.n1892 3.1505
R1976 VDD.n1960 VDD.n1959 3.1505
R1977 VDD.n1917 VDD.n1911 3.1505
R1978 VDD.n1921 VDD.n1911 3.1505
R1979 VDD.n1923 VDD.n1912 3.1505
R1980 VDD.n1923 VDD.n1922 3.1505
R1981 VDD.n1924 VDD.n1910 3.1505
R1982 VDD.n1924 VDD.n1905 3.1505
R1983 VDD.n1926 VDD.n1925 3.1505
R1984 VDD.n1925 VDD.n1906 3.1505
R1985 VDD.n1927 VDD.n1908 3.1505
R1986 VDD.n1908 VDD.n1907 3.1505
R1987 VDD.n1930 VDD.n1929 3.1505
R1988 VDD.n1931 VDD.n1930 3.1505
R1989 VDD.n1901 VDD.n1899 3.1505
R1990 VDD.n1899 VDD.n1897 3.1505
R1991 VDD.n1953 VDD.n1952 3.1505
R1992 VDD.n1954 VDD.n1953 3.1505
R1993 VDD.n1950 VDD.n1900 3.1505
R1994 VDD.n1900 VDD.n1898 3.1505
R1995 VDD.n1949 VDD.n1948 3.1505
R1996 VDD.n1948 VDD.n1947 3.1505
R1997 VDD.n1904 VDD.n1903 3.1505
R1998 VDD.n1945 VDD.n1904 3.1505
R1999 VDD.n1943 VDD.n1942 3.1505
R2000 VDD.n1944 VDD.n1943 3.1505
R2001 VDD.n1940 VDD.n1933 3.1505
R2002 VDD.n1933 VDD.n1932 3.1505
R2003 VDD.n1939 VDD.n1938 3.1505
R2004 VDD.n1938 VDD.n1937 3.1505
R2005 VDD.n1936 VDD.n1935 3.1505
R2006 VDD.n1936 VDD.n1896 3.1505
R2007 VDD.n1919 VDD.n1918 3.1505
R2008 VDD.n1914 VDD.n1913 3.1505
R2009 VDD.n1887 VDD.n1886 3.1505
R2010 VDD.n1890 VDD.n1887 3.1505
R2011 VDD.n422 VDD.n419 3.1505
R2012 VDD.n429 VDD.n422 3.1505
R2013 VDD.n435 VDD.n433 3.1505
R2014 VDD.n433 VDD.n431 3.1505
R2015 VDD.n2000 VDD.n1999 3.1505
R2016 VDD.n2001 VDD.n2000 3.1505
R2017 VDD.n1998 VDD.n434 3.1505
R2018 VDD.n438 VDD.n434 3.1505
R2019 VDD.n1997 VDD.n1996 3.1505
R2020 VDD.n1996 VDD.n1995 3.1505
R2021 VDD.n437 VDD.n436 3.1505
R2022 VDD.n448 VDD.n437 3.1505
R2023 VDD.n454 VDD.n452 3.1505
R2024 VDD.n452 VDD.n450 3.1505
R2025 VDD.n1985 VDD.n1984 3.1505
R2026 VDD.n1986 VDD.n1985 3.1505
R2027 VDD.n1983 VDD.n453 3.1505
R2028 VDD.n458 VDD.n453 3.1505
R2029 VDD.n1982 VDD.n1981 3.1505
R2030 VDD.n1981 VDD.n1980 3.1505
R2031 VDD.n1884 VDD.n456 3.1505
R2032 VDD.n457 VDD.n456 3.1505
R2033 VDD.n1885 VDD.n1882 3.1505
R2034 VDD.n1882 VDD.n1880 3.1505
R2035 VDD.n1970 VDD.n1969 3.1505
R2036 VDD.n1971 VDD.n1970 3.1505
R2037 VDD.n1968 VDD.n1883 3.1505
R2038 VDD.n1888 VDD.n1883 3.1505
R2039 VDD.n1967 VDD.n1966 3.1505
R2040 VDD.n1966 VDD.n1965 3.1505
R2041 VDD.n2011 VDD.n2010 3.1505
R2042 VDD.n2010 VDD.n2009 3.1505
R2043 VDD.n399 VDD.n398 3.1505
R2044 VDD.n400 VDD.n399 3.1505
R2045 VDD.n397 VDD.n365 3.1505
R2046 VDD.n379 VDD.n365 3.1505
R2047 VDD.n396 VDD.n395 3.1505
R2048 VDD.n395 VDD.n394 3.1505
R2049 VDD.n389 VDD.n380 3.1505
R2050 VDD.n384 VDD.n380 3.1505
R2051 VDD.n409 VDD.n408 3.1505
R2052 VDD.n410 VDD.n409 3.1505
R2053 VDD.n388 VDD.n387 3.1505
R2054 VDD.n387 VDD.n386 3.1505
R2055 VDD.n383 VDD.n358 3.1505
R2056 VDD.n385 VDD.n383 3.1505
R2057 VDD.n392 VDD.n391 3.1505
R2058 VDD.n393 VDD.n392 3.1505
R2059 VDD.n357 VDD.n356 3.1505
R2060 VDD.n411 VDD.n357 3.1505
R2061 VDD.n414 VDD.n413 3.1505
R2062 VDD.n413 VDD.n412 3.1505
R2063 VDD.n106 VDD.n66 3.1505
R2064 VDD.n2041 VDD.n66 3.1505
R2065 VDD.n2039 VDD.n2038 3.1505
R2066 VDD.n2040 VDD.n2039 3.1505
R2067 VDD.n2037 VDD.n67 3.1505
R2068 VDD.n112 VDD.n67 3.1505
R2069 VDD.n65 VDD.n60 3.1505
R2070 VDD.n2042 VDD.n65 3.1505
R2071 VDD.n83 VDD.n82 3.1505
R2072 VDD.n90 VDD.n83 3.1505
R2073 VDD.n92 VDD.n81 3.1505
R2074 VDD.n92 VDD.n91 3.1505
R2075 VDD.n94 VDD.n93 3.1505
R2076 VDD.n93 VDD.n74 3.1505
R2077 VDD.n88 VDD.n87 3.1505
R2078 VDD.n89 VDD.n88 3.1505
R2079 VDD.n84 VDD.n64 3.1505
R2080 VDD.n2044 VDD.n2043 3.1505
R2081 VDD.n2115 VDD.n2114 3.1505
R2082 VDD.n2114 VDD.n2113 3.1505
R2083 VDD.n2094 VDD.n2093 3.1505
R2084 VDD.n2093 VDD.n2092 3.1505
R2085 VDD.n2097 VDD.n2096 3.1505
R2086 VDD.n2096 VDD.n2095 3.1505
R2087 VDD VDD.n2105 3.1505
R2088 VDD.n2105 VDD.n2104 3.1505
R2089 VDD.n2103 VDD.n2101 3.1505
R2090 VDD.n2103 VDD.n2102 3.1505
R2091 VDD.n2100 VDD.n2099 3.1505
R2092 VDD.n2099 VDD.n2098 3.1505
R2093 VDD.n2088 VDD.n2087 3.1505
R2094 VDD.n2087 VDD.n2086 3.1505
R2095 VDD.n2075 VDD.n2074 3.1505
R2096 VDD.n2112 VDD.n2111 3.1505
R2097 VDD.n2148 VDD.n2147 3.1505
R2098 VDD.n2147 VDD.t54 3.1505
R2099 VDD.n2051 VDD.n2050 3.1505
R2100 VDD.n2146 VDD.n2145 3.1505
R2101 VDD.t54 VDD.n2146 3.1505
R2102 VDD.n1 VDD.n0 3.1505
R2103 VDD.n1176 VDD.n1175 3.14819
R2104 VDD.n220 VDD.n132 3.13854
R2105 VDD.n222 VDD.n129 3.13854
R2106 VDD.n223 VDD.n127 3.13854
R2107 VDD.n244 VDD.n237 3.13659
R2108 VDD.n250 VDD.n249 3.13659
R2109 VDD.n258 VDD.n247 3.13659
R2110 VDD.n1585 VDD.n626 3.09085
R2111 VDD.n1700 VDD.n1697 3.06224
R2112 VDD.n1654 VDD.n1653 3.06224
R2113 VDD.n666 VDD.n663 3.06224
R2114 VDD.n647 VDD.n644 3.06224
R2115 VDD.n885 VDD.n884 3.06224
R2116 VDD.n879 VDD.n876 3.06224
R2117 VDD.n1094 VDD.n1091 3.06224
R2118 VDD.n1050 VDD.n1047 3.06224
R2119 VDD.n1055 VDD.n1054 3.06224
R2120 VDD.n1195 VDD.n1192 3.06224
R2121 VDD.n618 VDD.n617 3.06224
R2122 VDD.n601 VDD.n600 3.06224
R2123 VDD.n2084 VDD.n2083 3.06224
R2124 VDD.n1744 VDD.n579 3.04049
R2125 VDD.n1724 VDD.n582 3.03982
R2126 VDD.n1559 VDD.n627 3.03982
R2127 VDD.n102 VDD.n69 2.98985
R2128 VDD.n73 VDD.n71 2.98985
R2129 VDD.n175 VDD.n167 2.98985
R2130 VDD.n171 VDD.n169 2.98985
R2131 VDD.n300 VDD.n298 2.98985
R2132 VDD.n305 VDD.n296 2.98985
R2133 VDD.n364 VDD.n362 2.98985
R2134 VDD.n404 VDD.n360 2.98985
R2135 VDD.n87 VDD.n86 2.98721
R2136 VDD.n63 VDD.n62 2.97811
R2137 VDD.n165 VDD.n160 2.97811
R2138 VDD.n163 VDD.n162 2.97811
R2139 VDD.n287 VDD.n286 2.97811
R2140 VDD.n330 VDD.n289 2.97811
R2141 VDD.n378 VDD.n377 2.97811
R2142 VDD.n390 VDD.n382 2.97811
R2143 VDD.n1294 VDD.t580 2.91474
R2144 VDD.n1395 VDD.t575 2.91474
R2145 VDD.n254 VDD.n252 2.88811
R2146 VDD.n934 VDD.n932 2.87637
R2147 VDD.n923 VDD.n921 2.87637
R2148 VDD.n1139 VDD.n1138 2.87637
R2149 VDD.n1134 VDD.n1133 2.87637
R2150 VDD.n2066 VDD.n2064 2.87637
R2151 VDD.n2119 VDD.n2118 2.87637
R2152 VDD.n78 VDD.t478 2.84673
R2153 VDD.n150 VDD.t16 2.84673
R2154 VDD.n278 VDD.t787 2.84631
R2155 VDD.n369 VDD.t309 2.84631
R2156 VDD.n37 VDD.n36 2.82741
R2157 VDD.n142 VDD.n136 2.78441
R2158 VDD.n141 VDD.n138 2.78441
R2159 VDD.n267 VDD.n261 2.78441
R2160 VDD.n266 VDD.n263 2.78441
R2161 VDD.n1807 VDD.n528 2.7478
R2162 VDD.n1805 VDD.n528 2.7478
R2163 VDD.n228 VDD.n118 2.74538
R2164 VDD.n2145 VDD.n2144 2.60854
R2165 VDD.n187 VDD.n184 2.6005
R2166 VDD.n143 VDD.n134 2.6005
R2167 VDD.n270 VDD.n269 2.6005
R2168 VDD.n314 VDD.n313 2.6005
R2169 VDD.n355 VDD.n354 2.6005
R2170 VDD.n478 VDD.n477 2.6005
R2171 VDD.n545 VDD.n544 2.6005
R2172 VDD.n551 VDD.n550 2.6005
R2173 VDD.n1700 VDD.n1699 2.6005
R2174 VDD.n1654 VDD.n1651 2.6005
R2175 VDD.n1464 VDD.n1461 2.6005
R2176 VDD.n1453 VDD.n1450 2.6005
R2177 VDD.n666 VDD.n665 2.6005
R2178 VDD.n647 VDD.n646 2.6005
R2179 VDD.n1331 VDD.n1330 2.6005
R2180 VDD.n1311 VDD.n1310 2.6005
R2181 VDD.n1317 VDD.n1313 2.6005
R2182 VDD.n1316 VDD.n1315 2.6005
R2183 VDD.n1320 VDD.n1319 2.6005
R2184 VDD.n776 VDD.n775 2.6005
R2185 VDD.n1356 VDD.n1355 2.6005
R2186 VDD.n1353 VDD.n1352 2.6005
R2187 VDD.n1359 VDD.n1358 2.6005
R2188 VDD.n1364 VDD.n1363 2.6005
R2189 VDD.n885 VDD.n882 2.6005
R2190 VDD.n879 VDD.n878 2.6005
R2191 VDD.n1094 VDD.n1093 2.6005
R2192 VDD.n1050 VDD.n1049 2.6005
R2193 VDD.n1055 VDD.n1052 2.6005
R2194 VDD.n1195 VDD.n1194 2.6005
R2195 VDD.n1323 VDD.n1322 2.6005
R2196 VDD.n1338 VDD.n1337 2.6005
R2197 VDD.n1335 VDD.n1334 2.6005
R2198 VDD.n1344 VDD.n1328 2.6005
R2199 VDD.n1345 VDD.n1326 2.6005
R2200 VDD.n1341 VDD.n1340 2.6005
R2201 VDD.n618 VDD.n615 2.6005
R2202 VDD.n601 VDD.n598 2.6005
R2203 VDD.n494 VDD.n493 2.6005
R2204 VDD.n484 VDD.n483 2.6005
R2205 VDD.n510 VDD.n509 2.6005
R2206 VDD.n500 VDD.n499 2.6005
R2207 VDD.n445 VDD.n444 2.6005
R2208 VDD.n1876 VDD.n1875 2.6005
R2209 VDD.n472 VDD.n471 2.6005
R2210 VDD.n466 VDD.n465 2.6005
R2211 VDD.n1869 VDD.n1868 2.6005
R2212 VDD.n1872 VDD.n1871 2.6005
R2213 VDD.n503 VDD.n502 2.6005
R2214 VDD.n475 VDD.n474 2.6005
R2215 VDD.n481 VDD.n480 2.6005
R2216 VDD.n497 VDD.n496 2.6005
R2217 VDD.n1860 VDD.n1859 2.6005
R2218 VDD.n111 VDD.n108 2.6005
R2219 VDD.n2084 VDD.n2081 2.6005
R2220 VDD.n1738 VDD.n590 2.59264
R2221 VDD.n1734 VDD.n588 2.59264
R2222 VDD.n1730 VDD.n586 2.59264
R2223 VDD.n1726 VDD.n584 2.59264
R2224 VDD.n1741 VDD.n590 2.59264
R2225 VDD.n1736 VDD.n588 2.59264
R2226 VDD.n1732 VDD.n586 2.59264
R2227 VDD.n1728 VDD.n584 2.59264
R2228 VDD.n1583 VDD.n1582 2.59264
R2229 VDD.n1577 VDD.n637 2.59264
R2230 VDD.n1573 VDD.n635 2.59264
R2231 VDD.n1569 VDD.n633 2.59264
R2232 VDD.n1565 VDD.n631 2.59264
R2233 VDD.n1561 VDD.n629 2.59264
R2234 VDD.n1583 VDD.n626 2.59264
R2235 VDD.n1579 VDD.n637 2.59264
R2236 VDD.n1575 VDD.n635 2.59264
R2237 VDD.n1571 VDD.n633 2.59264
R2238 VDD.n1567 VDD.n631 2.59264
R2239 VDD.n1563 VDD.n629 2.59264
R2240 VDD.n230 VDD.n228 2.588
R2241 VDD.n1955 VDD.n1954 2.58448
R2242 VDD.n1736 VDD.n589 2.5167
R2243 VDD.n1732 VDD.n587 2.5167
R2244 VDD.n1728 VDD.n585 2.5167
R2245 VDD.n1724 VDD.n583 2.5167
R2246 VDD.n1738 VDD.n589 2.5167
R2247 VDD.n1734 VDD.n587 2.5167
R2248 VDD.n1730 VDD.n585 2.5167
R2249 VDD.n1726 VDD.n583 2.5167
R2250 VDD.n1579 VDD.n638 2.5167
R2251 VDD.n1575 VDD.n636 2.5167
R2252 VDD.n1571 VDD.n634 2.5167
R2253 VDD.n1567 VDD.n632 2.5167
R2254 VDD.n1563 VDD.n630 2.5167
R2255 VDD.n1582 VDD.n638 2.5167
R2256 VDD.n1577 VDD.n636 2.5167
R2257 VDD.n1573 VDD.n634 2.5167
R2258 VDD.n1569 VDD.n632 2.5167
R2259 VDD.n1565 VDD.n630 2.5167
R2260 VDD.n1972 VDD.t347 2.49842
R2261 VDD.n1956 VDD.n1955 2.49842
R2262 VDD.n810 VDD.n809 2.49842
R2263 VDD.n1742 VDD.n1741 2.47755
R2264 VDD.n1742 VDD.n579 2.47755
R2265 VDD.n1559 VDD.n628 2.47755
R2266 VDD.n1561 VDD.n628 2.47755
R2267 VDD.n1239 VDD.n1238 2.37611
R2268 VDD.n2049 VDD.n2048 2.36122
R2269 VDD.n2138 VDD.n2077 2.35567
R2270 VDD.n1236 VDD.n1235 2.34319
R2271 VDD.n1235 VDD.n827 2.33916
R2272 VDD.n2143 VDD.n2142 2.32106
R2273 VDD.n1077 VDD.n1076 2.31932
R2274 VDD.n939 VDD.n938 2.29638
R2275 VDD.n939 VDD.n918 2.29115
R2276 VDD.n1235 VDD.n1234 2.28732
R2277 VDD.n945 VDD.n944 2.2804
R2278 VDD.n2015 VDD.n2014 2.27396
R2279 VDD.n1679 VDD.n1678 2.25904
R2280 VDD.n2056 VDD.n2055 2.25144
R2281 VDD.n2013 VDD.n417 2.25144
R2282 VDD.n951 VDD.n950 2.2505
R2283 VDD.n837 VDD.n835 2.2505
R2284 VDD.n846 VDD.n845 2.2505
R2285 VDD.n874 VDD.n873 2.2505
R2286 VDD.n1156 VDD.n993 2.2505
R2287 VDD.n1125 VDD.n1124 2.2505
R2288 VDD.n1006 VDD.n996 2.2505
R2289 VDD.n1146 VDD.n990 2.2505
R2290 VDD.n1151 VDD.n1150 2.2505
R2291 VDD.n48 VDD.n47 2.2505
R2292 VDD.n2137 VDD.n2136 2.2505
R2293 VDD.n1230 VDD.n828 2.24806
R2294 VDD.n932 VDD.t650 2.16717
R2295 VDD.n932 VDD.n931 2.16717
R2296 VDD.n921 VDD.t453 2.16717
R2297 VDD.n921 VDD.n920 2.16717
R2298 VDD.n1138 VDD.t646 2.16717
R2299 VDD.n1138 VDD.n1137 2.16717
R2300 VDD.n1133 VDD.t467 2.16717
R2301 VDD.n1133 VDD.n1132 2.16717
R2302 VDD.n2064 VDD.t90 2.16717
R2303 VDD.n2064 VDD.n2063 2.16717
R2304 VDD.n2118 VDD.t292 2.16717
R2305 VDD.n2118 VDD.n2117 2.16717
R2306 VDD.n2019 VDD.n2018 2.06447
R2307 VDD VDD.n371 2.06161
R2308 VDD.n980 VDD.n841 2.05248
R2309 VDD.t459 VDD.n894 2.05248
R2310 VDD.n964 VDD.t449 2.05248
R2311 VDD.n1043 VDD.t41 2.05248
R2312 VDD.n1490 VDD.n1441 2.04683
R2313 VDD.n1486 VDD.n1441 2.04625
R2314 VDD.n1781 VDD.n532 2.04615
R2315 VDD.n1785 VDD.n532 2.04615
R2316 VDD VDD.n75 2.01923
R2317 VDD.n1959 VDD.n1958 2.00622
R2318 VDD.n1958 VDD.n1895 2.00565
R2319 VDD.n1485 VDD.n1445 1.94801
R2320 VDD.n1482 VDD.n1445 1.94746
R2321 VDD.n1786 VDD.n533 1.94734
R2322 VDD.n1789 VDD.n533 1.94734
R2323 VDD.n940 VDD.n939 1.94241
R2324 VDD.n1214 VDD.n1180 1.9255
R2325 VDD.n1743 VDD.n1742 1.91272
R2326 VDD.n1584 VDD.n628 1.91272
R2327 VDD.n2045 VDD.n64 1.90984
R2328 VDD.n2045 VDD.n2044 1.90929
R2329 VDD.n1695 VDD.n1694 1.8985
R2330 VDD.n1743 VDD.n583 1.89315
R2331 VDD.n1743 VDD.n585 1.89315
R2332 VDD.n1743 VDD.n587 1.89315
R2333 VDD.n1743 VDD.n589 1.89315
R2334 VDD.n1584 VDD.n630 1.89315
R2335 VDD.n1584 VDD.n632 1.89315
R2336 VDD.n1584 VDD.n634 1.89315
R2337 VDD.n1584 VDD.n636 1.89315
R2338 VDD.n1584 VDD.n638 1.89315
R2339 VDD.n342 VDD.n274 1.87485
R2340 VDD.n572 VDD.n527 1.87282
R2341 VDD.n728 VDD.n725 1.87282
R2342 VDD.n1811 VDD.n527 1.87228
R2343 VDD.n725 VDD.n724 1.87228
R2344 VDD.n1717 VDD.n580 1.8617
R2345 VDD.n1719 VDD.n580 1.8617
R2346 VDD.n1743 VDD.n584 1.85518
R2347 VDD.n1743 VDD.n586 1.85518
R2348 VDD.n1743 VDD.n588 1.85518
R2349 VDD.n1743 VDD.n590 1.85518
R2350 VDD.n1584 VDD.n629 1.85518
R2351 VDD.n1584 VDD.n631 1.85518
R2352 VDD.n1584 VDD.n633 1.85518
R2353 VDD.n1584 VDD.n635 1.85518
R2354 VDD.n1584 VDD.n637 1.85518
R2355 VDD.n1584 VDD.n1583 1.85518
R2356 VDD.n910 VDD.n908 1.85344
R2357 VDD.n952 VDD.n908 1.85344
R2358 VDD.n1070 VDD.n1069 1.85344
R2359 VDD.n1071 VDD.n1070 1.85344
R2360 VDD.n1477 VDD.n1455 1.83567
R2361 VDD.n1473 VDD.n1455 1.83513
R2362 VDD.n1794 VDD.n535 1.835
R2363 VDD.n1798 VDD.n535 1.835
R2364 VDD.n1472 VDD.n1471 1.82979
R2365 VDD.n1471 VDD.n1470 1.82925
R2366 VDD.n1799 VDD.n536 1.82912
R2367 VDD.n537 VDD.n536 1.82912
R2368 VDD VDD.n926 1.82452
R2369 VDD.n1634 VDD.n603 1.80965
R2370 VDD.n1634 VDD.n1633 1.80912
R2371 VDD.n892 VDD.n869 1.7505
R2372 VDD.n2141 VDD.n2140 1.71333
R2373 VDD.n1492 VDD.n1491 1.69304
R2374 VDD.n1481 VDD.n1448 1.69304
R2375 VDD.n1459 VDD.n1458 1.69304
R2376 VDD.n1458 VDD.n732 1.69252
R2377 VDD.n1478 VDD.n1448 1.69252
R2378 VDD.n1493 VDD.n1492 1.69252
R2379 VDD.n1790 VDD.n534 1.69238
R2380 VDD.n1777 VDD.n531 1.69238
R2381 VDD.n1793 VDD.n534 1.69238
R2382 VDD.n1780 VDD.n531 1.69238
R2383 VDD.n1273 VDD.n1272 1.66029
R2384 VDD.n1272 VDD.n1271 1.65977
R2385 VDD.n1266 VDD.n815 1.65963
R2386 VDD.n1264 VDD.n1263 1.65963
R2387 VDD.n1258 VDD.n819 1.65963
R2388 VDD.n1256 VDD.n1255 1.65963
R2389 VDD.n1250 VDD.n823 1.65963
R2390 VDD.n1248 VDD.n1247 1.65963
R2391 VDD.n1242 VDD.n1241 1.65963
R2392 VDD.n815 VDD.n812 1.65963
R2393 VDD.n1265 VDD.n1264 1.65963
R2394 VDD.n819 VDD.n816 1.65963
R2395 VDD.n1257 VDD.n1256 1.65963
R2396 VDD.n823 VDD.n820 1.65963
R2397 VDD.n1249 VDD.n1248 1.65963
R2398 VDD.n1241 VDD.n824 1.65963
R2399 VDD.n125 VDD.n122 1.64018
R2400 VDD.n242 VDD.n239 1.64018
R2401 VDD.n62 VDD.t254 1.6255
R2402 VDD.n62 VDD.n61 1.6255
R2403 VDD.n77 VDD.t482 1.6255
R2404 VDD.n77 VDD.n76 1.6255
R2405 VDD.n69 VDD.t789 1.6255
R2406 VDD.n69 VDD.n68 1.6255
R2407 VDD.n71 VDD.t388 1.6255
R2408 VDD.n71 VDD.n70 1.6255
R2409 VDD.n167 VDD.t794 1.6255
R2410 VDD.n167 VDD.n166 1.6255
R2411 VDD.n169 VDD.t544 1.6255
R2412 VDD.n169 VDD.n168 1.6255
R2413 VDD.n184 VDD.t524 1.6255
R2414 VDD.n184 VDD.n183 1.6255
R2415 VDD.n186 VDD.t659 1.6255
R2416 VDD.n186 VDD.n185 1.6255
R2417 VDD.n160 VDD.t726 1.6255
R2418 VDD.n160 VDD.n159 1.6255
R2419 VDD.n162 VDD.t98 1.6255
R2420 VDD.n162 VDD.n161 1.6255
R2421 VDD.n149 VDD.t14 1.6255
R2422 VDD.n149 VDD.n148 1.6255
R2423 VDD.n298 VDD.t734 1.6255
R2424 VDD.n298 VDD.n297 1.6255
R2425 VDD.n296 VDD.t840 1.6255
R2426 VDD.n296 VDD.n295 1.6255
R2427 VDD.n277 VDD.t782 1.6255
R2428 VDD.n277 VDD.n276 1.6255
R2429 VDD.n286 VDD.t759 1.6255
R2430 VDD.n286 VDD.n285 1.6255
R2431 VDD.n289 VDD.t305 1.6255
R2432 VDD.n289 VDD.n288 1.6255
R2433 VDD.n313 VDD.t771 1.6255
R2434 VDD.n313 VDD.n312 1.6255
R2435 VDD.n311 VDD.t775 1.6255
R2436 VDD.n311 VDD.n310 1.6255
R2437 VDD.n362 VDD.t103 1.6255
R2438 VDD.n362 VDD.n361 1.6255
R2439 VDD.n360 VDD.t256 1.6255
R2440 VDD.n360 VDD.n359 1.6255
R2441 VDD.n368 VDD.t307 1.6255
R2442 VDD.n368 VDD.n367 1.6255
R2443 VDD.n377 VDD.t386 1.6255
R2444 VDD.n377 VDD.n376 1.6255
R2445 VDD.n382 VDD.t27 1.6255
R2446 VDD.n382 VDD.n381 1.6255
R2447 VDD.n354 VDD.t803 1.6255
R2448 VDD.n354 VDD.n353 1.6255
R2449 VDD.n352 VDD.t804 1.6255
R2450 VDD.n352 VDD.n351 1.6255
R2451 VDD.n108 VDD.t607 1.6255
R2452 VDD.n108 VDD.n107 1.6255
R2453 VDD.n110 VDD.t121 1.6255
R2454 VDD.n110 VDD.n109 1.6255
R2455 VDD.n86 VDD.t828 1.6255
R2456 VDD.n86 VDD.n85 1.6255
R2457 VDD.n1332 VDD.n784 1.5755
R2458 VDD.n1222 VDD.n1167 1.5755
R2459 VDD.n1864 VDD.n1863 1.5755
R2460 VDD.n1348 VDD.n1347 1.57159
R2461 VDD.n505 VDD.n504 1.57159
R2462 VDD.n1586 VDD.n1585 1.54574
R2463 VDD.n1745 VDD.n1744 1.52056
R2464 VDD.n1722 VDD.n582 1.52041
R2465 VDD.n1557 VDD.n627 1.52041
R2466 VDD.n1219 VDD.n1181 1.5005
R2467 VDD.n1365 VDD.n761 1.49724
R2468 VDD.n469 VDD.n420 1.49724
R2469 VDD.n1176 VDD.n1169 1.488
R2470 VDD.n214 VDD.n146 1.44912
R2471 VDD.n1162 VDD.n1161 1.42211
R2472 VDD.n1130 VDD.n1129 1.42018
R2473 VDD.n867 VDD.n842 1.4005
R2474 VDD.n1808 VDD.n1807 1.3744
R2475 VDD.n1805 VDD.n1804 1.3744
R2476 VDD.n1213 VDD.n1212 1.36849
R2477 VDD.n1721 VDD.n1702 1.35142
R2478 VDD.n2139 VDD.n2138 1.25782
R2479 VDD.t218 VDD.t152 1.24946
R2480 VDD.t147 VDD.t191 1.24946
R2481 VDD.n1128 VDD.n1080 1.2474
R2482 VDD.n79 VDD.n77 1.23637
R2483 VDD.n151 VDD.n149 1.23637
R2484 VDD.n279 VDD.n277 1.23591
R2485 VDD.n370 VDD.n368 1.23591
R2486 VDD.n2142 VDD.n2141 1.19777
R2487 VDD.n1807 VDD.n1806 1.1854
R2488 VDD.n1806 VDD.n1805 1.1854
R2489 VDD.n2032 VDD.n2031 1.17953
R2490 VDD.n1238 VDD.n1237 1.14837
R2491 VDD.n950 VDD.n949 1.1255
R2492 VDD.n872 VDD.n835 1.1255
R2493 VDD.n1006 VDD.n1005 1.1255
R2494 VDD.n1156 VDD.n1155 1.1255
R2495 VDD.n1219 VDD.n1218 1.1255
R2496 VDD.n1231 VDD.n1230 1.1255
R2497 VDD.n1010 VDD.n999 1.12549
R2498 VDD.n2014 VDD.n416 1.11762
R2499 VDD.n1744 VDD.n1743 1.08825
R2500 VDD.n1743 VDD.n582 1.08806
R2501 VDD.n1584 VDD.n627 1.08806
R2502 VDD.n1585 VDD.n1584 1.07146
R2503 VDD.n2031 VDD.n2024 1.06955
R2504 VDD.n1350 VDD.n1349 1.06485
R2505 VDD.n1361 VDD.n1360 1.06485
R2506 VDD.n1346 VDD.n1324 1.06485
R2507 VDD.n1343 VDD.n1342 1.06485
R2508 VDD.n507 VDD.n506 1.06485
R2509 VDD.n1873 VDD.n463 1.06485
R2510 VDD.n1866 VDD.n1865 1.06485
R2511 VDD.n1862 VDD.n1861 1.06485
R2512 VDD.n902 VDD.n889 1.0505
R2513 VDD.n1119 VDD.n1084 1.0505
R2514 VDD.n1365 VDD.n783 1.01789
R2515 VDD.n761 VDD.n751 1.01789
R2516 VDD.n469 VDD.n468 1.01789
R2517 VDD.n1857 VDD.n420 1.01789
R2518 VDD.n1589 VDD.n1588 0.984049
R2519 VDD.n897 VDD.n889 0.963
R2520 VDD.n1131 VDD.n1130 0.950899
R2521 VDD.n38 VDD.n37 0.93487
R2522 VDD.n1240 VDD.n1239 0.931466
R2523 VDD.n974 VDD.n973 0.927241
R2524 VDD.n831 VDD.n826 0.92659
R2525 VDD.n1081 VDD.n1079 0.925561
R2526 VDD.n989 VDD.n832 0.904541
R2527 VDD.n1078 VDD.n1077 0.899617
R2528 VDD.n945 VDD.n940 0.898206
R2529 VDD.n1151 VDD.n1131 0.897926
R2530 VDD.n1160 VDD.n990 0.897926
R2531 VDD.n57 VDD.n22 0.873239
R2532 VDD.n56 VDD.n55 0.847535
R2533 VDD.t200 VDD.t243 0.833139
R2534 VDD.t188 VDD.t200 0.833139
R2535 VDD.t206 VDD.t194 0.833139
R2536 VDD.t197 VDD.t238 0.833139
R2537 VDD.t238 VDD.t185 0.833139
R2538 VDD.n1237 VDD 0.830218
R2539 VDD.n1317 VDD.n1316 0.802674
R2540 VDD.n1356 VDD.n1353 0.802674
R2541 VDD.n1338 VDD.n1335 0.802674
R2542 VDD.n1345 VDD.n1344 0.802674
R2543 VDD.n494 VDD.n484 0.802674
R2544 VDD.n1872 VDD.n1869 0.802674
R2545 VDD.n503 VDD.n475 0.802674
R2546 VDD.n497 VDD.n481 0.802674
R2547 VDD.n142 VDD.n141 0.798761
R2548 VDD.n267 VDD.n266 0.798761
R2549 VDD.n345 VDD.n344 0.795258
R2550 VDD.n714 VDD.n713 0.795217
R2551 VDD.n1161 VDD.n1160 0.792748
R2552 VDD.n1272 VDD.n811 0.746922
R2553 VDD.n815 VDD.n811 0.746686
R2554 VDD.n1264 VDD.n811 0.746686
R2555 VDD.n819 VDD.n811 0.746686
R2556 VDD.n1256 VDD.n811 0.746686
R2557 VDD.n823 VDD.n811 0.746686
R2558 VDD.n1248 VDD.n811 0.746686
R2559 VDD.n1241 VDD.n811 0.746686
R2560 VDD.n46 VDD.n45 0.735716
R2561 VDD.n1448 VDD.n726 0.730547
R2562 VDD.n1458 VDD.n726 0.730547
R2563 VDD.n1492 VDD.n726 0.730547
R2564 VDD.n1806 VDD.n534 0.73031
R2565 VDD.n1806 VDD.n531 0.73031
R2566 VDD.n935 VDD.n934 0.7187
R2567 VDD.n1635 VDD.n1634 0.674731
R2568 VDD.n1471 VDD.n726 0.662176
R2569 VDD.n1806 VDD.n536 0.661938
R2570 VDD.n2017 VDD.n417 0.660673
R2571 VDD.n1455 VDD.n726 0.659239
R2572 VDD.n1806 VDD.n535 0.659
R2573 VDD.n1743 VDD.n580 0.645651
R2574 VDD VDD.n2 0.642616
R2575 VDD.n924 VDD.n923 0.6395
R2576 VDD.n1141 VDD.n1139 0.6395
R2577 VDD.n1136 VDD.n1134 0.6395
R2578 VDD.n2067 VDD.n2066 0.6395
R2579 VDD.n2121 VDD.n2119 0.6395
R2580 VDD.n346 VDD.n345 0.626871
R2581 VDD.n2046 VDD.n2045 0.622154
R2582 VDD.n862 VDD.n842 0.613
R2583 VDD.n1445 VDD.n726 0.60307
R2584 VDD.n1806 VDD.n533 0.602829
R2585 VDD.n2130 VDD.n2129 0.597767
R2586 VDD.n1747 VDD.n1746 0.593699
R2587 VDD.n2018 VDD.n416 0.587674
R2588 VDD VDD.n2047 0.582694
R2589 VDD.n1311 VDD.n1308 0.581587
R2590 VDD.n1320 VDD.n756 0.581587
R2591 VDD.n1373 VDD.n776 0.581587
R2592 VDD.n1323 VDD.n746 0.581587
R2593 VDD.n1838 VDD.n510 0.581587
R2594 VDD.n500 VDD.n426 0.581587
R2595 VDD.n1990 VDD.n445 0.581587
R2596 VDD.n1976 VDD.n1876 0.581587
R2597 VDD.n45 VDD.n43 0.576883
R2598 VDD.n1958 VDD.n1957 0.573969
R2599 VDD.n1701 VDD.n1695 0.569476
R2600 VDD.n1441 VDD.n726 0.553668
R2601 VDD.n1806 VDD.n532 0.553425
R2602 VDD.n22 VDD.n21 0.5405
R2603 VDD.n21 VDD.n20 0.5405
R2604 VDD.n1161 VDD.n989 0.539532
R2605 VDD.n273 VDD.n272 0.539417
R2606 VDD.n216 VDD.n145 0.538543
R2607 VDD.n218 VDD.n143 0.538543
R2608 VDD.n271 VDD.n270 0.536587
R2609 VDD.n1802 VDD.n545 0.536587
R2610 VDD.n552 VDD.n551 0.536587
R2611 VDD.n558 VDD.n557 0.536587
R2612 VDD.n1468 VDD.n1464 0.536587
R2613 VDD.n1454 VDD.n1453 0.536587
R2614 VDD.n1444 VDD.n1443 0.536587
R2615 VDD.n1176 VDD.n1166 0.5255
R2616 VDD.n347 VDD.n346 0.50421
R2617 VDD.n224 VDD.n125 0.502171
R2618 VDD.n243 VDD.n242 0.500214
R2619 VDD.n1718 VDD.n1703 0.495796
R2620 VDD.n2148 VDD.n2052 0.489544
R2621 VDD VDD.n879 0.485717
R2622 VDD VDD.n885 0.485717
R2623 VDD.n96 VDD.n79 0.476034
R2624 VDD.n212 VDD.n151 0.476034
R2625 VDD.n340 VDD.n279 0.475523
R2626 VDD.n374 VDD.n370 0.475523
R2627 VDD VDD.n601 0.474784
R2628 VDD.n1365 VDD.n1364 0.467817
R2629 VDD.n472 VDD.n469 0.467817
R2630 VDD.n1341 VDD.n751 0.466777
R2631 VDD.n1860 VDD.n1857 0.466777
R2632 VDD.n318 VDD.n317 0.464945
R2633 VDD.n191 VDD.n190 0.463664
R2634 VDD.n103 VDD.n102 0.463032
R2635 VDD.n176 VDD.n175 0.463032
R2636 VDD.n306 VDD.n305 0.463032
R2637 VDD.n405 VDD.n404 0.463032
R2638 VDD.n1129 VDD.n1128 0.462817
R2639 VDD.n9 VDD.n8 0.446529
R2640 VDD.n342 VDD 0.44179
R2641 VDD.n1353 VDD.n1350 0.440717
R2642 VDD.n1873 VDD.n1872 0.440717
R2643 VDD.n1226 VDD.n1167 0.438
R2644 VDD.n214 VDD 0.437942
R2645 VDD.n143 VDD.n142 0.430935
R2646 VDD.n270 VDD.n267 0.430935
R2647 VDD.n478 VDD.n420 0.430935
R2648 VDD.n1331 VDD.n761 0.430935
R2649 VDD.n1359 VDD.n783 0.430935
R2650 VDD.n468 VDD.n466 0.430935
R2651 VDD.n8 VDD.n7 0.429324
R2652 VDD.n7 VDD.n6 0.429324
R2653 VDD.n2048 VDD.n59 0.428242
R2654 VDD.n1360 VDD.n1356 0.421152
R2655 VDD.n1342 VDD.n1341 0.421152
R2656 VDD.n1869 VDD.n1866 0.421152
R2657 VDD.n1861 VDD.n1860 0.421152
R2658 VDD.n2135 VDD.n2091 0.419346
R2659 VDD.n2133 VDD.n2107 0.419346
R2660 VDD.n2131 VDD.n2130 0.419346
R2661 VDD.n2077 VDD.n2072 0.419346
R2662 VDD.n192 VDD.n187 0.419196
R2663 VDD.n319 VDD.n314 0.419196
R2664 VDD.n415 VDD.n355 0.419196
R2665 VDD.n349 VDD.n348 0.419196
R2666 VDD.n2034 VDD.n115 0.419196
R2667 VDD.n2036 VDD.n111 0.419196
R2668 VDD.t221 VDD.t149 0.41682
R2669 VDD.t149 VDD.t213 0.41682
R2670 VDD.t231 VDD.t182 0.41682
R2671 VDD.t572 VDD.n749 0.41682
R2672 VDD.t155 VDD.t203 0.41682
R2673 VDD.t226 VDD.t155 0.41682
R2674 VDD.n1523 VDD.n1522 0.405977
R2675 VDD.n1774 VDD.n560 0.405977
R2676 VDD.n2048 VDD 0.40579
R2677 VDD.n1366 VDD.n1365 0.394968
R2678 VDD.n1416 VDD.n751 0.394968
R2679 VDD.n469 VDD.n467 0.394968
R2680 VDD.n1857 VDD.n1856 0.394968
R2681 VDD.n2011 VDD.n420 0.39039
R2682 VDD.n1324 VDD.n1323 0.389848
R2683 VDD.n510 VDD.n507 0.389848
R2684 VDD.n672 VDD.n671 0.389323
R2685 VDD.n1201 VDD.n1200 0.389323
R2686 VDD.n1625 VDD.n1622 0.389323
R2687 VDD.n2112 VDD.n2110 0.389323
R2688 VDD.n2072 VDD.n2071 0.388557
R2689 VDD.n1678 VDD.n1644 0.376152
R2690 VDD.n1679 VDD.n1641 0.376152
R2691 VDD.n690 VDD.n652 0.376152
R2692 VDD.n914 VDD.n913 0.376152
R2693 VDD.n857 VDD.n852 0.376152
R2694 VDD.n1123 VDD.n1082 0.376152
R2695 VDD.n1034 VDD.n1030 0.376152
R2696 VDD.n1034 VDD.n1033 0.376152
R2697 VDD.n1612 VDD.n609 0.376152
R2698 VDD.n1670 VDD.n1654 0.374196
R2699 VDD.n679 VDD.n666 0.374196
R2700 VDD.n648 VDD.n647 0.374196
R2701 VDD.n1109 VDD.n1094 0.374196
R2702 VDD.n1056 VDD.n1050 0.374196
R2703 VDD.n1056 VDD.n1055 0.374196
R2704 VDD.n1208 VDD.n1195 0.374196
R2705 VDD.n619 VDD.n618 0.374196
R2706 VDD.n1688 VDD.n1635 0.372931
R2707 VDD.n1558 VDD.n714 0.359918
R2708 VDD.n1300 VDD.n783 0.358543
R2709 VDD.n1399 VDD.n761 0.358543
R2710 VDD.n468 VDD.n455 0.358543
R2711 VDD.n343 VDD.n342 0.357597
R2712 VDD.n1169 VDD.n1168 0.350287
R2713 VDD.n340 VDD.n339 0.334371
R2714 VDD.n344 VDD.n343 0.332919
R2715 VDD.n1348 VDD.n1317 0.327239
R2716 VDD.n504 VDD.n503 0.327239
R2717 VDD.n1335 VDD.n1324 0.323326
R2718 VDD.n1346 VDD.n1345 0.323326
R2719 VDD.n507 VDD.n494 0.323326
R2720 VDD.n506 VDD.n497 0.323326
R2721 VDD.n212 VDD.n211 0.32143
R2722 VDD.n690 VDD.n689 0.312794
R2723 VDD.n1863 VDD.n478 0.311587
R2724 VDD.n1332 VDD.n1331 0.311587
R2725 VDD.n1613 VDD.n1612 0.306039
R2726 VDD.n215 VDD.n214 0.305384
R2727 VDD.n58 VDD.n15 0.3007
R2728 VDD.n344 VDD.n259 0.292274
R2729 VDD.n345 VDD.n245 0.292274
R2730 VDD.n346 VDD.n235 0.292274
R2731 VDD.n347 VDD.n234 0.292274
R2732 VDD.n343 VDD.n273 0.292274
R2733 VDD.n1245 VDD.n825 0.292144
R2734 VDD.n1253 VDD.n821 0.292144
R2735 VDD.n1260 VDD.n817 0.292144
R2736 VDD.n1360 VDD.n1359 0.292022
R2737 VDD.n1364 VDD.n1361 0.292022
R2738 VDD.n1342 VDD.n1338 0.292022
R2739 VDD.n1344 VDD.n1343 0.292022
R2740 VDD.n1861 VDD.n484 0.292022
R2741 VDD.n1865 VDD.n472 0.292022
R2742 VDD.n1866 VDD.n466 0.292022
R2743 VDD.n1862 VDD.n481 0.292022
R2744 VDD.n1916 VDD.n1915 0.291683
R2745 VDD.n1928 VDD.n1909 0.291683
R2746 VDD.n1951 VDD.n1902 0.291683
R2747 VDD.n1268 VDD.n813 0.288544
R2748 VDD.n1941 VDD.n1934 0.288083
R2749 VDD.n1918 VDD.n1914 0.284207
R2750 VDD.n1316 VDD.n784 0.278326
R2751 VDD.n1864 VDD.n475 0.278326
R2752 VDD.n1350 VDD.n1311 0.272457
R2753 VDD.n1349 VDD.n776 0.272457
R2754 VDD.n463 VDD.n445 0.272457
R2755 VDD.n1876 VDD.n1873 0.272457
R2756 VDD.n1347 VDD.n1320 0.266587
R2757 VDD.n505 VDD.n500 0.266587
R2758 VDD.n1783 VDD.n559 0.266523
R2759 VDD.n1488 VDD.n1442 0.26536
R2760 VDD.n540 VDD.n538 0.264528
R2761 VDD.n1466 VDD.n1465 0.263373
R2762 VDD.n979 VDD.n869 0.263
R2763 VDD.n554 VDD.n553 0.262011
R2764 VDD.n1447 VDD.n1446 0.260887
R2765 VDD.n1796 VDD.n546 0.257984
R2766 VDD.n1475 VDD.n1456 0.257526
R2767 VDD.n1749 VDD.n1748 0.25389
R2768 VDD.n1175 VDD.n1174 0.253803
R2769 VDD.n1240 VDD.n805 0.252505
R2770 VDD.n937 VDD.n936 0.252091
R2771 VDD.n2024 VDD.n2023 0.251788
R2772 VDD.n1588 VDD.n623 0.248505
R2773 VDD.n101 VDD.n73 0.246576
R2774 VDD.n174 VDD.n171 0.246576
R2775 VDD.n304 VDD.n300 0.246576
R2776 VDD.n403 VDD.n364 0.246576
R2777 VDD.n102 VDD 0.245437
R2778 VDD.n175 VDD 0.245437
R2779 VDD.n305 VDD 0.245437
R2780 VDD.n404 VDD 0.245437
R2781 VDD.n1762 VDD.n573 0.238241
R2782 VDD.n1542 VDD.n1541 0.238069
R2783 VDD.n1540 VDD.n722 0.237294
R2784 VDD.n1661 VDD.n1659 0.237044
R2785 VDD.n1102 VDD.n1100 0.237044
R2786 VDD.n1593 VDD.n1592 0.237044
R2787 VDD.n856 VDD.n855 0.233429
R2788 VDD.n689 VDD.n655 0.229786
R2789 VDD.n944 VDD.n941 0.229786
R2790 VDD.n998 VDD.n997 0.229786
R2791 VDD.n1613 VDD.n608 0.229786
R2792 VDD.n221 VDD.n130 0.228829
R2793 VDD.n2023 VDD.n347 0.228403
R2794 VDD.n1507 VDD.n1506 0.221442
R2795 VDD.n1711 VDD.n1708 0.220495
R2796 VDD VDD.n2148 0.218882
R2797 VDD.n1130 VDD.n1078 0.217222
R2798 VDD.n2107 VDD 0.215115
R2799 VDD.n1276 VDD.n1275 0.209826
R2800 VDD.n1960 VDD.n1894 0.209826
R2801 VDD.n215 VDD.n144 0.209105
R2802 VDD.n228 VDD.n227 0.208053
R2803 VDD.n144 VDD.n130 0.19985
R2804 VDD.n2023 VDD.n2022 0.188845
R2805 VDD VDD.n318 0.186339
R2806 VDD.n1920 VDD.n1919 0.183919
R2807 VDD.n1103 VDD.n1097 0.182274
R2808 VDD.n2074 VDD.n2073 0.182274
R2809 VDD.n1660 VDD.n1658 0.182033
R2810 VDD.n687 VDD.n686 0.182033
R2811 VDD.n708 VDD.n640 0.182033
R2812 VDD.n1595 VDD.n1594 0.182033
R2813 VDD.n1616 VDD.n1615 0.182033
R2814 VDD VDD.n191 0.178694
R2815 VDD.n1773 VDD.n562 0.178585
R2816 VDD.n1499 VDD.n1495 0.17667
R2817 VDD.n1764 VDD.n526 0.176655
R2818 VDD.n1538 VDD.n723 0.176655
R2819 VDD.n2070 VDD 0.174184
R2820 VDD VDD.n2069 0.174184
R2821 VDD.n2128 VDD.n2126 0.174184
R2822 VDD.n713 VDD.n709 0.174122
R2823 VDD.n2123 VDD 0.173395
R2824 VDD.n1524 VDD.n1439 0.17241
R2825 VDD.n1822 VDD.n520 0.17241
R2826 VDD.n1816 VDD.n1815 0.171399
R2827 VDD.n1432 VDD.n730 0.171399
R2828 VDD.n1788 VDD.n1787 0.163357
R2829 VDD.n1484 VDD.n1483 0.163357
R2830 VDD.n2071 VDD.n2070 0.158395
R2831 VDD.n2129 VDD.n2128 0.158395
R2832 VDD.n1816 VDD.n515 0.157434
R2833 VDD.n331 VDD.n287 0.157274
R2834 VDD.n1433 VDD.n1432 0.15672
R2835 VDD VDD.n330 0.156548
R2836 VDD.n1277 VDD.n799 0.153197
R2837 VDD.n1962 VDD.n1961 0.153197
R2838 VDD.n164 VDD.n163 0.151198
R2839 VDD.n165 VDD 0.1505
R2840 VDD.n1914 VDD.n1886 0.146319
R2841 VDD.n1783 VDD.n1782 0.146214
R2842 VDD.n1489 VDD.n1488 0.146214
R2843 VDD.n1277 VDD.n1276 0.146118
R2844 VDD.n1961 VDD.n1960 0.146118
R2845 VDD.n1283 VDD.n805 0.146022
R2846 VDD.n1076 VDD.n1074 0.143441
R2847 VDD.n1533 VDD.n729 0.143084
R2848 VDD.n1784 VDD.n558 0.143
R2849 VDD.n1524 VDD.n1523 0.142944
R2850 VDD.n560 VDD.n520 0.142944
R2851 VDD.n2033 VDD.n2032 0.14289
R2852 VDD.n1500 VDD.n1499 0.142202
R2853 VDD.n564 VDD.n562 0.142202
R2854 VDD.n1813 VDD.n1812 0.142073
R2855 VDD.n1487 VDD.n1444 0.141929
R2856 VDD.n375 VDD.n374 0.141797
R2857 VDD.n1812 VDD.n526 0.141062
R2858 VDD.n729 VDD.n723 0.141062
R2859 VDD.n1800 VDD.n1797 0.140857
R2860 VDD.n1474 VDD.n1457 0.140857
R2861 VDD.n2143 VDD.n2058 0.140627
R2862 VDD.n1275 VDD.n808 0.14038
R2863 VDD.n1935 VDD.n1894 0.14038
R2864 VDD.n1801 VDD.n1800 0.139786
R2865 VDD.n1782 VDD.n1779 0.139786
R2866 VDD.n1489 VDD.n1440 0.139786
R2867 VDD.n1469 VDD.n1457 0.139786
R2868 VDD VDD.n935 0.139763
R2869 VDD.n1588 VDD.n1587 0.139295
R2870 VDD.n2031 VDD.n2030 0.1385
R2871 VDD.n1587 VDD.n624 0.138211
R2872 VDD.n1720 VDD.n1718 0.138211
R2873 VDD.n1796 VDD.n1795 0.137643
R2874 VDD.n1476 VDD.n1475 0.137643
R2875 VDD.n1823 VDD.n1822 0.137017
R2876 VDD.n1439 VDD.n1438 0.136006
R2877 VDD.n2123 VDD.n2122 0.1355
R2878 VDD.n2137 VDD.n2079 0.1355
R2879 VDD.n2069 VDD.n2068 0.134711
R2880 VDD.n1746 VDD.n578 0.133873
R2881 VDD.n1740 VDD.n1739 0.133873
R2882 VDD.n1737 VDD.n1735 0.133873
R2883 VDD.n1733 VDD.n1731 0.133873
R2884 VDD.n1729 VDD.n1727 0.133873
R2885 VDD.n1725 VDD.n1723 0.133873
R2886 VDD.n1581 VDD.n624 0.133873
R2887 VDD.n1580 VDD.n1578 0.133873
R2888 VDD.n1576 VDD.n1574 0.133873
R2889 VDD.n1572 VDD.n1570 0.133873
R2890 VDD.n1568 VDD.n1566 0.133873
R2891 VDD.n1564 VDD.n1562 0.133873
R2892 VDD.n1560 VDD.n1558 0.133873
R2893 VDD.n1751 VDD.n1750 0.133833
R2894 VDD.n576 VDD.n574 0.133833
R2895 VDD.n1761 VDD.n574 0.133833
R2896 VDD.n1764 VDD.n1763 0.133833
R2897 VDD.n1539 VDD.n1538 0.133833
R2898 VDD.n1545 VDD.n1544 0.133833
R2899 VDD.n1544 VDD.n1543 0.133833
R2900 VDD.n1554 VDD.n716 0.133833
R2901 VDD.n1810 VDD.n525 0.133132
R2902 VDD.n971 VDD 0.131587
R2903 VDD.n1517 VDD.n1500 0.131498
R2904 VDD.n565 VDD.n564 0.13055
R2905 VDD.n1476 VDD.n1454 0.130143
R2906 VDD.n970 VDD 0.12963
R2907 VDD.n1270 VDD.n808 0.129536
R2908 VDD.n1270 VDD.n1269 0.129536
R2909 VDD.n1267 VDD.n814 0.129536
R2910 VDD.n1262 VDD.n814 0.129536
R2911 VDD.n1262 VDD.n1261 0.129536
R2912 VDD.n1259 VDD.n818 0.129536
R2913 VDD.n1254 VDD.n818 0.129536
R2914 VDD.n1252 VDD.n1251 0.129536
R2915 VDD.n1251 VDD.n822 0.129536
R2916 VDD.n1246 VDD.n822 0.129536
R2917 VDD.n1244 VDD.n1243 0.129536
R2918 VDD.n1918 VDD.n1917 0.129536
R2919 VDD.n1912 VDD.n1910 0.129536
R2920 VDD.n1926 VDD.n1910 0.129536
R2921 VDD.n1927 VDD.n1926 0.129536
R2922 VDD.n1929 VDD.n1901 0.129536
R2923 VDD.n1952 VDD.n1901 0.129536
R2924 VDD.n1950 VDD.n1949 0.129536
R2925 VDD.n1949 VDD.n1903 0.129536
R2926 VDD.n1942 VDD.n1903 0.129536
R2927 VDD.n1940 VDD.n1939 0.129536
R2928 VDD.n1939 VDD.n1935 0.129536
R2929 VDD.n1121 VDD.n1084 0.129141
R2930 VDD.n1795 VDD.n552 0.129071
R2931 VDD.n2079 VDD.n2078 0.128577
R2932 VDD.n1500 VDD.n1498 0.128395
R2933 VDD.n564 VDD.n563 0.128395
R2934 VDD.n1739 VDD.n1737 0.127367
R2935 VDD.n1735 VDD.n1733 0.127367
R2936 VDD.n1731 VDD.n1729 0.127367
R2937 VDD.n1727 VDD.n1725 0.127367
R2938 VDD.n1245 VDD.n1244 0.127367
R2939 VDD.n1581 VDD.n1580 0.127367
R2940 VDD.n1578 VDD.n1576 0.127367
R2941 VDD.n1574 VDD.n1572 0.127367
R2942 VDD.n1570 VDD.n1568 0.127367
R2943 VDD.n1566 VDD.n1564 0.127367
R2944 VDD.n1917 VDD.n1916 0.127367
R2945 VDD.n2140 VDD.n2139 0.12616
R2946 VDD.n1073 VDD.n996 0.126143
R2947 VDD.n1740 VDD.n578 0.124114
R2948 VDD.n1562 VDD.n1560 0.124114
R2949 VDD.n1516 VDD.n1515 0.123227
R2950 VDD.n1515 VDD.n1501 0.123227
R2951 VDD.n1509 VDD.n1508 0.123227
R2952 VDD.n1508 VDD.n623 0.123227
R2953 VDD.n1707 VDD.n1703 0.123227
R2954 VDD.n1712 VDD.n1707 0.123227
R2955 VDD.n1710 VDD.n1709 0.123227
R2956 VDD.n1709 VDD.n567 0.123227
R2957 VDD.n1260 VDD.n1259 0.12303
R2958 VDD.n1952 VDD.n1951 0.12303
R2959 VDD.n1507 VDD.n1501 0.122205
R2960 VDD.n1711 VDD.n1710 0.122205
R2961 VDD.n1290 VDD.n799 0.120837
R2962 VDD.n1291 VDD.n1290 0.120837
R2963 VDD.n1292 VDD.n1291 0.120837
R2964 VDD.n1292 VDD.n785 0.120837
R2965 VDD.n1307 VDD.n786 0.120837
R2966 VDD.n786 VDD.n777 0.120837
R2967 VDD.n1372 VDD.n777 0.120837
R2968 VDD.n1375 VDD.n1374 0.120837
R2969 VDD.n1375 VDD.n766 0.120837
R2970 VDD.n1388 VDD.n766 0.120837
R2971 VDD.n1389 VDD.n1388 0.120837
R2972 VDD.n1391 VDD.n1389 0.120837
R2973 VDD.n1391 VDD.n1390 0.120837
R2974 VDD.n1406 VDD.n1405 0.120837
R2975 VDD.n1408 VDD.n1406 0.120837
R2976 VDD.n1408 VDD.n1407 0.120837
R2977 VDD.n1423 VDD.n1422 0.120837
R2978 VDD.n1424 VDD.n1423 0.120837
R2979 VDD.n1424 VDD.n737 0.120837
R2980 VDD.n1438 VDD.n737 0.120837
R2981 VDD.n1824 VDD.n1823 0.120837
R2982 VDD.n1824 VDD.n511 0.120837
R2983 VDD.n1836 VDD.n511 0.120837
R2984 VDD.n1837 VDD.n1836 0.120837
R2985 VDD.n1850 VDD.n1849 0.120837
R2986 VDD.n1849 VDD.n1848 0.120837
R2987 VDD.n1848 VDD.n1839 0.120837
R2988 VDD.n2006 VDD.n2005 0.120837
R2989 VDD.n2005 VDD.n2004 0.120837
R2990 VDD.n2004 VDD.n427 0.120837
R2991 VDD.n442 VDD.n427 0.120837
R2992 VDD.n1992 VDD.n442 0.120837
R2993 VDD.n1992 VDD.n1991 0.120837
R2994 VDD.n1989 VDD.n446 0.120837
R2995 VDD.n462 VDD.n446 0.120837
R2996 VDD.n1977 VDD.n462 0.120837
R2997 VDD.n1975 VDD.n1974 0.120837
R2998 VDD.n1974 VDD.n1877 0.120837
R2999 VDD.n1893 VDD.n1877 0.120837
R3000 VDD.n1962 VDD.n1893 0.120837
R3001 VDD.n1555 VDD.n714 0.119037
R3002 VDD.n539 VDD.n524 0.117286
R3003 VDD.n1792 VDD.n1791 0.117286
R3004 VDD.n1779 VDD.n1778 0.117286
R3005 VDD.n1494 VDD.n1440 0.117286
R3006 VDD.n1480 VDD.n1479 0.117286
R3007 VDD.n1531 VDD.n731 0.117286
R3008 VDD.n254 VDD.n253 0.115972
R3009 VDD.n244 VDD.n243 0.115972
R3010 VDD.n2057 VDD.n2056 0.115087
R3011 VDD.n273 VDD.n271 0.113142
R3012 VDD.n309 VDD.n308 0.113
R3013 VDD.n1518 VDD.n1517 0.113
R3014 VDD.n1772 VDD.n565 0.111977
R3015 VDD.n1308 VDD.n1307 0.110725
R3016 VDD.n243 VDD.n235 0.109745
R3017 VDD.n96 VDD.n95 0.109735
R3018 VDD.n1977 VDD.n1976 0.109713
R3019 VDD.n1814 VDD.n524 0.108714
R3020 VDD.n182 VDD.n181 0.10864
R3021 VDD.n2135 VDD.n2134 0.108385
R3022 VDD.n2144 VDD.n2143 0.108044
R3023 VDD.n1468 VDD.n1467 0.107643
R3024 VDD.n1532 VDD.n1531 0.107643
R3025 VDD.n1128 VDD.n1127 0.106797
R3026 VDD.n1803 VDD.n1802 0.106571
R3027 VDD.n1850 VDD.n1838 0.103646
R3028 VDD.n287 VDD.n282 0.103565
R3029 VDD.n1407 VDD.n746 0.102635
R3030 VDD.n2013 VDD.n2012 0.101533
R3031 VDD.n1232 VDD.n831 0.101088
R3032 VDD.n1284 VDD.n1283 0.1005
R3033 VDD.n1967 VDD.n1886 0.1005
R3034 VDD.n163 VDD.n154 0.0995698
R3035 VDD.n259 VDD.n258 0.0989906
R3036 VDD.n2133 VDD.n2132 0.0985769
R3037 VDD.n1763 VDD.n1762 0.0971667
R3038 VDD.n1540 VDD.n1539 0.0971667
R3039 VDD.n250 VDD.n245 0.0964434
R3040 VDD.n341 VDD.n340 0.0955806
R3041 VDD.n540 VDD.n539 0.0947857
R3042 VDD.n1466 VDD.n731 0.0947857
R3043 VDD.n1533 VDD.n1532 0.0945449
R3044 VDD.n1751 VDD.n1747 0.0938198
R3045 VDD.n1555 VDD.n1554 0.0938198
R3046 VDD.n1814 VDD.n1813 0.0935337
R3047 VDD.n338 VDD.n337 0.0919516
R3048 VDD.n337 VDD.n282 0.0919516
R3049 VDD.n329 VDD.n328 0.0919516
R3050 VDD.n328 VDD.n290 0.0919516
R3051 VDD.n321 VDD.n309 0.0919516
R3052 VDD.n321 VDD.n320 0.0919516
R3053 VDD.n213 VDD.n212 0.0918953
R3054 VDD.n12 VDD.n11 0.0914091
R3055 VDD.n11 VDD.n10 0.0914091
R3056 VDD.n36 VDD.n35 0.0914091
R3057 VDD.n35 VDD.n34 0.0914091
R3058 VDD.n34 VDD.n33 0.0914091
R3059 VDD.n33 VDD.n32 0.0914091
R3060 VDD.n32 VDD.n31 0.0914091
R3061 VDD.n31 VDD.n30 0.0914091
R3062 VDD VDD.n14 0.0900455
R3063 VDD.n925 VDD.n924 0.0893158
R3064 VDD.n1142 VDD.n1136 0.0893158
R3065 VDD.n1142 VDD.n1141 0.0893158
R3066 VDD.n2068 VDD.n2067 0.0893158
R3067 VDD.n2122 VDD.n2121 0.0893158
R3068 VDD.n1522 VDD.n1495 0.0884545
R3069 VDD.n210 VDD.n209 0.088407
R3070 VDD.n209 VDD.n154 0.088407
R3071 VDD.n202 VDD.n201 0.088407
R3072 VDD.n201 VDD.n200 0.088407
R3073 VDD.n194 VDD.n182 0.088407
R3074 VDD.n194 VDD.n193 0.088407
R3075 VDD.n1214 VDD.n1188 0.088
R3076 VDD.n307 VDD.n290 0.0875968
R3077 VDD.n1405 VDD.n756 0.0874663
R3078 VDD.n1774 VDD.n1773 0.0874318
R3079 VDD.n2056 VDD.n2053 0.0865195
R3080 VDD.n1839 VDD.n426 0.0864551
R3081 VDD.n1749 VDD.n576 0.0860556
R3082 VDD.n1543 VDD.n1542 0.0860556
R3083 VDD.n1829 VDD.n515 0.0855
R3084 VDD.n1830 VDD.n1829 0.0855
R3085 VDD.n1831 VDD.n1830 0.0855
R3086 VDD.n1831 VDD.n485 0.0855
R3087 VDD.n1855 VDD.n486 0.0855
R3088 VDD.n1842 VDD.n486 0.0855
R3089 VDD.n1842 VDD.n418 0.0855
R3090 VDD.n1285 VDD.n1284 0.0855
R3091 VDD.n1285 VDD.n796 0.0855
R3092 VDD.n1298 VDD.n796 0.0855
R3093 VDD.n1299 VDD.n1298 0.0855
R3094 VDD.n1302 VDD.n1301 0.0855
R3095 VDD.n1301 VDD.n782 0.0855
R3096 VDD.n1367 VDD.n782 0.0855
R3097 VDD.n1381 VDD.n771 0.0855
R3098 VDD.n1382 VDD.n1381 0.0855
R3099 VDD.n1383 VDD.n762 0.0855
R3100 VDD.n1397 VDD.n762 0.0855
R3101 VDD.n1398 VDD.n1397 0.0855
R3102 VDD.n1400 VDD.n752 0.0855
R3103 VDD.n1414 VDD.n752 0.0855
R3104 VDD.n1415 VDD.n1414 0.0855
R3105 VDD.n1417 VDD.n742 0.0855
R3106 VDD.n1430 VDD.n742 0.0855
R3107 VDD.n1431 VDD.n1430 0.0855
R3108 VDD.n1433 VDD.n1431 0.0855
R3109 VDD.n435 VDD.n419 0.0855
R3110 VDD.n1999 VDD.n435 0.0855
R3111 VDD.n1998 VDD.n1997 0.0855
R3112 VDD.n1997 VDD.n436 0.0855
R3113 VDD.n1984 VDD.n454 0.0855
R3114 VDD.n1984 VDD.n1983 0.0855
R3115 VDD.n1983 VDD.n1982 0.0855
R3116 VDD.n1885 VDD.n1884 0.0855
R3117 VDD.n1969 VDD.n1885 0.0855
R3118 VDD.n1969 VDD.n1968 0.0855
R3119 VDD.n1968 VDD.n1967 0.0855
R3120 VDD.n225 VDD.n224 0.0853962
R3121 VDD.n1269 VDD.n1268 0.0850783
R3122 VDD.n1941 VDD.n1940 0.0850783
R3123 VDD.n1302 VDD.n1300 0.0847857
R3124 VDD.n200 VDD.n177 0.0842209
R3125 VDD.n1982 VDD.n455 0.0840714
R3126 VDD.n928 VDD 0.0836933
R3127 VDD.n319 VDD 0.0832419
R3128 VDD.n1723 VDD.n1721 0.0818253
R3129 VDD.n224 VDD.n223 0.0817389
R3130 VDD.n223 VDD.n222 0.0817389
R3131 VDD.n258 VDD 0.0811604
R3132 VDD.n1990 VDD.n1989 0.0803876
R3133 VDD.n192 VDD 0.0800349
R3134 VDD VDD.n2027 0.0798636
R3135 VDD.n1373 VDD.n1372 0.0793764
R3136 VDD.n1152 VDD.n992 0.0790106
R3137 VDD.n2029 VDD 0.0778182
R3138 VDD.n1143 VDD 0.0774922
R3139 VDD.n1815 VDD.n1814 0.0773539
R3140 VDD.n1532 VDD.n730 0.0773539
R3141 VDD.n1788 VDD.n554 0.0765714
R3142 VDD.n1483 VDD.n1447 0.0765714
R3143 VDD.n1753 VDD.n1752 0.0752312
R3144 VDD.n10 VDD.n9 0.0750455
R3145 VDD.n1553 VDD.n715 0.074985
R3146 VDD.n1254 VDD.n1253 0.0742349
R3147 VDD.n1929 VDD.n1928 0.0742349
R3148 VDD.n1076 VDD.n1075 0.07388
R3149 VDD.n1721 VDD.n1720 0.0731506
R3150 VDD.n948 VDD.n917 0.0717174
R3151 VDD.n947 VDD.n946 0.0717174
R3152 VDD.n1672 VDD.n1645 0.0714756
R3153 VDD.n1681 VDD.n1636 0.0714756
R3154 VDD.n677 VDD.n668 0.0714756
R3155 VDD.n696 VDD.n695 0.0714756
R3156 VDD.n1117 VDD.n1116 0.0714756
R3157 VDD.n1199 VDD.n1196 0.0714756
R3158 VDD.n1606 VDD.n610 0.0714756
R3159 VDD.n1627 VDD.n1626 0.0714756
R3160 VDD.n1689 VDD.n592 0.0714756
R3161 VDD.n2101 VDD.n2100 0.0714756
R3162 VDD.n1154 VDD.n1153 0.0714615
R3163 VDD.n1671 VDD 0.0713871
R3164 VDD VDD.n678 0.0713871
R3165 VDD.n697 VDD 0.0713871
R3166 VDD VDD.n1086 0.0713871
R3167 VDD VDD.n1207 0.0713871
R3168 VDD.n1605 VDD 0.0713871
R3169 VDD.n1669 VDD.n1655 0.0709032
R3170 VDD.n1663 VDD.n1662 0.0709032
R3171 VDD.n658 VDD.n656 0.0709032
R3172 VDD.n680 VDD.n661 0.0709032
R3173 VDD.n705 VDD.n639 0.0709032
R3174 VDD.n704 VDD.n703 0.0709032
R3175 VDD.n1101 VDD.n1095 0.0709032
R3176 VDD.n1108 VDD.n1107 0.0709032
R3177 VDD.n1597 VDD.n1596 0.0709032
R3178 VDD.n1599 VDD.n1598 0.0709032
R3179 VDD.n605 VDD.n602 0.0709032
R3180 VDD.n1209 VDD.n1187 0.0701774
R3181 VDD.n1677 VDD.n1645 0.0692805
R3182 VDD.n1672 VDD.n1671 0.0692805
R3183 VDD.n1681 VDD.n1680 0.0692805
R3184 VDD.n1687 VDD.n1636 0.0692805
R3185 VDD.n678 VDD.n677 0.0692805
R3186 VDD.n672 VDD.n668 0.0692805
R3187 VDD.n697 VDD.n696 0.0692805
R3188 VDD.n695 VDD.n691 0.0692805
R3189 VDD.n1116 VDD.n1086 0.0692805
R3190 VDD.n1207 VDD.n1196 0.0692805
R3191 VDD.n1201 VDD.n1199 0.0692805
R3192 VDD.n1606 VDD.n1605 0.0692805
R3193 VDD.n1611 VDD.n610 0.0692805
R3194 VDD.n1627 VDD.n596 0.0692805
R3195 VDD.n1626 VDD.n1625 0.0692805
R3196 VDD.n1689 VDD 0.0692805
R3197 VDD.n2115 VDD.n2112 0.0692805
R3198 VDD.n2097 VDD.n2094 0.0692805
R3199 VDD VDD.n2101 0.0692805
R3200 VDD.n2052 VDD.n2049 0.0692083
R3201 VDD.n1663 VDD.n1655 0.0687258
R3202 VDD.n1662 VDD.n1661 0.0687258
R3203 VDD.n688 VDD.n656 0.0687258
R3204 VDD.n661 VDD.n658 0.0687258
R3205 VDD.n709 VDD.n639 0.0687258
R3206 VDD.n705 VDD.n704 0.0687258
R3207 VDD.n1102 VDD.n1101 0.0687258
R3208 VDD.n1107 VDD.n1095 0.0687258
R3209 VDD.n1599 VDD.n1597 0.0687258
R3210 VDD.n1614 VDD.n605 0.0687258
R3211 VDD.n2138 VDD.n2137 0.0685545
R3212 VDD.n1400 VDD.n1399 0.0683571
R3213 VDD.n226 VDD.n225 0.0676691
R3214 VDD.n2019 VDD.n350 0.0674625
R3215 VDD.n2142 VDD.n2059 0.0669557
R3216 VDD.n976 VDD.n871 0.0669486
R3217 VDD.n975 VDD.n974 0.0669486
R3218 VDD.n391 VDD.n378 0.0668481
R3219 VDD.n1534 VDD.n727 0.0668158
R3220 VDD VDD.n390 0.066541
R3221 VDD.n1856 VDD.n1855 0.0662143
R3222 VDD.n1416 VDD.n1415 0.0662143
R3223 VDD.n987 VDD.n986 0.0661075
R3224 VDD.n988 VDD.n833 0.0661075
R3225 VDD.n928 VDD.n925 0.0647857
R3226 VDD.n1158 VDD.n1157 0.0646489
R3227 VDD.n222 VDD.n221 0.0643765
R3228 VDD.n2131 VDD.n2116 0.0639615
R3229 VDD.n2133 VDD.n2106 0.0639615
R3230 VDD.n2135 VDD.n2090 0.0639615
R3231 VDD.n2077 VDD.n2076 0.0639615
R3232 VDD.n1670 VDD.n1669 0.0629194
R3233 VDD.n680 VDD.n679 0.0629194
R3234 VDD.n703 VDD.n648 0.0629194
R3235 VDD.n1109 VDD.n1108 0.0629194
R3236 VDD.n1209 VDD.n1208 0.0629194
R3237 VDD.n1598 VDD.n619 0.0629194
R3238 VDD VDD.n2091 0.0616538
R3239 VDD.n1143 VDD.n1142 0.0606172
R3240 VDD.n1118 VDD.n1117 0.0605
R3241 VDD.n1635 VDD.n596 0.0605
R3242 VDD.n216 VDD.n215 0.0603822
R3243 VDD.n2055 VDD.n2054 0.0593952
R3244 VDD.n1159 VDD.n991 0.0584808
R3245 VDD VDD.n234 0.0582358
R3246 VDD VDD.n2035 0.0570172
R3247 VDD.n2106 VDD.n2097 0.0561098
R3248 VDD.n1253 VDD.n1252 0.0558012
R3249 VDD.n1928 VDD.n1927 0.0558012
R3250 VDD VDD.n1688 0.055378
R3251 VDD.n2076 VDD.n2075 0.055378
R3252 VDD.n219 VDD.n130 0.0549355
R3253 VDD.n217 VDD.n144 0.0542097
R3254 VDD.n217 VDD.n216 0.0538628
R3255 VDD.n1185 VDD.n1184 0.0534412
R3256 VDD.n1182 VDD.n1163 0.0534412
R3257 VDD.n1361 VDD.n784 0.0533261
R3258 VDD.n1865 VDD.n1864 0.0533261
R3259 VDD.n220 VDD.n219 0.0530664
R3260 VDD.n1523 VDD.n1494 0.053
R3261 VDD.n1701 VDD.n592 0.0524512
R3262 VDD.n234 VDD.n233 0.0522925
R3263 VDD.n1778 VDD.n560 0.0519286
R3264 VDD.n59 VDD.n14 0.0518636
R3265 VDD.n919 VDD.n918 0.0509
R3266 VDD.n1150 VDD.n993 0.0504219
R3267 VDD.n1635 VDD.n602 0.0498548
R3268 VDD.n1367 VDD.n1366 0.0497857
R3269 VDD.n467 VDD.n454 0.0497857
R3270 VDD.n1999 VDD 0.0483571
R3271 VDD.n1750 VDD.n1749 0.0482778
R3272 VDD.n1542 VDD.n716 0.0482778
R3273 VDD.n408 VDD.n407 0.0481109
R3274 VDD.n1383 VDD 0.0462143
R3275 VDD.n937 VDD.n919 0.0458103
R3276 VDD.n1268 VDD.n1267 0.0449578
R3277 VDD.n1942 VDD.n1941 0.0449578
R3278 VDD.n396 VDD.n378 0.0441177
R3279 VDD.n231 VDD 0.0440029
R3280 VDD.n1374 VDD.n1373 0.0419607
R3281 VDD.n2016 VDD.n416 0.0414381
R3282 VDD.n2012 VDD.n418 0.0412143
R3283 VDD.n1791 VDD.n554 0.0412143
R3284 VDD.n1784 VDD.n1783 0.0412143
R3285 VDD.n1488 VDD.n1487 0.0412143
R3286 VDD.n1480 VDD.n1447 0.0412143
R3287 VDD.n1228 VDD.n1227 0.0411452
R3288 VDD.n1991 VDD.n1990 0.0409494
R3289 VDD.n1234 VDD.n829 0.0408043
R3290 VDD.n374 VDD.n373 0.0407389
R3291 VDD.n2032 VDD.n231 0.0401282
R3292 VDD VDD.n1382 0.0397857
R3293 VDD.n1243 VDD.n1240 0.0395361
R3294 VDD.n1239 VDD 0.0393983
R3295 VDD.n398 VDD.n397 0.0392031
R3296 VDD.n397 VDD.n396 0.0392031
R3297 VDD.n389 VDD.n388 0.0392031
R3298 VDD.n388 VDD.n358 0.0392031
R3299 VDD.n408 VDD.n356 0.0392031
R3300 VDD.n414 VDD.n356 0.0392031
R3301 VDD.n227 VDD.n226 0.0391413
R3302 VDD.n320 VDD.n319 0.0389677
R3303 VDD VDD.n1998 0.0376429
R3304 VDD.n1076 VDD.n996 0.0375588
R3305 VDD.n1593 VDD.n1589 0.0375161
R3306 VDD.n193 VDD.n192 0.0374767
R3307 VDD.n406 VDD.n358 0.0373601
R3308 VDD.n106 VDD.n105 0.0373074
R3309 VDD.n1762 VDD.n1761 0.0371667
R3310 VDD.n1545 VDD.n1540 0.0371667
R3311 VDD.n2012 VDD.n419 0.0369286
R3312 VDD.n713 VDD.n712 0.0369005
R3313 VDD.n1146 VDD.n1145 0.0367109
R3314 VDD.n2030 VDD.n2029 0.0363784
R3315 VDD.n1773 VDD.n1772 0.0362955
R3316 VDD.n1366 VDD.n771 0.0362143
R3317 VDD.n467 VDD.n436 0.0362143
R3318 VDD.n1039 VDD.n1024 0.0359878
R3319 VDD VDD.n1045 0.0359436
R3320 VDD.n1021 VDD.n1018 0.0357016
R3321 VDD.n1066 VDD.n1065 0.0357016
R3322 VDD.n2047 VDD.n63 0.0356451
R3323 VDD VDD.n415 0.0355171
R3324 VDD.n2024 VDD.n233 0.0353113
R3325 VDD VDD.n250 0.0353113
R3326 VDD.n1518 VDD.n1495 0.0352727
R3327 VDD.n1039 VDD.n1035 0.0348902
R3328 VDD.n1045 VDD.n1024 0.0348902
R3329 VDD.n2006 VDD.n426 0.034882
R3330 VDD.n1802 VDD.n1801 0.0347857
R3331 VDD.n1065 VDD.n1018 0.0346129
R3332 VDD.n82 VDD.n63 0.0342203
R3333 VDD.n1008 VDD.n1007 0.0340503
R3334 VDD.n1390 VDD.n756 0.0338708
R3335 VDD.n1347 VDD.n1346 0.0337609
R3336 VDD.n506 VDD.n505 0.0337609
R3337 VDD.n1469 VDD.n1468 0.0337143
R3338 VDD.n1003 VDD.n995 0.0335178
R3339 VDD.n1160 VDD.n1159 0.0331389
R3340 VDD.n2132 VDD.n2131 0.0328077
R3341 VDD.n2090 VDD.n2089 0.0326951
R3342 VDD.n1153 VDD.n1131 0.0322736
R3343 VDD.n1056 VDD.n1021 0.0317097
R3344 VDD.n1596 VDD.n1589 0.0317097
R3345 VDD.n97 VDD.n96 0.0316082
R3346 VDD.n2116 VDD.n2115 0.0305
R3347 VDD.n2134 VDD.n2133 0.0305
R3348 VDD.n2038 VDD.n106 0.0304208
R3349 VDD.n2038 VDD.n2037 0.0304208
R3350 VDD.n94 VDD.n81 0.0304208
R3351 VDD.n82 VDD.n81 0.0304208
R3352 VDD.n1158 VDD.n990 0.0301809
R3353 VDD.n940 VDD.n917 0.0299176
R3354 VDD.n1152 VDD.n1151 0.0292234
R3355 VDD.n1156 VDD.n992 0.0292234
R3356 VDD.n1157 VDD.n1156 0.0292234
R3357 VDD.n1520 VDD.n1519 0.0291956
R3358 VDD.n1505 VDD.n1504 0.0291956
R3359 VDD.n1715 VDD.n1704 0.0291956
R3360 VDD.n1771 VDD.n561 0.0291956
R3361 VDD.n219 VDD.n218 0.0291726
R3362 VDD.n104 VDD.n60 0.028996
R3363 VDD.n961 VDD.n904 0.0289211
R3364 VDD.n960 VDD.n959 0.0289211
R3365 VDD.n39 VDD.n38 0.028625
R3366 VDD.n218 VDD.n217 0.0283761
R3367 VDD.n339 VDD.n338 0.0280806
R3368 VDD.n1232 VDD.n1231 0.0278529
R3369 VDD.n1218 VDD.n1185 0.0278529
R3370 VDD.n1009 VDD.n1002 0.0277596
R3371 VDD.n2136 VDD.n2135 0.0276154
R3372 VDD.n2036 VDD 0.0275712
R3373 VDD.n2047 VDD.n2046 0.0274032
R3374 VDD.n1004 VDD.n994 0.0273269
R3375 VDD.n1702 VDD.n591 0.0270909
R3376 VDD.n211 VDD.n210 0.0270116
R3377 VDD.n872 VDD.n833 0.0265748
R3378 VDD.n1155 VDD.n1154 0.0264615
R3379 VDD.n1155 VDD.n991 0.0264615
R3380 VDD.n54 VDD.n48 0.026375
R3381 VDD.n975 VDD.n872 0.0257336
R3382 VDD.n958 VDD.n907 0.0256417
R3383 VDD.n2047 VDD.n60 0.025434
R3384 VDD.n330 VDD.n329 0.0251774
R3385 VDD.n1066 VDD.n1000 0.0251774
R3386 VDD.n350 VDD.n349 0.0250734
R3387 VDD.n1235 VDD.n828 0.0247707
R3388 VDD.n946 VDD.n945 0.0247609
R3389 VDD.n202 VDD.n165 0.0242209
R3390 VDD.n1349 VDD.n1348 0.0239783
R3391 VDD.n949 VDD.n948 0.0239783
R3392 VDD.n504 VDD.n463 0.0239783
R3393 VDD.n2014 VDD.n2013 0.0237036
R3394 VDD.n1012 VDD.n1011 0.0235488
R3395 VDD.n970 VDD.n880 0.0234555
R3396 VDD.n1231 VDD.n1162 0.0234412
R3397 VDD.n1803 VDD.n540 0.023
R3398 VDD.n1484 VDD.n1444 0.023
R3399 VDD.n1467 VDD.n1466 0.023
R3400 VDD.n984 VDD.n836 0.0227267
R3401 VDD.n1220 VDD.n1219 0.0225588
R3402 VDD.n1217 VDD.n1183 0.0225588
R3403 VDD.n857 VDD.n856 0.0223623
R3404 VDD.n1787 VDD.n558 0.0219286
R3405 VDD.n891 VDD.n890 0.0216336
R3406 VDD.n989 VDD.n988 0.0206869
R3407 VDD.n2100 VDD.n2090 0.0202561
R3408 VDD.n916 VDD.n912 0.0200652
R3409 VDD.n950 VDD.n915 0.0200652
R3410 VDD.n1343 VDD.n1332 0.0200652
R3411 VDD.n1863 VDD.n1862 0.0200652
R3412 VDD.n245 VDD.n244 0.0200283
R3413 VDD.n987 VDD.n834 0.0198458
R3414 VDD.n1856 VDD.n485 0.0197857
R3415 VDD.n1417 VDD.n1416 0.0197857
R3416 VDD.n2035 VDD.n2034 0.0194974
R3417 VDD.n308 VDD.n307 0.019371
R3418 VDD.n1150 VDD.n1149 0.0191328
R3419 VDD.n938 VDD.n937 0.0191207
R3420 VDD.n943 VDD.n942 0.019083
R3421 VDD.n1129 VDD.n1079 0.0190047
R3422 VDD.n1422 VDD.n746 0.0187022
R3423 VDD.n1221 VDD.n1181 0.0186452
R3424 VDD.n1216 VDD.n1186 0.0186452
R3425 VDD.n181 VDD.n177 0.0186395
R3426 VDD.n253 VDD.n235 0.0180472
R3427 VDD.n1838 VDD.n1837 0.017691
R3428 VDD.n1399 VDD.n1398 0.0176429
R3429 VDD.n271 VDD.n259 0.0174811
R3430 VDD.n2089 VDD.n2088 0.0173293
R3431 VDD.n985 VDD.n835 0.0173224
R3432 VDD.n977 VDD.n976 0.0173224
R3433 VDD.n415 VDD.n414 0.0167799
R3434 VDD.n2016 VDD.n2015 0.0167254
R3435 VDD.n1688 VDD.n1687 0.0165976
R3436 VDD.n1216 VDD.n1215 0.0164677
R3437 VDD.n1078 VDD.n994 0.0160453
R3438 VDD.n1007 VDD.n1006 0.0159438
R3439 VDD.n1006 VDD.n1003 0.0159438
R3440 VDD.n1077 VDD.n995 0.0159438
R3441 VDD.n2106 VDD 0.0158659
R3442 VDD.n1236 VDD.n826 0.0157992
R3443 VDD.n900 VDD.n873 0.0156402
R3444 VDD.n1127 VDD.n1126 0.0156402
R3445 VDD.n1230 VDD.n1229 0.015009
R3446 VDD.n936 VDD.n918 0.0149
R3447 VDD VDD.n230 0.0147661
R3448 VDD.n2022 VDD.n349 0.0146297
R3449 VDD.n935 VDD.n919 0.014
R3450 VDD.n2018 VDD.n2017 0.0136831
R3451 VDD.n1678 VDD.n1677 0.0136707
R3452 VDD.n1680 VDD.n1679 0.0136707
R3453 VDD.n691 VDD.n690 0.0136707
R3454 VDD.n1612 VDD.n1611 0.0136707
R3455 VDD.n1221 VDD.n1165 0.0135645
R3456 VDD.n58 VDD.n57 0.0134677
R3457 VDD.n2037 VDD.n2036 0.0130858
R3458 VDD.n1010 VDD.n1009 0.0130481
R3459 VDD.n1005 VDD.n1002 0.0130481
R3460 VDD.n1005 VDD.n1004 0.0130481
R3461 VDD.n2012 VDD.n2011 0.0122692
R3462 VDD.n829 VDD.n827 0.0122391
R3463 VDD.n398 VDD.n375 0.0121724
R3464 VDD.n844 VDD.n843 0.0121599
R3465 VDD.n1228 VDD.n1164 0.0121129
R3466 VDD.n1229 VDD.n1163 0.0119706
R3467 VDD.n930 VDD.n925 0.0118445
R3468 VDD.n567 VDD.n565 0.01175
R3469 VDD.n1976 VDD.n1975 0.0116236
R3470 VDD.n900 VDD.n871 0.0114346
R3471 VDD.n2034 VDD.n2033 0.0114235
R3472 VDD.n1792 VDD.n552 0.0112143
R3473 VDD.n390 VDD.n389 0.0109437
R3474 VDD.n1517 VDD.n1516 0.0107273
R3475 VDD.n1308 VDD.n785 0.0106124
R3476 VDD.n1126 VDD.n1125 0.0105935
R3477 VDD.n59 VDD.n12 0.0105
R3478 VDD.n221 VDD.n220 0.0104739
R3479 VDD.n52 VDD.n51 0.0103544
R3480 VDD.n1479 VDD.n1454 0.0101429
R3481 VDD.n1008 VDD.n1001 0.0100858
R3482 VDD.n1071 VDD.n1000 0.00993548
R3483 VDD.n986 VDD.n985 0.00975234
R3484 VDD.n95 VDD.n94 0.00952375
R3485 VDD.n1635 VDD 0.00932353
R3486 VDD.n1145 VDD.n993 0.00928906
R3487 VDD.n1118 VDD.n1083 0.00928049
R3488 VDD.n1124 VDD.n1080 0.00928049
R3489 VDD.n977 VDD.n835 0.00891121
R3490 VDD.n847 VDD.n846 0.00888057
R3491 VDD.n1122 VDD.n1083 0.00854878
R3492 VDD.n1124 VDD.n1123 0.00854878
R3493 VDD.n1072 VDD.n999 0.00853674
R3494 VDD.n972 VDD.n971 0.00851619
R3495 VDD.n407 VDD.n406 0.00848635
R3496 VDD.n935 VDD.n930 0.00806303
R3497 VDD.n891 VDD.n870 0.00778745
R3498 VDD.n689 VDD.n688 0.00775806
R3499 VDD.n1614 VDD.n1613 0.00775806
R3500 VDD.n1233 VDD.n830 0.00754348
R3501 VDD.n904 VDD.n880 0.00742308
R3502 VDD.n959 VDD.n958 0.00742308
R3503 VDD.n843 VDD.n836 0.00742308
R3504 VDD.n1164 VDD.n828 0.00738437
R3505 VDD.n53 VDD.n49 0.00725
R3506 VDD.n53 VDD.n52 0.00725
R3507 VDD.n1035 VDD.n1034 0.00708537
R3508 VDD.n859 VDD.n857 0.0070587
R3509 VDD.n901 VDD.n874 0.0070587
R3510 VDD.n1261 VDD.n1260 0.00700602
R3511 VDD.n1951 VDD.n1950 0.00700602
R3512 VDD.n984 VDD.n983 0.00669433
R3513 VDD.n105 VDD.n104 0.00667414
R3514 VDD VDD.n2019 0.00664335
R3515 VDD.n1175 VDD.n1171 0.00661998
R3516 VDD.n845 VDD.n834 0.00638785
R3517 VDD.n961 VDD.n960 0.00632996
R3518 VDD.n953 VDD.n952 0.00632996
R3519 VDD.n951 VDD.n914 0.00632996
R3520 VDD.n860 VDD.n847 0.00632996
R3521 VDD VDD.n1670 0.00630645
R3522 VDD.n679 VDD 0.00630645
R3523 VDD VDD.n648 0.00630645
R3524 VDD VDD.n1109 0.00630645
R3525 VDD.n1208 VDD 0.00630645
R3526 VDD VDD.n619 0.00630645
R3527 VDD.n1012 VDD.n1001 0.00582544
R3528 VDD.n1220 VDD.n1182 0.00579412
R3529 VDD.n845 VDD.n832 0.00572908
R3530 VDD.n2058 VDD.n2057 0.00562658
R3531 VDD.n1123 VDD.n1122 0.00562195
R3532 VDD.n1230 VDD.n830 0.00558696
R3533 VDD.n255 VDD.n254 0.00531132
R3534 VDD.n1125 VDD.n1081 0.00489628
R3535 VDD.n901 VDD.n899 0.00487247
R3536 VDD.n1234 VDD.n1233 0.00480435
R3537 VDD.n899 VDD.n898 0.0045081
R3538 VDD.n972 VDD.n874 0.0045081
R3539 VDD.n947 VDD.n915 0.00441304
R3540 VDD.n944 VDD.n943 0.00414372
R3541 VDD.n978 VDD.n837 0.00414372
R3542 VDD.n1074 VDD.n998 0.00412903
R3543 VDD.n1227 VDD.n1165 0.00412903
R3544 VDD.n1184 VDD.n1162 0.00402941
R3545 VDD.n1219 VDD.n1183 0.00402941
R3546 VDD.n40 VDD.n39 0.003875
R3547 VDD.n226 VDD.n120 0.00380882
R3548 VDD.n953 VDD.n907 0.00377935
R3549 VDD.n942 VDD.n914 0.00377935
R3550 VDD.n861 VDD.n859 0.00377935
R3551 VDD.n1014 VDD.n998 0.00376613
R3552 VDD.n1797 VDD.n1796 0.00371429
R3553 VDD.n1475 VDD.n1474 0.00371429
R3554 VDD.n827 VDD.n826 0.00360796
R3555 VDD.n1013 VDD.n999 0.00350186
R3556 VDD.n898 VDD.n890 0.00341498
R3557 VDD VDD.n1056 0.00340323
R3558 VDD.n1186 VDD.n1181 0.00340323
R3559 VDD.n861 VDD.n860 0.00305061
R3560 VDD.n846 VDD.n844 0.00305061
R3561 VDD.n1074 VDD.n1073 0.00304032
R3562 VDD.n47 VDD.n41 0.00283766
R3563 VDD.n973 VDD.n873 0.00283401
R3564 VDD.n48 VDD.n40 0.00275
R3565 VDD.n1246 VDD.n1245 0.00266867
R3566 VDD.n1916 VDD.n1912 0.00266867
R3567 VDD.n936 VDD 0.00254545
R3568 VDD.n1170 VDD.n1164 0.00254545
R3569 VDD.n971 VDD.n970 0.00245652
R3570 VDD.n950 VDD.n912 0.00206522
R3571 VDD.n1884 VDD.n455 0.00192857
R3572 VDD.n30 VDD 0.00186364
R3573 VDD VDD.n101 0.00163924
R3574 VDD VDD.n174 0.00163924
R3575 VDD VDD.n304 0.00163924
R3576 VDD VDD.n403 0.00163924
R3577 VDD.n983 VDD.n837 0.00159312
R3578 VDD.n978 VDD.n870 0.00159312
R3579 VDD.n1509 VDD.n1507 0.00152273
R3580 VDD.n1712 VDD.n1711 0.00152273
R3581 VDD.n1237 VDD 0.00151695
R3582 VDD.n255 VDD 0.00134906
R3583 VDD.n2015 VDD.n417 0.00132534
R3584 VDD.n2126 VDD 0.00128947
R3585 VDD.n952 VDD.n951 0.00122874
R3586 VDD VDD.n341 0.00122581
R3587 VDD.n331 VDD 0.00122581
R3588 VDD.n1215 VDD.n1187 0.00122581
R3589 VDD.n1300 VDD.n1299 0.00121429
R3590 VDD VDD.n213 0.00119767
R3591 VDD VDD.n164 0.00119767
R3592 VDD.n1013 VDD.n1012 0.00103254
R3593 VDD.n1171 VDD.n1170 0.00101136
R3594 VDD.n2046 VDD 0.000887097
R3595 VDD.n1071 VDD.n1014 0.000862903
R3596 VDD.n1149 VDD 0.000851563
R3597 VDD.n373 VDD 0.000807167
R3598 VDD.n391 VDD 0.000807167
R3599 VDD.n97 VDD 0.000737467
R3600 VDD.n87 VDD 0.000693548
R3601 VDD.n59 VDD.n58 0.000693548
R3602 VDD.n120 VDD.n116 0.000665441
R3603 VSS.n4304 VSS.n4303 5.941e+06
R3604 VSS.n5684 VSS.n5681 5.941e+06
R3605 VSS.n5684 VSS.n5683 3.75375e+06
R3606 VSS.n5735 VSS.n5734 3.75375e+06
R3607 VSS.n4762 VSS.n4761 1.21542e+06
R3608 VSS.n4761 VSS.n4760 558796
R3609 VSS.n5926 VSS.t593 148432
R3610 VSS.t692 VSS.t18 44337.9
R3611 VSS.n5877 VSS.n4762 28016
R3612 VSS.n4494 VSS.n4493 16684.1
R3613 VSS.n4305 VSS.n4304 15212.8
R3614 VSS.n4494 VSS.t43 13601.5
R3615 VSS.n5876 VSS.n5736 10655.7
R3616 VSS.n5014 VSS.n5013 10552.3
R3617 VSS.n5926 VSS.n5925 9445.69
R3618 VSS.n5779 VSS.t112 8953.91
R3619 VSS.n5854 VSS.n5769 8778.74
R3620 VSS.n5779 VSS.t578 7394.69
R3621 VSS.n4760 VSS.n4759 7304.73
R3622 VSS.t732 VSS.n5845 7210.65
R3623 VSS.n5814 VSS.t633 6204.1
R3624 VSS.n5013 VSS.n5012 6119.25
R3625 VSS.n5736 VSS.n5735 5553.02
R3626 VSS.t424 VSS.n5857 4486.13
R3627 VSS.n6019 VSS.n6018 4143.89
R3628 VSS.t51 VSS.t713 3685.04
R3629 VSS.n5844 VSS.t142 3621.08
R3630 VSS.n4303 VSS.n4302 3301.18
R3631 VSS.n5735 VSS.n4764 3000.68
R3632 VSS.n5355 VSS.n5354 2891.56
R3633 VSS.t662 VSS.t58 2166.67
R3634 VSS.t54 VSS.t94 2166.67
R3635 VSS.t141 VSS.t143 2166.67
R3636 VSS.n4735 VSS.n4734 1890.45
R3637 VSS.t55 VSS.t587 1842.52
R3638 VSS.t587 VSS.t52 1842.52
R3639 VSS.t116 VSS.t57 1822.88
R3640 VSS.t221 VSS.t89 1805.06
R3641 VSS.t237 VSS.t90 1778.39
R3642 VSS.n5855 VSS.n5854 1752.01
R3643 VSS.n959 VSS.t116 1720.94
R3644 VSS.t39 VSS.t46 1717.16
R3645 VSS.t43 VSS.t41 1707.46
R3646 VSS.t633 VSS.t120 1707.46
R3647 VSS.t246 VSS.t501 1657.99
R3648 VSS.t229 VSS.t503 1649.75
R3649 VSS.n5815 VSS.t576 1629.85
R3650 VSS.n4248 VSS.t647 1557.29
R3651 VSS.n6072 VSS.n6071 1536.82
R3652 VSS.n4858 VSS.n4857 1514.17
R3653 VSS.t663 VSS.n5931 1469.82
R3654 VSS.n4572 VSS.t237 1404.92
R3655 VSS.n48 VSS.t221 1316.01
R3656 VSS.n4591 VSS.t229 1303.3
R3657 VSS.n4392 VSS.t258 1229.06
R3658 VSS.n4670 VSS.t255 1229.06
R3659 VSS.n4591 VSS.t181 1224.94
R3660 VSS.n5800 VSS.t23 1216.04
R3661 VSS.t90 VSS.t87 1209.3
R3662 VSS.t89 VSS.t91 1209.3
R3663 VSS.n5926 VSS.t661 1153.55
R3664 VSS.n5845 VSS.t53 1153.55
R3665 VSS.t503 VSS.t86 1121.83
R3666 VSS.t501 VSS.t88 1121.83
R3667 VSS.t659 VSS.t39 1086.57
R3668 VSS.t122 VSS.t659 1086.57
R3669 VSS.t120 VSS.t122 1086.57
R3670 VSS.t687 VSS.t689 1083.33
R3671 VSS.t689 VSS.t661 1083.33
R3672 VSS.t762 VSS.t759 1083.33
R3673 VSS.t759 VSS.t53 1083.33
R3674 VSS.t25 VSS.t28 1083.33
R3675 VSS.t142 VSS.t25 1083.33
R3676 VSS.n5760 VSS.t166 1074.31
R3677 VSS.n5768 VSS.t84 1061.73
R3678 VSS.t723 VSS.t611 1060.11
R3679 VSS.t112 VSS.t574 1047.76
R3680 VSS.n5762 VSS.t472 967.024
R3681 VSS.n860 VSS.n859 953.981
R3682 VSS.n424 VSS.n423 944.048
R3683 VSS.n1479 VSS.n1478 929.726
R3684 VSS.n5925 VSS.t51 921.26
R3685 VSS.n5925 VSS.t55 921.26
R3686 VSS.n5736 VSS.n4763 914.569
R3687 VSS.t196 VSS.t428 855.827
R3688 VSS.n5857 VSS.t8 797.606
R3689 VSS.t578 VSS.t0 781.737
R3690 VSS.n5916 VSS.t687 767.361
R3691 VSS.n5784 VSS.t762 767.361
R3692 VSS.t28 VSS.n5843 767.361
R3693 VSS.t718 VSS.n5877 756.434
R3694 VSS.n5876 VSS.t701 750.444
R3695 VSS.t748 VSS.t146 727.73
R3696 VSS.n5878 VSS.t135 658.784
R3697 VSS.t101 VSS.n5875 650.385
R3698 VSS.n114 VSS.t226 617.99
R3699 VSS.t155 VSS.t153 581.962
R3700 VSS.t533 VSS.t155 581.962
R3701 VSS.t434 VSS.t533 581.962
R3702 VSS.t446 VSS.t448 581.962
R3703 VSS.t448 VSS.t466 581.962
R3704 VSS.n4971 VSS.n4970 572.302
R3705 VSS.n939 VSS.t62 561.086
R3706 VSS.n5925 VSS 552.953
R3707 VSS.t733 VSS.t263 522.588
R3708 VSS.t735 VSS.t722 522.588
R3709 VSS.n5853 VSS.t685 515.361
R3710 VSS.n5858 VSS.t424 481.087
R3711 VSS.n5336 VSS.n5335 477.231
R3712 VSS.n4468 VSS.t434 421.495
R3713 VSS.t726 VSS.t613 419.226
R3714 VSS.n591 VSS.n590 407.524
R3715 VSS.t146 VSS.t60 399.077
R3716 VSS.t96 VSS.t665 399.077
R3717 VSS.t98 VSS.t729 399.077
R3718 VSS.t743 VSS.t732 399.077
R3719 VSS.t468 VSS.t420 390.616
R3720 VSS.t471 VSS.t417 390.616
R3721 VSS.t103 VSS.t705 390.616
R3722 VSS.t139 VSS.t702 390.616
R3723 VSS.t2 VSS.t416 390.344
R3724 VSS.t11 VSS.t696 390.154
R3725 VSS.t140 VSS.t699 388.692
R3726 VSS.n5905 VSS.t267 365.812
R3727 VSS.n5859 VSS.n5858 352.084
R3728 VSS.n5916 VSS.t662 315.973
R3729 VSS.n5784 VSS.t54 315.973
R3730 VSS.n5843 VSS.t141 315.973
R3731 VSS.n162 VSS.t426 297.88
R3732 VSS.n199 VSS.t160 288.988
R3733 VSS.n5856 VSS.t14 282.526
R3734 VSS.n5015 VSS.n5014 281.462
R3735 VSS.n5769 VSS.n5768 279.142
R3736 VSS.n4612 VSS.t187 266.759
R3737 VSS.n202 VSS.t162 253.421
R3738 VSS.t724 VSS.n5926 248.296
R3739 VSS.n165 VSS.t528 244.529
R3740 VSS.n5854 VSS.n5853 240.343
R3741 VSS.t590 VSS.t172 232.776
R3742 VSS.n5930 VSS.t594 231.668
R3743 VSS.t576 VSS.n5814 223.135
R3744 VSS.t60 VSS.n5779 200.844
R3745 VSS.n4636 VSS.t92 191.177
R3746 VSS.n5683 VSS.n5682 187.726
R3747 VSS.n149 VSS.t202 186.731
R3748 VSS.t746 VSS.t683 182.947
R3749 VSS.n4618 VSS.t93 182.286
R3750 VSS.n5851 VSS.t740 181.751
R3751 VSS.t21 VSS.n5903 179.668
R3752 VSS.n121 VSS.t437 164.501
R3753 VSS.n5780 VSS.t748 164.327
R3754 VSS.t96 VSS.t764 164.327
R3755 VSS.t665 VSS.t98 164.327
R3756 VSS.t729 VSS.t743 164.327
R3757 VSS.n4468 VSS.t446 160.468
R3758 VSS.n5858 VSS.n5855 160.02
R3759 VSS.n5852 VSS.t744 156.163
R3760 VSS.n410 VSS.t648 154.649
R3761 VSS.n1526 VSS.n1525 145.089
R3762 VSS.n5904 VSS.t596 141.845
R3763 VSS.n465 VSS.t496 137.732
R3764 VSS.t482 VSS.t485 134.906
R3765 VSS.n456 VSS.n455 132.9
R3766 VSS.n5734 VSS.n5733 130.788
R3767 VSS.n206 VSS.t572 128.934
R3768 VSS.n1201 VSS.n1200 127.87
R3769 VSS.n4697 VSS.t125 127.856
R3770 VSS.n5001 VSS.n5000 127.537
R3771 VSS.n189 VSS.t525 120.041
R3772 VSS.n568 VSS.n567 116.502
R3773 VSS.n4210 VSS.t653 115.596
R3774 VSS.n391 VSS.n390 109.445
R3775 VSS.t5 VSS.n5856 107.629
R3776 VSS.n5989 VSS.n5988 98.3336
R3777 VSS.n5855 VSS.t49 92.842
R3778 VSS.t615 VSS.t675 88.6679
R3779 VSS.n5685 VSS.n5684 82.9732
R3780 VSS.n4957 VSS.t73 81.8473
R3781 VSS.n5710 VSS.n5709 81.5669
R3782 VSS.n5845 VSS.n5844 80.7206
R3783 VSS.t744 VSS.t715 75.3316
R3784 VSS.t683 VSS.n5782 74.1359
R3785 VSS.n569 VSS.n568 71.3171
R3786 VSS.n4725 VSS.t133 70.1147
R3787 VSS.n804 VSS.t636 68.7194
R3788 VSS.n854 VSS.t644 68.7194
R3789 VSS.n1432 VSS.t630 68.7194
R3790 VSS.n1489 VSS.t30 68.7194
R3791 VSS.n4630 VSS.t500 66.69
R3792 VSS.n325 VSS.t646 64.2392
R3793 VSS.n4714 VSS.t131 61.866
R3794 VSS.n474 VSS.t488 60.4094
R3795 VSS.n4864 VSS.t622 57.9753
R3796 VSS.n4939 VSS.t756 57.9753
R3797 VSS.n4898 VSS.t75 57.9753
R3798 VSS.n4624 VSS.t502 57.798
R3799 VSS.n4645 VSS.t190 57.798
R3800 VSS.n6065 VSS.n6064 55.1928
R3801 VSS.n5520 VSS.t178 51.6521
R3802 VSS.n4835 VSS.t669 51.1548
R3803 VSS.n4948 VSS.t751 51.1548
R3804 VSS.n4907 VSS.t70 51.1548
R3805 VSS.n5434 VSS.t275 49.6265
R3806 VSS.n4249 VSS.n4248 49.1159
R3807 VSS.n4914 VSS.n4913 44.3342
R3808 VSS.t776 VSS.t775 44.058
R3809 VSS.n5356 VSS.n5355 43.5499
R3810 VSS.n1226 VSS.n1225 42.6234
R3811 VSS.n5052 VSS.t80 41.5243
R3812 VSS.n5150 VSS.t175 41.5243
R3813 VSS.n5910 VSS.t266 38.8649
R3814 VSS.n4835 VSS.t617 37.5136
R3815 VSS.n5496 VSS.t83 35.4477
R3816 VSS.n4103 VSS.n4102 32.9568
R3817 VSS.n4495 VSS.n4494 31.0858
R3818 VSS.n4864 VSS.t672 30.6931
R3819 VSS.n1295 VSS.n1294 29.9489
R3820 VSS.n3932 VSS.n3931 29.0184
R3821 VSS.n1285 VSS.t650 28.751
R3822 VSS.n1389 VSS.n1388 28.7316
R3823 VSS.t266 VSS.t776 28.6791
R3824 VSS.n5592 VSS.t148 28.3582
R3825 VSS.n4915 VSS.t749 27.2828
R3826 VSS.n5199 VSS.t457 26.3327
R3827 VSS.n4113 VSS.n4112 26.1965
R3828 VSS.n414 VSS.t651 26.1718
R3829 VSS.n495 VSS.n494 26.0884
R3830 VSS.n4102 VSS.t482 25.3911
R3831 VSS.n953 VSS.t480 25.3179
R3832 VSS.n480 VSS.t478 24.1641
R3833 VSS.n4915 VSS.n4914 23.8725
R3834 VSS.n4077 VSS.t107 21.9714
R3835 VSS.n5846 VSS.n5781 21.6
R3836 VSS.n4306 VSS.n4305 20.5962
R3837 VSS.n5863 VSS.n5862 19.7293
R3838 VSS.n913 VSS.t108 19.4363
R3839 VSS.n425 VSS.n424 19.0342
R3840 VSS.n5934 VSS.n5933 18.6126
R3841 VSS.n5413 VSS.t517 18.2305
R3842 VSS.t685 VSS.n5852 17.9365
R3843 VSS.n5592 VSS.n5591 17.2177
R3844 VSS.n4841 VSS.t615 17.0519
R3845 VSS.n5929 VSS.t173 16.2066
R3846 VSS.n4086 VSS.n4085 15.2111
R3847 VSS.n4109 VSS.t491 15.2111
R3848 VSS.n5457 VSS.t451 15.1921
R3849 VSS.t611 VSS.t692 14.9316
R3850 VSS.t596 VSS.t723 14.9316
R3851 VSS.n5905 VSS.n5904 14.9316
R3852 VSS.t267 VSS.t733 14.9316
R3853 VSS.t263 VSS.t735 14.9316
R3854 VSS.t722 VSS.t593 14.9316
R3855 VSS.n5025 VSS.t218 13.1666
R3856 VSS.n5046 VSS.t81 13.1666
R3857 VSS.n5451 VSS.t504 13.1666
R3858 VSS.n5863 VSS.n5757 12.9101
R3859 VSS.n6063 VSS.n6062 12.8022
R3860 VSS.t135 VSS.t718 11.9784
R3861 VSS.t613 VSS.t21 11.9784
R3862 VSS.t18 VSS.t726 11.9784
R3863 VSS.n5929 VSS.n5928 11.769
R3864 VSS.n1010 VSS.t40 11.3982
R3865 VSS.n3991 VSS.t34 11.0483
R3866 VSS.n5844 VSS.t746 10.9931
R3867 VSS.n1015 VSS.n1014 10.7852
R3868 VSS.n4051 VSS.t771 10.3984
R3869 VSS.n4188 VSS.t65 10.315
R3870 VSS.n5557 VSS.t442 10.1283
R3871 VSS.n4017 VSS.t32 9.74855
R3872 VSS.n5875 VSS.t475 9.62158
R3873 VSS.n508 VSS.n507 9.61182
R3874 VSS.n5077 VSS.t215 9.55913
R3875 VSS.n4511 VSS.t236 9.55885
R3876 VSS.n76 VSS.t272 9.54136
R3877 VSS.n5064 VSS.t250 9.54089
R3878 VSS.n5065 VSS.t177 9.51568
R3879 VSS.n94 VSS.t228 9.5154
R3880 VSS.n5063 VSS.t281 9.5085
R3881 VSS.n63 VSS.t186 9.50824
R3882 VSS.n4510 VSS.t248 9.49457
R3883 VSS.n33 VSS.t220 9.49428
R3884 VSS.n32 VSS.t239 9.49428
R3885 VSS.n31 VSS.t254 9.49428
R3886 VSS.n58 VSS.t245 9.49428
R3887 VSS.n4965 VSS.t269 9.49403
R3888 VSS.n4964 VSS.t277 9.49403
R3889 VSS.n4925 VSS.t233 9.49403
R3890 VSS.n4807 VSS.t217 9.49403
R3891 VSS.n5066 VSS.t223 9.49372
R3892 VSS.n59 VSS.t189 9.45083
R3893 VSS.n4806 VSS.t279 9.45057
R3894 VSS.n92 VSS.t243 9.43205
R3895 VSS.n4508 VSS.t180 9.43205
R3896 VSS.n82 VSS.t206 9.43205
R3897 VSS.n74 VSS.t260 9.43205
R3898 VSS.n65 VSS.t201 9.43205
R3899 VSS.n5075 VSS.t204 9.43205
R3900 VSS.n5110 VSS.t252 9.43205
R3901 VSS.n5131 VSS.t231 9.43205
R3902 VSS.n5103 VSS.t241 9.43205
R3903 VSS.n5122 VSS.t174 9.43205
R3904 VSS.n4378 VSS.t198 9.3886
R3905 VSS.n5298 VSS.t213 9.3886
R3906 VSS.n5322 VSS.t274 9.3886
R3907 VSS.n4409 VSS.t195 9.3886
R3908 VSS.n243 VSS.t225 9.34514
R3909 VSS.n4382 VSS.t257 9.34514
R3910 VSS.n108 VSS.t192 9.34514
R3911 VSS.n5253 VSS.t211 9.34514
R3912 VSS.n5274 VSS.t183 9.34514
R3913 VSS.n5258 VSS.t208 9.34514
R3914 VSS.n1460 VSS.n1458 9.13939
R3915 VSS.n4717 VSS.n4715 9.13939
R3916 VSS.n4719 VSS.n4717 9.13939
R3917 VSS.n4712 VSS.n4711 9.13939
R3918 VSS.n4711 VSS.n4710 9.13939
R3919 VSS.n839 VSS.n837 9.13939
R3920 VSS.n4947 VSS.n4930 9.13939
R3921 VSS.n4949 VSS.n4947 9.13939
R3922 VSS.n4834 VSS.n4818 9.13939
R3923 VSS.n4836 VSS.n4834 9.13939
R3924 VSS.n4872 VSS.n4855 9.13939
R3925 VSS.n4874 VSS.n4872 9.13939
R3926 VSS.n4906 VSS.n4812 9.13939
R3927 VSS.n4908 VSS.n4906 9.13939
R3928 VSS.n5025 VSS.n5024 9.11549
R3929 VSS.n6096 VSS.t635 8.89703
R3930 VSS.n26 VSS.n25 8.78137
R3931 VSS.n27 VSS.t145 8.5505
R3932 VSS.n28 VSS.t121 8.5505
R3933 VSS.n6096 VSS.t634 8.5505
R3934 VSS.n1010 VSS.n1009 8.5505
R3935 VSS.t255 VSS.t246 8.24923
R3936 VSS.n4157 VSS.n4155 8.16717
R3937 VSS.n1078 VSS.n1077 7.61323
R3938 VSS.n1468 VSS.n1466 7.58383
R3939 VSS.n957 VSS.n956 7.50194
R3940 VSS.n830 VSS.n828 7.48661
R3941 VSS.n5910 VSS.t262 7.3005
R3942 VSS.n5502 VSS.t82 7.08994
R3943 VSS.n5866 VSS.n5742 6.8902
R3944 VSS.n5867 VSS.n5741 6.87063
R3945 VSS.n5862 VSS.t425 6.80709
R3946 VSS.n1382 VSS.n1381 6.76077
R3947 VSS.n5757 VSS.t473 6.68867
R3948 VSS.n924 VSS.n923 6.65541
R3949 VSS.n948 VSS.t117 6.65541
R3950 VSS.n1425 VSS.n1418 6.65541
R3951 VSS.n1425 VSS.n1419 6.65541
R3952 VSS.n1482 VSS.t629 6.65541
R3953 VSS.n1482 VSS.t31 6.65541
R3954 VSS.n1405 VSS.t35 6.65541
R3955 VSS.n3981 VSS.n1524 6.65541
R3956 VSS.n797 VSS.n790 6.65541
R3957 VSS.n797 VSS.n791 6.65541
R3958 VSS.n863 VSS.t645 6.65541
R3959 VSS.n863 VSS.t682 6.65541
R3960 VSS.n4885 VSS.t616 6.65541
R3961 VSS.n4860 VSS.n4856 6.65541
R3962 VSS.n4822 VSS.n4819 6.65541
R3963 VSS.n4847 VSS.t676 6.65541
R3964 VSS.n4894 VSS.n4813 6.65541
R3965 VSS.n4921 VSS.t74 6.65541
R3966 VSS.n4960 VSS.t750 6.65541
R3967 VSS.n4935 VSS.n4931 6.65541
R3968 VSS.n4198 VSS.t481 6.65541
R3969 VSS.n4138 VSS.n890 6.65541
R3970 VSS.n4692 VSS.n29 6.65541
R3971 VSS.n4692 VSS.n30 6.65541
R3972 VSS.n4733 VSS.t134 6.65541
R3973 VSS.n4733 VSS.t581 6.65541
R3974 VSS.t594 VSS.t724 6.65125
R3975 VSS.t172 VSS.t663 6.65125
R3976 VSS.n4509 VSS.t182 6.63905
R3977 VSS.n5076 VSS.t205 6.63905
R3978 VSS.n4379 VSS.t200 6.63522
R3979 VSS.n5323 VSS.t276 6.63522
R3980 VSS.n5299 VSS.t214 6.63522
R3981 VSS.n4410 VSS.t197 6.63522
R3982 VSS.n4383 VSS.t259 6.63331
R3983 VSS.n5275 VSS.t185 6.63331
R3984 VSS.n5746 VSS.t12 6.62607
R3985 VSS.n5754 VSS.t15 6.62607
R3986 VSS.n5747 VSS.n5743 6.6202
R3987 VSS.n5755 VSS.n5751 6.6202
R3988 VSS.n244 VSS.t227 6.5165
R3989 VSS.n5254 VSS.t212 6.5165
R3990 VSS.n109 VSS.t194 6.50525
R3991 VSS.n5259 VSS.t210 6.50525
R3992 VSS.n5749 VSS.n5748 6.4265
R3993 VSS.n5756 VSS.n5750 6.4265
R3994 VSS.n148 VSS.t427 6.4265
R3995 VSS.n146 VSS.t597 6.4265
R3996 VSS.n141 VSS.t538 6.4265
R3997 VSS.n84 VSS.t244 6.4265
R3998 VSS.n77 VSS.t207 6.4265
R3999 VSS.n64 VSS.t261 6.4265
R4000 VSS.n66 VSS.t203 6.4265
R4001 VSS.n4357 VSS.n4356 6.4265
R4002 VSS.n105 VSS.n104 6.4265
R4003 VSS.n103 VSS.n102 6.4265
R4004 VSS.n5121 VSS.t232 6.4265
R4005 VSS.n5168 VSS.n5163 6.4265
R4006 VSS.n5098 VSS.n5097 6.4265
R4007 VSS.n5319 VSS.t165 6.4265
R4008 VSS.n5250 VSS.t431 6.4265
R4009 VSS.n5255 VSS.t520 6.4265
R4010 VSS.n5096 VSS.t242 6.4265
R4011 VSS.n5105 VSS.t253 6.4265
R4012 VSS.n5170 VSS.n5162 6.4265
R4013 VSS.n5123 VSS.t176 6.4265
R4014 VSS.n3738 VSS.n3737 6.39416
R4015 VSS.n4123 VSS.n4122 5.91574
R4016 VSS.n1176 VSS.n1175 5.84933
R4017 VSS.n259 VSS.n258 5.80511
R4018 VSS.n5839 VSS.n5838 5.60567
R4019 VSS.n528 VSS.n527 5.60395
R4020 VSS.n5932 VSS.t169 5.54279
R4021 VSS.n1028 VSS.n1027 5.4005
R4022 VSS.n1028 VSS.t42 5.4005
R4023 VSS.n24 VSS.n23 5.4005
R4024 VSS.n24 VSS.t660 5.4005
R4025 VSS.n5899 VSS.t136 5.35216
R4026 VSS VSS.t686 5.34447
R4027 VSS VSS.t664 5.34447
R4028 VSS VSS.t745 5.34447
R4029 VSS VSS.n5910 5.27587
R4030 VSS.n5920 VSS.n5919 5.27322
R4031 VSS.n5788 VSS.n5787 5.27322
R4032 VSS.n5922 VSS.n5921 5.27266
R4033 VSS.n270 VSS.n269 5.26318
R4034 VSS.n6098 VSS.n6097 5.24323
R4035 VSS.n5915 VSS.t59 5.23126
R4036 VSS.n4749 VSS.t714 5.23126
R4037 VSS.n4750 VSS.t612 5.23126
R4038 VSS.n5887 VSS.t693 5.23126
R4039 VSS.n5783 VSS.t95 5.23126
R4040 VSS.n5839 VSS.t144 5.23126
R4041 VSS.n5789 VSS.t147 5.23126
R4042 VSS.n5792 VSS.t61 5.23126
R4043 VSS.n1012 VSS.n1011 5.20095
R4044 VSS VSS.n5916 5.2005
R4045 VSS.n952 VSS.n951 5.2005
R4046 VSS.n954 VSS.n953 5.2005
R4047 VSS.n3998 VSS.n3997 5.2005
R4048 VSS.n4022 VSS.n4021 5.2005
R4049 VSS.n4016 VSS.n4015 5.2005
R4050 VSS.n4015 VSS.n4014 5.2005
R4051 VSS.n1516 VSS.n1515 5.2005
R4052 VSS.n286 VSS.n285 5.2005
R4053 VSS.n285 VSS.n284 5.2005
R4054 VSS.n289 VSS.n288 5.2005
R4055 VSS.n288 VSS.n287 5.2005
R4056 VSS.n293 VSS.n291 5.2005
R4057 VSS.n293 VSS.n292 5.2005
R4058 VSS.n278 VSS.n277 5.2005
R4059 VSS.n466 VSS.n465 5.2005
R4060 VSS.n830 VSS.n820 5.2005
R4061 VSS.n830 VSS.n829 5.2005
R4062 VSS.n359 VSS.n338 5.2005
R4063 VSS.n330 VSS.n329 5.2005
R4064 VSS.n329 VSS.n328 5.2005
R4065 VSS.n333 VSS.n332 5.2005
R4066 VSS.n332 VSS.n331 5.2005
R4067 VSS.n341 VSS.n340 5.2005
R4068 VSS.n4134 VSS.n4133 5.2005
R4069 VSS.n4192 VSS.n4191 5.2005
R4070 VSS.n4157 VSS.n4156 5.2005
R4071 VSS.n4178 VSS.n4177 5.2005
R4072 VSS.n4218 VSS.n4217 5.2005
R4073 VSS.n4217 VSS.n4216 5.2005
R4074 VSS.n4215 VSS.n4214 5.2005
R4075 VSS.n4214 VSS.n4213 5.2005
R4076 VSS.n4687 VSS.n4686 5.2005
R4077 VSS VSS.n5932 5.2005
R4078 VSS.n5930 VSS 5.2005
R4079 VSS VSS.n5905 5.2005
R4080 VSS VSS.n5904 5.2005
R4081 VSS.n5879 VSS.n5878 5.2005
R4082 VSS.n5903 VSS.n5902 5.2005
R4083 VSS.n5875 VSS 5.2005
R4084 VSS VSS.n5784 5.2005
R4085 VSS.n5843 VSS 5.2005
R4086 VSS.n1466 VSS.n1465 5.2005
R4087 VSS.n1395 VSS.n1394 5.2005
R4088 VSS.n4122 VSS.n4121 5.2005
R4089 VSS.n4120 VSS.n917 5.2005
R4090 VSS.n1397 VSS.n1396 5.2005
R4091 VSS.n914 VSS.n913 5.2005
R4092 VSS.n4129 VSS.n4128 5.2005
R4093 VSS.n4132 VSS.n4131 5.2005
R4094 VSS.n916 VSS.n915 5.2005
R4095 VSS.n960 VSS.n959 5.2005
R4096 VSS.n964 VSS.n963 5.2005
R4097 VSS.n4203 VSS.n4202 5.2005
R4098 VSS.n4205 VSS.n4204 5.2005
R4099 VSS.n4207 VSS.n4206 5.2005
R4100 VSS.n5851 VSS 5.2005
R4101 VSS.n5782 VSS 5.2005
R4102 VSS.n5801 VSS.n5800 5.2005
R4103 VSS.n5818 VSS.n5815 5.2005
R4104 VSS.n1030 VSS.n1026 5.2005
R4105 VSS.n999 VSS.n0 5.2005
R4106 VSS VSS.n1 5.2005
R4107 VSS.n6106 VSS.n2 5.2005
R4108 VSS.n6105 VSS.n18 5.2005
R4109 VSS.n6104 VSS.n19 5.2005
R4110 VSS.n6102 VSS.n22 5.2005
R4111 VSS.n6100 VSS.n6094 5.2005
R4112 VSS.n6099 VSS.n6095 5.2005
R4113 VSS.n1024 VSS.n1023 5.2005
R4114 VSS.n1031 VSS.n1025 5.2005
R4115 VSS.n144 VSS.t506 5.1234
R4116 VSS.n4503 VSS.t467 5.12337
R4117 VSS.n5545 VSS.n5544 5.12337
R4118 VSS.n4406 VSS.n4395 5.12334
R4119 VSS.n5318 VSS.t149 5.12332
R4120 VSS.n5166 VSS.n5164 5.12328
R4121 VSS.n5282 VSS.t559 5.12118
R4122 VSS.n4360 VSS.n4359 5.12105
R4123 VSS.n4756 VSS.t719 5.06496
R4124 VSS.n5820 VSS.t24 5.06496
R4125 VSS.n5812 VSS.t577 5.06496
R4126 VSS.n4088 VSS.n1393 4.88533
R4127 VSS.n327 VSS.n324 4.88449
R4128 VSS.n283 VSS.n280 4.88277
R4129 VSS.n4212 VSS.n4209 4.88215
R4130 VSS.n4177 VSS.t493 4.6889
R4131 VSS.n2795 VSS.n2794 4.50764
R4132 VSS.n2662 VSS.n2661 4.50764
R4133 VSS.n2791 VSS.n2790 4.50622
R4134 VSS.n2724 VSS.n2723 4.50622
R4135 VSS.n2562 VSS.n2561 4.50565
R4136 VSS.n2658 VSS.n2657 4.50564
R4137 VSS.n2197 VSS.n2195 4.50554
R4138 VSS.n2881 VSS.n2880 4.50542
R4139 VSS.n2582 VSS.n2581 4.50495
R4140 VSS.n2493 VSS.n2492 4.5026
R4141 VSS.n2492 VSS.n2491 4.50224
R4142 VSS.n2882 VSS.n2881 4.50095
R4143 VSS.n2794 VSS.n2793 4.50095
R4144 VSS.n2792 VSS.n2791 4.50095
R4145 VSS.n2726 VSS.n2197 4.50095
R4146 VSS.n2725 VSS.n2724 4.50095
R4147 VSS.n2661 VSS.n2660 4.50095
R4148 VSS.n2563 VSS.n2562 4.50089
R4149 VSS.n2659 VSS.n2658 4.50089
R4150 VSS.n2582 VSS.n2564 4.50089
R4151 VSS.n4011 VSS.n4008 4.5005
R4152 VSS.n4011 VSS.n4010 4.5005
R4153 VSS.n4001 VSS.n4000 4.5005
R4154 VSS.n1519 VSS.n1518 4.5005
R4155 VSS.n296 VSS.n295 4.5005
R4156 VSS.n295 VSS.n294 4.5005
R4157 VSS.n468 VSS.n467 4.5005
R4158 VSS.n283 VSS.n282 4.5005
R4159 VSS.n282 VSS.n281 4.5005
R4160 VSS.n833 VSS.n826 4.5005
R4161 VSS.n833 VSS.n832 4.5005
R4162 VSS.n262 VSS.n261 4.5005
R4163 VSS.n261 VSS.n260 4.5005
R4164 VSS.n327 VSS.n326 4.5005
R4165 VSS.n326 VSS.n325 4.5005
R4166 VSS.n346 VSS.n345 4.5005
R4167 VSS.n345 VSS.n344 4.5005
R4168 VSS.n2001 VSS.n1996 4.5005
R4169 VSS.n2018 VSS.n2004 4.5005
R4170 VSS.n2015 VSS.n2014 4.5005
R4171 VSS.n2019 VSS.n2005 4.5005
R4172 VSS.n2070 VSS.n2069 4.5005
R4173 VSS.n2083 VSS.n2082 4.5005
R4174 VSS.n2842 VSS.n2841 4.5005
R4175 VSS.n2025 VSS.n2023 4.5005
R4176 VSS.n2804 VSS.n2803 4.5005
R4177 VSS.n2817 VSS.n2816 4.5005
R4178 VSS.n2829 VSS.n2828 4.5005
R4179 VSS.n2878 VSS.n2877 4.5005
R4180 VSS.n2815 VSS.n2814 4.5005
R4181 VSS.n2827 VSS.n2826 4.5005
R4182 VSS.n2068 VSS.n2067 4.5005
R4183 VSS.n2031 VSS.n2016 4.5005
R4184 VSS.n2858 VSS.n2857 4.5005
R4185 VSS.n2039 VSS.n2038 4.5005
R4186 VSS.n2876 VSS.n2875 4.5005
R4187 VSS.n2867 VSS.n2866 4.5005
R4188 VSS.n2037 VSS.n2027 4.5005
R4189 VSS.n2840 VSS.n2839 4.5005
R4190 VSS.n2831 VSS.n2830 4.5005
R4191 VSS.n2081 VSS.n2078 4.5005
R4192 VSS.n2046 VSS.n2045 4.5005
R4193 VSS.n2041 VSS.n2040 4.5005
R4194 VSS.n2000 VSS.n1997 4.5005
R4195 VSS.n2088 VSS.n2085 4.5005
R4196 VSS.n2806 VSS.n2805 4.5005
R4197 VSS.n2825 VSS.n2824 4.5005
R4198 VSS.n2012 VSS.n2008 4.5005
R4199 VSS.n2813 VSS.n2812 4.5005
R4200 VSS.n2846 VSS.n2845 4.5005
R4201 VSS.n2036 VSS.n2035 4.5005
R4202 VSS.n2860 VSS.n2859 4.5005
R4203 VSS.n2065 VSS.n2063 4.5005
R4204 VSS.n2071 VSS.n2066 4.5005
R4205 VSS.n2869 VSS.n2868 4.5005
R4206 VSS.n2187 VSS.n2178 4.5005
R4207 VSS.n2732 VSS.n2175 4.5005
R4208 VSS.n2133 VSS.n2132 4.5005
R4209 VSS.n2138 VSS.n2117 4.5005
R4210 VSS.n2106 VSS.n2103 4.5005
R4211 VSS.n2136 VSS.n2135 4.5005
R4212 VSS.n2107 VSS.n2105 4.5005
R4213 VSS.n2139 VSS.n2118 4.5005
R4214 VSS.n2176 VSS.n2174 4.5005
R4215 VSS.n2184 VSS.n2165 4.5005
R4216 VSS.n2186 VSS.n2185 4.5005
R4217 VSS.n2731 VSS.n2730 4.5005
R4218 VSS.n2101 VSS.n2095 4.5005
R4219 VSS.n2788 VSS.n2787 4.5005
R4220 VSS.n2734 VSS.n2733 4.5005
R4221 VSS.n2164 VSS.n2129 4.5005
R4222 VSS.n2099 VSS.n2096 4.5005
R4223 VSS.n2776 VSS.n2775 4.5005
R4224 VSS.n2745 VSS.n2744 4.5005
R4225 VSS.n2145 VSS.n2128 4.5005
R4226 VSS.n2196 VSS.n2194 4.5005
R4227 VSS.n2778 VSS.n2777 4.5005
R4228 VSS.n2113 VSS.n2109 4.5005
R4229 VSS.n2758 VSS.n2757 4.5005
R4230 VSS.n2183 VSS.n2182 4.5005
R4231 VSS.n2200 VSS.n2199 4.5005
R4232 VSS.n2147 VSS.n2144 4.5005
R4233 VSS.n2124 VSS.n2120 4.5005
R4234 VSS.n2736 VSS.n2735 4.5005
R4235 VSS.n2786 VSS.n2785 4.5005
R4236 VSS.n2134 VSS.n2114 4.5005
R4237 VSS.n2181 VSS.n2180 4.5005
R4238 VSS.n2767 VSS.n2766 4.5005
R4239 VSS.n2747 VSS.n2746 4.5005
R4240 VSS.n2202 VSS.n2201 4.5005
R4241 VSS.n2765 VSS.n2764 4.5005
R4242 VSS.n2721 VSS.n2720 4.5005
R4243 VSS.n2702 VSS.n2701 4.5005
R4244 VSS.n2282 VSS.n2278 4.5005
R4245 VSS.n2218 VSS.n2213 4.5005
R4246 VSS.n2246 VSS.n2237 4.5005
R4247 VSS.n2233 VSS.n2229 4.5005
R4248 VSS.n2291 VSS.n2290 4.5005
R4249 VSS.n2305 VSS.n2304 4.5005
R4250 VSS.n2302 VSS.n2270 4.5005
R4251 VSS.n2283 VSS.n2280 4.5005
R4252 VSS.n2700 VSS.n2699 4.5005
R4253 VSS.n2301 VSS.n2269 4.5005
R4254 VSS.n2300 VSS.n2299 4.5005
R4255 VSS.n2285 VSS.n2248 4.5005
R4256 VSS.n2231 VSS.n2221 4.5005
R4257 VSS.n2287 VSS.n2286 4.5005
R4258 VSS.n2665 VSS.n2664 4.5005
R4259 VSS.n2232 VSS.n2222 4.5005
R4260 VSS.n2710 VSS.n2709 4.5005
R4261 VSS.n2239 VSS.n2236 4.5005
R4262 VSS.n2313 VSS.n2281 4.5005
R4263 VSS.n2303 VSS.n2272 4.5005
R4264 VSS.n2217 VSS.n2214 4.5005
R4265 VSS.n2712 VSS.n2711 4.5005
R4266 VSS.n2677 VSS.n2676 4.5005
R4267 VSS.n2289 VSS.n2251 4.5005
R4268 VSS.n2298 VSS.n2254 4.5005
R4269 VSS.n2669 VSS.n2668 4.5005
R4270 VSS.n2690 VSS.n2689 4.5005
R4271 VSS.n2667 VSS.n2666 4.5005
R4272 VSS.n2228 VSS.n2224 4.5005
R4273 VSS.n2698 VSS.n2697 4.5005
R4274 VSS.n2288 VSS.n2249 4.5005
R4275 VSS.n2679 VSS.n2678 4.5005
R4276 VSS.n2244 VSS.n2238 4.5005
R4277 VSS.n2719 VSS.n2718 4.5005
R4278 VSS.n2655 VSS.n2654 4.5005
R4279 VSS.n2345 VSS.n2344 4.5005
R4280 VSS.n2631 VSS.n2630 4.5005
R4281 VSS.n2343 VSS.n2333 4.5005
R4282 VSS.n2391 VSS.n2390 4.5005
R4283 VSS.n2591 VSS.n2590 4.5005
R4284 VSS.n2566 VSS.n2404 4.5005
R4285 VSS.n2328 VSS.n2321 4.5005
R4286 VSS.n2643 VSS.n2642 4.5005
R4287 VSS.n2629 VSS.n2628 4.5005
R4288 VSS.n2403 VSS.n2401 4.5005
R4289 VSS.n2606 VSS.n2605 4.5005
R4290 VSS.n2622 VSS.n2621 4.5005
R4291 VSS.n2350 VSS.n2348 4.5005
R4292 VSS.n2604 VSS.n2603 4.5005
R4293 VSS.n2593 VSS.n2592 4.5005
R4294 VSS.n2618 VSS.n2363 4.5005
R4295 VSS.n2389 VSS.n2388 4.5005
R4296 VSS.n2620 VSS.n2619 4.5005
R4297 VSS.n2641 VSS.n2330 4.5005
R4298 VSS.n2645 VSS.n2644 4.5005
R4299 VSS.n2342 VSS.n2340 4.5005
R4300 VSS.n2347 VSS.n2341 4.5005
R4301 VSS.n2339 VSS.n2335 4.5005
R4302 VSS.n2386 VSS.n2384 4.5005
R4303 VSS.n2589 VSS.n2588 4.5005
R4304 VSS.n2565 VSS.n2405 4.5005
R4305 VSS.n2355 VSS.n2349 4.5005
R4306 VSS.n2608 VSS.n2607 4.5005
R4307 VSS.n2595 VSS.n2594 4.5005
R4308 VSS.n2334 VSS.n2327 4.5005
R4309 VSS.n2324 VSS.n2322 4.5005
R4310 VSS.n2406 VSS.n2402 4.5005
R4311 VSS.n2392 VSS.n2387 4.5005
R4312 VSS.n2617 VSS.n2616 4.5005
R4313 VSS.n2627 VSS.n2626 4.5005
R4314 VSS.n2602 VSS.n2601 4.5005
R4315 VSS.n2653 VSS.n2652 4.5005
R4316 VSS.n2529 VSS.n2528 4.5005
R4317 VSS.n2518 VSS.n2517 4.5005
R4318 VSS.n2428 VSS.n2427 4.5005
R4319 VSS.n2532 VSS.n2531 4.5005
R4320 VSS.n2520 VSS.n2519 4.5005
R4321 VSS.n2472 VSS.n2453 4.5005
R4322 VSS.n2489 VSS.n2481 4.5005
R4323 VSS.n2437 VSS.n2430 4.5005
R4324 VSS.n2557 VSS.n2414 4.5005
R4325 VSS.n2450 VSS.n2442 4.5005
R4326 VSS.n2506 VSS.n2505 4.5005
R4327 VSS.n2494 VSS.n2493 4.5005
R4328 VSS.n2559 VSS.n2558 4.5005
R4329 VSS.n2504 VSS.n2503 4.5005
R4330 VSS.n2417 VSS.n2415 4.5005
R4331 VSS.n2424 VSS.n2422 4.5005
R4332 VSS.n2508 VSS.n2507 4.5005
R4333 VSS.n2534 VSS.n2533 4.5005
R4334 VSS.n2476 VSS.n2473 4.5005
R4335 VSS.n2443 VSS.n2441 4.5005
R4336 VSS.n2452 VSS.n2448 4.5005
R4337 VSS.n2556 VSS.n2555 4.5005
R4338 VSS.n2470 VSS.n2454 4.5005
R4339 VSS.n2496 VSS.n2495 4.5005
R4340 VSS.n2449 VSS.n2444 4.5005
R4341 VSS.n2435 VSS.n2431 4.5005
R4342 VSS.n2490 VSS.n2482 4.5005
R4343 VSS.n2516 VSS.n2515 4.5005
R4344 VSS.n2420 VSS.n2419 4.5005
R4345 VSS.n2457 VSS.n2455 4.5005
R4346 VSS.n2536 VSS.n2535 4.5005
R4347 VSS.n2524 VSS.n2523 4.5005
R4348 VSS.n2537 VSS.n2432 4.5005
R4349 VSS.n2511 VSS.n2456 4.5005
R4350 VSS.n2480 VSS.n2478 4.5005
R4351 VSS.n2554 VSS.n2553 4.5005
R4352 VSS.n2510 VSS.n2509 4.5005
R4353 VSS.n2514 VSS.n2513 4.5005
R4354 VSS.n2446 VSS.n2445 4.5005
R4355 VSS.n2471 VSS.n2469 4.5005
R4356 VSS.n2551 VSS.n2550 4.5005
R4357 VSS.n2358 VSS.n2351 4.5005
R4358 VSS.n2615 VSS.n2614 4.5005
R4359 VSS.n2585 VSS.n2408 4.5005
R4360 VSS.n2409 VSS.n2407 4.5005
R4361 VSS.n2396 VSS.n2385 4.5005
R4362 VSS.n2647 VSS.n2646 4.5005
R4363 VSS.n2354 VSS.n2353 4.5005
R4364 VSS.n2636 VSS.n2337 4.5005
R4365 VSS.n2397 VSS.n2393 4.5005
R4366 VSS.n2587 VSS.n2586 4.5005
R4367 VSS.n2611 VSS.n2610 4.5005
R4368 VSS.n2370 VSS.n2369 4.5005
R4369 VSS.n2371 VSS.n2365 4.5005
R4370 VSS.n2336 VSS.n2326 4.5005
R4371 VSS.n2649 VSS.n2323 4.5005
R4372 VSS.n2400 VSS.n2398 4.5005
R4373 VSS.n2609 VSS.n2383 4.5005
R4374 VSS.n2357 VSS.n2356 4.5005
R4375 VSS.n2635 VSS.n2634 4.5005
R4376 VSS.n2651 VSS.n2650 4.5005
R4377 VSS.n2311 VSS.n2276 4.5005
R4378 VSS.n2245 VSS.n2243 4.5005
R4379 VSS.n2681 VSS.n2680 4.5005
R4380 VSS.n2717 VSS.n2716 4.5005
R4381 VSS.n2242 VSS.n2240 4.5005
R4382 VSS.n2315 VSS.n2314 4.5005
R4383 VSS.n2675 VSS.n2674 4.5005
R4384 VSS.n2688 VSS.n2687 4.5005
R4385 VSS.n2268 VSS.n2267 4.5005
R4386 VSS.n2708 VSS.n2707 4.5005
R4387 VSS.n2696 VSS.n2695 4.5005
R4388 VSS.n2273 VSS.n2271 4.5005
R4389 VSS.n2312 VSS.n2279 4.5005
R4390 VSS.n2686 VSS.n2685 4.5005
R4391 VSS.n2694 VSS.n2241 4.5005
R4392 VSS.n2715 VSS.n2215 4.5005
R4393 VSS.n2220 VSS.n2216 4.5005
R4394 VSS.n2225 VSS.n2223 4.5005
R4395 VSS.n2741 VSS.n2167 4.5005
R4396 VSS.n2206 VSS.n2198 4.5005
R4397 VSS.n2163 VSS.n2162 4.5005
R4398 VSS.n2759 VSS.n2123 4.5005
R4399 VSS.n2771 VSS.n2110 4.5005
R4400 VSS.n2121 VSS.n2116 4.5005
R4401 VSS.n2100 VSS.n2098 4.5005
R4402 VSS.n2770 VSS.n2769 4.5005
R4403 VSS.n2122 VSS.n2119 4.5005
R4404 VSS.n2160 VSS.n2146 4.5005
R4405 VSS.n2782 VSS.n2097 4.5005
R4406 VSS.n2203 VSS.n2173 4.5005
R4407 VSS.n2168 VSS.n2166 4.5005
R4408 VSS.n2749 VSS.n2748 4.5005
R4409 VSS.n2208 VSS.n2207 4.5005
R4410 VSS.n2743 VSS.n2742 4.5005
R4411 VSS.n2763 VSS.n2762 4.5005
R4412 VSS.n2111 VSS.n2104 4.5005
R4413 VSS.n2784 VSS.n2783 4.5005
R4414 VSS.n2205 VSS.n2204 4.5005
R4415 VSS.n2009 VSS.n2006 4.5005
R4416 VSS.n2863 VSS.n2862 4.5005
R4417 VSS.n2838 VSS.n2837 4.5005
R4418 VSS.n2043 VSS.n2042 4.5005
R4419 VSS.n2030 VSS.n2029 4.5005
R4420 VSS.n2049 VSS.n2044 4.5005
R4421 VSS.n2003 VSS.n1999 4.5005
R4422 VSS.n2872 VSS.n1998 4.5005
R4423 VSS.n2861 VSS.n2010 4.5005
R4424 VSS.n2075 VSS.n2064 4.5005
R4425 VSS.n2807 VSS.n2086 4.5005
R4426 VSS.n2832 VSS.n2062 4.5005
R4427 VSS.n2809 VSS.n2808 4.5005
R4428 VSS.n2076 VSS.n2072 4.5005
R4429 VSS.n2034 VSS.n2033 4.5005
R4430 VSS.n2834 VSS.n2833 4.5005
R4431 VSS.n2848 VSS.n2847 4.5005
R4432 VSS.n2084 VSS.n2077 4.5005
R4433 VSS.n2811 VSS.n2810 4.5005
R4434 VSS.n2874 VSS.n2873 4.5005
R4435 VSS.n4189 VSS.n4188 4.5005
R4436 VSS.n4149 VSS.n4148 4.5005
R4437 VSS.n4212 VSS.n4211 4.5005
R4438 VSS.n4211 VSS.n4210 4.5005
R4439 VSS.n4685 VSS.n4684 4.5005
R4440 VSS.n1416 VSS.n1415 4.5005
R4441 VSS.n4088 VSS.n4087 4.5005
R4442 VSS.n4087 VSS.n4086 4.5005
R4443 VSS.n4125 VSS.n4124 4.5005
R4444 VSS.n4124 VSS.n4123 4.5005
R4445 VSS.n966 VSS.n965 4.5005
R4446 VSS.n212 VSS.t514 4.44646
R4447 VSS.t196 VSS.t199 4.44646
R4448 VSS.n4137 VSS.n4136 4.25879
R4449 VSS.n919 VSS.n918 4.25822
R4450 VSS.n5935 VSS.n5934 4.22638
R4451 VSS.t258 VSS.t193 4.12487
R4452 VSS.t193 VSS.t196 4.12487
R4453 VSS.n4718 VSS.t128 4.12487
R4454 VSS.n5874 VSS.n5871 4.11115
R4455 VSS.n5874 VSS.n5873 4.0918
R4456 VSS VSS.n5918 4.0484
R4457 VSS VSS.n5924 4.0484
R4458 VSS VSS.n5786 4.0484
R4459 VSS VSS.n5842 4.0484
R4460 VSS.n816 VSS.t639 4.04279
R4461 VSS.n841 VSS.t641 4.04279
R4462 VSS.n1457 VSS.t625 4.04279
R4463 VSS.n1473 VSS.t36 4.04279
R4464 VSS.n911 VSS.n910 3.95365
R4465 VSS.n971 VSS.n970 3.95358
R4466 VSS VSS.n5901 3.86981
R4467 VSS.n5913 VSS.n5909 3.76876
R4468 VSS.n5914 VSS.n5907 3.76876
R4469 VSS.n5848 VSS.n5776 3.76876
R4470 VSS.n5847 VSS.n5778 3.76876
R4471 VSS.n4199 VSS.t67 3.75122
R4472 VSS.n26 VSS.n24 3.68267
R4473 VSS.n5850 VSS.n5771 3.66898
R4474 VSS.n5933 VSS.n4748 3.66898
R4475 VSS.n5774 VSS.n5773 3.66898
R4476 VSS.n5868 VSS.n5740 3.60687
R4477 VSS.n5884 VSS.n5883 3.60246
R4478 VSS.n5798 VSS.n5797 3.60246
R4479 VSS.n5832 VSS.n5831 3.60246
R4480 VSS.n4274 VSS.n4273 3.59971
R4481 VSS.n5869 VSS.n5738 3.5873
R4482 VSS.n1029 VSS.n1028 3.48846
R4483 VSS.n1719 VSS.t707 3.45416
R4484 VSS.n1728 VSS.t710 3.45416
R4485 VSS.n1720 VSS.t708 3.45416
R4486 VSS.n1754 VSS.t333 3.41655
R4487 VSS.n2458 VSS.t387 3.41655
R4488 VSS.n2372 VSS.t309 3.41655
R4489 VSS.n2255 VSS.t339 3.41655
R4490 VSS.n2148 VSS.t292 3.41655
R4491 VSS.n2051 VSS.t369 3.41655
R4492 VSS.n1981 VSS.t368 3.41655
R4493 VSS.n1826 VSS.t365 3.41655
R4494 VSS.n1792 VSS.t320 3.41655
R4495 VSS.n1771 VSS.t316 3.41655
R4496 VSS.n1743 VSS.t343 3.41655
R4497 VSS.n4854 VSS.t620 3.41078
R4498 VSS.n4817 VSS.t667 3.41078
R4499 VSS.n4929 VSS.t754 3.41078
R4500 VSS.n4811 VSS.t78 3.41078
R4501 VSS VSS.n5759 3.41059
R4502 VSS.n5766 VSS.n5765 3.40289
R4503 VSS.n1382 VSS.t106 3.38064
R4504 VSS.n4094 VSS.t479 3.38064
R4505 VSS.n922 VSS.n921 3.37941
R4506 VSS.n1414 VSS.n1411 3.37941
R4507 VSS.n1414 VSS.n1413 3.37941
R4508 VSS.n4013 VSS.n3986 3.37941
R4509 VSS.n835 VSS.n822 3.37941
R4510 VSS.n835 VSS.n824 3.37941
R4511 VSS.n4853 VSS.n4852 3.37941
R4512 VSS.n4816 VSS.n4815 3.37941
R4513 VSS.n4810 VSS.n4809 3.37941
R4514 VSS.n4928 VSS.n4927 3.37941
R4515 VSS.n4153 VSS.n4152 3.37941
R4516 VSS.n4709 VSS.n4706 3.37941
R4517 VSS.n4709 VSS.n4708 3.37941
R4518 VSS.n4116 VSS.n4115 3.3685
R4519 VSS.n4108 VSS.n4107 3.35882
R4520 VSS.n5746 VSS.n5745 3.3442
R4521 VSS.n5754 VSS.n5753 3.3442
R4522 VSS.n4510 VSS.t249 3.333
R4523 VSS.n5066 VSS.t224 3.33271
R4524 VSS.n76 VSS.t273 3.33057
R4525 VSS.n5064 VSS.t251 3.33036
R4526 VSS.n4965 VSS.t271 3.32608
R4527 VSS.n4964 VSS.t278 3.32608
R4528 VSS.n4925 VSS.t235 3.32608
R4529 VSS.n4807 VSS.t219 3.32608
R4530 VSS.n33 VSS.t222 3.32582
R4531 VSS.n32 VSS.t240 3.32582
R4532 VSS.n31 VSS.t256 3.32582
R4533 VSS.n58 VSS.t247 3.32582
R4534 VSS.n4806 VSS.t280 3.32512
R4535 VSS.n59 VSS.t191 3.32486
R4536 VSS.n4511 VSS.t238 3.31238
R4537 VSS.n5077 VSS.t216 3.31209
R4538 VSS.n63 VSS.t188 3.31186
R4539 VSS.n5063 VSS.t283 3.3116
R4540 VSS.n94 VSS.t230 3.31143
R4541 VSS.n5065 VSS.t179 3.31114
R4542 VSS.n6064 VSS.n6063 3.30479
R4543 VSS.n5745 VSS.t13 3.2765
R4544 VSS.n5745 VSS.n5744 3.2765
R4545 VSS.n5738 VSS.t474 3.2765
R4546 VSS.n5738 VSS.n5737 3.2765
R4547 VSS.n5873 VSS.t706 3.2765
R4548 VSS.n5873 VSS.n5872 3.2765
R4549 VSS.n5871 VSS.t102 3.2765
R4550 VSS.n5871 VSS.n5870 3.2765
R4551 VSS.n5740 VSS.t421 3.2765
R4552 VSS.n5740 VSS.n5739 3.2765
R4553 VSS.n5753 VSS.t700 3.2765
R4554 VSS.n5753 VSS.n5752 3.2765
R4555 VSS.n5765 VSS.t85 3.2765
R4556 VSS.n5765 VSS.n5764 3.2765
R4557 VSS.n5759 VSS.t50 3.2765
R4558 VSS.n5759 VSS.n5758 3.2765
R4559 VSS.n231 VSS.t460 3.2765
R4560 VSS.n231 VSS.n230 3.2765
R4561 VSS.n234 VSS.t560 3.2765
R4562 VSS.n234 VSS.n233 3.2765
R4563 VSS.n237 VSS.t161 3.2765
R4564 VSS.n237 VSS.n236 3.2765
R4565 VSS.n179 VSS.t454 3.2765
R4566 VSS.n179 VSS.n178 3.2765
R4567 VSS.n182 VSS.t526 3.2765
R4568 VSS.n182 VSS.n181 3.2765
R4569 VSS.n176 VSS.t565 3.2765
R4570 VSS.n176 VSS.n175 3.2765
R4571 VSS.n172 VSS.t521 3.2765
R4572 VSS.n172 VSS.n171 3.2765
R4573 VSS.n169 VSS.t447 3.2765
R4574 VSS.n169 VSS.n168 3.2765
R4575 VSS.n125 VSS.t534 3.2765
R4576 VSS.n125 VSS.n124 3.2765
R4577 VSS.n129 VSS.t568 3.2765
R4578 VSS.n129 VSS.n128 3.2765
R4579 VSS.n133 VSS.t547 3.2765
R4580 VSS.n133 VSS.n132 3.2765
R4581 VSS.n136 VSS.t537 3.2765
R4582 VSS.n136 VSS.n135 3.2765
R4583 VSS.n139 VSS.t573 3.2765
R4584 VSS.n139 VSS.n138 3.2765
R4585 VSS.n223 VSS.t553 3.2765
R4586 VSS.n223 VSS.n222 3.2765
R4587 VSS.n227 VSS.t154 3.2765
R4588 VSS.n227 VSS.n226 3.2765
R4589 VSS.n921 VSS.t115 3.2765
R4590 VSS.n921 VSS.n920 3.2765
R4591 VSS.n1413 VSS.t765 3.2765
R4592 VSS.n1413 VSS.n1412 3.2765
R4593 VSS.n1411 VSS.t626 3.2765
R4594 VSS.n1411 VSS.n1410 3.2765
R4595 VSS.n3986 VSS.t33 3.2765
R4596 VSS.n3986 VSS.n3985 3.2765
R4597 VSS.n824 VSS.t679 3.2765
R4598 VSS.n824 VSS.n823 3.2765
R4599 VSS.n822 VSS.t640 3.2765
R4600 VSS.n822 VSS.n821 3.2765
R4601 VSS.n5183 VSS.t556 3.2765
R4602 VSS.n5183 VSS.n5182 3.2765
R4603 VSS.n5185 VSS.t443 3.2765
R4604 VSS.n5185 VSS.n5184 3.2765
R4605 VSS.n5187 VSS.t603 3.2765
R4606 VSS.n5187 VSS.n5186 3.2765
R4607 VSS.n5212 VSS.t445 3.2765
R4608 VSS.n5212 VSS.n5211 3.2765
R4609 VSS.n5210 VSS.t524 3.2765
R4610 VSS.n5210 VSS.n5209 3.2765
R4611 VSS.n5208 VSS.t569 3.2765
R4612 VSS.n5208 VSS.n5207 3.2765
R4613 VSS.n5204 VSS.t159 3.2765
R4614 VSS.n5204 VSS.n5203 3.2765
R4615 VSS.n5206 VSS.t463 3.2765
R4616 VSS.n5206 VSS.n5205 3.2765
R4617 VSS.n5179 VSS.t604 3.2765
R4618 VSS.n5179 VSS.n5178 3.2765
R4619 VSS.n5181 VSS.t444 3.2765
R4620 VSS.n5181 VSS.n5180 3.2765
R4621 VSS.n4792 VSS.t507 3.2765
R4622 VSS.n4792 VSS.n4791 3.2765
R4623 VSS.n4790 VSS.t552 3.2765
R4624 VSS.n4790 VSS.n4789 3.2765
R4625 VSS.n4788 VSS.t598 3.2765
R4626 VSS.n4788 VSS.n4787 3.2765
R4627 VSS.n4786 VSS.t505 3.2765
R4628 VSS.n4786 VSS.n4785 3.2765
R4629 VSS.n4784 VSS.t527 3.2765
R4630 VSS.n4784 VSS.n4783 3.2765
R4631 VSS.n4852 VSS.t621 3.2765
R4632 VSS.n4852 VSS.n4851 3.2765
R4633 VSS.n4815 VSS.t668 3.2765
R4634 VSS.n4815 VSS.n4814 3.2765
R4635 VSS.n4809 VSS.t79 3.2765
R4636 VSS.n4809 VSS.n4808 3.2765
R4637 VSS.n4927 VSS.t755 3.2765
R4638 VSS.n4927 VSS.n4926 3.2765
R4639 VSS.n4152 VSS.t499 3.2765
R4640 VSS.n4152 VSS.n4151 3.2765
R4641 VSS.n4708 VSS.t586 3.2765
R4642 VSS.n4708 VSS.n4707 3.2765
R4643 VSS.n4706 VSS.t132 3.2765
R4644 VSS.n4706 VSS.n4705 3.2765
R4645 VSS.n4745 VSS.n4743 3.17523
R4646 VSS.n140 VSS.n139 3.1505
R4647 VSS.n137 VSS.n136 3.1505
R4648 VSS.n130 VSS.n129 3.1505
R4649 VSS.n228 VSS.n227 3.1505
R4650 VSS.n173 VSS.n172 3.1505
R4651 VSS.n183 VSS.n182 3.1505
R4652 VSS.n180 VSS.n179 3.1505
R4653 VSS.n238 VSS.n237 3.1505
R4654 VSS.n235 VSS.n234 3.1505
R4655 VSS.n5192 VSS.n5181 3.1505
R4656 VSS.n5193 VSS.n5179 3.1505
R4657 VSS.n5218 VSS.n5206 3.1505
R4658 VSS.n5219 VSS.n5204 3.1505
R4659 VSS.n5215 VSS.n5210 3.1505
R4660 VSS.n4799 VSS.n4784 3.1505
R4661 VSS.n4798 VSS.n4786 3.1505
R4662 VSS.n4795 VSS.n4790 3.1505
R4663 VSS.n5189 VSS.n5185 3.1505
R4664 VSS.n5985 VSS.n5984 3.08765
R4665 VSS.n4682 VSS.n4681 3.07743
R4666 VSS.n4124 VSS.n916 2.9883
R4667 VSS.n4087 VSS.n1397 2.9883
R4668 VSS.n4745 VSS.n4744 2.91648
R4669 VSS.n4993 VSS.n4992 2.83943
R4670 VSS.n4989 VSS.n4988 2.83943
R4671 VSS.n4985 VSS.n4984 2.83943
R4672 VSS.n4679 VSS.n4678 2.83943
R4673 VSS.n4676 VSS.n4675 2.83943
R4674 VSS.n4662 VSS.n4661 2.83943
R4675 VSS.n4584 VSS.n4583 2.83943
R4676 VSS.n4588 VSS.n4587 2.83943
R4677 VSS.n1311 VSS.n1310 2.81354
R4678 VSS.n3914 VSS.n3908 2.7874
R4679 VSS.n4236 VSS.n4235 2.75024
R4680 VSS.n1021 VSS.n1017 2.65705
R4681 VSS.n1021 VSS.n1020 2.65638
R4682 VSS.n4860 VSS.n4859 2.64393
R4683 VSS.n4822 VSS.n4821 2.64393
R4684 VSS.n134 VSS.n133 2.6255
R4685 VSS.n170 VSS.n169 2.6255
R4686 VSS.n177 VSS.n176 2.6255
R4687 VSS.n232 VSS.n231 2.6255
R4688 VSS.n5217 VSS.n5208 2.6255
R4689 VSS.n4797 VSS.n4788 2.6255
R4690 VSS.n5188 VSS.n5187 2.6255
R4691 VSS.n5191 VSS.n5183 2.6255
R4692 VSS.n5460 VSS.n5420 2.61042
R4693 VSS.n5444 VSS.n5422 2.61042
R4694 VSS.n5555 VSS.n5474 2.61042
R4695 VSS.n5619 VSS.n5618 2.60873
R4696 VSS.n4064 VSS.n1399 2.60616
R4697 VSS.n4040 VSS.n4039 2.60562
R4698 VSS.n1424 VSS.n1421 2.60491
R4699 VSS.n1481 VSS.n1480 2.60491
R4700 VSS.n796 VSS.n793 2.60491
R4701 VSS.n862 VSS.n861 2.60491
R4702 VSS.n4778 VSS.n4777 2.60246
R4703 VSS.n5325 VSS.n5324 2.60244
R4704 VSS.n5304 VSS.n5300 2.60244
R4705 VSS.n117 VSS.n110 2.60148
R4706 VSS.n4411 VSS.n4394 2.60147
R4707 VSS.n5767 VSS 2.6005
R4708 VSS.n5768 VSS.n5767 2.6005
R4709 VSS VSS.n5763 2.6005
R4710 VSS.n5763 VSS.n5762 2.6005
R4711 VSS.n5861 VSS.n5860 2.6005
R4712 VSS.n5860 VSS.n5859 2.6005
R4713 VSS.n5761 VSS 2.6005
R4714 VSS.n5761 VSS.n5760 2.6005
R4715 VSS.n1308 VSS.n958 2.6005
R4716 VSS.n958 VSS.n957 2.6005
R4717 VSS.n1324 VSS.n1323 2.6005
R4718 VSS.n1323 VSS.n1322 2.6005
R4719 VSS.n1320 VSS.n1319 2.6005
R4720 VSS.n1319 VSS.n1318 2.6005
R4721 VSS.n1316 VSS.n1315 2.6005
R4722 VSS.n1315 VSS.n1314 2.6005
R4723 VSS.n1313 VSS.n1312 2.6005
R4724 VSS.n1312 VSS.n1311 2.6005
R4725 VSS.n1326 VSS.n1325 2.6005
R4726 VSS.n926 VSS.n925 2.6005
R4727 VSS.n929 VSS.n928 2.6005
R4728 VSS.n931 VSS.n930 2.6005
R4729 VSS.n933 VSS.n932 2.6005
R4730 VSS VSS.n935 2.6005
R4731 VSS.n937 VSS.n936 2.6005
R4732 VSS.n942 VSS.n941 2.6005
R4733 VSS.n945 VSS.n944 2.6005
R4734 VSS.n947 VSS.n946 2.6005
R4735 VSS.n950 VSS.n949 2.6005
R4736 VSS.n1340 VSS.n1339 2.6005
R4737 VSS.n1338 VSS.n1337 2.6005
R4738 VSS.n1336 VSS.n1335 2.6005
R4739 VSS.n1332 VSS.n1331 2.6005
R4740 VSS.n1330 VSS.n1329 2.6005
R4741 VSS.n1403 VSS.n1400 2.6005
R4742 VSS.n1520 VSS.n1517 2.6005
R4743 VSS.n4002 VSS.n3999 2.6005
R4744 VSS.n4012 VSS.n4009 2.6005
R4745 VSS.n4025 VSS.n4023 2.6005
R4746 VSS.n3984 VSS.n3983 2.6005
R4747 VSS.n3983 VSS.n3982 2.6005
R4748 VSS.n4030 VSS.n4029 2.6005
R4749 VSS.n4029 VSS.n4028 2.6005
R4750 VSS.n4026 VSS.n4025 2.6005
R4751 VSS.n4019 VSS.n4018 2.6005
R4752 VSS.n4018 VSS.n4017 2.6005
R4753 VSS VSS.n4012 2.6005
R4754 VSS.n4007 VSS.n4006 2.6005
R4755 VSS.n4006 VSS.n4005 2.6005
R4756 VSS.n4003 VSS.n4002 2.6005
R4757 VSS.n3993 VSS.n3992 2.6005
R4758 VSS.n3992 VSS.n3991 2.6005
R4759 VSS.n1521 VSS.n1520 2.6005
R4760 VSS.n3980 VSS.n3979 2.6005
R4761 VSS.n3979 VSS.n3978 2.6005
R4762 VSS.n5011 VSS.n4805 2.6005
R4763 VSS.n4805 VSS.n4804 2.6005
R4764 VSS.n5003 VSS.n5002 2.6005
R4765 VSS.n5002 VSS.n5001 2.6005
R4766 VSS.n5006 VSS.n5005 2.6005
R4767 VSS.n5005 VSS.n5004 2.6005
R4768 VSS.n5010 VSS.n5009 2.6005
R4769 VSS.n5009 VSS.n5008 2.6005
R4770 VSS.n5017 VSS.n5016 2.6005
R4771 VSS.n5016 VSS.n5015 2.6005
R4772 VSS.n4973 VSS.n4972 2.6005
R4773 VSS.n5486 VSS.n5485 2.6005
R4774 VSS.n5485 VSS.n5484 2.6005
R4775 VSS.n5483 VSS.n5482 2.6005
R4776 VSS.n5482 VSS.n5481 2.6005
R4777 VSS.n4969 VSS.n4968 2.6005
R4778 VSS.n4968 VSS.n4967 2.6005
R4779 VSS.n4972 VSS.n4971 2.6005
R4780 VSS.n5489 VSS.n5488 2.6005
R4781 VSS.n5488 VSS.n5487 2.6005
R4782 VSS.n4976 VSS.n4975 2.6005
R4783 VSS.n4975 VSS.n4974 2.6005
R4784 VSS.n4980 VSS.n4979 2.6005
R4785 VSS.n4982 VSS.n4981 2.6005
R4786 VSS.n4986 VSS.n4985 2.6005
R4787 VSS.n4990 VSS.n4989 2.6005
R4788 VSS.n4893 VSS.n4892 2.6005
R4789 VSS.n4892 VSS.n4891 2.6005
R4790 VSS.n4897 VSS.n4896 2.6005
R4791 VSS.n4896 VSS.n4895 2.6005
R4792 VSS.n4900 VSS.n4899 2.6005
R4793 VSS.n4899 VSS.n4898 2.6005
R4794 VSS.n4903 VSS.n4902 2.6005
R4795 VSS.n4902 VSS.n4901 2.6005
R4796 VSS.n4904 VSS.n4812 2.6005
R4797 VSS.n4812 VSS.n4811 2.6005
R4798 VSS.n4906 VSS 2.6005
R4799 VSS.n4906 VSS.n4905 2.6005
R4800 VSS.n4909 VSS.n4908 2.6005
R4801 VSS.n4908 VSS.n4907 2.6005
R4802 VSS.n4912 VSS.n4911 2.6005
R4803 VSS.n4911 VSS.n4910 2.6005
R4804 VSS.n4917 VSS.n4916 2.6005
R4805 VSS.n4916 VSS.n4915 2.6005
R4806 VSS.n4920 VSS.n4919 2.6005
R4807 VSS.n4919 VSS.n4918 2.6005
R4808 VSS.n4924 VSS.n4923 2.6005
R4809 VSS.n4923 VSS.n4922 2.6005
R4810 VSS.n4994 VSS.n4993 2.6005
R4811 VSS.n4999 VSS.n4998 2.6005
R4812 VSS.n4888 VSS.n4887 2.6005
R4813 VSS.n4887 VSS.n4886 2.6005
R4814 VSS.n4863 VSS.n4862 2.6005
R4815 VSS.n4862 VSS.n4861 2.6005
R4816 VSS.n4866 VSS.n4865 2.6005
R4817 VSS.n4865 VSS.n4864 2.6005
R4818 VSS.n4869 VSS.n4868 2.6005
R4819 VSS.n4868 VSS.n4867 2.6005
R4820 VSS.n4870 VSS.n4855 2.6005
R4821 VSS.n4855 VSS.n4854 2.6005
R4822 VSS.n4872 VSS 2.6005
R4823 VSS.n4872 VSS.n4871 2.6005
R4824 VSS.n4875 VSS.n4874 2.6005
R4825 VSS.n4874 VSS.n4873 2.6005
R4826 VSS.n4878 VSS.n4877 2.6005
R4827 VSS.n4877 VSS.n4876 2.6005
R4828 VSS.n4881 VSS.n4880 2.6005
R4829 VSS.n4880 VSS.n4879 2.6005
R4830 VSS.n4884 VSS.n4883 2.6005
R4831 VSS.n4883 VSS.n4882 2.6005
R4832 VSS.n4859 VSS.n4858 2.6005
R4833 VSS.n4821 VSS.n4820 2.6005
R4834 VSS.n4825 VSS.n4824 2.6005
R4835 VSS.n4824 VSS.n4823 2.6005
R4836 VSS.n4828 VSS.n4827 2.6005
R4837 VSS.n4827 VSS.n4826 2.6005
R4838 VSS.n4831 VSS.n4830 2.6005
R4839 VSS.n4830 VSS.n4829 2.6005
R4840 VSS.n4832 VSS.n4818 2.6005
R4841 VSS.n4818 VSS.n4817 2.6005
R4842 VSS.n4834 VSS 2.6005
R4843 VSS.n4834 VSS.n4833 2.6005
R4844 VSS.n4837 VSS.n4836 2.6005
R4845 VSS.n4836 VSS.n4835 2.6005
R4846 VSS.n4840 VSS.n4839 2.6005
R4847 VSS.n4839 VSS.n4838 2.6005
R4848 VSS.n4843 VSS.n4842 2.6005
R4849 VSS.n4842 VSS.n4841 2.6005
R4850 VSS.n4846 VSS.n4845 2.6005
R4851 VSS.n4845 VSS.n4844 2.6005
R4852 VSS.n4850 VSS.n4849 2.6005
R4853 VSS.n4849 VSS.n4848 2.6005
R4854 VSS.n4934 VSS.n4933 2.6005
R4855 VSS.n4933 VSS.n4932 2.6005
R4856 VSS.n4938 VSS.n4937 2.6005
R4857 VSS.n4937 VSS.n4936 2.6005
R4858 VSS.n4941 VSS.n4940 2.6005
R4859 VSS.n4940 VSS.n4939 2.6005
R4860 VSS.n4944 VSS.n4943 2.6005
R4861 VSS.n4943 VSS.n4942 2.6005
R4862 VSS.n4945 VSS.n4930 2.6005
R4863 VSS.n4930 VSS.n4929 2.6005
R4864 VSS.n4947 VSS 2.6005
R4865 VSS.n4947 VSS.n4946 2.6005
R4866 VSS.n4950 VSS.n4949 2.6005
R4867 VSS.n4949 VSS.n4948 2.6005
R4868 VSS.n4953 VSS.n4952 2.6005
R4869 VSS.n4952 VSS.n4951 2.6005
R4870 VSS.n4956 VSS.n4955 2.6005
R4871 VSS.n4955 VSS.n4954 2.6005
R4872 VSS.n4959 VSS.n4958 2.6005
R4873 VSS.n4958 VSS.n4957 2.6005
R4874 VSS.n4963 VSS.n4962 2.6005
R4875 VSS.n4962 VSS.n4961 2.6005
R4876 VSS.n470 VSS.n469 2.6005
R4877 VSS.n862 VSS.n858 2.6005
R4878 VSS.n858 VSS.n857 2.6005
R4879 VSS.n800 VSS.n799 2.6005
R4880 VSS.n799 VSS.n798 2.6005
R4881 VSS.n806 VSS.n805 2.6005
R4882 VSS.n805 VSS.n804 2.6005
R4883 VSS.n812 VSS.n811 2.6005
R4884 VSS.n811 VSS.n810 2.6005
R4885 VSS.n818 VSS.n817 2.6005
R4886 VSS.n817 VSS.n816 2.6005
R4887 VSS.n837 VSS 2.6005
R4888 VSS.n837 VSS.n836 2.6005
R4889 VSS.n840 VSS.n839 2.6005
R4890 VSS.n839 VSS.n838 2.6005
R4891 VSS.n846 VSS.n845 2.6005
R4892 VSS.n845 VSS.n844 2.6005
R4893 VSS.n853 VSS.n852 2.6005
R4894 VSS.n852 VSS.n851 2.6005
R4895 VSS.n869 VSS.n868 2.6005
R4896 VSS.n868 VSS.n867 2.6005
R4897 VSS.n793 VSS.n792 2.6005
R4898 VSS.n834 VSS.n831 2.6005
R4899 VSS.n803 VSS.n802 2.6005
R4900 VSS.n802 VSS.n801 2.6005
R4901 VSS.n809 VSS.n808 2.6005
R4902 VSS.n808 VSS.n807 2.6005
R4903 VSS.n815 VSS.n814 2.6005
R4904 VSS.n814 VSS.n813 2.6005
R4905 VSS.n828 VSS.n827 2.6005
R4906 VSS VSS.n834 2.6005
R4907 VSS.n843 VSS.n842 2.6005
R4908 VSS.n842 VSS.n841 2.6005
R4909 VSS.n850 VSS.n849 2.6005
R4910 VSS.n849 VSS.n848 2.6005
R4911 VSS.n856 VSS.n855 2.6005
R4912 VSS.n855 VSS.n854 2.6005
R4913 VSS.n866 VSS.n865 2.6005
R4914 VSS.n865 VSS.n864 2.6005
R4915 VSS.n861 VSS.n860 2.6005
R4916 VSS.n796 VSS.n795 2.6005
R4917 VSS.n795 VSS.n794 2.6005
R4918 VSS.n257 VSS.n256 2.6005
R4919 VSS.n342 VSS.n339 2.6005
R4920 VSS.n343 VSS.n342 2.6005
R4921 VSS.n4049 VSS.n4048 2.6005
R4922 VSS.n4067 VSS.n4066 2.6005
R4923 VSS.n4066 VSS.n4065 2.6005
R4924 VSS.n1399 VSS.n1398 2.6005
R4925 VSS.n4063 VSS.n4062 2.6005
R4926 VSS.n4062 VSS.n4061 2.6005
R4927 VSS.n4060 VSS.n4059 2.6005
R4928 VSS.n4059 VSS.n4058 2.6005
R4929 VSS.n4057 VSS.n4056 2.6005
R4930 VSS.n4056 VSS.n4055 2.6005
R4931 VSS.n4053 VSS.n4052 2.6005
R4932 VSS.n4052 VSS.n4051 2.6005
R4933 VSS.n4048 VSS.n4047 2.6005
R4934 VSS.n371 VSS.n370 2.6005
R4935 VSS.n370 VSS.n369 2.6005
R4936 VSS.n374 VSS.n373 2.6005
R4937 VSS.n373 VSS.n372 2.6005
R4938 VSS.n377 VSS.n376 2.6005
R4939 VSS.n376 VSS.n375 2.6005
R4940 VSS.n380 VSS.n379 2.6005
R4941 VSS.n379 VSS.n378 2.6005
R4942 VSS.n383 VSS.n382 2.6005
R4943 VSS.n382 VSS.n381 2.6005
R4944 VSS.n386 VSS.n385 2.6005
R4945 VSS.n385 VSS.n384 2.6005
R4946 VSS.n389 VSS.n388 2.6005
R4947 VSS.n388 VSS.n387 2.6005
R4948 VSS.n393 VSS.n392 2.6005
R4949 VSS.n392 VSS.n391 2.6005
R4950 VSS.n396 VSS.n395 2.6005
R4951 VSS.n395 VSS.n394 2.6005
R4952 VSS.n399 VSS.n398 2.6005
R4953 VSS.n398 VSS.n397 2.6005
R4954 VSS.n402 VSS.n401 2.6005
R4955 VSS.n401 VSS.n400 2.6005
R4956 VSS.n405 VSS.n404 2.6005
R4957 VSS.n404 VSS.n403 2.6005
R4958 VSS.n409 VSS.n408 2.6005
R4959 VSS.n408 VSS.n407 2.6005
R4960 VSS.n412 VSS.n411 2.6005
R4961 VSS.n411 VSS.n410 2.6005
R4962 VSS.n416 VSS.n415 2.6005
R4963 VSS.n415 VSS.n414 2.6005
R4964 VSS.n419 VSS.n418 2.6005
R4965 VSS.n418 VSS.n417 2.6005
R4966 VSS.n422 VSS.n421 2.6005
R4967 VSS.n421 VSS.n420 2.6005
R4968 VSS.n427 VSS.n426 2.6005
R4969 VSS.n426 VSS.n425 2.6005
R4970 VSS.n430 VSS.n429 2.6005
R4971 VSS.n429 VSS.n428 2.6005
R4972 VSS.n433 VSS.n432 2.6005
R4973 VSS.n432 VSS.n431 2.6005
R4974 VSS.n436 VSS.n435 2.6005
R4975 VSS.n435 VSS.n434 2.6005
R4976 VSS.n439 VSS.n438 2.6005
R4977 VSS.n438 VSS.n437 2.6005
R4978 VSS.n442 VSS.n441 2.6005
R4979 VSS.n441 VSS.n440 2.6005
R4980 VSS.n445 VSS.n444 2.6005
R4981 VSS.n444 VSS.n443 2.6005
R4982 VSS.n448 VSS.n447 2.6005
R4983 VSS.n447 VSS.n446 2.6005
R4984 VSS.n451 VSS.n450 2.6005
R4985 VSS.n450 VSS.n449 2.6005
R4986 VSS.n454 VSS.n453 2.6005
R4987 VSS.n453 VSS.n452 2.6005
R4988 VSS.n458 VSS.n457 2.6005
R4989 VSS.n457 VSS.n456 2.6005
R4990 VSS.n461 VSS.n460 2.6005
R4991 VSS.n460 VSS.n459 2.6005
R4992 VSS.n464 VSS.n463 2.6005
R4993 VSS.n463 VSS.n462 2.6005
R4994 VSS.n473 VSS.n472 2.6005
R4995 VSS.n472 VSS.n471 2.6005
R4996 VSS.n476 VSS.n475 2.6005
R4997 VSS.n475 VSS.n474 2.6005
R4998 VSS.n479 VSS.n478 2.6005
R4999 VSS.n478 VSS.n477 2.6005
R5000 VSS.n482 VSS.n481 2.6005
R5001 VSS.n481 VSS.n480 2.6005
R5002 VSS.n485 VSS.n484 2.6005
R5003 VSS.n484 VSS.n483 2.6005
R5004 VSS.n487 VSS.n486 2.6005
R5005 VSS.n491 VSS.n490 2.6005
R5006 VSS.n493 VSS.n492 2.6005
R5007 VSS.n763 VSS.n762 2.6005
R5008 VSS.n716 VSS.n715 2.6005
R5009 VSS.n715 VSS.n714 2.6005
R5010 VSS.n762 VSS.n761 2.6005
R5011 VSS.n760 VSS.n759 2.6005
R5012 VSS.n759 VSS.n758 2.6005
R5013 VSS.n757 VSS.n756 2.6005
R5014 VSS.n756 VSS.n755 2.6005
R5015 VSS.n754 VSS.n753 2.6005
R5016 VSS.n753 VSS.n752 2.6005
R5017 VSS.n732 VSS.n731 2.6005
R5018 VSS.n731 VSS.n730 2.6005
R5019 VSS.n728 VSS.n727 2.6005
R5020 VSS.n727 VSS.n726 2.6005
R5021 VSS.n725 VSS.n724 2.6005
R5022 VSS.n724 VSS.n723 2.6005
R5023 VSS.n722 VSS.n721 2.6005
R5024 VSS.n721 VSS.n720 2.6005
R5025 VSS.n719 VSS.n718 2.6005
R5026 VSS.n718 VSS.n717 2.6005
R5027 VSS.n497 VSS.n496 2.6005
R5028 VSS.n496 VSS.n495 2.6005
R5029 VSS.n500 VSS.n499 2.6005
R5030 VSS.n502 VSS.n501 2.6005
R5031 VSS.n5353 VSS.n5352 2.6005
R5032 VSS.n5349 VSS.n5348 2.6005
R5033 VSS.n5346 VSS.n5345 2.6005
R5034 VSS.n5343 VSS.n5342 2.6005
R5035 VSS.n5341 VSS.n5340 2.6005
R5036 VSS.n5338 VSS.n5337 2.6005
R5037 VSS.n5337 VSS.n5336 2.6005
R5038 VSS.n5334 VSS.n5333 2.6005
R5039 VSS.n5333 VSS.n5332 2.6005
R5040 VSS.n514 VSS.n513 2.6005
R5041 VSS.n513 VSS.n512 2.6005
R5042 VSS.n517 VSS.n516 2.6005
R5043 VSS.n516 VSS.n515 2.6005
R5044 VSS.n520 VSS.n519 2.6005
R5045 VSS.n519 VSS.n518 2.6005
R5046 VSS.n523 VSS.n522 2.6005
R5047 VSS.n522 VSS.n521 2.6005
R5048 VSS.n526 VSS.n525 2.6005
R5049 VSS.n525 VSS.n524 2.6005
R5050 VSS.n530 VSS.n529 2.6005
R5051 VSS.n529 VSS.n528 2.6005
R5052 VSS.n533 VSS.n532 2.6005
R5053 VSS.n532 VSS.n531 2.6005
R5054 VSS.n536 VSS.n535 2.6005
R5055 VSS.n535 VSS.n534 2.6005
R5056 VSS.n539 VSS.n538 2.6005
R5057 VSS.n538 VSS.n537 2.6005
R5058 VSS.n542 VSS.n541 2.6005
R5059 VSS.n541 VSS.n540 2.6005
R5060 VSS.n545 VSS.n544 2.6005
R5061 VSS.n544 VSS.n543 2.6005
R5062 VSS.n548 VSS.n547 2.6005
R5063 VSS.n547 VSS.n546 2.6005
R5064 VSS.n551 VSS.n550 2.6005
R5065 VSS.n550 VSS.n549 2.6005
R5066 VSS.n554 VSS.n553 2.6005
R5067 VSS.n556 VSS.n555 2.6005
R5068 VSS.n559 VSS.n558 2.6005
R5069 VSS.n562 VSS.n561 2.6005
R5070 VSS.n566 VSS.n565 2.6005
R5071 VSS.n571 VSS.n570 2.6005
R5072 VSS.n570 VSS.n569 2.6005
R5073 VSS.n574 VSS.n573 2.6005
R5074 VSS.n573 VSS.n572 2.6005
R5075 VSS.n577 VSS.n576 2.6005
R5076 VSS.n576 VSS.n575 2.6005
R5077 VSS.n580 VSS.n579 2.6005
R5078 VSS.n579 VSS.n578 2.6005
R5079 VSS.n583 VSS.n582 2.6005
R5080 VSS.n582 VSS.n581 2.6005
R5081 VSS.n586 VSS.n585 2.6005
R5082 VSS.n585 VSS.n584 2.6005
R5083 VSS.n589 VSS.n588 2.6005
R5084 VSS.n588 VSS.n587 2.6005
R5085 VSS.n593 VSS.n592 2.6005
R5086 VSS.n592 VSS.n591 2.6005
R5087 VSS.n595 VSS.n594 2.6005
R5088 VSS.n598 VSS.n597 2.6005
R5089 VSS.n601 VSS.n600 2.6005
R5090 VSS.n600 VSS.n599 2.6005
R5091 VSS.n604 VSS.n603 2.6005
R5092 VSS.n603 VSS.n602 2.6005
R5093 VSS.n607 VSS.n606 2.6005
R5094 VSS.n606 VSS.n605 2.6005
R5095 VSS.n610 VSS.n609 2.6005
R5096 VSS.n609 VSS.n608 2.6005
R5097 VSS.n613 VSS.n612 2.6005
R5098 VSS.n612 VSS.n611 2.6005
R5099 VSS.n616 VSS.n615 2.6005
R5100 VSS.n615 VSS.n614 2.6005
R5101 VSS.n619 VSS.n618 2.6005
R5102 VSS.n618 VSS.n617 2.6005
R5103 VSS.n622 VSS.n621 2.6005
R5104 VSS.n621 VSS.n620 2.6005
R5105 VSS.n625 VSS.n624 2.6005
R5106 VSS.n624 VSS.n623 2.6005
R5107 VSS.n628 VSS.n627 2.6005
R5108 VSS.n627 VSS.n626 2.6005
R5109 VSS.n631 VSS.n630 2.6005
R5110 VSS.n630 VSS.n629 2.6005
R5111 VSS.n634 VSS.n633 2.6005
R5112 VSS.n633 VSS.n632 2.6005
R5113 VSS.n637 VSS.n636 2.6005
R5114 VSS.n636 VSS.n635 2.6005
R5115 VSS.n640 VSS.n639 2.6005
R5116 VSS.n639 VSS.n638 2.6005
R5117 VSS.n643 VSS.n642 2.6005
R5118 VSS.n642 VSS.n641 2.6005
R5119 VSS.n646 VSS.n645 2.6005
R5120 VSS.n645 VSS.n644 2.6005
R5121 VSS.n649 VSS.n648 2.6005
R5122 VSS.n648 VSS.n647 2.6005
R5123 VSS.n652 VSS.n651 2.6005
R5124 VSS.n651 VSS.n650 2.6005
R5125 VSS.n655 VSS.n654 2.6005
R5126 VSS.n654 VSS.n653 2.6005
R5127 VSS.n658 VSS.n657 2.6005
R5128 VSS.n657 VSS.n656 2.6005
R5129 VSS.n661 VSS.n660 2.6005
R5130 VSS.n660 VSS.n659 2.6005
R5131 VSS.n664 VSS.n663 2.6005
R5132 VSS.n663 VSS.n662 2.6005
R5133 VSS.n667 VSS.n666 2.6005
R5134 VSS.n666 VSS.n665 2.6005
R5135 VSS.n670 VSS.n669 2.6005
R5136 VSS.n669 VSS.n668 2.6005
R5137 VSS.n673 VSS.n672 2.6005
R5138 VSS.n675 VSS.n674 2.6005
R5139 VSS.n678 VSS.n677 2.6005
R5140 VSS.n681 VSS.n680 2.6005
R5141 VSS.n685 VSS.n684 2.6005
R5142 VSS.n691 VSS.n690 2.6005
R5143 VSS.n687 VSS.n686 2.6005
R5144 VSS.n735 VSS.n734 2.6005
R5145 VSS.n734 VSS.n733 2.6005
R5146 VSS.n713 VSS.n712 2.6005
R5147 VSS.n712 VSS.n711 2.6005
R5148 VSS.n710 VSS.n709 2.6005
R5149 VSS.n709 VSS.n708 2.6005
R5150 VSS.n707 VSS.n706 2.6005
R5151 VSS.n706 VSS.n705 2.6005
R5152 VSS.n704 VSS.n703 2.6005
R5153 VSS.n703 VSS.n702 2.6005
R5154 VSS.n506 VSS.n505 2.6005
R5155 VSS.n509 VSS.n508 2.6005
R5156 VSS.n700 VSS.n699 2.6005
R5157 VSS.n699 VSS.n698 2.6005
R5158 VSS.n697 VSS.n696 2.6005
R5159 VSS.n696 VSS.n695 2.6005
R5160 VSS.n694 VSS.n693 2.6005
R5161 VSS.n693 VSS.n692 2.6005
R5162 VSS.n775 VSS.n255 2.6005
R5163 VSS.n255 VSS.n254 2.6005
R5164 VSS.n787 VSS.n786 2.6005
R5165 VSS.n786 VSS.n785 2.6005
R5166 VSS.n784 VSS.n783 2.6005
R5167 VSS.n783 VSS.n782 2.6005
R5168 VSS.n781 VSS.n780 2.6005
R5169 VSS.n780 VSS.n779 2.6005
R5170 VSS.n778 VSS.n777 2.6005
R5171 VSS.n777 VSS.n776 2.6005
R5172 VSS.n751 VSS.n750 2.6005
R5173 VSS.n750 VSS.n749 2.6005
R5174 VSS.n748 VSS.n747 2.6005
R5175 VSS.n747 VSS.n746 2.6005
R5176 VSS.n745 VSS.n744 2.6005
R5177 VSS.n744 VSS.n743 2.6005
R5178 VSS.n742 VSS.n741 2.6005
R5179 VSS.n741 VSS.n740 2.6005
R5180 VSS.n739 VSS.n738 2.6005
R5181 VSS.n738 VSS.n737 2.6005
R5182 VSS.n770 VSS.n769 2.6005
R5183 VSS.n769 VSS.n768 2.6005
R5184 VSS.n773 VSS.n772 2.6005
R5185 VSS.n772 VSS.n771 2.6005
R5186 VSS.n766 VSS.n765 2.6005
R5187 VSS.n765 VSS.n764 2.6005
R5188 VSS.n4298 VSS.n4297 2.6005
R5189 VSS.n4297 VSS.n4296 2.6005
R5190 VSS.n4295 VSS.n4294 2.6005
R5191 VSS.n4294 VSS.n4293 2.6005
R5192 VSS.n4292 VSS.n4291 2.6005
R5193 VSS.n4291 VSS.n4290 2.6005
R5194 VSS.n4289 VSS.n4288 2.6005
R5195 VSS.n4288 VSS.n4287 2.6005
R5196 VSS.n4301 VSS.n4300 2.6005
R5197 VSS.n4312 VSS.n4311 2.6005
R5198 VSS.n4307 VSS.n4306 2.6005
R5199 VSS.n1174 VSS.n1173 2.6005
R5200 VSS.n1173 VSS.n1172 2.6005
R5201 VSS.n1178 VSS.n1177 2.6005
R5202 VSS.n1177 VSS.n1176 2.6005
R5203 VSS.n1181 VSS.n1180 2.6005
R5204 VSS.n1180 VSS.n1179 2.6005
R5205 VSS.n1184 VSS.n1183 2.6005
R5206 VSS.n1183 VSS.n1182 2.6005
R5207 VSS.n1187 VSS.n1186 2.6005
R5208 VSS.n1186 VSS.n1185 2.6005
R5209 VSS.n1190 VSS.n1189 2.6005
R5210 VSS.n1189 VSS.n1188 2.6005
R5211 VSS.n1193 VSS.n1192 2.6005
R5212 VSS.n1192 VSS.n1191 2.6005
R5213 VSS.n1196 VSS.n1195 2.6005
R5214 VSS.n1195 VSS.n1194 2.6005
R5215 VSS.n1199 VSS.n1198 2.6005
R5216 VSS.n1198 VSS.n1197 2.6005
R5217 VSS.n1171 VSS.n1170 2.6005
R5218 VSS.n1342 VSS.n1341 2.6005
R5219 VSS.n1345 VSS.n1344 2.6005
R5220 VSS.n1347 VSS.n1346 2.6005
R5221 VSS.n1350 VSS.n1349 2.6005
R5222 VSS.n1352 VSS.n1351 2.6005
R5223 VSS.n1355 VSS.n1354 2.6005
R5224 VSS.n1357 VSS.n1356 2.6005
R5225 VSS.n1360 VSS.n1359 2.6005
R5226 VSS.n1362 VSS.n1361 2.6005
R5227 VSS.n1365 VSS.n1364 2.6005
R5228 VSS.n1367 VSS.n1366 2.6005
R5229 VSS.n1371 VSS.n1370 2.6005
R5230 VSS.n1377 VSS.n1376 2.6005
R5231 VSS.n1376 VSS.n1375 2.6005
R5232 VSS.n1374 VSS.n1373 2.6005
R5233 VSS.n1373 VSS.n1372 2.6005
R5234 VSS.n4193 VSS.n4190 2.6005
R5235 VSS.n4158 VSS.n4150 2.6005
R5236 VSS.n4140 VSS.n4139 2.6005
R5237 VSS.n4143 VSS.n4142 2.6005
R5238 VSS.n4145 VSS.n4144 2.6005
R5239 VSS.n4159 VSS.n4158 2.6005
R5240 VSS.n4155 VSS 2.6005
R5241 VSS.n4155 VSS.n4154 2.6005
R5242 VSS.n4180 VSS.n4179 2.6005
R5243 VSS.n4184 VSS.n4183 2.6005
R5244 VSS.n4183 VSS.n4182 2.6005
R5245 VSS.n4194 VSS.n4193 2.6005
R5246 VSS.n4197 VSS.n4196 2.6005
R5247 VSS.n4201 VSS.n4200 2.6005
R5248 VSS.n4200 VSS.n4199 2.6005
R5249 VSS.n4229 VSS.n4228 2.6005
R5250 VSS.n4228 VSS.n4227 2.6005
R5251 VSS.n4226 VSS.n4225 2.6005
R5252 VSS.n4225 VSS.n4224 2.6005
R5253 VSS.n4223 VSS.n4222 2.6005
R5254 VSS.n4222 VSS.n4221 2.6005
R5255 VSS.n893 VSS.n892 2.6005
R5256 VSS.n892 VSS.n891 2.6005
R5257 VSS.n895 VSS.n894 2.6005
R5258 VSS.n897 VSS.n896 2.6005
R5259 VSS.n899 VSS.n898 2.6005
R5260 VSS.n902 VSS.n901 2.6005
R5261 VSS.n905 VSS.n904 2.6005
R5262 VSS.n907 VSS.n906 2.6005
R5263 VSS.n4255 VSS.n4254 2.6005
R5264 VSS.n4349 VSS.n4348 2.6005
R5265 VSS.n4345 VSS.n4344 2.6005
R5266 VSS.n4343 VSS.n4342 2.6005
R5267 VSS.n4340 VSS.n4339 2.6005
R5268 VSS.n4337 VSS.n4336 2.6005
R5269 VSS.n4270 VSS.n4269 2.6005
R5270 VSS.n4269 VSS.n4268 2.6005
R5271 VSS.n4267 VSS.n4266 2.6005
R5272 VSS.n4266 VSS.n4265 2.6005
R5273 VSS.n4264 VSS.n4263 2.6005
R5274 VSS.n4263 VSS.n4262 2.6005
R5275 VSS.n4261 VSS.n4260 2.6005
R5276 VSS.n4260 VSS.n4259 2.6005
R5277 VSS.n4258 VSS.n4257 2.6005
R5278 VSS.n4257 VSS.n4256 2.6005
R5279 VSS.n4254 VSS.n4253 2.6005
R5280 VSS.n4319 VSS.n4318 2.6005
R5281 VSS.n4315 VSS.n4314 2.6005
R5282 VSS.n4286 VSS.n4285 2.6005
R5283 VSS.n4285 VSS.n4284 2.6005
R5284 VSS.n4334 VSS.n4333 2.6005
R5285 VSS.n4330 VSS.n4329 2.6005
R5286 VSS.n4327 VSS.n4326 2.6005
R5287 VSS.n4324 VSS.n4323 2.6005
R5288 VSS.n4321 VSS.n4320 2.6005
R5289 VSS.n4278 VSS.n4277 2.6005
R5290 VSS.n4280 VSS.n4279 2.6005
R5291 VSS.n4283 VSS.n4282 2.6005
R5292 VSS.n4614 VSS.n4613 2.6005
R5293 VSS.n4613 VSS.n4612 2.6005
R5294 VSS.n4617 VSS.n4616 2.6005
R5295 VSS.n4616 VSS.n4615 2.6005
R5296 VSS.n4620 VSS.n4619 2.6005
R5297 VSS.n4619 VSS.n4618 2.6005
R5298 VSS.n4623 VSS.n4622 2.6005
R5299 VSS.n4622 VSS.n4621 2.6005
R5300 VSS.n4626 VSS.n4625 2.6005
R5301 VSS.n4625 VSS.n4624 2.6005
R5302 VSS.n4629 VSS.n4628 2.6005
R5303 VSS.n4628 VSS.n4627 2.6005
R5304 VSS.n4632 VSS.n4631 2.6005
R5305 VSS.n4631 VSS.n4630 2.6005
R5306 VSS.n4635 VSS.n4634 2.6005
R5307 VSS.n4634 VSS.n4633 2.6005
R5308 VSS.n4638 VSS.n4637 2.6005
R5309 VSS.n4637 VSS.n4636 2.6005
R5310 VSS.n4641 VSS.n4640 2.6005
R5311 VSS.n4640 VSS.n4639 2.6005
R5312 VSS.n4644 VSS.n4643 2.6005
R5313 VSS.n4643 VSS.n4642 2.6005
R5314 VSS.n4647 VSS.n4646 2.6005
R5315 VSS.n4646 VSS.n4645 2.6005
R5316 VSS.n4650 VSS.n4649 2.6005
R5317 VSS.n4649 VSS.n4648 2.6005
R5318 VSS.n4653 VSS.n4652 2.6005
R5319 VSS.n4652 VSS.n4651 2.6005
R5320 VSS.n116 VSS.n115 2.6005
R5321 VSS.n115 VSS.n114 2.6005
R5322 VSS.n113 VSS.n112 2.6005
R5323 VSS.n112 VSS.n111 2.6005
R5324 VSS.n123 VSS.n122 2.6005
R5325 VSS.n122 VSS.n121 2.6005
R5326 VSS.n198 VSS.n197 2.6005
R5327 VSS.n197 VSS.n196 2.6005
R5328 VSS.n201 VSS.n200 2.6005
R5329 VSS.n200 VSS.n199 2.6005
R5330 VSS.n204 VSS.n203 2.6005
R5331 VSS.n203 VSS.n202 2.6005
R5332 VSS.n194 VSS.n193 2.6005
R5333 VSS.n193 VSS.n192 2.6005
R5334 VSS.n208 VSS.n207 2.6005
R5335 VSS.n207 VSS.n206 2.6005
R5336 VSS.n211 VSS.n210 2.6005
R5337 VSS.n210 VSS.n209 2.6005
R5338 VSS.n214 VSS.n213 2.6005
R5339 VSS.n213 VSS.n212 2.6005
R5340 VSS.n218 VSS.n217 2.6005
R5341 VSS.n217 VSS.n216 2.6005
R5342 VSS.n191 VSS.n190 2.6005
R5343 VSS.n190 VSS.n189 2.6005
R5344 VSS.n187 VSS.n186 2.6005
R5345 VSS.n186 VSS.n185 2.6005
R5346 VSS.n167 VSS.n166 2.6005
R5347 VSS.n166 VSS.n165 2.6005
R5348 VSS.n164 VSS.n163 2.6005
R5349 VSS.n163 VSS.n162 2.6005
R5350 VSS.n251 VSS.n250 2.6005
R5351 VSS.n247 VSS.n246 2.6005
R5352 VSS.n120 VSS.n119 2.6005
R5353 VSS.n4391 VSS.n4390 2.6005
R5354 VSS.n4389 VSS.n4388 2.6005
R5355 VSS.n4385 VSS.n4384 2.6005
R5356 VSS.n101 VSS.n100 2.6005
R5357 VSS.n160 VSS.n159 2.6005
R5358 VSS.n159 VSS.n158 2.6005
R5359 VSS.n157 VSS.n156 2.6005
R5360 VSS.n156 VSS.n155 2.6005
R5361 VSS.n154 VSS.n153 2.6005
R5362 VSS.n153 VSS.n152 2.6005
R5363 VSS.n151 VSS.n150 2.6005
R5364 VSS.n150 VSS.n149 2.6005
R5365 VSS.n62 VSS.n61 2.6005
R5366 VSS.n61 VSS.n60 2.6005
R5367 VSS.n4611 VSS.n4610 2.6005
R5368 VSS.n4605 VSS.n4604 2.6005
R5369 VSS.n4600 VSS.n4599 2.6005
R5370 VSS.n4608 VSS.n4607 2.6005
R5371 VSS.n4597 VSS.n4596 2.6005
R5372 VSS.n4594 VSS.n4593 2.6005
R5373 VSS.n4589 VSS.n4588 2.6005
R5374 VSS.n4585 VSS.n4584 2.6005
R5375 VSS.n4581 VSS.n4580 2.6005
R5376 VSS.n4578 VSS.n4577 2.6005
R5377 VSS.n4656 VSS.n4655 2.6005
R5378 VSS.n4655 VSS.n4654 2.6005
R5379 VSS.n4660 VSS.n4659 2.6005
R5380 VSS.n4663 VSS.n4662 2.6005
R5381 VSS.n4666 VSS.n4665 2.6005
R5382 VSS.n4669 VSS.n4668 2.6005
R5383 VSS.n4673 VSS.n4672 2.6005
R5384 VSS.n4677 VSS.n4676 2.6005
R5385 VSS.n4680 VSS.n4679 2.6005
R5386 VSS.n54 VSS.n53 2.6005
R5387 VSS.n56 VSS.n55 2.6005
R5388 VSS.n4738 VSS.n4736 2.6005
R5389 VSS.n4736 VSS.n4735 2.6005
R5390 VSS.n4696 VSS.n4694 2.6005
R5391 VSS.n4694 VSS.n4693 2.6005
R5392 VSS.n4700 VSS.n4698 2.6005
R5393 VSS.n4698 VSS.n4697 2.6005
R5394 VSS.n4704 VSS.n4702 2.6005
R5395 VSS.n4702 VSS.n4701 2.6005
R5396 VSS.n4715 VSS.n4713 2.6005
R5397 VSS.n4715 VSS.n4714 2.6005
R5398 VSS.n4717 VSS 2.6005
R5399 VSS.n4717 VSS.n4716 2.6005
R5400 VSS.n4720 VSS.n4719 2.6005
R5401 VSS.n4719 VSS.n4718 2.6005
R5402 VSS.n4724 VSS.n4721 2.6005
R5403 VSS.n4728 VSS.n4726 2.6005
R5404 VSS.n4726 VSS.n4725 2.6005
R5405 VSS.n4732 VSS.n4729 2.6005
R5406 VSS.n4690 VSS.n4683 2.6005
R5407 VSS.n4696 VSS.n4695 2.6005
R5408 VSS.n4700 VSS.n4699 2.6005
R5409 VSS.n4704 VSS.n4703 2.6005
R5410 VSS.n4713 VSS.n4712 2.6005
R5411 VSS.n4711 VSS 2.6005
R5412 VSS.n4724 VSS.n4723 2.6005
R5413 VSS.n4723 VSS.n4722 2.6005
R5414 VSS.n4728 VSS.n4727 2.6005
R5415 VSS.n4732 VSS.n4731 2.6005
R5416 VSS.n4731 VSS.n4730 2.6005
R5417 VSS.n4738 VSS.n4737 2.6005
R5418 VSS.n4690 VSS.n4689 2.6005
R5419 VSS.n4689 VSS.n4688 2.6005
R5420 VSS.n5993 VSS.n5992 2.6005
R5421 VSS.n5995 VSS.n5994 2.6005
R5422 VSS.n5998 VSS.n5997 2.6005
R5423 VSS.n6000 VSS.n5999 2.6005
R5424 VSS.n6003 VSS.n6002 2.6005
R5425 VSS.n6005 VSS.n6004 2.6005
R5426 VSS.n6009 VSS.n6008 2.6005
R5427 VSS.n6012 VSS.n6011 2.6005
R5428 VSS.n6014 VSS.n6013 2.6005
R5429 VSS.n6017 VSS.n6016 2.6005
R5430 VSS.n6022 VSS.n6021 2.6005
R5431 VSS.n6025 VSS.n6024 2.6005
R5432 VSS.n6027 VSS.n6026 2.6005
R5433 VSS.n6030 VSS.n6029 2.6005
R5434 VSS.n6033 VSS.n6032 2.6005
R5435 VSS.n6036 VSS.n6035 2.6005
R5436 VSS.n6040 VSS.n6039 2.6005
R5437 VSS.n1531 VSS.n1530 2.6005
R5438 VSS.n1530 VSS.n1529 2.6005
R5439 VSS.n1534 VSS.n1533 2.6005
R5440 VSS.n1533 VSS.n1532 2.6005
R5441 VSS.n3910 VSS.n3909 2.6005
R5442 VSS.n3912 VSS.n3911 2.6005
R5443 VSS.n3918 VSS.n3917 2.6005
R5444 VSS.n3917 VSS.n3916 2.6005
R5445 VSS.n3921 VSS.n3920 2.6005
R5446 VSS.n3920 VSS.n3919 2.6005
R5447 VSS.n3924 VSS.n3923 2.6005
R5448 VSS.n3923 VSS.n3922 2.6005
R5449 VSS.n3927 VSS.n3926 2.6005
R5450 VSS.n3926 VSS.n3925 2.6005
R5451 VSS.n3930 VSS.n3929 2.6005
R5452 VSS.n3929 VSS.n3928 2.6005
R5453 VSS.n3934 VSS.n3933 2.6005
R5454 VSS.n3933 VSS.n3932 2.6005
R5455 VSS.n3937 VSS.n3936 2.6005
R5456 VSS.n3936 VSS.n3935 2.6005
R5457 VSS.n3940 VSS.n3939 2.6005
R5458 VSS.n3939 VSS.n3938 2.6005
R5459 VSS.n3943 VSS.n3942 2.6005
R5460 VSS.n3942 VSS.n3941 2.6005
R5461 VSS.n3946 VSS.n3945 2.6005
R5462 VSS.n3945 VSS.n3944 2.6005
R5463 VSS.n3949 VSS.n3948 2.6005
R5464 VSS.n3948 VSS.n3947 2.6005
R5465 VSS.n3952 VSS.n3951 2.6005
R5466 VSS.n3951 VSS.n3950 2.6005
R5467 VSS.n3955 VSS.n3954 2.6005
R5468 VSS.n3954 VSS.n3953 2.6005
R5469 VSS.n3958 VSS.n3957 2.6005
R5470 VSS.n3957 VSS.n3956 2.6005
R5471 VSS.n3961 VSS.n3960 2.6005
R5472 VSS.n3960 VSS.n3959 2.6005
R5473 VSS.n3964 VSS.n3963 2.6005
R5474 VSS.n3963 VSS.n3962 2.6005
R5475 VSS.n3967 VSS.n3966 2.6005
R5476 VSS.n3966 VSS.n3965 2.6005
R5477 VSS.n3970 VSS.n3969 2.6005
R5478 VSS.n3969 VSS.n3968 2.6005
R5479 VSS.n3973 VSS.n3972 2.6005
R5480 VSS.n3972 VSS.n3971 2.6005
R5481 VSS.n3976 VSS.n3975 2.6005
R5482 VSS.n3975 VSS.n3974 2.6005
R5483 VSS.n4039 VSS.n4038 2.6005
R5484 VSS.n4046 VSS.n4045 2.6005
R5485 VSS.n4042 VSS.n4041 2.6005
R5486 VSS.n4037 VSS.n4036 2.6005
R5487 VSS.n4036 VSS.n4035 2.6005
R5488 VSS.n4034 VSS.n4033 2.6005
R5489 VSS.n4033 VSS.n4032 2.6005
R5490 VSS.n1528 VSS.n1527 2.6005
R5491 VSS.n1527 VSS.n1526 2.6005
R5492 VSS.n366 VSS.n365 2.6005
R5493 VSS.n368 VSS.n367 2.6005
R5494 VSS.n362 VSS.n361 2.6005
R5495 VSS.n1481 VSS.n1477 2.6005
R5496 VSS.n1477 VSS.n1476 2.6005
R5497 VSS.n1428 VSS.n1427 2.6005
R5498 VSS.n1427 VSS.n1426 2.6005
R5499 VSS.n1434 VSS.n1433 2.6005
R5500 VSS.n1433 VSS.n1432 2.6005
R5501 VSS.n1440 VSS.n1439 2.6005
R5502 VSS.n1439 VSS.n1438 2.6005
R5503 VSS.n1458 VSS.n1456 2.6005
R5504 VSS.n1458 VSS.n1457 2.6005
R5505 VSS VSS.n1460 2.6005
R5506 VSS.n1460 VSS.n1459 2.6005
R5507 VSS.n1472 VSS.n1471 2.6005
R5508 VSS.n1471 VSS.n1470 2.6005
R5509 VSS.n1500 VSS.n1499 2.6005
R5510 VSS.n1499 VSS.n1498 2.6005
R5511 VSS.n1494 VSS.n1493 2.6005
R5512 VSS.n1493 VSS.n1492 2.6005
R5513 VSS.n1488 VSS.n1487 2.6005
R5514 VSS.n1487 VSS.n1486 2.6005
R5515 VSS.n1421 VSS.n1420 2.6005
R5516 VSS VSS.n1468 2.6005
R5517 VSS.n1468 VSS.n1467 2.6005
R5518 VSS.n1475 VSS.n1474 2.6005
R5519 VSS.n1474 VSS.n1473 2.6005
R5520 VSS.n1497 VSS.n1496 2.6005
R5521 VSS.n1496 VSS.n1495 2.6005
R5522 VSS.n1491 VSS.n1490 2.6005
R5523 VSS.n1490 VSS.n1489 2.6005
R5524 VSS.n1485 VSS.n1484 2.6005
R5525 VSS.n1484 VSS.n1483 2.6005
R5526 VSS.n1480 VSS.n1479 2.6005
R5527 VSS.n1424 VSS.n1423 2.6005
R5528 VSS.n1423 VSS.n1422 2.6005
R5529 VSS.n1431 VSS.n1430 2.6005
R5530 VSS.n1430 VSS.n1429 2.6005
R5531 VSS.n1437 VSS.n1436 2.6005
R5532 VSS.n1436 VSS.n1435 2.6005
R5533 VSS.n1443 VSS.n1442 2.6005
R5534 VSS.n1442 VSS.n1441 2.6005
R5535 VSS.n1464 VSS.n1462 2.6005
R5536 VSS.n1464 VSS.n1463 2.6005
R5537 VSS.n1380 VSS.n1379 2.6005
R5538 VSS.n1379 VSS.n1378 2.6005
R5539 VSS.n1384 VSS.n1383 2.6005
R5540 VSS.n1383 VSS.n1382 2.6005
R5541 VSS.n1387 VSS.n1386 2.6005
R5542 VSS.n1386 VSS.n1385 2.6005
R5543 VSS.n1391 VSS.n1390 2.6005
R5544 VSS.n1390 VSS.n1389 2.6005
R5545 VSS.n4096 VSS.n4095 2.6005
R5546 VSS.n4095 VSS.n4094 2.6005
R5547 VSS.n4099 VSS.n4098 2.6005
R5548 VSS.n4098 VSS.n4097 2.6005
R5549 VSS.n4117 VSS.n4101 2.6005
R5550 VSS.n4101 VSS.n4100 2.6005
R5551 VSS.n4114 VSS.n4113 2.6005
R5552 VSS.n4104 VSS.n4103 2.6005
R5553 VSS.n4111 VSS.n4110 2.6005
R5554 VSS.n4110 VSS.n4109 2.6005
R5555 VSS.n4073 VSS.n4072 2.6005
R5556 VSS.n4072 VSS.n4071 2.6005
R5557 VSS.n4076 VSS.n4075 2.6005
R5558 VSS.n4075 VSS.n4074 2.6005
R5559 VSS.n4079 VSS.n4078 2.6005
R5560 VSS.n4078 VSS.n4077 2.6005
R5561 VSS.n4082 VSS.n4081 2.6005
R5562 VSS.n4081 VSS.n4080 2.6005
R5563 VSS.n4084 VSS.n4083 2.6005
R5564 VSS.n4085 VSS.n4084 2.6005
R5565 VSS.n4070 VSS.n4069 2.6005
R5566 VSS.n4069 VSS.n4068 2.6005
R5567 VSS.n1203 VSS.n1202 2.6005
R5568 VSS.n1202 VSS.n1201 2.6005
R5569 VSS.n1206 VSS.n1205 2.6005
R5570 VSS.n1205 VSS.n1204 2.6005
R5571 VSS.n1209 VSS.n1208 2.6005
R5572 VSS.n1208 VSS.n1207 2.6005
R5573 VSS.n1212 VSS.n1211 2.6005
R5574 VSS.n1211 VSS.n1210 2.6005
R5575 VSS.n1215 VSS.n1214 2.6005
R5576 VSS.n1214 VSS.n1213 2.6005
R5577 VSS.n1218 VSS.n1217 2.6005
R5578 VSS.n1217 VSS.n1216 2.6005
R5579 VSS.n1221 VSS.n1220 2.6005
R5580 VSS.n1220 VSS.n1219 2.6005
R5581 VSS.n1224 VSS.n1223 2.6005
R5582 VSS.n1223 VSS.n1222 2.6005
R5583 VSS.n1228 VSS.n1227 2.6005
R5584 VSS.n1227 VSS.n1226 2.6005
R5585 VSS.n1231 VSS.n1230 2.6005
R5586 VSS.n1230 VSS.n1229 2.6005
R5587 VSS.n1234 VSS.n1233 2.6005
R5588 VSS.n1233 VSS.n1232 2.6005
R5589 VSS.n1237 VSS.n1236 2.6005
R5590 VSS.n1236 VSS.n1235 2.6005
R5591 VSS.n1240 VSS.n1239 2.6005
R5592 VSS.n1239 VSS.n1238 2.6005
R5593 VSS.n1243 VSS.n1242 2.6005
R5594 VSS.n1242 VSS.n1241 2.6005
R5595 VSS.n1246 VSS.n1245 2.6005
R5596 VSS.n1245 VSS.n1244 2.6005
R5597 VSS.n1249 VSS.n1248 2.6005
R5598 VSS.n1248 VSS.n1247 2.6005
R5599 VSS.n1307 VSS.n1306 2.6005
R5600 VSS.n1304 VSS.n1303 2.6005
R5601 VSS.n1301 VSS.n1300 2.6005
R5602 VSS.n4241 VSS.n4240 2.6005
R5603 VSS.n4237 VSS.n4236 2.6005
R5604 VSS.n4234 VSS.n4233 2.6005
R5605 VSS.n4232 VSS.n4231 2.6005
R5606 VSS.n1283 VSS.n1282 2.6005
R5607 VSS.n1280 VSS.n1279 2.6005
R5608 VSS.n1277 VSS.n1276 2.6005
R5609 VSS.n1274 VSS.n1273 2.6005
R5610 VSS.n1271 VSS.n1270 2.6005
R5611 VSS.n1268 VSS.n1267 2.6005
R5612 VSS.n1265 VSS.n1264 2.6005
R5613 VSS.n1262 VSS.n1261 2.6005
R5614 VSS.n1259 VSS.n1258 2.6005
R5615 VSS.n1257 VSS.n1256 2.6005
R5616 VSS.n1251 VSS.n1250 2.6005
R5617 VSS.n1250 VSS.t652 2.6005
R5618 VSS.n1254 VSS.n1253 2.6005
R5619 VSS.n1253 VSS.n1252 2.6005
R5620 VSS.n1284 VSS.n974 2.6005
R5621 VSS.n1290 VSS.n1289 2.6005
R5622 VSS.n1297 VSS.n1296 2.6005
R5623 VSS.n1296 VSS.n1295 2.6005
R5624 VSS.n1293 VSS.n1292 2.6005
R5625 VSS.n1292 VSS.n1291 2.6005
R5626 VSS.n4251 VSS.n4250 2.6005
R5627 VSS.n4250 VSS.n4249 2.6005
R5628 VSS.n4247 VSS.n4246 2.6005
R5629 VSS.n4246 VSS.n4245 2.6005
R5630 VSS.n4244 VSS.n4243 2.6005
R5631 VSS.n4243 VSS.n4242 2.6005
R5632 VSS.n1288 VSS.n1287 2.6005
R5633 VSS.n38 VSS.n37 2.6005
R5634 VSS.n41 VSS.n40 2.6005
R5635 VSS.n44 VSS.n43 2.6005
R5636 VSS.n46 VSS.n45 2.6005
R5637 VSS.n51 VSS.n50 2.6005
R5638 VSS.n4575 VSS.n4574 2.6005
R5639 VSS.n4569 VSS.n4568 2.6005
R5640 VSS.n4564 VSS.n4563 2.6005
R5641 VSS.n4567 VSS.n4566 2.6005
R5642 VSS.n4560 VSS.n4559 2.6005
R5643 VSS.n4427 VSS.n4426 2.6005
R5644 VSS.n4424 VSS.n4423 2.6005
R5645 VSS.n4422 VSS.n4421 2.6005
R5646 VSS.n99 VSS.n98 2.6005
R5647 VSS.n976 VSS.n975 2.6005
R5648 VSS.n980 VSS.n979 2.6005
R5649 VSS.n4354 VSS.n4353 2.6005
R5650 VSS.n4418 VSS.n4417 2.6005
R5651 VSS.n4413 VSS.n4412 2.6005
R5652 VSS.n4351 VSS.n4350 2.6005
R5653 VSS.n4430 VSS.n4429 2.6005
R5654 VSS.n4429 VSS.n4428 2.6005
R5655 VSS.n4439 VSS.n4438 2.6005
R5656 VSS.n4438 VSS.n4437 2.6005
R5657 VSS.n4443 VSS.n4442 2.6005
R5658 VSS.n4442 VSS.n4441 2.6005
R5659 VSS.n4446 VSS.n4445 2.6005
R5660 VSS.n4445 VSS.n4444 2.6005
R5661 VSS.n4449 VSS.n4448 2.6005
R5662 VSS.n4448 VSS.n4447 2.6005
R5663 VSS.n4452 VSS.n4451 2.6005
R5664 VSS.n4451 VSS.n4450 2.6005
R5665 VSS.n4455 VSS.n4454 2.6005
R5666 VSS.n4454 VSS.n4453 2.6005
R5667 VSS.n4458 VSS.n4457 2.6005
R5668 VSS.n4457 VSS.n4456 2.6005
R5669 VSS.n4461 VSS.n4460 2.6005
R5670 VSS.n4460 VSS.n4459 2.6005
R5671 VSS.n4464 VSS.n4463 2.6005
R5672 VSS.n4463 VSS.n4462 2.6005
R5673 VSS.n4467 VSS.n4466 2.6005
R5674 VSS.n4466 VSS.n4465 2.6005
R5675 VSS.n4471 VSS.n4470 2.6005
R5676 VSS.n4470 VSS.n4469 2.6005
R5677 VSS.n4474 VSS.n4473 2.6005
R5678 VSS.n4473 VSS.n4472 2.6005
R5679 VSS.n4477 VSS.n4476 2.6005
R5680 VSS.n4476 VSS.n4475 2.6005
R5681 VSS.n4480 VSS.n4479 2.6005
R5682 VSS.n4479 VSS.n4478 2.6005
R5683 VSS.n4483 VSS.n4482 2.6005
R5684 VSS.n4482 VSS.n4481 2.6005
R5685 VSS.n4486 VSS.n4485 2.6005
R5686 VSS.n4485 VSS.n4484 2.6005
R5687 VSS.n4500 VSS.n4499 2.6005
R5688 VSS.n4499 VSS.n4498 2.6005
R5689 VSS.n4497 VSS.n4496 2.6005
R5690 VSS.n4496 VSS.n4495 2.6005
R5691 VSS.n4492 VSS.n4491 2.6005
R5692 VSS.n4491 VSS.n4490 2.6005
R5693 VSS.n4489 VSS.n4488 2.6005
R5694 VSS.n4488 VSS.n4487 2.6005
R5695 VSS.n4558 VSS.n4557 2.6005
R5696 VSS.n4555 VSS.n4554 2.6005
R5697 VSS.n4554 VSS.n4553 2.6005
R5698 VSS.n4552 VSS.n4551 2.6005
R5699 VSS.n4551 VSS.n4550 2.6005
R5700 VSS.n4549 VSS.n4548 2.6005
R5701 VSS.n4548 VSS.n4547 2.6005
R5702 VSS.n4546 VSS.n4545 2.6005
R5703 VSS.n4545 VSS.n4544 2.6005
R5704 VSS.n4543 VSS.n4542 2.6005
R5705 VSS.n4542 VSS.n4541 2.6005
R5706 VSS.n4540 VSS.n4539 2.6005
R5707 VSS.n4539 VSS.n4538 2.6005
R5708 VSS.n4537 VSS.n4536 2.6005
R5709 VSS.n4536 VSS.n4535 2.6005
R5710 VSS.n4534 VSS.n4533 2.6005
R5711 VSS.n4533 VSS.n4532 2.6005
R5712 VSS.n4531 VSS.n4530 2.6005
R5713 VSS.n4530 VSS.n4529 2.6005
R5714 VSS.n4528 VSS.n4527 2.6005
R5715 VSS.n4527 VSS.n4526 2.6005
R5716 VSS.n4525 VSS.n4524 2.6005
R5717 VSS.n4524 VSS.n4523 2.6005
R5718 VSS.n4522 VSS.n4521 2.6005
R5719 VSS.n4521 VSS.n4520 2.6005
R5720 VSS.n4519 VSS.n4518 2.6005
R5721 VSS.n4518 VSS.n4517 2.6005
R5722 VSS.n4516 VSS.n4515 2.6005
R5723 VSS.n4515 VSS.n4514 2.6005
R5724 VSS.n4513 VSS.n4512 2.6005
R5725 VSS.n35 VSS.n34 2.6005
R5726 VSS.n4433 VSS.n4432 2.6005
R5727 VSS.n4432 VSS.n4431 2.6005
R5728 VSS.n4436 VSS.n4435 2.6005
R5729 VSS.n4435 VSS.n4434 2.6005
R5730 VSS.n983 VSS.n982 2.6005
R5731 VSS.n985 VSS.n984 2.6005
R5732 VSS.n988 VSS.n987 2.6005
R5733 VSS.n992 VSS.n991 2.6005
R5734 VSS.n6067 VSS.n6066 2.6005
R5735 VSS.n6066 VSS.n6065 2.6005
R5736 VSS.n6070 VSS.n6069 2.6005
R5737 VSS.n6069 VSS.n6068 2.6005
R5738 VSS.n6074 VSS.n6073 2.6005
R5739 VSS.n6073 VSS.n6072 2.6005
R5740 VSS.n6078 VSS.n6077 2.6005
R5741 VSS.n6077 VSS.n6076 2.6005
R5742 VSS.n6081 VSS.n6080 2.6005
R5743 VSS.n6080 VSS.n6079 2.6005
R5744 VSS.n6084 VSS.n6083 2.6005
R5745 VSS.n6083 VSS.n6082 2.6005
R5746 VSS.n6087 VSS.n6086 2.6005
R5747 VSS.n6086 VSS.n6085 2.6005
R5748 VSS.n6090 VSS.n6089 2.6005
R5749 VSS.n6089 VSS.n6088 2.6005
R5750 VSS.n6092 VSS.n6091 2.6005
R5751 VSS.n6093 VSS.n6092 2.6005
R5752 VSS.n8 VSS.n7 2.6005
R5753 VSS.n7 VSS.n6 2.6005
R5754 VSS.n11 VSS.n10 2.6005
R5755 VSS.n10 VSS.n9 2.6005
R5756 VSS.n14 VSS.n13 2.6005
R5757 VSS.n13 VSS.n12 2.6005
R5758 VSS.n16 VSS.n15 2.6005
R5759 VSS.n17 VSS.n16 2.6005
R5760 VSS.n5 VSS.n4 2.6005
R5761 VSS.n4 VSS.n3 2.6005
R5762 VSS.n995 VSS.n994 2.6005
R5763 VSS.n994 VSS.n993 2.6005
R5764 VSS.n998 VSS.n997 2.6005
R5765 VSS.n997 VSS.n996 2.6005
R5766 VSS.n1002 VSS.n1001 2.6005
R5767 VSS.n1001 VSS.n1000 2.6005
R5768 VSS.n1005 VSS.n1004 2.6005
R5769 VSS.n1004 VSS.n1003 2.6005
R5770 VSS.n1008 VSS.n1007 2.6005
R5771 VSS.n1007 VSS.n1006 2.6005
R5772 VSS.n1037 VSS.n1036 2.6005
R5773 VSS.n1036 VSS.n1035 2.6005
R5774 VSS.n1040 VSS.n1039 2.6005
R5775 VSS.n1039 VSS.n1038 2.6005
R5776 VSS.n1043 VSS.n1042 2.6005
R5777 VSS.n1042 VSS.n1041 2.6005
R5778 VSS.n1046 VSS.n1045 2.6005
R5779 VSS.n1045 VSS.n1044 2.6005
R5780 VSS.n1049 VSS.n1048 2.6005
R5781 VSS.n1048 VSS.n1047 2.6005
R5782 VSS.n1052 VSS.n1051 2.6005
R5783 VSS.n1051 VSS.n1050 2.6005
R5784 VSS.n1055 VSS.n1054 2.6005
R5785 VSS.n1054 VSS.n1053 2.6005
R5786 VSS.n1058 VSS.n1057 2.6005
R5787 VSS.n1057 VSS.n1056 2.6005
R5788 VSS.n1061 VSS.n1060 2.6005
R5789 VSS.n1060 VSS.n1059 2.6005
R5790 VSS.n1064 VSS.n1063 2.6005
R5791 VSS.n1063 VSS.n1062 2.6005
R5792 VSS.n1067 VSS.n1066 2.6005
R5793 VSS.n1066 VSS.n1065 2.6005
R5794 VSS.n1070 VSS.n1069 2.6005
R5795 VSS.n1069 VSS.n1068 2.6005
R5796 VSS.n1073 VSS.n1072 2.6005
R5797 VSS.n1072 VSS.n1071 2.6005
R5798 VSS.n1076 VSS.n1075 2.6005
R5799 VSS.n1075 VSS.n1074 2.6005
R5800 VSS.n1080 VSS.n1079 2.6005
R5801 VSS.n1079 VSS.n1078 2.6005
R5802 VSS.n1083 VSS.n1082 2.6005
R5803 VSS.n1082 VSS.n1081 2.6005
R5804 VSS.n1086 VSS.n1085 2.6005
R5805 VSS.n1085 VSS.n1084 2.6005
R5806 VSS.n1089 VSS.n1088 2.6005
R5807 VSS.n1088 VSS.n1087 2.6005
R5808 VSS.n1092 VSS.n1091 2.6005
R5809 VSS.n1091 VSS.n1090 2.6005
R5810 VSS.n1095 VSS.n1094 2.6005
R5811 VSS.n1094 VSS.n1093 2.6005
R5812 VSS.n1098 VSS.n1097 2.6005
R5813 VSS.n1097 VSS.n1096 2.6005
R5814 VSS.n1101 VSS.n1100 2.6005
R5815 VSS.n1100 VSS.n1099 2.6005
R5816 VSS.n1104 VSS.n1103 2.6005
R5817 VSS.n1103 VSS.n1102 2.6005
R5818 VSS.n1107 VSS.n1106 2.6005
R5819 VSS.n1106 VSS.n1105 2.6005
R5820 VSS.n1110 VSS.n1109 2.6005
R5821 VSS.n1109 VSS.n1108 2.6005
R5822 VSS.n1113 VSS.n1112 2.6005
R5823 VSS.n1112 VSS.n1111 2.6005
R5824 VSS.n1116 VSS.n1115 2.6005
R5825 VSS.n1115 VSS.n1114 2.6005
R5826 VSS.n1119 VSS.n1118 2.6005
R5827 VSS.n1118 VSS.n1117 2.6005
R5828 VSS.n1122 VSS.n1121 2.6005
R5829 VSS.n1121 VSS.n1120 2.6005
R5830 VSS.n1125 VSS.n1124 2.6005
R5831 VSS.n1124 VSS.n1123 2.6005
R5832 VSS.n1128 VSS.n1127 2.6005
R5833 VSS.n1127 VSS.n1126 2.6005
R5834 VSS.n1131 VSS.n1130 2.6005
R5835 VSS.n1130 VSS.n1129 2.6005
R5836 VSS.n1134 VSS.n1133 2.6005
R5837 VSS.n1133 VSS.n1132 2.6005
R5838 VSS.n1137 VSS.n1136 2.6005
R5839 VSS.n1136 VSS.n1135 2.6005
R5840 VSS.n1140 VSS.n1139 2.6005
R5841 VSS.n1139 VSS.n1138 2.6005
R5842 VSS.n1143 VSS.n1142 2.6005
R5843 VSS.n1142 VSS.n1141 2.6005
R5844 VSS.n1146 VSS.n1145 2.6005
R5845 VSS.n1145 VSS.n1144 2.6005
R5846 VSS.n1149 VSS.n1148 2.6005
R5847 VSS.n1148 VSS.n1147 2.6005
R5848 VSS.n1152 VSS.n1151 2.6005
R5849 VSS.n1151 VSS.n1150 2.6005
R5850 VSS.n1155 VSS.n1154 2.6005
R5851 VSS.n1154 VSS.n1153 2.6005
R5852 VSS.n1158 VSS.n1157 2.6005
R5853 VSS.n1157 VSS.n1156 2.6005
R5854 VSS.n1161 VSS.n1160 2.6005
R5855 VSS.n1160 VSS.n1159 2.6005
R5856 VSS.n1168 VSS.n1167 2.6005
R5857 VSS.n1164 VSS.n1163 2.6005
R5858 VSS.n1163 VSS.n1162 2.6005
R5859 VSS.n6043 VSS.n6042 2.6005
R5860 VSS.n6045 VSS.n6044 2.6005
R5861 VSS.n6048 VSS.n6047 2.6005
R5862 VSS.n6051 VSS.n6050 2.6005
R5863 VSS.n6054 VSS.n6053 2.6005
R5864 VSS.n6057 VSS.n6056 2.6005
R5865 VSS.n6061 VSS.n6060 2.6005
R5866 VSS.n5622 VSS.n5621 2.6005
R5867 VSS.n5624 VSS.n5623 2.6005
R5868 VSS.n5626 VSS.n5625 2.6005
R5869 VSS.n5629 VSS.n5628 2.6005
R5870 VSS.n5632 VSS.n5631 2.6005
R5871 VSS.n5530 VSS.n5529 2.6005
R5872 VSS.n5436 VSS.n5435 2.6005
R5873 VSS.n5435 VSS.n5434 2.6005
R5874 VSS.n5433 VSS.n5432 2.6005
R5875 VSS.n5432 VSS.n5431 2.6005
R5876 VSS.n5430 VSS.n5429 2.6005
R5877 VSS.n5429 VSS.n5428 2.6005
R5878 VSS.n5426 VSS.n5425 2.6005
R5879 VSS.n5331 VSS.n5330 2.6005
R5880 VSS.n5062 VSS.n5061 2.6005
R5881 VSS.n5020 VSS.n5019 2.6005
R5882 VSS.n5019 VSS.n5018 2.6005
R5883 VSS.n5023 VSS.n5022 2.6005
R5884 VSS.n5022 VSS.n5021 2.6005
R5885 VSS.n5027 VSS.n5026 2.6005
R5886 VSS.n5026 VSS.n5025 2.6005
R5887 VSS.n5030 VSS.n5029 2.6005
R5888 VSS.n5029 VSS.n5028 2.6005
R5889 VSS.n5033 VSS.n5032 2.6005
R5890 VSS.n5032 VSS.n5031 2.6005
R5891 VSS.n5036 VSS.n5035 2.6005
R5892 VSS.n5035 VSS.n5034 2.6005
R5893 VSS.n5039 VSS.n5038 2.6005
R5894 VSS.n5038 VSS.n5037 2.6005
R5895 VSS.n5042 VSS.n5041 2.6005
R5896 VSS.n5041 VSS.n5040 2.6005
R5897 VSS.n5045 VSS.n5044 2.6005
R5898 VSS.n5044 VSS.n5043 2.6005
R5899 VSS.n5048 VSS.n5047 2.6005
R5900 VSS.n5047 VSS.n5046 2.6005
R5901 VSS.n5051 VSS.n5050 2.6005
R5902 VSS.n5050 VSS.n5049 2.6005
R5903 VSS.n5054 VSS.n5053 2.6005
R5904 VSS.n5053 VSS.n5052 2.6005
R5905 VSS.n5057 VSS.n5056 2.6005
R5906 VSS.n5056 VSS.n5055 2.6005
R5907 VSS.n5060 VSS.n5059 2.6005
R5908 VSS.n5059 VSS.n5058 2.6005
R5909 VSS.n5279 VSS.n5278 2.6005
R5910 VSS.n5649 VSS.n5648 2.6005
R5911 VSS.n5329 VSS.n5328 2.6005
R5912 VSS.n5307 VSS.n5306 2.6005
R5913 VSS.n5303 VSS.n5302 2.6005
R5914 VSS.n5639 VSS.n5638 2.6005
R5915 VSS.n5641 VSS.n5640 2.6005
R5916 VSS.n5644 VSS.n5643 2.6005
R5917 VSS.n5647 VSS.n5646 2.6005
R5918 VSS.n5636 VSS.n5635 2.6005
R5919 VSS.n4782 VSS.n4781 2.6005
R5920 VSS.n5667 VSS.n5666 2.6005
R5921 VSS.n5669 VSS.n5668 2.6005
R5922 VSS.n5672 VSS.n5671 2.6005
R5923 VSS.n5677 VSS.n5676 2.6005
R5924 VSS.n5663 VSS.n5662 2.6005
R5925 VSS.n5660 VSS.n5659 2.6005
R5926 VSS.n5658 VSS.n5657 2.6005
R5927 VSS.n5655 VSS.n5654 2.6005
R5928 VSS.n5653 VSS.n5652 2.6005
R5929 VSS.n5267 VSS.n5266 2.6005
R5930 VSS.n5269 VSS.n5268 2.6005
R5931 VSS.n5263 VSS.n5262 2.6005
R5932 VSS.n5261 VSS.n5260 2.6005
R5933 VSS.n5080 VSS.n5079 2.6005
R5934 VSS.n5082 VSS.n5081 2.6005
R5935 VSS.n5069 VSS.n5068 2.6005
R5936 VSS.n5085 VSS.n5084 2.6005
R5937 VSS.n5088 VSS.n5087 2.6005
R5938 VSS.n5091 VSS.n5090 2.6005
R5939 VSS.n5095 VSS.n5094 2.6005
R5940 VSS.n5114 VSS.n5113 2.6005
R5941 VSS.n5118 VSS.n5117 2.6005
R5942 VSS.n5120 VSS.n5119 2.6005
R5943 VSS.n5139 VSS.n5138 2.6005
R5944 VSS.n5142 VSS.n5141 2.6005
R5945 VSS.n5476 VSS.n5475 2.6005
R5946 VSS.n5145 VSS.n5144 2.6005
R5947 VSS.n5149 VSS.n5148 2.6005
R5948 VSS.n5148 VSS.n5147 2.6005
R5949 VSS.n5152 VSS.n5151 2.6005
R5950 VSS.n5151 VSS.n5150 2.6005
R5951 VSS.n5155 VSS.n5154 2.6005
R5952 VSS.n5154 VSS.n5153 2.6005
R5953 VSS.n5158 VSS.n5157 2.6005
R5954 VSS.n5157 VSS.n5156 2.6005
R5955 VSS.n5161 VSS.n5160 2.6005
R5956 VSS.n5160 VSS.n5159 2.6005
R5957 VSS.n5174 VSS.n5173 2.6005
R5958 VSS.n5173 VSS.n5172 2.6005
R5959 VSS.n5177 VSS.n5176 2.6005
R5960 VSS.n5176 VSS.n5175 2.6005
R5961 VSS.n5197 VSS.n5196 2.6005
R5962 VSS.n5196 VSS.n5195 2.6005
R5963 VSS.n5201 VSS.n5200 2.6005
R5964 VSS.n5200 VSS.n5199 2.6005
R5965 VSS.n5224 VSS.n5223 2.6005
R5966 VSS.n5223 VSS.n5222 2.6005
R5967 VSS.n5228 VSS.n5227 2.6005
R5968 VSS.n5227 VSS.n5226 2.6005
R5969 VSS.n5231 VSS.n5230 2.6005
R5970 VSS.n5230 VSS.n5229 2.6005
R5971 VSS.n5234 VSS.n5233 2.6005
R5972 VSS.n5233 VSS.n5232 2.6005
R5973 VSS.n4803 VSS.n4802 2.6005
R5974 VSS.n4802 VSS.n4801 2.6005
R5975 VSS.n5238 VSS.n5237 2.6005
R5976 VSS.n5237 VSS.n5236 2.6005
R5977 VSS.n5241 VSS.n5240 2.6005
R5978 VSS.n5240 VSS.n5239 2.6005
R5979 VSS.n5244 VSS.n5243 2.6005
R5980 VSS.n5243 VSS.n5242 2.6005
R5981 VSS.n5248 VSS.n5247 2.6005
R5982 VSS.n5247 VSS.n5246 2.6005
R5983 VSS.n4772 VSS.n4771 2.6005
R5984 VSS.n4771 VSS.n4770 2.6005
R5985 VSS.n4775 VSS.n4774 2.6005
R5986 VSS.n4774 VSS.n4773 2.6005
R5987 VSS.n5439 VSS.n5438 2.6005
R5988 VSS.n5438 VSS.n5437 2.6005
R5989 VSS.n5443 VSS.n5442 2.6005
R5990 VSS.n5442 VSS.n5441 2.6005
R5991 VSS.n5422 VSS.n5421 2.6005
R5992 VSS.n5447 VSS.n5446 2.6005
R5993 VSS.n5446 VSS.n5445 2.6005
R5994 VSS.n5450 VSS.n5449 2.6005
R5995 VSS.n5449 VSS.n5448 2.6005
R5996 VSS.n5453 VSS.n5452 2.6005
R5997 VSS.n5452 VSS.n5451 2.6005
R5998 VSS.n5456 VSS.n5455 2.6005
R5999 VSS.n5455 VSS.n5454 2.6005
R6000 VSS.n5459 VSS.n5458 2.6005
R6001 VSS.n5458 VSS.n5457 2.6005
R6002 VSS.n5420 VSS.n5419 2.6005
R6003 VSS.n5463 VSS.n5462 2.6005
R6004 VSS.n5462 VSS.n5461 2.6005
R6005 VSS.n5466 VSS.n5465 2.6005
R6006 VSS.n5465 VSS.n5464 2.6005
R6007 VSS.n5469 VSS.n5468 2.6005
R6008 VSS.n5468 VSS.n5467 2.6005
R6009 VSS.n5472 VSS.n5471 2.6005
R6010 VSS.n5471 VSS.n5470 2.6005
R6011 VSS.n5474 VSS.n5473 2.6005
R6012 VSS.n5554 VSS.n5553 2.6005
R6013 VSS.n5553 VSS.n5552 2.6005
R6014 VSS.n5551 VSS.n5550 2.6005
R6015 VSS.n5550 VSS.n5549 2.6005
R6016 VSS.n5543 VSS.n5542 2.6005
R6017 VSS.n5542 VSS.n5541 2.6005
R6018 VSS.n5540 VSS.n5539 2.6005
R6019 VSS.n5539 VSS.n5538 2.6005
R6020 VSS.n5537 VSS.n5536 2.6005
R6021 VSS.n5536 VSS.n5535 2.6005
R6022 VSS.n5534 VSS.n5533 2.6005
R6023 VSS.n5533 VSS.n5532 2.6005
R6024 VSS.n5480 VSS.n5479 2.6005
R6025 VSS.n5479 VSS.n5478 2.6005
R6026 VSS.n5495 VSS.n5494 2.6005
R6027 VSS.n5494 VSS.n5493 2.6005
R6028 VSS.n5498 VSS.n5497 2.6005
R6029 VSS.n5497 VSS.n5496 2.6005
R6030 VSS.n5501 VSS.n5500 2.6005
R6031 VSS.n5500 VSS.n5499 2.6005
R6032 VSS.n5504 VSS.n5503 2.6005
R6033 VSS.n5503 VSS.n5502 2.6005
R6034 VSS.n5507 VSS.n5506 2.6005
R6035 VSS.n5506 VSS.n5505 2.6005
R6036 VSS.n5510 VSS.n5509 2.6005
R6037 VSS.n5509 VSS.n5508 2.6005
R6038 VSS.n5513 VSS.n5512 2.6005
R6039 VSS.n5512 VSS.n5511 2.6005
R6040 VSS.n5516 VSS.n5515 2.6005
R6041 VSS.n5515 VSS.n5514 2.6005
R6042 VSS.n5519 VSS.n5518 2.6005
R6043 VSS.n5518 VSS.n5517 2.6005
R6044 VSS.n5522 VSS.n5521 2.6005
R6045 VSS.n5521 VSS.n5520 2.6005
R6046 VSS.n5525 VSS.n5524 2.6005
R6047 VSS.n5524 VSS.n5523 2.6005
R6048 VSS.n5528 VSS.n5527 2.6005
R6049 VSS.n5527 VSS.n5526 2.6005
R6050 VSS.n5492 VSS.n5491 2.6005
R6051 VSS.n5491 VSS.n5490 2.6005
R6052 VSS.n5616 VSS.n5615 2.6005
R6053 VSS.n5615 VSS.n5614 2.6005
R6054 VSS.n5613 VSS.n5612 2.6005
R6055 VSS.n5612 VSS.n5611 2.6005
R6056 VSS.n5610 VSS.n5609 2.6005
R6057 VSS.n5609 VSS.n5608 2.6005
R6058 VSS.n5606 VSS.n5605 2.6005
R6059 VSS.n5605 VSS.n5604 2.6005
R6060 VSS.n5603 VSS.n5602 2.6005
R6061 VSS.n5602 VSS.n5601 2.6005
R6062 VSS.n5600 VSS.n5599 2.6005
R6063 VSS.n5599 VSS.n5598 2.6005
R6064 VSS.n5597 VSS.n5596 2.6005
R6065 VSS.n5596 VSS.n5595 2.6005
R6066 VSS.n5594 VSS.n5593 2.6005
R6067 VSS.n5593 VSS.n5592 2.6005
R6068 VSS.n5590 VSS.n5589 2.6005
R6069 VSS.n5589 VSS.n5588 2.6005
R6070 VSS.n5586 VSS.n5585 2.6005
R6071 VSS.n5585 VSS.t150 2.6005
R6072 VSS.n5584 VSS.n5583 2.6005
R6073 VSS.n5583 VSS.n5582 2.6005
R6074 VSS.n5581 VSS.n5580 2.6005
R6075 VSS.n5580 VSS.n5579 2.6005
R6076 VSS.n5578 VSS.n5577 2.6005
R6077 VSS.n5577 VSS.n5576 2.6005
R6078 VSS.n5575 VSS.n5574 2.6005
R6079 VSS.n5574 VSS.n5573 2.6005
R6080 VSS.n5571 VSS.n5570 2.6005
R6081 VSS.n5570 VSS.n5569 2.6005
R6082 VSS.n5568 VSS.n5567 2.6005
R6083 VSS.n5567 VSS.n5566 2.6005
R6084 VSS.n5565 VSS.n5564 2.6005
R6085 VSS.n5564 VSS.n5563 2.6005
R6086 VSS.n5562 VSS.n5561 2.6005
R6087 VSS.n5561 VSS.n5560 2.6005
R6088 VSS.n5559 VSS.n5558 2.6005
R6089 VSS.n5558 VSS.n5557 2.6005
R6090 VSS.n5418 VSS.n5417 2.6005
R6091 VSS.n5417 VSS.n5416 2.6005
R6092 VSS.n5415 VSS.n5414 2.6005
R6093 VSS.n5414 VSS.n5413 2.6005
R6094 VSS.n5412 VSS.n5411 2.6005
R6095 VSS.n5411 VSS.n5410 2.6005
R6096 VSS.n5409 VSS.n5408 2.6005
R6097 VSS.n5408 VSS.n5407 2.6005
R6098 VSS.n5406 VSS.n5405 2.6005
R6099 VSS.n5405 VSS.n5404 2.6005
R6100 VSS.n5403 VSS.n5402 2.6005
R6101 VSS.n5402 VSS.n5401 2.6005
R6102 VSS.n5400 VSS.n5399 2.6005
R6103 VSS.n5399 VSS.n5398 2.6005
R6104 VSS.n5397 VSS.n5396 2.6005
R6105 VSS.n5396 VSS.n5395 2.6005
R6106 VSS.n5394 VSS.n5393 2.6005
R6107 VSS.n5393 VSS.n5392 2.6005
R6108 VSS.n5391 VSS.n5390 2.6005
R6109 VSS.n5390 VSS.n5389 2.6005
R6110 VSS.n5388 VSS.n5387 2.6005
R6111 VSS.n5387 VSS.n5386 2.6005
R6112 VSS.n5385 VSS.n5384 2.6005
R6113 VSS.n5384 VSS.n5383 2.6005
R6114 VSS.n5382 VSS.n5381 2.6005
R6115 VSS.n5381 VSS.n5380 2.6005
R6116 VSS.n5379 VSS.n5378 2.6005
R6117 VSS.n5378 VSS.n5377 2.6005
R6118 VSS.n5376 VSS.n5375 2.6005
R6119 VSS.n5375 VSS.n5374 2.6005
R6120 VSS.n5373 VSS.n5372 2.6005
R6121 VSS.n5372 VSS.n5371 2.6005
R6122 VSS.n5370 VSS.n5369 2.6005
R6123 VSS.n5369 VSS.n5368 2.6005
R6124 VSS.n5367 VSS.n5366 2.6005
R6125 VSS.n5366 VSS.n5365 2.6005
R6126 VSS.n5364 VSS.n5363 2.6005
R6127 VSS.n5363 VSS.n5362 2.6005
R6128 VSS.n5361 VSS.n5360 2.6005
R6129 VSS.n5360 VSS.n5359 2.6005
R6130 VSS.n5358 VSS.n5357 2.6005
R6131 VSS.n5357 VSS.n5356 2.6005
R6132 VSS.n5680 VSS.n5679 2.6005
R6133 VSS.n5679 VSS.n5678 2.6005
R6134 VSS.n5687 VSS.n5686 2.6005
R6135 VSS.n5686 VSS.n5685 2.6005
R6136 VSS.n5690 VSS.n5689 2.6005
R6137 VSS.n5689 VSS.n5688 2.6005
R6138 VSS.n5693 VSS.n5692 2.6005
R6139 VSS.n5692 VSS.n5691 2.6005
R6140 VSS.n5696 VSS.n5695 2.6005
R6141 VSS.n5695 VSS.n5694 2.6005
R6142 VSS.n5699 VSS.n5698 2.6005
R6143 VSS.n5698 VSS.n5697 2.6005
R6144 VSS.n5702 VSS.n5701 2.6005
R6145 VSS.n5701 VSS.n5700 2.6005
R6146 VSS.n5705 VSS.n5704 2.6005
R6147 VSS.n5704 VSS.n5703 2.6005
R6148 VSS.n5708 VSS.n5707 2.6005
R6149 VSS.n5707 VSS.n5706 2.6005
R6150 VSS.n5712 VSS.n5711 2.6005
R6151 VSS.n5711 VSS.n5710 2.6005
R6152 VSS.n5715 VSS.n5714 2.6005
R6153 VSS.n5714 VSS.n5713 2.6005
R6154 VSS.n5718 VSS.n5717 2.6005
R6155 VSS.n5717 VSS.n5716 2.6005
R6156 VSS.n5721 VSS.n5720 2.6005
R6157 VSS.n5720 VSS.n5719 2.6005
R6158 VSS.n5724 VSS.n5723 2.6005
R6159 VSS.n5723 VSS.n5722 2.6005
R6160 VSS.n5727 VSS.n5726 2.6005
R6161 VSS.n5726 VSS.n5725 2.6005
R6162 VSS.n5730 VSS.n5729 2.6005
R6163 VSS.n5729 VSS.n5728 2.6005
R6164 VSS.n5732 VSS.n5731 2.6005
R6165 VSS.n5733 VSS.n5732 2.6005
R6166 VSS.n5941 VSS.n5940 2.6005
R6167 VSS.n5940 VSS.n5939 2.6005
R6168 VSS.n5944 VSS.n5943 2.6005
R6169 VSS.n5943 VSS.n5942 2.6005
R6170 VSS.n5947 VSS.n5946 2.6005
R6171 VSS.n5946 VSS.n5945 2.6005
R6172 VSS.n5950 VSS.n5949 2.6005
R6173 VSS.n5949 VSS.n5948 2.6005
R6174 VSS.n5953 VSS.n5952 2.6005
R6175 VSS.n5952 VSS.n5951 2.6005
R6176 VSS.n5956 VSS.n5955 2.6005
R6177 VSS.n5955 VSS.n5954 2.6005
R6178 VSS.n5959 VSS.n5958 2.6005
R6179 VSS.n5958 VSS.n5957 2.6005
R6180 VSS.n5962 VSS.n5961 2.6005
R6181 VSS.n5961 VSS.n5960 2.6005
R6182 VSS.n5965 VSS.n5964 2.6005
R6183 VSS.n5964 VSS.n5963 2.6005
R6184 VSS.n5968 VSS.n5967 2.6005
R6185 VSS.n5967 VSS.n5966 2.6005
R6186 VSS.n5971 VSS.n5970 2.6005
R6187 VSS.n5970 VSS.n5969 2.6005
R6188 VSS.n5974 VSS.n5973 2.6005
R6189 VSS.n5973 VSS.n5972 2.6005
R6190 VSS.n5977 VSS.n5976 2.6005
R6191 VSS.n5976 VSS.n5975 2.6005
R6192 VSS.n5980 VSS.n5979 2.6005
R6193 VSS.n5979 VSS.n5978 2.6005
R6194 VSS.n5983 VSS.n5982 2.6005
R6195 VSS.n5982 VSS.n5981 2.6005
R6196 VSS.n5987 VSS.n5986 2.6005
R6197 VSS.n5986 VSS.n5985 2.6005
R6198 VSS.n5991 VSS.n5990 2.6005
R6199 VSS.n5990 VSS.n5989 2.6005
R6200 VSS.n4769 VSS.n4768 2.6005
R6201 VSS.n4766 VSS.n4765 2.6005
R6202 VSS.n4741 VSS.n4740 2.6005
R6203 VSS.n5938 VSS.n5937 2.6005
R6204 VSS VSS.n5846 2.6005
R6205 VSS.n5846 VSS.t96 2.6005
R6206 VSS.n5781 VSS 2.6005
R6207 VSS.n5781 VSS.n5780 2.6005
R6208 VSS.n1019 VSS.n1018 2.6005
R6209 VSS.n1022 VSS.n1021 2.6005
R6210 VSS.n1016 VSS.n1015 2.6005
R6211 VSS.n4055 VSS.n4054 2.59998
R6212 VSS.n1566 VSS.n1565 2.53192
R6213 VSS.n1261 VSS.n1260 2.48961
R6214 VSS.n1264 VSS.n1263 2.48961
R6215 VSS.n1267 VSS.n1266 2.48961
R6216 VSS.n1270 VSS.n1269 2.48961
R6217 VSS.n1273 VSS.n1272 2.48961
R6218 VSS.n1276 VSS.n1275 2.48961
R6219 VSS.n1279 VSS.n1278 2.48961
R6220 VSS.n471 VSS.n470 2.41686
R6221 VSS.n5828 VSS.n5827 2.36862
R6222 VSS.n1646 VSS.n1554 2.3405
R6223 VSS.n1647 VSS.n1544 2.33208
R6224 VSS.n1566 VSS.n1561 2.33079
R6225 VSS.n5807 VSS.n21 2.30179
R6226 VSS.n987 VSS.n986 2.29396
R6227 VSS.n5827 VSS.n5826 2.29248
R6228 VSS.n2802 VSS.n2801 2.28632
R6229 VSS.n5345 VSS.n5344 2.28399
R6230 VSS.n5348 VSS.n5347 2.28399
R6231 VSS.n558 VSS.n557 2.28399
R6232 VSS.n561 VSS.n560 2.28399
R6233 VSS.n677 VSS.n676 2.28399
R6234 VSS.n680 VSS.n679 2.28399
R6235 VSS.n6016 VSS.n6015 2.28399
R6236 VSS.n6029 VSS.n6028 2.28399
R6237 VSS.n6032 VSS.n6031 2.28399
R6238 VSS.n6035 VSS.n6034 2.28399
R6239 VSS.n6047 VSS.n6046 2.28399
R6240 VSS.n6050 VSS.n6049 2.28399
R6241 VSS.n6053 VSS.n6052 2.28399
R6242 VSS.n6056 VSS.n6055 2.28399
R6243 VSS.n5671 VSS.n5670 2.28399
R6244 VSS.n5643 VSS.n5642 2.28399
R6245 VSS.n5631 VSS.n5630 2.28399
R6246 VSS.n5628 VSS.n5627 2.28399
R6247 VSS.n4740 VSS.n4739 2.28399
R6248 VSS.n5911 VSS 2.28174
R6249 VSS.n2722 VSS.n2212 2.2791
R6250 VSS.n2580 VSS.n2579 2.27836
R6251 VSS.n2193 VSS.n2192 2.27834
R6252 VSS.n2879 VSS.n1995 2.27413
R6253 VSS.n2789 VSS.n2094 2.27187
R6254 VSS.n2656 VSS.n2320 2.26934
R6255 VSS.n2663 VSS.n2308 2.25712
R6256 VSS.n4371 VSS.n4370 2.25676
R6257 VSS.n5292 VSS.n5291 2.25635
R6258 VSS.n2560 VSS.n2413 2.25613
R6259 VSS.n874 VSS.n870 2.25575
R6260 VSS.n1754 VSS.t341 2.25428
R6261 VSS.n1755 VSS.t321 2.25428
R6262 VSS.n1756 VSS.t393 2.25428
R6263 VSS.n1757 VSS.t402 2.25428
R6264 VSS.n1758 VSS.t319 2.25428
R6265 VSS.n1759 VSS.t328 2.25428
R6266 VSS.n1760 VSS.t306 2.25428
R6267 VSS.n1761 VSS.t386 2.25428
R6268 VSS.n1762 VSS.t389 2.25428
R6269 VSS.n1763 VSS.t367 2.25428
R6270 VSS.n1764 VSS.t312 2.25428
R6271 VSS.n2458 VSS.t396 2.25428
R6272 VSS.n2459 VSS.t378 2.25428
R6273 VSS.n2460 VSS.t314 2.25428
R6274 VSS.n2461 VSS.t323 2.25428
R6275 VSS.n2462 VSS.t374 2.25428
R6276 VSS.n2463 VSS.t385 2.25428
R6277 VSS.n2464 VSS.t359 2.25428
R6278 VSS.n2465 VSS.t305 2.25428
R6279 VSS.n2466 VSS.t308 2.25428
R6280 VSS.n2467 VSS.t412 2.25428
R6281 VSS.n2468 VSS.t366 2.25428
R6282 VSS.n2372 VSS.t317 2.25428
R6283 VSS.n2373 VSS.t294 2.25428
R6284 VSS.n2374 VSS.t371 2.25428
R6285 VSS.n2375 VSS.t383 2.25428
R6286 VSS.n2376 VSS.t291 2.25428
R6287 VSS.n2377 VSS.t300 2.25428
R6288 VSS.n2378 VSS.t407 2.25428
R6289 VSS.n2379 VSS.t361 2.25428
R6290 VSS.n2380 VSS.t363 2.25428
R6291 VSS.n2381 VSS.t338 2.25428
R6292 VSS.n2382 VSS.t284 2.25428
R6293 VSS.n2255 VSS.t349 2.25428
R6294 VSS.n2256 VSS.t327 2.25428
R6295 VSS.n2257 VSS.t401 2.25428
R6296 VSS.n2258 VSS.t405 2.25428
R6297 VSS.n2259 VSS.t325 2.25428
R6298 VSS.n2260 VSS.t332 2.25428
R6299 VSS.n2261 VSS.t311 2.25428
R6300 VSS.n2262 VSS.t391 2.25428
R6301 VSS.n2263 VSS.t392 2.25428
R6302 VSS.n2264 VSS.t375 2.25428
R6303 VSS.n2265 VSS.t318 2.25428
R6304 VSS.n2148 VSS.t301 2.25428
R6305 VSS.n2149 VSS.t408 2.25428
R6306 VSS.n2150 VSS.t357 2.25428
R6307 VSS.n2151 VSS.t364 2.25428
R6308 VSS.n2152 VSS.t406 2.25428
R6309 VSS.n2153 VSS.t285 2.25428
R6310 VSS.n2154 VSS.t398 2.25428
R6311 VSS.n2155 VSS.t344 2.25428
R6312 VSS.n2156 VSS.t346 2.25428
R6313 VSS.n2157 VSS.t324 2.25428
R6314 VSS.n2158 VSS.t404 2.25428
R6315 VSS.n2051 VSS.t381 2.25428
R6316 VSS.n2052 VSS.t356 2.25428
R6317 VSS.n2053 VSS.t293 2.25428
R6318 VSS.n2054 VSS.t302 2.25428
R6319 VSS.n2055 VSS.t353 2.25428
R6320 VSS.n2056 VSS.t362 2.25428
R6321 VSS.n2057 VSS.t337 2.25428
R6322 VSS.n2058 VSS.t414 2.25428
R6323 VSS.n2059 VSS.t286 2.25428
R6324 VSS.n2060 VSS.t400 2.25428
R6325 VSS.n2061 VSS.t345 2.25428
R6326 VSS.n1981 VSS.t379 2.25428
R6327 VSS.n1982 VSS.t354 2.25428
R6328 VSS.n1983 VSS.t290 2.25428
R6329 VSS.n1984 VSS.t298 2.25428
R6330 VSS.n1985 VSS.t350 2.25428
R6331 VSS.n1986 VSS.t360 2.25428
R6332 VSS.n1987 VSS.t335 2.25428
R6333 VSS.n1988 VSS.t411 2.25428
R6334 VSS.n1989 VSS.t415 2.25428
R6335 VSS.n1990 VSS.t397 2.25428
R6336 VSS.n1991 VSS.t342 2.25428
R6337 VSS.n1826 VSS.t377 2.25428
R6338 VSS.n1827 VSS.t352 2.25428
R6339 VSS.n1828 VSS.t289 2.25428
R6340 VSS.n1829 VSS.t297 2.25428
R6341 VSS.n1830 VSS.t347 2.25428
R6342 VSS.n1831 VSS.t358 2.25428
R6343 VSS.n1832 VSS.t334 2.25428
R6344 VSS.n1833 VSS.t410 2.25428
R6345 VSS.n1834 VSS.t413 2.25428
R6346 VSS.n1835 VSS.t394 2.25428
R6347 VSS.n1836 VSS.t340 2.25428
R6348 VSS.n1792 VSS.t329 2.25428
R6349 VSS.n1793 VSS.t307 2.25428
R6350 VSS.n1794 VSS.t384 2.25428
R6351 VSS.n1795 VSS.t390 2.25428
R6352 VSS.n1796 VSS.t303 2.25428
R6353 VSS.n1797 VSS.t313 2.25428
R6354 VSS.n1798 VSS.t288 2.25428
R6355 VSS.n1799 VSS.t372 2.25428
R6356 VSS.n1800 VSS.t376 2.25428
R6357 VSS.n1801 VSS.t351 2.25428
R6358 VSS.n1802 VSS.t296 2.25428
R6359 VSS.n1771 VSS.t326 2.25428
R6360 VSS.n1772 VSS.t304 2.25428
R6361 VSS.n1773 VSS.t382 2.25428
R6362 VSS.n1774 VSS.t388 2.25428
R6363 VSS.n1775 VSS.t299 2.25428
R6364 VSS.n1776 VSS.t310 2.25428
R6365 VSS.n1777 VSS.t287 2.25428
R6366 VSS.n1778 VSS.t370 2.25428
R6367 VSS.n1779 VSS.t373 2.25428
R6368 VSS.n1780 VSS.t348 2.25428
R6369 VSS.n1781 VSS.t295 2.25428
R6370 VSS.n1743 VSS.t355 2.25428
R6371 VSS.n1744 VSS.t331 2.25428
R6372 VSS.n1745 VSS.t403 2.25428
R6373 VSS.n1746 VSS.t409 2.25428
R6374 VSS.n1747 VSS.t330 2.25428
R6375 VSS.n1748 VSS.t336 2.25428
R6376 VSS.n1749 VSS.t315 2.25428
R6377 VSS.n1750 VSS.t395 2.25428
R6378 VSS.n1751 VSS.t399 2.25428
R6379 VSS.n1752 VSS.t380 2.25428
R6380 VSS.n1753 VSS.t322 2.25428
R6381 VSS.n1719 VSS.t712 2.25416
R6382 VSS.n1728 VSS.t711 2.25416
R6383 VSS.n1720 VSS.t709 2.25416
R6384 VSS.n1662 VSS.n1661 2.2531
R6385 VSS.n1669 VSS.n1665 2.2531
R6386 VSS.n3907 VSS.n3906 2.25293
R6387 VSS.n1402 VSS.n1401 2.25285
R6388 VSS.n1656 VSS.n1654 2.25253
R6389 VSS.n2491 VSS.n2478 2.25113
R6390 VSS.n1686 VSS.n1685 2.25077
R6391 VSS.n319 VSS.n318 2.2505
R6392 VSS.n1455 VSS.n1454 2.2505
R6393 VSS.n1513 VSS.n1512 2.2505
R6394 VSS.n3995 VSS.n3990 2.2505
R6395 VSS.n1502 VSS.n1501 2.2505
R6396 VSS.n337 VSS.n336 2.2505
R6397 VSS.n357 VSS.n356 2.2505
R6398 VSS.n1645 VSS.n1644 2.2505
R6399 VSS.n1579 VSS.n1578 2.2505
R6400 VSS.n1571 VSS.n1570 2.2505
R6401 VSS.n1569 VSS.n1568 2.2505
R6402 VSS.n1577 VSS.n1576 2.2505
R6403 VSS.n3397 VSS.n3369 2.2505
R6404 VSS.n3388 VSS.n3372 2.2505
R6405 VSS.n3403 VSS.n3367 2.2505
R6406 VSS.n3396 VSS.n3370 2.2505
R6407 VSS.n3386 VSS.n3373 2.2505
R6408 VSS.n3398 VSS.n3368 2.2505
R6409 VSS.n3379 VSS.n3375 2.2505
R6410 VSS.n3382 VSS.n3374 2.2505
R6411 VSS.n3390 VSS.n3371 2.2505
R6412 VSS.n3078 VSS.n3077 2.2505
R6413 VSS.n3229 VSS.n3206 2.2505
R6414 VSS.n3074 VSS.n3073 2.2505
R6415 VSS.n3082 VSS.n3081 2.2505
R6416 VSS.n3213 VSS.n3212 2.2505
R6417 VSS.n3224 VSS.n3223 2.2505
R6418 VSS.n3219 VSS.n3208 2.2505
R6419 VSS.n3225 VSS.n3207 2.2505
R6420 VSS.n3216 VSS.n3209 2.2505
R6421 VSS.n2923 VSS.n2922 2.2505
R6422 VSS.n2952 VSS.n2951 2.2505
R6423 VSS.n2938 VSS.n2937 2.2505
R6424 VSS.n2927 VSS.n2926 2.2505
R6425 VSS.n2948 VSS.n2947 2.2505
R6426 VSS.n2942 VSS.n2941 2.2505
R6427 VSS.n2931 VSS.n2930 2.2505
R6428 VSS.n2950 VSS.n2949 2.2505
R6429 VSS.n2936 VSS.n2935 2.2505
R6430 VSS.n1858 VSS.n1857 2.2505
R6431 VSS.n1847 VSS.n1843 2.2505
R6432 VSS.n1854 VSS.n1840 2.2505
R6433 VSS.n1870 VSS.n1837 2.2505
R6434 VSS.n1859 VSS.n1839 2.2505
R6435 VSS.n1849 VSS.n1841 2.2505
R6436 VSS.n1864 VSS.n1863 2.2505
R6437 VSS.n1848 VSS.n1842 2.2505
R6438 VSS.n1867 VSS.n1838 2.2505
R6439 VSS.n2798 VSS.n2797 2.2505
R6440 VSS.n2017 VSS.n1995 2.2505
R6441 VSS.n2801 VSS.n2080 2.2505
R6442 VSS.n2024 VSS.n2022 2.2505
R6443 VSS.n2021 VSS.n2020 2.2505
R6444 VSS.n2844 VSS.n2843 2.2505
R6445 VSS.n2796 VSS.n2047 2.2505
R6446 VSS.n2856 VSS.n2855 2.2505
R6447 VSS.n2800 VSS.n2799 2.2505
R6448 VSS.n2854 VSS.n2853 2.2505
R6449 VSS.n2130 VSS.n2108 2.2505
R6450 VSS.n2192 VSS.n2191 2.2505
R6451 VSS.n2753 VSS.n2143 2.2505
R6452 VSS.n2137 VSS.n2131 2.2505
R6453 VSS.n2190 VSS.n2177 2.2505
R6454 VSS.n2189 VSS.n2179 2.2505
R6455 VSS.n2141 VSS.n2140 2.2505
R6456 VSS.n2755 VSS.n2754 2.2505
R6457 VSS.n2142 VSS.n2127 2.2505
R6458 VSS.n2102 VSS.n2094 2.2505
R6459 VSS.n2293 VSS.n2235 2.2505
R6460 VSS.n2292 VSS.n2234 2.2505
R6461 VSS.n2308 VSS.n2277 2.2505
R6462 VSS.n2307 VSS.n2306 2.2505
R6463 VSS.n2297 VSS.n2284 2.2505
R6464 VSS.n2296 VSS.n2295 2.2505
R6465 VSS.n2230 VSS.n2212 2.2505
R6466 VSS.n2294 VSS.n2247 2.2505
R6467 VSS.n2571 VSS.n2361 2.2505
R6468 VSS.n2579 VSS.n2578 2.2505
R6469 VSS.n2570 VSS.n2360 2.2505
R6470 VSS.n2331 VSS.n2320 2.2505
R6471 VSS.n2575 VSS.n2574 2.2505
R6472 VSS.n2577 VSS.n2568 2.2505
R6473 VSS.n2573 VSS.n2572 2.2505
R6474 VSS.n2569 VSS.n2346 2.2505
R6475 VSS.n2640 VSS.n2332 2.2505
R6476 VSS.n2368 VSS.n2362 2.2505
R6477 VSS.n2485 VSS.n2451 2.2505
R6478 VSS.n2484 VSS.n2440 2.2505
R6479 VSS.n2486 VSS.n2474 2.2505
R6480 VSS.n2546 VSS.n2545 2.2505
R6481 VSS.n2530 VSS.n2439 2.2505
R6482 VSS.n2543 VSS.n2542 2.2505
R6483 VSS.n2426 VSS.n2413 2.2505
R6484 VSS.n2541 VSS.n2540 2.2505
R6485 VSS.n2548 VSS.n2547 2.2505
R6486 VSS.n2549 VSS.n2421 2.2505
R6487 VSS.n2539 VSS.n2538 2.2505
R6488 VSS.n3908 VSS.n3907 2.2505
R6489 VSS.n1673 VSS.n1672 2.2505
R6490 VSS.n1687 VSS.n1686 2.2505
R6491 VSS.n4162 VSS.n4161 2.2505
R6492 VSS.n4174 VSS.n4173 2.2505
R6493 VSS.n5794 VSS.n5793 2.2505
R6494 VSS.n5791 VSS.n5790 2.2505
R6495 VSS.n3845 VSS.n1727 2.24994
R6496 VSS.n1678 VSS.n1677 2.24918
R6497 VSS.n972 VSS.n971 2.24654
R6498 VSS.n912 VSS.n911 2.24654
R6499 VSS.n3844 VSS.n3843 2.24495
R6500 VSS.n1662 VSS.n1660 2.24449
R6501 VSS.n1656 VSS.n1655 2.24449
R6502 VSS.n1669 VSS.n1668 2.24449
R6503 VSS.n3907 VSS.n1690 2.24449
R6504 VSS.n469 VSS.n468 2.22001
R6505 VSS.n295 VSS.n293 2.04928
R6506 VSS.n910 VSS.t492 2.02838
R6507 VSS.n1393 VSS.t111 2.02837
R6508 VSS.n324 VSS.t649 2.02837
R6509 VSS.t234 VSS.t270 2.02605
R6510 VSS.t218 VSS.t234 2.02605
R6511 VSS.n5226 VSS.t158 2.02605
R6512 VSS.n4209 VSS.n4208 2.0097
R6513 VSS.n970 VSS.n969 2.00969
R6514 VSS.n280 VSS.n279 2.00969
R6515 VSS.n293 VSS.n278 1.96391
R6516 VSS VSS.n4738 1.9362
R6517 VSS.t416 VSS.t468 1.92472
R6518 VSS.t420 VSS.t471 1.92472
R6519 VSS.t417 VSS.t475 1.92472
R6520 VSS.t705 VSS.t101 1.92472
R6521 VSS.t702 VSS.t103 1.92472
R6522 VSS.t138 VSS.t139 1.92472
R6523 VSS.t699 VSS.t138 1.92472
R6524 VSS.t137 VSS.t140 1.92472
R6525 VSS.t701 VSS.t137 1.92472
R6526 VSS.t8 VSS.t5 1.92244
R6527 VSS.t14 VSS.t11 1.92244
R6528 VSS.t696 VSS.t2 1.92244
R6529 VSS.n4469 VSS.n4468 1.90368
R6530 VSS.n1318 VSS.n1317 1.87586
R6531 VSS.n4221 VSS.n4220 1.87586
R6532 VSS.n224 VSS.n223 1.85787
R6533 VSS.n126 VSS.n125 1.85767
R6534 VSS.n5213 VSS.n5212 1.85765
R6535 VSS.n4793 VSS.n4792 1.85765
R6536 VSS.n5877 VSS.n5876 1.85285
R6537 VSS.n250 VSS.n249 1.83785
R6538 VSS.n4388 VSS.n4387 1.83785
R6539 VSS.n4563 VSS.n4562 1.83785
R6540 VSS.n4394 VSS.n4393 1.83724
R6541 VSS.n5278 VSS.n5277 1.83716
R6542 VSS.n50 VSS.n49 1.83716
R6543 VSS.n4417 VSS.n4416 1.83716
R6544 VSS.n5328 VSS.n5327 1.83716
R6545 VSS.n5306 VSS.n5305 1.83716
R6546 VSS.n4781 VSS.n4780 1.83716
R6547 VSS.n5266 VSS.n5265 1.83716
R6548 VSS.n5068 VSS.n5067 1.83716
R6549 VSS.n5087 VSS.n5086 1.83716
R6550 VSS.n5094 VSS.n5093 1.83716
R6551 VSS.n5117 VSS.n5116 1.83716
R6552 VSS.n5138 VSS.n5137 1.83716
R6553 VSS.n884 VSS.n883 1.82536
R6554 VSS.n970 VSS.t66 1.82525
R6555 VSS.n280 VSS.t497 1.82525
R6556 VSS.n4209 VSS.t656 1.82525
R6557 VSS.n1507 VSS.n1506 1.82479
R6558 VSS.n5827 VSS.n5809 1.80764
R6559 VSS.n1393 VSS.n1392 1.80405
R6560 VSS.n324 VSS.n323 1.80405
R6561 VSS.n910 VSS.n909 1.80404
R6562 VSS.n503 VSS.n500 1.8001
R6563 VSS.n4308 VSS.n4301 1.8001
R6564 VSS.n3913 VSS.n3910 1.8001
R6565 VSS.n4045 VSS.n4044 1.8001
R6566 VSS.n365 VSS.n364 1.8001
R6567 VSS.n490 VSS.n489 1.79951
R6568 VSS.n503 VSS.n502 1.79951
R6569 VSS.n4308 VSS.n4307 1.79951
R6570 VSS.n4274 VSS.n4271 1.79951
R6571 VSS.n3913 VSS.n3912 1.79951
R6572 VSS.n4108 VSS.n4104 1.79951
R6573 VSS.n4282 VSS.n4281 1.79942
R6574 VSS.n901 VSS.n900 1.79942
R6575 VSS.n469 VSS.n466 1.79318
R6576 VSS.n4025 VSS.n4022 1.7505
R6577 VSS.n119 VSS.n118 1.7445
R6578 VSS.n1329 VSS.n1328 1.68421
R6579 VSS.n1335 VSS.n1334 1.68421
R6580 VSS.n4116 VSS.n4114 1.68421
R6581 VSS.n1349 VSS.n1348 1.68411
R6582 VSS.n1354 VSS.n1353 1.68411
R6583 VSS.n1359 VSS.n1358 1.68411
R6584 VSS.n1364 VSS.n1363 1.68411
R6585 VSS.n1370 VSS.n1369 1.68411
R6586 VSS.n1287 VSS.n1286 1.68411
R6587 VSS.n928 VSS.n927 1.65879
R6588 VSS.n934 VSS.n933 1.65879
R6589 VSS.n944 VSS.n943 1.65879
R6590 VSS.n935 VSS.n934 1.65822
R6591 VSS.n941 VSS.n940 1.65822
R6592 VSS.n4142 VSS.n4141 1.65811
R6593 VSS.n834 VSS.n830 1.65328
R6594 VSS.n342 VSS.n341 1.62245
R6595 VSS.n4998 VSS.n4997 1.60209
R6596 VSS.n4596 VSS.n4595 1.60209
R6597 VSS.n4577 VSS.n4576 1.60209
R6598 VSS.n4668 VSS.n4667 1.60209
R6599 VSS.n4566 VSS.n4565 1.60209
R6600 VSS.n5302 VSS.n5301 1.60209
R6601 VSS.n5425 VSS.n5424 1.60199
R6602 VSS.n4979 VSS.n4978 1.60199
R6603 VSS.n37 VSS.n36 1.60199
R6604 VSS.n43 VSS.n42 1.60199
R6605 VSS.n53 VSS.n52 1.60199
R6606 VSS.n4672 VSS.n4671 1.60199
R6607 VSS.n4659 VSS.n4658 1.60199
R6608 VSS.n4574 VSS.n4573 1.60199
R6609 VSS.n4593 VSS.n4592 1.60199
R6610 VSS.n4604 VSS.n4603 1.60199
R6611 VSS.n4426 VSS.n4425 1.60199
R6612 VSS.n4421 VSS.n4420 1.60199
R6613 VSS.n510 VSS.n506 1.59295
R6614 VSS.n4318 VSS.n4317 1.59295
R6615 VSS.n510 VSS.n509 1.5924
R6616 VSS.n4339 VSS.n4338 1.59228
R6617 VSS.n4323 VSS.n4322 1.59228
R6618 VSS.n4353 VSS.n4352 1.59228
R6619 VSS.n690 VSS.n689 1.58814
R6620 VSS.n597 VSS.n596 1.58759
R6621 VSS.n5652 VSS.n5651 1.58759
R6622 VSS.n6008 VSS.n6007 1.58747
R6623 VSS.n6002 VSS.n6001 1.58747
R6624 VSS.n5997 VSS.n5996 1.58747
R6625 VSS.n5662 VSS.n5661 1.58747
R6626 VSS.n5657 VSS.n5656 1.58747
R6627 VSS.n262 VSS.n259 1.56241
R6628 VSS.n4231 VSS.n4230 1.55933
R6629 VSS.n904 VSS.n903 1.55922
R6630 VSS.n4240 VSS.n4239 1.55922
R6631 VSS.n1466 VSS.n1464 1.55606
R6632 VSS.n1648 VSS.n1647 1.50717
R6633 VSS.n1647 VSS.n1646 1.50266
R6634 VSS.n3906 VSS.n3905 1.5016
R6635 VSS.n299 VSS.n297 1.5005
R6636 VSS.n1552 VSS.n1551 1.5005
R6637 VSS.n3897 VSS.n3896 1.5005
R6638 VSS.n3902 VSS.n3901 1.5005
R6639 VSS.n1726 VSS.n1725 1.5005
R6640 VSS.n3838 VSS.n3837 1.5005
R6641 VSS.n3752 VSS.n3751 1.5005
R6642 VSS.n3805 VSS.n3804 1.5005
R6643 VSS.n3825 VSS.n3824 1.5005
R6644 VSS.n3769 VSS.n3768 1.5005
R6645 VSS.n3789 VSS.n3788 1.5005
R6646 VSS.n1542 VSS.n1541 1.5005
R6647 VSS.n5771 VSS.t684 1.463
R6648 VSS.n5771 VSS.n5770 1.463
R6649 VSS.n5918 VSS.t688 1.463
R6650 VSS.n5918 VSS.n5917 1.463
R6651 VSS.n5924 VSS.t56 1.463
R6652 VSS.n5924 VSS.n5923 1.463
R6653 VSS.n5901 VSS.t614 1.463
R6654 VSS.n5901 VSS.n5900 1.463
R6655 VSS.n5883 VSS.t22 1.463
R6656 VSS.n5883 VSS.n5882 1.463
R6657 VSS.n5909 VSS.t734 1.463
R6658 VSS.n5909 VSS.n5908 1.463
R6659 VSS.n5907 VSS.t268 1.463
R6660 VSS.n5907 VSS.n5906 1.463
R6661 VSS.n5928 VSS.t725 1.463
R6662 VSS.n5928 VSS.n5927 1.463
R6663 VSS.n4748 VSS.t595 1.463
R6664 VSS.n4748 VSS.n4747 1.463
R6665 VSS.n5786 VSS.t763 1.463
R6666 VSS.n5786 VSS.n5785 1.463
R6667 VSS.n5842 VSS.t29 1.463
R6668 VSS.n5842 VSS.n5841 1.463
R6669 VSS.n5773 VSS.t747 1.463
R6670 VSS.n5773 VSS.n5772 1.463
R6671 VSS.n5776 VSS.t666 1.463
R6672 VSS.n5776 VSS.n5775 1.463
R6673 VSS.n5778 VSS.t97 1.463
R6674 VSS.n5778 VSS.n5777 1.463
R6675 VSS.n5797 VSS.t1 1.463
R6676 VSS.n5797 VSS.n5796 1.463
R6677 VSS.n5831 VSS.t575 1.463
R6678 VSS.n5831 VSS.n5830 1.463
R6679 VSS.n5674 VSS.n5673 1.4595
R6680 VSS.n4689 VSS.n4687 1.45883
R6681 VSS.n1520 VSS.n1516 1.45883
R6682 VSS.n5547 VSS.n5546 1.43813
R6683 VSS.n1256 VSS.n1255 1.43195
R6684 VSS.n1170 VSS.n1169 1.43182
R6685 VSS.n1344 VSS.n1343 1.43182
R6686 VSS.n1282 VSS.n1281 1.43182
R6687 VSS.n1306 VSS.n1305 1.43182
R6688 VSS.n1300 VSS.n1299 1.43182
R6689 VSS.n4193 VSS.n4192 1.36161
R6690 VSS.n979 VSS.n978 1.33389
R6691 VSS.n991 VSS.n990 1.33389
R6692 VSS.n982 VSS.n981 1.33375
R6693 VSS.n98 VSS.n97 1.33375
R6694 VSS.n4348 VSS.n4347 1.33375
R6695 VSS.n4342 VSS.n4341 1.33375
R6696 VSS.n4333 VSS.n4332 1.33375
R6697 VSS.n4326 VSS.n4325 1.33375
R6698 VSS.n5340 VSS.n5339 1.32883
R6699 VSS.n565 VSS.n564 1.32883
R6700 VSS.n684 VSS.n683 1.32883
R6701 VSS.n6021 VSS.n6020 1.32883
R6702 VSS.n6039 VSS.n6038 1.32883
R6703 VSS.n6060 VSS.n6059 1.32883
R6704 VSS.n5676 VSS.n5675 1.32883
R6705 VSS.n5646 VSS.n5645 1.32883
R6706 VSS.n5635 VSS.n5634 1.32883
R6707 VSS.n1017 VSS.n1016 1.32883
R6708 VSS.n672 VSS.n671 1.32869
R6709 VSS.n553 VSS.n552 1.32869
R6710 VSS.n5352 VSS.n5351 1.32869
R6711 VSS.n4768 VSS.n4767 1.32869
R6712 VSS.n5666 VSS.n5665 1.32869
R6713 VSS.n5638 VSS.n5637 1.32869
R6714 VSS.n5621 VSS.n5620 1.32869
R6715 VSS.n1020 VSS.n1019 1.32869
R6716 VSS.n6042 VSS.n6041 1.32869
R6717 VSS.n6024 VSS.n6023 1.32869
R6718 VSS.n6011 VSS.n6010 1.32869
R6719 VSS.n5317 VSS.n5316 1.27022
R6720 VSS.n4405 VSS.n4404 1.26985
R6721 VSS.n1023 VSS.n1022 1.26929
R6722 VSS.n1000 VSS.n999 1.26929
R6723 VSS.n18 VSS.n17 1.26929
R6724 VSS.n6094 VSS.n6093 1.26929
R6725 VSS.n4158 VSS.n4149 1.26439
R6726 VSS.n4179 VSS.n4176 1.26439
R6727 VSS.n4983 VSS.n4963 1.22037
R6728 VSS.n5782 VSS.t740 1.19623
R6729 VSS.t715 VSS.n5851 1.19623
R6730 VSS.n4002 VSS.n3998 1.16717
R6731 VSS.n1764 VSS.n1763 1.16276
R6732 VSS.n1763 VSS.n1762 1.16276
R6733 VSS.n1762 VSS.n1761 1.16276
R6734 VSS.n1761 VSS.n1760 1.16276
R6735 VSS.n1760 VSS.n1759 1.16276
R6736 VSS.n1759 VSS.n1758 1.16276
R6737 VSS.n1758 VSS.n1757 1.16276
R6738 VSS.n1757 VSS.n1756 1.16276
R6739 VSS.n1756 VSS.n1755 1.16276
R6740 VSS.n1755 VSS.n1754 1.16276
R6741 VSS.n2468 VSS.n2467 1.16276
R6742 VSS.n2467 VSS.n2466 1.16276
R6743 VSS.n2466 VSS.n2465 1.16276
R6744 VSS.n2465 VSS.n2464 1.16276
R6745 VSS.n2464 VSS.n2463 1.16276
R6746 VSS.n2463 VSS.n2462 1.16276
R6747 VSS.n2462 VSS.n2461 1.16276
R6748 VSS.n2461 VSS.n2460 1.16276
R6749 VSS.n2460 VSS.n2459 1.16276
R6750 VSS.n2459 VSS.n2458 1.16276
R6751 VSS.n2382 VSS.n2381 1.16276
R6752 VSS.n2381 VSS.n2380 1.16276
R6753 VSS.n2380 VSS.n2379 1.16276
R6754 VSS.n2379 VSS.n2378 1.16276
R6755 VSS.n2378 VSS.n2377 1.16276
R6756 VSS.n2377 VSS.n2376 1.16276
R6757 VSS.n2376 VSS.n2375 1.16276
R6758 VSS.n2375 VSS.n2374 1.16276
R6759 VSS.n2374 VSS.n2373 1.16276
R6760 VSS.n2373 VSS.n2372 1.16276
R6761 VSS.n2265 VSS.n2264 1.16276
R6762 VSS.n2264 VSS.n2263 1.16276
R6763 VSS.n2263 VSS.n2262 1.16276
R6764 VSS.n2262 VSS.n2261 1.16276
R6765 VSS.n2261 VSS.n2260 1.16276
R6766 VSS.n2260 VSS.n2259 1.16276
R6767 VSS.n2259 VSS.n2258 1.16276
R6768 VSS.n2258 VSS.n2257 1.16276
R6769 VSS.n2257 VSS.n2256 1.16276
R6770 VSS.n2256 VSS.n2255 1.16276
R6771 VSS.n2158 VSS.n2157 1.16276
R6772 VSS.n2157 VSS.n2156 1.16276
R6773 VSS.n2156 VSS.n2155 1.16276
R6774 VSS.n2155 VSS.n2154 1.16276
R6775 VSS.n2154 VSS.n2153 1.16276
R6776 VSS.n2153 VSS.n2152 1.16276
R6777 VSS.n2152 VSS.n2151 1.16276
R6778 VSS.n2151 VSS.n2150 1.16276
R6779 VSS.n2150 VSS.n2149 1.16276
R6780 VSS.n2149 VSS.n2148 1.16276
R6781 VSS.n2061 VSS.n2060 1.16276
R6782 VSS.n2060 VSS.n2059 1.16276
R6783 VSS.n2059 VSS.n2058 1.16276
R6784 VSS.n2058 VSS.n2057 1.16276
R6785 VSS.n2057 VSS.n2056 1.16276
R6786 VSS.n2056 VSS.n2055 1.16276
R6787 VSS.n2055 VSS.n2054 1.16276
R6788 VSS.n2054 VSS.n2053 1.16276
R6789 VSS.n2053 VSS.n2052 1.16276
R6790 VSS.n2052 VSS.n2051 1.16276
R6791 VSS.n1991 VSS.n1990 1.16276
R6792 VSS.n1990 VSS.n1989 1.16276
R6793 VSS.n1989 VSS.n1988 1.16276
R6794 VSS.n1988 VSS.n1987 1.16276
R6795 VSS.n1987 VSS.n1986 1.16276
R6796 VSS.n1986 VSS.n1985 1.16276
R6797 VSS.n1985 VSS.n1984 1.16276
R6798 VSS.n1984 VSS.n1983 1.16276
R6799 VSS.n1983 VSS.n1982 1.16276
R6800 VSS.n1982 VSS.n1981 1.16276
R6801 VSS.n1836 VSS.n1835 1.16276
R6802 VSS.n1835 VSS.n1834 1.16276
R6803 VSS.n1834 VSS.n1833 1.16276
R6804 VSS.n1833 VSS.n1832 1.16276
R6805 VSS.n1832 VSS.n1831 1.16276
R6806 VSS.n1831 VSS.n1830 1.16276
R6807 VSS.n1830 VSS.n1829 1.16276
R6808 VSS.n1829 VSS.n1828 1.16276
R6809 VSS.n1828 VSS.n1827 1.16276
R6810 VSS.n1827 VSS.n1826 1.16276
R6811 VSS.n1802 VSS.n1801 1.16276
R6812 VSS.n1801 VSS.n1800 1.16276
R6813 VSS.n1800 VSS.n1799 1.16276
R6814 VSS.n1799 VSS.n1798 1.16276
R6815 VSS.n1798 VSS.n1797 1.16276
R6816 VSS.n1797 VSS.n1796 1.16276
R6817 VSS.n1796 VSS.n1795 1.16276
R6818 VSS.n1795 VSS.n1794 1.16276
R6819 VSS.n1794 VSS.n1793 1.16276
R6820 VSS.n1793 VSS.n1792 1.16276
R6821 VSS.n1781 VSS.n1780 1.16276
R6822 VSS.n1780 VSS.n1779 1.16276
R6823 VSS.n1779 VSS.n1778 1.16276
R6824 VSS.n1778 VSS.n1777 1.16276
R6825 VSS.n1777 VSS.n1776 1.16276
R6826 VSS.n1776 VSS.n1775 1.16276
R6827 VSS.n1775 VSS.n1774 1.16276
R6828 VSS.n1774 VSS.n1773 1.16276
R6829 VSS.n1773 VSS.n1772 1.16276
R6830 VSS.n1772 VSS.n1771 1.16276
R6831 VSS.n1753 VSS.n1752 1.16276
R6832 VSS.n1752 VSS.n1751 1.16276
R6833 VSS.n1751 VSS.n1750 1.16276
R6834 VSS.n1750 VSS.n1749 1.16276
R6835 VSS.n1749 VSS.n1748 1.16276
R6836 VSS.n1748 VSS.n1747 1.16276
R6837 VSS.n1747 VSS.n1746 1.16276
R6838 VSS.n1746 VSS.n1745 1.16276
R6839 VSS.n1745 VSS.n1744 1.16276
R6840 VSS.n1744 VSS.n1743 1.16276
R6841 VSS.n4991 VSS.n4924 1.15537
R6842 VSS.n3589 VSS.n3588 1.13934
R6843 VSS.n2487 VSS.n2486 1.12652
R6844 VSS.n353 VSS.n349 1.12642
R6845 VSS.n1447 VSS.n1446 1.1255
R6846 VSS.n318 VSS.n317 1.1255
R6847 VSS.n3822 VSS.n3821 1.1255
R6848 VSS.n3835 VSS.n3831 1.1255
R6849 VSS.n3749 VSS.n3748 1.1255
R6850 VSS.n3802 VSS.n3797 1.1255
R6851 VSS.n3766 VSS.n3761 1.1255
R6852 VSS.n3786 VSS.n3785 1.1255
R6853 VSS.n1742 VSS.n1741 1.1255
R6854 VSS.n3529 VSS.n3506 1.1255
R6855 VSS.n1770 VSS.n1769 1.1255
R6856 VSS.n1791 VSS.n1790 1.1255
R6857 VSS.n1825 VSS.n1824 1.1255
R6858 VSS.n1964 VSS.n1963 1.1255
R6859 VSS.n2026 VSS.n2024 1.1255
R6860 VSS.n2798 VSS.n2073 1.1255
R6861 VSS.n2853 VSS.n2852 1.1255
R6862 VSS.n2818 VSS.n2080 1.1255
R6863 VSS.n2020 VSS.n2007 1.1255
R6864 VSS.n2856 VSS.n2013 1.1255
R6865 VSS.n2048 VSS.n2047 1.1255
R6866 VSS.n2799 VSS.n2079 1.1255
R6867 VSS.n2017 VSS.n2002 1.1255
R6868 VSS.n1994 VSS.n1993 1.1255
R6869 VSS.n2779 VSS.n2102 1.1255
R6870 VSS.n2756 VSS.n2127 1.1255
R6871 VSS.n2188 VSS.n2169 1.1255
R6872 VSS.n2189 VSS.n2188 1.1255
R6873 VSS.n2774 VSS.n2108 1.1255
R6874 VSS.n2190 VSS.n2171 1.1255
R6875 VSS.n2137 VSS.n2115 1.1255
R6876 VSS.n2191 VSS.n2172 1.1255
R6877 VSS.n2704 VSS.n2234 1.1255
R6878 VSS.n2230 VSS.n2219 1.1255
R6879 VSS.n2691 VSS.n2247 1.1255
R6880 VSS.n2296 VSS.n2252 1.1255
R6881 VSS.n2306 VSS.n2275 1.1255
R6882 VSS.n2703 VSS.n2235 1.1255
R6883 VSS.n2297 VSS.n2253 1.1255
R6884 VSS.n2670 VSS.n2277 1.1255
R6885 VSS.n2640 VSS.n2639 1.1255
R6886 VSS.n2572 VSS.n2364 1.1255
R6887 VSS.n2575 VSS.n2395 1.1255
R6888 VSS.n2331 VSS.n2329 1.1255
R6889 VSS.n2329 VSS.n2325 1.1255
R6890 VSS.n2624 VSS.n2360 1.1255
R6891 VSS.n2577 VSS.n2576 1.1255
R6892 VSS.n2623 VSS.n2361 1.1255
R6893 VSS.n2578 VSS.n2399 1.1255
R6894 VSS.n2632 VSS.n2346 1.1255
R6895 VSS.n2544 VSS.n2429 1.1255
R6896 VSS.n2426 VSS.n2416 1.1255
R6897 VSS.n2530 VSS.n2438 1.1255
R6898 VSS.n2502 VSS.n2474 1.1255
R6899 VSS.n2483 VSS.n2475 1.1255
R6900 VSS.n2527 VSS.n2440 1.1255
R6901 VSS.n2488 VSS.n2479 1.1255
R6902 VSS.n2521 VSS.n2451 1.1255
R6903 VSS.n2418 VSS.n2416 1.1255
R6904 VSS.n2552 VSS.n2418 1.1255
R6905 VSS.n2502 VSS.n2501 1.1255
R6906 VSS.n2501 VSS.n2500 1.1255
R6907 VSS.n2436 VSS.n2434 1.1255
R6908 VSS.n2438 VSS.n2436 1.1255
R6909 VSS.n2411 VSS.n2410 1.1255
R6910 VSS.n2412 VSS.n2411 1.1255
R6911 VSS.n2477 VSS.n2475 1.1255
R6912 VSS.n2499 VSS.n2477 1.1255
R6913 VSS.n2526 VSS.n2525 1.1255
R6914 VSS.n2527 VSS.n2526 1.1255
R6915 VSS.n2497 VSS.n2479 1.1255
R6916 VSS.n2498 VSS.n2497 1.1255
R6917 VSS.n2522 VSS.n2447 1.1255
R6918 VSS.n2522 VSS.n2521 1.1255
R6919 VSS.n2648 VSS.n2325 1.1255
R6920 VSS.n2623 VSS.n2352 1.1255
R6921 VSS.n2319 VSS.n2318 1.1255
R6922 VSS.n2583 VSS.n2567 1.1255
R6923 VSS.n2576 VSS.n2394 1.1255
R6924 VSS.n2596 VSS.n2399 1.1255
R6925 VSS.n2600 VSS.n2395 1.1255
R6926 VSS.n2600 VSS.n2599 1.1255
R6927 VSS.n2625 VSS.n2359 1.1255
R6928 VSS.n2625 VSS.n2624 1.1255
R6929 VSS.n2366 VSS.n2364 1.1255
R6930 VSS.n2613 VSS.n2366 1.1255
R6931 VSS.n2597 VSS.n2596 1.1255
R6932 VSS.n2633 VSS.n2338 1.1255
R6933 VSS.n2633 VSS.n2632 1.1255
R6934 VSS.n2639 VSS.n2638 1.1255
R6935 VSS.n2598 VSS.n2394 1.1255
R6936 VSS.n2584 VSS.n2583 1.1255
R6937 VSS.n2638 VSS.n2637 1.1255
R6938 VSS.n2318 VSS.n2317 1.1255
R6939 VSS.n2367 VSS.n2352 1.1255
R6940 VSS.n2310 VSS.n2309 1.1255
R6941 VSS.n2684 VSS.n2252 1.1255
R6942 VSS.n2211 VSS.n2210 1.1255
R6943 VSS.n2683 VSS.n2253 1.1255
R6944 VSS.n2703 VSS.n2227 1.1255
R6945 VSS.n2672 VSS.n2275 1.1255
R6946 VSS.n2692 VSS.n2691 1.1255
R6947 VSS.n2713 VSS.n2219 1.1255
R6948 VSS.n2714 VSS.n2713 1.1255
R6949 VSS.n2693 VSS.n2692 1.1255
R6950 VSS.n2673 VSS.n2672 1.1255
R6951 VSS.n2227 VSS.n2226 1.1255
R6952 VSS.n2683 VSS.n2682 1.1255
R6953 VSS.n2671 VSS.n2274 1.1255
R6954 VSS.n2671 VSS.n2670 1.1255
R6955 VSS.n2705 VSS.n2704 1.1255
R6956 VSS.n2210 VSS.n2209 1.1255
R6957 VSS.n2706 VSS.n2705 1.1255
R6958 VSS.n2684 VSS.n2250 1.1255
R6959 VSS.n2316 VSS.n2310 1.1255
R6960 VSS.n2740 VSS.n2169 1.1255
R6961 VSS.n2737 VSS.n2172 1.1255
R6962 VSS.n2752 VSS.n2751 1.1255
R6963 VSS.n2768 VSS.n2115 1.1255
R6964 VSS.n2738 VSS.n2171 1.1255
R6965 VSS.n2774 VSS.n2773 1.1255
R6966 VSS.n2093 VSS.n2092 1.1255
R6967 VSS.n2760 VSS.n2125 1.1255
R6968 VSS.n2729 VSS.n2728 1.1255
R6969 VSS.n2159 VSS.n2126 1.1255
R6970 VSS.n2756 VSS.n2126 1.1255
R6971 VSS.n2781 VSS.n2780 1.1255
R6972 VSS.n2780 VSS.n2779 1.1255
R6973 VSS.n2761 VSS.n2760 1.1255
R6974 VSS.n2728 VSS.n2727 1.1255
R6975 VSS.n2092 VSS.n2091 1.1255
R6976 VSS.n2773 VSS.n2772 1.1255
R6977 VSS.n2739 VSS.n2738 1.1255
R6978 VSS.n2768 VSS.n2112 1.1255
R6979 VSS.n2751 VSS.n2750 1.1255
R6980 VSS.n2737 VSS.n2170 1.1255
R6981 VSS.n1993 VSS.n1992 1.1255
R6982 VSS.n2865 VSS.n2007 1.1255
R6983 VSS.n2852 VSS.n2851 1.1255
R6984 VSS.n2870 VSS.n2002 1.1255
R6985 VSS.n2079 VSS.n2074 1.1255
R6986 VSS.n2089 VSS.n2087 1.1255
R6987 VSS.n2820 VSS.n2819 1.1255
R6988 VSS.n2819 VSS.n2818 1.1255
R6989 VSS.n2032 VSS.n2011 1.1255
R6990 VSS.n2013 VSS.n2011 1.1255
R6991 VSS.n2050 VSS.n2048 1.1255
R6992 VSS.n2823 VSS.n2073 1.1255
R6993 VSS.n2823 VSS.n2822 1.1255
R6994 VSS.n2090 VSS.n2087 1.1255
R6995 VSS.n2836 VSS.n2050 1.1255
R6996 VSS.n2821 VSS.n2074 1.1255
R6997 VSS.n2871 VSS.n2870 1.1255
R6998 VSS.n2851 VSS.n2850 1.1255
R6999 VSS.n2849 VSS.n2028 1.1255
R7000 VSS.n2028 VSS.n2026 1.1255
R7001 VSS.n2865 VSS.n2864 1.1255
R7002 VSS.n1920 VSS.n1905 1.1255
R7003 VSS.n1945 VSS.n1944 1.1255
R7004 VSS.n1932 VSS.n1895 1.1255
R7005 VSS.n1923 VSS.n1896 1.1255
R7006 VSS.n1911 VSS.n1910 1.1255
R7007 VSS.n1947 VSS.n1946 1.1255
R7008 VSS.n1974 VSS.n1973 1.1255
R7009 VSS.n1954 VSS.n1886 1.1255
R7010 VSS.n1922 VSS.n1921 1.1255
R7011 VSS.n1979 VSS.n1879 1.1255
R7012 VSS.n3052 VSS.n1825 1.1255
R7013 VSS.n3027 VSS.n3022 1.1255
R7014 VSS.n3068 VSS.n3063 1.1255
R7015 VSS.n2961 VSS.n2959 1.1255
R7016 VSS.n2980 VSS.n2973 1.1255
R7017 VSS.n2981 VSS.n2980 1.1255
R7018 VSS.n2999 VSS.n2998 1.1255
R7019 VSS.n2998 VSS.n2997 1.1255
R7020 VSS.n2962 VSS.n2961 1.1255
R7021 VSS.n3014 VSS.n3011 1.1255
R7022 VSS.n3048 VSS.n3044 1.1255
R7023 VSS.n3049 VSS.n3048 1.1255
R7024 VSS.n3015 VSS.n3014 1.1255
R7025 VSS.n2984 VSS.n2983 1.1255
R7026 VSS.n2983 VSS.n2982 1.1255
R7027 VSS.n3037 VSS.n3036 1.1255
R7028 VSS.n3038 VSS.n3037 1.1255
R7029 VSS.n3069 VSS.n3068 1.1255
R7030 VSS.n3028 VSS.n3027 1.1255
R7031 VSS.n1812 VSS.n1808 1.1255
R7032 VSS.n3188 VSS.n1791 1.1255
R7033 VSS.n3102 VSS.n3097 1.1255
R7034 VSS.n3146 VSS.n3145 1.1255
R7035 VSS.n3186 VSS.n3181 1.1255
R7036 VSS.n3239 VSS.n3238 1.1255
R7037 VSS.n3115 VSS.n3110 1.1255
R7038 VSS.n3153 VSS.n3152 1.1255
R7039 VSS.n3089 VSS.n3087 1.1255
R7040 VSS.n3130 VSS.n3129 1.1255
R7041 VSS.n3170 VSS.n3165 1.1255
R7042 VSS.n3171 VSS.n3170 1.1255
R7043 VSS.n3131 VSS.n3130 1.1255
R7044 VSS.n3090 VSS.n3089 1.1255
R7045 VSS.n3198 VSS.n3197 1.1255
R7046 VSS.n3197 VSS.n3196 1.1255
R7047 VSS.n3154 VSS.n3153 1.1255
R7048 VSS.n3116 VSS.n3115 1.1255
R7049 VSS.n3240 VSS.n3239 1.1255
R7050 VSS.n3187 VSS.n3186 1.1255
R7051 VSS.n3147 VSS.n3146 1.1255
R7052 VSS.n3103 VSS.n3102 1.1255
R7053 VSS.n3359 VSS.n1770 1.1255
R7054 VSS.n3294 VSS.n3288 1.1255
R7055 VSS.n3335 VSS.n3328 1.1255
R7056 VSS.n3251 VSS.n3250 1.1255
R7057 VSS.n3298 VSS.n3297 1.1255
R7058 VSS.n3414 VSS.n3413 1.1255
R7059 VSS.n3413 VSS.n3412 1.1255
R7060 VSS.n3353 VSS.n3352 1.1255
R7061 VSS.n3354 VSS.n3353 1.1255
R7062 VSS.n3299 VSS.n3298 1.1255
R7063 VSS.n3252 VSS.n3251 1.1255
R7064 VSS.n3259 VSS.n3258 1.1255
R7065 VSS.n3258 VSS.n3257 1.1255
R7066 VSS.n3338 VSS.n3337 1.1255
R7067 VSS.n3314 VSS.n3311 1.1255
R7068 VSS.n3274 VSS.n3273 1.1255
R7069 VSS.n3339 VSS.n3338 1.1255
R7070 VSS.n3315 VSS.n3314 1.1255
R7071 VSS.n3275 VSS.n3274 1.1255
R7072 VSS.n3336 VSS.n3335 1.1255
R7073 VSS.n3295 VSS.n3294 1.1255
R7074 VSS.n3726 VSS.n1742 1.1255
R7075 VSS.n3662 VSS.n3657 1.1255
R7076 VSS.n3701 VSS.n3695 1.1255
R7077 VSS.n3647 VSS.n3646 1.1255
R7078 VSS.n3622 VSS.n3620 1.1255
R7079 VSS.n3636 VSS.n3631 1.1255
R7080 VSS.n3734 VSS.n3733 1.1255
R7081 VSS.n3721 VSS.n3717 1.1255
R7082 VSS.n3685 VSS.n3684 1.1255
R7083 VSS.n3684 VSS.n3683 1.1255
R7084 VSS.n3665 VSS.n3664 1.1255
R7085 VSS.n3709 VSS.n3708 1.1255
R7086 VSS.n3735 VSS.n3734 1.1255
R7087 VSS.n3710 VSS.n3709 1.1255
R7088 VSS.n3666 VSS.n3665 1.1255
R7089 VSS.n3637 VSS.n3636 1.1255
R7090 VSS.n3623 VSS.n3622 1.1255
R7091 VSS.n3722 VSS.n3721 1.1255
R7092 VSS.n3648 VSS.n3647 1.1255
R7093 VSS.n3702 VSS.n3701 1.1255
R7094 VSS.n3663 VSS.n3662 1.1255
R7095 VSS.n3787 VSS.n3786 1.1255
R7096 VSS.n3767 VSS.n3766 1.1255
R7097 VSS.n3750 VSS.n3749 1.1255
R7098 VSS.n3836 VSS.n3835 1.1255
R7099 VSS.n3803 VSS.n3802 1.1255
R7100 VSS.n3823 VSS.n3822 1.1255
R7101 VSS.n1642 VSS.n1641 1.1255
R7102 VSS.n1503 VSS.n1502 1.1234
R7103 VSS.n1814 VSS.n1813 1.12321
R7104 VSS.n1554 VSS.n1553 1.12277
R7105 VSS.n1544 VSS.n1543 1.12277
R7106 VSS.t169 VSS.n5930 1.10896
R7107 VSS.n5932 VSS.t590 1.10896
R7108 VSS.n316 VSS.n315 1.09796
R7109 VSS.n4012 VSS.n4011 1.06994
R7110 VSS.n4002 VSS.n4001 1.06994
R7111 VSS.n690 VSS.n688 1.03151
R7112 VSS.n916 VSS.n914 1.02489
R7113 VSS.n1397 VSS.n1395 1.02489
R7114 VSS.t178 VSS.t282 1.01328
R7115 VSS.n5136 VSS.n5134 1.01328
R7116 VSS.t275 VSS.t209 1.01328
R7117 VSS.t209 VSS.t184 1.01328
R7118 VSS.n1284 VSS.n1168 1.0102
R7119 VSS.n4158 VSS.n4157 0.972722
R7120 VSS.n4179 VSS.n4178 0.972722
R7121 VSS.n27 VSS.n26 0.967979
R7122 VSS.n2915 VSS.n1980 0.96059
R7123 VSS.n4150 VSS.t498 0.93818
R7124 VSS.n1322 VSS.n1321 0.93818
R7125 VSS.n1511 VSS.n1510 0.931667
R7126 VSS.n889 VSS.n888 0.929276
R7127 VSS.n879 VSS.n878 0.928071
R7128 VSS.n1450 VSS.n1449 0.925894
R7129 VSS.n4335 VSS.n253 0.919029
R7130 VSS.n4419 VSS.n4355 0.919029
R7131 VSS.n1012 VSS.n1010 0.910283
R7132 VSS.n5862 VSS.n5861 0.908479
R7133 VSS.n3086 VSS.n3085 0.900727
R7134 VSS.n2802 VSS.n2795 0.900647
R7135 VSS.n2663 VSS.n2662 0.900647
R7136 VSS.n2140 VSS.n2125 0.9005
R7137 VSS.n2753 VSS.n2752 0.9005
R7138 VSS.n3619 VSS.n3618 0.900467
R7139 VSS.n2958 VSS.n2957 0.900467
R7140 VSS.n2581 VSS.n2580 0.900467
R7141 VSS.n3407 VSS.n3406 0.900443
R7142 VSS.n3233 VSS.n3232 0.900443
R7143 VSS.n2657 VSS.n2656 0.900443
R7144 VSS.n2561 VSS.n2560 0.900442
R7145 VSS.n2880 VSS.n2879 0.900405
R7146 VSS.n2195 VSS.n2193 0.900387
R7147 VSS.n1909 VSS.n1908 0.900368
R7148 VSS.n2790 VSS.n2789 0.900365
R7149 VSS.n2723 VSS.n2722 0.900365
R7150 VSS.n1874 VSS.n1873 0.900347
R7151 VSS.n1556 VSS.n1555 0.900305
R7152 VSS.n1644 VSS.n1643 0.90028
R7153 VSS.n336 VSS.n335 0.898922
R7154 VSS.n1807 VSS.n1806 0.898321
R7155 VSS.n314 VSS.n308 0.897993
R7156 VSS.n1646 VSS.n1645 0.891062
R7157 VSS.n4193 VSS.n4189 0.8755
R7158 VSS.n564 VSS.n563 0.849401
R7159 VSS.n683 VSS.n682 0.849401
R7160 VSS.n6020 VSS.n6019 0.849401
R7161 VSS.n6038 VSS.n6037 0.849401
R7162 VSS.n6059 VSS.n6058 0.849401
R7163 VSS.n5675 VSS.n5674 0.849401
R7164 VSS.n5351 VSS.n5350 0.849205
R7165 VSS.n978 VSS.n977 0.846031
R7166 VSS.n990 VSS.n989 0.846031
R7167 VSS.n4347 VSS.n4346 0.845835
R7168 VSS.n4332 VSS.n4331 0.845835
R7169 VSS.n882 VSS.n874 0.829906
R7170 VSS VSS.n4746 0.805351
R7171 VSS.n5850 VSS.n5849 0.801258
R7172 VSS.n4137 VSS.n4134 0.79929
R7173 VSS.n5911 VSS 0.793969
R7174 VSS.n5747 VSS.n5746 0.781777
R7175 VSS.n5755 VSS.n5754 0.781777
R7176 VSS.n1299 VSS.n1298 0.780455
R7177 VSS.n4689 VSS.n4685 0.778278
R7178 VSS.n1520 VSS.n1519 0.778278
R7179 VSS.n5808 VSS.n5807 0.772481
R7180 VSS.n315 VSS.n314 0.768418
R7181 VSS.n4203 VSS.n4201 0.726531
R7182 VSS.n5849 VSS.n5774 0.722141
R7183 VSS.n4107 VSS.n4106 0.69552
R7184 VSS.n4239 VSS.n4238 0.69552
R7185 VSS.n1033 VSS 0.683795
R7186 VSS.n1464 VSS.n1416 0.681056
R7187 VSS.n4997 VSS.n4996 0.66722
R7188 VSS.n4603 VSS.n4602 0.66701
R7189 VSS.n4592 VSS.n4591 0.66701
R7190 VSS.n4658 VSS.n4657 0.66701
R7191 VSS.n4671 VSS.n4670 0.66701
R7192 VSS.n4573 VSS.n4572 0.66701
R7193 VSS.n3893 VSS.n1719 0.652915
R7194 VSS.n4005 VSS.t768 0.65037
R7195 VSS.n3858 VSS.n1720 0.643803
R7196 VSS.n140 VSS.n137 0.642239
R7197 VSS.n183 VSS.n180 0.642239
R7198 VSS.n238 VSS.n235 0.642239
R7199 VSS.n5193 VSS.n5192 0.642239
R7200 VSS.n5219 VSS.n5218 0.642239
R7201 VSS.n4799 VSS.n4798 0.642239
R7202 VSS.n2835 VSS.n2061 0.615498
R7203 VSS.n2161 VSS.n2158 0.614262
R7204 VSS.n4502 VSS.n4501 0.611348
R7205 VSS.n5548 VSS.n5547 0.610998
R7206 VSS.n2266 VSS.n2265 0.609999
R7207 VSS.n3431 VSS.n1764 0.609008
R7208 VSS.n3003 VSS.n1836 0.608439
R7209 VSS.n3703 VSS.n1753 0.606848
R7210 VSS.n2612 VSS.n2382 0.606843
R7211 VSS.n3156 VSS.n1802 0.606489
R7212 VSS.n3316 VSS.n1781 0.605607
R7213 VSS.n2896 VSS.n1991 0.601243
R7214 VSS.n235 VSS.n232 0.597879
R7215 VSS.n4798 VSS.n4797 0.597879
R7216 VSS.n137 VSS.n134 0.596788
R7217 VSS.n5218 VSS.n5217 0.596788
R7218 VSS.n180 VSS.n177 0.595696
R7219 VSS.n5192 VSS.n5191 0.595696
R7220 VSS.n2512 VSS.n2468 0.593624
R7221 VSS.n174 VSS.n173 0.587994
R7222 VSS.n5190 VSS.n5189 0.587128
R7223 VSS.n131 VSS.n130 0.586903
R7224 VSS.n5216 VSS.n5215 0.586037
R7225 VSS.n229 VSS.n228 0.585812
R7226 VSS.n4796 VSS.n4795 0.584946
R7227 VSS.n834 VSS.n833 0.583833
R7228 VSS.n5215 VSS.n5214 0.574718
R7229 VSS.n130 VSS.n127 0.574288
R7230 VSS.n4795 VSS.n4794 0.573627
R7231 VSS.n228 VSS.n225 0.573197
R7232 VSS.n3530 VSS.n3529 0.563
R7233 VSS.n2544 VSS.n2425 0.563
R7234 VSS.n2425 VSS.n2423 0.563
R7235 VSS.n2433 VSS.n2423 0.563
R7236 VSS.n3566 VSS.n3530 0.563
R7237 VSS.n3567 VSS.n3566 0.563
R7238 VSS.n1567 VSS.n1566 0.551597
R7239 VSS.n173 VSS.n170 0.550283
R7240 VSS.n5189 VSS.n5188 0.550283
R7241 VSS.n4363 VSS.n4362 0.54076
R7242 VSS.n5898 VSS.n5897 0.5405
R7243 VSS.n3738 VSS.n1728 0.534462
R7244 VSS.n5935 VSS.n4745 0.508005
R7245 VSS.n4743 VSS.n4742 0.508005
R7246 VSS.n6007 VSS.n6006 0.507764
R7247 VSS.n511 VSS.n510 0.505601
R7248 VSS.n4317 VSS.n4316 0.505601
R7249 VSS.n963 VSS.n962 0.502377
R7250 VSS.n4366 VSS.n4365 0.502362
R7251 VSS.n5286 VSS.n5285 0.502362
R7252 VSS.n4369 VSS.n4368 0.497425
R7253 VSS.n5289 VSS.n5288 0.497402
R7254 VSS.n4025 VSS.n4024 0.486611
R7255 VSS.n5864 VSS.n5756 0.477891
R7256 VSS.n3242 VSS.n3241 0.473104
R7257 VSS.n940 VSS.n939 0.472687
R7258 VSS.n4136 VSS.n4135 0.472687
R7259 VSS.n2660 VSS.n2659 0.467151
R7260 VSS.n3416 VSS.n3415 0.465504
R7261 VSS.n1328 VSS.n1327 0.459689
R7262 VSS.n4117 VSS.n4116 0.459689
R7263 VSS.n1369 VSS.n1368 0.459446
R7264 VSS.n1286 VSS.n1285 0.459446
R7265 VSS.n3842 VSS.n3841 0.459227
R7266 VSS.n2916 VSS.n2915 0.458913
R7267 VSS.n5865 VSS.n5749 0.458326
R7268 VSS.n2726 VSS.n2725 0.456584
R7269 VSS.n2793 VSS.n2792 0.451624
R7270 VSS.n2564 VSS.n2563 0.449946
R7271 VSS.n1403 VSS 0.449668
R7272 VSS.n3072 VSS.n3071 0.443676
R7273 VSS.n3574 VSS.n3573 0.441768
R7274 VSS.n66 VSS.n65 0.435547
R7275 VSS.n5123 VSS.n5122 0.434956
R7276 VSS.n5934 VSS.n4746 0.434362
R7277 VSS.n4117 VSS.n4111 0.4313
R7278 VSS.n117 VSS.n116 0.427022
R7279 VSS.n4778 VSS.n4775 0.426043
R7280 VSS VSS.n1402 0.405813
R7281 VSS.n489 VSS.n488 0.402035
R7282 VSS.n4044 VSS.n4043 0.402035
R7283 VSS.n364 VSS.n363 0.402035
R7284 VSS.n504 VSS.n503 0.402035
R7285 VSS.n4309 VSS.n4308 0.402035
R7286 VSS.n4111 VSS.n4108 0.402035
R7287 VSS.n4275 VSS.n4274 0.402035
R7288 VSS.n4273 VSS.n4272 0.402035
R7289 VSS.n3914 VSS.n3913 0.402035
R7290 VSS.n4106 VSS.n4105 0.401791
R7291 VSS.n5492 VSS.n5489 0.393137
R7292 VSS.n4516 VSS.n4513 0.393137
R7293 VSS.n5556 VSS.n5555 0.391771
R7294 VSS.n735 VSS.n732 0.390642
R7295 VSS.n511 VSS.n504 0.390642
R7296 VSS.n773 VSS.n770 0.390642
R7297 VSS.n4312 VSS.n4309 0.390642
R7298 VSS.n28 VSS.n27 0.383479
R7299 VSS.n249 VSS.n248 0.383166
R7300 VSS.n4393 VSS.n4392 0.383166
R7301 VSS.n1014 VSS.n1013 0.383166
R7302 VSS.n49 VSS.n48 0.382921
R7303 VSS.n4416 VSS.n4415 0.382921
R7304 VSS.n4780 VSS.n4779 0.382921
R7305 VSS.n5137 VSS.n5136 0.382921
R7306 VSS.n5136 VSS.n5135 0.382921
R7307 VSS.n4561 VSS.n4511 0.376519
R7308 VSS.n4582 VSS.n94 0.376518
R7309 VSS.n5078 VSS.n5077 0.37489
R7310 VSS.n5092 VSS.n5065 0.374889
R7311 VSS.n5171 VSS.n5170 0.372135
R7312 VSS.n161 VSS.n148 0.372135
R7313 VSS.n4402 VSS.n4401 0.371392
R7314 VSS.n5314 VSS.n5313 0.371022
R7315 VSS.n4399 VSS.n4398 0.370645
R7316 VSS.n5311 VSS.n5310 0.370645
R7317 VSS.n5062 VSS.n5060 0.358977
R7318 VSS.n4614 VSS.n4611 0.358977
R7319 VSS.n4601 VSS.n63 0.356537
R7320 VSS.n5140 VSS.n5063 0.354994
R7321 VSS.n6101 VSS.n28 0.350926
R7322 VSS.n5919 VSS 0.347643
R7323 VSS VSS.n5922 0.347643
R7324 VSS.n5787 VSS 0.347643
R7325 VSS VSS.n5840 0.347643
R7326 VSS.n5069 VSS.n5066 0.347591
R7327 VSS.n6098 VSS.n6096 0.342028
R7328 VSS.n147 VSS.n146 0.341179
R7329 VSS.n5169 VSS.n5168 0.340476
R7330 VSS.n106 VSS.n105 0.338978
R7331 VSS.n5650 VSS.n5329 0.331895
R7332 VSS.n5633 VSS.n5331 0.331895
R7333 VSS.n3980 VSS.n3977 0.327038
R7334 VSS.n5618 VSS.n5617 0.326081
R7335 VSS.n5115 VSS.n5064 0.321363
R7336 VSS.n4590 VSS.n76 0.320022
R7337 VSS.n5824 VSS.n5813 0.3191
R7338 VSS.n5823 VSS.n5819 0.3191
R7339 VSS.n5817 VSS.n5816 0.3191
R7340 VSS.n5892 VSS.n5886 0.3191
R7341 VSS.n5894 VSS.n5881 0.3191
R7342 VSS.n5897 VSS.n5896 0.3191
R7343 VSS.n4754 VSS.n4751 0.3191
R7344 VSS.n4758 VSS.n4755 0.3191
R7345 VSS.n5895 VSS.n5880 0.3191
R7346 VSS.n5893 VSS.n5885 0.3191
R7347 VSS.n5835 VSS.n5795 0.3191
R7348 VSS.n5167 VSS.n5166 0.31827
R7349 VSS.n145 VSS.n144 0.318076
R7350 VSS.n5834 VSS.n5833 0.315513
R7351 VSS.n4570 VSS.n4510 0.313628
R7352 VSS VSS.n2882 0.307487
R7353 VSS.n259 VSS.n257 0.302495
R7354 VSS.n5664 VSS.n5271 0.301198
R7355 VSS.n1167 VSS.n1166 0.3005
R7356 VSS.n5829 VSS.n5799 0.2957
R7357 VSS.n5803 VSS.n5802 0.2957
R7358 VSS.n5822 VSS.n5821 0.2957
R7359 VSS.n5825 VSS.n5811 0.2957
R7360 VSS.n4995 VSS.n4807 0.292445
R7361 VSS.n80 VSS.n79 0.291512
R7362 VSS.n4674 VSS.n58 0.290903
R7363 VSS.n5007 VSS.n4806 0.289506
R7364 VSS.n4987 VSS.n4925 0.288772
R7365 VSS.n4664 VSS.n59 0.287963
R7366 VSS.n57 VSS.n31 0.287229
R7367 VSS.n4966 VSS.n4965 0.285098
R7368 VSS.n4977 VSS.n4964 0.285098
R7369 VSS.n39 VSS.n33 0.283556
R7370 VSS.n47 VSS.n32 0.283556
R7371 VSS.n4275 VSS 0.281962
R7372 VSS.n5849 VSS.n5848 0.281211
R7373 VSS.n240 VSS.n239 0.2753
R7374 VSS.n5249 VSS.n4800 0.2753
R7375 VSS.n3877 VSS.n3876 0.274296
R7376 VSS.n221 VSS.n220 0.2729
R7377 VSS.n5220 VSS.n5202 0.2729
R7378 VSS.n184 VSS.n183 0.272046
R7379 VSS.n5194 VSS.n5193 0.27149
R7380 VSS.n241 VSS.n240 0.269479
R7381 VSS.n5251 VSS.n5249 0.269479
R7382 VSS.n3874 VSS.n3873 0.266088
R7383 VSS.n4504 VSS.n4503 0.254764
R7384 VSS.n220 VSS.n140 0.250935
R7385 VSS.n239 VSS.n238 0.250935
R7386 VSS.n5220 VSS.n5219 0.250935
R7387 VSS.n4800 VSS.n4799 0.250935
R7388 VSS.n5144 VSS.n5143 0.2505
R7389 VSS.n4607 VSS.n4606 0.2505
R7390 VSS.n142 VSS.n141 0.24562
R7391 VSS.n5101 VSS.n5098 0.244911
R7392 VSS.n952 VSS 0.243106
R7393 VSS.n5860 VSS.n5761 0.241879
R7394 VSS.n5320 VSS.n5319 0.241152
R7395 VSS.n5101 VSS.n5100 0.239887
R7396 VSS.n4376 VSS.n4357 0.235283
R7397 VSS.n4252 VSS.n4219 0.224214
R7398 VSS.n83 VSS.n77 0.213053
R7399 VSS.n93 VSS.n84 0.213053
R7400 VSS.n75 VSS.n64 0.213053
R7401 VSS.n5132 VSS.n5121 0.213053
R7402 VSS.n5111 VSS.n5105 0.213053
R7403 VSS.n5104 VSS.n5096 0.213053
R7404 VSS.n5108 VSS.n5107 0.211098
R7405 VSS.n4130 VSS.n908 0.205426
R7406 VSS.n5251 VSS.n5250 0.205144
R7407 VSS.n4890 VSS.n4889 0.205045
R7408 VSS.n5749 VSS.n5747 0.200065
R7409 VSS.n5756 VSS.n5755 0.200065
R7410 VSS.n143 VSS.n142 0.199702
R7411 VSS.n406 VSS.n360 0.1985
R7412 VSS.n4893 VSS.n4890 0.196574
R7413 VSS.n72 VSS.n71 0.196132
R7414 VSS.n5129 VSS.n5128 0.196132
R7415 VSS VSS.n1032 0.195846
R7416 VSS.n4050 VSS.n4031 0.193921
R7417 VSS.n4064 VSS.n1523 0.193087
R7418 VSS.n5767 VSS.n5763 0.188841
R7419 VSS.n413 VSS.n322 0.188079
R7420 VSS.n1174 VSS.n1171 0.188
R7421 VSS.n239 VSS.n221 0.1865
R7422 VSS.n5202 VSS.n4800 0.1865
R7423 VSS.n351 VSS.n350 0.185092
R7424 VSS.n220 VSS.n219 0.1805
R7425 VSS.n5221 VSS.n5220 0.1805
R7426 VSS.n4552 VSS.n4549 0.174181
R7427 VSS.n5528 VSS.n5525 0.17414
R7428 VSS.n4407 VSS.n4406 0.174137
R7429 VSS.n5320 VSS.n5318 0.172819
R7430 VSS.n90 VSS.n89 0.170926
R7431 VSS.n4120 VSS.n4119 0.169688
R7432 VSS.n21 VSS.n20 0.167572
R7433 VSS.n4311 VSS.n4310 0.164562
R7434 VSS.n3871 VSS.n3870 0.163308
R7435 VSS.n5170 VSS.n5169 0.163136
R7436 VSS.n148 VSS.n147 0.162433
R7437 VSS.n4205 VSS.n4203 0.161214
R7438 VSS.n954 VSS.n952 0.161214
R7439 VSS.n4121 VSS.n4120 0.161214
R7440 VSS.n4134 VSS.n4132 0.161214
R7441 VSS.n497 VSS.n493 0.160198
R7442 VSS.n5806 VSS.n5805 0.159119
R7443 VSS.n5912 VSS.n5911 0.157743
R7444 VSS.n4411 VSS.n4410 0.157329
R7445 VSS.n5325 VSS.n5323 0.15648
R7446 VSS.n5913 VSS.n5912 0.156251
R7447 VSS VSS.n4205 0.155589
R7448 VSS.n5304 VSS.n5299 0.155512
R7449 VSS.n4386 VSS.n4383 0.153637
R7450 VSS.n5168 VSS.n5167 0.153513
R7451 VSS.n4505 VSS.n4504 0.152808
R7452 VSS.n1293 VSS.n1290 0.15275
R7453 VSS.n146 VSS.n145 0.152738
R7454 VSS.n4557 VSS.n4556 0.152674
R7455 VSS.n4091 VSS.n4090 0.151571
R7456 VSS.n4129 VSS.n4127 0.151571
R7457 VSS.n961 VSS.n960 0.150768
R7458 VSS.n5017 VSS.n5011 0.150235
R7459 VSS.n4660 VSS.n4656 0.150235
R7460 VSS.n5036 VSS.n5033 0.148852
R7461 VSS.n5039 VSS.n5036 0.148852
R7462 VSS.n5042 VSS.n5039 0.148852
R7463 VSS.n5045 VSS.n5042 0.148852
R7464 VSS.n5048 VSS.n5045 0.148852
R7465 VSS.n5051 VSS.n5048 0.148852
R7466 VSS.n5054 VSS.n5051 0.148852
R7467 VSS.n5057 VSS.n5054 0.148852
R7468 VSS.n5060 VSS.n5057 0.148852
R7469 VSS.n5495 VSS.n5492 0.148852
R7470 VSS.n5498 VSS.n5495 0.148852
R7471 VSS.n5501 VSS.n5498 0.148852
R7472 VSS.n5504 VSS.n5501 0.148852
R7473 VSS.n5507 VSS.n5504 0.148852
R7474 VSS.n5510 VSS.n5507 0.148852
R7475 VSS.n5513 VSS.n5510 0.148852
R7476 VSS.n5516 VSS.n5513 0.148852
R7477 VSS.n5519 VSS.n5516 0.148852
R7478 VSS.n5522 VSS.n5519 0.148852
R7479 VSS.n4617 VSS.n4614 0.148852
R7480 VSS.n4620 VSS.n4617 0.148852
R7481 VSS.n4623 VSS.n4620 0.148852
R7482 VSS.n4626 VSS.n4623 0.148852
R7483 VSS.n4629 VSS.n4626 0.148852
R7484 VSS.n4632 VSS.n4629 0.148852
R7485 VSS.n4635 VSS.n4632 0.148852
R7486 VSS.n4638 VSS.n4635 0.148852
R7487 VSS.n4641 VSS.n4638 0.148852
R7488 VSS.n4546 VSS.n4543 0.148852
R7489 VSS.n4543 VSS.n4540 0.148852
R7490 VSS.n4540 VSS.n4537 0.148852
R7491 VSS.n4537 VSS.n4534 0.148852
R7492 VSS.n4534 VSS.n4531 0.148852
R7493 VSS.n4531 VSS.n4528 0.148852
R7494 VSS.n4528 VSS.n4525 0.148852
R7495 VSS.n4525 VSS.n4522 0.148852
R7496 VSS.n4522 VSS.n4519 0.148852
R7497 VSS.n4519 VSS.n4516 0.148852
R7498 VSS.n4119 VSS.n919 0.148402
R7499 VSS.n4391 VSS.n4389 0.147239
R7500 VSS.n167 VSS.n164 0.147239
R7501 VSS.n211 VSS.n208 0.147239
R7502 VSS.n214 VSS.n211 0.147239
R7503 VSS.n201 VSS.n198 0.147239
R7504 VSS.n204 VSS.n201 0.147239
R7505 VSS.n116 VSS.n113 0.147239
R7506 VSS.n251 VSS.n247 0.147239
R7507 VSS.n5177 VSS.n5174 0.147239
R7508 VSS.n5241 VSS.n5238 0.147239
R7509 VSS.n5244 VSS.n5241 0.147239
R7510 VSS.n5231 VSS.n5228 0.147239
R7511 VSS.n5234 VSS.n5231 0.147239
R7512 VSS.n4775 VSS.n4772 0.147239
R7513 VSS.n5269 VSS.n5267 0.147239
R7514 VSS.n5263 VSS.n5261 0.147239
R7515 VSS.n4427 VSS.n4424 0.147239
R7516 VSS.n4424 VSS.n4422 0.147239
R7517 VSS.n2883 VSS 0.145448
R7518 VSS.n4758 VSS.n4757 0.144944
R7519 VSS.n5433 VSS.n5430 0.144304
R7520 VSS.n4433 VSS.n4430 0.144304
R7521 VSS.n5325 VSS.n5307 0.142348
R7522 VSS.n4414 VSS.n4413 0.142348
R7523 VSS.n4413 VSS.n4411 0.14137
R7524 VSS.n5525 VSS.n5522 0.139951
R7525 VSS.n4549 VSS.n4546 0.139951
R7526 VSS.n1302 VSS.n973 0.139082
R7527 VSS.n5296 VSS.n5295 0.137463
R7528 VSS.n4376 VSS.n4375 0.136472
R7529 VSS.n3739 VSS.n3738 0.133072
R7530 VSS.n290 VSS.n289 0.132286
R7531 VSS.n245 VSS.n244 0.131851
R7532 VSS.n5866 VSS.n5865 0.131118
R7533 VSS.n160 VSS.n157 0.130588
R7534 VSS.n109 VSS.n108 0.130302
R7535 VSS.n5161 VSS.n5158 0.130084
R7536 VSS.n5259 VSS.n5258 0.129374
R7537 VSS.n1374 VSS.n1371 0.12841
R7538 VSS.n1257 VSS.n1254 0.128
R7539 VSS.n5257 VSS.n5256 0.125349
R7540 VSS.n4171 VSS.n4170 0.12483
R7541 VSS.n107 VSS.n106 0.124421
R7542 VSS.n5297 VSS.n5296 0.123458
R7543 VSS.n244 VSS.n243 0.122817
R7544 VSS.n4430 VSS.n4427 0.122783
R7545 VSS.n5273 VSS.n5272 0.122669
R7546 VSS.n4377 VSS.n4376 0.122609
R7547 VSS.n1510 VSS.n1509 0.1225
R7548 VSS.n5321 VSS.n5320 0.12249
R7549 VSS.n5254 VSS.n5253 0.121959
R7550 VSS.n4379 VSS.n4378 0.121915
R7551 VSS.n5323 VSS.n5322 0.121915
R7552 VSS.n5299 VSS.n5298 0.121915
R7553 VSS.n4410 VSS.n4409 0.121915
R7554 VSS.n4381 VSS.n4380 0.121893
R7555 VSS.n106 VSS.n103 0.121804
R7556 VSS.n5256 VSS.n5255 0.121804
R7557 VSS.n4408 VSS.n4407 0.121641
R7558 VSS.n5799 VSS.n5798 0.121611
R7559 VSS.n215 VSS.n191 0.120826
R7560 VSS.n4782 VSS.n4778 0.120826
R7561 VSS.n5088 VSS.n5085 0.119969
R7562 VSS.n5145 VSS.n5142 0.119969
R7563 VSS.n5082 VSS.n5080 0.119969
R7564 VSS.n5011 VSS.n5010 0.119969
R7565 VSS.n5006 VSS.n5003 0.119969
R7566 VSS.n5003 VSS.n4999 0.119969
R7567 VSS.n4982 VSS.n4980 0.119969
R7568 VSS.n4976 VSS.n4973 0.119969
R7569 VSS.n4973 VSS.n4969 0.119969
R7570 VSS.n5486 VSS.n5483 0.119969
R7571 VSS.n5489 VSS.n5486 0.119969
R7572 VSS.n4608 VSS.n4605 0.119969
R7573 VSS.n4567 VSS.n4564 0.119969
R7574 VSS.n4569 VSS.n4567 0.119969
R7575 VSS.n4578 VSS.n4575 0.119969
R7576 VSS.n38 VSS.n35 0.119969
R7577 VSS.n44 VSS.n41 0.119969
R7578 VSS.n46 VSS.n44 0.119969
R7579 VSS.n54 VSS.n51 0.119969
R7580 VSS.n56 VSS.n54 0.119969
R7581 VSS.n4680 VSS.n4677 0.119969
R7582 VSS.n4673 VSS.n4669 0.119969
R7583 VSS.n4669 VSS.n4666 0.119969
R7584 VSS.n4663 VSS.n4660 0.119969
R7585 VSS.n120 VSS.n117 0.119848
R7586 VSS.n5225 VSS.n5201 0.119848
R7587 VSS.n4165 VSS.n4164 0.119263
R7588 VSS.n888 VSS.n887 0.119263
R7589 VSS.n4558 VSS.n4555 0.119173
R7590 VSS.n5472 VSS.n5469 0.118921
R7591 VSS.n5469 VSS.n5466 0.118921
R7592 VSS.n5459 VSS.n5456 0.118921
R7593 VSS.n5456 VSS.n5453 0.118921
R7594 VSS.n5453 VSS.n5450 0.118921
R7595 VSS.n5450 VSS.n5447 0.118921
R7596 VSS.n5554 VSS.n5551 0.118921
R7597 VSS.n4446 VSS.n4443 0.118921
R7598 VSS.n4449 VSS.n4446 0.118921
R7599 VSS.n4452 VSS.n4449 0.118921
R7600 VSS.n4455 VSS.n4452 0.118921
R7601 VSS.n4458 VSS.n4455 0.118921
R7602 VSS.n4461 VSS.n4458 0.118921
R7603 VSS.n4464 VSS.n4461 0.118921
R7604 VSS.n4467 VSS.n4464 0.118921
R7605 VSS.n4474 VSS.n4471 0.118921
R7606 VSS.n4477 VSS.n4474 0.118921
R7607 VSS.n4480 VSS.n4477 0.118921
R7608 VSS.n4483 VSS.n4480 0.118921
R7609 VSS.n4486 VSS.n4483 0.118921
R7610 VSS.n108 VSS.n107 0.118335
R7611 VSS.n5258 VSS.n5257 0.118335
R7612 VSS.n4555 VSS.n4552 0.116783
R7613 VSS.n5444 VSS.n5443 0.116553
R7614 VSS.n5436 VSS.n5433 0.115403
R7615 VSS.n5531 VSS.n5530 0.115328
R7616 VSS.n4436 VSS.n4433 0.115214
R7617 VSS.n1340 VSS.n1338 0.113945
R7618 VSS.n1338 VSS.n1336 0.113945
R7619 VSS.n1332 VSS.n1330 0.113945
R7620 VSS.n1330 VSS.n1326 0.113945
R7621 VSS.n1326 VSS.n1324 0.113945
R7622 VSS.n1324 VSS.n1320 0.113945
R7623 VSS.n1320 VSS.n1316 0.113945
R7624 VSS.n1316 VSS.n1313 0.113945
R7625 VSS.n1308 VSS.n1307 0.113945
R7626 VSS.n1307 VSS.n1304 0.113945
R7627 VSS.n1377 VSS.n1374 0.113945
R7628 VSS.n1380 VSS.n1377 0.113945
R7629 VSS.n1384 VSS.n1380 0.113945
R7630 VSS.n1387 VSS.n1384 0.113945
R7631 VSS.n1391 VSS.n1387 0.113945
R7632 VSS.n4099 VSS.n4096 0.113945
R7633 VSS.n1301 VSS.n1297 0.113933
R7634 VSS.n5530 VSS.n5528 0.113776
R7635 VSS.n5083 VSS.n5082 0.113597
R7636 VSS.n874 VSS.n873 0.113103
R7637 VSS.n1290 VSS.n1288 0.113
R7638 VSS.n1297 VSS.n1293 0.113
R7639 VSS.n687 VSS.n685 0.113
R7640 VSS.n1259 VSS.n1257 0.113
R7641 VSS.n1262 VSS.n1259 0.113
R7642 VSS.n1265 VSS.n1262 0.113
R7643 VSS.n1268 VSS.n1265 0.113
R7644 VSS.n1271 VSS.n1268 0.113
R7645 VSS.n1274 VSS.n1271 0.113
R7646 VSS.n1277 VSS.n1274 0.113
R7647 VSS.n1280 VSS.n1277 0.113
R7648 VSS.n1283 VSS.n1280 0.113
R7649 VSS.n1178 VSS.n1174 0.113
R7650 VSS.n1181 VSS.n1178 0.113
R7651 VSS.n1184 VSS.n1181 0.113
R7652 VSS.n1187 VSS.n1184 0.113
R7653 VSS.n1190 VSS.n1187 0.113
R7654 VSS.n1193 VSS.n1190 0.113
R7655 VSS.n1196 VSS.n1193 0.113
R7656 VSS.n1199 VSS.n1196 0.113
R7657 VSS.n1203 VSS.n1199 0.113
R7658 VSS.n1206 VSS.n1203 0.113
R7659 VSS.n1209 VSS.n1206 0.113
R7660 VSS.n1212 VSS.n1209 0.113
R7661 VSS.n1215 VSS.n1212 0.113
R7662 VSS.n1218 VSS.n1215 0.113
R7663 VSS.n1221 VSS.n1218 0.113
R7664 VSS.n1224 VSS.n1221 0.113
R7665 VSS.n1228 VSS.n1224 0.113
R7666 VSS.n1231 VSS.n1228 0.113
R7667 VSS.n1234 VSS.n1231 0.113
R7668 VSS.n1237 VSS.n1234 0.113
R7669 VSS.n1240 VSS.n1237 0.113
R7670 VSS.n1243 VSS.n1240 0.113
R7671 VSS.n1246 VSS.n1243 0.113
R7672 VSS.n1249 VSS.n1246 0.113
R7673 VSS.n1251 VSS.n1249 0.113
R7674 VSS.n1254 VSS.n1251 0.113
R7675 VSS.n1345 VSS.n1342 0.113
R7676 VSS.n1347 VSS.n1345 0.113
R7677 VSS.n1350 VSS.n1347 0.113
R7678 VSS.n1352 VSS.n1350 0.113
R7679 VSS.n1355 VSS.n1352 0.113
R7680 VSS.n1357 VSS.n1355 0.113
R7681 VSS.n1360 VSS.n1357 0.113
R7682 VSS.n1362 VSS.n1360 0.113
R7683 VSS.n1365 VSS.n1362 0.113
R7684 VSS.n1367 VSS.n1365 0.113
R7685 VSS.n1371 VSS.n1367 0.113
R7686 VSS.n1164 VSS.n1161 0.112367
R7687 VSS.n4414 VSS.n4379 0.111845
R7688 VSS.n4383 VSS.n4382 0.111448
R7689 VSS.n5275 VSS.n5274 0.111448
R7690 VSS.n491 VSS.n487 0.111156
R7691 VSS.n493 VSS.n491 0.111156
R7692 VSS.n487 VSS.n485 0.11043
R7693 VSS.n763 VSS.n760 0.110256
R7694 VSS.n760 VSS.n757 0.110256
R7695 VSS.n757 VSS.n754 0.110256
R7696 VSS.n4070 VSS.n4067 0.110256
R7697 VSS.n4083 VSS.n4070 0.110256
R7698 VSS.n4083 VSS.n4082 0.110256
R7699 VSS.n4082 VSS.n4079 0.110256
R7700 VSS.n4079 VSS.n4076 0.110256
R7701 VSS.n4076 VSS.n4073 0.110256
R7702 VSS.n366 VSS.n362 0.110256
R7703 VSS.n368 VSS.n366 0.110256
R7704 VSS.n371 VSS.n368 0.110256
R7705 VSS.n374 VSS.n371 0.110256
R7706 VSS.n377 VSS.n374 0.110256
R7707 VSS.n380 VSS.n377 0.110256
R7708 VSS.n383 VSS.n380 0.110256
R7709 VSS.n386 VSS.n383 0.110256
R7710 VSS.n389 VSS.n386 0.110256
R7711 VSS.n393 VSS.n389 0.110256
R7712 VSS.n396 VSS.n393 0.110256
R7713 VSS.n399 VSS.n396 0.110256
R7714 VSS.n402 VSS.n399 0.110256
R7715 VSS.n405 VSS.n402 0.110256
R7716 VSS.n412 VSS.n409 0.110256
R7717 VSS.n419 VSS.n416 0.110256
R7718 VSS.n422 VSS.n419 0.110256
R7719 VSS.n427 VSS.n422 0.110256
R7720 VSS.n430 VSS.n427 0.110256
R7721 VSS.n433 VSS.n430 0.110256
R7722 VSS.n436 VSS.n433 0.110256
R7723 VSS.n439 VSS.n436 0.110256
R7724 VSS.n442 VSS.n439 0.110256
R7725 VSS.n445 VSS.n442 0.110256
R7726 VSS.n448 VSS.n445 0.110256
R7727 VSS.n451 VSS.n448 0.110256
R7728 VSS.n454 VSS.n451 0.110256
R7729 VSS.n458 VSS.n454 0.110256
R7730 VSS.n461 VSS.n458 0.110256
R7731 VSS.n464 VSS.n461 0.110256
R7732 VSS.n473 VSS.n464 0.110256
R7733 VSS.n476 VSS.n473 0.110256
R7734 VSS.n479 VSS.n476 0.110256
R7735 VSS.n482 VSS.n479 0.110256
R7736 VSS.n485 VSS.n482 0.110256
R7737 VSS.n1534 VSS.n1531 0.110256
R7738 VSS.n1531 VSS.n1528 0.110256
R7739 VSS.n4037 VSS.n4034 0.110256
R7740 VSS.n3976 VSS.n3973 0.110256
R7741 VSS.n3973 VSS.n3970 0.110256
R7742 VSS.n3970 VSS.n3967 0.110256
R7743 VSS.n3967 VSS.n3964 0.110256
R7744 VSS.n3964 VSS.n3961 0.110256
R7745 VSS.n3961 VSS.n3958 0.110256
R7746 VSS.n3958 VSS.n3955 0.110256
R7747 VSS.n3955 VSS.n3952 0.110256
R7748 VSS.n3952 VSS.n3949 0.110256
R7749 VSS.n3949 VSS.n3946 0.110256
R7750 VSS.n3946 VSS.n3943 0.110256
R7751 VSS.n3943 VSS.n3940 0.110256
R7752 VSS.n3940 VSS.n3937 0.110256
R7753 VSS.n3937 VSS.n3934 0.110256
R7754 VSS.n3934 VSS.n3930 0.110256
R7755 VSS.n3930 VSS.n3927 0.110256
R7756 VSS.n3927 VSS.n3924 0.110256
R7757 VSS.n3924 VSS.n3921 0.110256
R7758 VSS.n3921 VSS.n3918 0.110256
R7759 VSS.n4046 VSS.n4042 0.110256
R7760 VSS.n4049 VSS.n4046 0.110256
R7761 VSS.n4057 VSS.n4053 0.110256
R7762 VSS.n4060 VSS.n4057 0.110256
R7763 VSS.n4063 VSS.n4060 0.110256
R7764 VSS.n728 VSS.n725 0.110256
R7765 VSS.n725 VSS.n722 0.110256
R7766 VSS.n722 VSS.n719 0.110256
R7767 VSS.n4280 VSS.n4278 0.110256
R7768 VSS.n4283 VSS.n4280 0.110256
R7769 VSS.n4286 VSS.n4283 0.110256
R7770 VSS.n4298 VSS.n4295 0.110256
R7771 VSS.n4295 VSS.n4292 0.110256
R7772 VSS.n4292 VSS.n4289 0.110256
R7773 VSS.n907 VSS.n905 0.110256
R7774 VSS.n905 VSS.n902 0.110256
R7775 VSS.n902 VSS.n899 0.110256
R7776 VSS.n899 VSS.n897 0.110256
R7777 VSS.n897 VSS.n895 0.110256
R7778 VSS.n895 VSS.n893 0.110256
R7779 VSS.n4226 VSS.n4223 0.110256
R7780 VSS.n4229 VSS.n4226 0.110256
R7781 VSS.n4232 VSS.n4229 0.110256
R7782 VSS.n4234 VSS.n4232 0.110256
R7783 VSS.n4237 VSS.n4234 0.110256
R7784 VSS.n4241 VSS.n4237 0.110256
R7785 VSS.n4244 VSS.n4241 0.110256
R7786 VSS.n4247 VSS.n4244 0.110256
R7787 VSS.n4251 VSS.n4247 0.110256
R7788 VSS.n4258 VSS.n4255 0.110256
R7789 VSS.n4261 VSS.n4258 0.110256
R7790 VSS.n4264 VSS.n4261 0.110256
R7791 VSS.n4267 VSS.n4264 0.110256
R7792 VSS.n4270 VSS.n4267 0.110256
R7793 VSS.n5807 VSS.n5806 0.110211
R7794 VSS.n243 VSS.n242 0.109357
R7795 VSS.n5253 VSS.n5252 0.109357
R7796 VSS.n6075 VSS 0.109087
R7797 VSS.n5276 VSS.n5275 0.108345
R7798 VSS.n5322 VSS.n5321 0.10833
R7799 VSS.n5298 VSS.n5297 0.10833
R7800 VSS.n4378 VSS.n4377 0.10833
R7801 VSS.n4409 VSS.n4408 0.10833
R7802 VSS.n4492 VSS.n4489 0.108109
R7803 VSS.n5537 VSS.n5534 0.108109
R7804 VSS.n4050 VSS.n4049 0.108061
R7805 VSS.n498 VSS.n497 0.108061
R7806 VSS.n1336 VSS.n1333 0.107895
R7807 VSS.n5304 VSS.n5303 0.10713
R7808 VSS.n5463 VSS.n5460 0.107079
R7809 VSS VSS.n358 0.107055
R7810 VSS.n4990 VSS.n4987 0.106429
R7811 VSS.n4299 VSS.n4298 0.105134
R7812 VSS.n5439 VSS.n5436 0.104711
R7813 VSS.n4439 VSS.n4436 0.104711
R7814 VSS.n252 VSS.n251 0.104196
R7815 VSS.n5267 VSS.n5264 0.104196
R7816 VSS.n5880 VSS 0.103833
R7817 VSS VSS.n5799 0.103833
R7818 VSS VSS.n5817 0.103833
R7819 VSS.n5120 VSS.n5118 0.10383
R7820 VSS.n4597 VSS.n4594 0.103507
R7821 VSS.n5920 VSS 0.10345
R7822 VSS.n4611 VSS.n4609 0.103243
R7823 VSS.n5155 VSS.n5152 0.103217
R7824 VSS.n154 VSS.n151 0.103217
R7825 VSS.n4118 VSS.n4099 0.102601
R7826 VSS.n5146 VSS.n5062 0.102447
R7827 VSS.n4986 VSS.n4983 0.102447
R7828 VSS.n5152 VSS.n5149 0.102239
R7829 VSS.n5158 VSS.n5155 0.102239
R7830 VSS.n157 VSS.n154 0.102239
R7831 VSS.n151 VSS.n62 0.102239
R7832 VSS.n3846 VSS.n3845 0.100173
R7833 VSS.n187 VSS.n184 0.0999444
R7834 VSS.n240 VSS.n123 0.0999444
R7835 VSS.n5197 VSS.n5194 0.0999444
R7836 VSS.n5249 VSS.n5248 0.0999444
R7837 VSS VSS.n5850 0.0997784
R7838 VSS.n5933 VSS 0.0997784
R7839 VSS VSS.n5774 0.0997784
R7840 VSS.n4585 VSS.n4582 0.0992611
R7841 VSS.n4382 VSS.n4381 0.0990345
R7842 VSS.n5274 VSS.n5273 0.0990345
R7843 VSS.n96 VSS.n95 0.0986818
R7844 VSS.n5095 VSS.n5092 0.0984646
R7845 VSS.n5083 VSS.n5076 0.0978681
R7846 VSS.n5023 VSS.n5020 0.0974231
R7847 VSS.n5030 VSS.n5027 0.0974231
R7848 VSS.n5033 VSS.n5030 0.0974231
R7849 VSS.n4644 VSS.n4641 0.0974231
R7850 VSS.n4647 VSS.n4644 0.0974231
R7851 VSS.n4653 VSS.n4650 0.0974231
R7852 VSS.n5427 VSS.n5426 0.0973478
R7853 VSS.n1165 VSS.n1164 0.0968905
R7854 VSS.n5027 VSS.n5023 0.0964341
R7855 VSS.n4650 VSS.n4647 0.0964341
R7856 VSS.n5307 VSS.n5304 0.0963696
R7857 VSS.n3915 VSS.n1534 0.0956219
R7858 VSS.n4980 VSS.n4977 0.0952788
R7859 VSS.n51 VSS.n47 0.0952788
R7860 VSS.n5071 VSS.n5070 0.0945909
R7861 VSS VSS.n5874 0.0945618
R7862 VSS.n5270 VSS.n5254 0.0945541
R7863 VSS.n4497 VSS.n4492 0.0942929
R7864 VSS.n5540 VSS.n5537 0.0941041
R7865 VSS.n4119 VSS.n4118 0.09365
R7866 VSS.n5252 VSS.n5251 0.0922143
R7867 VSS.n4561 VSS.n4560 0.0920929
R7868 VSS.n1031 VSS.n1030 0.0914091
R7869 VSS VSS.n0 0.0914091
R7870 VSS VSS.n6106 0.0914091
R7871 VSS.n6106 VSS.n6105 0.0914091
R7872 VSS.n6105 VSS.n6104 0.0914091
R7873 VSS.n6100 VSS.n6099 0.0914091
R7874 VSS.n242 VSS.n241 0.0913571
R7875 VSS.n1284 VSS.n1283 0.09125
R7876 VSS.n1024 VSS.n1012 0.0909545
R7877 VSS.n321 VSS.n320 0.0907679
R7878 VSS.n252 VSS.n109 0.0905
R7879 VSS.n5264 VSS.n5259 0.0905
R7880 VSS.n4995 VSS.n4994 0.0905
R7881 VSS.n4419 VSS.n4418 0.0905
R7882 VSS.n4677 VSS.n4674 0.0905
R7883 VSS.n4073 VSS.n908 0.0897683
R7884 VSS.n4042 VSS.n4040 0.0897683
R7885 VSS.n5149 VSS.n5146 0.0895217
R7886 VSS.n5140 VSS.n5139 0.0889071
R7887 VSS.n4609 VSS.n62 0.0885435
R7888 VSS.n4601 VSS.n4600 0.0881106
R7889 VSS.n5868 VSS.n5867 0.0877209
R7890 VSS.n5543 VSS.n5540 0.0873421
R7891 VSS.n4500 VSS.n4497 0.0873421
R7892 VSS.n1452 VSS.n1451 0.0862944
R7893 VSS.n1449 VSS.n1448 0.0862944
R7894 VSS.n5379 VSS.n5376 0.0854057
R7895 VSS.n5382 VSS.n5379 0.0854057
R7896 VSS.n5385 VSS.n5382 0.0854057
R7897 VSS.n5388 VSS.n5385 0.0854057
R7898 VSS.n5391 VSS.n5388 0.0854057
R7899 VSS.n5394 VSS.n5391 0.0854057
R7900 VSS.n5397 VSS.n5394 0.0854057
R7901 VSS.n5400 VSS.n5397 0.0854057
R7902 VSS.n5403 VSS.n5400 0.0854057
R7903 VSS.n5406 VSS.n5403 0.0854057
R7904 VSS.n5409 VSS.n5406 0.0854057
R7905 VSS.n5412 VSS.n5409 0.0854057
R7906 VSS.n5415 VSS.n5412 0.0854057
R7907 VSS.n5418 VSS.n5415 0.0854057
R7908 VSS.n5562 VSS.n5559 0.0854057
R7909 VSS.n5565 VSS.n5562 0.0854057
R7910 VSS.n5568 VSS.n5565 0.0854057
R7911 VSS.n5571 VSS.n5568 0.0854057
R7912 VSS.n5578 VSS.n5575 0.0854057
R7913 VSS.n5581 VSS.n5578 0.0854057
R7914 VSS.n5584 VSS.n5581 0.0854057
R7915 VSS.n5586 VSS.n5584 0.0854057
R7916 VSS.n5594 VSS.n5590 0.0854057
R7917 VSS.n5597 VSS.n5594 0.0854057
R7918 VSS.n5600 VSS.n5597 0.0854057
R7919 VSS.n5603 VSS.n5600 0.0854057
R7920 VSS.n5606 VSS.n5603 0.0854057
R7921 VSS.n5613 VSS.n5610 0.0854057
R7922 VSS.n5616 VSS.n5613 0.0854057
R7923 VSS.n1032 VSS.n1031 0.0850455
R7924 VSS.n4360 VSS.n4358 0.0846795
R7925 VSS.n5279 VSS.n5276 0.0846304
R7926 VSS.n5376 VSS.n5373 0.0843639
R7927 VSS.n4560 VSS.n4558 0.0841283
R7928 VSS.n39 VSS.n38 0.0841283
R7929 VSS.n5112 VSS.n5095 0.0838349
R7930 VSS.n4777 VSS.n4776 0.0838333
R7931 VSS.n5115 VSS.n5114 0.0837469
R7932 VSS.n4590 VSS.n4589 0.0832732
R7933 VSS.n5480 VSS.n5476 0.0832014
R7934 VSS.n5373 VSS.n5370 0.0830864
R7935 VSS VSS.n5914 0.083054
R7936 VSS.n4586 VSS.n4585 0.0830384
R7937 VSS.n4345 VSS.n4343 0.0828171
R7938 VSS.n1161 VSS.n1158 0.0828171
R7939 VSS.n1158 VSS.n1155 0.0828171
R7940 VSS.n1155 VSS.n1152 0.0828171
R7941 VSS.n1152 VSS.n1149 0.0828171
R7942 VSS.n1149 VSS.n1146 0.0828171
R7943 VSS.n1146 VSS.n1143 0.0828171
R7944 VSS.n1143 VSS.n1140 0.0828171
R7945 VSS.n1140 VSS.n1137 0.0828171
R7946 VSS.n1137 VSS.n1134 0.0828171
R7947 VSS.n1134 VSS.n1131 0.0828171
R7948 VSS.n1131 VSS.n1128 0.0828171
R7949 VSS.n1128 VSS.n1125 0.0828171
R7950 VSS.n1125 VSS.n1122 0.0828171
R7951 VSS.n1122 VSS.n1119 0.0828171
R7952 VSS.n1119 VSS.n1116 0.0828171
R7953 VSS.n1116 VSS.n1113 0.0828171
R7954 VSS.n1113 VSS.n1110 0.0828171
R7955 VSS.n1110 VSS.n1107 0.0828171
R7956 VSS.n1107 VSS.n1104 0.0828171
R7957 VSS.n1104 VSS.n1101 0.0828171
R7958 VSS.n1101 VSS.n1098 0.0828171
R7959 VSS.n1098 VSS.n1095 0.0828171
R7960 VSS.n1095 VSS.n1092 0.0828171
R7961 VSS.n1092 VSS.n1089 0.0828171
R7962 VSS.n1089 VSS.n1086 0.0828171
R7963 VSS.n1086 VSS.n1083 0.0828171
R7964 VSS.n1083 VSS.n1080 0.0828171
R7965 VSS.n1080 VSS.n1076 0.0828171
R7966 VSS.n1076 VSS.n1073 0.0828171
R7967 VSS.n1073 VSS.n1070 0.0828171
R7968 VSS.n1070 VSS.n1067 0.0828171
R7969 VSS.n1067 VSS.n1064 0.0828171
R7970 VSS.n1064 VSS.n1061 0.0828171
R7971 VSS.n1061 VSS.n1058 0.0828171
R7972 VSS.n1058 VSS.n1055 0.0828171
R7973 VSS.n1055 VSS.n1052 0.0828171
R7974 VSS.n1052 VSS.n1049 0.0828171
R7975 VSS.n1049 VSS.n1046 0.0828171
R7976 VSS.n1046 VSS.n1043 0.0828171
R7977 VSS.n1043 VSS.n1040 0.0828171
R7978 VSS.n1040 VSS.n1037 0.0828171
R7979 VSS.n713 VSS.n710 0.0828171
R7980 VSS.n710 VSS.n707 0.0828171
R7981 VSS.n707 VSS.n704 0.0828171
R7982 VSS.n700 VSS.n697 0.0828171
R7983 VSS.n697 VSS.n694 0.0828171
R7984 VSS.n691 VSS.n687 0.0828171
R7985 VSS.n685 VSS.n681 0.0828171
R7986 VSS.n681 VSS.n678 0.0828171
R7987 VSS.n678 VSS.n675 0.0828171
R7988 VSS.n675 VSS.n673 0.0828171
R7989 VSS.n673 VSS.n670 0.0828171
R7990 VSS.n670 VSS.n667 0.0828171
R7991 VSS.n667 VSS.n664 0.0828171
R7992 VSS.n664 VSS.n661 0.0828171
R7993 VSS.n661 VSS.n658 0.0828171
R7994 VSS.n658 VSS.n655 0.0828171
R7995 VSS.n655 VSS.n652 0.0828171
R7996 VSS.n652 VSS.n649 0.0828171
R7997 VSS.n649 VSS.n646 0.0828171
R7998 VSS.n646 VSS.n643 0.0828171
R7999 VSS.n643 VSS.n640 0.0828171
R8000 VSS.n640 VSS.n637 0.0828171
R8001 VSS.n637 VSS.n634 0.0828171
R8002 VSS.n634 VSS.n631 0.0828171
R8003 VSS.n631 VSS.n628 0.0828171
R8004 VSS.n628 VSS.n625 0.0828171
R8005 VSS.n625 VSS.n622 0.0828171
R8006 VSS.n622 VSS.n619 0.0828171
R8007 VSS.n619 VSS.n616 0.0828171
R8008 VSS.n616 VSS.n613 0.0828171
R8009 VSS.n613 VSS.n610 0.0828171
R8010 VSS.n610 VSS.n607 0.0828171
R8011 VSS.n607 VSS.n604 0.0828171
R8012 VSS.n604 VSS.n601 0.0828171
R8013 VSS.n601 VSS.n598 0.0828171
R8014 VSS.n598 VSS.n595 0.0828171
R8015 VSS.n595 VSS.n593 0.0828171
R8016 VSS.n593 VSS.n589 0.0828171
R8017 VSS.n589 VSS.n586 0.0828171
R8018 VSS.n586 VSS.n583 0.0828171
R8019 VSS.n583 VSS.n580 0.0828171
R8020 VSS.n580 VSS.n577 0.0828171
R8021 VSS.n577 VSS.n574 0.0828171
R8022 VSS.n574 VSS.n571 0.0828171
R8023 VSS.n571 VSS.n566 0.0828171
R8024 VSS.n566 VSS.n562 0.0828171
R8025 VSS.n562 VSS.n559 0.0828171
R8026 VSS.n559 VSS.n556 0.0828171
R8027 VSS.n556 VSS.n554 0.0828171
R8028 VSS.n554 VSS.n551 0.0828171
R8029 VSS.n551 VSS.n548 0.0828171
R8030 VSS.n548 VSS.n545 0.0828171
R8031 VSS.n545 VSS.n542 0.0828171
R8032 VSS.n542 VSS.n539 0.0828171
R8033 VSS.n539 VSS.n536 0.0828171
R8034 VSS.n536 VSS.n533 0.0828171
R8035 VSS.n533 VSS.n530 0.0828171
R8036 VSS.n530 VSS.n526 0.0828171
R8037 VSS.n526 VSS.n523 0.0828171
R8038 VSS.n523 VSS.n520 0.0828171
R8039 VSS.n520 VSS.n517 0.0828171
R8040 VSS.n517 VSS.n514 0.0828171
R8041 VSS.n5338 VSS.n5334 0.0828171
R8042 VSS.n5341 VSS.n5338 0.0828171
R8043 VSS.n5343 VSS.n5341 0.0828171
R8044 VSS.n5346 VSS.n5343 0.0828171
R8045 VSS.n5349 VSS.n5346 0.0828171
R8046 VSS.n5353 VSS.n5349 0.0828171
R8047 VSS.n5358 VSS.n5353 0.0828171
R8048 VSS.n5361 VSS.n5358 0.0828171
R8049 VSS.n5364 VSS.n5361 0.0828171
R8050 VSS.n5367 VSS.n5364 0.0828171
R8051 VSS.n5370 VSS.n5367 0.0828171
R8052 VSS.n787 VSS.n784 0.0828171
R8053 VSS.n784 VSS.n781 0.0828171
R8054 VSS.n781 VSS.n778 0.0828171
R8055 VSS.n778 VSS.n775 0.0828171
R8056 VSS.n751 VSS.n748 0.0828171
R8057 VSS.n748 VSS.n745 0.0828171
R8058 VSS.n745 VSS.n742 0.0828171
R8059 VSS.n742 VSS.n739 0.0828171
R8060 VSS.n992 VSS.n988 0.0828171
R8061 VSS.n988 VSS.n985 0.0828171
R8062 VSS.n985 VSS.n983 0.0828171
R8063 VSS.n983 VSS.n980 0.0828171
R8064 VSS.n980 VSS.n976 0.0828171
R8065 VSS.n976 VSS.n99 0.0828171
R8066 VSS.n4354 VSS.n4351 0.0828171
R8067 VSS.n4351 VSS.n4349 0.0828171
R8068 VSS.n4349 VSS.n4345 0.0828171
R8069 VSS.n4343 VSS.n4340 0.0828171
R8070 VSS.n4340 VSS.n4337 0.0828171
R8071 VSS.n4334 VSS.n4330 0.0828171
R8072 VSS.n4327 VSS.n4324 0.0828171
R8073 VSS.n4324 VSS.n4321 0.0828171
R8074 VSS.n4321 VSS.n4319 0.0828171
R8075 VSS.n4319 VSS.n4315 0.0828171
R8076 VSS.n1008 VSS.n1005 0.0828171
R8077 VSS.n1005 VSS.n1002 0.0828171
R8078 VSS.n1002 VSS.n998 0.0828171
R8079 VSS.n998 VSS.n995 0.0828171
R8080 VSS.n15 VSS.n5 0.0828171
R8081 VSS.n15 VSS.n14 0.0828171
R8082 VSS.n14 VSS.n11 0.0828171
R8083 VSS.n11 VSS.n8 0.0828171
R8084 VSS.n6091 VSS.n6090 0.0828171
R8085 VSS.n6090 VSS.n6087 0.0828171
R8086 VSS.n6087 VSS.n6084 0.0828171
R8087 VSS.n6084 VSS.n6081 0.0828171
R8088 VSS.n6081 VSS.n6078 0.0828171
R8089 VSS.n6074 VSS.n6070 0.0828171
R8090 VSS.n6070 VSS.n6067 0.0828171
R8091 VSS.n6067 VSS.n6061 0.0828171
R8092 VSS.n6061 VSS.n6057 0.0828171
R8093 VSS.n6057 VSS.n6054 0.0828171
R8094 VSS.n6054 VSS.n6051 0.0828171
R8095 VSS.n6051 VSS.n6048 0.0828171
R8096 VSS.n6048 VSS.n6045 0.0828171
R8097 VSS.n6045 VSS.n6043 0.0828171
R8098 VSS.n6043 VSS.n6040 0.0828171
R8099 VSS.n6040 VSS.n6036 0.0828171
R8100 VSS.n6036 VSS.n6033 0.0828171
R8101 VSS.n6033 VSS.n6030 0.0828171
R8102 VSS.n6030 VSS.n6027 0.0828171
R8103 VSS.n6027 VSS.n6025 0.0828171
R8104 VSS.n6025 VSS.n6022 0.0828171
R8105 VSS.n6022 VSS.n6017 0.0828171
R8106 VSS.n6017 VSS.n6014 0.0828171
R8107 VSS.n6014 VSS.n6012 0.0828171
R8108 VSS.n6012 VSS.n6009 0.0828171
R8109 VSS.n6009 VSS.n6005 0.0828171
R8110 VSS.n6005 VSS.n6003 0.0828171
R8111 VSS.n6003 VSS.n6000 0.0828171
R8112 VSS.n6000 VSS.n5998 0.0828171
R8113 VSS.n5998 VSS.n5995 0.0828171
R8114 VSS.n5995 VSS.n5993 0.0828171
R8115 VSS.n5993 VSS.n5991 0.0828171
R8116 VSS.n5991 VSS.n5987 0.0828171
R8117 VSS.n5987 VSS.n5983 0.0828171
R8118 VSS.n5983 VSS.n5980 0.0828171
R8119 VSS.n5980 VSS.n5977 0.0828171
R8120 VSS.n5977 VSS.n5974 0.0828171
R8121 VSS.n5974 VSS.n5971 0.0828171
R8122 VSS.n5971 VSS.n5968 0.0828171
R8123 VSS.n5968 VSS.n5965 0.0828171
R8124 VSS.n5965 VSS.n5962 0.0828171
R8125 VSS.n5962 VSS.n5959 0.0828171
R8126 VSS.n5959 VSS.n5956 0.0828171
R8127 VSS.n5956 VSS.n5953 0.0828171
R8128 VSS.n5953 VSS.n5950 0.0828171
R8129 VSS.n5950 VSS.n5947 0.0828171
R8130 VSS.n5947 VSS.n5944 0.0828171
R8131 VSS.n5944 VSS.n5941 0.0828171
R8132 VSS.n4766 VSS.n4741 0.0828171
R8133 VSS.n4769 VSS.n4766 0.0828171
R8134 VSS.n5731 VSS.n4769 0.0828171
R8135 VSS.n5731 VSS.n5730 0.0828171
R8136 VSS.n5730 VSS.n5727 0.0828171
R8137 VSS.n5727 VSS.n5724 0.0828171
R8138 VSS.n5724 VSS.n5721 0.0828171
R8139 VSS.n5721 VSS.n5718 0.0828171
R8140 VSS.n5718 VSS.n5715 0.0828171
R8141 VSS.n5715 VSS.n5712 0.0828171
R8142 VSS.n5712 VSS.n5708 0.0828171
R8143 VSS.n5708 VSS.n5705 0.0828171
R8144 VSS.n5705 VSS.n5702 0.0828171
R8145 VSS.n5702 VSS.n5699 0.0828171
R8146 VSS.n5699 VSS.n5696 0.0828171
R8147 VSS.n5696 VSS.n5693 0.0828171
R8148 VSS.n5693 VSS.n5690 0.0828171
R8149 VSS.n5690 VSS.n5687 0.0828171
R8150 VSS.n5687 VSS.n5680 0.0828171
R8151 VSS.n5680 VSS.n5677 0.0828171
R8152 VSS.n5677 VSS.n5672 0.0828171
R8153 VSS.n5672 VSS.n5669 0.0828171
R8154 VSS.n5669 VSS.n5667 0.0828171
R8155 VSS.n5663 VSS.n5660 0.0828171
R8156 VSS.n5660 VSS.n5658 0.0828171
R8157 VSS.n5658 VSS.n5655 0.0828171
R8158 VSS.n5655 VSS.n5653 0.0828171
R8159 VSS.n5649 VSS.n5647 0.0828171
R8160 VSS.n5647 VSS.n5644 0.0828171
R8161 VSS.n5644 VSS.n5641 0.0828171
R8162 VSS.n5641 VSS.n5639 0.0828171
R8163 VSS.n5639 VSS.n5636 0.0828171
R8164 VSS.n5632 VSS.n5629 0.0828171
R8165 VSS.n5629 VSS.n5626 0.0828171
R8166 VSS.n5626 VSS.n5624 0.0828171
R8167 VSS.n5624 VSS.n5622 0.0828171
R8168 VSS.n5426 VSS.n5423 0.0826739
R8169 VSS.n4600 VSS.n4598 0.082242
R8170 VSS.n704 VSS.n701 0.0817195
R8171 VSS.n188 VSS.n167 0.0816957
R8172 VSS.n271 VSS.n270 0.0816607
R8173 VSS.n4889 VSS.n4888 0.0815383
R8174 VSS.n5139 VSS.n5133 0.0814455
R8175 VSS.n6078 VSS.n6075 0.0811707
R8176 VSS.n5089 VSS.n5088 0.0809425
R8177 VSS.n955 VSS.n954 0.0808571
R8178 VSS.n4132 VSS.n4130 0.0808571
R8179 VSS.n4219 VSS.n4207 0.0808571
R8180 VSS.n5198 VSS.n5177 0.0807174
R8181 VSS.n4328 VSS 0.0803113
R8182 VSS.n4501 VSS.n4500 0.0802368
R8183 VSS.n4579 VSS.n4578 0.080146
R8184 VSS.n307 VSS.n306 0.079766
R8185 VSS.n5548 VSS.n5543 0.0794474
R8186 VSS.n313 VSS.n312 0.0794283
R8187 VSS VSS.n950 0.07925
R8188 VSS.n5912 VSS.n4746 0.0790301
R8189 VSS.n4040 VSS.n4037 0.0787927
R8190 VSS.n5936 VSS.n4741 0.0784268
R8191 VSS.n5007 VSS.n5006 0.0777566
R8192 VSS.n4064 VSS.n4063 0.0773293
R8193 VSS.n84 VSS.n83 0.0770957
R8194 VSS.n5105 VSS.n5104 0.0770957
R8195 VSS.n5555 VSS.n5472 0.077079
R8196 VSS.n4666 VSS.n4664 0.0769602
R8197 VSS.n5587 VSS.n5586 0.0769151
R8198 VSS.n5479 VSS.n5477 0.076587
R8199 VSS.n5892 VSS.n5891 0.0763268
R8200 VSS.n4328 VSS.n4327 0.0762317
R8201 VSS.n4092 VSS 0.0760357
R8202 VSS.n4130 VSS 0.0760357
R8203 VSS.n908 VSS.n907 0.0758658
R8204 VSS.n5238 VSS.n5235 0.0758261
R8205 VSS.n1333 VSS.n938 0.0755
R8206 VSS VSS.n955 0.0752321
R8207 VSS.n882 VSS.n879 0.0752
R8208 VSS.n205 VSS.n204 0.0748478
R8209 VSS.n5622 VSS.n5619 0.0745854
R8210 VSS.n5890 VSS.n5889 0.0744082
R8211 VSS VSS.n5463 0.0739211
R8212 VSS.n5270 VSS.n5269 0.0738696
R8213 VSS VSS.n4467 0.0731316
R8214 VSS.n276 VSS.n275 0.0728214
R8215 VSS.n4681 VSS.n57 0.0721814
R8216 VSS.n1304 VSS.n1302 0.0715924
R8217 VSS.n4575 VSS.n4571 0.071385
R8218 VSS.n5837 VSS.n5836 0.0712072
R8219 VSS.n5835 VSS.n5834 0.0711439
R8220 VSS.n5788 VSS 0.0710963
R8221 VSS.n6102 VSS.n6101 0.0709545
R8222 VSS.n4991 VSS.n4990 0.0705885
R8223 VSS.n337 VSS.n333 0.0704107
R8224 VSS.n360 VSS.n359 0.0704107
R8225 VSS.n4219 VSS.n4218 0.0704107
R8226 VSS.n3977 VSS.n3976 0.0700122
R8227 VSS.n4299 VSS.n4286 0.0700122
R8228 VSS VSS.n5929 0.0696579
R8229 VSS.n5633 VSS.n5632 0.0696463
R8230 VSS.n4508 VSS.n4507 0.0687418
R8231 VSS.n5075 VSS.n5074 0.0687418
R8232 VSS.n4118 VSS.n1340 0.0685672
R8233 VSS.n3918 VSS.n3915 0.0685488
R8234 VSS.n5653 VSS.n5650 0.0685488
R8235 VSS.n5919 VSS.n5915 0.068
R8236 VSS.n5922 VSS.n4749 0.068
R8237 VSS.n5787 VSS.n5783 0.068
R8238 VSS.n5840 VSS.n5839 0.068
R8239 VSS.n1309 VSS.n1308 0.0678109
R8240 VSS.n5555 VSS.n5554 0.0676053
R8241 VSS.n75 VSS.n66 0.0675213
R8242 VSS.n5132 VSS.n5123 0.0675213
R8243 VSS.n5440 VSS.n5439 0.0673304
R8244 VSS.n4440 VSS.n4439 0.067297
R8245 VSS.n5534 VSS.n5531 0.0670217
R8246 VSS.n92 VSS.n91 0.0666326
R8247 VSS.n5110 VSS.n5109 0.0661354
R8248 VSS.n4093 VSS.n4092 0.0656429
R8249 VSS.n4278 VSS.n4276 0.0656219
R8250 VSS.n5559 VSS.n5556 0.0655943
R8251 VSS.n5610 VSS.n5607 0.0655943
R8252 VSS.n74 VSS.n73 0.0649262
R8253 VSS.n5131 VSS.n5130 0.0644344
R8254 VSS.n87 VSS.n86 0.0640294
R8255 VSS.n4096 VSS.n4093 0.0640294
R8256 VSS.n1309 VSS.n955 0.0639286
R8257 VSS.n5848 VSS.n5847 0.0636651
R8258 VSS.n5111 VSS.n5110 0.0636492
R8259 VSS.n93 VSS.n92 0.0636492
R8260 VSS.n5076 VSS.n5075 0.0633022
R8261 VSS.n4509 VSS.n4508 0.0633022
R8262 VSS.n75 VSS.n74 0.062959
R8263 VSS.n5132 VSS.n5131 0.062959
R8264 VSS.n729 VSS.n728 0.0626951
R8265 VSS.n5104 VSS.n5103 0.0622838
R8266 VSS.n83 VSS.n82 0.0622838
R8267 VSS.n4411 VSS.n4391 0.0621304
R8268 VSS.n5282 VSS.n5281 0.0618391
R8269 VSS.n5879 VSS.n4758 0.0616111
R8270 VSS.n5802 VSS.n5801 0.0616111
R8271 VSS.n5819 VSS.n5818 0.0616111
R8272 VSS.n310 VSS.n309 0.0616009
R8273 VSS.n302 VSS.n301 0.0616009
R8274 VSS.n4571 VSS.n4509 0.0613736
R8275 VSS.n208 VSS.n205 0.0611522
R8276 VSS.n4252 VSS.n4251 0.0605
R8277 VSS.n5174 VSS.n5171 0.0603902
R8278 VSS.n5235 VSS.n5234 0.0601739
R8279 VSS.n929 VSS.n926 0.0596608
R8280 VSS.n931 VSS.n929 0.0596608
R8281 VSS.n932 VSS.n931 0.0596608
R8282 VSS.n937 VSS 0.0596608
R8283 VSS.n945 VSS.n942 0.0596608
R8284 VSS.n947 VSS.n945 0.0596608
R8285 VSS.n4866 VSS.n4863 0.0596608
R8286 VSS.n4869 VSS.n4866 0.0596608
R8287 VSS.n4870 VSS.n4869 0.0596608
R8288 VSS VSS.n4870 0.0596608
R8289 VSS.n4878 VSS.n4875 0.0596608
R8290 VSS.n4881 VSS.n4878 0.0596608
R8291 VSS.n4884 VSS.n4881 0.0596608
R8292 VSS.n4828 VSS.n4825 0.0596608
R8293 VSS.n4831 VSS.n4828 0.0596608
R8294 VSS.n4832 VSS.n4831 0.0596608
R8295 VSS VSS.n4832 0.0596608
R8296 VSS.n4840 VSS.n4837 0.0596608
R8297 VSS.n4843 VSS.n4840 0.0596608
R8298 VSS.n4846 VSS.n4843 0.0596608
R8299 VSS.n4900 VSS.n4897 0.0596608
R8300 VSS.n4903 VSS.n4900 0.0596608
R8301 VSS.n4904 VSS.n4903 0.0596608
R8302 VSS VSS.n4904 0.0596608
R8303 VSS.n4912 VSS.n4909 0.0596608
R8304 VSS.n4917 VSS.n4912 0.0596608
R8305 VSS.n4920 VSS.n4917 0.0596608
R8306 VSS.n4941 VSS.n4938 0.0596608
R8307 VSS.n4944 VSS.n4941 0.0596608
R8308 VSS.n4945 VSS.n4944 0.0596608
R8309 VSS VSS.n4945 0.0596608
R8310 VSS.n4953 VSS.n4950 0.0596608
R8311 VSS.n4956 VSS.n4953 0.0596608
R8312 VSS.n4959 VSS.n4956 0.0596608
R8313 VSS.n4143 VSS.n4140 0.0596608
R8314 VSS.n4145 VSS.n4143 0.0596608
R8315 VSS.n164 VSS.n161 0.0594119
R8316 VSS.n5888 VSS.n5887 0.0587734
R8317 VSS.n4753 VSS.n4752 0.0584651
R8318 VSS.n767 VSS.n763 0.0583049
R8319 VSS.n5833 VSS.n5832 0.0581418
R8320 VSS.n4020 VSS.n4019 0.0574719
R8321 VSS.n4422 VSS.n4419 0.0572391
R8322 VSS.n5885 VSS.n5884 0.0571667
R8323 VSS.n5824 VSS.n5823 0.0570217
R8324 VSS.n5020 VSS.n5017 0.0568736
R8325 VSS.n4656 VSS.n4653 0.0568736
R8326 VSS.n5619 VSS.n5616 0.0559717
R8327 VSS.n406 VSS.n405 0.055378
R8328 VSS.n409 VSS.n406 0.055378
R8329 VSS.n413 VSS.n412 0.055378
R8330 VSS.n416 VSS.n413 0.055378
R8331 VSS.n5201 VSS.n5198 0.0552826
R8332 VSS.n932 VSS.n922 0.0552552
R8333 VSS.n4875 VSS.n4853 0.0552552
R8334 VSS.n4837 VSS.n4816 0.0552552
R8335 VSS.n4909 VSS.n4810 0.0552552
R8336 VSS.n4950 VSS.n4928 0.0552552
R8337 VSS.n5894 VSS.n5893 0.0550669
R8338 VSS VSS.n218 0.0549444
R8339 VSS.n5224 VSS 0.0543889
R8340 VSS.n191 VSS.n188 0.0543043
R8341 VSS.n4008 VSS.n4007 0.0536953
R8342 VSS VSS.n4147 0.0533671
R8343 VSS.n4184 VSS.n4181 0.0533671
R8344 VSS.n4443 VSS.n4440 0.0530777
R8345 VSS.n5443 VSS.n5440 0.0530398
R8346 VSS.n1037 VSS.n1034 0.0526341
R8347 VSS.n4019 VSS.n4016 0.0521084
R8348 VSS.n4007 VSS.n4004 0.0521084
R8349 VSS.n5896 VSS.n5895 0.0515236
R8350 VSS.n5102 VSS.n5101 0.0514211
R8351 VSS.n4890 VSS.n4850 0.0513891
R8352 VSS.n5271 VSS.n4782 0.0513696
R8353 VSS.n4197 VSS.n4195 0.0508497
R8354 VSS.n4355 VSS.n99 0.050439
R8355 VSS.n4093 VSS.n1391 0.050416
R8356 VSS.n4255 VSS.n4252 0.0502561
R8357 VSS.n701 VSS.n700 0.0498902
R8358 VSS.n4335 VSS.n4334 0.0498902
R8359 VSS.n4994 VSS.n4991 0.0498805
R8360 VSS.n885 VSS.n884 0.0496753
R8361 VSS.n1030 VSS.n1029 0.0486818
R8362 VSS.n6099 VSS.n6098 0.0486818
R8363 VSS.n5572 VSS.n5571 0.0486132
R8364 VSS.n4030 VSS.n4027 0.0483322
R8365 VSS.n4757 VSS.n4756 0.0482778
R8366 VSS.n5821 VSS.n5820 0.0482778
R8367 VSS.n5813 VSS.n5812 0.0482778
R8368 VSS.n4313 VSS.n787 0.0476951
R8369 VSS.n5829 VSS.n5828 0.0474565
R8370 VSS.n1313 VSS.n1309 0.0466345
R8371 VSS.n4471 VSS 0.0462895
R8372 VSS VSS.n5221 0.0460556
R8373 VSS.n6104 VSS.n6103 0.0459545
R8374 VSS.n6103 VSS.n6102 0.0459545
R8375 VSS.n4276 VSS.n4270 0.0458659
R8376 VSS.n5809 VSS.n5808 0.0457506
R8377 VSS.n82 VSS.n81 0.0457432
R8378 VSS.n219 VSS 0.0455
R8379 VSS.n5466 VSS 0.0455
R8380 VSS.n5326 VSS.n5325 0.0455
R8381 VSS.n5103 VSS.n5102 0.0452568
R8382 VSS.n5847 VSS 0.0450872
R8383 VSS.n4755 VSS.n4754 0.044437
R8384 VSS.n73 VSS.n68 0.04425
R8385 VSS.n5130 VSS.n5125 0.04425
R8386 VSS.n1650 VSS.n1649 0.044243
R8387 VSS.n950 VSS.n948 0.0439266
R8388 VSS.n4894 VSS.n4893 0.0439266
R8389 VSS.n4935 VSS.n4934 0.0439266
R8390 VSS.n4138 VSS.n4137 0.0439266
R8391 VSS.n5264 VSS.n5263 0.0435435
R8392 VSS.n4664 VSS.n4663 0.0435088
R8393 VSS.n1029 VSS.n0 0.0432273
R8394 VSS.n1302 VSS.n1301 0.0428529
R8395 VSS.n5010 VSS.n5007 0.0427124
R8396 VSS.n89 VSS.n88 0.0426277
R8397 VSS.n1505 VSS.n1408 0.0425561
R8398 VSS.n5664 VSS.n5663 0.0422073
R8399 VSS.n5826 VSS.n5810 0.0413696
R8400 VSS.n5667 VSS.n5664 0.0411098
R8401 VSS.n1687 VSS.n1673 0.0404721
R8402 VSS.n4581 VSS.n4579 0.040323
R8403 VSS.n1523 VSS.n1522 0.0401503
R8404 VSS.n5091 VSS.n5089 0.0395266
R8405 VSS.n1034 VSS.n1008 0.0394634
R8406 VSS.n4389 VSS.n4386 0.0386522
R8407 VSS.n4067 VSS.n4064 0.0385488
R8408 VSS.n5805 VSS.n5804 0.0377928
R8409 VSS.n5791 VSS.n5789 0.037656
R8410 VSS.n938 VSS.n937 0.0376329
R8411 VSS.n5460 VSS.n5459 0.0376053
R8412 VSS.n5575 VSS.n5572 0.0372925
R8413 VSS.n6103 VSS.n21 0.0372105
R8414 VSS.n1564 VSS.n1563 0.0368785
R8415 VSS.n1568 VSS.n1567 0.0368564
R8416 VSS.n775 VSS.n774 0.0367195
R8417 VSS.n5326 VSS.n5279 0.0366957
R8418 VSS.n4969 VSS.n4966 0.0363407
R8419 VSS.n41 VSS.n39 0.0363407
R8420 VSS.n1404 VSS.n1403 0.0357448
R8421 VSS.n4375 VSS.n4374 0.0352779
R8422 VSS.n5295 VSS.n5294 0.0352465
R8423 VSS.n924 VSS.n919 0.0351154
R8424 VSS.n3981 VSS.n3980 0.0351154
R8425 VSS.n4888 VSS.n4885 0.0351154
R8426 VSS.n4850 VSS.n4847 0.0351154
R8427 VSS.n4924 VSS.n4921 0.0351154
R8428 VSS.n4963 VSS.n4960 0.0351154
R8429 VSS.n4185 VSS.n4184 0.0351154
R8430 VSS.n4201 VSS.n4198 0.0351154
R8431 VSS.n4681 VSS.n4680 0.0347478
R8432 VSS.n3994 VSS.n3993 0.034486
R8433 VSS.n4125 VSS.n912 0.0334464
R8434 VSS.n739 VSS.n736 0.0334268
R8435 VSS.n4337 VSS.n4335 0.0334268
R8436 VSS.n4570 VSS.n4569 0.0331549
R8437 VSS.n4355 VSS.n4354 0.032878
R8438 VSS.n4146 VSS.n4145 0.0325979
R8439 VSS.n4605 VSS.n4601 0.0323584
R8440 VSS.n3071 VSS.n1815 0.0323182
R8441 VSS.n1645 VSS.n1579 0.0320446
R8442 VSS.n1551 VSS.n1550 0.032
R8443 VSS.n1726 VSS.n1721 0.032
R8444 VSS.n1541 VSS.n1540 0.032
R8445 VSS.n4031 VSS.n4030 0.0319685
R8446 VSS.n4700 VSS.n4696 0.0318333
R8447 VSS.n4704 VSS.n4700 0.0318333
R8448 VSS.n4713 VSS.n4704 0.0318333
R8449 VSS.n4720 VSS 0.0318333
R8450 VSS.n4724 VSS.n4720 0.0318333
R8451 VSS.n4728 VSS.n4724 0.0318333
R8452 VSS.n4732 VSS.n4728 0.0318333
R8453 VSS.n5836 VSS.n5835 0.0315825
R8454 VSS.n5142 VSS.n5140 0.0315619
R8455 VSS.n1558 VSS.n1557 0.0309839
R8456 VSS.n314 VSS.n313 0.0305726
R8457 VSS.n1679 VSS.n1678 0.0302848
R8458 VSS.n4999 VSS.n4995 0.029969
R8459 VSS.n4674 VSS.n4673 0.029969
R8460 VSS.n1664 VSS.n1663 0.0299134
R8461 VSS.n4713 VSS.n4709 0.0295
R8462 VSS.n887 VSS.n886 0.0292629
R8463 VSS.n1586 VSS.n1585 0.0291175
R8464 VSS.n2439 VSS.n2429 0.0289279
R8465 VSS.n4153 VSS.n788 0.0288217
R8466 VSS.n966 VSS.n964 0.028625
R8467 VSS.n286 VSS.n283 0.028625
R8468 VSS.n330 VSS.n327 0.028625
R8469 VSS.n3506 VSS.n3500 0.028625
R8470 VSS.n4089 VSS.n4088 0.028625
R8471 VSS.n4126 VSS.n4125 0.028625
R8472 VSS.n4215 VSS.n4212 0.028625
R8473 VSS.n1165 VSS.n992 0.0284878
R8474 VSS.n872 VSS.n871 0.0284
R8475 VSS.n4564 VSS.n4561 0.0283761
R8476 VSS.n886 VSS.n885 0.0283351
R8477 VSS.n5766 VSS.n5757 0.0282695
R8478 VSS.n4031 VSS.n3984 0.0281923
R8479 VSS.n5447 VSS.n5444 0.0281316
R8480 VSS.n1613 VSS.n1612 0.0276659
R8481 VSS.n5080 VSS.n5078 0.0275796
R8482 VSS.n873 VSS.n872 0.0275
R8483 VSS.n1574 VSS.n1573 0.0274585
R8484 VSS.n79 VSS.n78 0.0273085
R8485 VSS.n5100 VSS.n5099 0.0273085
R8486 VSS.n253 VSS.n101 0.026913
R8487 VSS.n1677 VSS.n1676 0.0266
R8488 VSS.n1682 VSS.n1681 0.0266
R8489 VSS.n4370 VSS.n4369 0.0265939
R8490 VSS.n1502 VSS.n1409 0.0265748
R8491 VSS.n1448 VSS.n1447 0.0265748
R8492 VSS.n5792 VSS.n5791 0.0265092
R8493 VSS.n5789 VSS.n5788 0.0265092
R8494 VSS.n2803 VSS.n2082 0.0262358
R8495 VSS.n5291 VSS.n5289 0.0261799
R8496 VSS.n1899 VSS.n1898 0.0261034
R8497 VSS.n312 VSS.n311 0.0260963
R8498 VSS.n4368 VSS.n4367 0.0259717
R8499 VSS.n5288 VSS.n5287 0.0259717
R8500 VSS.n1703 VSS.n1702 0.0258911
R8501 VSS.n1446 VSS.n1445 0.0257336
R8502 VSS.n1447 VSS.n1408 0.0257336
R8503 VSS.n1547 VSS.n1546 0.0257
R8504 VSS.n1723 VSS.n1722 0.0257
R8505 VSS.n1537 VSS.n1536 0.0257
R8506 VSS.n1434 VSS.n1431 0.0256748
R8507 VSS.n1440 VSS.n1437 0.0256748
R8508 VSS.n1497 VSS.n1494 0.0256748
R8509 VSS.n1491 VSS.n1488 0.0256748
R8510 VSS.n806 VSS.n803 0.0256748
R8511 VSS.n812 VSS.n809 0.0256748
R8512 VSS.n818 VSS.n815 0.0256748
R8513 VSS.n846 VSS.n843 0.0256748
R8514 VSS.n853 VSS.n850 0.0256748
R8515 VSS.n1596 VSS.n1595 0.0255922
R8516 VSS.n2179 VSS.n2143 0.0254833
R8517 VSS.n1582 VSS.n1581 0.0253848
R8518 VSS.n2805 VSS.n2088 0.0253328
R8519 VSS.n2307 VSS.n2284 0.0253328
R8520 VSS.n311 VSS.n310 0.0252706
R8521 VSS.n308 VSS.n307 0.0252706
R8522 VSS.n4977 VSS.n4976 0.0251903
R8523 VSS.n47 VSS.n46 0.0251903
R8524 VSS.n2797 VSS.n2796 0.0251823
R8525 VSS.n1914 VSS.n1913 0.0251724
R8526 VSS.n926 VSS.n924 0.0250455
R8527 VSS.n1501 VSS.n1475 0.0250455
R8528 VSS.n3984 VSS.n3981 0.0250455
R8529 VSS.n4885 VSS.n4884 0.0250455
R8530 VSS.n4847 VSS.n4846 0.0250455
R8531 VSS.n4921 VSS.n4920 0.0250455
R8532 VSS.n4960 VSS.n4959 0.0250455
R8533 VSS.n4198 VSS.n4197 0.0250455
R8534 VSS.n2429 VSS.n2413 0.0249978
R8535 VSS.n1570 VSS 0.0247376
R8536 VSS.n820 VSS.n819 0.0247308
R8537 VSS.n5294 VSS.n5280 0.0247308
R8538 VSS.n335 VSS.n334 0.024574
R8539 VSS.n2808 VSS.n2807 0.0244298
R8540 VSS.n1811 VSS.n1810 0.0243636
R8541 VSS.n1625 VSS.n1624 0.0241406
R8542 VSS.n694 VSS.n691 0.0240976
R8543 VSS.n5941 VSS.n5938 0.0240976
R8544 VSS.n5430 VSS.n5427 0.0239783
R8545 VSS.n1806 VSS.n1805 0.0236818
R8546 VSS.n1808 VSS.n1804 0.0236818
R8547 VSS.n1606 VSS.n1605 0.0235184
R8548 VSS.n4738 VSS.n4733 0.0235
R8549 VSS.n5284 VSS.n5283 0.0234789
R8550 VSS.n3583 VSS.n3582 0.0233924
R8551 VSS.n161 VSS.n160 0.0232368
R8552 VSS VSS.n5869 0.0231603
R8553 VSS.n4364 VSS.n4363 0.0230525
R8554 VSS.n5271 VSS.n5270 0.023
R8555 VSS.n3505 VSS.n3504 0.0228692
R8556 VSS.n2956 VSS.n2955 0.0228692
R8557 VSS.n5838 VSS.n5794 0.0227936
R8558 VSS.n5171 VSS.n5161 0.0227632
R8559 VSS.n942 VSS.n938 0.022528
R8560 VSS.n2486 VSS.n2485 0.0225087
R8561 VSS.n1715 VSS.n1714 0.0221201
R8562 VSS.n4398 VSS.n4397 0.0220702
R8563 VSS.n1637 VSS.n1636 0.0220668
R8564 VSS.n5092 VSS.n5091 0.0220044
R8565 VSS.n346 VSS.n343 0.0217195
R8566 VSS.n273 VSS.n272 0.0213929
R8567 VSS.n4401 VSS.n4400 0.0213264
R8568 VSS.n5310 VSS.n5309 0.0213264
R8569 VSS.n5313 VSS.n5312 0.0213264
R8570 VSS.n4374 VSS.n4373 0.0212692
R8571 VSS.n4582 VSS.n4581 0.021208
R8572 VSS.n4507 VSS.n96 0.0209545
R8573 VSS.n5074 VSS.n5071 0.0209545
R8574 VSS.n6101 VSS.n6100 0.0209545
R8575 VSS.n4365 VSS.n4364 0.0208774
R8576 VSS.n2915 VSS.n2914 0.020815
R8577 VSS.n349 VSS.n347 0.0207174
R8578 VSS.n317 VSS.n268 0.0207174
R8579 VSS.n1461 VSS 0.0206399
R8580 VSS.n2141 VSS.n2131 0.0205167
R8581 VSS.n2294 VSS.n2293 0.0205167
R8582 VSS.n4594 VSS.n4590 0.0204115
R8583 VSS.n2574 VSS.n2573 0.0203837
R8584 VSS.n300 VSS.n299 0.0203165
R8585 VSS.n5556 VSS.n5418 0.0203113
R8586 VSS.n5607 VSS.n5606 0.0203113
R8587 VSS.n2543 VSS.n2430 0.0201507
R8588 VSS.n245 VSS.n120 0.0200652
R8589 VSS.n349 VSS.n348 0.0200652
R8590 VSS.n317 VSS.n316 0.0200652
R8591 VSS.n5547 VSS.n5545 0.0200447
R8592 VSS.n5285 VSS.n5284 0.0200283
R8593 VSS.n4166 VSS.n4165 0.0199845
R8594 VSS.n3499 VSS.n3498 0.0198605
R8595 VSS.n4404 VSS.n4403 0.0198388
R8596 VSS.n297 VSS.n276 0.0197857
R8597 VSS.n4503 VSS.n4502 0.0197025
R8598 VSS.n5118 VSS.n5115 0.019615
R8599 VSS.n144 VSS.n143 0.0196091
R8600 VSS.n2591 VSS.n2404 0.0195988
R8601 VSS.n353 VSS.n352 0.0195947
R8602 VSS.n5214 VSS.n5213 0.019555
R8603 VSS.n4794 VSS.n4793 0.019555
R8604 VSS.n2541 VSS.n2431 0.0193646
R8605 VSS.n5166 VSS.n5165 0.0193395
R8606 VSS.n127 VSS.n126 0.0191251
R8607 VSS.n225 VSS.n224 0.0191251
R8608 VSS.n5316 VSS.n5315 0.019095
R8609 VSS.n247 VSS.n245 0.019087
R8610 VSS.n3457 VSS.n3456 0.0190756
R8611 VSS.n4163 VSS.n4162 0.0190567
R8612 VSS.n2721 VSS.n2213 0.0190117
R8613 VSS.n291 VSS.n290 0.0189821
R8614 VSS.n5921 VSS.n4750 0.0189532
R8615 VSS.n3617 VSS.n3616 0.0189448
R8616 VSS.n355 VSS.n354 0.0188673
R8617 VSS.n2589 VSS.n2405 0.018814
R8618 VSS.n5828 VSS.n5803 0.0187609
R8619 VSS.n5217 VSS.n5216 0.0186836
R8620 VSS.n4797 VSS.n4796 0.0186836
R8621 VSS.n5191 VSS.n5190 0.0186836
R8622 VSS.n306 VSS.n305 0.0186651
R8623 VSS.n2539 VSS.n2432 0.0185786
R8624 VSS.n3989 VSS.n3988 0.0185
R8625 VSS.n883 VSS.n882 0.0185
R8626 VSS.n4406 VSS.n4405 0.018485
R8627 VSS.n5315 VSS.n5314 0.0184602
R8628 VSS.n1444 VSS.n1443 0.0184371
R8629 VSS.n3446 VSS.n3445 0.0182907
R8630 VSS.n2732 VSS.n2731 0.0182592
R8631 VSS.n4173 VSS.n4172 0.0181289
R8632 VSS.n4386 VSS.n4385 0.0181087
R8633 VSS.n2719 VSS.n2214 0.0181087
R8634 VSS.n5318 VSS.n5317 0.0181073
R8635 VSS.n4403 VSS.n4402 0.0180867
R8636 VSS.n2587 VSS.n2408 0.0180291
R8637 VSS.n5146 VSS.n5145 0.0180221
R8638 VSS.n4983 VSS.n4982 0.0180221
R8639 VSS.n304 VSS.n303 0.0178394
R8640 VSS.n134 VSS.n131 0.0178182
R8641 VSS.n177 VSS.n174 0.0178182
R8642 VSS.n232 VSS.n229 0.0178182
R8643 VSS.n1425 VSS.n1424 0.0178077
R8644 VSS.n1482 VSS.n1481 0.0178077
R8645 VSS.n797 VSS.n796 0.0178077
R8646 VSS.n863 VSS.n862 0.0178077
R8647 VSS.n2855 VSS.n2021 0.0178077
R8648 VSS.n2292 VSS.n2212 0.0176572
R8649 VSS.n3502 VSS.n3501 0.0176366
R8650 VSS.n1549 VSS.n1548 0.0175923
R8651 VSS.n1539 VSS.n1538 0.0175923
R8652 VSS.n3990 VSS.n3987 0.0175
R8653 VSS.n870 VSS.n856 0.017493
R8654 VSS.n972 VSS.n967 0.0174458
R8655 VSS.n967 VSS.n966 0.0173807
R8656 VSS.n272 VSS.n271 0.017375
R8657 VSS.n275 VSS.n274 0.017375
R8658 VSS.n2570 VSS.n2569 0.017375
R8659 VSS.n2201 VSS.n2194 0.0173562
R8660 VSS.n4609 VSS.n4608 0.0172257
R8661 VSS.n2717 VSS.n2215 0.0172057
R8662 VSS.n971 VSS.n968 0.0171955
R8663 VSS.n253 VSS.n252 0.0171304
R8664 VSS.n264 VSS.n263 0.0170306
R8665 VSS.n3071 VSS.n3070 0.0167984
R8666 VSS.n2855 VSS.n2854 0.0167542
R8667 VSS.n1407 VSS.n1406 0.0165
R8668 VSS.n2021 VSS.n1995 0.0164532
R8669 VSS.n2207 VSS.n2206 0.0164532
R8670 VSS.n4571 VSS.n4570 0.0164292
R8671 VSS.n4170 VSS.n4169 0.0162732
R8672 VSS.n948 VSS.n947 0.0162343
R8673 VSS.n4863 VSS.n4860 0.0162343
R8674 VSS.n4825 VSS.n4822 0.0162343
R8675 VSS.n4897 VSS.n4894 0.0162343
R8676 VSS.n4938 VSS.n4935 0.0162343
R8677 VSS.n4140 VSS.n4138 0.0162343
R8678 VSS.n2545 VSS.n2428 0.0162205
R8679 VSS.n5228 VSS.n5225 0.0161522
R8680 VSS.n318 VSS.n267 0.0161122
R8681 VSS.n3402 VSS.n3401 0.0160669
R8682 VSS.n736 VSS.n713 0.0158659
R8683 VSS.n5312 VSS.n5311 0.015852
R8684 VSS.n877 VSS.n876 0.0158
R8685 VSS.n1469 VSS 0.0156049
R8686 VSS.n1853 VSS.n1852 0.0155517
R8687 VSS.n1512 VSS.n1407 0.0155
R8688 VSS.n2547 VSS.n2424 0.0154345
R8689 VSS.n2184 VSS.n2129 0.0153997
R8690 VSS.n5287 VSS.n5286 0.015398
R8691 VSS.n2302 VSS.n2301 0.0152492
R8692 VSS.n215 VSS.n214 0.0151739
R8693 VSS.n4400 VSS.n4399 0.0151082
R8694 VSS.n5309 VSS.n5308 0.0151082
R8695 VSS.n2828 VSS.n2068 0.0150987
R8696 VSS.n5902 VSS.n5899 0.0150588
R8697 VSS.n3586 VSS.n3585 0.0150203
R8698 VSS.n3393 VSS.n3392 0.0148895
R8699 VSS.n5085 VSS.n5083 0.0148363
R8700 VSS.n5292 VSS.n5282 0.0148234
R8701 VSS.n4371 VSS.n4360 0.0148073
R8702 VSS.n5650 VSS.n5649 0.0147683
R8703 VSS.n4397 VSS.n4396 0.0147345
R8704 VSS.n840 VSS.n789 0.0146608
R8705 VSS.n2550 VSS.n2549 0.0146485
R8706 VSS.n3611 VSS.n3610 0.0146279
R8707 VSS.n1893 VSS.n1892 0.0146207
R8708 VSS.n4367 VSS.n4366 0.014549
R8709 VSS.n2746 VSS.n2745 0.0144967
R8710 VSS.n1872 VSS.n1871 0.0144655
R8711 VSS.n358 VSS.n357 0.0144024
R8712 VSS.n2678 VSS.n2677 0.0143462
R8713 VSS.n2830 VSS.n2065 0.0141957
R8714 VSS.n5864 VSS.n5863 0.0141817
R8715 VSS.n296 VSS 0.0141607
R8716 VSS.n319 VSS.n262 0.0141607
R8717 VSS.n1505 VSS.n1504 0.0141607
R8718 VSS.n5794 VSS.n5792 0.0141239
R8719 VSS.n3525 VSS.n3524 0.0141047
R8720 VSS.n2878 VSS.n1996 0.0140452
R8721 VSS.n4987 VSS.n4986 0.0140398
R8722 VSS.n57 VSS.n56 0.0140398
R8723 VSS.n1660 VSS.n1659 0.0140123
R8724 VSS.n1690 VSS.n1689 0.0140123
R8725 VSS.n1668 VSS.n1667 0.0140123
R8726 VSS.n1453 VSS.n1452 0.0139579
R8727 VSS.n4692 VSS.n4691 0.0138333
R8728 VSS.n2518 VSS.n2453 0.0137314
R8729 VSS.n1930 VSS.n1929 0.0136897
R8730 VSS.n5636 VSS.n5633 0.0136707
R8731 VSS.n2166 VSS.n2163 0.0135936
R8732 VSS.n1877 VSS.n1876 0.0135345
R8733 VSS.n4696 VSS.n4692 0.0135
R8734 VSS.n4169 VSS.n4168 0.0134897
R8735 VSS.n2271 VSS.n2268 0.0134431
R8736 VSS.n3487 VSS.n3486 0.0133198
R8737 VSS.n2833 VSS.n2832 0.0132926
R8738 VSS.n1815 VSS.n1814 0.0132273
R8739 VSS.n2944 VSS.n2943 0.013189
R8740 VSS.n2876 VSS.n1997 0.0131421
R8741 VSS.n4161 VSS.n4160 0.0130874
R8742 VSS.n2516 VSS.n2454 0.0129454
R8743 VSS.n1977 VSS.n1976 0.0126034
R8744 VSS.n3850 VSS.n3849 0.0125737
R8745 VSS.n774 VSS.n751 0.0125732
R8746 VSS.n3559 VSS.n3558 0.0125349
R8747 VSS.n3990 VSS.n3989 0.0125
R8748 VSS.n4175 VSS.n4174 0.012458
R8749 VSS.n267 VSS.n266 0.0124388
R8750 VSS.n90 VSS.n85 0.0124337
R8751 VSS.n5112 VSS.n5111 0.0124337
R8752 VSS.n4506 VSS.n4505 0.0123681
R8753 VSS.n72 VSS.n69 0.0123033
R8754 VSS.n5133 VSS.n5132 0.0123033
R8755 VSS.n1454 VSS.n1453 0.0122757
R8756 VSS.n2874 VSS.n1998 0.0122391
R8757 VSS.n876 VSS.n875 0.0122
R8758 VSS.n2514 VSS.n2456 0.0121594
R8759 VSS.n88 VSS.n87 0.0119894
R8760 VSS.n4586 VSS.n93 0.0119365
R8761 VSS.n5108 VSS.n5106 0.0119365
R8762 VSS.n5073 VSS.n5072 0.0118736
R8763 VSS.n4027 VSS.n4026 0.0118287
R8764 VSS.n4598 VSS.n75 0.0118115
R8765 VSS.n5129 VSS.n5126 0.0118115
R8766 VSS.n5826 VSS.n5825 0.0118043
R8767 VSS.n2788 VSS.n2095 0.0117876
R8768 VSS.n360 VSS.n337 0.01175
R8769 VSS.n2605 VSS.n2389 0.0116192
R8770 VSS.n352 VSS.n351 0.0115204
R8771 VSS.n71 VSS.n70 0.0113172
R8772 VSS.n5128 VSS.n5127 0.0113172
R8773 VSS.n3996 VSS.n3995 0.0111993
R8774 VSS.n2809 VSS.n2086 0.0111355
R8775 VSS.n964 VSS.n961 0.0109464
R8776 VSS.n289 VSS.n286 0.0109464
R8777 VSS.n320 VSS.n319 0.0109464
R8778 VSS.n4218 VSS.n4215 0.0109464
R8779 VSS.n2786 VSS.n2096 0.0108846
R8780 VSS.n2607 VSS.n2386 0.0108343
R8781 VSS.n5838 VSS.n5837 0.0107901
R8782 VSS.n4172 VSS.n4171 0.0107062
R8783 VSS.n1653 VSS.n1652 0.0106256
R8784 VSS.n2655 VSS.n2321 0.0105727
R8785 VSS.n1472 VSS.n1469 0.0105699
R8786 VSS.n3993 VSS.n1523 0.0105699
R8787 VSS.n4187 VSS.n4186 0.0105699
R8788 VSS.n5823 VSS.n5822 0.0105
R8789 VSS.n2139 VSS.n2138 0.0104331
R8790 VSS.n2700 VSS.n2237 0.0104331
R8791 VSS.n1684 VSS.n1683 0.0102906
R8792 VSS.n973 VSS.n972 0.0101429
R8793 VSS.n1506 VSS.n1505 0.0101429
R8794 VSS.n333 VSS.n330 0.0101429
R8795 VSS.n4090 VSS.n4089 0.0101429
R8796 VSS.n4127 VSS.n4126 0.0101429
R8797 VSS.n3867 VSS.n3866 0.0100852
R8798 VSS.n3588 VSS.n3587 0.0100494
R8799 VSS.n2610 VSS.n2609 0.0100494
R8800 VSS.n343 VSS.n322 0.0100122
R8801 VSS.n2784 VSS.n2097 0.00998161
R8802 VSS.n5133 VSS.n5120 0.00997368
R8803 VSS.n1522 VSS.n1521 0.00994056
R8804 VSS.n1514 VSS.n1513 0.00994056
R8805 VSS.n3885 VSS.n3884 0.00989535
R8806 VSS.n3809 VSS.n3808 0.00982401
R8807 VSS.n2653 VSS.n2322 0.00978779
R8808 VSS.n4164 VSS.n4163 0.00977835
R8809 VSS.n4173 VSS.n4166 0.00977835
R8810 VSS.n2964 VSS.n2963 0.00974419
R8811 VSS.n356 VSS.n355 0.00968367
R8812 VSS.n2131 VSS.n2130 0.0096806
R8813 VSS.n1577 VSS 0.00958911
R8814 VSS.n881 VSS.n880 0.00958707
R8815 VSS.n2766 VSS.n2765 0.0095301
R8816 VSS.n2698 VSS.n2238 0.0095301
R8817 VSS.n2332 VSS.n2320 0.00952616
R8818 VSS.n4598 VSS.n4597 0.0095
R8819 VSS.n3585 VSS.n3584 0.00939535
R8820 VSS.n4186 VSS.n4185 0.00931119
R8821 VSS.n4195 VSS.n4194 0.00931119
R8822 VSS.n3384 VSS.n3383 0.00926454
R8823 VSS.n68 VSS.n67 0.00925
R8824 VSS.n5125 VSS.n5124 0.00925
R8825 VSS.n4589 VSS.n4586 0.00902632
R8826 VSS.n2651 VSS.n2323 0.00900291
R8827 VSS.n5590 VSS.n5587 0.00899057
R8828 VSS.n3516 VSS.n3515 0.00887209
R8829 VSS.n4733 VSS.n4732 0.00883333
R8830 VSS.n1405 VSS.n1404 0.00868182
R8831 VSS.n870 VSS.n869 0.00868182
R8832 VSS.n4160 VSS.n4159 0.00868182
R8833 VSS.n4180 VSS.n4175 0.00868182
R8834 VSS.n2130 VSS.n2094 0.00862709
R8835 VSS.n2119 VSS.n2116 0.00862709
R8836 VSS.n2295 VSS.n2294 0.00862709
R8837 VSS.n2696 VSS.n2241 0.00862709
R8838 VSS.n3858 VSS.n3857 0.0086106
R8839 VSS.n2630 VSS.n2629 0.00861047
R8840 VSS.n5114 VSS.n5112 0.00855263
R8841 VSS.n2886 VSS.n2885 0.00855063
R8842 VSS.n3284 VSS.n3283 0.00847965
R8843 VSS.n3569 VSS.n3568 0.00840698
R8844 VSS.n2538 VSS.n2537 0.00838571
R8845 VSS.n1553 VSS.n1552 0.00836872
R8846 VSS.n1725 VSS.n1724 0.00836872
R8847 VSS.n1543 VSS.n1542 0.00836872
R8848 VSS.n1428 VSS.n1425 0.00836713
R8849 VSS.n1485 VSS.n1482 0.00836713
R8850 VSS.n800 VSS.n797 0.00836713
R8851 VSS.n866 VSS.n863 0.00836713
R8852 VSS.n2569 VSS.n2332 0.00834884
R8853 VSS.n3773 VSS.n3772 0.00833217
R8854 VSS.n198 VSS.n195 0.00832609
R8855 VSS.n2586 VSS.n2585 0.0082907
R8856 VSS.n3473 VSS.n3472 0.00808721
R8857 VSS.n3228 VSS.n3227 0.00808721
R8858 VSS.n4004 VSS.n4003 0.00805245
R8859 VSS.n3995 VSS.n3994 0.00805245
R8860 VSS.n3905 VSS.n3904 0.0080419
R8861 VSS.n1673 VSS.n1650 0.0080419
R8862 VSS.n2796 VSS.n2022 0.00802508
R8863 VSS.n1288 VSS.n1284 0.008
R8864 VSS.n3625 VSS.n3624 0.00797826
R8865 VSS.n1168 VSS.n1165 0.00795562
R8866 VSS.n1866 VSS.n1865 0.00794828
R8867 VSS.n305 VSS.n304 0.00793119
R8868 VSS.n303 VSS.n302 0.00793119
R8869 VSS.n265 VSS.n264 0.00784694
R8870 VSS.n2349 VSS.n2347 0.00782558
R8871 VSS.n357 VSS.n346 0.00781707
R8872 VSS.n1663 VSS.n1662 0.0077905
R8873 VSS.n1709 VSS.n1708 0.0077905
R8874 VSS.n3897 VSS.n1718 0.0077905
R8875 VSS.n1649 VSS.n1648 0.0077905
R8876 VSS.n274 VSS.n273 0.00773214
R8877 VSS.n2857 VSS.n2015 0.00772408
R8878 VSS.n3290 VSS.n3289 0.00769477
R8879 VSS.n5551 VSS.n5548 0.00760526
R8880 VSS.n2232 VSS.n2231 0.00757358
R8881 VSS.n1508 VSS.n1507 0.00757142
R8882 VSS.n1662 VSS.n1657 0.00753911
R8883 VSS.n1669 VSS.n1664 0.00753911
R8884 VSS.n1697 VSS.n1696 0.00753911
R8885 VSS.n2716 VSS.n2715 0.00748113
R8886 VSS.n1504 VSS.n1503 0.00743371
R8887 VSS VSS.n4008 0.00742308
R8888 VSS.n4003 VSS.n3996 0.00742308
R8889 VSS.n882 VSS.n881 0.00735714
R8890 VSS.n5245 VSS.n5244 0.00734783
R8891 VSS.n1611 VSS.n1610 0.00734332
R8892 VSS.n1641 VSS.n1640 0.00734332
R8893 VSS.n2208 VSS.n2198 0.0073277
R8894 VSS.n3545 VSS.n3544 0.00730233
R8895 VSS.n1671 VSS.n1670 0.00728771
R8896 VSS.n1713 VSS.n1712 0.00728771
R8897 VSS.n1813 VSS.n1812 0.00726364
R8898 VSS.n1609 VSS.n1608 0.00713594
R8899 VSS.n1639 VSS.n1638 0.00713594
R8900 VSS.n767 VSS.n766 0.00708537
R8901 VSS.n4330 VSS.n4328 0.00708537
R8902 VSS.n2356 VSS.n2354 0.0070407
R8903 VSS.n3907 VSS.n1691 0.00703631
R8904 VSS.n1701 VSS.n1700 0.00703631
R8905 VSS.n1705 VSS.n1704 0.00703631
R8906 VSS.n3803 VSS.n3794 0.00701869
R8907 VSS.n1961 VSS.n1960 0.00701724
R8908 VSS.n5130 VSS.n5129 0.00689344
R8909 VSS.n1032 VSS.n1024 0.00686364
R8910 VSS.n1862 VSS.n1861 0.00686207
R8911 VSS.n2859 VSS.n2012 0.00682107
R8912 VSS.n4501 VSS.n4486 0.00681579
R8913 VSS.n3788 VSS.n3778 0.00680841
R8914 VSS.n4161 VSS.n4146 0.00679371
R8915 VSS.n4159 VSS.n4147 0.00679371
R8916 VSS.n4174 VSS.n788 0.00679371
R8917 VSS.n4181 VSS.n4180 0.00679371
R8918 VSS.n1686 VSS.n1680 0.00678492
R8919 VSS.n1693 VSS.n1692 0.00678492
R8920 VSS.n2929 VSS.n2928 0.00677907
R8921 VSS.n3358 VSS.n3357 0.00668497
R8922 VSS.n2551 VSS.n2421 0.00667143
R8923 VSS.n2038 VSS.n2016 0.00667057
R8924 VSS.n2711 VSS.n2710 0.00667057
R8925 VSS.n1869 VSS.n1868 0.00655172
R8926 VSS.n1333 VSS.n1332 0.00655042
R8927 VSS.n5938 VSS.n5936 0.00653659
R8928 VSS VSS.n5766 0.00652231
R8929 VSS.n1557 VSS.n1556 0.00651383
R8930 VSS.n1584 VSS.n1583 0.00651383
R8931 VSS.n1509 VSS.n1508 0.0065
R8932 VSS.n736 VSS.n735 0.0064434
R8933 VSS.n701 VSS.n511 0.0064434
R8934 VSS.n774 VSS.n773 0.0064434
R8935 VSS.n4313 VSS.n4312 0.0064434
R8936 VSS.n73 VSS.n72 0.00640164
R8937 VSS.n2019 VSS.n2018 0.00636957
R8938 VSS.n1644 VSS.n1582 0.00630645
R8939 VSS.n1642 VSS.n1607 0.00630645
R8940 VSS.n301 VSS.n300 0.00627982
R8941 VSS.n3602 VSS.n3601 0.00625581
R8942 VSS.n2573 VSS.n2571 0.00625581
R8943 VSS.n1979 VSS.n1978 0.00624138
R8944 VSS.n1974 VSS.n1968 0.00624138
R8945 VSS.n1964 VSS.n1958 0.00624138
R8946 VSS.n1954 VSS.n1953 0.00624138
R8947 VSS.n1932 VSS.n1931 0.00624138
R8948 VSS.n1911 VSS.n1906 0.00624138
R8949 VSS.n1402 VSS.n912 0.00622751
R8950 VSS.n2834 VSS.n2062 0.00618562
R8951 VSS.n1565 VSS.n1564 0.00617757
R8952 VSS.n3797 VSS.n3796 0.00617757
R8953 VSS.n3820 VSS.n3819 0.00617757
R8954 VSS.n3802 VSS.n3801 0.00617757
R8955 VSS.n3767 VSS.n3757 0.00617757
R8956 VSS.n3319 VSS.n3318 0.00616474
R8957 VSS.n4194 VSS.n4187 0.00616434
R8958 VSS.n960 VSS 0.006125
R8959 VSS.n291 VSS 0.006125
R8960 VSS.n4207 VSS 0.006125
R8961 VSS.n2168 VSS.n2162 0.00610386
R8962 VSS.n1975 VSS.n1974 0.00608621
R8963 VSS.n1965 VSS.n1964 0.00608621
R8964 VSS.n1957 VSS.n1956 0.00608621
R8965 VSS.n1955 VSS.n1954 0.00608621
R8966 VSS.n1912 VSS.n1911 0.00608621
R8967 VSS.n2875 VSS.n1993 0.00606856
R8968 VSS.n2870 VSS.n2869 0.00606856
R8969 VSS.n2865 VSS.n2008 0.00606856
R8970 VSS.n2035 VSS.n2011 0.00606856
R8971 VSS.n2063 VSS.n2050 0.00606856
R8972 VSS.n2794 VSS.n2087 0.00606856
R8973 VSS.n2785 VSS.n2092 0.00606856
R8974 VSS.n2768 VSS.n2767 0.00606856
R8975 VSS.n2728 VSS.n2197 0.00606856
R8976 VSS.n2718 VSS.n2210 0.00606856
R8977 VSS.n2713 VSS.n2712 0.00606856
R8978 VSS.n2661 VSS.n2310 0.00606856
R8979 VSS.n3651 VSS.n3650 0.00606522
R8980 VSS.n3506 VSS.n3505 0.00599419
R8981 VSS.n1822 VSS.n1821 0.00599419
R8982 VSS.n5109 VSS.n5108 0.00596961
R8983 VSS.n3785 VSS.n3784 0.00596729
R8984 VSS.n3786 VSS.n3782 0.00596729
R8985 VSS.n3751 VSS.n3743 0.00596729
R8986 VSS.n1884 VSS.n1883 0.00593103
R8987 VSS.n2881 VSS.n1993 0.00591806
R8988 VSS.n2870 VSS.n2000 0.00591806
R8989 VSS.n2866 VSS.n2865 0.00591806
R8990 VSS.n2862 VSS.n2861 0.00591806
R8991 VSS.n2860 VSS.n2011 0.00591806
R8992 VSS.n2806 VSS.n2087 0.00591806
R8993 VSS.n2791 VSS.n2092 0.00591806
R8994 VSS.n2780 VSS.n2099 0.00591806
R8995 VSS.n2728 VSS.n2196 0.00591806
R8996 VSS.n2724 VSS.n2210 0.00591806
R8997 VSS.n2713 VSS.n2217 0.00591806
R8998 VSS.n2692 VSS.n2244 0.00591806
R8999 VSS.n2273 VSS.n2267 0.0059088
R9000 VSS.n1621 VSS.n1620 0.0058917
R9001 VSS.n1633 VSS.n1632 0.0058917
R9002 VSS.n1675 VSS.n1674 0.00588013
R9003 VSS.n2933 VSS.n2932 0.00586337
R9004 VSS.n825 VSS.n789 0.00584965
R9005 VSS.n3434 VSS.n3433 0.00584884
R9006 VSS.n1873 VSS.n1872 0.00577586
R9007 VSS.n1870 VSS.n1869 0.00577586
R9008 VSS.n1867 VSS.n1866 0.00577586
R9009 VSS.n1864 VSS.n1862 0.00577586
R9010 VSS.n1854 VSS.n1853 0.00577586
R9011 VSS.n1879 VSS.n1878 0.00577586
R9012 VSS.n1973 VSS.n1972 0.00577586
R9013 VSS.n1963 VSS.n1962 0.00577586
R9014 VSS.n1886 VSS.n1885 0.00577586
R9015 VSS.n1895 VSS.n1894 0.00577586
R9016 VSS.n2040 VSS.n2036 0.00576756
R9017 VSS.n2223 VSS.n2220 0.00576756
R9018 VSS.n2873 VSS.n2872 0.00571739
R9019 VSS.n1617 VSS.n1616 0.00568433
R9020 VSS.n1629 VSS.n1628 0.00568433
R9021 VSS.n1871 VSS.n1870 0.00562069
R9022 VSS.n1868 VSS.n1867 0.00562069
R9023 VSS.n1865 VSS.n1864 0.00562069
R9024 VSS.n1908 VSS.n1907 0.00562069
R9025 VSS.n1971 VSS.n1970 0.00562069
R9026 VSS.n2879 VSS.n2878 0.00561706
R9027 VSS.n2018 VSS.n2017 0.00561706
R9028 VSS.n2020 VSS.n2015 0.00561706
R9029 VSS.n2856 VSS.n2016 0.00561706
R9030 VSS.n2068 VSS.n2047 0.00561706
R9031 VSS.n2877 VSS.n1994 0.00561706
R9032 VSS.n2004 VSS.n2002 0.00561706
R9033 VSS.n2014 VSS.n2007 0.00561706
R9034 VSS.n2031 VSS.n2013 0.00561706
R9035 VSS.n2067 VSS.n2048 0.00561706
R9036 VSS.n2143 VSS.n2142 0.00561706
R9037 VSS.n2789 VSS.n2788 0.00561706
R9038 VSS.n2138 VSS.n2137 0.00561706
R9039 VSS.n2753 VSS.n2129 0.00561706
R9040 VSS.n2787 VSS.n2093 0.00561706
R9041 VSS.n2117 VSS.n2115 0.00561706
R9042 VSS.n2722 VSS.n2721 0.00561706
R9043 VSS.n2231 VSS.n2230 0.00561706
R9044 VSS.n2720 VSS.n2211 0.00561706
R9045 VSS.n2221 VSS.n2219 0.00561706
R9046 VSS.n2925 VSS.n2924 0.00560174
R9047 VSS.n3828 VSS.n3827 0.00554673
R9048 VSS.n1455 VSS.n1444 0.00553496
R9049 VSS.n1462 VSS.n1461 0.00553496
R9050 VSS.n1521 VSS.n1514 0.00553496
R9051 VSS.n3894 VSS.n3893 0.00552326
R9052 VSS.n4691 VSS.n4690 0.0055
R9053 VSS.n91 VSS.n90 0.00547238
R9054 VSS.n3691 VSS.n3690 0.00547093
R9055 VSS.n2017 VSS.n1996 0.00546656
R9056 VSS.n2020 VSS.n2019 0.00546656
R9057 VSS.n2857 VSS.n2856 0.00546656
R9058 VSS.n2803 VSS.n2802 0.00546656
R9059 VSS.n2002 VSS.n2001 0.00546656
R9060 VSS.n2868 VSS.n2867 0.00546656
R9061 VSS.n2007 VSS.n2005 0.00546656
R9062 VSS.n2858 VSS.n2013 0.00546656
R9063 VSS.n2804 VSS.n2089 0.00546656
R9064 VSS.n2142 VSS.n2141 0.00546656
R9065 VSS.n2102 VSS.n2095 0.00546656
R9066 VSS.n2140 VSS.n2139 0.00546656
R9067 VSS.n2140 VSS.n2127 0.00546656
R9068 VSS.n2754 VSS.n2753 0.00546656
R9069 VSS.n2731 VSS.n2193 0.00546656
R9070 VSS.n2779 VSS.n2101 0.00546656
R9071 VSS.n2730 VSS.n2729 0.00546656
R9072 VSS.n2230 VSS.n2213 0.00546656
R9073 VSS.n2247 VSS.n2237 0.00546656
R9074 VSS.n2219 VSS.n2218 0.00546656
R9075 VSS.n2691 VSS.n2246 0.00546656
R9076 VSS.n1808 VSS.n1807 0.00546429
R9077 VSS.n2512 VSS.n2511 0.00541429
R9078 VSS.n4418 VSS.n4414 0.0053913
R9079 VSS.n3004 VSS.n3003 0.00538372
R9080 VSS.n2422 VSS.n2418 0.00534716
R9081 VSS.n2540 VSS.n2423 0.00534716
R9082 VSS.n3622 VSS.n3621 0.00534012
R9083 VSS.n3503 VSS.n3502 0.00534012
R9084 VSS.n3561 VSS.n3560 0.00534012
R9085 VSS.n3542 VSS.n3541 0.00534012
R9086 VSS.n1770 VSS.n1766 0.00534012
R9087 VSS.n3274 VSS.n3267 0.00534012
R9088 VSS.n3239 VSS.n3205 0.00534012
R9089 VSS.n3197 VSS.n3193 0.00534012
R9090 VSS.n3170 VSS.n3169 0.00534012
R9091 VSS.n3130 VSS.n3123 0.00534012
R9092 VSS.n3089 VSS.n3088 0.00534012
R9093 VSS.n3068 VSS.n3067 0.00534012
R9094 VSS.n1825 VSS.n1819 0.00534012
R9095 VSS.n3048 VSS.n3047 0.00534012
R9096 VSS.n3014 VSS.n3013 0.00534012
R9097 VSS.n2961 VSS.n2960 0.00534012
R9098 VSS.n2652 VSS.n2318 0.00534012
R9099 VSS.n2633 VSS.n2341 0.00534012
R9100 VSS.n2384 VSS.n2366 0.00534012
R9101 VSS.n2583 VSS.n2582 0.00534012
R9102 VSS.n3761 VSS.n3760 0.00533645
R9103 VSS.n3766 VSS.n3765 0.00533645
R9104 VSS.n3833 VSS.n3832 0.00533645
R9105 VSS.n3813 VSS.n3812 0.00533645
R9106 VSS.n297 VSS.n296 0.00532143
R9107 VSS.n359 VSS 0.00532143
R9108 VSS VSS.n4091 0.00532143
R9109 VSS VSS.n4129 0.00532143
R9110 VSS.n1810 VSS.n1809 0.00527273
R9111 VSS.n2562 VSS.n2411 0.00521616
R9112 VSS.n2548 VSS.n2423 0.00521616
R9113 VSS.n3684 VSS.n3670 0.0052093
R9114 VSS.n3622 VSS.n3576 0.0052093
R9115 VSS.n3439 VSS.n3438 0.0052093
R9116 VSS.n3444 VSS.n3443 0.0052093
R9117 VSS.n3566 VSS.n3447 0.0052093
R9118 VSS.n3543 VSS.n3542 0.0052093
R9119 VSS.n3413 VSS.n3362 0.0052093
R9120 VSS.n3413 VSS.n3366 0.0052093
R9121 VSS.n3274 VSS.n3263 0.0052093
R9122 VSS.n3239 VSS.n3201 0.0052093
R9123 VSS.n3115 VSS.n3114 0.0052093
R9124 VSS.n3068 VSS.n3056 0.0052093
R9125 VSS.n1818 VSS.n1817 0.0052093
R9126 VSS.n2961 VSS.n2918 0.0052093
R9127 VSS.n2658 VSS.n2318 0.0052093
R9128 VSS.n2325 VSS.n2324 0.0052093
R9129 VSS.n2583 VSS.n2565 0.0052093
R9130 VSS.n2757 VSS.n2125 0.00516555
R9131 VSS.n2164 VSS.n2144 0.00516555
R9132 VSS.n2748 VSS.n2747 0.00516555
R9133 VSS.n3748 VSS.n3747 0.00512617
R9134 VSS.n3749 VSS.n3746 0.00512617
R9135 VSS.n3817 VSS.n3816 0.00512617
R9136 VSS.n5293 VSS.n5292 0.00511538
R9137 VSS.n4372 VSS.n4371 0.00511538
R9138 VSS.n318 VSS.n265 0.00509184
R9139 VSS.n3593 VSS.n3592 0.00507849
R9140 VSS.n1572 VSS.n1571 0.00506221
R9141 VSS.n1592 VSS.n1591 0.00506221
R9142 VSS.n1602 VSS.n1601 0.00506221
R9143 VSS.n5936 VSS.n5935 0.00504545
R9144 VSS.n2124 VSS.n2118 0.00501505
R9145 VSS.n2752 VSS.n2128 0.00501505
R9146 VSS.n2764 VSS.n2763 0.00501505
R9147 VSS.n1952 VSS.n1951 0.005
R9148 VSS.n2428 VSS.n2426 0.00495415
R9149 VSS.n2544 VSS.n2543 0.00495415
R9150 VSS.n2427 VSS.n2416 0.00495415
R9151 VSS.n2542 VSS.n2425 0.00495415
R9152 VSS.n3595 VSS.n3594 0.00494767
R9153 VSS.n3604 VSS.n3603 0.00494767
R9154 VSS.n3717 VSS.n3716 0.00494767
R9155 VSS.n3721 VSS.n3720 0.00494767
R9156 VSS.n3498 VSS.n3497 0.00494767
R9157 VSS.n3526 VSS.n3525 0.00494767
R9158 VSS.n3517 VSS.n3516 0.00494767
R9159 VSS.n3514 VSS.n3513 0.00494767
R9160 VSS.n3455 VSS.n3454 0.00494767
R9161 VSS.n3489 VSS.n3488 0.00494767
R9162 VSS.n3475 VSS.n3474 0.00494767
R9163 VSS.n3470 VSS.n3469 0.00494767
R9164 VSS.n3441 VSS.n3440 0.00494767
R9165 VSS.n3547 VSS.n3546 0.00494767
R9166 VSS.n3406 VSS.n3405 0.00494767
R9167 VSS.n3403 VSS.n3402 0.00494767
R9168 VSS.n3382 VSS.n3381 0.00494767
R9169 VSS.n3412 VSS.n3411 0.00494767
R9170 VSS.n1769 VSS.n1768 0.00494767
R9171 VSS.n3273 VSS.n3272 0.00494767
R9172 VSS.n3232 VSS.n3231 0.00494767
R9173 VSS.n3229 VSS.n3228 0.00494767
R9174 VSS.n3219 VSS.n3218 0.00494767
R9175 VSS.n3075 VSS.n3074 0.00494767
R9176 VSS.n3079 VSS.n3078 0.00494767
R9177 VSS.n3238 VSS.n3237 0.00494767
R9178 VSS.n3196 VSS.n3195 0.00494767
R9179 VSS.n3165 VSS.n3164 0.00494767
R9180 VSS.n3129 VSS.n3128 0.00494767
R9181 VSS.n3110 VSS.n3109 0.00494767
R9182 VSS.n2924 VSS.n2923 0.00494767
R9183 VSS.n2928 VSS.n2927 0.00494767
R9184 VSS.n2932 VSS.n2931 0.00494767
R9185 VSS.n2943 VSS.n2942 0.00494767
R9186 VSS.n3063 VSS.n3062 0.00494767
R9187 VSS.n1824 VSS.n1823 0.00494767
R9188 VSS.n3044 VSS.n3043 0.00494767
R9189 VSS.n3011 VSS.n3010 0.00494767
R9190 VSS.n2656 VSS.n2655 0.00494767
R9191 VSS.n2642 VSS.n2331 0.00494767
R9192 VSS.n2630 VSS.n2346 0.00494767
R9193 VSS.n2572 VSS.n2389 0.00494767
R9194 VSS.n2654 VSS.n2319 0.00494767
R9195 VSS.n2632 VSS.n2631 0.00494767
R9196 VSS.n2388 VSS.n2364 0.00494767
R9197 VSS VSS.n922 0.00490559
R9198 VSS.n1431 VSS.n1428 0.00490559
R9199 VSS.n1437 VSS.n1434 0.00490559
R9200 VSS.n1443 VSS.n1440 0.00490559
R9201 VSS.n1475 VSS.n1472 0.00490559
R9202 VSS.n1500 VSS.n1497 0.00490559
R9203 VSS.n1494 VSS.n1491 0.00490559
R9204 VSS.n1488 VSS.n1485 0.00490559
R9205 VSS.n4013 VSS 0.00490559
R9206 VSS.n803 VSS.n800 0.00490559
R9207 VSS.n809 VSS.n806 0.00490559
R9208 VSS.n815 VSS.n812 0.00490559
R9209 VSS.n819 VSS.n818 0.00490559
R9210 VSS.n843 VSS.n840 0.00490559
R9211 VSS.n856 VSS.n853 0.00490559
R9212 VSS.n869 VSS.n866 0.00490559
R9213 VSS VSS.n4853 0.00490559
R9214 VSS VSS.n4816 0.00490559
R9215 VSS VSS.n4810 0.00490559
R9216 VSS VSS.n4928 0.00490559
R9217 VSS VSS.n4153 0.00490559
R9218 VSS.n322 VSS.n321 0.00489024
R9219 VSS.n2034 VSS.n2030 0.00486455
R9220 VSS.n1512 VSS.n1511 0.00486421
R9221 VSS.n1569 VSS.n1559 0.00485484
R9222 VSS.n1576 VSS.n1575 0.00485484
R9223 VSS.n1590 VSS.n1589 0.00485484
R9224 VSS.n1600 VSS.n1599 0.00485484
R9225 VSS.n2545 VSS.n2544 0.00482314
R9226 VSS.n2546 VSS.n2425 0.00482314
R9227 VSS.n3594 VSS.n3593 0.00481686
R9228 VSS.n3603 VSS.n3602 0.00481686
R9229 VSS.n3618 VSS.n3617 0.00481686
R9230 VSS.n3620 VSS.n3578 0.00481686
R9231 VSS.n3636 VSS.n3635 0.00481686
R9232 VSS.n3529 VSS.n3499 0.00481686
R9233 VSS.n3515 VSS.n3514 0.00481686
R9234 VSS.n3530 VSS.n3458 0.00481686
R9235 VSS.n3471 VSS.n3470 0.00481686
R9236 VSS.n3404 VSS.n3403 0.00481686
R9237 VSS.n3383 VSS.n3382 0.00481686
R9238 VSS.n3380 VSS.n3379 0.00481686
R9239 VSS.n3273 VSS.n3268 0.00481686
R9240 VSS.n3230 VSS.n3229 0.00481686
R9241 VSS.n3218 VSS.n3217 0.00481686
R9242 VSS.n3217 VSS.n3216 0.00481686
R9243 VSS.n3078 VSS.n3076 0.00481686
R9244 VSS.n3082 VSS.n3080 0.00481686
R9245 VSS.n2923 VSS.n2921 0.00481686
R9246 VSS.n2927 VSS.n2925 0.00481686
R9247 VSS.n2931 VSS.n2929 0.00481686
R9248 VSS.n2957 VSS.n2956 0.00481686
R9249 VSS.n3063 VSS.n3058 0.00481686
R9250 VSS.n3061 VSS.n3060 0.00481686
R9251 VSS.n2959 VSS.n2920 0.00481686
R9252 VSS.n2331 VSS.n2321 0.00481686
R9253 VSS.n2641 VSS.n2640 0.00481686
R9254 VSS.n2580 VSS.n2404 0.00481686
R9255 VSS.n2329 VSS.n2328 0.00481686
R9256 VSS.n2644 VSS.n2329 0.00481686
R9257 VSS.n2567 VSS.n2566 0.00481686
R9258 VSS.n2895 VSS.n2894 0.0048038
R9259 VSS.n3844 VSS.n3842 0.00476036
R9260 VSS.n3872 VSS.n3871 0.00476036
R9261 VSS.n3875 VSS.n3874 0.00476036
R9262 VSS.n2611 VSS.n2383 0.00474419
R9263 VSS.n2132 VSS.n2108 0.00471405
R9264 VSS.n2760 VSS.n2759 0.00471405
R9265 VSS.n1967 VSS.n1966 0.00468966
R9266 VSS.n3683 VSS.n3682 0.00468605
R9267 VSS.n3697 VSS.n3696 0.00468605
R9268 VSS.n3647 VSS.n3641 0.00468605
R9269 VSS.n3378 VSS.n3377 0.00468605
R9270 VSS.n3249 VSS.n3248 0.00468605
R9271 VSS.n3245 VSS.n3244 0.00468605
R9272 VSS.n3215 VSS.n3214 0.00468605
R9273 VSS.n2639 VSS.n2334 0.00468605
R9274 VSS.n2006 VSS.n2003 0.00456355
R9275 VSS.n2137 VSS.n2136 0.00456355
R9276 VSS.n2751 VSS.n2146 0.00456355
R9277 VSS.n1454 VSS.n1450 0.00456316
R9278 VSS.n2783 VSS.n2782 0.00455797
R9279 VSS.n3564 VSS.n3563 0.00455523
R9280 VSS.n2914 VSS.n2913 0.00444937
R9281 VSS.n2555 VSS.n2417 0.00443013
R9282 VSS.n3615 VSS.n3614 0.00442442
R9283 VSS.n3631 VSS.n3630 0.00442442
R9284 VSS.n3083 VSS.n3082 0.00442442
R9285 VSS.n2646 VSS.n2325 0.00442442
R9286 VSS.n2485 VSS.n2484 0.00429913
R9287 VSS.n2519 VSS.n2518 0.00429913
R9288 VSS.n3592 VSS.n3591 0.0042936
R9289 VSS.n3613 VSS.n3612 0.0042936
R9290 VSS.n1737 VSS.n1736 0.0042936
R9291 VSS.n3646 VSS.n3645 0.0042936
R9292 VSS.n3684 VSS.n3676 0.0042936
R9293 VSS.n3512 VSS.n3511 0.0042936
R9294 VSS.n3463 VSS.n3462 0.0042936
R9295 VSS.n3535 VSS.n3534 0.0042936
R9296 VSS.n3227 VSS.n3226 0.0042936
R9297 VSS.n3225 VSS.n3224 0.0042936
R9298 VSS.n3085 VSS.n3084 0.0042936
R9299 VSS.n3046 VSS.n3045 0.0042936
R9300 VSS.n2571 VSS.n2570 0.0042936
R9301 VSS.n2629 VSS.n2348 0.0042936
R9302 VSS.n2361 VSS.n2360 0.0042936
R9303 VSS.n2624 VSS.n2623 0.0042936
R9304 VSS.n2638 VSS.n2336 0.0042936
R9305 VSS.n2625 VSS.n2352 0.0042936
R9306 VSS.n2650 VSS.n2649 0.00427907
R9307 VSS.n826 VSS.n825 0.00427622
R9308 VSS.n850 VSS.n847 0.00427622
R9309 VSS.n5834 VSS.n5829 0.00426459
R9310 VSS.n2774 VSS.n2109 0.00426254
R9311 VSS.n3662 VSS.n3661 0.00416279
R9312 VSS.n3496 VSS.n3495 0.00416279
R9313 VSS.n3452 VSS.n3451 0.00416279
R9314 VSS.n81 VSS.n80 0.00414865
R9315 VSS.n2134 VSS.n2115 0.00411204
R9316 VSS.n2239 VSS.n2227 0.00411204
R9317 VSS.n3587 VSS.n3586 0.00403198
R9318 VSS.n3597 VSS.n3596 0.00403198
R9319 VSS.n3599 VSS.n3598 0.00403198
R9320 VSS.n3601 VSS.n3600 0.00403198
R9321 VSS.n3231 VSS.n3230 0.00403198
R9322 VSS.n3163 VSS.n3162 0.00403198
R9323 VSS.n3097 VSS.n3096 0.00403198
R9324 VSS.n3066 VSS.n3065 0.00403198
R9325 VSS.n2640 VSS.n2333 0.00403198
R9326 VSS.n2122 VSS.n2121 0.00397826
R9327 VSS.n4168 VSS.n4167 0.00396895
R9328 VSS.n5294 VSS.n5293 0.00396154
R9329 VSS.n2705 VSS.n2224 0.00396154
R9330 VSS.n2517 VSS.n2452 0.00390611
R9331 VSS.n2515 VSS.n2455 0.00390611
R9332 VSS.n3731 VSS.n3730 0.00390116
R9333 VSS.n1739 VSS.n1738 0.00390116
R9334 VSS.n3728 VSS.n3727 0.00390116
R9335 VSS.n1733 VSS.n1732 0.00390116
R9336 VSS.n3466 VSS.n3465 0.00390116
R9337 VSS.n3460 VSS.n3459 0.00390116
R9338 VSS.n3538 VSS.n3537 0.00390116
R9339 VSS.n3532 VSS.n3531 0.00390116
R9340 VSS.n1788 VSS.n1787 0.00390116
R9341 VSS.n1784 VSS.n1783 0.00390116
R9342 VSS.n2346 VSS.n2345 0.00390116
R9343 VSS.n2628 VSS.n2627 0.00390116
R9344 VSS.n2355 VSS.n2351 0.00390116
R9345 VSS.n2616 VSS.n2365 0.00390116
R9346 VSS.n2695 VSS.n2694 0.00389623
R9347 VSS.n3847 VSS.n3846 0.00381797
R9348 VSS.n3849 VSS.n3848 0.00381797
R9349 VSS.n3868 VSS.n3867 0.00381797
R9350 VSS.n3870 VSS.n3869 0.00381797
R9351 VSS.n2773 VSS.n2110 0.00381104
R9352 VSS.n2737 VSS.n2736 0.00381104
R9353 VSS.n3609 VSS.n3608 0.00377035
R9354 VSS.n3657 VSS.n3656 0.00377035
R9355 VSS.n3504 VSS.n3503 0.00377035
R9356 VSS.n3528 VSS.n3527 0.00377035
R9357 VSS.n3524 VSS.n3523 0.00377035
R9358 VSS.n3522 VSS.n3521 0.00377035
R9359 VSS.n3519 VSS.n3518 0.00377035
R9360 VSS.n3492 VSS.n3491 0.00377035
R9361 VSS.n3482 VSS.n3481 0.00377035
R9362 VSS.n5083 VSS.n5069 0.00371429
R9363 VSS.n3277 VSS.n3276 0.00367919
R9364 VSS.n3789 VSS.n3774 0.00367016
R9365 VSS.n3807 VSS.n3806 0.00367016
R9366 VSS.n2106 VSS.n2102 0.00366054
R9367 VSS.n2769 VSS.n2768 0.00366054
R9368 VSS.n2182 VSS.n2169 0.00366054
R9369 VSS.n2701 VSS.n2235 0.00366054
R9370 VSS.n2285 VSS.n2247 0.00366054
R9371 VSS.n2703 VSS.n2702 0.00366054
R9372 VSS.n4026 VSS.n4020 0.00364685
R9373 VSS.n4016 VSS.n4013 0.00364685
R9374 VSS.n2559 VSS.n2414 0.0036441
R9375 VSS.n2558 VSS.n2557 0.0036441
R9376 VSS.n3607 VSS.n3606 0.00363953
R9377 VSS.n3693 VSS.n3692 0.00363953
R9378 VSS.n3699 VSS.n3698 0.00363953
R9379 VSS.n3213 VSS.n3211 0.00363953
R9380 VSS.n3102 VSS.n3101 0.00363953
R9381 VSS.n2639 VSS.n2335 0.00363953
R9382 VSS.n3896 VSS.n3895 0.00356977
R9383 VSS.n5825 VSS.n5824 0.00354348
R9384 VSS.n3425 VSS.n3424 0.00352326
R9385 VSS.n2108 VSS.n2107 0.00351003
R9386 VSS.n2234 VSS.n2233 0.00351003
R9387 VSS.n2704 VSS.n2229 0.00351003
R9388 VSS.n2683 VSS.n2254 0.00351003
R9389 VSS.n2672 VSS.n2272 0.00351003
R9390 VSS.n1731 VSS.n1730 0.00350872
R9391 VSS.n3513 VSS.n3512 0.00350872
R9392 VSS.n3554 VSS.n3553 0.00350872
R9393 VSS.n3385 VSS.n3384 0.00350872
R9394 VSS.n2620 VSS.n2363 0.00350872
R9395 VSS.n2632 VSS.n2342 0.00350872
R9396 VSS.n2619 VSS.n2618 0.00350872
R9397 VSS.n3893 VSS.n3892 0.00347674
R9398 VSS.n732 VSS.n729 0.0034717
R9399 VSS.n504 VSS.n498 0.0034717
R9400 VSS.n770 VSS.n767 0.0034717
R9401 VSS.n4276 VSS.n4275 0.0034717
R9402 VSS.n4309 VSS.n4299 0.0034717
R9403 VSS.n1948 VSS.n1947 0.00344828
R9404 VSS.n2357 VSS.n2353 0.00340698
R9405 VSS.n3485 VSS.n3484 0.00337791
R9406 VSS.n3477 VSS.n3476 0.00337791
R9407 VSS.n3557 VSS.n3556 0.00337791
R9408 VSS.n3549 VSS.n3548 0.00337791
R9409 VSS.n2851 VSS.n2027 0.00335953
R9410 VSS.n2191 VSS.n2176 0.00335953
R9411 VSS.n2174 VSS.n2172 0.00335953
R9412 VSS.n2777 VSS.n2776 0.00335953
R9413 VSS.n3752 VSS.n3740 0.0032972
R9414 VSS.n3771 VSS.n3770 0.0032972
R9415 VSS.n3886 VSS.n3885 0.0032907
R9416 VSS.n3892 VSS.n3891 0.0032907
R9417 VSS.n3915 VSS.n3914 0.00327533
R9418 VSS.n3845 VSS.n3844 0.00324751
R9419 VSS.n3876 VSS.n3875 0.00324751
R9420 VSS.n3873 VSS.n3872 0.00324751
R9421 VSS.n3236 VSS.n3235 0.00324709
R9422 VSS.n3168 VSS.n3167 0.00324709
R9423 VSS.n2638 VSS.n2337 0.00324709
R9424 VSS.n1804 VSS.n1803 0.00322727
R9425 VSS.n2189 VSS.n2178 0.00320903
R9426 VSS.n2779 VSS.n2778 0.00320903
R9427 VSS.n2188 VSS.n2187 0.00320903
R9428 VSS.n2691 VSS.n2690 0.00320903
R9429 VSS.n3878 VSS.n3877 0.00319767
R9430 VSS.n3884 VSS.n3883 0.00319767
R9431 VSS.n3889 VSS.n3888 0.00319767
R9432 VSS.n2873 VSS.n1992 0.00317559
R9433 VSS.n2871 VSS.n1999 0.00317559
R9434 VSS.n2864 VSS.n2863 0.00317559
R9435 VSS.n2033 VSS.n2032 0.00317559
R9436 VSS.n2793 VSS.n2090 0.00317559
R9437 VSS.n3852 VSS.n3851 0.00317281
R9438 VSS.n3856 VSS.n3855 0.00317281
R9439 VSS.n3861 VSS.n3860 0.00317281
R9440 VSS.n3865 VSS.n3864 0.00317281
R9441 VSS.n4690 VSS.n4682 0.00316667
R9442 VSS.n3191 VSS.n3190 0.00315896
R9443 VSS.n5902 VSS 0.00314706
R9444 VSS.n878 VSS.n877 0.00313878
R9445 VSS.n1861 VSS.n1860 0.00313793
R9446 VSS.n1859 VSS.n1858 0.00313793
R9447 VSS.n1858 VSS.n1856 0.00313793
R9448 VSS.n1856 VSS.n1855 0.00313793
R9449 VSS.n1852 VSS.n1851 0.00313793
R9450 VSS.n1849 VSS.n1848 0.00313793
R9451 VSS.n1846 VSS.n1845 0.00313793
R9452 VSS.n1947 VSS.n1945 0.00313793
R9453 VSS.n1923 VSS.n1922 0.00313793
R9454 VSS.n2526 VSS.n2444 0.00312009
R9455 VSS.n3286 VSS.n3285 0.00311628
R9456 VSS.n3292 VSS.n3291 0.00311628
R9457 VSS.n3220 VSS.n3219 0.00311628
R9458 VSS.n3076 VSS.n3075 0.00311628
R9459 VSS.n3129 VSS.n3124 0.00311628
R9460 VSS.n2634 VSS.n2633 0.00311628
R9461 VSS.n2882 VSS.n1992 0.0031087
R9462 VSS.n2872 VSS.n2871 0.0031087
R9463 VSS.n2864 VSS.n2009 0.0031087
R9464 VSS.n2032 VSS.n2010 0.0031087
R9465 VSS.n2090 VSS.n2086 0.0031087
R9466 VSS.n3881 VSS.n3880 0.00310465
R9467 VSS.n2783 VSS.n2091 0.00307649
R9468 VSS.n2121 VSS.n2112 0.00307649
R9469 VSS.n2727 VSS.n2726 0.00307649
R9470 VSS.n2854 VSS.n2022 0.00305853
R9471 VSS.n2800 VSS.n2797 0.00305853
R9472 VSS.n2038 VSS.n2023 0.00305853
R9473 VSS.n2853 VSS.n2024 0.00305853
R9474 VSS.n2843 VSS.n2024 0.00305853
R9475 VSS.n2843 VSS.n2842 0.00305853
R9476 VSS.n2828 VSS.n2827 0.00305853
R9477 VSS.n2799 VSS.n2798 0.00305853
R9478 VSS.n2816 VSS.n2815 0.00305853
R9479 VSS.n2852 VSS.n2026 0.00305853
R9480 VSS.n2079 VSS.n2073 0.00305853
R9481 VSS.n2851 VSS.n2028 0.00305853
R9482 VSS.n2823 VSS.n2074 0.00305853
R9483 VSS.n2775 VSS.n2774 0.00305853
R9484 VSS.n2295 VSS.n2284 0.00305853
R9485 VSS.n2297 VSS.n2296 0.00305853
R9486 VSS.n2300 VSS.n2297 0.00305853
R9487 VSS.n2301 VSS.n2300 0.00305853
R9488 VSS.n2306 VSS.n2305 0.00305853
R9489 VSS.n2253 VSS.n2252 0.00305853
R9490 VSS.n2299 VSS.n2253 0.00305853
R9491 VSS.n2304 VSS.n2275 0.00305853
R9492 VSS.n2684 VSS.n2683 0.00305853
R9493 VSS.n3810 VSS.n3809 0.00301748
R9494 VSS.n3841 VSS.n3840 0.00301748
R9495 VSS.n2716 VSS.n2209 0.00301572
R9496 VSS.n2714 VSS.n2216 0.00301572
R9497 VSS.n2660 VSS.n2316 0.00301572
R9498 VSS.n2792 VSS.n2091 0.00301208
R9499 VSS.n2782 VSS.n2781 0.00301208
R9500 VSS.n2727 VSS.n2208 0.00301208
R9501 VSS.n2534 VSS.n2436 0.00298908
R9502 VSS.n3144 VSS.n3143 0.00298547
R9503 VSS.n3037 VSS.n3031 0.00298547
R9504 VSS.n2579 VSS.n2568 0.00298547
R9505 VSS.n2604 VSS.n2390 0.00298547
R9506 VSS.n2578 VSS.n2577 0.00298547
R9507 VSS.n2592 VSS.n2591 0.00298547
R9508 VSS.n2576 VSS.n2399 0.00298547
R9509 VSS.n2596 VSS.n2394 0.00298547
R9510 VSS.n1860 VSS.n1859 0.00298276
R9511 VSS.n1855 VSS.n1854 0.00298276
R9512 VSS.n1920 VSS.n1919 0.00298276
R9513 VSS.n4507 VSS.n4506 0.00297253
R9514 VSS.n5074 VSS.n5073 0.00297253
R9515 VSS.n2725 VSS.n2209 0.00295283
R9516 VSS.n2715 VSS.n2714 0.00295283
R9517 VSS.n2694 VSS.n2693 0.00295283
R9518 VSS.n3838 VSS.n3826 0.00292424
R9519 VSS.n2795 VSS.n2089 0.00292012
R9520 VSS.n2662 VSS.n2309 0.00292012
R9521 VSS.n2853 VSS.n2023 0.00290803
R9522 VSS.n2842 VSS.n2047 0.00290803
R9523 VSS.n2852 VSS.n2025 0.00290803
R9524 VSS.n2819 VSS.n2078 0.00290803
R9525 VSS.n2308 VSS.n2307 0.00290803
R9526 VSS.n2296 VSS.n2291 0.00290803
R9527 VSS.n2305 VSS.n2302 0.00290803
R9528 VSS.n2306 VSS.n2277 0.00290803
R9529 VSS.n2664 VSS.n2283 0.00290803
R9530 VSS.n2290 VSS.n2252 0.00290803
R9531 VSS.n2670 VSS.n2275 0.00290803
R9532 VSS.n2672 VSS.n2671 0.00290803
R9533 VSS.n2863 VSS.n2010 0.00290803
R9534 VSS.n3589 VSS.n3580 0.0028968
R9535 VSS.n3509 VSS.n3508 0.0028968
R9536 VSS.n3859 VSS.n3858 0.00289631
R9537 VSS.n3590 VSS.n3589 0.00289361
R9538 VSS.n3510 VSS.n3509 0.00289361
R9539 VSS.n299 VSS.n298 0.00287973
R9540 VSS.n3392 VSS.n3391 0.00285465
R9541 VSS.n3314 VSS.n3304 0.00285465
R9542 VSS.n2835 VSS.n2834 0.00284114
R9543 VSS.n4162 VSS.n889 0.00283689
R9544 VSS.n4709 VSS 0.00283333
R9545 VSS.n1924 VSS.n1923 0.00282759
R9546 VSS.n2650 VSS.n2317 0.00282558
R9547 VSS.n2353 VSS.n2338 0.00282558
R9548 VSS.n2584 VSS.n2564 0.00282558
R9549 VSS.n3069 VSS.n3054 0.00282558
R9550 VSS.n3052 VSS.n3051 0.00282558
R9551 VSS.n3049 VSS.n3041 0.00282558
R9552 VSS.n3015 VSS.n3004 0.00282558
R9553 VSS.n2962 VSS.n2916 0.00282558
R9554 VSS.n3435 VSS.n3434 0.00282558
R9555 VSS.n3423 VSS.n3422 0.00282558
R9556 VSS.n3623 VSS.n3574 0.00281884
R9557 VSS.n3240 VSS.n3200 0.00281214
R9558 VSS.n3198 VSS.n3191 0.00281214
R9559 VSS.n3171 VSS.n3158 0.00281214
R9560 VSS.n3131 VSS.n3118 0.00281214
R9561 VSS.n3090 VSS.n3072 0.00281214
R9562 VSS.n3359 VSS.n3358 0.00281214
R9563 VSS.n3275 VSS.n3262 0.00281214
R9564 VSS.n4374 VSS.n4372 0.00280769
R9565 VSS.n3087 VSS.n3086 0.00278682
R9566 VSS.n2552 VSS.n2551 0.00278571
R9567 VSS.n2538 VSS.n2433 0.00278571
R9568 VSS.n2659 VSS.n2317 0.00276744
R9569 VSS.n2649 VSS.n2648 0.00276744
R9570 VSS.n2585 VSS.n2584 0.00276744
R9571 VSS.n3070 VSS.n3069 0.00276744
R9572 VSS.n3053 VSS.n3052 0.00276744
R9573 VSS.n3050 VSS.n3049 0.00276744
R9574 VSS.n2963 VSS.n2962 0.00276744
R9575 VSS.n3573 VSS.n3572 0.00276744
R9576 VSS.n3572 VSS.n3571 0.00276744
R9577 VSS.n3570 VSS.n3569 0.00276744
R9578 VSS.n3568 VSS.n3567 0.00276744
R9579 VSS.n3424 VSS.n3423 0.00276744
R9580 VSS.n3723 VSS.n3722 0.00276087
R9581 VSS.n3686 VSS.n3685 0.00276087
R9582 VSS.n3624 VSS.n3623 0.00276087
R9583 VSS.n2824 VSS.n2823 0.00275752
R9584 VSS.n2780 VSS.n2100 0.00275752
R9585 VSS.n2692 VSS.n2245 0.00275752
R9586 VSS.n3241 VSS.n3240 0.00275434
R9587 VSS.n3199 VSS.n3198 0.00275434
R9588 VSS.n3117 VSS.n3116 0.00275434
R9589 VSS.n3415 VSS.n3414 0.00275434
R9590 VSS.n3276 VSS.n3275 0.00275434
R9591 VSS.n2563 VSS.n2410 0.00272857
R9592 VSS.n2433 VSS.n2421 0.00272857
R9593 VSS.n2484 VSS.n2439 0.00272707
R9594 VSS.n2531 VSS.n2430 0.00272707
R9595 VSS.n2450 VSS.n2440 0.00272707
R9596 VSS.n2527 VSS.n2442 0.00272707
R9597 VSS.n2497 VSS.n2496 0.00272707
R9598 VSS.n3468 VSS.n3467 0.00272384
R9599 VSS.n3130 VSS.n3119 0.00272384
R9600 VSS.n2934 VSS.n2933 0.00272384
R9601 VSS.n2938 VSS.n2936 0.00272384
R9602 VSS.n2939 VSS.n2938 0.00272384
R9603 VSS.n2940 VSS.n2939 0.00272384
R9604 VSS.n2945 VSS.n2944 0.00272384
R9605 VSS.n2950 VSS.n2948 0.00272384
R9606 VSS.n2954 VSS.n2953 0.00272384
R9607 VSS VSS.n5879 0.00272222
R9608 VSS.n5801 VSS 0.00272222
R9609 VSS.n5818 VSS 0.00272222
R9610 VSS.n1980 VSS.n1979 0.00270985
R9611 VSS.n1456 VSS.n1455 0.0027028
R9612 VSS.n1456 VSS.n1417 0.0027028
R9613 VSS.n1462 VSS.n1417 0.0027028
R9614 VSS VSS.n1414 0.0027028
R9615 VSS VSS.n1414 0.0027028
R9616 VSS VSS.n835 0.0027028
R9617 VSS.n835 VSS 0.0027028
R9618 VSS.n2225 VSS.n2216 0.00270126
R9619 VSS.n729 VSS.n716 0.00269512
R9620 VSS.n4053 VSS.n4050 0.00269512
R9621 VSS.n2749 VSS.n2162 0.00269002
R9622 VSS.n1882 VSS.n1881 0.00267241
R9623 VSS.n1944 VSS.n1943 0.00267241
R9624 VSS.n1941 VSS.n1940 0.00267241
R9625 VSS.n1891 VSS.n1890 0.00267241
R9626 VSS.n1903 VSS.n1902 0.00267241
R9627 VSS.n1950 VSS.n1949 0.00267241
R9628 VSS.n1935 VSS.n1934 0.00267241
R9629 VSS.n1928 VSS.n1927 0.00267241
R9630 VSS.n1918 VSS.n1917 0.00267241
R9631 VSS.n4111 VSS.n908 0.00266
R9632 VSS.n3437 VSS.n3436 0.00265116
R9633 VSS.n3426 VSS.n3425 0.00265116
R9634 VSS.n4754 VSS.n4753 0.00262598
R9635 VSS.n5896 VSS.n4755 0.00262598
R9636 VSS.n5895 VSS.n5894 0.00262598
R9637 VSS.n5893 VSS.n5892 0.00262598
R9638 VSS.n5891 VSS.n5890 0.00262598
R9639 VSS.n2762 VSS.n2122 0.0026256
R9640 VSS.n2039 VSS.n2037 0.00260702
R9641 VSS.n2845 VSS.n2026 0.00260702
R9642 VSS.n2841 VSS.n2046 0.00260702
R9643 VSS.n2829 VSS.n2066 0.00260702
R9644 VSS.n2814 VSS.n2081 0.00260702
R9645 VSS.n2042 VSS.n2041 0.00260702
R9646 VSS.n2839 VSS.n2049 0.00260702
R9647 VSS.n2831 VSS.n2064 0.00260702
R9648 VSS.n2812 VSS.n2084 0.00260702
R9649 VSS.n2773 VSS.n2104 0.00260702
R9650 VSS.n2298 VSS.n2269 0.00260702
R9651 VSS.n2689 VSS.n2688 0.00260702
R9652 VSS.n2685 VSS.n2684 0.00260702
R9653 VSS.n2680 VSS.n2679 0.00260702
R9654 VSS.n2531 VSS.n2530 0.00259607
R9655 VSS.n2505 VSS.n2504 0.00259607
R9656 VSS.n2532 VSS.n2438 0.00259607
R9657 VSS.n2479 VSS.n2475 0.00259607
R9658 VSS.n2501 VSS.n2476 0.00259607
R9659 VSS.n2497 VSS.n2477 0.00259607
R9660 VSS.n3388 VSS.n3387 0.00259302
R9661 VSS.n3222 VSS.n3221 0.00259302
R9662 VSS.n3136 VSS.n3135 0.00259302
R9663 VSS.n2936 VSS.n2934 0.00259302
R9664 VSS.n2942 VSS.n2940 0.00259302
R9665 VSS.n3036 VSS.n3035 0.00259302
R9666 VSS.n2980 VSS.n2979 0.00259302
R9667 VSS.n2603 VSS.n2602 0.00259302
R9668 VSS.n2590 VSS.n2402 0.00259302
R9669 VSS.n2393 VSS.n2392 0.00259302
R9670 VSS.n2588 VSS.n2407 0.00259302
R9671 VSS.n3051 VSS.n3050 0.00259302
R9672 VSS.n3637 VSS.n3626 0.00258696
R9673 VSS.n3116 VSS.n3105 0.00258092
R9674 VSS.n3414 VSS.n3361 0.00258092
R9675 VSS.n2553 VSS.n2420 0.00255714
R9676 VSS.n1812 VSS.n1811 0.00254545
R9677 VSS.n3649 VSS.n3648 0.00252899
R9678 VSS.n2912 VSS.n2911 0.00252532
R9679 VSS.n2909 VSS.n2908 0.00252532
R9680 VSS.n2906 VSS.n2905 0.00252532
R9681 VSS.n2884 VSS.n2883 0.00252532
R9682 VSS.n3154 VSS.n3147 0.00252312
R9683 VSS.n3104 VSS.n3103 0.00252312
R9684 VSS.n3360 VSS.n3359 0.00252312
R9685 VSS.n3261 VSS.n3260 0.00252312
R9686 VSS.n3259 VSS.n3252 0.00252312
R9687 VSS.n3243 VSS.n3242 0.00252312
R9688 VSS.n1847 VSS.n1846 0.00251724
R9689 VSS.n1905 VSS.n1904 0.00251724
R9690 VSS.n2913 VSS.n2912 0.00247468
R9691 VSS.n2910 VSS.n2909 0.00247468
R9692 VSS.n2907 VSS.n2906 0.00247468
R9693 VSS.n2897 VSS.n2896 0.00247468
R9694 VSS.n2885 VSS.n2884 0.00247468
R9695 VSS.n3722 VSS.n3713 0.00247101
R9696 VSS.n3391 VSS.n3390 0.00246221
R9697 VSS.n3307 VSS.n3306 0.00246221
R9698 VSS.n3311 VSS.n3308 0.00246221
R9699 VSS.n3303 VSS.n3302 0.00246221
R9700 VSS.n3204 VSS.n3203 0.00246221
R9701 VSS.n2998 VSS.n2990 0.00246221
R9702 VSS.n2816 VSS.n2080 0.00245652
R9703 VSS.n2840 VSS.n2048 0.00245652
R9704 VSS.n2818 VSS.n2817 0.00245652
R9705 VSS.n2179 VSS.n2177 0.00245652
R9706 VSS.n2107 VSS.n2106 0.00245652
R9707 VSS.n2185 VSS.n2184 0.00245652
R9708 VSS.n2190 VSS.n2189 0.00245652
R9709 VSS.n2733 VSS.n2176 0.00245652
R9710 VSS.n2105 VSS.n2103 0.00245652
R9711 VSS.n2188 VSS.n2171 0.00245652
R9712 VSS.n2738 VSS.n2169 0.00245652
R9713 VSS.n2293 VSS.n2292 0.00245652
R9714 VSS.n2233 VSS.n2232 0.00245652
R9715 VSS.n2235 VSS.n2234 0.00245652
R9716 VSS.n2701 VSS.n2700 0.00245652
R9717 VSS.n2286 VSS.n2285 0.00245652
R9718 VSS.n2704 VSS.n2703 0.00245652
R9719 VSS.n2287 VSS.n2248 0.00245652
R9720 VSS.n2303 VSS.n2270 0.00245652
R9721 VSS.n2666 VSS.n2665 0.00245652
R9722 VSS.n2705 VSS.n2227 0.00245652
R9723 VSS.n2676 VSS.n2675 0.00245652
R9724 VSS.n2668 VSS.n2667 0.00245652
R9725 VSS.n2313 VSS.n2279 0.00245652
R9726 VSS.n5889 VSS.n5888 0.00244245
R9727 VSS.n5887 VSS.n4750 0.00244245
R9728 VSS.n5921 VSS.n5920 0.00244245
R9729 VSS.n5914 VSS.n5913 0.00244245
R9730 VSS.n2033 VSS.n2029 0.0024398
R9731 VSS VSS.n826 0.00238811
R9732 VSS.n1850 VSS.n1849 0.00236207
R9733 VSS.n3687 VSS.n3686 0.00235507
R9734 VSS.n2489 VSS.n2488 0.00233406
R9735 VSS.n2533 VSS.n2437 0.00233406
R9736 VSS.n2481 VSS.n2479 0.00233406
R9737 VSS.n2535 VSS.n2435 0.00233406
R9738 VSS.n3381 VSS.n3380 0.0023314
R9739 VSS.n3294 VSS.n3293 0.0023314
R9740 VSS.n3127 VSS.n3126 0.0023314
R9741 VSS.n3170 VSS.n3160 0.0023314
R9742 VSS.n3034 VSS.n3033 0.0023314
R9743 VSS.n3022 VSS.n3021 0.0023314
R9744 VSS.n2993 VSS.n2992 0.0023314
R9745 VSS.n2971 VSS.n2970 0.0023314
R9746 VSS.n3030 VSS.n3029 0.0023314
R9747 VSS.n2987 VSS.n2986 0.0023314
R9748 VSS.n2978 VSS.n2977 0.0023314
R9749 VSS.n2596 VSS.n2595 0.0023314
R9750 VSS.n2908 VSS.n2907 0.00232278
R9751 VSS.n2798 VSS.n2069 0.00230602
R9752 VSS.n2073 VSS.n2070 0.00230602
R9753 VSS.n2114 VSS.n2113 0.00230602
R9754 VSS.n2009 VSS.n1999 0.00230602
R9755 VSS.n2761 VSS.n2123 0.00230354
R9756 VSS.n3663 VSS.n3652 0.0022971
R9757 VSS.n2491 VSS.n2490 0.00224426
R9758 VSS.n2648 VSS.n2647 0.00224419
R9759 VSS.n5291 VSS.n5290 0.00224148
R9760 VSS.n1879 VSS.n1874 0.00222181
R9761 VSS.n1945 VSS.n1938 0.0022069
R9762 VSS.n2530 VSS.n2529 0.00220306
R9763 VSS.n2504 VSS.n2474 0.00220306
R9764 VSS.n2506 VSS.n2473 0.00220306
R9765 VSS.n2503 VSS.n2502 0.00220306
R9766 VSS.n2492 VSS.n2482 0.00220306
R9767 VSS.n2508 VSS.n2471 0.00220306
R9768 VSS.n3400 VSS.n3399 0.00220058
R9769 VSS.n3397 VSS.n3396 0.00220058
R9770 VSS.n3394 VSS.n3393 0.00220058
R9771 VSS.n3221 VSS.n3220 0.00220058
R9772 VSS.n3177 VSS.n3176 0.00220058
R9773 VSS.n3138 VSS.n3137 0.00220058
R9774 VSS.n2953 VSS.n2952 0.00220058
R9775 VSS.n3011 VSS.n3008 0.00220058
R9776 VSS.n2973 VSS.n2972 0.00220058
R9777 VSS.n2340 VSS.n2339 0.00220058
R9778 VSS.n2601 VSS.n2600 0.00220058
R9779 VSS.n1643 VSS.n1642 0.0022002
R9780 VSS.n2242 VSS.n2226 0.00219811
R9781 VSS.n2790 VSS.n2093 0.00219111
R9782 VSS.n2723 VSS.n2211 0.00219111
R9783 VSS.n2637 VSS.n2326 0.00218605
R9784 VSS.n2358 VSS.n2357 0.00218605
R9785 VSS.n2367 VSS.n2359 0.00218605
R9786 VSS.n2614 VSS.n2371 0.00218605
R9787 VSS.n3041 VSS.n3040 0.00218605
R9788 VSS.n3421 VSS.n3420 0.00218605
R9789 VSS.n3419 VSS.n3418 0.00218605
R9790 VSS.n3417 VSS.n3416 0.00218605
R9791 VSS.n3737 VSS.n3736 0.00218116
R9792 VSS.n3735 VSS.n3726 0.00218116
R9793 VSS.n3725 VSS.n3724 0.00218116
R9794 VSS.n3685 VSS.n3669 0.00218116
R9795 VSS.n3190 VSS.n3189 0.0021763
R9796 VSS.n3188 VSS.n3187 0.0021763
R9797 VSS.n5198 VSS.n5197 0.00216667
R9798 VSS.n5235 VSS.n4803 0.00216667
R9799 VSS.n5225 VSS.n5224 0.00216667
R9800 VSS.n5248 VSS.n5245 0.00216667
R9801 VSS.n2513 VSS.n2457 0.00215714
R9802 VSS.n2847 VSS.n2028 0.00215552
R9803 VSS.n2282 VSS.n2277 0.00215552
R9804 VSS.n6075 VSS.n6074 0.00214634
R9805 VSS.n2707 VSS.n2706 0.00213522
R9806 VSS.n3667 VSS.n3666 0.00212319
R9807 VSS.n3157 VSS.n3156 0.0021185
R9808 VSS.n2111 VSS.n2098 0.00211031
R9809 VSS.n2203 VSS.n2170 0.00211031
R9810 VSS.n2451 VSS.n2450 0.00207205
R9811 VSS.n3401 VSS.n3400 0.00206977
R9812 VSS.n3398 VSS.n3397 0.00206977
R9813 VSS.n3395 VSS.n3394 0.00206977
R9814 VSS.n3335 VSS.n3334 0.00206977
R9815 VSS.n2948 VSS.n2946 0.00206977
R9816 VSS.n2997 VSS.n2996 0.00206977
R9817 VSS.n3054 VSS.n3053 0.00206977
R9818 VSS.n3688 VSS.n3687 0.00206522
R9819 VSS.n2561 VSS.n2412 0.0020629
R9820 VSS.n3449 VSS.n3448 0.00206165
R9821 VSS.n3412 VSS.n3407 0.00206165
R9822 VSS.n3238 VSS.n3233 0.00206165
R9823 VSS.n2657 VSS.n2319 0.00206165
R9824 VSS.n1910 VSS.n1909 0.0020532
R9825 VSS.n1933 VSS.n1932 0.00205172
R9826 VSS.n2488 VSS.n2487 0.00204803
R9827 VSS.n2487 VSS.n2483 0.00204706
R9828 VSS.n2741 VSS.n2740 0.00204589
R9829 VSS.n2729 VSS.n2195 0.00202155
R9830 VSS.n2838 VSS.n2050 0.00200502
R9831 VSS.n2180 VSS.n2165 0.00200502
R9832 VSS.n2735 VSS.n2734 0.00200502
R9833 VSS.n2744 VSS.n2743 0.00200502
R9834 VSS.n2199 VSS.n2173 0.00200502
R9835 VSS.n2664 VSS.n2663 0.00200502
R9836 VSS.n2228 VSS.n2222 0.00200502
R9837 VSS.n2699 VSS.n2236 0.00200502
R9838 VSS.n2709 VSS.n2708 0.00200502
R9839 VSS.n2697 VSS.n2240 0.00200502
R9840 VSS.n2880 VSS.n1994 0.00199156
R9841 VSS.n2850 VSS.n2043 0.00197157
R9842 VSS.n2905 VSS.n2904 0.00196835
R9843 VSS.n3433 VSS.n3432 0.00195349
R9844 VSS.n1559 VSS.n1558 0.00195161
R9845 VSS.n1571 VSS.n1569 0.00195161
R9846 VSS.n1573 VSS.n1572 0.00195161
R9847 VSS.n1575 VSS.n1574 0.00195161
R9848 VSS.n1581 VSS.n1580 0.00195161
R9849 VSS.n1591 VSS.n1590 0.00195161
R9850 VSS.n1601 VSS.n1600 0.00195161
R9851 VSS.n2682 VSS.n2681 0.00194654
R9852 VSS.n2674 VSS.n2673 0.00194654
R9853 VSS.n3173 VSS.n3172 0.00194509
R9854 VSS.n3555 VSS.n3554 0.00193895
R9855 VSS.n3551 VSS.n3550 0.00193895
R9856 VSS.n3540 VSS.n3539 0.00193895
R9857 VSS.n3386 VSS.n3385 0.00193895
R9858 VSS.n3288 VSS.n3287 0.00193895
R9859 VSS.n3353 VSS.n3345 0.00193895
R9860 VSS.n3027 VSS.n3026 0.00193895
R9861 VSS.n2578 VSS.n2403 0.00193895
R9862 VSS.n2401 VSS.n2399 0.00193895
R9863 VSS.n2772 VSS.n2771 0.00191707
R9864 VSS.n5329 VSS.n5326 0.00189535
R9865 VSS.n5423 VSS.n5331 0.00189535
R9866 VSS.n3620 VSS.n3619 0.00188813
R9867 VSS.n2959 VSS.n2958 0.00188813
R9868 VSS.n2581 VSS.n2567 0.00188813
R9869 VSS.n3103 VSS.n3092 0.00188728
R9870 VSS.n2911 VSS.n2910 0.00186709
R9871 VSS.n356 VSS.n353 0.00185388
R9872 VSS.n2770 VSS.n2112 0.00185266
R9873 VSS.n3431 VSS.n3430 0.00183721
R9874 VSS.n3724 VSS.n3723 0.00183333
R9875 VSS.n3091 VSS.n3090 0.00182948
R9876 VSS.n3278 VSS.n3277 0.00182948
R9877 VSS.n4370 VSS.n4361 0.0018278
R9878 VSS.n2525 VSS.n2524 0.00181429
R9879 VSS.n2560 VSS.n2559 0.00181004
R9880 VSS.n2441 VSS.n2438 0.00181004
R9881 VSS.n3701 VSS.n3700 0.00180814
R9882 VSS.n3389 VSS.n3388 0.00180814
R9883 VSS.n3350 VSS.n3349 0.00180814
R9884 VSS.n3324 VSS.n3323 0.00180814
R9885 VSS.n3344 VSS.n3343 0.00180814
R9886 VSS.n3331 VSS.n3330 0.00180814
R9887 VSS.n3211 VSS.n3210 0.00180814
R9888 VSS.n3179 VSS.n3178 0.00180814
R9889 VSS.n3142 VSS.n3141 0.00180814
R9890 VSS.n3100 VSS.n3099 0.00180814
R9891 VSS.n3014 VSS.n3006 0.00180814
R9892 VSS.n2572 VSS.n2363 0.00180814
R9893 VSS.n2575 VSS.n2390 0.00180814
R9894 VSS.n2395 VSS.n2391 0.00180814
R9895 VSS.n5816 VSS.n5803 0.00180435
R9896 VSS.n2612 VSS.n2611 0.00177907
R9897 VSS.n3039 VSS.n3038 0.00177907
R9898 VSS.n3428 VSS.n3427 0.00177907
R9899 VSS.n3133 VSS.n3132 0.00177168
R9900 VSS.n3299 VSS.n3296 0.00177168
R9901 VSS.n2820 VSS.n2077 0.0017709
R9902 VSS.n3760 VSS.n3759 0.00176168
R9903 VSS.n3836 VSS.n3829 0.00176168
R9904 VSS.n1513 VSS.n1405 0.00175874
R9905 VSS.n2536 VSS.n2434 0.00175714
R9906 VSS.n1579 VSS.n1577 0.00174752
R9907 VSS.n1619 VSS.n1618 0.00174424
R9908 VSS.n1631 VSS.n1630 0.00174424
R9909 VSS.n2637 VSS.n2636 0.00172093
R9910 VSS.n3712 VSS.n3711 0.00171739
R9911 VSS.n3158 VSS.n3157 0.00171387
R9912 VSS.n2670 VSS.n2669 0.00170401
R9913 VSS.n2822 VSS.n2076 0.00170401
R9914 VSS.n2312 VSS.n2311 0.00169497
R9915 VSS.n5862 VSS 0.00168421
R9916 VSS.n2426 VSS.n2414 0.00167904
R9917 VSS.n2521 VSS.n2449 0.00167904
R9918 VSS.n3584 VSS.n3583 0.00167733
R9919 VSS.n3606 VSS.n3605 0.00167733
R9920 VSS.n3608 VSS.n3607 0.00167733
R9921 VSS.n3610 VSS.n3609 0.00167733
R9922 VSS.n3709 VSS.n3705 0.00167733
R9923 VSS.n3529 VSS.n3528 0.00167733
R9924 VSS.n3396 VSS.n3395 0.00167733
R9925 VSS.n3348 VSS.n3347 0.00167733
R9926 VSS.n3328 VSS.n3327 0.00167733
R9927 VSS.n3326 VSS.n3325 0.00167733
R9928 VSS.n3342 VSS.n3341 0.00167733
R9929 VSS.n3333 VSS.n3332 0.00167733
R9930 VSS.n2635 VSS.n2338 0.00166279
R9931 VSS.n2771 VSS.n2770 0.00165942
R9932 VSS.n2161 VSS.n2160 0.00165942
R9933 VSS.n3316 VSS.n3315 0.00165607
R9934 VSS.n2498 VSS.n2478 0.00164286
R9935 VSS.n2043 VSS.n2029 0.00163712
R9936 VSS.n2850 VSS.n2849 0.00163712
R9937 VSS.n2837 VSS.n2044 0.00163712
R9938 VSS.n2075 VSS.n2062 0.00163712
R9939 VSS.n2822 VSS.n2821 0.00163712
R9940 VSS.n2810 VSS.n2077 0.00163712
R9941 VSS.n3761 VSS.n3758 0.00163049
R9942 VSS.n2903 VSS.n2902 0.00161392
R9943 VSS.n188 VSS.n187 0.00161111
R9944 VSS.n218 VSS.n215 0.00161111
R9945 VSS.n205 VSS.n194 0.00161111
R9946 VSS.n195 VSS.n123 0.00161111
R9947 VSS.n2636 VSS.n2635 0.00160465
R9948 VSS.n2397 VSS.n2396 0.00160465
R9949 VSS.n2598 VSS.n2597 0.00160465
R9950 VSS.n2586 VSS.n2409 0.00160465
R9951 VSS.n2981 VSS.n2966 0.00160465
R9952 VSS.n3710 VSS.n3703 0.00160145
R9953 VSS.n4315 VSS.n4313 0.00159756
R9954 VSS.n2500 VSS.n2469 0.00158571
R9955 VSS.n2687 VSS.n2243 0.00156918
R9956 VSS.n2681 VSS.n2267 0.00156918
R9957 VSS.n2283 VSS.n2282 0.00155351
R9958 VSS.n2280 VSS.n2278 0.00155351
R9959 VSS.n2309 VSS.n2281 0.00155351
R9960 VSS.n3746 VSS.n3745 0.0015514
R9961 VSS.n3816 VSS.n3815 0.0015514
R9962 VSS.n3818 VSS.n3817 0.0015514
R9963 VSS.n3824 VSS.n3814 0.0015514
R9964 VSS.n2522 VSS.n2448 0.00154803
R9965 VSS.n1742 VSS.n1734 0.00154651
R9966 VSS.n3527 VSS.n3526 0.00154651
R9967 VSS.n3523 VSS.n3522 0.00154651
R9968 VSS.n3483 VSS.n3482 0.00154651
R9969 VSS.n3534 VSS.n3533 0.00154651
R9970 VSS.n3405 VSS.n3404 0.00154651
R9971 VSS.n3399 VSS.n3398 0.00154651
R9972 VSS.n3390 VSS.n3389 0.00154651
R9973 VSS.n3352 VSS.n3351 0.00154651
R9974 VSS.n3271 VSS.n3270 0.00154651
R9975 VSS.n3080 VSS.n3079 0.00154651
R9976 VSS.n3186 VSS.n3185 0.00154651
R9977 VSS.n3122 VSS.n3121 0.00154651
R9978 VSS.n2613 VSS.n2612 0.00154651
R9979 VSS.n3000 VSS.n2999 0.00154651
R9980 VSS.n3318 VSS.n3317 0.00154046
R9981 VSS.n1587 VSS.n1586 0.00153687
R9982 VSS.n1589 VSS.n1588 0.00153687
R9983 VSS.n1597 VSS.n1596 0.00153687
R9984 VSS.n1599 VSS.n1598 0.00153687
R9985 VSS.n1607 VSS.n1606 0.00153687
R9986 VSS.n2674 VSS.n2273 0.00150629
R9987 VSS.n2673 VSS.n2274 0.00150629
R9988 VSS.n2315 VSS.n2312 0.00150629
R9989 VSS.n1694 VSS.n1693 0.00150559
R9990 VSS.n1699 VSS.n1698 0.00150559
R9991 VSS.n1704 VSS.n1703 0.00150559
R9992 VSS.n1706 VSS.n1705 0.00150559
R9993 VSS.n2597 VSS.n2398 0.00148837
R9994 VSS.n3040 VSS.n3039 0.00148837
R9995 VSS.n3038 VSS.n3028 0.00148837
R9996 VSS.n3017 VSS.n3016 0.00148837
R9997 VSS.n3002 VSS.n3001 0.00148837
R9998 VSS.n2999 VSS.n2984 0.00148837
R9999 VSS.n2966 VSS.n2965 0.00148837
R10000 VSS.n3132 VSS.n3131 0.00148266
R10001 VSS.n3295 VSS.n3278 0.00148266
R10002 VSS.n2537 VSS.n2536 0.00147143
R10003 VSS.n2781 VSS.n2098 0.00146618
R10004 VSS.n2889 VSS.n2888 0.00146203
R10005 VSS.n1654 VSS.n1651 0.00145031
R10006 VSS.n1685 VSS.n1682 0.00144995
R10007 VSS.n1685 VSS.n1684 0.00144995
R10008 VSS.n1654 VSS.n1653 0.0014496
R10009 VSS VSS.n820 0.00144406
R10010 VSS.n2693 VSS.n2243 0.0014434
R10011 VSS.n2266 VSS.n2250 0.0014434
R10012 VSS.n1937 VSS.n1936 0.00143104
R10013 VSS.n2599 VSS.n2397 0.00143023
R10014 VSS.n3092 VSS.n3091 0.00142485
R10015 VSS.n3300 VSS.n3299 0.00142485
R10016 VSS.n2415 VSS.n2412 0.00141703
R10017 VSS.n2445 VSS.n2436 0.00141703
R10018 VSS.n2526 VSS.n2443 0.00141703
R10019 VSS.n3600 VSS.n3599 0.0014157
R10020 VSS.n3695 VSS.n3694 0.0014157
R10021 VSS.n3734 VSS.n3729 0.0014157
R10022 VSS.n3536 VSS.n3535 0.0014157
R10023 VSS.n3387 VSS.n3386 0.0014157
R10024 VSS.n1791 VSS.n1785 0.0014157
R10025 VSS.n2345 VSS.n2333 0.0014157
R10026 VSS.n2344 VSS.n2343 0.0014157
R10027 VSS.n2617 VSS.n2364 0.0014157
R10028 VSS.n2626 VSS.n2625 0.0014157
R10029 VSS.n2510 VSS.n2469 0.00141429
R10030 VSS.n2499 VSS.n2498 0.00141429
R10031 VSS.n2892 VSS.n2891 0.00141139
R10032 VSS.n2846 VSS.n2045 0.00140301
R10033 VSS.n2136 VSS.n2132 0.00140301
R10034 VSS.n2135 VSS.n2133 0.00140301
R10035 VSS.n2772 VSS.n2111 0.00140177
R10036 VSS.n1554 VSS.n1545 0.0014
R10037 VSS.n1552 VSS.n1547 0.0014
R10038 VSS.n1551 VSS.n1549 0.0014
R10039 VSS.n1667 VSS.n1666 0.0014
R10040 VSS.n1689 VSS.n1688 0.0014
R10041 VSS.n1659 VSS.n1658 0.0014
R10042 VSS.n1677 VSS.n1675 0.0014
R10043 VSS.n1727 VSS.n1726 0.0014
R10044 VSS.n1725 VSS.n1723 0.0014
R10045 VSS.n1561 VSS.n1560 0.0014
R10046 VSS.n1541 VSS.n1539 0.0014
R10047 VSS.n1542 VSS.n1537 0.0014
R10048 VSS.n1544 VSS.n1535 0.0014
R10049 VSS.n2686 VSS.n2250 0.0013805
R10050 VSS.n3429 VSS.n3428 0.00137209
R10051 VSS.n3200 VSS.n3199 0.00136705
R10052 VSS.n3336 VSS.n3321 0.00136705
R10053 VSS.n2904 VSS.n2903 0.00136076
R10054 VSS.n2902 VSS.n2901 0.00136076
R10055 VSS.n2899 VSS.n2898 0.00136076
R10056 VSS.n2894 VSS.n2893 0.00136076
R10057 VSS.n2891 VSS.n2890 0.00136076
R10058 VSS.n2888 VSS.n2887 0.00136076
R10059 VSS.n3765 VSS.n3764 0.00134112
R10060 VSS.n3763 VSS.n3762 0.00134112
R10061 VSS.n3834 VSS.n3833 0.00134112
R10062 VSS.n3743 VSS.n3742 0.00134112
R10063 VSS.n3812 VSS.n3811 0.00134112
R10064 VSS.n3814 VSS.n3813 0.00134112
R10065 VSS.n3825 VSS.n3810 0.00133916
R10066 VSS.n3840 VSS.n3839 0.00133916
R10067 VSS.n2742 VSS.n2168 0.00133736
R10068 VSS.n2740 VSS.n2739 0.00133736
R10069 VSS.n2204 VSS.n2203 0.00133736
R10070 VSS.n1614 VSS.n1613 0.00132949
R10071 VSS.n1616 VSS.n1615 0.00132949
R10072 VSS.n1623 VSS.n1622 0.00132949
R10073 VSS.n1626 VSS.n1625 0.00132949
R10074 VSS.n1628 VSS.n1627 0.00132949
R10075 VSS.n1635 VSS.n1634 0.00132949
R10076 VSS.n1638 VSS.n1637 0.00132949
R10077 VSS.n1585 VSS.n1584 0.00132949
R10078 VSS.n1593 VSS.n1592 0.00132949
R10079 VSS.n1595 VSS.n1594 0.00132949
R10080 VSS.n1603 VSS.n1602 0.00132949
R10081 VSS.n1605 VSS.n1604 0.00132949
R10082 VSS.n2707 VSS.n2225 0.00131761
R10083 VSS.n2706 VSS.n2226 0.00131761
R10084 VSS.n2695 VSS.n2242 0.00131761
R10085 VSS.n3432 VSS.n3431 0.00131395
R10086 VSS.n3172 VSS.n3171 0.00130925
R10087 VSS.n3355 VSS.n3354 0.00130925
R10088 VSS.n2848 VSS.n2044 0.00130268
R10089 VSS.n2556 VSS.n2416 0.00128603
R10090 VSS.n2523 VSS.n2522 0.00128603
R10091 VSS.n3596 VSS.n3595 0.00128488
R10092 VSS.n3598 VSS.n3597 0.00128488
R10093 VSS.n3708 VSS.n3707 0.00128488
R10094 VSS.n3655 VSS.n3654 0.00128488
R10095 VSS.n3660 VSS.n3659 0.00128488
R10096 VSS.n3495 VSS.n3494 0.00128488
R10097 VSS.n3530 VSS.n3493 0.00128488
R10098 VSS.n3025 VSS.n3024 0.00128488
R10099 VSS.n2621 VSS.n2620 0.00128488
R10100 VSS.n5531 VSS.n5480 0.00127586
R10101 VSS.n1680 VSS.n1679 0.00125419
R10102 VSS.n1695 VSS.n1694 0.00125419
R10103 VSS.n1700 VSS.n1699 0.00125419
R10104 VSS.n1702 VSS.n1701 0.00125419
R10105 VSS.n1711 VSS.n1710 0.00125419
R10106 VSS.n1712 VSS.n1711 0.00125419
R10107 VSS.n1714 VSS.n1713 0.00125419
R10108 VSS.n1716 VSS.n1715 0.00125419
R10109 VSS.n1718 VSS.n1717 0.00125419
R10110 VSS.n3904 VSS.n3903 0.00125419
R10111 VSS.n3908 VSS.n1687 0.00125419
R10112 VSS.n3702 VSS.n3688 0.00125362
R10113 VSS.n2671 VSS.n2276 0.00125251
R10114 VSS.n3134 VSS.n3133 0.00125145
R10115 VSS.n3356 VSS.n3355 0.00125145
R10116 VSS.n3339 VSS.n3336 0.00125145
R10117 VSS.n3320 VSS.n3319 0.00125145
R10118 VSS.n2849 VSS.n2848 0.00123579
R10119 VSS.n3018 VSS.n3017 0.00119767
R10120 VSS.n3711 VSS.n3710 0.00119565
R10121 VSS.n3357 VSS.n3356 0.00119364
R10122 VSS.n3354 VSS.n3339 0.00119364
R10123 VSS.n3321 VSS.n3320 0.00119364
R10124 VSS.n2837 VSS.n2836 0.0011689
R10125 VSS.n2519 VSS.n2451 0.00115502
R10126 VSS.n2521 VSS.n2520 0.00115502
R10127 VSS.n3591 VSS.n3590 0.00115407
R10128 VSS.n1741 VSS.n1740 0.00115407
R10129 VSS.n3675 VSS.n3674 0.00115407
R10130 VSS.n3497 VSS.n3496 0.00115407
R10131 VSS.n3520 VSS.n3519 0.00115407
R10132 VSS.n3508 VSS.n3507 0.00115407
R10133 VSS.n3490 VSS.n3489 0.00115407
R10134 VSS.n3479 VSS.n3478 0.00115407
R10135 VSS.n3462 VSS.n3461 0.00115407
R10136 VSS.n3311 VSS.n3310 0.00115407
R10137 VSS.n3224 VSS.n3222 0.00115407
R10138 VSS.n3181 VSS.n3180 0.00115407
R10139 VSS.n2621 VSS.n2361 0.00115407
R10140 VSS.n2623 VSS.n2622 0.00115407
R10141 VSS.n2369 VSS.n2352 0.00115407
R10142 VSS.n3879 VSS.n3878 0.00115116
R10143 VSS.n3883 VSS.n3882 0.00115116
R10144 VSS.n3851 VSS.n3850 0.00114516
R10145 VSS.n3857 VSS.n3856 0.00114516
R10146 VSS.n3860 VSS.n3859 0.00114516
R10147 VSS.n3866 VSS.n3865 0.00114516
R10148 VSS.n3028 VSS.n3018 0.00113953
R10149 VSS.n3422 VSS.n3421 0.00113953
R10150 VSS.n3418 VSS.n3417 0.00113953
R10151 VSS.n3726 VSS.n3725 0.00113768
R10152 VSS.n3187 VSS.n3174 0.00113584
R10153 VSS.n3781 VSS.n3780 0.00113084
R10154 VSS.n3757 VSS.n3756 0.00113084
R10155 VSS.n3756 VSS.n3755 0.00113084
R10156 VSS.n3755 VSS.n3754 0.00113084
R10157 VSS.n3829 VSS.n3828 0.00113084
R10158 VSS.n1501 VSS.n1500 0.00112937
R10159 VSS.n847 VSS.n846 0.00112937
R10160 VSS.n2457 VSS.n2447 0.00112857
R10161 VSS.n1612 VSS.n1611 0.00112212
R10162 VSS.n1615 VSS.n1614 0.00112212
R10163 VSS.n1622 VSS.n1621 0.00112212
R10164 VSS.n1624 VSS.n1623 0.00112212
R10165 VSS.n1627 VSS.n1626 0.00112212
R10166 VSS.n1634 VSS.n1633 0.00112212
R10167 VSS.n1636 VSS.n1635 0.00112212
R10168 VSS.n1594 VSS.n1593 0.00112212
R10169 VSS.n1604 VSS.n1603 0.00112212
R10170 VSS.n1851 VSS.n1850 0.00112069
R10171 VSS.n1848 VSS.n1847 0.00112069
R10172 VSS.n1845 VSS.n1844 0.00112069
R10173 VSS.n1922 VSS.n1920 0.00112069
R10174 VSS.n2900 VSS.n2899 0.00110759
R10175 VSS.n2801 VSS.n2800 0.00110201
R10176 VSS.n2827 VSS.n2069 0.00110201
R10177 VSS.n2799 VSS.n2080 0.00110201
R10178 VSS.n2815 VSS.n2082 0.00110201
R10179 VSS.n2818 VSS.n2079 0.00110201
R10180 VSS.n2819 VSS.n2074 0.00110201
R10181 VSS.n2145 VSS.n2126 0.00110201
R10182 VSS.n2291 VSS.n2286 0.00110201
R10183 VSS.n2314 VSS.n2310 0.00110201
R10184 VSS.n2647 VSS.n2326 0.0010814
R10185 VSS.n2359 VSS.n2358 0.0010814
R10186 VSS.n3016 VSS.n3015 0.0010814
R10187 VSS.n3420 VSS.n3419 0.0010814
R10188 VSS.n2750 VSS.n2161 0.00107971
R10189 VSS.n3736 VSS.n3735 0.00107971
R10190 VSS.n3189 VSS.n3188 0.00107803
R10191 VSS.n2525 VSS.n2446 0.00107143
R10192 VSS.n3740 VSS.n3739 0.00105944
R10193 VSS.n3772 VSS.n3771 0.00105944
R10194 VSS.n3887 VSS.n3886 0.00105814
R10195 VSS.n3891 VSS.n3890 0.00105814
R10196 VSS.n2901 VSS.n2900 0.00105696
R10197 VSS.n3854 VSS.n3853 0.00105299
R10198 VSS.n3863 VSS.n3862 0.00105299
R10199 VSS.n2529 VSS.n2440 0.00102402
R10200 VSS.n2505 VSS.n2453 0.00102402
R10201 VSS.n2483 VSS.n2474 0.00102402
R10202 VSS.n2493 VSS.n2489 0.00102402
R10203 VSS.n2528 VSS.n2527 0.00102402
R10204 VSS.n2502 VSS.n2475 0.00102402
R10205 VSS.n2419 VSS.n2411 0.00102402
R10206 VSS.n2501 VSS.n2477 0.00102402
R10207 VSS.n3582 VSS.n3581 0.00102326
R10208 VSS.n3580 VSS.n3579 0.00102326
R10209 VSS.n3612 VSS.n3611 0.00102326
R10210 VSS.n3614 VSS.n3613 0.00102326
R10211 VSS.n3616 VSS.n3615 0.00102326
R10212 VSS.n3733 VSS.n3732 0.00102326
R10213 VSS.n3679 VSS.n3678 0.00102326
R10214 VSS.n3521 VSS.n3520 0.00102326
R10215 VSS.n3511 VSS.n3510 0.00102326
R10216 VSS.n3464 VSS.n3463 0.00102326
R10217 VSS.n3288 VSS.n3282 0.00102326
R10218 VSS.n3226 VSS.n3225 0.00102326
R10219 VSS.n3084 VSS.n3083 0.00102326
R10220 VSS.n1790 VSS.n1789 0.00102326
R10221 VSS.n3095 VSS.n3094 0.00102326
R10222 VSS.n3184 VSS.n3183 0.00102326
R10223 VSS.n2946 VSS.n2945 0.00102326
R10224 VSS.n2952 VSS.n2950 0.00102326
R10225 VSS.n2955 VSS.n2954 0.00102326
R10226 VSS.n2574 VSS.n2568 0.00102326
R10227 VSS.n2360 VSS.n2348 0.00102326
R10228 VSS.n2605 VSS.n2604 0.00102326
R10229 VSS.n2577 VSS.n2575 0.00102326
R10230 VSS.n2592 VSS.n2403 0.00102326
R10231 VSS.n2624 VSS.n2350 0.00102326
R10232 VSS.n2576 VSS.n2395 0.00102326
R10233 VSS.n2645 VSS.n2327 0.00102326
R10234 VSS.n2615 VSS.n2366 0.00102326
R10235 VSS.n2600 VSS.n2394 0.00102326
R10236 VSS.n3669 VSS.n3668 0.00102174
R10237 VSS.n3666 VSS.n3663 0.00102174
R10238 VSS.n3652 VSS.n3651 0.00102174
R10239 VSS.n2898 VSS.n2897 0.00100633
R10240 VSS.n2687 VSS.n2686 0.00100314
R10241 VSS.n1670 VSS.n1669 0.00100279
R10242 VSS.n1707 VSS.n1706 0.00100279
R10243 VSS.n3902 VSS.n3898 0.00100279
R10244 VSS.n3769 VSS.n3753 0.0009662
R10245 VSS.n1878 VSS.n1877 0.000965517
R10246 VSS.n1876 VSS.n1875 0.000965517
R10247 VSS.n1972 VSS.n1971 0.000965517
R10248 VSS.n1970 VSS.n1969 0.000965517
R10249 VSS.n1962 VSS.n1961 0.000965517
R10250 VSS.n1960 VSS.n1959 0.000965517
R10251 VSS.n1885 VSS.n1884 0.000965517
R10252 VSS.n1883 VSS.n1882 0.000965517
R10253 VSS.n1881 VSS.n1880 0.000965517
R10254 VSS.n1943 VSS.n1942 0.000965517
R10255 VSS.n1942 VSS.n1941 0.000965517
R10256 VSS.n1940 VSS.n1939 0.000965517
R10257 VSS.n1894 VSS.n1893 0.000965517
R10258 VSS.n1892 VSS.n1891 0.000965517
R10259 VSS.n1890 VSS.n1889 0.000965517
R10260 VSS.n1888 VSS.n1887 0.000965517
R10261 VSS.n1904 VSS.n1903 0.000965517
R10262 VSS.n1902 VSS.n1901 0.000965517
R10263 VSS.n1900 VSS.n1899 0.000965517
R10264 VSS.n1898 VSS.n1897 0.000965517
R10265 VSS.n1978 VSS.n1977 0.000965517
R10266 VSS.n1976 VSS.n1975 0.000965517
R10267 VSS.n1968 VSS.n1967 0.000965517
R10268 VSS.n1966 VSS.n1965 0.000965517
R10269 VSS.n1958 VSS.n1957 0.000965517
R10270 VSS.n1956 VSS.n1955 0.000965517
R10271 VSS.n1953 VSS.n1952 0.000965517
R10272 VSS.n1951 VSS.n1950 0.000965517
R10273 VSS.n1949 VSS.n1948 0.000965517
R10274 VSS.n1938 VSS.n1937 0.000965517
R10275 VSS.n1936 VSS.n1935 0.000965517
R10276 VSS.n1934 VSS.n1933 0.000965517
R10277 VSS.n1931 VSS.n1930 0.000965517
R10278 VSS.n1929 VSS.n1928 0.000965517
R10279 VSS.n1927 VSS.n1926 0.000965517
R10280 VSS.n1925 VSS.n1924 0.000965517
R10281 VSS.n1919 VSS.n1918 0.000965517
R10282 VSS.n1917 VSS.n1916 0.000965517
R10283 VSS.n1915 VSS.n1914 0.000965517
R10284 VSS.n1913 VSS.n1912 0.000965517
R10285 VSS.n3703 VSS.n3702 0.000963768
R10286 VSS.n3118 VSS.n3117 0.000962428
R10287 VSS.n2877 VSS.n2876 0.000951505
R10288 VSS.n2001 VSS.n1997 0.000951505
R10289 VSS.n2868 VSS.n2004 0.000951505
R10290 VSS.n2867 VSS.n2005 0.000951505
R10291 VSS.n2014 VSS.n2012 0.000951505
R10292 VSS.n2859 VSS.n2858 0.000951505
R10293 VSS.n2036 VSS.n2031 0.000951505
R10294 VSS.n2040 VSS.n2039 0.000951505
R10295 VSS.n2037 VSS.n2025 0.000951505
R10296 VSS.n2845 VSS.n2844 0.000951505
R10297 VSS.n2844 VSS.n2046 0.000951505
R10298 VSS.n2841 VSS.n2840 0.000951505
R10299 VSS.n2067 VSS.n2065 0.000951505
R10300 VSS.n2830 VSS.n2829 0.000951505
R10301 VSS.n2826 VSS.n2066 0.000951505
R10302 VSS.n2825 VSS.n2070 0.000951505
R10303 VSS.n2817 VSS.n2081 0.000951505
R10304 VSS.n2814 VSS.n2813 0.000951505
R10305 VSS.n2088 VSS.n2083 0.000951505
R10306 VSS.n2805 VSS.n2804 0.000951505
R10307 VSS.n2875 VSS.n2874 0.000951505
R10308 VSS.n2000 VSS.n1998 0.000951505
R10309 VSS.n2869 VSS.n2003 0.000951505
R10310 VSS.n2866 VSS.n2006 0.000951505
R10311 VSS.n2862 VSS.n2008 0.000951505
R10312 VSS.n2861 VSS.n2860 0.000951505
R10313 VSS.n2035 VSS.n2034 0.000951505
R10314 VSS.n2041 VSS.n2030 0.000951505
R10315 VSS.n2042 VSS.n2027 0.000951505
R10316 VSS.n2847 VSS.n2846 0.000951505
R10317 VSS.n2049 VSS.n2045 0.000951505
R10318 VSS.n2839 VSS.n2838 0.000951505
R10319 VSS.n2833 VSS.n2063 0.000951505
R10320 VSS.n2832 VSS.n2831 0.000951505
R10321 VSS.n2071 VSS.n2064 0.000951505
R10322 VSS.n2824 VSS.n2072 0.000951505
R10323 VSS.n2084 VSS.n2078 0.000951505
R10324 VSS.n2812 VSS.n2811 0.000951505
R10325 VSS.n2808 VSS.n2085 0.000951505
R10326 VSS.n2807 VSS.n2806 0.000951505
R10327 VSS.n2787 VSS.n2786 0.000951505
R10328 VSS.n2101 VSS.n2096 0.000951505
R10329 VSS.n2778 VSS.n2103 0.000951505
R10330 VSS.n2775 VSS.n2105 0.000951505
R10331 VSS.n2133 VSS.n2109 0.000951505
R10332 VSS.n2135 VSS.n2134 0.000951505
R10333 VSS.n2766 VSS.n2117 0.000951505
R10334 VSS.n2765 VSS.n2118 0.000951505
R10335 VSS.n2125 VSS.n2124 0.000951505
R10336 VSS.n2755 VSS.n2128 0.000951505
R10337 VSS.n2752 VSS.n2144 0.000951505
R10338 VSS.n2746 VSS.n2164 0.000951505
R10339 VSS.n2745 VSS.n2165 0.000951505
R10340 VSS.n2735 VSS.n2174 0.000951505
R10341 VSS.n2730 VSS.n2194 0.000951505
R10342 VSS.n2785 VSS.n2784 0.000951505
R10343 VSS.n2099 VSS.n2097 0.000951505
R10344 VSS.n2777 VSS.n2100 0.000951505
R10345 VSS.n2776 VSS.n2104 0.000951505
R10346 VSS.n2113 VSS.n2110 0.000951505
R10347 VSS.n2769 VSS.n2114 0.000951505
R10348 VSS.n2767 VSS.n2116 0.000951505
R10349 VSS.n2764 VSS.n2119 0.000951505
R10350 VSS.n2763 VSS.n2120 0.000951505
R10351 VSS.n2760 VSS.n2120 0.000951505
R10352 VSS.n2759 VSS.n2758 0.000951505
R10353 VSS.n2146 VSS.n2145 0.000951505
R10354 VSS.n2751 VSS.n2147 0.000951505
R10355 VSS.n2748 VSS.n2147 0.000951505
R10356 VSS.n2747 VSS.n2163 0.000951505
R10357 VSS.n2744 VSS.n2166 0.000951505
R10358 VSS.n2736 VSS.n2173 0.000951505
R10359 VSS.n2207 VSS.n2196 0.000951505
R10360 VSS.n2720 VSS.n2719 0.000951505
R10361 VSS.n2218 VSS.n2214 0.000951505
R10362 VSS.n2711 VSS.n2221 0.000951505
R10363 VSS.n2710 VSS.n2222 0.000951505
R10364 VSS.n2229 VSS.n2228 0.000951505
R10365 VSS.n2702 VSS.n2236 0.000951505
R10366 VSS.n2699 VSS.n2698 0.000951505
R10367 VSS.n2246 VSS.n2238 0.000951505
R10368 VSS.n2690 VSS.n2248 0.000951505
R10369 VSS.n2299 VSS.n2298 0.000951505
R10370 VSS.n2678 VSS.n2269 0.000951505
R10371 VSS.n2677 VSS.n2270 0.000951505
R10372 VSS.n2304 VSS.n2303 0.000951505
R10373 VSS.n2669 VSS.n2278 0.000951505
R10374 VSS.n2666 VSS.n2280 0.000951505
R10375 VSS.n2665 VSS.n2281 0.000951505
R10376 VSS.n2718 VSS.n2717 0.000951505
R10377 VSS.n2217 VSS.n2215 0.000951505
R10378 VSS.n2712 VSS.n2220 0.000951505
R10379 VSS.n2709 VSS.n2223 0.000951505
R10380 VSS.n2708 VSS.n2224 0.000951505
R10381 VSS.n2240 VSS.n2239 0.000951505
R10382 VSS.n2697 VSS.n2696 0.000951505
R10383 VSS.n2244 VSS.n2241 0.000951505
R10384 VSS.n2689 VSS.n2245 0.000951505
R10385 VSS.n2688 VSS.n2249 0.000951505
R10386 VSS.n2685 VSS.n2251 0.000951505
R10387 VSS.n2680 VSS.n2254 0.000951505
R10388 VSS.n2679 VSS.n2268 0.000951505
R10389 VSS.n2676 VSS.n2271 0.000951505
R10390 VSS.n2675 VSS.n2272 0.000951505
R10391 VSS.n2668 VSS.n2276 0.000951505
R10392 VSS.n2667 VSS.n2279 0.000951505
R10393 VSS.n2314 VSS.n2313 0.000951505
R10394 VSS.n2160 VSS.n2159 0.000950886
R10395 VSS.n5899 VSS.n5898 0.000940313
R10396 VSS.n1563 VSS.n1562 0.000920561
R10397 VSS.n3784 VSS.n3783 0.000920561
R10398 VSS.n3796 VSS.n3795 0.000920561
R10399 VSS.n3831 VSS.n3830 0.000920561
R10400 VSS.n3764 VSS.n3763 0.000920561
R10401 VSS.n3780 VSS.n3779 0.000920561
R10402 VSS.n3782 VSS.n3781 0.000920561
R10403 VSS.n3801 VSS.n3800 0.000920561
R10404 VSS.n3800 VSS.n3799 0.000920561
R10405 VSS.n3799 VSS.n3798 0.000920561
R10406 VSS.n3835 VSS.n3834 0.000920561
R10407 VSS.n3742 VSS.n3741 0.000920561
R10408 VSS.n3776 VSS.n3775 0.000920561
R10409 VSS.n3777 VSS.n3776 0.000920561
R10410 VSS.n3778 VSS.n3777 0.000920561
R10411 VSS.n3794 VSS.n3793 0.000920561
R10412 VSS.n3792 VSS.n3791 0.000920561
R10413 VSS.n1588 VSS.n1587 0.000914747
R10414 VSS.n1598 VSS.n1597 0.000914747
R10415 VSS.n1034 VSS.n1033 0.000914747
R10416 VSS.n3156 VSS.n3155 0.000904624
R10417 VSS.n2446 VSS.n2434 0.0009
R10418 VSS.n2558 VSS.n2415 0.000893013
R10419 VSS.n2557 VSS.n2556 0.000893013
R10420 VSS.n2427 VSS.n2424 0.000893013
R10421 VSS.n2547 VSS.n2546 0.000893013
R10422 VSS.n2542 VSS.n2541 0.000893013
R10423 VSS.n2437 VSS.n2431 0.000893013
R10424 VSS.n2533 VSS.n2532 0.000893013
R10425 VSS.n2528 VSS.n2441 0.000893013
R10426 VSS.n2449 VSS.n2442 0.000893013
R10427 VSS.n2520 VSS.n2452 0.000893013
R10428 VSS.n2517 VSS.n2516 0.000893013
R10429 VSS.n2472 VSS.n2454 0.000893013
R10430 VSS.n2507 VSS.n2506 0.000893013
R10431 VSS.n2503 VSS.n2473 0.000893013
R10432 VSS.n2495 VSS.n2481 0.000893013
R10433 VSS.n2494 VSS.n2482 0.000893013
R10434 VSS.n2419 VSS.n2417 0.000893013
R10435 VSS.n2555 VSS.n2554 0.000893013
R10436 VSS.n2554 VSS.n2418 0.000893013
R10437 VSS.n2550 VSS.n2422 0.000893013
R10438 VSS.n2549 VSS.n2548 0.000893013
R10439 VSS.n2540 VSS.n2539 0.000893013
R10440 VSS.n2435 VSS.n2432 0.000893013
R10441 VSS.n2535 VSS.n2534 0.000893013
R10442 VSS.n2445 VSS.n2443 0.000893013
R10443 VSS.n2523 VSS.n2444 0.000893013
R10444 VSS.n2455 VSS.n2448 0.000893013
R10445 VSS.n2515 VSS.n2514 0.000893013
R10446 VSS.n2470 VSS.n2456 0.000893013
R10447 VSS.n2509 VSS.n2508 0.000893013
R10448 VSS.n2476 VSS.n2471 0.000893013
R10449 VSS.n2496 VSS.n2480 0.000893013
R10450 VSS.n3732 VSS.n3731 0.000892442
R10451 VSS.n1740 VSS.n1739 0.000892442
R10452 VSS.n1738 VSS.n1737 0.000892442
R10453 VSS.n1736 VSS.n1735 0.000892442
R10454 VSS.n3716 VSS.n3715 0.000892442
R10455 VSS.n3715 VSS.n3714 0.000892442
R10456 VSS.n3707 VSS.n3706 0.000892442
R10457 VSS.n3694 VSS.n3693 0.000892442
R10458 VSS.n3692 VSS.n3691 0.000892442
R10459 VSS.n3690 VSS.n3689 0.000892442
R10460 VSS.n3678 VSS.n3677 0.000892442
R10461 VSS.n3656 VSS.n3655 0.000892442
R10462 VSS.n3654 VSS.n3653 0.000892442
R10463 VSS.n3643 VSS.n3642 0.000892442
R10464 VSS.n3645 VSS.n3644 0.000892442
R10465 VSS.n3630 VSS.n3629 0.000892442
R10466 VSS.n3628 VSS.n3627 0.000892442
R10467 VSS.n3578 VSS.n3577 0.000892442
R10468 VSS.n3729 VSS.n3728 0.000892442
R10469 VSS.n1734 VSS.n1733 0.000892442
R10470 VSS.n1732 VSS.n1731 0.000892442
R10471 VSS.n1730 VSS.n1729 0.000892442
R10472 VSS.n3720 VSS.n3719 0.000892442
R10473 VSS.n3719 VSS.n3718 0.000892442
R10474 VSS.n3705 VSS.n3704 0.000892442
R10475 VSS.n3700 VSS.n3699 0.000892442
R10476 VSS.n3698 VSS.n3697 0.000892442
R10477 VSS.n3676 VSS.n3675 0.000892442
R10478 VSS.n3661 VSS.n3660 0.000892442
R10479 VSS.n3659 VSS.n3658 0.000892442
R10480 VSS.n3639 VSS.n3638 0.000892442
R10481 VSS.n3641 VSS.n3640 0.000892442
R10482 VSS.n3635 VSS.n3634 0.000892442
R10483 VSS.n3633 VSS.n3632 0.000892442
R10484 VSS.n3576 VSS.n3575 0.000892442
R10485 VSS.n3518 VSS.n3517 0.000892442
R10486 VSS.n3450 VSS.n3449 0.000892442
R10487 VSS.n3451 VSS.n3450 0.000892442
R10488 VSS.n3453 VSS.n3452 0.000892442
R10489 VSS.n3456 VSS.n3455 0.000892442
R10490 VSS.n3458 VSS.n3457 0.000892442
R10491 VSS.n3493 VSS.n3492 0.000892442
R10492 VSS.n3491 VSS.n3490 0.000892442
R10493 VSS.n3488 VSS.n3487 0.000892442
R10494 VSS.n3486 VSS.n3485 0.000892442
R10495 VSS.n3484 VSS.n3483 0.000892442
R10496 VSS.n3480 VSS.n3479 0.000892442
R10497 VSS.n3478 VSS.n3477 0.000892442
R10498 VSS.n3476 VSS.n3475 0.000892442
R10499 VSS.n3474 VSS.n3473 0.000892442
R10500 VSS.n3472 VSS.n3471 0.000892442
R10501 VSS.n3469 VSS.n3468 0.000892442
R10502 VSS.n3467 VSS.n3466 0.000892442
R10503 VSS.n3465 VSS.n3464 0.000892442
R10504 VSS.n3461 VSS.n3460 0.000892442
R10505 VSS.n3440 VSS.n3439 0.000892442
R10506 VSS.n3445 VSS.n3444 0.000892442
R10507 VSS.n3447 VSS.n3446 0.000892442
R10508 VSS.n3566 VSS.n3565 0.000892442
R10509 VSS.n3565 VSS.n3564 0.000892442
R10510 VSS.n3563 VSS.n3562 0.000892442
R10511 VSS.n3560 VSS.n3559 0.000892442
R10512 VSS.n3558 VSS.n3557 0.000892442
R10513 VSS.n3556 VSS.n3555 0.000892442
R10514 VSS.n3550 VSS.n3549 0.000892442
R10515 VSS.n3548 VSS.n3547 0.000892442
R10516 VSS.n3546 VSS.n3545 0.000892442
R10517 VSS.n3544 VSS.n3543 0.000892442
R10518 VSS.n3541 VSS.n3540 0.000892442
R10519 VSS.n3539 VSS.n3538 0.000892442
R10520 VSS.n3537 VSS.n3536 0.000892442
R10521 VSS.n3533 VSS.n3532 0.000892442
R10522 VSS.n3411 VSS.n3410 0.000892442
R10523 VSS.n3409 VSS.n3408 0.000892442
R10524 VSS.n1768 VSS.n1767 0.000892442
R10525 VSS.n3347 VSS.n3346 0.000892442
R10526 VSS.n3349 VSS.n3348 0.000892442
R10527 VSS.n3351 VSS.n3350 0.000892442
R10528 VSS.n3327 VSS.n3326 0.000892442
R10529 VSS.n3325 VSS.n3324 0.000892442
R10530 VSS.n3323 VSS.n3322 0.000892442
R10531 VSS.n3306 VSS.n3305 0.000892442
R10532 VSS.n3308 VSS.n3307 0.000892442
R10533 VSS.n3310 VSS.n3309 0.000892442
R10534 VSS.n3282 VSS.n3281 0.000892442
R10535 VSS.n3287 VSS.n3286 0.000892442
R10536 VSS.n3285 VSS.n3284 0.000892442
R10537 VSS.n3272 VSS.n3271 0.000892442
R10538 VSS.n3270 VSS.n3269 0.000892442
R10539 VSS.n1766 VSS.n1765 0.000892442
R10540 VSS.n3341 VSS.n3340 0.000892442
R10541 VSS.n3343 VSS.n3342 0.000892442
R10542 VSS.n3345 VSS.n3344 0.000892442
R10543 VSS.n3334 VSS.n3333 0.000892442
R10544 VSS.n3332 VSS.n3331 0.000892442
R10545 VSS.n3330 VSS.n3329 0.000892442
R10546 VSS.n3302 VSS.n3301 0.000892442
R10547 VSS.n3304 VSS.n3303 0.000892442
R10548 VSS.n3313 VSS.n3312 0.000892442
R10549 VSS.n3280 VSS.n3279 0.000892442
R10550 VSS.n3293 VSS.n3292 0.000892442
R10551 VSS.n3291 VSS.n3290 0.000892442
R10552 VSS.n3267 VSS.n3266 0.000892442
R10553 VSS.n3265 VSS.n3264 0.000892442
R10554 VSS.n3254 VSS.n3253 0.000892442
R10555 VSS.n3246 VSS.n3245 0.000892442
R10556 VSS.n3237 VSS.n3236 0.000892442
R10557 VSS.n3235 VSS.n3234 0.000892442
R10558 VSS.n3195 VSS.n3194 0.000892442
R10559 VSS.n1787 VSS.n1786 0.000892442
R10560 VSS.n1789 VSS.n1788 0.000892442
R10561 VSS.n3180 VSS.n3179 0.000892442
R10562 VSS.n3178 VSS.n3177 0.000892442
R10563 VSS.n3176 VSS.n3175 0.000892442
R10564 VSS.n3164 VSS.n3163 0.000892442
R10565 VSS.n3162 VSS.n3161 0.000892442
R10566 VSS.n3143 VSS.n3142 0.000892442
R10567 VSS.n3128 VSS.n3127 0.000892442
R10568 VSS.n3126 VSS.n3125 0.000892442
R10569 VSS.n3109 VSS.n3108 0.000892442
R10570 VSS.n3107 VSS.n3106 0.000892442
R10571 VSS.n3096 VSS.n3095 0.000892442
R10572 VSS.n3094 VSS.n3093 0.000892442
R10573 VSS.n3205 VSS.n3204 0.000892442
R10574 VSS.n3203 VSS.n3202 0.000892442
R10575 VSS.n3193 VSS.n3192 0.000892442
R10576 VSS.n1783 VSS.n1782 0.000892442
R10577 VSS.n1785 VSS.n1784 0.000892442
R10578 VSS.n3185 VSS.n3184 0.000892442
R10579 VSS.n3183 VSS.n3182 0.000892442
R10580 VSS.n3160 VSS.n3159 0.000892442
R10581 VSS.n3169 VSS.n3168 0.000892442
R10582 VSS.n3167 VSS.n3166 0.000892442
R10583 VSS.n3149 VSS.n3148 0.000892442
R10584 VSS.n3139 VSS.n3138 0.000892442
R10585 VSS.n3137 VSS.n3136 0.000892442
R10586 VSS.n3123 VSS.n3122 0.000892442
R10587 VSS.n3121 VSS.n3120 0.000892442
R10588 VSS.n3101 VSS.n3100 0.000892442
R10589 VSS.n3099 VSS.n3098 0.000892442
R10590 VSS.n3058 VSS.n3057 0.000892442
R10591 VSS.n3062 VSS.n3061 0.000892442
R10592 VSS.n3060 VSS.n3059 0.000892442
R10593 VSS.n1823 VSS.n1822 0.000892442
R10594 VSS.n1821 VSS.n1820 0.000892442
R10595 VSS.n3043 VSS.n3042 0.000892442
R10596 VSS.n3033 VSS.n3032 0.000892442
R10597 VSS.n3035 VSS.n3034 0.000892442
R10598 VSS.n3021 VSS.n3020 0.000892442
R10599 VSS.n3020 VSS.n3019 0.000892442
R10600 VSS.n3008 VSS.n3007 0.000892442
R10601 VSS.n3010 VSS.n3009 0.000892442
R10602 VSS.n2992 VSS.n2991 0.000892442
R10603 VSS.n2994 VSS.n2993 0.000892442
R10604 VSS.n2996 VSS.n2995 0.000892442
R10605 VSS.n2972 VSS.n2971 0.000892442
R10606 VSS.n2970 VSS.n2969 0.000892442
R10607 VSS.n2968 VSS.n2967 0.000892442
R10608 VSS.n2920 VSS.n2919 0.000892442
R10609 VSS.n3056 VSS.n3055 0.000892442
R10610 VSS.n3067 VSS.n3066 0.000892442
R10611 VSS.n3065 VSS.n3064 0.000892442
R10612 VSS.n1819 VSS.n1818 0.000892442
R10613 VSS.n1817 VSS.n1816 0.000892442
R10614 VSS.n3047 VSS.n3046 0.000892442
R10615 VSS.n3031 VSS.n3030 0.000892442
R10616 VSS.n3026 VSS.n3025 0.000892442
R10617 VSS.n3024 VSS.n3023 0.000892442
R10618 VSS.n3006 VSS.n3005 0.000892442
R10619 VSS.n3013 VSS.n3012 0.000892442
R10620 VSS.n2986 VSS.n2985 0.000892442
R10621 VSS.n2988 VSS.n2987 0.000892442
R10622 VSS.n2990 VSS.n2989 0.000892442
R10623 VSS.n2979 VSS.n2978 0.000892442
R10624 VSS.n2977 VSS.n2976 0.000892442
R10625 VSS.n2975 VSS.n2974 0.000892442
R10626 VSS.n2918 VSS.n2917 0.000892442
R10627 VSS.n2654 VSS.n2653 0.000892442
R10628 VSS.n2328 VSS.n2322 0.000892442
R10629 VSS.n2343 VSS.n2335 0.000892442
R10630 VSS.n2344 VSS.n2342 0.000892442
R10631 VSS.n2631 VSS.n2347 0.000892442
R10632 VSS.n2628 VSS.n2349 0.000892442
R10633 VSS.n2627 VSS.n2350 0.000892442
R10634 VSS.n2622 VSS.n2362 0.000892442
R10635 VSS.n2619 VSS.n2362 0.000892442
R10636 VSS.n2618 VSS.n2617 0.000892442
R10637 VSS.n2388 VSS.n2386 0.000892442
R10638 VSS.n2607 VSS.n2606 0.000892442
R10639 VSS.n2603 VSS.n2387 0.000892442
R10640 VSS.n2602 VSS.n2391 0.000892442
R10641 VSS.n2594 VSS.n2401 0.000892442
R10642 VSS.n2593 VSS.n2402 0.000892442
R10643 VSS.n2590 VSS.n2589 0.000892442
R10644 VSS.n2566 VSS.n2405 0.000892442
R10645 VSS.n2652 VSS.n2651 0.000892442
R10646 VSS.n2324 VSS.n2323 0.000892442
R10647 VSS.n2646 VSS.n2645 0.000892442
R10648 VSS.n2336 VSS.n2327 0.000892442
R10649 VSS.n2339 VSS.n2337 0.000892442
R10650 VSS.n2634 VSS.n2340 0.000892442
R10651 VSS.n2354 VSS.n2341 0.000892442
R10652 VSS.n2356 VSS.n2355 0.000892442
R10653 VSS.n2626 VSS.n2351 0.000892442
R10654 VSS.n2369 VSS.n2368 0.000892442
R10655 VSS.n2368 VSS.n2365 0.000892442
R10656 VSS.n2616 VSS.n2615 0.000892442
R10657 VSS.n2610 VSS.n2384 0.000892442
R10658 VSS.n2609 VSS.n2608 0.000892442
R10659 VSS.n2392 VSS.n2385 0.000892442
R10660 VSS.n2601 VSS.n2393 0.000892442
R10661 VSS.n2595 VSS.n2400 0.000892442
R10662 VSS.n2407 VSS.n2406 0.000892442
R10663 VSS.n2588 VSS.n2587 0.000892442
R10664 VSS.n2565 VSS.n2408 0.000892442
R10665 VSS.n2762 VSS.n2761 0.000886473
R10666 VSS.n2750 VSS.n2749 0.000886473
R10667 VSS.n2371 VSS.n2370 0.000848837
R10668 VSS.n3713 VSS.n3712 0.000847826
R10669 VSS.n2524 VSS.n2447 0.000842857
R10670 VSS.n2836 VSS.n2835 0.000834448
R10671 VSS.n2159 VSS.n2123 0.000822061
R10672 VSS.n2311 VSS.n2274 0.000814465
R10673 VSS.n2192 VSS.n2177 0.000801003
R10674 VSS.n2185 VSS.n2178 0.000801003
R10675 VSS.n2191 VSS.n2190 0.000801003
R10676 VSS.n2733 VSS.n2732 0.000801003
R10677 VSS.n2757 VSS.n2756 0.000801003
R10678 VSS.n2183 VSS.n2180 0.000801003
R10679 VSS.n2187 VSS.n2186 0.000801003
R10680 VSS.n2172 VSS.n2171 0.000801003
R10681 VSS.n2734 VSS.n2175 0.000801003
R10682 VSS.n2201 VSS.n2200 0.000801003
R10683 VSS.n2758 VSS.n2126 0.000801003
R10684 VSS.n2743 VSS.n2167 0.000801003
R10685 VSS.n2182 VSS.n2181 0.000801003
R10686 VSS.n2738 VSS.n2737 0.000801003
R10687 VSS.n2202 VSS.n2199 0.000801003
R10688 VSS.n2206 VSS.n2205 0.000801003
R10689 VSS.n2289 VSS.n2288 0.000801003
R10690 VSS.n2251 VSS.n2249 0.000801003
R10691 VSS.n2370 VSS.n2367 0.000790698
R10692 VSS.n3147 VSS.n3134 0.000789017
R10693 VSS.n3252 VSS.n3243 0.000789017
R10694 VSS.n3895 VSS.n3894 0.00077907
R10695 VSS.n2076 VSS.n2075 0.000767559
R10696 VSS.n2821 VSS.n2820 0.000767559
R10697 VSS.n2810 VSS.n2809 0.000767559
R10698 VSS.n3682 VSS.n3681 0.000761628
R10699 VSS.n3680 VSS.n3679 0.000761628
R10700 VSS.n3673 VSS.n3672 0.000761628
R10701 VSS.n3454 VSS.n3453 0.000761628
R10702 VSS.n3442 VSS.n3441 0.000761628
R10703 VSS.n3562 VSS.n3561 0.000761628
R10704 VSS.n3553 VSS.n3552 0.000761628
R10705 VSS.n3379 VSS.n3378 0.000761628
R10706 VSS.n3410 VSS.n3409 0.000761628
R10707 VSS.n3257 VSS.n3256 0.000761628
R10708 VSS.n3250 VSS.n3249 0.000761628
R10709 VSS.n3365 VSS.n3364 0.000761628
R10710 VSS.n3314 VSS.n3313 0.000761628
R10711 VSS.n3266 VSS.n3265 0.000761628
R10712 VSS.n3251 VSS.n3246 0.000761628
R10713 VSS.n3216 VSS.n3215 0.000761628
R10714 VSS.n3152 VSS.n3151 0.000761628
R10715 VSS.n3145 VSS.n3144 0.000761628
R10716 VSS.n3108 VSS.n3107 0.000761628
R10717 VSS.n3146 VSS.n3139 0.000761628
R10718 VSS.n3113 VSS.n3112 0.000761628
R10719 VSS.n2642 VSS.n2641 0.000761628
R10720 VSS.n2643 VSS.n2330 0.000761628
R10721 VSS.n2316 VSS.n2315 0.000751572
R10722 VSS.n1657 VSS.n1656 0.000751397
R10723 VSS.n1672 VSS.n1671 0.000751397
R10724 VSS.n1696 VSS.n1695 0.000751397
R10725 VSS.n1698 VSS.n1697 0.000751397
R10726 VSS.n1708 VSS.n1707 0.000751397
R10727 VSS.n1710 VSS.n1709 0.000751397
R10728 VSS.n1717 VSS.n1716 0.000751397
R10729 VSS.n3898 VSS.n3897 0.000751397
R10730 VSS.n3905 VSS.n3902 0.000751397
R10731 VSS.n4118 VSS.n4117 0.00074
R10732 VSS.n2614 VSS.n2613 0.000732558
R10733 VSS.n2396 VSS.n2383 0.000732558
R10734 VSS.n2599 VSS.n2598 0.000732558
R10735 VSS.n2409 VSS.n2398 0.000732558
R10736 VSS.n3001 VSS.n3000 0.000732558
R10737 VSS.n2984 VSS.n2981 0.000732558
R10738 VSS.n2965 VSS.n2964 0.000732558
R10739 VSS.n3650 VSS.n3649 0.000731884
R10740 VSS.n3648 VSS.n3637 0.000731884
R10741 VSS.n3626 VSS.n3625 0.000731884
R10742 VSS.n3174 VSS.n3173 0.000731214
R10743 VSS.n3155 VSS.n3154 0.000731214
R10744 VSS.n3105 VSS.n3104 0.000731214
R10745 VSS.n3361 VSS.n3360 0.000731214
R10746 VSS.n3260 VSS.n3259 0.000731214
R10747 VSS.n2420 VSS.n2410 0.000728571
R10748 VSS.n2511 VSS.n2510 0.000728571
R10749 VSS.n2500 VSS.n2499 0.000728571
R10750 VSS.n5865 VSS.n5864 0.000713777
R10751 VSS.n5867 VSS.n5866 0.000713777
R10752 VSS.n5869 VSS.n5868 0.000713777
R10753 VSS.n3821 VSS.n3820 0.00071028
R10754 VSS.n3745 VSS.n3744 0.00071028
R10755 VSS.n3822 VSS.n3818 0.00071028
R10756 VSS.n3751 VSS.n3750 0.00071028
R10757 VSS.n3768 VSS.n3767 0.00071028
R10758 VSS.n3788 VSS.n3787 0.00071028
R10759 VSS.n3804 VSS.n3803 0.00071028
R10760 VSS.n3793 VSS.n3792 0.00071028
R10761 VSS.n3824 VSS.n3823 0.00071028
R10762 VSS.n3837 VSS.n3836 0.00071028
R10763 VSS.n1610 VSS.n1609 0.000707373
R10764 VSS.n1618 VSS.n1617 0.000707373
R10765 VSS.n1620 VSS.n1619 0.000707373
R10766 VSS.n1630 VSS.n1629 0.000707373
R10767 VSS.n1632 VSS.n1631 0.000707373
R10768 VSS.n1641 VSS.n1639 0.000707373
R10769 VSS.n2893 VSS.n2892 0.000702532
R10770 VSS.n2890 VSS.n2889 0.000702532
R10771 VSS.n2887 VSS.n2886 0.000702532
R10772 VSS.n3774 VSS.n3773 0.00068648
R10773 VSS.n3808 VSS.n3807 0.00068648
R10774 VSS.n3901 VSS.n3899 0.000686047
R10775 VSS.n3567 VSS.n3437 0.000674419
R10776 VSS.n3427 VSS.n3426 0.000674419
R10777 VSS.n2553 VSS.n2552 0.000671429
R10778 VSS.n2513 VSS.n2512 0.000671429
R10779 VSS.n1889 VSS.n1888 0.000655172
R10780 VSS.n1901 VSS.n1900 0.000655172
R10781 VSS.n1926 VSS.n1925 0.000655172
R10782 VSS.n1916 VSS.n1915 0.000655172
R10783 VSS.n2826 VSS.n2825 0.000650502
R10784 VSS.n2813 VSS.n2083 0.000650502
R10785 VSS.n2072 VSS.n2071 0.000650502
R10786 VSS.n2811 VSS.n2085 0.000650502
R10787 VSS.n2754 VSS.n2127 0.000650502
R10788 VSS.n2756 VSS.n2755 0.000650502
R10789 VSS.n2186 VSS.n2183 0.000650502
R10790 VSS.n2200 VSS.n2175 0.000650502
R10791 VSS.n2181 VSS.n2167 0.000650502
R10792 VSS.n2205 VSS.n2202 0.000650502
R10793 VSS.n2288 VSS.n2287 0.000650502
R10794 VSS.n2290 VSS.n2289 0.000650502
R10795 VSS.n2507 VSS.n2472 0.000631004
R10796 VSS.n2495 VSS.n2494 0.000631004
R10797 VSS.n2509 VSS.n2470 0.000631004
R10798 VSS.n2490 VSS.n2480 0.000631004
R10799 VSS.n3605 VSS.n3604 0.000630814
R10800 VSS.n3681 VSS.n3680 0.000630814
R10801 VSS.n3644 VSS.n3643 0.000630814
R10802 VSS.n3629 VSS.n3628 0.000630814
R10803 VSS.n3674 VSS.n3673 0.000630814
R10804 VSS.n3672 VSS.n3671 0.000630814
R10805 VSS.n3640 VSS.n3639 0.000630814
R10806 VSS.n3634 VSS.n3633 0.000630814
R10807 VSS.n3481 VSS.n3480 0.000630814
R10808 VSS.n3443 VSS.n3442 0.000630814
R10809 VSS.n3552 VSS.n3551 0.000630814
R10810 VSS.n3377 VSS.n3376 0.000630814
R10811 VSS.n3257 VSS.n3255 0.000630814
R10812 VSS.n3250 VSS.n3247 0.000630814
R10813 VSS.n3366 VSS.n3365 0.000630814
R10814 VSS.n3364 VSS.n3363 0.000630814
R10815 VSS.n3294 VSS.n3280 0.000630814
R10816 VSS.n3258 VSS.n3254 0.000630814
R10817 VSS.n3214 VSS.n3213 0.000630814
R10818 VSS.n3152 VSS.n3150 0.000630814
R10819 VSS.n3145 VSS.n3140 0.000630814
R10820 VSS.n3153 VSS.n3149 0.000630814
R10821 VSS.n3114 VSS.n3113 0.000630814
R10822 VSS.n3112 VSS.n3111 0.000630814
R10823 VSS.n2995 VSS.n2994 0.000630814
R10824 VSS.n2969 VSS.n2968 0.000630814
R10825 VSS.n2989 VSS.n2988 0.000630814
R10826 VSS.n2976 VSS.n2975 0.000630814
R10827 VSS.n2644 VSS.n2643 0.000630814
R10828 VSS.n2334 VSS.n2330 0.000630814
R10829 VSS.n2606 VSS.n2387 0.000630814
R10830 VSS.n2594 VSS.n2593 0.000630814
R10831 VSS.n2608 VSS.n2385 0.000630814
R10832 VSS.n2406 VSS.n2400 0.000630814
R10833 VSS.n2742 VSS.n2741 0.000628824
R10834 VSS.n2739 VSS.n2170 0.000628824
R10835 VSS.n2204 VSS.n2198 0.000628824
R10836 VSS.n2682 VSS.n2266 0.000625786
R10837 VSS.n3436 VSS.n3435 0.000616279
R10838 VSS.n3430 VSS.n3429 0.000616279
R10839 VSS.n3668 VSS.n3667 0.000615942
R10840 VSS.n3315 VSS.n3300 0.000615607
R10841 VSS.n3262 VSS.n3261 0.000615607
R10842 VSS.n3753 VSS.n3752 0.00059324
R10843 VSS.n3770 VSS.n3769 0.00059324
R10844 VSS.n3790 VSS.n3789 0.00059324
R10845 VSS.n3805 VSS.n3790 0.00059324
R10846 VSS.n3806 VSS.n3805 0.00059324
R10847 VSS.n3826 VSS.n3825 0.00059324
R10848 VSS.n3839 VSS.n3838 0.00059324
R10849 VSS.n3880 VSS.n3879 0.000593023
R10850 VSS.n3882 VSS.n3881 0.000593023
R10851 VSS.n3888 VSS.n3887 0.000593023
R10852 VSS.n3890 VSS.n3889 0.000593023
R10853 VSS.n3901 VSS.n3900 0.000593023
R10854 VSS.n5861 VSS 0.000592784
R10855 VSS.n3848 VSS.n3847 0.000592166
R10856 VSS.n3853 VSS.n3852 0.000592166
R10857 VSS.n3855 VSS.n3854 0.000592166
R10858 VSS.n3862 VSS.n3861 0.000592166
R10859 VSS.n3864 VSS.n3863 0.000592166
R10860 VSS.n3869 VSS.n3868 0.000592166
R10861 VSS.n3003 VSS.n3002 0.00055814
R10862 VSS.n3571 VSS.n3570 0.00055814
R10863 VSS.n3317 VSS.n3316 0.000557804
R10864 VSS.n3296 VSS.n3295 0.000557804
R10865 VSS.n2896 VSS.n2895 0.000550633
R10866 VCTRL2.n124 VCTRL2.n123 10.0043
R10867 VCTRL2.n124 VCTRL2.n61 9.34779
R10868 VCTRL2.n53 VCTRL2.t66 8.213
R10869 VCTRL2.n26 VCTRL2.t30 8.213
R10870 VCTRL2.n112 VCTRL2.t12 8.16955
R10871 VCTRL2.n99 VCTRL2.t36 8.16955
R10872 VCTRL2.n33 VCTRL2.t23 8.16955
R10873 VCTRL2.n18 VCTRL2.t16 8.16955
R10874 VCTRL2.n22 VCTRL2.t24 8.16955
R10875 VCTRL2.n58 VCTRL2.t34 8.16955
R10876 VCTRL2.n88 VCTRL2.t22 8.1261
R10877 VCTRL2.n81 VCTRL2.t26 8.1261
R10878 VCTRL2.n95 VCTRL2.t17 8.1261
R10879 VCTRL2.n117 VCTRL2.t0 8.1261
R10880 VCTRL2.n44 VCTRL2.t11 8.1261
R10881 VCTRL2.n13 VCTRL2.t67 8.1261
R10882 VCTRL2.n75 VCTRL2.t9 8.08264
R10883 VCTRL2.n67 VCTRL2.t72 8.08264
R10884 VCTRL2.n49 VCTRL2.t15 7.51776
R10885 VCTRL2.n24 VCTRL2.t70 7.51776
R10886 VCTRL2.n108 VCTRL2.t13 7.47431
R10887 VCTRL2.n97 VCTRL2.t44 7.47431
R10888 VCTRL2.n56 VCTRL2.t74 7.47431
R10889 VCTRL2.n29 VCTRL2.t60 7.47431
R10890 VCTRL2.n15 VCTRL2.t54 7.47431
R10891 VCTRL2.n51 VCTRL2.t2 7.47431
R10892 VCTRL2.n20 VCTRL2.t61 7.47431
R10893 VCTRL2.n25 VCTRL2.t48 7.47431
R10894 VCTRL2.n85 VCTRL2.t49 7.43086
R10895 VCTRL2.n78 VCTRL2.t59 7.43086
R10896 VCTRL2.n111 VCTRL2.t1 7.43086
R10897 VCTRL2.n92 VCTRL2.t75 7.43086
R10898 VCTRL2.n115 VCTRL2.t19 7.43086
R10899 VCTRL2.n98 VCTRL2.t27 7.43086
R10900 VCTRL2.n30 VCTRL2.t38 7.43086
R10901 VCTRL2.n16 VCTRL2.t32 7.43086
R10902 VCTRL2.n41 VCTRL2.t45 7.43086
R10903 VCTRL2.n5 VCTRL2.t18 7.43086
R10904 VCTRL2.n21 VCTRL2.t39 7.43086
R10905 VCTRL2.n57 VCTRL2.t51 7.43086
R10906 VCTRL2.n87 VCTRL2.t33 7.3874
R10907 VCTRL2.n80 VCTRL2.t40 7.3874
R10908 VCTRL2.n72 VCTRL2.t8 7.3874
R10909 VCTRL2.n65 VCTRL2.t31 7.3874
R10910 VCTRL2.n93 VCTRL2.t57 7.3874
R10911 VCTRL2.n116 VCTRL2.t7 7.3874
R10912 VCTRL2.n42 VCTRL2.t25 7.3874
R10913 VCTRL2.n11 VCTRL2.t3 7.3874
R10914 VCTRL2.n74 VCTRL2.t73 7.34395
R10915 VCTRL2.n66 VCTRL2.t14 7.34395
R10916 VCTRL2.n76 VCTRL2.t62 7.3005
R10917 VCTRL2.n68 VCTRL2.t42 7.3005
R10918 VCTRL2.n96 VCTRL2.t76 7.25705
R10919 VCTRL2.n89 VCTRL2.t79 7.25705
R10920 VCTRL2.n82 VCTRL2.t4 7.25705
R10921 VCTRL2.t9 VCTRL2.n74 7.25705
R10922 VCTRL2.t72 VCTRL2.n66 7.25705
R10923 VCTRL2.n118 VCTRL2.t52 7.25705
R10924 VCTRL2.n45 VCTRL2.t28 7.25705
R10925 VCTRL2.n14 VCTRL2.t6 7.25705
R10926 VCTRL2.n100 VCTRL2.t10 7.2136
R10927 VCTRL2.t22 VCTRL2.n87 7.2136
R10928 VCTRL2.t26 VCTRL2.n80 7.2136
R10929 VCTRL2.t73 VCTRL2.n72 7.2136
R10930 VCTRL2.t14 VCTRL2.n65 7.2136
R10931 VCTRL2.n113 VCTRL2.t69 7.2136
R10932 VCTRL2.t17 VCTRL2.n93 7.2136
R10933 VCTRL2.t0 VCTRL2.n116 7.2136
R10934 VCTRL2.n34 VCTRL2.t41 7.2136
R10935 VCTRL2.n19 VCTRL2.t35 7.2136
R10936 VCTRL2.t11 VCTRL2.n42 7.2136
R10937 VCTRL2.t67 VCTRL2.n11 7.2136
R10938 VCTRL2.n23 VCTRL2.t43 7.2136
R10939 VCTRL2.n59 VCTRL2.t55 7.2136
R10940 VCTRL2.t33 VCTRL2.n85 7.17014
R10941 VCTRL2.t40 VCTRL2.n78 7.17014
R10942 VCTRL2.t12 VCTRL2.n111 7.17014
R10943 VCTRL2.t57 VCTRL2.n92 7.17014
R10944 VCTRL2.t7 VCTRL2.n115 7.17014
R10945 VCTRL2.t36 VCTRL2.n98 7.17014
R10946 VCTRL2.t23 VCTRL2.n30 7.17014
R10947 VCTRL2.t16 VCTRL2.n16 7.17014
R10948 VCTRL2.t25 VCTRL2.n41 7.17014
R10949 VCTRL2.t3 VCTRL2.n5 7.17014
R10950 VCTRL2.n54 VCTRL2.t5 7.17014
R10951 VCTRL2.t24 VCTRL2.n21 7.17014
R10952 VCTRL2.t34 VCTRL2.n57 7.17014
R10953 VCTRL2.n27 VCTRL2.t50 7.17014
R10954 VCTRL2.t1 VCTRL2.n108 7.12669
R10955 VCTRL2.t27 VCTRL2.n97 7.12669
R10956 VCTRL2.t38 VCTRL2.n29 7.12669
R10957 VCTRL2.t32 VCTRL2.n15 7.12669
R10958 VCTRL2.t66 VCTRL2.n51 7.12669
R10959 VCTRL2.t39 VCTRL2.n20 7.12669
R10960 VCTRL2.t51 VCTRL2.n56 7.12669
R10961 VCTRL2.t30 VCTRL2.n25 7.12669
R10962 VCTRL2.t2 VCTRL2.n49 7.08324
R10963 VCTRL2.n54 VCTRL2.t20 7.08324
R10964 VCTRL2.t48 VCTRL2.n24 7.08324
R10965 VCTRL2.n27 VCTRL2.t71 7.08324
R10966 VCTRL2.n113 VCTRL2.t53 7.03979
R10967 VCTRL2.n100 VCTRL2.t78 7.03979
R10968 VCTRL2.n34 VCTRL2.t63 7.03979
R10969 VCTRL2.n19 VCTRL2.t56 7.03979
R10970 VCTRL2.n23 VCTRL2.t64 7.03979
R10971 VCTRL2.n59 VCTRL2.t77 7.03979
R10972 VCTRL2.n96 VCTRL2.t58 6.99633
R10973 VCTRL2.n89 VCTRL2.t65 6.99633
R10974 VCTRL2.n82 VCTRL2.t68 6.99633
R10975 VCTRL2.n118 VCTRL2.t37 6.99633
R10976 VCTRL2.n45 VCTRL2.t47 6.99633
R10977 VCTRL2.n14 VCTRL2.t21 6.99633
R10978 VCTRL2.n76 VCTRL2.t46 6.95288
R10979 VCTRL2.n68 VCTRL2.t29 6.95288
R10980 VCTRL2.t46 VCTRL2.n75 6.51836
R10981 VCTRL2.t29 VCTRL2.n67 6.51836
R10982 VCTRL2.t58 VCTRL2.n95 6.4749
R10983 VCTRL2.t65 VCTRL2.n88 6.4749
R10984 VCTRL2.t68 VCTRL2.n81 6.4749
R10985 VCTRL2.t37 VCTRL2.n117 6.4749
R10986 VCTRL2.t47 VCTRL2.n44 6.4749
R10987 VCTRL2.t21 VCTRL2.n13 6.4749
R10988 VCTRL2.t53 VCTRL2.n112 6.43145
R10989 VCTRL2.t78 VCTRL2.n99 6.43145
R10990 VCTRL2.t63 VCTRL2.n33 6.43145
R10991 VCTRL2.t56 VCTRL2.n18 6.43145
R10992 VCTRL2.t64 VCTRL2.n22 6.43145
R10993 VCTRL2.t77 VCTRL2.n58 6.43145
R10994 VCTRL2.t20 VCTRL2.n53 6.388
R10995 VCTRL2.t71 VCTRL2.n26 6.388
R10996 VCTRL2.n28 VCTRL2.n27 4.03166
R10997 VCTRL2.n101 VCTRL2.n100 4.0306
R10998 VCTRL2.n119 VCTRL2.n118 3.63007
R10999 VCTRL2.n60 VCTRL2.n59 3.62933
R11000 VCTRL2.n11 VCTRL2.n10 3.62499
R11001 VCTRL2.n102 VCTRL2.n89 3.62466
R11002 VCTRL2.n88 VCTRL2.n83 3.62466
R11003 VCTRL2.n108 VCTRL2.n107 3.62466
R11004 VCTRL2.n5 VCTRL2.n4 3.62466
R11005 VCTRL2.n41 VCTRL2.n40 3.62466
R11006 VCTRL2.n28 VCTRL2.n23 3.62466
R11007 VCTRL2.n36 VCTRL2.n19 3.62466
R11008 VCTRL2.n47 VCTRL2.n14 3.62466
R11009 VCTRL2.n85 VCTRL2.n84 3.62466
R11010 VCTRL2.n87 VCTRL2.n86 3.62466
R11011 VCTRL2.n112 VCTRL2.n106 3.62466
R11012 VCTRL2.n114 VCTRL2.n113 3.62466
R11013 VCTRL2.n111 VCTRL2.n110 3.62466
R11014 VCTRL2.n18 VCTRL2.n17 3.62466
R11015 VCTRL2.n44 VCTRL2.n43 3.62466
R11016 VCTRL2.n46 VCTRL2.n45 3.62466
R11017 VCTRL2.n13 VCTRL2.n12 3.62466
R11018 VCTRL2.n101 VCTRL2.n96 3.62462
R11019 VCTRL2.n103 VCTRL2.n82 3.62462
R11020 VCTRL2.n78 VCTRL2.n77 3.62462
R11021 VCTRL2.n80 VCTRL2.n79 3.62462
R11022 VCTRL2.n75 VCTRL2.n70 3.62462
R11023 VCTRL2.n104 VCTRL2.n76 3.62462
R11024 VCTRL2.n72 VCTRL2.n71 3.62462
R11025 VCTRL2.n74 VCTRL2.n73 3.62462
R11026 VCTRL2.n67 VCTRL2.n63 3.62462
R11027 VCTRL2.n105 VCTRL2.n68 3.62462
R11028 VCTRL2.n65 VCTRL2.n64 3.62462
R11029 VCTRL2.n93 VCTRL2.n90 3.62462
R11030 VCTRL2.n92 VCTRL2.n91 3.62462
R11031 VCTRL2.n95 VCTRL2.n94 3.62462
R11032 VCTRL2.n33 VCTRL2.n32 3.62462
R11033 VCTRL2.n35 VCTRL2.n34 3.62462
R11034 VCTRL2.n49 VCTRL2.n48 3.62462
R11035 VCTRL2.n53 VCTRL2.n52 3.62462
R11036 VCTRL2.n55 VCTRL2.n54 3.62462
R11037 VCTRL2.n51 VCTRL2.n50 3.62462
R11038 VCTRL2.n122 VCTRL2.n121 2.2505
R11039 VCTRL2.n3 VCTRL2.n2 2.2505
R11040 VCTRL2.n125 VCTRL2.n124 1.5049
R11041 VCTRL2 VCTRL2.n0 1.16594
R11042 VCTRL2 VCTRL2.n62 1.16341
R11043 VCTRL2.n122 VCTRL2.n119 1.05045
R11044 VCTRL2.n61 VCTRL2.n60 0.984409
R11045 VCTRL2.n120 VCTRL2 0.936261
R11046 VCTRL2.n1 VCTRL2 0.936261
R11047 VCTRL2.n125 VCTRL2 0.61117
R11048 VCTRL2.n119 VCTRL2.n114 0.442081
R11049 VCTRL2.n60 VCTRL2.n55 0.441056
R11050 VCTRL2.n8 VCTRL2.n7 0.404715
R11051 VCTRL2.n36 VCTRL2.n35 0.404715
R11052 VCTRL2.n103 VCTRL2.n102 0.404539
R11053 VCTRL2.n39 VCTRL2.n38 0.404539
R11054 VCTRL2.n46 VCTRL2.n36 0.401155
R11055 VCTRL2.n9 VCTRL2.n8 0.401155
R11056 VCTRL2.n40 VCTRL2.n39 0.401155
R11057 VCTRL2.n104 VCTRL2.n103 0.400353
R11058 VCTRL2.n70 VCTRL2.n69 0.400178
R11059 VCTRL2.n47 VCTRL2.n46 0.398905
R11060 VCTRL2.n10 VCTRL2.n9 0.398484
R11061 VCTRL2.n55 VCTRL2.n47 0.397919
R11062 VCTRL2.n114 VCTRL2.n105 0.397919
R11063 VCTRL2.n105 VCTRL2.n104 0.397753
R11064 VCTRL2.n110 VCTRL2.n109 0.397744
R11065 VCTRL2.n7 VCTRL2.n6 0.389969
R11066 VCTRL2.n102 VCTRL2.n101 0.389723
R11067 VCTRL2.n38 VCTRL2.n37 0.389723
R11068 VCTRL2.n35 VCTRL2.n28 0.389547
R11069 VCTRL2.n32 VCTRL2.n31 0.389547
R11070 VCTRL2 VCTRL2.n125 0.10046
R11071 VCTRL2.n123 VCTRL2.n62 0.0698976
R11072 VCTRL2.n3 VCTRL2.n0 0.0695909
R11073 VCTRL2.n121 VCTRL2 0.0362534
R11074 VCTRL2.n2 VCTRL2 0.0362534
R11075 VCTRL2.n123 VCTRL2.n122 0.0124277
R11076 VCTRL2.n61 VCTRL2.n3 0.00395428
R11077 VCTRL2.n121 VCTRL2.n120 0.00173288
R11078 VCTRL2.n2 VCTRL2.n1 0.00173288
R11079 DN_INPUT.t0 DN_INPUT.t3 44.058
R11080 DN_INPUT.n0 DN_INPUT.t1 38.8649
R11081 DN_INPUT.t1 DN_INPUT.t0 28.6791
R11082 DN_INPUT.n0 DN_INPUT.t2 7.3005
R11083 DN_INPUT DN_INPUT.n0 5.27587
R11084 S6.t5 S6.t9 144.929
R11085 S6.t2 S6.t11 44.058
R11086 S6.n6 S6.t12 25.9486
R11087 S6.t12 S6 15.8807
R11088 S6.n1 S6.n0 15.8172
R11089 S6.n2 S6.n1 15.8172
R11090 S6.n5 S6.t5 14.796
R11091 S6.n5 S6.t2 13.8835
R11092 S6.n3 S6.t1 13.7188
R11093 S6.n8 S6.n6 13.2388
R11094 S6.n7 S6.t3 12.3193
R11095 S6.n0 S6.t7 11.7326
R11096 S6.n0 S6.t4 11.7326
R11097 S6.n1 S6.t8 11.7326
R11098 S6.n1 S6.t6 11.7326
R11099 S6.n2 S6.t10 11.7326
R11100 S6.t1 S6.n2 11.7326
R11101 S6 S6.n5 9.83964
R11102 S6.n6 S6.t0 7.3005
R11103 S6.n10 S6.n9 2.87402
R11104 S6.n4 S6.n3 2.3068
R11105 S6.n9 S6.n8 1.43443
R11106 S6.n8 S6.n7 0.391571
R11107 S6 S6.n10 0.176591
R11108 S6.n10 S6.n4 0.0139921
R11109 OUT.n7 OUT.t27 23.6945
R11110 OUT.t31 OUT.n8 23.6945
R11111 OUT.n34 OUT.t20 23.6945
R11112 OUT.t15 OUT.n35 23.6945
R11113 OUT.n8 OUT.n7 18.8035
R11114 OUT.n35 OUT.n34 18.8035
R11115 OUT.n5 OUT.n3 15.8172
R11116 OUT.n4 OUT.n0 15.8172
R11117 OUT.n5 OUT.n4 15.8172
R11118 OUT.n32 OUT.n30 15.8172
R11119 OUT.n32 OUT.n31 15.8172
R11120 OUT.n31 OUT.n27 15.8172
R11121 OUT.n3 OUT.t16 14.8925
R11122 OUT.t22 OUT.n5 14.8925
R11123 OUT.n4 OUT.t35 14.8925
R11124 OUT.n30 OUT.t34 14.8925
R11125 OUT.t21 OUT.n32 14.8925
R11126 OUT.n31 OUT.t32 14.8925
R11127 OUT.n9 OUT.n1 12.2457
R11128 OUT.n6 OUT.n1 12.2457
R11129 OUT.n6 OUT.n2 12.2457
R11130 OUT.n36 OUT.n28 12.2457
R11131 OUT.n33 OUT.n28 12.2457
R11132 OUT.n33 OUT.n29 12.2457
R11133 OUT.n10 OUT.t23 11.6285
R11134 OUT.n37 OUT.t28 11.6285
R11135 OUT.n2 OUT.t27 8.9065
R11136 OUT.t29 OUT.n6 8.9065
R11137 OUT.t18 OUT.n1 8.9065
R11138 OUT.n9 OUT.t31 8.9065
R11139 OUT.n29 OUT.t20 8.9065
R11140 OUT.t33 OUT.n33 8.9065
R11141 OUT.t19 OUT.n28 8.9065
R11142 OUT.n36 OUT.t15 8.9065
R11143 OUT.n5 OUT.t25 8.6145
R11144 OUT.n3 OUT.t17 8.6145
R11145 OUT.n4 OUT.t14 8.6145
R11146 OUT.n32 OUT.t30 8.6145
R11147 OUT.n30 OUT.t24 8.6145
R11148 OUT.n31 OUT.t12 8.6145
R11149 OUT.n0 OUT.t26 8.59715
R11150 OUT.n27 OUT.t13 8.59715
R11151 OUT.t16 OUT.n2 8.3225
R11152 OUT.n6 OUT.t22 8.3225
R11153 OUT.t35 OUT.n1 8.3225
R11154 OUT.t23 OUT.n9 8.3225
R11155 OUT.t34 OUT.n29 8.3225
R11156 OUT.n33 OUT.t21 8.3225
R11157 OUT.t32 OUT.n28 8.3225
R11158 OUT.t28 OUT.n36 8.3225
R11159 OUT.n40 OUT 4.9636
R11160 OUT OUT.n10 4.223
R11161 OUT OUT.n37 4.223
R11162 OUT.n7 OUT.t29 3.6505
R11163 OUT.n8 OUT.t18 3.6505
R11164 OUT.n34 OUT.t33 3.6505
R11165 OUT.n35 OUT.t19 3.6505
R11166 OUT.n14 OUT.t0 3.6405
R11167 OUT.n14 OUT.n13 3.6405
R11168 OUT.n12 OUT.t6 3.6405
R11169 OUT.n12 OUT.n11 3.6405
R11170 OUT.n21 OUT.t2 3.6405
R11171 OUT.n21 OUT.n20 3.6405
R11172 OUT.n19 OUT.t7 3.6405
R11173 OUT.n19 OUT.n18 3.6405
R11174 OUT.n26 OUT.n17 3.50463
R11175 OUT.n25 OUT.n24 3.50463
R11176 OUT.n17 OUT.t11 3.2765
R11177 OUT.n17 OUT.n16 3.2765
R11178 OUT.n24 OUT.t9 3.2765
R11179 OUT.n24 OUT.n23 3.2765
R11180 OUT.n10 OUT.n0 3.1807
R11181 OUT.n37 OUT.n27 3.1807
R11182 OUT.n15 OUT.n12 3.06224
R11183 OUT.n22 OUT.n19 3.06224
R11184 OUT.n15 OUT.n14 2.6005
R11185 OUT.n22 OUT.n21 2.6005
R11186 OUT OUT.n40 1.41493
R11187 OUT.n38 OUT 1.24006
R11188 OUT.n26 OUT.n25 0.798761
R11189 OUT.n39 OUT.n38 0.611422
R11190 OUT OUT.n26 0.562022
R11191 OUT.n38 OUT 0.247022
R11192 OUT.n40 OUT.n39 0.202264
R11193 OUT.n39 OUT 0.19218
R11194 OUT.n26 OUT.n15 0.18637
R11195 OUT.n25 OUT.n22 0.18637
R11196 S3.t5 S3.t12 144.929
R11197 S3.t0 S3.t1 44.058
R11198 S3.n6 S3.t9 25.9486
R11199 S3.t9 S3 15.8807
R11200 S3.n1 S3.n0 15.8172
R11201 S3.n2 S3.n1 15.8172
R11202 S3.n5 S3.t5 14.796
R11203 S3.n5 S3.t0 13.8835
R11204 S3.n3 S3.t3 13.7188
R11205 S3.n8 S3.n6 13.2388
R11206 S3.n7 S3.t6 12.3193
R11207 S3.n0 S3.t7 11.7326
R11208 S3.n0 S3.t4 11.7326
R11209 S3.n1 S3.t10 11.7326
R11210 S3.n1 S3.t8 11.7326
R11211 S3.n2 S3.t11 11.7326
R11212 S3.t3 S3.n2 11.7326
R11213 S3 S3.n5 9.83964
R11214 S3.n6 S3.t2 7.3005
R11215 S3.n10 S3.n9 2.87402
R11216 S3.n4 S3.n3 2.3068
R11217 S3.n9 S3.n8 1.43443
R11218 S3.n8 S3.n7 0.391571
R11219 S3 S3.n10 0.176591
R11220 S3.n10 S3.n4 0.0139921
R11221 ITAIL1.n5 ITAIL1.n4 28.0418
R11222 ITAIL1.n3 ITAIL1.n2 14.6005
R11223 ITAIL1.n1 ITAIL1.n0 7.61735
R11224 ITAIL1.n1 ITAIL1.t7 7.20135
R11225 ITAIL1.n8 ITAIL1.n7 6.82463
R11226 ITAIL1.n10 ITAIL1.t4 6.77907
R11227 ITAIL1.n5 ITAIL1.t0 6.71389
R11228 ITAIL1.n2 ITAIL1.t11 6.51836
R11229 ITAIL1.n2 ITAIL1.t2 6.51836
R11230 ITAIL1.n3 ITAIL1.t10 6.51836
R11231 ITAIL1.n10 ITAIL1.t12 6.25764
R11232 ITAIL1.n4 ITAIL1.t6 6.25764
R11233 ITAIL1.n6 ITAIL1.t13 6.19246
R11234 ITAIL1.n11 ITAIL1.t5 5.89613
R11235 ITAIL1.n11 ITAIL1.n10 4.23548
R11236 ITAIL1.n8 ITAIL1.n6 4.21461
R11237 ITAIL1.n13 ITAIL1 2.59768
R11238 ITAIL1 ITAIL1.n13 2.36014
R11239 ITAIL1.n9 ITAIL1.n8 1.42665
R11240 ITAIL1.n12 ITAIL1.n11 1.13763
R11241 ITAIL1.n13 ITAIL1.n12 0.501708
R11242 ITAIL1.n12 ITAIL1.n9 0.474918
R11243 ITAIL1.n4 ITAIL1.n3 0.261214
R11244 ITAIL1.n9 ITAIL1.n1 0.2105
R11245 ITAIL1.n6 ITAIL1.n5 0.130857
R11246 UP.n1 UP.n0 14.6005
R11247 UP.n3 UP.n2 12.8446
R11248 UP.n0 UP.t3 6.51836
R11249 UP.n0 UP.t7 6.51836
R11250 UP.n1 UP.t5 6.51836
R11251 UP.n3 UP.t4 6.388
R11252 UP.n2 UP.t6 6.19246
R11253 UP.n10 UP.n9 5.47387
R11254 UP.n4 UP.n3 5.03263
R11255 UP.n11 UP.n7 4.65398
R11256 UP.n10 UP.n8 4.2255
R11257 UP.n5 UP 2.32152
R11258 UP.n6 UP 2.0124
R11259 UP UP.n4 1.20571
R11260 UP.n6 UP.n5 0.85728
R11261 UP.n12 UP.n6 0.515191
R11262 UP.n11 UP.n10 0.427022
R11263 UP.n2 UP.n1 0.326393
R11264 UP.n12 UP 0.283382
R11265 UP UP.n11 0.257096
R11266 UP.n5 UP.n4 0.124995
R11267 UP UP.n12 0.00534345
R11268 DIV_OUT.t3 DIV_OUT.t2 44.058
R11269 DIV_OUT.n0 DIV_OUT.t0 38.8649
R11270 DIV_OUT.t0 DIV_OUT.t3 28.6791
R11271 DIV_OUT.n0 DIV_OUT.t1 7.3005
R11272 DIV_OUT DIV_OUT.n0 5.27587
R11273 S4.n16 S4.t18 45.6363
R11274 S4.n12 S4.t13 29.6446
R11275 S4.t14 S4.n13 29.6446
R11276 S4.n11 S4.t20 24.6117
R11277 S4.n5 S4.t6 23.6945
R11278 S4.n6 S4.t12 23.6945
R11279 S4.n13 S4.n12 22.2047
R11280 S4.t18 S4.t3 22.1925
R11281 S4.n17 S4.n16 20.9314
R11282 S4.n6 S4.n5 18.8035
R11283 S4 S4.t14 18.5175
R11284 S4.n3 S4.n0 15.8172
R11285 S4.n9 S4.n8 15.8172
R11286 S4.n8 S4.n0 15.8172
R11287 S4.t9 S4.n3 14.8925
R11288 S4.t15 S4.n0 14.8925
R11289 S4.n8 S4.t4 14.8925
R11290 S4.n7 S4.n1 12.2457
R11291 S4.n7 S4.n2 12.2457
R11292 S4.n4 S4.n2 12.2457
R11293 S4.n10 S4.t16 11.6285
R11294 S4.t6 S4.n4 8.9065
R11295 S4.t11 S4.n2 8.9065
R11296 S4.n7 S4.t0 8.9065
R11297 S4.t12 S4.n1 8.9065
R11298 S4.n3 S4.t10 8.6145
R11299 S4.n0 S4.t17 8.6145
R11300 S4.n8 S4.t5 8.6145
R11301 S4.n9 S4.t19 8.59715
R11302 S4.n4 S4.t9 8.3225
R11303 S4.n2 S4.t15 8.3225
R11304 S4.t4 S4.n7 8.3225
R11305 S4.n1 S4.t16 8.3225
R11306 S4.n11 S4.t7 6.1325
R11307 S4.n12 S4.t1 6.1325
R11308 S4.n13 S4.t2 6.1325
R11309 S4.n16 S4.t8 6.1325
R11310 S4.n17 S4.t21 6.1325
R11311 S4.n18 S4.n17 4.86779
R11312 S4.n14 S4.n11 4.79907
R11313 S4 S4.n10 4.223
R11314 S4.n5 S4.t11 3.6505
R11315 S4.t0 S4.n6 3.6505
R11316 S4.n10 S4.n9 3.1807
R11317 S4.n19 S4.n18 2.65123
R11318 S4.n14 S4 0.640368
R11319 S4.n15 S4 0.1655
R11320 S4.n18 S4.n15 0.109537
R11321 S4.n19 S4 0.0733182
R11322 S4.n15 S4.n14 0.0592755
R11323 S4 S4.n19 0.0318393
R11324 S2.t1 S2.t0 144.929
R11325 S2.t6 S2.t2 44.058
R11326 S2.n4 S2.t10 25.8834
R11327 S2.t10 S2 15.9445
R11328 S2.n1 S2.n0 15.8172
R11329 S2.n2 S2.n1 15.8172
R11330 S2.n3 S2.t1 14.7309
R11331 S2.n3 S2.t6 13.9487
R11332 S2.n8 S2.t4 13.7337
R11333 S2.n6 S2.n4 13.2388
R11334 S2.n5 S2.t11 12.2541
R11335 S2.n0 S2.t7 11.7326
R11336 S2.n0 S2.t3 11.7326
R11337 S2.n1 S2.t12 11.7326
R11338 S2.n1 S2.t9 11.7326
R11339 S2.n2 S2.t8 11.7326
R11340 S2.t4 S2.n2 11.7326
R11341 S2 S2.n3 9.83964
R11342 S2.n4 S2.t5 7.3005
R11343 S2.n9 S2.n8 2.30789
R11344 S2.n7 S2.n6 1.49961
R11345 S2.n8 S2.n7 0.546054
R11346 S2.n6 S2.n5 0.391571
R11347 S2 S2.n10 0.176591
R11348 S2.n10 S2.n9 0.0139921
R11349 S1.t1 S1.t7 144.929
R11350 S1.t9 S1.t11 44.058
R11351 S1.n4 S1.t6 25.8834
R11352 S1.t6 S1 15.9445
R11353 S1.n1 S1.n0 15.8172
R11354 S1.n2 S1.n1 15.8172
R11355 S1.n3 S1.t1 14.7309
R11356 S1.n3 S1.t9 13.9487
R11357 S1.n8 S1.t3 13.7337
R11358 S1.n6 S1.n4 13.2388
R11359 S1.n5 S1.t12 12.2541
R11360 S1.n0 S1.t2 11.7326
R11361 S1.n0 S1.t10 11.7326
R11362 S1.n1 S1.t8 11.7326
R11363 S1.n1 S1.t4 11.7326
R11364 S1.n2 S1.t5 11.7326
R11365 S1.t3 S1.n2 11.7326
R11366 S1 S1.n3 9.83964
R11367 S1.n4 S1.t0 7.3005
R11368 S1.n9 S1.n8 2.30789
R11369 S1.n7 S1.n6 1.49961
R11370 S1.n8 S1.n7 0.546054
R11371 S1.n6 S1.n5 0.391571
R11372 S1 S1.n10 0.176591
R11373 S1.n10 S1.n9 0.0139921
R11374 PRE_SCALAR.t0 PRE_SCALAR.t2 44.058
R11375 PRE_SCALAR.n0 PRE_SCALAR.t1 38.8649
R11376 PRE_SCALAR.t1 PRE_SCALAR.t0 28.6791
R11377 PRE_SCALAR.n0 PRE_SCALAR.t3 7.3005
R11378 PRE_SCALAR PRE_SCALAR.n0 5.27587
R11379 ITAIL.n7 ITAIL.t10 10.9054
R11380 ITAIL.n0 ITAIL.t17 10.8613
R11381 ITAIL.n17 ITAIL.t23 10.773
R11382 ITAIL.n13 ITAIL.t26 10.6003
R11383 ITAIL.n0 ITAIL.t0 10.5984
R11384 ITAIL.n17 ITAIL.t8 10.5336
R11385 ITAIL.n7 ITAIL.t18 10.5336
R11386 ITAIL.n1 ITAIL.t21 10.5334
R11387 ITAIL.n35 ITAIL.t22 10.533
R11388 ITAIL.n34 ITAIL.t4 10.5098
R11389 ITAIL.n18 ITAIL.t27 10.4686
R11390 ITAIL.n16 ITAIL.t12 10.0514
R11391 ITAIL.n10 ITAIL.t2 9.72546
R11392 ITAIL.n4 ITAIL.t6 9.65907
R11393 ITAIL.n36 ITAIL.t14 9.29485
R11394 ITAIL.n37 ITAIL.t19 8.47237
R11395 ITAIL.n29 ITAIL.t7 8.17686
R11396 ITAIL.n24 ITAIL.t13 8.07837
R11397 ITAIL.n25 ITAIL.n23 7.98962
R11398 ITAIL.n30 ITAIL.n28 7.84993
R11399 ITAIL.n29 ITAIL.t1 7.79699
R11400 ITAIL.n32 ITAIL.n26 7.73548
R11401 ITAIL.n24 ITAIL.t9 7.72811
R11402 ITAIL.n31 ITAIL.n27 7.58076
R11403 ITAIL.n39 ITAIL.n38 3.7682
R11404 ITAIL.n32 ITAIL.n31 1.75757
R11405 ITAIL.n20 ITAIL.n16 1.50725
R11406 ITAIL.n11 ITAIL.n10 1.50717
R11407 ITAIL.n6 ITAIL.n5 1.49748
R11408 ITAIL.n39 ITAIL 1.10761
R11409 ITAIL.n31 ITAIL.n30 0.661924
R11410 ITAIL.n14 ITAIL.n6 0.490305
R11411 ITAIL.n21 ITAIL.n14 0.446994
R11412 ITAIL.n37 ITAIL.n36 0.413008
R11413 ITAIL.n1 ITAIL.n0 0.390708
R11414 ITAIL.n36 ITAIL.n35 0.375243
R11415 ITAIL.n18 ITAIL.n17 0.365503
R11416 ITAIL.n19 ITAIL.n18 0.357915
R11417 ITAIL.n2 ITAIL.n1 0.357771
R11418 ITAIL.n13 ITAIL.n12 0.356995
R11419 ITAIL.n8 ITAIL.n7 0.341087
R11420 ITAIL.n33 ITAIL.n32 0.31096
R11421 ITAIL.n25 ITAIL.n24 0.301864
R11422 ITAIL.n30 ITAIL.n29 0.285711
R11423 ITAIL.n38 ITAIL.n22 0.278
R11424 ITAIL.n38 ITAIL.n37 0.244031
R11425 ITAIL.n33 ITAIL.n25 0.2255
R11426 ITAIL.n35 ITAIL.n34 0.201238
R11427 ITAIL.n34 ITAIL.n33 0.1493
R11428 ITAIL ITAIL.n39 0.0489615
R11429 ITAIL.n11 ITAIL.n8 0.028981
R11430 ITAIL.n14 ITAIL.n13 0.0236995
R11431 ITAIL.n21 ITAIL.n20 0.017375
R11432 ITAIL.n12 ITAIL.n11 0.0163348
R11433 ITAIL.n20 ITAIL.n19 0.0150187
R11434 ITAIL.n6 ITAIL.n3 0.013491
R11435 ITAIL.n3 ITAIL.n2 0.0117754
R11436 ITAIL.n22 ITAIL.n21 0.003875
R11437 ITAIL.n16 ITAIL.n15 0.00243623
R11438 ITAIL.n10 ITAIL.n9 0.00242648
R11439 ITAIL.n5 ITAIL.n4 0.00155882
R11440 OUTB.n27 OUTB 6.6528
R11441 OUTB.n6 OUTB.n5 5.81586
R11442 OUTB.n2 OUTB.t19 5.10151
R11443 OUTB.n8 OUTB.t16 5.1005
R11444 OUTB.n7 OUTB.t13 5.08021
R11445 OUTB.n2 OUTB.n1 4.66164
R11446 OUTB.n13 OUTB.t7 3.6405
R11447 OUTB.n13 OUTB.n12 3.6405
R11448 OUTB.n15 OUTB.t3 3.6405
R11449 OUTB.n15 OUTB.n14 3.6405
R11450 OUTB.n20 OUTB.t0 3.6405
R11451 OUTB.n20 OUTB.n19 3.6405
R11452 OUTB.n22 OUTB.t6 3.6405
R11453 OUTB.n22 OUTB.n21 3.6405
R11454 OUTB.n25 OUTB.n11 3.50463
R11455 OUTB.n24 OUTB.n18 3.50463
R11456 OUTB.n11 OUTB.t10 3.2765
R11457 OUTB.n11 OUTB.n10 3.2765
R11458 OUTB.n18 OUTB.t11 3.2765
R11459 OUTB.n18 OUTB.n17 3.2765
R11460 OUTB.n16 OUTB.n15 3.06224
R11461 OUTB.n23 OUTB.n22 3.06224
R11462 OUTB.n6 OUTB.n4 2.85093
R11463 OUTB.n16 OUTB.n13 2.6005
R11464 OUTB.n23 OUTB.n20 2.6005
R11465 OUTB.n4 OUTB.t14 2.16717
R11466 OUTB.n4 OUTB.n3 2.16717
R11467 OUTB.n1 OUTB.t18 1.9505
R11468 OUTB.n1 OUTB.n0 1.9505
R11469 OUTB.n27 OUTB.n26 1.47848
R11470 OUTB OUTB.n27 1.06887
R11471 OUTB.n25 OUTB.n24 0.798761
R11472 OUTB.n7 OUTB.n6 0.644196
R11473 OUTB OUTB.n25 0.562022
R11474 OUTB.n8 OUTB.n7 0.447229
R11475 OUTB.n9 OUTB.n2 0.308586
R11476 OUTB.n9 OUTB.n8 0.277162
R11477 OUTB.n25 OUTB.n16 0.18637
R11478 OUTB.n24 OUTB.n23 0.18637
R11479 OUTB.n26 OUTB 0.161224
R11480 OUTB OUTB.n9 0.115935
R11481 OUTB.n26 OUTB 0.0483126
R11482 DN.t7 DN.t5 12.5148
R11483 DN.n3 DN.t7 10.2564
R11484 DN.n0 DN.t4 10.1117
R11485 DN.n1 DN.t6 9.54068
R11486 DN.n2 DN.t8 9.4755
R11487 DN.n0 DN.t3 9.4755
R11488 DN.n7 DN.n5 5.47387
R11489 DN.n9 DN.n8 4.65398
R11490 DN.n7 DN.n6 4.2255
R11491 DN.n4 DN 1.15322
R11492 DN.n4 DN 0.960106
R11493 DN.n2 DN.n1 0.50481
R11494 DN.n1 DN.n0 0.501707
R11495 DN.n9 DN.n7 0.427022
R11496 DN.n3 DN.n2 0.332569
R11497 DN DN.n9 0.257096
R11498 DN DN.n3 0.2505
R11499 DN DN.n4 0.0373182
R11500 F_IN.t3 F_IN.t1 44.058
R11501 F_IN.n0 F_IN.t0 38.8649
R11502 F_IN.t0 F_IN.t3 28.6791
R11503 F_IN.n0 F_IN.t2 7.3005
R11504 F_IN F_IN.n0 5.27587
R11505 F_IN.n1 F_IN 2.02926
R11506 F_IN.n1 F_IN 1.4172
R11507 F_IN F_IN.n1 0.00465837
R11508 VCTRL_IN.n3 VCTRL_IN.n2 5.81586
R11509 VCTRL_IN.n5 VCTRL_IN.t7 5.10208
R11510 VCTRL_IN.n8 VCTRL_IN.t5 5.10194
R11511 VCTRL_IN.n4 VCTRL_IN.t1 5.08021
R11512 VCTRL_IN.n8 VCTRL_IN.n7 4.66114
R11513 VCTRL_IN.n3 VCTRL_IN.n1 2.85093
R11514 VCTRL_IN.n1 VCTRL_IN.t2 2.16717
R11515 VCTRL_IN.n1 VCTRL_IN.n0 2.16717
R11516 VCTRL_IN.n7 VCTRL_IN.t4 1.9505
R11517 VCTRL_IN.n7 VCTRL_IN.n6 1.9505
R11518 VCTRL_IN.n4 VCTRL_IN.n3 0.644196
R11519 VCTRL_IN.n5 VCTRL_IN.n4 0.449473
R11520 VCTRL_IN.n9 VCTRL_IN.n8 0.21214
R11521 VCTRL_IN.n9 VCTRL_IN.n5 0.198571
R11522 VCTRL_IN VCTRL_IN.n9 0.0718949
R11523 UP_INPUT.t2 UP_INPUT.t1 44.058
R11524 UP_INPUT.n0 UP_INPUT.t0 38.8649
R11525 UP_INPUT.t0 UP_INPUT.t2 28.6791
R11526 UP_INPUT.n0 UP_INPUT.t3 7.3005
R11527 UP_INPUT UP_INPUT.n0 5.27587
C0 a_20097_10547# PRE_SCALAR 0.002f
C1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 1.21f
C2 a_44716_1837# OUT 0.00801f
C3 PFD_T2_0.INV_mag_0.IN S2 0.0531f
C4 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_1284# 0.893f
C5 PFD_T2_0.Buffer_V_2_0.IN a_25557_8739# 0.182f
C6 VCO_DFF_C_0.VCO_C_0.OUT VCTRL2 0.0145f
C7 a_20097_10547# F_IN 0.123f
C8 a_27722_10564# UP_INPUT 0.23f
C9 mux_magic_0.OR_magic_0.B mux_magic_1.OR_magic_0.B 4.14e-20
C10 PFD_T2_0.INV_mag_0.IN a_22880_9797# 0.0939f
C11 a_46528_12082# VDD 0.257f
C12 a_43228_11254# a_43528_10426# 8.33e-21
C13 PFD_T2_0.UP S2 0.235f
C14 mux_magic_2.OR_magic_0.A mux_magic_3.OR_magic_0.A 0.00129f
C15 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCTRL2 0.344f
C16 a_43828_9804# VDD 0.257f
C17 a_42763_5679# VCTRL_IN 0.269f
C18 mux_magic_1.OR_magic_0.B UP 4.52e-19
C19 a_42928_8976# a_43228_9598# 0.0149f
C20 a_45628_9804# a_45328_8976# 8.33e-21
C21 a_45928_8976# VDD 0.257f
C22 PFD_T2_0.INV_mag_1.OUT a_22879_10704# 0.0502f
C23 a_27722_10564# a_27922_10564# 0.298f
C24 a_19897_10547# a_20103_9637# 4.68e-20
C25 a_22880_10947# PFD_T2_0.INV_mag_0.OUT 0.00145f
C26 PFD_T2_0.INV_mag_1.IN mux_magic_3.OR_magic_0.B 4.1e-19
C27 PFD_T2_0.FIN a_22967_8787# 2.04e-19
C28 a_31468_10271# VDD 1.1f
C29 S6 DIV_OUT 0.296f
C30 a_45328_8770# a_45628_8148# 0.0149f
C31 VDD ITAIL1 0.775f
C32 a_27922_11758# S2 0.00329f
C33 VDD PRE_SCALAR 0.898f
C34 mux_magic_1.AND2_magic_0.A a_28075_8520# 0.029f
C35 a_19903_8443# a_20103_8443# 0.296f
C36 a_29415_8145# a_27875_8520# 7.98e-19
C37 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN m1_33892_1807# 0.00112f
C38 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 0.624f
C39 PFD_T2_0.Buffer_V_2_0.IN a_24437_9224# 0.603f
C40 mux_magic_3.AND2_magic_0.A a_21443_8068# 3.58e-20
C41 a_29415_9553# DN 0.127f
C42 UP_INPUT S3 8.12e-19
C43 a_44728_12082# a_44428_11254# 8.33e-21
C44 VDD F_IN 0.364f
C45 PFD_T2_0.FIN S2 9.36e-19
C46 a_43228_11254# a_43228_9804# 0.00239f
C47 a_46228_11460# VDD 0.255f
C48 mux_magic_1.OR_magic_0.A PFD_T2_0.DOWN 0.00118f
C49 a_27922_10564# S3 0.00562f
C50 RES_74k_1.P a_42628_11254# 0.0457f
C51 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_0.OUT 0.479f
C52 PFD_T2_0.FIN a_22880_9797# 3.78e-20
C53 a_19897_10547# a_19903_9637# 0.00402f
C54 mux_magic_0.OR_magic_0.A mux_magic_1.OR_magic_0.B 9.11e-20
C55 mux_magic_2.OR_magic_0.B S2 0.00863f
C56 RES_74k_1.P a_44728_10426# 0.00241f
C57 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUTB 0.0234f
C58 a_23836_10693# VDD 0.0011f
C59 a_44428_9598# a_44128_8770# 8.33e-21
C60 a_45028_8148# a_45628_8148# 0.0415f
C61 a_25556_11637# S2 0.00926f
C62 VCO_DFF_C_0.VCO_C_0.OUTB OUT 0.00703f
C63 mux_magic_1.AND2_magic_0.A a_27875_8520# 0.251f
C64 a_43228_11460# a_43528_12082# 0.0149f
C65 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.OUTB 0.0222f
C66 a_44428_11460# a_44428_11254# 0.227f
C67 PFD_T2_0.Buffer_V_2_1.IN a_22967_8787# 7.01e-23
C68 a_42928_10632# a_43228_9804# 8.33e-21
C69 a_45328_10632# a_45628_11254# 0.0149f
C70 a_44128_10426# a_44728_10426# 0.0415f
C71 a_19897_10547# S6 1.08e-19
C72 a_22966_11778# a_22881_9554# 4.4e-22
C73 a_45328_10426# a_45628_9598# 8.33e-21
C74 a_24436_11277# a_22879_10704# 0.00339f
C75 a_44128_8976# a_44128_8770# 0.227f
C76 RES_74k_1.P a_44428_9804# 0.0106f
C77 a_22880_10947# VDD 0.0329f
C78 S4 OUTB 0.0286f
C79 a_44428_8148# VCO_DFF_C_0.VCTRL 0.00231f
C80 RES_74k_1.P a_46528_8976# 0.0572f
C81 a_21437_10708# a_21443_9476# 0.0202f
C82 PFD_T2_0.Buffer_V_2_1.IN S2 0.0205f
C83 mux_magic_2.OR_magic_0.A S2 0.00163f
C84 RES_74k_1.M a_43528_12082# 0.00176f
C85 VCO_DFF_C_0.VCTRL a_25706_n567# 6.1e-19
C86 a_44428_11460# a_44128_10632# 8.33e-21
C87 mux_magic_2.OR_magic_0.B mux_magic_3.OR_magic_0.B 0.00142f
C88 a_31940_9626# DN 2.33e-20
C89 a_43528_10426# VDD 0.257f
C90 a_44128_10426# a_44428_9804# 0.0149f
C91 a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.00276f
C92 a_45628_9598# VDD 0.257f
C93 a_45328_10426# a_45328_8976# 0.00239f
C94 RES_74k_1.P a_46828_11254# 0.096f
C95 PFD_T2_0.INV_mag_1.OUT VDD 0.708f
C96 a_46228_9598# a_46528_8976# 0.0149f
C97 a_44128_8976# a_43828_8148# 8.33e-21
C98 mux_magic_0.AND2_magic_0.A S2 0.593f
C99 a_27875_9714# DN 1.68e-19
C100 PFD_T2_0.INV_mag_0.IN UP_INPUT 4.06e-19
C101 a_29262_10725# ITAIL 0.00132f
C102 a_45928_12082# VDD 0.257f
C103 a_21437_10708# mux_magic_3.OR_magic_0.A 7e-19
C104 a_22966_11778# a_22967_8787# 0.0253f
C105 a_43228_11254# a_42928_10426# 8.33e-21
C106 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT 0.385f
C107 a_27875_9714# DN_INPUT 0.223f
C108 a_43828_9804# a_44428_9804# 0.0415f
C109 a_46528_10632# a_46528_10426# 0.227f
C110 a_43228_9804# VDD 0.257f
C111 a_41879_n196# VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.277f
C112 a_45328_8976# VDD 0.257f
C113 a_45028_9804# a_45328_8976# 8.33e-21
C114 a_42628_8770# a_42928_8976# 0.0415f
C115 PFD_T2_0.INV_mag_1.IN a_22879_10704# 0.0588f
C116 a_27722_10564# VDD 0.871f
C117 PFD_T2_0.UP UP_INPUT 0.127f
C118 a_45928_8976# a_46528_8976# 0.0415f
C119 mux_magic_2.OR_magic_0.A mux_magic_3.OR_magic_0.B 3.55e-21
C120 a_28075_9714# PFD_T2_0.DOWN 0.002f
C121 mux_magic_1.OR_magic_0.B DN 0.00106f
C122 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.00342f
C123 a_45028_8148# a_45328_8770# 0.0149f
C124 VDD DIV_OUT 0.899f
C125 mux_magic_0.OR_magic_0.B ITAIL 5.71e-19
C126 a_22966_11778# S2 0.00706f
C127 mux_magic_1.AND2_magic_0.A a_29415_8145# 3.58e-20
C128 PFD_T2_0.UP a_27922_10564# 0.002f
C129 a_42928_12082# a_43528_12082# 0.0415f
C130 PFD_T2_0.FDIV a_21443_8068# 1.35e-20
C131 mux_magic_1.OR_magic_0.B DN_INPUT 0.00118f
C132 UP ITAIL 0.634f
C133 a_46528_12082# a_46828_11254# 0.0149f
C134 a_44128_12082# a_44428_11254# 8.33e-21
C135 a_27922_11758# UP_INPUT 0.00693f
C136 a_22966_11778# a_22880_9797# 3.25e-19
C137 a_42928_10632# a_42928_10426# 0.227f
C138 a_45028_11254# a_45628_11254# 0.0415f
C139 a_45628_11460# VDD 0.255f
C140 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 3.61e-20
C141 mux_magic_2.OR_magic_0.B a_19903_9637# 2.99e-21
C142 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 3.46e-19
C143 a_46528_10632# a_46228_9804# 8.33e-21
C144 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 3.19f
C145 VDD S3 2.58f
C146 a_42628_9598# a_43228_9598# 0.0415f
C147 a_19897_10547# a_20097_10547# 0.298f
C148 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_0.OUT 0.218f
C149 a_27922_11758# a_27922_10564# 0.0206f
C150 PFD_T2_0.INV_mag_0.IN a_22879_10704# 0.251f
C151 RES_74k_1.P a_44128_10426# 0.00241f
C152 a_24436_11277# VDD 0.275f
C153 a_43828_9598# a_44128_8770# 8.33e-21
C154 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD 2.87f
C155 RES_74k_1.P a_46228_9598# 0.0323f
C156 a_31732_10267# RES_74k_1.P 0.478f
C157 mux_magic_2.OR_magic_0.B UP_INPUT 1.47e-19
C158 mux_magic_0.OR_magic_0.A S2 1.1e-20
C159 a_42928_12082# a_43228_11460# 0.0149f
C160 a_28075_9714# DN_INPUT 0.12f
C161 PFD_T2_0.FDIV mux_magic_3.AND2_magic_0.A 8.78e-21
C162 a_44128_12082# a_44128_10632# 0.00239f
C163 a_46228_11460# a_46828_11254# 0.0415f
C164 a_25556_11637# UP_INPUT 4.14e-19
C165 a_45028_11254# a_45328_10632# 0.0149f
C166 a_42928_10632# a_42628_9804# 8.33e-21
C167 a_44716_1837# a_44716_n517# 7.6e-20
C168 RES_74k_1.P a_46528_12082# 0.272f
C169 a_42628_9598# a_42928_8976# 0.0149f
C170 a_45328_10426# a_45028_9598# 8.33e-21
C171 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.OUT 0.318f
C172 RES_74k_1.P a_43828_9804# 0.0108f
C173 a_43828_9598# a_43828_8148# 0.00239f
C174 a_19897_10547# VDD 0.871f
C175 a_43828_8148# VCO_DFF_C_0.VCTRL 0.00369f
C176 RES_74k_1.P a_45928_8976# 0.0103f
C177 a_31468_10271# RES_74k_1.P 5.88e-19
C178 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 7.97e-19
C179 PFD_T2_0.FIN a_22879_10704# 0.0578f
C180 a_21437_10708# S2 0.00407f
C181 a_42628_11460# a_43228_11460# 0.0415f
C182 PFD_T2_0.FDIV PFD_T2_0.Buffer_V_2_0.IN 0.00929f
C183 a_21443_9476# a_21443_8068# 0.475f
C184 RES_74k_1.M a_42928_12082# 0.0504f
C185 RES_74k_1.P ITAIL1 1.67f
C186 a_43828_11460# a_44128_10632# 8.33e-21
C187 PFD_T2_0.Buffer_V_2_1.IN UP_INPUT 1.54e-20
C188 a_28075_8520# S3 0.00329f
C189 a_44728_10632# a_45328_10632# 0.0415f
C190 mux_magic_2.OR_magic_0.B a_22879_10704# 1.09e-19
C191 mux_magic_1.OR_magic_0.A a_29415_9553# 0.0334f
C192 a_22967_8787# PFD_T2_0.DOWN 3.31e-20
C193 a_42928_10426# VDD 0.257f
C194 VCO_DFF_C_0.VCTRL VCTRL2 0.227f
C195 VDD OUTB 0.781f
C196 a_43828_9804# a_44128_10426# 0.0149f
C197 a_46228_11254# a_46528_10426# 8.33e-21
C198 RES_74k_1.P a_46228_11460# 0.00579f
C199 a_45028_9598# VDD 0.257f
C200 a_45028_9804# a_45028_9598# 0.227f
C201 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.765f
C202 PFD_T2_0.INV_mag_1.IN VDD 5f
C203 a_43528_8976# a_43828_8148# 8.33e-21
C204 a_45928_8976# a_46228_9598# 0.0149f
C205 A_MUX_0.Tr_Gate_1.CLK OUTB 0.00188f
C206 a_44728_8770# a_45328_8770# 0.0415f
C207 a_31468_10271# a_31732_10267# 0.492f
C208 a_21437_12116# S2 0.00468f
C209 PFD_T2_0.FIN PFD_T2_0.INV_mag_0.OUT 0.0515f
C210 a_21443_9476# mux_magic_3.AND2_magic_0.A 2.4e-20
C211 PFD_T2_0.DOWN S2 1.31e-20
C212 RES_74k_1.M a_42628_11460# 0.0167f
C213 a_31732_10267# ITAIL1 0.0371f
C214 VCO_DFF_C_0.VCO_C_0.OUT VDD 0.723f
C215 a_45328_12082# VDD 0.257f
C216 mux_magic_0.AND2_magic_0.A UP_INPUT 0.0757f
C217 a_27875_8520# S3 6.67e-19
C218 a_42628_10426# a_42928_10426# 0.0415f
C219 a_22967_8787# a_25557_8739# 4.4e-19
C220 mux_magic_3.OR_magic_0.A a_21443_8068# 0.397f
C221 a_42628_9804# VDD 0.257f
C222 a_46228_11254# a_46228_9804# 0.00239f
C223 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD 12.5f
C224 a_44728_8976# VDD 0.257f
C225 a_45028_9804# a_44728_8976# 8.33e-21
C226 a_21437_10708# mux_magic_3.OR_magic_0.B 7.12e-19
C227 PFD_T2_0.Buffer_V_2_1.IN a_22879_10704# 0.0325f
C228 a_25556_11637# PFD_T2_0.INV_mag_0.OUT 5.66e-19
C229 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.306f
C230 VCO_DFF_C_0.VCO_C_0.OUTB a_44716_n517# 9.39e-20
C231 mux_magic_0.AND2_magic_0.A a_27922_10564# 0.00103f
C232 PFD_T2_0.INV_mag_0.IN VDD 4.75f
C233 a_20103_8443# DIV_OUT 0.12f
C234 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.915f
C235 a_44728_8770# a_45028_8148# 0.0149f
C236 mux_magic_0.OR_magic_0.B UP_INPUT 0.00118f
C237 VCO_DFF_C_0.VCO_C_0.OUTB VCTRL_IN 0.00272f
C238 a_27722_11758# S2 6.67e-19
C239 a_21443_9476# PFD_T2_0.Buffer_V_2_0.IN 2.15e-20
C240 PFD_T2_0.UP VDD 0.981f
C241 a_27875_9714# a_29415_9553# 0.00114f
C242 a_31468_10271# ITAIL1 2.45e-19
C243 a_44128_12082# a_43828_11254# 8.33e-21
C244 a_46228_11460# a_46528_12082# 0.0149f
C245 a_42628_10426# a_42628_9804# 0.0149f
C246 a_45028_11460# VDD 0.255f
C247 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.419f
C248 a_22967_8787# a_24437_9224# 0.00175f
C249 mux_magic_3.OR_magic_0.A mux_magic_3.AND2_magic_0.A 0.00108f
C250 a_45928_10632# a_46228_9804# 8.33e-21
C251 S2 DN_INPUT 0.784f
C252 ITAIL DN 0.0315f
C253 a_42628_9598# a_42628_8770# 0.0149f
C254 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT OUT 0.577f
C255 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.OUT 0.00184f
C256 VCO_DFF_C_0.VCO_C_0.OUTB a_41879_n196# 0.72f
C257 a_27922_11758# VDD 0.0671f
C258 a_19903_8443# DIV_OUT 0.325f
C259 RES_74k_1.P a_43528_10426# 0.00282f
C260 a_43828_9598# a_43528_8770# 8.33e-21
C261 mux_magic_1.OR_magic_0.B a_29415_9553# 0.411f
C262 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN a_25706_n567# 0.854f
C263 PRE_SCALAR F_IN 0.0249f
C264 RES_74k_1.P a_45628_9598# 0.0313f
C265 a_44428_8148# a_45028_8148# 0.0415f
C266 a_20097_11741# a_20097_10547# 0.0206f
C267 PFD_T2_0.FIN VDD 0.802f
C268 a_42628_11460# a_42928_12082# 0.0149f
C269 a_43828_11460# a_43828_11254# 0.227f
C270 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK OUTB 0.493f
C271 a_42628_11254# a_42928_10426# 8.33e-21
C272 a_44728_10632# a_45028_11254# 0.0149f
C273 a_22880_9797# a_24437_9224# 0.00315f
C274 a_22967_8787# a_21443_8068# 9.91e-20
C275 a_27875_9714# mux_magic_1.OR_magic_0.A 0.00184f
C276 mux_magic_2.OR_magic_0.B VDD 1.19f
C277 a_43528_10426# a_44128_10426# 0.0415f
C278 RES_74k_1.P a_45928_12082# 0.228f
C279 VCO_DFF_C_0.VCO_C_0.OUTB a_44716_1837# 0.71f
C280 a_22966_11778# a_22879_10704# 0.372f
C281 a_44728_10426# a_45028_9598# 8.33e-21
C282 mux_magic_0.OR_magic_0.A a_27922_10564# 1.77e-19
C283 RES_74k_1.P a_43228_9804# 0.0113f
C284 a_25556_11637# VDD 0.501f
C285 a_45628_9598# a_46228_9598# 0.0415f
C286 mux_magic_2.OR_magic_0.A a_20097_10547# 1.77e-19
C287 a_43528_8976# a_43528_8770# 0.227f
C288 a_43228_8148# VCO_DFF_C_0.VCTRL 0.00368f
C289 a_22881_9554# PFD_T2_0.Buffer_V_2_0.IN 0.0369f
C290 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.OUT 9.22e-19
C291 VCO_DFF_C_0.VCTRL S4 0.523f
C292 RES_74k_1.P a_45328_8976# 0.00953f
C293 a_20097_11741# VDD 0.0578f
C294 mux_magic_1.OR_magic_0.B mux_magic_1.OR_magic_0.A 0.178f
C295 m1_33892_1807# VDD 0.0434f
C296 a_43828_11460# a_43528_10632# 8.33e-21
C297 a_42628_11254# a_42628_9804# 0.00239f
C298 a_43528_10426# a_43828_9804# 0.0149f
C299 a_23837_9553# PFD_T2_0.Buffer_V_2_0.IN 0.262f
C300 a_46228_11254# a_45928_10426# 8.33e-21
C301 RES_74k_1.P a_45628_11460# 0.00482f
C302 a_44428_9598# VDD 0.257f
C303 a_44728_10426# a_44728_8976# 0.00239f
C304 a_22966_11778# PFD_T2_0.INV_mag_0.OUT 0.0613f
C305 VCO_DFF_C_0.VCO_C_0.OUTB a_41879_1284# 0.121f
C306 PFD_T2_0.Buffer_V_2_1.IN VDD 1.18f
C307 a_45628_9598# a_45928_8976# 0.0149f
C308 a_43528_8976# a_43228_8148# 8.33e-21
C309 a_45158_5339# S4 0.0148f
C310 mux_magic_2.OR_magic_0.A VDD 1.23f
C311 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.13f
C312 a_22880_10947# a_23836_10693# 0.0514f
C313 a_29262_12133# VDD 1.6f
C314 m1_30034_1474# VDD 0.0163f
C315 a_28075_9714# mux_magic_1.OR_magic_0.A 1.77e-19
C316 a_21443_9476# PFD_T2_0.FDIV 0.133f
C317 a_20103_9637# S1 0.00147f
C318 a_45928_12082# a_46528_12082# 0.0415f
C319 a_44728_12082# VDD 0.257f
C320 PFD_T2_0.DOWN UP_INPUT 0.00739f
C321 mux_magic_1.AND2_magic_0.A S3 0.59f
C322 a_22967_8787# PFD_T2_0.Buffer_V_2_0.IN 0.0311f
C323 a_43228_9804# a_43828_9804# 0.0415f
C324 a_45928_10632# a_45928_10426# 0.227f
C325 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 0.391f
C326 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT 0.02f
C327 a_44128_8976# VDD 0.257f
C328 a_44428_9804# a_44728_8976# 8.33e-21
C329 a_21437_10708# a_22879_10704# 3.4e-19
C330 a_29262_10725# VDD 0.929f
C331 mux_magic_0.AND2_magic_0.A VDD 1.3f
C332 a_45328_8976# a_45928_8976# 0.0415f
C333 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.389f
C334 a_27875_9714# mux_magic_1.OR_magic_0.B 0.125f
C335 a_42763_5679# S4 0.719f
C336 mux_magic_3.OR_magic_0.B a_21443_8068# 0.173f
C337 a_44428_8148# a_44728_8770# 0.0149f
C338 PFD_T2_0.INV_mag_1.OUT a_23836_10693# 0.00331f
C339 a_43528_12082# a_43828_11254# 8.33e-21
C340 a_45928_12082# a_46228_11460# 0.0149f
C341 a_19903_9637# S1 1.08e-19
C342 a_27722_11758# UP_INPUT 0.00635f
C343 a_44428_11460# VDD 0.255f
C344 a_44428_11254# a_45028_11254# 0.0415f
C345 mux_magic_0.OR_magic_0.B VDD 1.2f
C346 a_22880_9797# PFD_T2_0.Buffer_V_2_0.IN 0.038f
C347 a_46528_10632# VDD 0.257f
C348 a_45928_10632# a_45628_9804# 8.33e-21
C349 VDD UP 0.998f
C350 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN m1_33892_1807# 0.106f
C351 a_21437_10708# PFD_T2_0.INV_mag_0.OUT 7.29e-19
C352 RES_74k_1.P a_42928_10426# 0.00384f
C353 a_46528_8770# VDD 0.255f
C354 a_43228_9598# a_43528_8770# 8.33e-21
C355 a_25706_n567# VCO_DFF_C_0.VCO_C_0.OUTB 1.54f
C356 a_22966_11778# VDD 2.85f
C357 mux_magic_2.AND2_magic_0.A a_20097_10547# 0.00103f
C358 UP_INPUT DN_INPUT 0.95f
C359 a_19897_11741# VDD 0.986f
C360 RES_74k_1.P OUTB 0.168f
C361 PFD_T2_0.FDIV a_22881_9554# 0.0955f
C362 a_27875_9714# a_28075_9714# 0.298f
C363 RES_74k_1.P a_45028_9598# 0.0309f
C364 PFD_T2_0.INV_mag_1.OUT a_22880_10947# 7.65e-19
C365 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCTRL2 0.321f
C366 a_27922_10564# DN_INPUT 0.00289f
C367 S1 S6 0.0283f
C368 a_45628_11460# a_46228_11460# 0.0415f
C369 a_43528_12082# a_43528_10632# 0.00239f
C370 a_44428_11254# a_44728_10632# 0.0149f
C371 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD 2.74f
C372 a_44728_10426# a_44428_9598# 8.33e-21
C373 RES_74k_1.P a_45328_12082# 0.227f
C374 RES_74k_1.P a_42628_9804# 0.0563f
C375 mux_magic_0.OR_magic_0.A VDD 1.24f
C376 a_46228_8148# VDD 0.261f
C377 a_42628_8148# VCO_DFF_C_0.VCTRL 0.00293f
C378 a_43228_9598# a_43228_8148# 0.00239f
C379 mux_magic_2.AND2_magic_0.A VDD 1.27f
C380 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.DOWN 7.95e-19
C381 a_20103_9637# mux_magic_3.AND2_magic_0.A 0.00103f
C382 a_19903_9637# a_21443_8068# 1.14e-19
C383 RES_74k_1.P a_44728_8976# 0.00937f
C384 a_22879_10704# DN_INPUT 6.16e-20
C385 a_43228_11460# a_43528_10632# 8.33e-21
C386 a_44128_10632# a_44728_10632# 0.0415f
C387 a_22967_8787# PFD_T2_0.FDIV 0.174f
C388 a_45628_11254# a_45928_10426# 8.33e-21
C389 a_43228_9804# a_43528_10426# 0.0149f
C390 VDD OUT 4.42f
C391 mux_magic_3.OR_magic_0.A a_21443_9476# 0.0334f
C392 a_19897_10547# F_IN 0.32f
C393 a_44428_9804# a_44428_9598# 0.227f
C394 a_43828_9598# VDD 0.257f
C395 RES_74k_1.P a_45028_11460# 0.00442f
C396 VCO_DFF_C_0.VCTRL VDD 12.8f
C397 a_21437_10708# VDD 0.931f
C398 a_42928_8976# a_43228_8148# 8.33e-21
C399 a_45328_8976# a_45628_9598# 0.0149f
C400 PFD_T2_0.INV_mag_0.OUT a_25557_8739# 0.00304f
C401 a_19903_9637# mux_magic_3.AND2_magic_0.A 1.03e-19
C402 A_MUX_0.Tr_Gate_1.CLK VCO_DFF_C_0.VCTRL 0.422f
C403 a_44128_8770# a_44728_8770# 0.0415f
C404 a_27722_10564# PFD_T2_0.INV_mag_1.OUT 8.07e-19
C405 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.348f
C406 PFD_T2_0.INV_mag_0.OUT DN_INPUT 0.142f
C407 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_n517# 0.855f
C408 a_44128_12082# VDD 0.257f
C409 a_46228_11254# VDD 0.257f
C410 a_45628_11254# a_45628_9804# 0.00239f
C411 a_22880_9797# PFD_T2_0.FDIV 0.0427f
C412 a_43528_8976# VDD 0.257f
C413 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN OUT 0.382f
C414 a_45158_5339# VDD 1.37f
C415 a_44428_9804# a_44128_8976# 8.33e-21
C416 mux_magic_3.AND2_magic_0.A S6 0.589f
C417 a_21437_12116# VDD 1.6f
C418 a_31940_9626# ITAIL 0.00128f
C419 PFD_T2_0.INV_mag_0.OUT a_24437_9224# 0.371f
C420 a_44128_8770# a_44428_8148# 0.0149f
C421 PFD_T2_0.INV_mag_1.OUT S3 6.87e-19
C422 PFD_T2_0.DOWN VDD 1.07f
C423 A_MUX_0.Tr_Gate_1.CLK a_45158_5339# 0.706f
C424 PFD_T2_0.INV_mag_1.IN a_23836_10693# 0.017f
C425 a_24436_11277# PFD_T2_0.INV_mag_1.OUT 0.0143f
C426 a_27875_9714# S2 3.71e-19
C427 a_43528_12082# a_43228_11254# 8.33e-21
C428 a_20097_10547# S1 0.0292f
C429 a_45628_11460# a_45928_12082# 0.0149f
C430 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 0.546f
C431 a_43828_11460# VDD 0.255f
C432 a_45928_10632# VDD 0.257f
C433 a_45328_10632# a_45628_9804# 8.33e-21
C434 a_22967_8787# a_21443_9476# 0.0163f
C435 a_42763_5679# VDD 1.2f
C436 S4 VCTRL_IN 0.548f
C437 a_27722_11758# VDD 0.996f
C438 a_43228_9598# a_42928_8770# 8.33e-21
C439 a_45928_8770# VDD 0.255f
C440 mux_magic_3.OR_magic_0.B PFD_T2_0.FDIV 1.24e-20
C441 a_25557_8739# VDD 0.507f
C442 RES_74k_1.P a_44428_9598# 0.0309f
C443 a_46528_8976# a_46528_8770# 0.227f
C444 A_MUX_0.Tr_Gate_1.CLK a_42763_5679# 0.00257f
C445 a_27722_10564# S3 0.0013f
C446 a_43828_8148# a_44428_8148# 0.0415f
C447 VDD DN 2.35f
C448 PFD_T2_0.INV_mag_0.IN a_23836_10693# 0.145f
C449 PFD_T2_0.INV_mag_1.IN a_22880_10947# 0.00927f
C450 VCO_DFF_C_0.VCO_C_0.OUTB VCTRL2 0.00407f
C451 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 1.63f
C452 a_23837_9553# a_22881_9554# 0.0514f
C453 VDD DN_INPUT 0.853f
C454 a_43228_11460# a_43228_11254# 0.227f
C455 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_1837# 0.855f
C456 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK OUT 0.00102f
C457 VDD S1 1.97f
C458 a_46828_11254# a_46528_10632# 0.0149f
C459 a_44128_10632# a_44428_11254# 0.0149f
C460 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.00756f
C461 a_22880_9797# a_21443_9476# 5.39e-19
C462 a_42928_10426# a_43528_10426# 0.0415f
C463 RES_74k_1.P a_44728_12082# 0.227f
C464 a_44128_10426# a_44428_9598# 8.33e-21
C465 a_46528_10426# a_46828_9598# 0.0149f
C466 PFD_T2_0.DOWN a_28075_8520# 0.12f
C467 a_42928_8976# a_42928_8770# 0.227f
C468 a_45628_8148# VDD 0.257f
C469 a_45028_9598# a_45628_9598# 0.0415f
C470 a_28075_9714# S2 0.00478f
C471 a_24437_9224# VDD 0.272f
C472 a_22967_8787# mux_magic_3.OR_magic_0.A 0.0014f
C473 RES_74k_1.P a_44128_8976# 0.00937f
C474 a_46528_8976# a_46228_8148# 8.33e-21
C475 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.OUT 0.229f
C476 PFD_T2_0.INV_mag_0.IN a_22880_10947# 0.22f
C477 a_25706_n567# VCTRL2 5.69f
C478 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.0108f
C479 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 0.388f
C480 a_22967_8787# a_22881_9554# 0.306f
C481 VCO_DFF_C_0.VCTRL a_34443_2598# 6.1e-19
C482 mux_magic_0.OR_magic_0.B a_29415_8145# 4.38e-20
C483 a_43228_11460# a_42928_10632# 8.33e-21
C484 mux_magic_2.OR_magic_0.B F_IN 0.00118f
C485 a_42928_10426# a_43228_9804# 0.0149f
C486 a_45628_11254# a_45328_10426# 8.33e-21
C487 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT 0.00912f
C488 a_44128_10426# a_44128_8976# 0.00239f
C489 PFD_T2_0.DOWN a_27875_8520# 0.223f
C490 a_20097_11741# PRE_SCALAR 0.12f
C491 a_43228_9598# VDD 0.257f
C492 RES_74k_1.P a_44428_11460# 0.00442f
C493 a_46228_9804# a_46828_9598# 0.0415f
C494 a_45028_9598# a_45328_8976# 0.0149f
C495 RES_74k_1.P a_46528_10632# 0.047f
C496 a_42928_8976# a_42628_8148# 8.33e-21
C497 a_22967_8787# a_23837_9553# 0.0324f
C498 mux_magic_3.OR_magic_0.B a_21443_9476# 0.411f
C499 a_19903_9637# PFD_T2_0.FDIV 1.83e-19
C500 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.Buffer_V_2_0.IN 0.187f
C501 RES_74k_1.P UP 0.00276f
C502 a_21443_8068# VDD 1.6f
C503 a_20097_11741# F_IN 0.00449f
C504 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_1.OUT 0.405f
C505 RES_74k_1.P a_46528_8770# 0.0724f
C506 a_28075_8520# DN_INPUT 0.00449f
C507 a_22880_9797# a_22881_9554# 0.145f
C508 a_45328_12082# a_45928_12082# 0.0415f
C509 PFD_T2_0.FIN a_22880_10947# 0.0855f
C510 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.403f
C511 PFD_T2_0.UP PFD_T2_0.INV_mag_1.OUT 0.0222f
C512 mux_magic_2.OR_magic_0.A PRE_SCALAR 0.00118f
C513 a_43528_12082# VDD 0.257f
C514 a_42628_9804# a_43228_9804# 0.0415f
C515 a_45328_10632# a_45328_10426# 0.227f
C516 a_45628_11254# VDD 0.257f
C517 a_42928_8976# VDD 0.257f
C518 a_43828_9804# a_44128_8976# 8.33e-21
C519 a_27875_8520# DN 1.63e-20
C520 a_44728_8976# a_45328_8976# 0.0415f
C521 a_22880_9797# a_23837_9553# 0.0428f
C522 a_46228_9598# a_46528_8770# 8.33e-21
C523 a_43828_8148# a_44128_8770# 0.0149f
C524 a_31732_10267# UP 0.0189f
C525 mux_magic_3.AND2_magic_0.A VDD 1.27f
C526 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT OUTB 0.00852f
C527 PFD_T2_0.INV_mag_1.IN a_24436_11277# 0.0616f
C528 PFD_T2_0.Buffer_V_2_1.IN a_23836_10693# 0.262f
C529 a_29262_10725# a_31468_10271# 9.93e-20
C530 RES_74k_1.P a_46228_8148# 0.279f
C531 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD 0.958f
C532 mux_magic_3.OR_magic_0.B mux_magic_3.OR_magic_0.A 0.178f
C533 a_45328_12082# a_45628_11460# 0.0149f
C534 a_42928_12082# a_43228_11254# 8.33e-21
C535 VCO_DFF_C_0.VCO_C_0.OUTB S4 0.0152f
C536 a_46528_12082# a_46528_10632# 0.00239f
C537 a_43828_11254# a_44428_11254# 0.0415f
C538 a_43228_11460# VDD 0.255f
C539 a_46828_11254# a_46228_11254# 0.0415f
C540 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCTRL2 0.0917f
C541 a_45328_10632# VDD 0.257f
C542 a_45328_10632# a_45028_9804# 8.33e-21
C543 a_45328_8770# VDD 0.255f
C544 RES_74k_1.P OUT 0.0217f
C545 a_42628_8770# a_42928_8770# 0.0415f
C546 a_22879_10704# PFD_T2_0.FDIV 5.53e-20
C547 PFD_T2_0.Buffer_V_2_0.IN VDD 1.3f
C548 a_27922_10564# a_27875_9714# 7.59e-19
C549 a_22880_9797# a_22967_8787# 0.372f
C550 a_19903_9637# a_21443_9476# 0.00114f
C551 RES_74k_1.P a_43828_9598# 0.0311f
C552 a_46228_9598# a_46228_8148# 0.00239f
C553 RES_74k_1.P VCO_DFF_C_0.VCTRL 1.41f
C554 a_31468_10271# UP 0.0593f
C555 a_25556_11637# PFD_T2_0.INV_mag_1.OUT 0.00986f
C556 PFD_T2_0.Buffer_V_2_1.IN a_22880_10947# 0.0368f
C557 a_27922_11758# a_27722_10564# 0.00308f
C558 PFD_T2_0.INV_mag_0.IN a_24436_11277# 0.342f
C559 a_44716_n517# VDD 1.24f
C560 UP ITAIL1 0.079f
C561 a_20103_9637# mux_magic_3.OR_magic_0.A 1.77e-19
C562 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD 14.8f
C563 a_42928_12082# a_42928_10632# 0.00239f
C564 a_45028_11460# a_45628_11460# 0.0415f
C565 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.00204f
C566 a_19897_11741# PRE_SCALAR 0.323f
C567 a_43828_11254# a_44128_10632# 0.0149f
C568 a_46228_11460# a_46528_10632# 8.33e-21
C569 RES_74k_1.M VDD 0.826f
C570 VDD VCTRL_IN 0.112f
C571 RES_74k_1.P a_44128_12082# 0.227f
C572 a_44128_10426# a_43828_9598# 8.33e-21
C573 a_46228_9804# a_46528_10426# 0.0149f
C574 RES_74k_1.P a_46228_11254# 0.00138f
C575 a_42628_8770# a_42628_8148# 0.0149f
C576 a_45028_8148# VDD 0.257f
C577 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.FDIV 0.0514f
C578 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD 2.15f
C579 a_29415_9553# VDD 0.926f
C580 RES_74k_1.P a_43528_8976# 0.00978f
C581 a_45928_8976# a_46228_8148# 8.33e-21
C582 RES_74k_1.P a_45158_5339# 0.269f
C583 a_22966_11778# a_23836_10693# 0.0324f
C584 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.OUT 0.135f
C585 a_28075_9714# UP_INPUT 0.00341f
C586 a_41879_n196# VDD 1.17f
C587 a_19903_9637# mux_magic_3.OR_magic_0.A 0.00184f
C588 mux_magic_3.OR_magic_0.B a_22967_8787# 0.00306f
C589 a_44716_n517# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 0.269f
C590 a_42628_11460# a_42928_10632# 8.33e-21
C591 RES_74k_1.M a_42628_10426# 7.3e-19
C592 mux_magic_2.AND2_magic_0.A PRE_SCALAR 0.545f
C593 a_43528_10632# a_44128_10632# 0.0415f
C594 a_27922_10564# a_28075_9714# 0.0196f
C595 a_42628_9804# a_42928_10426# 0.0149f
C596 a_45028_11254# a_45328_10426# 8.33e-21
C597 a_43828_9804# a_43828_9598# 0.227f
C598 PFD_T2_0.DOWN mux_magic_1.AND2_magic_0.A 0.406f
C599 RES_74k_1.P a_43828_11460# 0.00458f
C600 a_42628_8770# VDD 0.289f
C601 mux_magic_2.AND2_magic_0.A F_IN 0.0189f
C602 RES_74k_1.P a_45928_10632# 0.00217f
C603 a_44728_8976# a_45028_9598# 0.0149f
C604 a_42628_9598# a_42928_8770# 8.33e-21
C605 a_43528_8770# a_44128_8770# 0.0415f
C606 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.00977f
C607 RES_74k_1.P a_45928_8770# 0.00968f
C608 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_1.IN 1.33f
C609 a_25556_11637# a_24436_11277# 0.00805f
C610 a_22966_11778# a_22880_10947# 0.306f
C611 mux_magic_3.OR_magic_0.A S6 1.1e-20
C612 a_44716_1837# VDD 1.26f
C613 RES_74k_1.P DN 1.07e-19
C614 mux_magic_1.OR_magic_0.A VDD 1.24f
C615 a_29262_12133# a_27722_10564# 1.14e-19
C616 PFD_T2_0.FIN a_19897_10547# 1.84e-19
C617 PFD_T2_0.UP PFD_T2_0.INV_mag_1.IN 4.12e-19
C618 a_46528_12082# a_46228_11254# 8.33e-21
C619 a_42928_12082# VDD 0.257f
C620 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUT 0.791f
C621 a_45028_11254# a_45028_9804# 0.00239f
C622 a_45028_11254# VDD 0.257f
C623 mux_magic_3.AND2_magic_0.A a_20103_8443# 0.029f
C624 a_21443_8068# a_19903_8443# 7.98e-19
C625 a_43828_9804# a_43528_8976# 8.33e-21
C626 a_25557_8739# mux_magic_1.AND2_magic_0.A 5.85e-20
C627 mux_magic_1.AND2_magic_0.A DN 8.78e-21
C628 mux_magic_2.OR_magic_0.B a_19897_10547# 0.125f
C629 a_42628_9598# a_42628_8148# 0.00239f
C630 a_43528_8770# a_43828_8148# 0.0149f
C631 a_46228_9598# a_45928_8770# 8.33e-21
C632 PFD_T2_0.FDIV VDD 0.825f
C633 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_44716_n517# 0.737f
C634 a_29262_10725# a_27722_10564# 0.00114f
C635 PFD_T2_0.Buffer_V_2_1.IN a_24436_11277# 0.619f
C636 a_22966_11778# PFD_T2_0.INV_mag_1.OUT 0.00225f
C637 a_21437_10708# a_23836_10693# 1.64e-20
C638 mux_magic_1.AND2_magic_0.A DN_INPUT 0.0174f
C639 RES_74k_1.P a_45628_8148# 0.23f
C640 mux_magic_0.AND2_magic_0.A a_27722_10564# 1.03e-19
C641 a_41879_1284# VDD 1.34f
C642 a_31732_10267# DN 0.00226f
C643 a_19903_9637# a_22967_8787# 1.59e-20
C644 a_44716_1837# VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 1.06e-20
C645 a_31940_9626# VDD 0.00834f
C646 a_45028_11460# a_45328_12082# 0.0149f
C647 RES_74k_1.M a_42628_11254# 8.18e-19
C648 a_20097_11741# a_19897_10547# 0.00308f
C649 a_42628_11460# VDD 0.255f
C650 PFD_T2_0.FIN PFD_T2_0.INV_mag_1.IN 0.00909f
C651 a_46228_11460# a_46228_11254# 0.227f
C652 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 7.5e-19
C653 PFD_T2_0.UP PFD_T2_0.INV_mag_0.IN 1.06e-19
C654 a_44728_10632# VDD 0.257f
C655 a_44728_10632# a_45028_9804# 8.33e-21
C656 a_45928_10426# a_46528_10426# 0.0415f
C657 a_42628_9598# VDD 0.257f
C658 mux_magic_0.OR_magic_0.B a_27722_10564# 0.125f
C659 a_29415_9553# a_27875_8520# 7.16e-20
C660 mux_magic_3.AND2_magic_0.A a_19903_8443# 0.227f
C661 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 2.23e-19
C662 a_44728_8770# VDD 0.255f
C663 RES_74k_1.P a_43228_9598# 0.0316f
C664 a_27875_9714# VDD 0.871f
C665 a_45928_8976# a_45928_8770# 0.227f
C666 a_43228_8148# a_43828_8148# 0.0415f
C667 a_27722_10564# UP 7.57e-20
C668 a_25556_11637# PFD_T2_0.INV_mag_1.IN 0.00255f
C669 mux_magic_1.OR_magic_0.A a_28075_8520# 9.27e-19
C670 a_21437_10708# a_22880_10947# 6.37e-19
C671 mux_magic_2.OR_magic_0.A a_19897_10547# 0.00184f
C672 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 3.46e-19
C673 a_31468_10271# DN 1.4f
C674 VCO_DFF_C_0.VCO_C_0.OUTB VDD 5.93f
C675 PFD_T2_0.FIN PFD_T2_0.INV_mag_0.IN 0.144f
C676 a_43528_10632# a_43828_11254# 0.0149f
C677 DN ITAIL1 5.59e-19
C678 PFD_T2_0.UP a_27922_11758# 0.12f
C679 a_46228_11460# a_45928_10632# 8.33e-21
C680 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 0.809f
C681 S2 UP_INPUT 0.437f
C682 PFD_T2_0.INV_mag_0.OUT a_22881_9554# 0.00219f
C683 mux_magic_1.OR_magic_0.B VDD 1.19f
C684 RES_74k_1.P a_43528_12082# 0.227f
C685 a_43528_10426# a_43828_9598# 8.33e-21
C686 a_45928_10426# a_46228_9804# 0.0149f
C687 a_44428_8148# VDD 0.257f
C688 mux_magic_2.OR_magic_0.B PFD_T2_0.INV_mag_0.IN 3.92e-19
C689 a_44428_9598# a_45028_9598# 0.0415f
C690 RES_74k_1.P a_45628_11254# 4.03e-19
C691 a_27922_10564# S2 0.0292f
C692 S1 PRE_SCALAR 0.455f
C693 a_21443_9476# VDD 0.933f
C694 RES_74k_1.P a_42928_8976# 0.0108f
C695 a_45928_8976# a_45628_8148# 8.33e-21
C696 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_44716_1837# 0.0017f
C697 mux_magic_1.OR_magic_0.A a_27875_8520# 0.128f
C698 mux_magic_0.OR_magic_0.A a_27722_10564# 0.00184f
C699 a_25556_11637# PFD_T2_0.INV_mag_0.IN 0.0258f
C700 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.IN 0.0388f
C701 a_22966_11778# a_24436_11277# 0.00177f
C702 a_25706_n567# VDD 3.74e-19
C703 S1 F_IN 0.526f
C704 a_22879_10704# a_22967_8787# 3.24e-19
C705 PFD_T2_0.INV_mag_0.OUT a_23837_9553# 0.0019f
C706 a_42928_12082# a_42628_11254# 8.33e-21
C707 PFD_T2_0.UP a_25556_11637# 0.136f
C708 a_28075_9714# VDD 0.0133f
C709 a_45028_11254# a_44728_10426# 8.33e-21
C710 a_19903_9637# mux_magic_3.OR_magic_0.B 0.125f
C711 a_46828_9598# VDD 0.289f
C712 RES_74k_1.P a_43228_11460# 0.00512f
C713 a_43528_10426# a_43528_8976# 0.00239f
C714 a_45628_9804# a_46228_9804# 0.0415f
C715 a_27875_9714# a_28075_8520# 0.00308f
C716 RES_74k_1.P a_45328_10632# 0.00164f
C717 a_44428_9598# a_44728_8976# 0.0149f
C718 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK a_41879_1284# 0.708f
C719 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.403f
C720 a_22966_11778# a_19897_10547# 1.74e-20
C721 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN 0.428f
C722 RES_74k_1.P a_45328_8770# 0.00888f
C723 mux_magic_2.OR_magic_0.A PFD_T2_0.INV_mag_0.IN 2.07e-19
C724 a_19897_11741# a_19897_10547# 0.00638f
C725 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.DOWN 0.0184f
C726 mux_magic_2.OR_magic_0.B PFD_T2_0.FIN 3.02e-21
C727 PFD_T2_0.INV_mag_0.OUT a_22967_8787# 0.0704f
C728 mux_magic_3.OR_magic_0.A VDD 1.23f
C729 a_44728_12082# a_45328_12082# 0.0415f
C730 a_42628_11460# a_42628_11254# 0.227f
C731 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN m1_30034_1474# 0.00112f
C732 PFD_T2_0.UP PFD_T2_0.Buffer_V_2_1.IN 0.00913f
C733 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCTRL2 0.0273f
C734 a_45928_12082# a_46228_11254# 8.33e-21
C735 a_44428_11254# VDD 0.257f
C736 a_22881_9554# VDD 0.0315f
C737 a_44728_10632# a_44728_10426# 0.227f
C738 a_19903_9637# a_20103_9637# 0.298f
C739 a_29415_9553# a_29415_8145# 0.475f
C740 a_27875_9714# a_27875_8520# 0.00638f
C741 RES_74k_1.P RES_74k_1.M 0.231f
C742 a_43228_9804# a_43528_8976# 8.33e-21
C743 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.0179f
C744 RES_74k_1.P VCTRL_IN 4.84e-20
C745 a_44128_8976# a_44728_8976# 0.0415f
C746 PFD_T2_0.INV_mag_0.OUT S2 1.77e-20
C747 a_43228_8148# a_43528_8770# 0.0149f
C748 a_45628_9598# a_45928_8770# 8.33e-21
C749 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT OUT 0.0191f
C750 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 0.703f
C751 a_22966_11778# PFD_T2_0.INV_mag_1.IN 0.0645f
C752 RES_74k_1.P a_45028_8148# 0.229f
C753 mux_magic_2.AND2_magic_0.A a_19897_10547# 1.03e-19
C754 PFD_T2_0.INV_mag_1.OUT a_25557_8739# 6.07e-19
C755 PFD_T2_0.INV_mag_0.OUT a_22880_9797# 0.304f
C756 a_23837_9553# VDD 0.0011f
C757 a_44728_12082# a_45028_11460# 0.0149f
C758 a_28075_9714# a_28075_8520# 0.0206f
C759 PFD_T2_0.FIN PFD_T2_0.Buffer_V_2_1.IN 0.00914f
C760 a_45928_12082# a_45928_10632# 0.00239f
C761 a_43228_11254# a_43828_11254# 0.0415f
C762 a_20103_9637# S6 0.0292f
C763 PFD_T2_0.INV_mag_1.OUT DN_INPUT 0.216f
C764 a_44128_10632# VDD 0.257f
C765 mux_magic_0.AND2_magic_0.A PFD_T2_0.UP 0.374f
C766 a_44728_10632# a_44428_9804# 8.33e-21
C767 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD 12.6f
C768 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN OUTB 1.27f
C769 PFD_T2_0.FDIV a_19903_8443# 3.51e-20
C770 a_29415_9553# mux_magic_1.AND2_magic_0.A 2.4e-20
C771 mux_magic_3.AND2_magic_0.A F_IN 5.44e-19
C772 a_44128_8770# VDD 0.255f
C773 mux_magic_2.OR_magic_0.A mux_magic_2.OR_magic_0.B 0.178f
C774 RES_74k_1.P a_42628_8770# 0.105f
C775 a_45628_9598# a_45628_8148# 0.00239f
C776 PFD_T2_0.DOWN S3 0.248f
C777 mux_magic_1.OR_magic_0.A a_29415_8145# 0.397f
C778 a_22966_11778# PFD_T2_0.INV_mag_0.IN 0.806f
C779 PFD_T2_0.Buffer_V_2_1.IN a_25556_11637# 0.172f
C780 a_27722_11758# a_27722_10564# 0.00638f
C781 a_21437_10708# a_19897_10547# 0.00114f
C782 mux_magic_0.AND2_magic_0.A a_27922_11758# 0.029f
C783 PFD_T2_0.INV_mag_1.OUT a_24437_9224# 4.79e-19
C784 a_22967_8787# VDD 2.84f
C785 a_44428_11460# a_45028_11460# 0.0415f
C786 a_43228_11254# a_43528_10632# 0.0149f
C787 PFD_T2_0.UP a_22966_11778# 8.04e-20
C788 mux_magic_2.OR_magic_0.A a_20097_11741# 9.27e-19
C789 a_45628_11460# a_45928_10632# 8.33e-21
C790 a_19903_9637# S6 0.195f
C791 a_27722_10564# DN_INPUT 0.00169f
C792 OUTB OUT 0.5f
C793 a_46528_10426# VDD 0.257f
C794 RES_74k_1.P a_42928_12082# 0.228f
C795 a_43528_10426# a_43228_9598# 8.33e-21
C796 a_45628_9804# a_45928_10426# 0.0149f
C797 VCO_DFF_C_0.VCTRL OUTB 0.0294f
C798 a_43828_8148# VDD 0.257f
C799 VDD S2 3.19f
C800 a_45328_8976# a_45628_8148# 8.33e-21
C801 a_25557_8739# S3 0.0043f
C802 a_21437_12116# a_19897_10547# 1.14e-19
C803 mux_magic_1.OR_magic_0.A mux_magic_1.AND2_magic_0.A 0.00108f
C804 mux_magic_0.AND2_magic_0.A a_25556_11637# 1.24e-19
C805 a_27922_10564# UP_INPUT 0.123f
C806 a_31468_10271# a_29415_9553# 1.05e-21
C807 VDD ITAIL 6.65f
C808 a_22880_9797# VDD 0.048f
C809 PFD_T2_0.FIN a_22966_11778# 0.175f
C810 a_42928_10632# a_43528_10632# 0.0415f
C811 S3 DN_INPUT 0.215f
C812 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.OUT 0.0471f
C813 a_19897_11741# PFD_T2_0.FIN 2.69e-20
C814 PFD_T2_0.UP mux_magic_0.OR_magic_0.A 0.00118f
C815 a_24436_11277# DN_INPUT 0.00219f
C816 RES_74k_1.P a_31940_9626# 0.511f
C817 VDD VCTRL2 1.23f
C818 a_44428_11254# a_44728_10426# 8.33e-21
C819 a_46228_9804# VDD 0.257f
C820 a_43228_9804# a_43228_9598# 0.227f
C821 RES_74k_1.P a_42628_11460# 0.0501f
C822 a_27875_9714# a_29415_8145# 1.14e-19
C823 a_21443_9476# a_19903_8443# 7.16e-20
C824 RES_74k_1.P a_44728_10632# 0.00149f
C825 mux_magic_2.OR_magic_0.B a_22966_11778# 0.00382f
C826 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 3.31f
C827 a_44128_8976# a_44428_9598# 0.0149f
C828 a_46828_9598# a_46528_8976# 0.0149f
C829 a_42928_8770# a_43528_8770# 0.0415f
C830 RES_74k_1.P a_42628_9598# 0.0766f
C831 mux_magic_3.OR_magic_0.A a_20103_8443# 9.27e-19
C832 RES_74k_1.P a_44728_8770# 0.00873f
C833 mux_magic_0.OR_magic_0.A a_27922_11758# 9.27e-19
C834 a_21437_10708# PFD_T2_0.INV_mag_0.IN 0.00177f
C835 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 10.3f
C836 mux_magic_0.AND2_magic_0.A PFD_T2_0.Buffer_V_2_1.IN 2.76e-20
C837 PFD_T2_0.INV_mag_1.IN PFD_T2_0.DOWN 0.0028f
C838 mux_magic_1.OR_magic_0.B a_29415_8145# 0.173f
C839 a_29262_12133# a_29262_10725# 0.475f
C840 a_45928_12082# a_45628_11254# 8.33e-21
C841 mux_magic_2.AND2_magic_0.A PFD_T2_0.FIN 9.36e-21
C842 a_19897_11741# a_20097_11741# 0.296f
C843 mux_magic_0.AND2_magic_0.A a_29262_12133# 3.58e-20
C844 a_31732_10267# a_31940_9626# 4.66e-20
C845 a_20097_10547# a_20103_9637# 0.026f
C846 a_43828_11254# VDD 0.257f
C847 a_44428_11254# a_44428_9804# 0.00239f
C848 a_19897_10547# S1 0.195f
C849 mux_magic_3.OR_magic_0.B VDD 1.19f
C850 a_27875_9714# mux_magic_1.AND2_magic_0.A 1.03e-19
C851 a_43228_9804# a_42928_8976# 8.33e-21
C852 a_42928_8770# a_43228_8148# 0.0149f
C853 a_45628_9598# a_45328_8770# 8.33e-21
C854 a_22966_11778# PFD_T2_0.Buffer_V_2_1.IN 0.0278f
C855 mux_magic_3.OR_magic_0.A a_19903_8443# 0.128f
C856 a_21443_8068# S3 8.01e-19
C857 mux_magic_0.OR_magic_0.B a_29262_12133# 0.173f
C858 a_21437_12116# PFD_T2_0.INV_mag_0.IN 4.7e-20
C859 RES_74k_1.P a_44428_8148# 0.228f
C860 mux_magic_0.AND2_magic_0.A a_29262_10725# 2.4e-20
C861 mux_magic_2.OR_magic_0.A a_22966_11778# 0.00196f
C862 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN a_34443_2598# 0.756f
C863 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.Buffer_V_2_0.IN 0.0183f
C864 PFD_T2_0.INV_mag_0.OUT UP_INPUT 8.05e-19
C865 a_19897_11741# mux_magic_2.OR_magic_0.A 0.128f
C866 PFD_T2_0.INV_mag_1.IN a_25557_8739# 0.0341f
C867 a_29262_12133# UP 0.00982f
C868 a_44428_11460# a_44728_12082# 0.0149f
C869 mux_magic_3.AND2_magic_0.A DIV_OUT 0.508f
C870 a_21437_10708# PFD_T2_0.FIN 0.171f
C871 mux_magic_2.AND2_magic_0.A a_20097_11741# 0.029f
C872 a_45628_11460# a_45628_11254# 0.227f
C873 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 0.674f
C874 a_43528_10632# VDD 0.257f
C875 PFD_T2_0.INV_mag_1.IN DN_INPUT 0.0154f
C876 a_20097_10547# a_19903_9637# 4.66e-20
C877 a_44128_10632# a_44428_9804# 8.33e-21
C878 a_20103_9637# VDD 0.0124f
C879 a_45328_10426# a_45928_10426# 0.0415f
C880 mux_magic_0.OR_magic_0.B a_29262_10725# 0.411f
C881 a_31940_9626# ITAIL1 0.655f
C882 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD 2.59f
C883 mux_magic_2.OR_magic_0.B a_21437_10708# 0.411f
C884 a_43528_8770# VDD 0.255f
C885 RES_74k_1.P a_46828_9598# 0.117f
C886 a_42628_8148# a_43228_8148# 0.0415f
C887 a_45328_8976# a_45328_8770# 0.227f
C888 a_29262_10725# UP 0.15f
C889 mux_magic_0.AND2_magic_0.A UP 8.78e-21
C890 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCTRL2 0.108f
C891 mux_magic_2.AND2_magic_0.A mux_magic_2.OR_magic_0.A 0.00108f
C892 PFD_T2_0.INV_mag_1.IN a_24437_9224# 0.354f
C893 a_28075_9714# mux_magic_1.AND2_magic_0.A 0.00103f
C894 VCO_DFF_C_0.VCTRL m1_33892_1807# 5.46e-20
C895 a_21437_12116# PFD_T2_0.FIN 3.99e-20
C896 a_42928_10632# a_43228_11254# 0.0149f
C897 a_45628_11460# a_45328_10632# 8.33e-21
C898 mux_magic_0.OR_magic_0.A a_29262_12133# 0.397f
C899 PFD_T2_0.UP a_27722_11758# 0.223f
C900 a_20097_10547# S6 0.00148f
C901 PFD_T2_0.INV_mag_0.OUT a_22879_10704# 0.305f
C902 PFD_T2_0.INV_mag_0.IN DN_INPUT 0.0495f
C903 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.381f
C904 a_19903_9637# VDD 0.871f
C905 mux_magic_0.OR_magic_0.B UP 0.0202f
C906 a_42928_10426# a_43228_9598# 8.33e-21
C907 a_45328_10426# a_45628_9804# 0.0149f
C908 a_45928_10426# VDD 0.257f
C909 a_43228_8148# VDD 0.257f
C910 mux_magic_2.OR_magic_0.B a_21437_12116# 0.173f
C911 a_43828_9598# a_44428_9598# 0.0415f
C912 a_46828_9598# a_46228_9598# 0.0415f
C913 a_46528_10426# a_46528_8976# 0.00239f
C914 VDD S4 2.92f
C915 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 1.27f
C916 PFD_T2_0.UP DN_INPUT 0.0335f
C917 a_45328_8976# a_45028_8148# 8.33e-21
C918 mux_magic_0.OR_magic_0.A a_29262_10725# 0.0334f
C919 a_21437_10708# PFD_T2_0.Buffer_V_2_1.IN 3.23e-22
C920 a_27722_11758# a_27922_11758# 0.296f
C921 a_34443_2598# VCTRL2 6.39f
C922 PFD_T2_0.Buffer_V_2_0.IN S3 0.00112f
C923 A_MUX_0.Tr_Gate_1.CLK S4 0.403f
C924 mux_magic_2.OR_magic_0.A a_21437_10708# 0.0334f
C925 PFD_T2_0.INV_mag_1.IN a_21443_8068# 1.56e-19
C926 PFD_T2_0.INV_mag_0.IN a_24437_9224# 0.0719f
C927 mux_magic_0.AND2_magic_0.A mux_magic_0.OR_magic_0.A 0.00108f
C928 a_22880_10947# PFD_T2_0.FDIV 3e-20
C929 VDD UP_INPUT 0.693f
C930 VCO_DFF_C_0.VCTRL m1_30034_1474# 0.0168f
C931 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCTRL2 0.198f
C932 VDD S6 1.99f
C933 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_44716_n517# 0.0175f
C934 a_44428_11254# a_44128_10426# 8.33e-21
C935 a_27922_10564# VDD 0.0144f
C936 a_45628_9804# VDD 0.257f
C937 a_42928_10426# a_42928_8976# 0.00239f
C938 a_45028_9804# a_45628_9804# 0.0415f
C939 mux_magic_0.OR_magic_0.A mux_magic_0.OR_magic_0.B 0.178f
C940 RES_74k_1.P a_44128_10632# 0.00149f
C941 a_46228_9804# a_46528_8976# 8.33e-21
C942 a_43828_9598# a_44128_8976# 0.0149f
C943 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD 2.16f
C944 mux_magic_0.OR_magic_0.A UP 0.00973f
C945 RES_74k_1.P a_44128_8770# 0.00873f
C946 a_46228_8148# a_46528_8770# 0.0149f
C947 mux_magic_2.OR_magic_0.A a_21437_12116# 0.397f
C948 mux_magic_2.AND2_magic_0.A a_19897_11741# 0.228f
C949 mux_magic_2.OR_magic_0.B DN_INPUT 7.17e-19
C950 a_44128_12082# a_44728_12082# 0.0415f
C951 a_45328_12082# a_45628_11254# 8.33e-21
C952 a_43228_11254# VDD 0.257f
C953 a_25556_11637# DN_INPUT 0.0195f
C954 a_22879_10704# VDD 0.05f
C955 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_41879_n196# 0.0136f
C956 a_44128_10632# a_44128_10426# 0.227f
C957 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VDD 0.893f
C958 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.39f
C959 a_42628_9804# a_42928_8976# 8.33e-21
C960 a_43528_8976# a_44128_8976# 0.0415f
C961 a_42628_8148# a_42928_8770# 0.0149f
C962 a_45028_9598# a_45328_8770# 8.33e-21
C963 a_20097_11741# S1 0.00329f
C964 RES_74k_1.P a_46528_10426# 0.0479f
C965 RES_74k_1.P a_43828_8148# 0.229f
C966 a_21437_10708# a_22966_11778# 0.0165f
C967 a_19897_11741# a_21437_10708# 7.16e-20
C968 PFD_T2_0.INV_mag_1.IN PFD_T2_0.Buffer_V_2_0.IN 0.595f
C969 PFD_T2_0.INV_mag_1.OUT a_27875_9714# 3.67e-19
C970 a_44128_12082# a_44428_11460# 0.0149f
C971 mux_magic_1.OR_magic_0.A S3 1.1e-20
C972 a_27722_11758# a_29262_12133# 7.98e-19
C973 a_20103_9637# a_20103_8443# 0.0206f
C974 a_45328_12082# a_45328_10632# 0.00239f
C975 RES_74k_1.P ITAIL 1.83f
C976 a_44128_10632# a_43828_9804# 8.33e-21
C977 a_42928_10632# VDD 0.257f
C978 PFD_T2_0.Buffer_V_2_1.IN DN_INPUT 0.0136f
C979 a_46228_11254# a_46528_10632# 0.0149f
C980 mux_magic_2.OR_magic_0.A DN_INPUT 2.66e-20
C981 PFD_T2_0.INV_mag_0.OUT VDD 0.674f
C982 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_44716_1837# 0.343f
C983 VCTRL_IN OUTB 0.0234f
C984 mux_magic_2.OR_magic_0.A S1 1.1e-20
C985 a_42928_8770# VDD 0.255f
C986 a_46528_10426# a_46228_9598# 8.33e-21
C987 RES_74k_1.P a_46228_9804# 0.012f
C988 a_45028_9598# a_45028_8148# 0.00239f
C989 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT 1.19f
C990 a_21437_12116# a_22966_11778# 8.19e-19
C991 a_27722_11758# a_29262_10725# 7.16e-20
C992 mux_magic_2.AND2_magic_0.A a_21437_10708# 2.4e-20
C993 mux_magic_0.AND2_magic_0.A a_27722_11758# 0.251f
C994 a_19897_11741# a_21437_12116# 7.98e-19
C995 a_27722_10564# a_27875_9714# 0.00228f
C996 PFD_T2_0.INV_mag_0.IN PFD_T2_0.Buffer_V_2_0.IN 0.0412f
C997 a_29262_10725# DN 0.00133f
C998 a_43828_11460# a_44428_11460# 0.0415f
C999 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 10.4f
C1000 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.4f
C1001 a_19903_9637# a_20103_8443# 0.00308f
C1002 a_42628_10426# a_42928_10632# 0.0415f
C1003 a_45028_11460# a_45328_10632# 8.33e-21
C1004 a_31732_10267# ITAIL 1.52f
C1005 a_45928_10632# a_46528_10632# 0.0415f
C1006 a_20097_10547# VDD 0.0124f
C1007 mux_magic_0.AND2_magic_0.A DN_INPUT 2.04e-19
C1008 a_45328_10426# VDD 0.257f
C1009 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 5.91e-19
C1010 a_45028_9804# a_45328_10426# 0.0149f
C1011 RES_74k_1.P a_43828_11254# 1.61e-19
C1012 a_42628_8148# VDD 0.257f
C1013 a_46228_9804# a_46228_9598# 0.227f
C1014 PFD_T2_0.INV_mag_1.OUT a_28075_9714# 0.00238f
C1015 a_44728_8976# a_45028_8148# 8.33e-21
C1016 a_27722_11758# UP 1.63e-20
C1017 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.00409f
C1018 a_27875_9714# S3 0.195f
C1019 a_45928_8770# a_46528_8770# 0.0415f
C1020 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 1.2f
C1021 UP DN 0.547f
C1022 mux_magic_2.AND2_magic_0.A a_21437_12116# 3.58e-20
C1023 a_44716_1837# OUTB 8.01e-19
C1024 a_20103_8443# S6 0.00329f
C1025 a_19903_9637# a_19903_8443# 0.00638f
C1026 a_42628_11254# a_43228_11254# 0.0415f
C1027 a_22966_11778# DN_INPUT 0.00319f
C1028 a_31468_10271# ITAIL 0.0368f
C1029 a_43828_11254# a_44128_10426# 8.33e-21
C1030 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.652f
C1031 a_45028_9804# VDD 0.257f
C1032 a_19897_11741# S1 3.96e-19
C1033 ITAIL ITAIL1 0.0176f
C1034 a_46228_9804# a_45928_8976# 8.33e-21
C1035 RES_74k_1.P a_43528_10632# 0.0019f
C1036 a_43528_8976# a_43828_9598# 0.0149f
C1037 a_27722_10564# a_28075_9714# 5.95e-19
C1038 a_45158_5339# VCO_DFF_C_0.VCTRL 0.939f
C1039 A_MUX_0.Tr_Gate_1.CLK VDD 1.93f
C1040 a_45928_8770# a_46228_8148# 0.0149f
C1041 RES_74k_1.P a_43528_8770# 0.00914f
C1042 a_21443_9476# S3 6.49e-19
C1043 a_21437_12116# a_21437_10708# 0.475f
C1044 a_27722_11758# mux_magic_0.OR_magic_0.A 0.128f
C1045 RES_74k_1.P VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 5.27e-19
C1046 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT a_34443_2598# 0.939f
C1047 PFD_T2_0.INV_mag_1.IN PFD_T2_0.FDIV 0.149f
C1048 a_41879_1284# OUTB 0.27f
C1049 a_19903_8443# S6 3.96e-19
C1050 a_42628_11254# a_42928_10632# 0.0149f
C1051 a_45328_12082# a_45028_11254# 8.33e-21
C1052 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT 1.64f
C1053 PFD_T2_0.INV_mag_1.OUT a_23837_9553# 1.35e-20
C1054 a_22880_10947# a_22967_8787# 6.22e-22
C1055 a_42628_10426# VDD 0.289f
C1056 a_43828_11254# a_43828_9804# 0.00239f
C1057 a_42928_10426# a_42628_9598# 8.33e-21
C1058 mux_magic_2.AND2_magic_0.A S1 0.586f
C1059 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD 0.921f
C1060 a_28075_9714# S3 0.0292f
C1061 mux_magic_3.OR_magic_0.A DIV_OUT 0.00118f
C1062 a_42763_5679# VCO_DFF_C_0.VCTRL 0.93f
C1063 a_45028_9598# a_44728_8770# 8.33e-21
C1064 RES_74k_1.P a_45928_10426# 0.00309f
C1065 RES_74k_1.P a_43228_8148# 0.229f
C1066 RES_74k_1.P S4 0.0112f
C1067 a_45628_8148# a_46228_8148# 0.0415f
C1068 VCO_DFF_C_0.VCTRL DN 0.109f
C1069 PFD_T2_0.INV_mag_0.IN PFD_T2_0.FDIV 3.6e-22
C1070 VCO_DFF_C_0.VCO_C_0.OUTB OUTB 0.725f
C1071 a_43828_11460# a_44128_12082# 0.0149f
C1072 a_28075_8520# VDD 0.0611f
C1073 a_45028_11460# a_45028_11254# 0.227f
C1074 PFD_T2_0.INV_mag_1.OUT a_22967_8787# 5.92e-19
C1075 a_45928_10632# a_46228_11254# 0.0149f
C1076 a_43528_10632# a_43828_9804# 8.33e-21
C1077 a_44728_10426# a_45328_10426# 0.0415f
C1078 a_42628_9804# a_42628_9598# 0.227f
C1079 a_45928_10426# a_46228_9598# 8.33e-21
C1080 a_42763_5679# a_45158_5339# 0.0097f
C1081 RES_74k_1.P a_45628_9804# 0.011f
C1082 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN m1_30034_1474# 0.103f
C1083 a_44728_8976# a_44728_8770# 0.227f
C1084 a_45628_8148# VCO_DFF_C_0.VCTRL 7.83e-19
C1085 mux_magic_1.AND2_magic_0.A UP_INPUT 7.89e-20
C1086 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.OUTB 1.64f
C1087 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD 14.9f
C1088 PFD_T2_0.INV_mag_1.IN a_21443_9476# 0.0018f
C1089 PFD_T2_0.INV_mag_1.OUT S2 0.0248f
C1090 a_25557_8739# PFD_T2_0.DOWN 0.137f
C1091 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.618f
C1092 a_27875_8520# VDD 0.994f
C1093 a_45028_11460# a_44728_10632# 8.33e-21
C1094 a_20103_9637# F_IN 0.00296f
C1095 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD 3.8f
C1096 PFD_T2_0.INV_mag_1.OUT a_22880_9797# 0.037f
C1097 a_42628_11254# VDD 0.257f
C1098 PFD_T2_0.FIN PFD_T2_0.FDIV 0.00835f
C1099 PFD_T2_0.DOWN DN_INPUT 0.0322f
C1100 a_44728_10426# VDD 0.257f
C1101 a_44728_10426# a_45028_9804# 0.0149f
C1102 RES_74k_1.P a_43228_11254# 6.97e-19
C1103 a_43228_9598# a_43828_9598# 0.0415f
C1104 a_45928_10426# a_45928_8976# 0.00239f
C1105 a_44728_8976# a_44428_8148# 8.33e-21
C1106 VCO_DFF_C_0.VCO_C_0.OUT a_25706_n567# 0.939f
C1107 RES_74k_1.M m1_53234_16109# 0.782f
C1108 a_29262_10725# a_29415_9553# 0.00851f
C1109 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 1.21f
C1110 a_27722_10564# S2 0.195f
C1111 a_34443_2598# VDD 3.74e-19
C1112 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN a_25706_n567# 0.756f
C1113 a_20103_8443# VDD 0.0577f
C1114 a_42628_11254# a_42628_10426# 0.0149f
C1115 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VDD 0.795f
C1116 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 0.488f
C1117 PFD_T2_0.INV_mag_1.IN mux_magic_3.OR_magic_0.A 2.08e-19
C1118 a_43828_11254# a_43528_10426# 8.33e-21
C1119 a_25557_8739# DN_INPUT 6.6e-19
C1120 a_44428_9804# VDD 0.257f
C1121 a_44428_9804# a_45028_9804# 0.0415f
C1122 RES_74k_1.P a_42928_10632# 0.00291f
C1123 a_46528_8976# VDD 0.257f
C1124 a_45628_9804# a_45928_8976# 8.33e-21
C1125 a_43228_9598# a_43528_8976# 0.0149f
C1126 mux_magic_0.OR_magic_0.B a_29415_9553# 5.06e-19
C1127 a_29262_12133# mux_magic_1.OR_magic_0.A 4.38e-20
C1128 PFD_T2_0.INV_mag_1.IN a_22881_9554# 0.231f
C1129 RES_74k_1.P a_42928_8770# 0.0102f
C1130 a_29415_9553# UP 0.0018f
C1131 S2 S3 0.0293f
C1132 a_45628_8148# a_45928_8770# 0.0149f
C1133 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_44716_n517# 2.57e-20
C1134 a_27875_8520# a_28075_8520# 0.296f
C1135 a_24436_11277# S2 1.78e-19
C1136 a_43528_12082# a_44128_12082# 0.0415f
C1137 F_IN S6 0.0089f
C1138 a_19903_8443# VDD 0.986f
C1139 a_44728_12082# a_45028_11254# 8.33e-21
C1140 a_29262_10725# mux_magic_1.OR_magic_0.A 7.77e-19
C1141 a_46828_11254# VDD 0.289f
C1142 PFD_T2_0.INV_mag_1.IN a_23837_9553# 0.155f
C1143 a_43528_10632# a_43528_10426# 0.227f
C1144 a_45628_11254# a_46228_11254# 0.0415f
C1145 a_42928_8976# a_43528_8976# 0.0415f
C1146 PFD_T2_0.INV_mag_0.IN a_22881_9554# 1.57e-19
C1147 mux_magic_2.OR_magic_0.B a_21443_9476# 7.06e-19
C1148 RES_74k_1.P a_45328_10426# 0.00257f
C1149 a_44428_9598# a_44728_8770# 8.33e-21
C1150 RES_74k_1.P a_42628_8148# 0.274f
C1151 mux_magic_0.OR_magic_0.B mux_magic_1.OR_magic_0.A 8.13e-19
C1152 mux_magic_0.OR_magic_0.A a_29415_9553# 3.44e-19
C1153 a_44716_n517# OUT 0.00245f
C1154 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_n196# 0.902f
C1155 a_43528_12082# a_43828_11460# 0.0149f
C1156 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 1.57f
C1157 mux_magic_1.OR_magic_0.A UP 3.03e-19
C1158 a_29415_8145# VDD 1.6f
C1159 a_44728_12082# a_44728_10632# 0.00239f
C1160 PFD_T2_0.INV_mag_1.IN a_22967_8787# 0.855f
C1161 PFD_T2_0.INV_mag_0.IN a_23837_9553# 0.00872f
C1162 a_45628_11254# a_45928_10632# 0.0149f
C1163 a_43528_10632# a_43228_9804# 8.33e-21
C1164 mux_magic_3.OR_magic_0.B S3 0.00168f
C1165 VCO_DFF_C_0.VCTRL VCTRL_IN 1.25f
C1166 a_34443_2598# VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 0.854f
C1167 a_45928_10426# a_45628_9598# 8.33e-21
C1168 a_23836_10693# a_22879_10704# 0.0428f
C1169 RES_74k_1.P VDD 23.1f
C1170 RES_74k_1.P a_45028_9804# 0.0106f
C1171 a_44428_9598# a_44428_8148# 0.00239f
C1172 a_45028_8148# VCO_DFF_C_0.VCTRL 8.04e-19
C1173 a_20103_9637# DIV_OUT 0.002f
C1174 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.0107f
C1175 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 0.915f
C1176 PFD_T2_0.INV_mag_1.IN S2 0.00119f
C1177 PFD_T2_0.FIN a_22881_9554# 2.24e-20
C1178 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_44716_1837# 0.00328f
C1179 a_22966_11778# PFD_T2_0.FDIV 1.88e-19
C1180 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK 0.496f
C1181 mux_magic_2.OR_magic_0.A a_21443_9476# 7.01e-19
C1182 mux_magic_2.OR_magic_0.B mux_magic_3.OR_magic_0.A 3.55e-21
C1183 a_43228_11460# a_43828_11460# 0.0415f
C1184 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.DOWN 0.014f
C1185 RES_74k_1.M a_44128_12082# 3.99e-19
C1186 a_31940_9626# UP 0.13f
C1187 a_44428_11460# a_44728_10632# 8.33e-21
C1188 mux_magic_1.AND2_magic_0.A VDD 1.29f
C1189 PFD_T2_0.INV_mag_1.OUT UP_INPUT 0.0197f
C1190 PFD_T2_0.INV_mag_0.IN a_22967_8787# 0.0259f
C1191 PFD_T2_0.INV_mag_1.IN a_22880_9797# 0.196f
C1192 a_45328_10632# a_45928_10632# 0.0415f
C1193 a_44128_10426# VDD 0.257f
C1194 a_45158_5339# VCTRL_IN 3.4e-22
C1195 a_44428_9804# a_44728_10426# 0.0149f
C1196 RES_74k_1.P a_42628_10426# 0.099f
C1197 a_46228_9598# VDD 0.257f
C1198 a_45628_9804# a_45628_9598# 0.227f
C1199 a_23836_10693# PFD_T2_0.INV_mag_0.OUT 7.19e-20
C1200 a_29262_10725# mux_magic_1.OR_magic_0.B 4.91e-19
C1201 a_22880_10947# a_22879_10704# 0.145f
C1202 PFD_T2_0.INV_mag_1.OUT a_27922_10564# 0.00279f
C1203 a_31732_10267# VDD 5.23f
C1204 mux_magic_0.OR_magic_0.B a_27875_9714# 3.31e-19
C1205 a_44128_8976# a_44428_8148# 8.33e-21
C1206 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT a_34443_2598# 1.53f
C1207 a_27875_9714# UP 1.04e-20
C1208 a_45328_8770# a_45928_8770# 0.0415f
.ends

