** sch_path:
*+ /home/shahid/GF180Projects/PGA_Decoder/Folded_OPAMP_nobias/Xschem/folded_single_TB_slew.sch
**.subckt folded_single_TB_slew
V5 VDD GND 3.3
.save i(v5)
V2 VINP GND pulse(0.2 1.6 0 100p 100p 50n 100n)
.save i(v2)
V1 VSS GND 0
.save i(v1)
I1 IBIAS VSS 50u
C1 OUTo VSS 20p m=1
x1 OUT VDD VSS OUTo VINP IBIAS VBS2 VBS3 VBIASN OUTo pex_fold_cascode_opamp_mag
**** begin user architecture code


.include pex_fold_cascode_opamp_mag.spice
.control
*save all
*.options savecurrents
save all

tran 100p 200n
*dc V4 0 3 10m
*plot v(IBIAS)
plot i(V5)
plot v(OUTo) v(VINP)

*write pmos_nmos.raw
*let vdiff = @m.xm1.m0[vdsat]+vds
*plot @m.xm1.m0[vdsat]
*tran 1u 2m
*let gain = (maximum(out1)-minimum(out2) )* 1000
*print vbb

*plot vdiff
*display all
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
* .lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_statistical

**** end user architecture code
**.ends
.GLOBAL GND
.end
