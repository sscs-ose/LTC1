* NGSPICE file created from TG_5x_Layout.ext - technology: gf180mcuC

.subckt nmos_3p3_FGGST2 a_n52_n50# a_n516_n50# a_428_n50# a_n428_n94# a_n212_n50#
+ a_n372_n50# a_52_n94# a_108_n50# a_268_n50# a_n108_n94# a_n268_n94# a_212_n94# a_372_n94#
+ VSUBS
X0 a_108_n50# a_52_n94# a_n52_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1 a_268_n50# a_212_n94# a_108_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 a_n372_n50# a_n428_n94# a_n516_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X3 a_428_n50# a_372_n94# a_268_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 a_n52_n50# a_n108_n94# a_n212_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 a_n212_n50# a_n268_n94# a_n372_n50# VSUBS nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
.ends

.subckt pmos_3p3_MN2VAR a_n292_n100# a_28_n100# a_n28_n144# a_132_n144# a_188_n100#
+ w_n522_n230# a_n188_n144# a_292_n144# a_348_n100# a_n348_n144# a_n436_n100# a_n132_n100#
X0 a_n132_n100# a_n188_n144# a_n292_n100# w_n522_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_188_n100# a_132_n144# a_28_n100# w_n522_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X2 a_n292_n100# a_n348_n144# a_n436_n100# w_n522_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 a_348_n100# a_292_n144# a_188_n100# w_n522_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X4 a_28_n100# a_n28_n144# a_n132_n100# w_n522_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_GGGST2 a_n28_n94# a_n116_n50# a_28_n50# VSUBS
X0 a_28_n50# a_n28_n94# a_n116_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt pmos_3p3_MNVUAR w_n202_n230# a_28_n100# a_n28_n144# a_n116_n100#
X0 a_28_n100# a_n28_n144# a_n116_n100# w_n202_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
.ends

.subckt Inverter_Layout IN OUT VSS VDD
Xnmos_3p3_GGGST2_0 IN VSS OUT VSS nmos_3p3_GGGST2
Xpmos_3p3_MNVUAR_0 VDD OUT IN VDD pmos_3p3_MNVUAR
.ends

.subckt TG_5x_Layout VIN VOUT VSS VDD CLK
Xnmos_3p3_FGGST2_0 VIN VOUT VOUT CLK VOUT VIN CLK VOUT VIN CLK CLK CLK CLK VSS nmos_3p3_FGGST2
Xpmos_3p3_MN2VAR_0 VIN VIN Inverter_Layout_0/OUT Inverter_Layout_0/OUT VOUT VDD Inverter_Layout_0/OUT
+ Inverter_Layout_0/OUT VIN Inverter_Layout_0/OUT VOUT VOUT pmos_3p3_MN2VAR
XInverter_Layout_0 CLK Inverter_Layout_0/OUT VSS VDD Inverter_Layout
.ends

