magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3367 -2147 14129 12917
<< polysilicon >>
rect 803 8900 1033 8996
rect 2677 8900 2907 8996
rect 3151 8900 3381 8996
rect 5025 8900 5255 8996
rect 5499 8900 5729 8996
rect 7373 8900 7603 8996
rect 7847 8900 8077 8996
rect 9721 8900 9951 8996
rect 803 1028 1033 1124
rect 2677 1028 2907 1124
rect 3151 1028 3381 1124
rect 5025 1028 5255 1124
rect 5499 1028 5729 1124
rect 7373 1028 7603 1124
rect 7847 1028 8077 1124
rect 9721 1028 9951 1124
<< metal1 >>
rect -440 9400 5218 9508
rect -440 9240 3344 9340
rect -440 9080 2870 9180
rect -440 8920 996 9020
rect 2708 8988 2870 9080
rect 3182 8988 3344 9240
rect 5056 8988 5218 9400
rect 5532 9400 11180 9508
rect 5532 8988 5694 9400
rect 7404 9240 11180 9340
rect 7404 8988 7566 9240
rect 7883 9080 11180 9180
rect 7883 8988 8045 9080
rect 893 1079 939 8920
rect 2772 1079 2818 8926
rect 3242 1079 3288 8926
rect 5114 1079 5160 8926
rect 5588 1079 5634 8926
rect 7462 1079 7508 8926
rect 7941 1079 7987 8926
rect 9756 8920 11180 9020
rect 9814 1079 9860 8920
use comp018green_out_drv_nleg_4T  comp018green_out_drv_nleg_4T_0
timestamp 1713338890
transform 1 0 597 0 1 680
box 48 444 2468 8220
use comp018green_out_drv_nleg_4T  comp018green_out_drv_nleg_4T_1
timestamp 1713338890
transform 1 0 2945 0 1 680
box 48 444 2468 8220
use comp018green_out_drv_nleg_4T  comp018green_out_drv_nleg_4T_2
timestamp 1713338890
transform 1 0 5293 0 1 680
box 48 444 2468 8220
use comp018green_out_drv_nleg_4T  comp018green_out_drv_nleg_4T_3
timestamp 1713338890
transform 1 0 7641 0 1 680
box 48 444 2468 8220
use GR_NMOS_4T  GR_NMOS_4T_0
timestamp 1713338890
transform 1 0 363 0 1 436
box -1730 -583 11766 10481
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform 0 1 915 1 0 8954
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform 0 1 915 1 0 1082
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_2
timestamp 1713338890
transform 0 1 2789 1 0 1082
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_3
timestamp 1713338890
transform 0 1 3263 1 0 8954
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_4
timestamp 1713338890
transform 0 1 2789 1 0 8954
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_5
timestamp 1713338890
transform 0 1 3263 1 0 1082
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_6
timestamp 1713338890
transform 0 1 5137 1 0 1082
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_7
timestamp 1713338890
transform 0 1 5137 1 0 8954
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_8
timestamp 1713338890
transform 0 1 7485 1 0 1082
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_9
timestamp 1713338890
transform 0 1 5611 1 0 1082
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_10
timestamp 1713338890
transform 0 1 7485 1 0 8954
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_11
timestamp 1713338890
transform 0 1 5611 1 0 8954
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_12
timestamp 1713338890
transform 0 1 9837 1 0 1082
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_13
timestamp 1713338890
transform 0 1 7964 1 0 1082
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_14
timestamp 1713338890
transform 0 1 7964 1 0 8954
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_15
timestamp 1713338890
transform 0 1 9837 1 0 8954
box -42 -89 42 89
use nmos_4T_metal_stack  nmos_4T_metal_stack_0
timestamp 1713338890
transform 1 0 603 0 1 812
box -44 400 2074 8000
use nmos_4T_metal_stack  nmos_4T_metal_stack_1
timestamp 1713338890
transform 1 0 2951 0 1 812
box -44 400 2074 8000
use nmos_4T_metal_stack  nmos_4T_metal_stack_2
timestamp 1713338890
transform 1 0 5299 0 1 812
box -44 400 2074 8000
use nmos_4T_metal_stack  nmos_4T_metal_stack_3
timestamp 1713338890
transform 1 0 7647 0 1 812
box -44 400 2074 8000
use nmos_4T_metal_stack  nmos_4T_metal_stack_4
timestamp 1713338890
transform -1 0 10151 0 1 812
box -44 400 2074 8000
<< end >>
