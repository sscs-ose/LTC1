* NGSPICE file created from CLK_div_93_mag_flat.ext - technology: gf180mcuC

.subckt CLK_div_93_mag_flat VSS Vdiv93 RST CLK VDD
X0 VDD CLK_div_31_mag_0.Q0.t3 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t432 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD.t181 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2 VDD CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t144 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 a_15342_208# CLK_div_3_mag_0.CLK a_15182_208# VSS.t212 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X4 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD.t104 VDD.t103 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X5 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t108 VSS.t107 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X6 VDD CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t136 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X7 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t140 VDD.t139 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 VDD VDD.t75 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X9 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t239 VDD.t238 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X10 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK VDD.t328 VDD.t327 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 VDD CLK_div_31_mag_0.Q1.t3 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t208 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X12 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD.t444 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 VDD CLK_div_31_mag_0.Q4.t2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t244 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X14 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t3 a_18365_1305# VSS.t89 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X15 VDD CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t271 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X16 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.Q4.t3 a_7249_360# VSS.t151 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X17 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VDD.t119 VDD.t118 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 VDD.t356 VDD.t355 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q2 a_9404_3954# VSS.t82 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X20 a_981_1449# VDD.t472 VSS.t51 VSS.t50 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X21 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VDD.t243 VDD.t242 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X22 a_7819_1501# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VSS.t153 VSS.t152 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X23 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 a_17194_252# VSS.t301 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X24 a_4023_1458# VDD.t473 VSS.t49 VSS.t48 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X25 a_18199_208# VDD.t474 VSS.t47 VSS.t46 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X26 a_5428_4226# CLK_div_31_mag_0.Q0.t4 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t285 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X27 VSS CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_1798_3130# VSS.t96 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X28 a_11989_2561# CLK_div_31_mag_0.Q4.t4 VDD.t406 VDD.t405 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X29 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_8383_1501# VSS.t126 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X30 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t252 VDD.t251 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X31 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VDD.t332 VDD.t331 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X32 a_4140_4226# CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t67 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X33 RST CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN VDD.t30 VDD.t29 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.QB a_4183_1458# VSS.t13 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X35 a_18365_1305# CLK_div_3_mag_0.CLK a_18205_1305# VSS.t211 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X36 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t32 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 VSS VDD.t475 a_2522_3130# VSS.t43 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X38 VSS CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_3730_3129# VSS.t258 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X39 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VDD.t412 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X40 a_16066_208# RST.t2 a_15906_208# VSS.t55 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X41 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VSS.t134 VSS.t133 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X42 VDD VDD.t71 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t72 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X43 VSS CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_1234_3130# VSS.t96 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X44 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q4.t5 a_7506_3203# VSS.t268 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X45 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X46 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT RST.t3 VDD.t91 VDD.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X47 VDD CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.Q4 VDD.t163 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X48 a_4183_1458# CLK_div_31_mag_0.Q2 a_4023_1458# VSS.t81 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X49 a_8383_1501# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VSS.t92 VSS.t91 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X50 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD.t68 VDD.t70 VDD.t69 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X51 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t287 VSS.t286 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X52 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.QB.t3 a_2833_1493# VSS.t272 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X53 a_4177_361# CLK_div_31_mag_0.Q2 a_4017_361# VSS.t80 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X54 a_1705_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t202 VSS.t201 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X55 VSS CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VSS.t273 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X56 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VDD.t440 VDD.t439 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X57 VSS VDD.t477 a_2528_4227# VSS.t40 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X58 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t100 VDD.t99 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X59 VDD CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t461 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X60 VDD CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t133 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X61 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t340 VDD.t339 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X62 a_1804_4227# RST.t4 a_1644_4227# VSS.t56 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X63 VDD CLK_div_31_mag_0.Q4.t6 CLK_div_31_mag_0.JK_FF_mag_4.QB VDD.t407 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X64 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 VDD.t438 VDD.t437 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X65 a_18923_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t17 VSS.t16 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X66 VDD RST.t5 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t184 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X67 VDD CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t268 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X68 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t254 VDD.t253 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X69 VDD CLK_div_31_mag_0.Q1.t4 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X70 a_16630_252# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t161 VSS.t160 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X71 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t93 VDD.t92 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X72 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VSS.t181 VSS.t180 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X73 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q2 a_8452_3208# VSS.t79 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X74 VDD CLK.t0 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD.t166 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X75 a_8453_3965# CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS.t234 VSS.t233 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X76 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t336 VDD.t335 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X77 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t387 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X78 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK VSS.t210 VSS.t209 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X79 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t352 VDD.t351 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X80 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD.t180 VDD.t179 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X81 VSS CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t175 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X82 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4747_1502# VSS.t195 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X83 a_4901_361# RST.t6 a_4741_361# VSS.t113 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X84 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0 a_19614_2684# VDD.t308 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X85 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t221 VDD.t220 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X86 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_16066_208# VSS.t222 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X87 VDD RST.t7 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t187 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X88 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.Q1.t5 VDD.t17 VDD.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X89 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t65 VDD.t67 VDD.t66 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X90 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.JK_FF_mag_1.QB a_5875_1502# VSS.t12 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X91 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t364 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X92 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t350 VDD.t349 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X93 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2423_396# VSS.t166 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X94 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 VDD.t460 VDD.t459 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X95 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_31_mag_0.Q2 VDD.t132 VDD.t131 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X96 a_8537_404# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VSS.t74 VSS.t73 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X97 a_1859_352# RST.t8 a_1699_352# VSS.t114 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X98 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5311_1502# VSS.t86 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X99 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_31_mag_0.Q3.t2 a_4177_361# VSS.t7 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X100 VDD CLK_div_31_mag_0.Q3.t3 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD.t79 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X101 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t160 VDD.t159 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X102 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t250 VDD.t249 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X103 a_5875_1502# CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t84 VSS.t83 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X104 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t4 VDD.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X105 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.Q0.t5 VDD.t431 VDD.t430 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X106 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t232 VDD.t231 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X107 VDD CLK.t1 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t169 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X108 CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t95 VDD.t94 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X109 VDD CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.Q0.t2 VDD.t392 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X110 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.Q1.t6 VSS.t9 VSS.t8 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X111 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t384 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X112 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q0.t6 VDD.t429 VDD.t428 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X113 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t147 VSS.t146 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X114 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD.t344 VDD.t343 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X115 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q0.t7 VDD.t427 VDD.t426 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X116 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.Q2 VSS.t78 VSS.t77 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X117 VSS CLK.t2 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS.t99 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X118 a_8947_1501# CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VSS.t150 VSS.t149 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X119 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VDD.t287 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X120 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK VSS.t208 VSS.t207 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X121 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 VDD.t458 VDD.t457 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X122 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VSS.t168 VSS.t167 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X123 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VDD.t368 VDD.t367 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X124 a_9404_3954# CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS.t288 VSS.t82 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X125 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t334 VDD.t333 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X126 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_31_mag_0.Q1.t0 VDD.t174 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X127 VDD CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD.t262 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X128 a_19083_208# RST.t9 a_18923_208# VSS.t115 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X129 VDD CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t1 VDD.t305 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X130 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 VDD.t373 VDD.t372 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X131 a_1798_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t96 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X132 VSS CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t198 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X133 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t257 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X134 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t217 VDD.t216 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X135 VSS CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_4858_3129# VSS.t162 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X136 CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_31_mag_0.or_2_mag_0.IN1 a_11989_2561# VDD.t282 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X137 a_18205_1305# CLK_div_3_mag_0.Q1 VSS.t300 VSS.t299 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X138 a_2522_3130# CLK_div_31_mag_0.Q0.t8 a_2362_3130# VSS.t43 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X139 a_3730_3129# CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.Q0.t0 VSS.t3 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X140 CLK_div_3_mag_0.CLK CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t284 VDD.t283 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X141 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q1 a_18641_2448# VSS.t298 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X142 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_31_mag_0.Q2 a_1135_352# VSS.t76 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X143 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t448 VDD.t447 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X144 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_31_mag_0.Q0.t9 VDD.t425 VDD.t424 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X145 a_1234_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t96 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X146 VSS VDD.t478 a_5582_3129# VSS.t37 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X147 a_7506_3203# CLK_div_31_mag_0.Q0.t10 VSS.t284 VSS.t268 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X148 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.QB VDD.t261 VDD.t260 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X149 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t330 VDD.t329 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X150 VSS CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VSS.t182 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X151 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.Q4.t7 a_9101_404# VSS.t269 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X152 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD.t156 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X153 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t441 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X154 VSS CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_4294_3129# VSS.t262 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X155 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_4.QB a_8947_1501# VSS.t98 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X156 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q3.t4 a_9403_3219# VSS.t52 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X157 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB a_15348_1305# VSS.t1 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X158 VDD CLK_div_3_mag_0.CLK CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t324 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X159 VDD CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t235 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X160 VSS CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_670_3130# VSS.t96 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X161 a_4858_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t130 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X162 VDD CLK_div_31_mag_0.Q3.t5 CLK_div_31_mag_0.JK_FF_mag_1.QB VDD.t82 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X163 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_4901_361# VSS.t156 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X164 a_2362_3130# CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t43 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X165 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2269_1493# VSS.t165 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X166 a_2833_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t158 VSS.t157 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X167 VDD CLK_div_31_mag_0.Q1.t7 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD.t18 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X168 a_5582_3129# CLK.t3 a_5422_3129# VSS.t102 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X169 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t281 VDD.t280 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X170 VDD CLK_div_3_mag_0.JK_FF_mag_1.K.t4 CLK_div_3_mag_0.Q0 VDD.t149 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 a_19647_252# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t242 VSS.t241 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X172 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t348 VDD.t347 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X173 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD.t342 VDD.t341 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X174 a_4294_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t66 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X175 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t88 VSS.t87 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X176 a_18929_1349# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t58 VSS.t57 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X177 VDD CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.QB.t0 VDD.t128 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X178 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 a_15342_208# VSS.t297 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X179 CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VSS.t236 VSS.t235 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X180 a_2528_4227# CLK_div_31_mag_0.Q0.t11 a_2368_4227# VSS.t283 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X181 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.CLK VDD.t323 VDD.t322 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X182 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_1859_352# VSS.t219 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X183 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t65 VSS.t64 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X184 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT RST.t10 VDD.t191 VDD.t190 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X185 a_670_3130# CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_31_mag_0.Q1.t2 VSS.t96 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X186 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VDD.t241 VDD.t240 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X187 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_19493_1349# VSS.t255 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X188 a_20211_252# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t189 VSS.t188 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X189 VSS CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_1080_4227# VSS.t93 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X190 a_1644_4227# CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t291 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X191 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_2.QB VDD.t359 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X192 a_2269_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t218 VSS.t217 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X193 a_7089_360# VDD.t479 VSS.t36 VSS.t35 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X194 a_6029_405# CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t230 VSS.t229 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X195 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t346 VDD.t345 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X196 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VDD.t219 VDD.t218 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X197 VSS CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_4864_4226# VSS.t143 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X198 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t354 VDD.t353 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X199 VDD CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VDD.t205 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X200 a_2368_4227# CLK_div_31_mag_0.Q1.t8 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t10 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X201 a_1080_4227# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t223 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X202 VDD CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VDD.t115 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X203 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_18929_1349# VSS.t240 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X204 a_19493_1349# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t228 VSS.t227 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X205 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK.t4 a_10368_3965# VSS.t70 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X206 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t214 VSS.t213 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X207 RST CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN VSS.t15 VSS.t14 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X208 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t465 VDD.t464 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X209 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.Q3.t6 VDD.t86 VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X210 a_18359_208# CLK_div_3_mag_0.CLK a_18199_208# VSS.t206 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X211 VSS CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_516_4227# VSS.t237 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X212 a_4864_4226# RST.t11 a_4704_4226# VSS.t137 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X213 a_8452_3208# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS.t148 VSS.t79 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X214 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_4.QB VDD.t162 VDD.t161 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X215 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q1.t9 a_7507_3970# VSS.t11 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X216 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t173 VDD.t172 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X217 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_19083_208# VSS.t226 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X218 a_4747_1502# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t136 VSS.t135 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X219 a_10368_3965# CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS.t248 VSS.t70 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X220 a_19614_2684# CLK_div_3_mag_0.or_2_mag_0.IN2 VDD.t148 VDD.t147 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X221 VDD CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t454 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X222 a_15912_1349# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t140 VSS.t139 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X223 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X224 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VSS.t253 VSS.t252 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X225 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 VDD.t304 VDD.t303 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X226 a_7813_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VSS.t110 VSS.t109 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X227 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VDD.t155 VDD.t154 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X228 a_5311_1502# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t155 VSS.t154 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X229 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X230 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_15912_1349# VSS.t159 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X231 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t302 VDD.t301 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X232 VDD CLK_div_3_mag_0.CLK CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t319 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X233 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t201 VDD.t200 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X234 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VDD.t286 VDD.t285 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X235 VDD CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD.t265 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X236 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_4.QB a_7255_1457# VSS.t97 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X237 VSS CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VSS.t18 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X238 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t62 VDD.t64 VDD.t63 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X239 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.QB VDD.t9 VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X240 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t470 VDD.t469 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X241 VDD VDD.t58 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t59 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X242 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t55 VDD.t57 VDD.t56 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X243 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_16630_252# VSS.t69 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X244 CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t60 VSS.t59 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X245 VDD CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD.t398 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X246 VDD CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t466 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X247 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t338 VDD.t337 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X248 a_7249_360# CLK_div_31_mag_0.Q3.t7 a_7089_360# VSS.t53 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X249 VDD CLK_div_31_mag_0.Q0.t12 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD.t421 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X250 VDD CLK_div_31_mag_0.Q3.t8 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X251 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VDD.t402 VDD.t401 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X252 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.Q3.t9 a_6029_405# VSS.t54 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X253 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t215 VDD.t214 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X254 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X255 VDD CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VDD.t295 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X256 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 a_20057_1349# VSS.t265 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X257 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.Q2 a_2987_396# VSS.t75 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X258 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK.t5 VDD.t112 VDD.t111 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X259 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 a_18359_208# VSS.t197 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X260 VDD RST.t12 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VDD.t222 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X261 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD.t102 VDD.t101 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X262 a_18641_2448# CLK_div_3_mag_0.CLK VSS.t205 VSS.t204 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X263 CLK_div_3_mag_0.CLK CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t179 VSS.t178 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X264 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t256 VDD.t255 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X265 VDD CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_3.QB VDD.t192 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X266 VDD VDD.t51 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD.t52 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X267 VSS CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VSS.t190 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X268 a_9403_3219# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS.t277 VSS.t52 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X269 a_15348_1305# CLK_div_3_mag_0.CLK a_15188_1305# VSS.t203 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X270 a_20057_1349# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t225 VSS.t224 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X271 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VSS.t216 VSS.t215 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X272 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_8537_404# VSS.t125 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X273 a_975_352# VDD.t482 VSS.t34 VSS.t33 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X274 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_0.QB.t4 a_1141_1449# VSS.t296 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X275 CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.Q0.t13 VDD.t420 VDD.t419 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X276 a_5422_3129# CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t2 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X277 VDD CLK_div_31_mag_0.Q1.t10 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t21 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X278 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t436 VDD.t435 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X279 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.Q4.t8 VDD.t411 VDD.t410 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X280 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK.t6 VDD.t114 VDD.t113 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X281 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VDD.t275 VDD.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X282 VDD CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD.t211 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X283 a_15188_1305# CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS.t267 VSS.t266 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X284 VSS CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_3576_4226# VSS.t116 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X285 VDD CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD.t395 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X286 Vdiv93 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t279 VDD.t278 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X287 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X288 a_2987_396# CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t104 VSS.t103 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X289 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VDD.t234 VDD.t233 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X290 VSS VDD.t483 a_5588_4226# VSS.t30 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X291 CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_31_mag_0.Q1.t11 VDD.t196 VDD.t195 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X292 VSS CLK_div_31_mag_0.Q0.t14 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS.t280 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X293 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VDD.t416 VDD.t415 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X294 VDD CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t141 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X295 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t48 VDD.t50 VDD.t49 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X296 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS.t290 VSS.t289 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X297 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t391 VDD.t390 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X298 VDD CLK_div_31_mag_0.Q3.t10 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t374 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X299 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q1.t12 a_10367_3208# VSS.t119 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X300 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_7819_1501# VSS.t72 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X301 a_3576_4226# CLK_div_31_mag_0.Q0.t15 CLK_div_31_mag_0.JK_FF_mag_3.QB VSS.t279 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X302 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD.t248 VDD.t247 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X303 a_5588_4226# CLK.t7 a_5428_4226# VSS.t71 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X304 VSS CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VSS.t4 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X305 VSS CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_4140_4226# VSS.t127 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X306 VDD CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VDD.t202 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X307 VDD CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t125 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X308 a_516_4227# CLK_div_31_mag_0.Q1.t13 CLK_div_31_mag_0.JK_FF_mag_2.QB VSS.t120 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X309 a_4704_4226# CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t261 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X310 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t303 VSS.t302 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X311 Vdiv93 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t172 VSS.t171 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X312 VDD CLK_div_31_mag_0.Q3.t11 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD.t377 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X313 a_7507_3970# CLK_div_31_mag_0.Q0.t16 VSS.t278 VSS.t11 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X314 a_10367_3208# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS.t276 VSS.t119 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X315 a_4741_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t232 VSS.t231 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X316 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD.t369 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X317 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_16476_1349# VSS.t68 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X318 a_17040_1349# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t124 VSS.t123 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X319 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t277 VDD.t276 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X320 CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VDD.t358 VDD.t357 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X321 a_5465_405# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t194 VSS.t193 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X322 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t174 VSS.t173 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X323 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VDD.t153 VDD.t152 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X324 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD.t45 VDD.t47 VDD.t46 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X325 a_2423_396# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t306 VSS.t305 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X326 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_1705_1493# VSS.t304 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X327 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_19647_252# VSS.t254 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X328 a_15182_208# VDD.t484 VSS.t29 VSS.t28 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X329 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.Q3.t12 VSS.t250 VSS.t249 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X330 a_16476_1349# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t221 VSS.t220 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X331 VDD CLK_div_31_mag_0.Q1.t14 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t197 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X332 a_1699_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t257 VSS.t256 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X333 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VDD.t36 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X334 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB a_17040_1349# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X335 VSS CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_1804_4227# VSS.t245 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X336 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0 a_20211_252# VSS.t196 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X337 VDD CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t122 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X338 a_17194_252# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t132 VSS.t131 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X339 a_7255_1457# CLK_div_31_mag_0.Q3.t13 a_7095_1457# VSS.t251 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X340 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t178 VDD.t177 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X341 VDD CLK_div_31_mag_0.JK_FF_mag_0.QB.t5 CLK_div_31_mag_0.Q2 VDD.t449 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X342 VDD RST.t13 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t225 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X343 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t363 VDD.t362 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X344 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_0.QB.t6 VDD.t453 VDD.t452 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X345 VSS CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VSS.t21 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X346 a_15906_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t170 VSS.t169 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X347 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_7973_360# VSS.t90 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X348 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t310 VDD.t309 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X349 VDD CLK_div_3_mag_0.CLK CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t316 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X350 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VDD.t418 VDD.t417 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X351 a_7095_1457# VDD.t485 VSS.t27 VSS.t26 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X352 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK VDD.t315 VDD.t314 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X353 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t294 VDD.t293 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X354 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q3.t14 a_8453_3965# VSS.t233 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X355 VDD CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD.t5 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X356 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VDD.t290 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X357 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VDD.t404 VDD.t403 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X358 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VDD.t96 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X359 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VDD.t383 VDD.t382 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X360 a_1135_352# CLK_div_31_mag_0.Q1.t15 a_975_352# VSS.t121 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X361 VDD CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t298 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X362 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_31_mag_0.Q3.t15 VDD.t381 VDD.t380 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X363 a_4017_361# VDD.t486 VSS.t25 VSS.t24 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X364 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.Q2 VDD.t121 VDD.t120 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X365 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VSS.t244 VSS.t243 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X366 a_9101_404# CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VSS.t142 VSS.t141 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X367 CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_31_mag_0.Q4.t9 VSS.t271 VSS.t270 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X368 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t42 VDD.t44 VDD.t43 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X369 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t39 VDD.t41 VDD.t40 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X370 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.QB VDD.t28 VDD.t27 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X371 VDD CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.Q3 VDD.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X372 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5465_405# VSS.t85 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X373 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t295 VSS.t294 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X374 VDD CLK_div_3_mag_0.CLK CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t311 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X375 a_7973_360# RST.t14 a_7813_360# VSS.t138 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X376 a_1141_1449# CLK_div_31_mag_0.Q1.t16 a_981_1449# VSS.t122 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X377 VSS CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS.t185 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X378 VSS CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VSS.t61 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X379 VDD RST.t15 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t228 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 CLK_div_31_mag_0.Q0.n14 CLK_div_31_mag_0.Q0.t8 36.935
R1 CLK_div_31_mag_0.Q0.n9 CLK_div_31_mag_0.Q0.t11 36.935
R2 CLK_div_31_mag_0.Q0.n20 CLK_div_31_mag_0.Q0.t4 36.935
R3 CLK_div_31_mag_0.Q0.n26 CLK_div_31_mag_0.Q0.t15 31.4332
R4 CLK_div_31_mag_0.Q0.n23 CLK_div_31_mag_0.Q0.t7 30.9379
R5 CLK_div_31_mag_0.Q0.n22 CLK_div_31_mag_0.Q0.t6 30.9379
R6 CLK_div_31_mag_0.Q0.n6 CLK_div_31_mag_0.Q0.t12 25.4744
R7 CLK_div_31_mag_0.Q0.n23 CLK_div_31_mag_0.Q0.t10 21.6422
R8 CLK_div_31_mag_0.Q0.n22 CLK_div_31_mag_0.Q0.t16 21.6422
R9 CLK_div_31_mag_0.Q0.n14 CLK_div_31_mag_0.Q0.t5 18.1962
R10 CLK_div_31_mag_0.Q0.n9 CLK_div_31_mag_0.Q0.t9 18.1962
R11 CLK_div_31_mag_0.Q0.n20 CLK_div_31_mag_0.Q0.t3 18.1962
R12 CLK_div_31_mag_0.Q0.n26 CLK_div_31_mag_0.Q0.t13 15.3826
R13 CLK_div_31_mag_0.Q0.n6 CLK_div_31_mag_0.Q0.t14 14.1417
R14 CLK_div_31_mag_0.Q0.n4 CLK_div_31_mag_0.Q0.t0 7.09905
R15 CLK_div_31_mag_0.Q0.n27 CLK_div_31_mag_0.Q0.n26 6.86029
R16 CLK_div_31_mag_0.Q0.n24 CLK_div_31_mag_0.Q0 6.54296
R17 CLK_div_31_mag_0.Q0.n25 CLK_div_31_mag_0.Q0.n24 4.54543
R18 CLK_div_31_mag_0.Q0.n1 CLK_div_31_mag_0.Q0.n0 1.50092
R19 CLK_div_31_mag_0.Q0.n11 CLK_div_31_mag_0.Q0.n8 4.5005
R20 CLK_div_31_mag_0.Q0.n13 CLK_div_31_mag_0.Q0.n12 4.5005
R21 CLK_div_31_mag_0.Q0.n17 CLK_div_31_mag_0.Q0.n15 4.5005
R22 CLK_div_31_mag_0.Q0.n17 CLK_div_31_mag_0.Q0.n16 4.5005
R23 CLK_div_31_mag_0.Q0.n19 CLK_div_31_mag_0.Q0.n5 4.5005
R24 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q0.n23 4.11094
R25 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q0.n22 4.11094
R26 CLK_div_31_mag_0.Q0.n28 CLK_div_31_mag_0.Q0.n25 3.5302
R27 CLK_div_31_mag_0.Q0.n4 CLK_div_31_mag_0.Q0.n3 3.25053
R28 CLK_div_31_mag_0.Q0.n3 CLK_div_31_mag_0.Q0.t2 2.2755
R29 CLK_div_31_mag_0.Q0.n3 CLK_div_31_mag_0.Q0.n2 2.2755
R30 CLK_div_31_mag_0.Q0.n29 CLK_div_31_mag_0.Q0 2.25167
R31 CLK_div_31_mag_0.Q0.n18 CLK_div_31_mag_0.Q0.n7 2.25107
R32 CLK_div_31_mag_0.Q0.n21 CLK_div_31_mag_0.Q0.n20 2.13459
R33 CLK_div_31_mag_0.Q0.n10 CLK_div_31_mag_0.Q0.n9 2.12444
R34 CLK_div_31_mag_0.Q0.n15 CLK_div_31_mag_0.Q0.n14 2.12188
R35 CLK_div_31_mag_0.Q0.n17 CLK_div_31_mag_0.Q0.n13 1.71671
R36 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q0.n28 1.52539
R37 CLK_div_31_mag_0.Q0.n10 CLK_div_31_mag_0.Q0.n8 1.50503
R38 CLK_div_31_mag_0.Q0.n25 CLK_div_31_mag_0.Q0.n21 1.37844
R39 CLK_div_31_mag_0.Q0.n28 CLK_div_31_mag_0.Q0.n27 1.12067
R40 CLK_div_31_mag_0.Q0.n0 CLK_div_31_mag_0.Q0.n18 0.932217
R41 CLK_div_31_mag_0.Q0.n24 CLK_div_31_mag_0.Q0 0.485557
R42 CLK_div_31_mag_0.Q0.n5 CLK_div_31_mag_0.Q0 0.1705
R43 CLK_div_31_mag_0.Q0.n29 CLK_div_31_mag_0.Q0.n4 0.0905
R44 CLK_div_31_mag_0.Q0.n27 CLK_div_31_mag_0.Q0 0.0857632
R45 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q0.n29 0.0834687
R46 CLK_div_31_mag_0.Q0.n21 CLK_div_31_mag_0.Q0 0.0800273
R47 CLK_div_31_mag_0.Q0.n16 CLK_div_31_mag_0.Q0 0.0457995
R48 CLK_div_31_mag_0.Q0.n11 CLK_div_31_mag_0.Q0 0.0457995
R49 CLK_div_31_mag_0.Q0.n13 CLK_div_31_mag_0.Q0.n8 0.0386356
R50 CLK_div_31_mag_0.Q0.n16 CLK_div_31_mag_0.Q0.n7 0.0377414
R51 CLK_div_31_mag_0.Q0.n12 CLK_div_31_mag_0.Q0.n11 0.0377414
R52 CLK_div_31_mag_0.Q0.n19 CLK_div_31_mag_0.Q0.n0 0.0322517
R53 CLK_div_31_mag_0.Q0.n5 CLK_div_31_mag_0.Q0.n1 0.0326665
R54 CLK_div_31_mag_0.Q0.n18 CLK_div_31_mag_0.Q0.n17 0.0122182
R55 CLK_div_31_mag_0.Q0.n15 CLK_div_31_mag_0.Q0.n7 0.00360345
R56 CLK_div_31_mag_0.Q0.n12 CLK_div_31_mag_0.Q0.n10 0.00203726
R57 CLK_div_31_mag_0.Q0.n1 CLK_div_31_mag_0.Q0.n6 1.42251
R58 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q0.n19 0.338856
R59 VDD.n141 VDD.t355 13882.6
R60 VDD.n188 VDD.t240 13882.6
R61 VDD.n138 VDD.t437 12382.6
R62 VDD.n176 VDD.t417 12382.6
R63 VDD.n293 VDD.n292 11185.2
R64 VDD.n134 VDD.t372 7208.33
R65 VDD.n165 VDD.t415 7041.67
R66 VDD.t268 VDD.t253 961.905
R67 VDD.t452 VDD.t309 961.905
R68 VDD.t435 VDD.n161 848.615
R69 VDD.t21 VDD.n162 809.492
R70 VDD.t345 VDD.t387 765.152
R71 VDD.t364 VDD.t349 765.152
R72 VDD.t92 VDD.t403 765.152
R73 VDD.t384 VDD.t293 765.152
R74 VDD.t347 VDD.t362 765.152
R75 VDD.t303 VDD.t31 765.152
R76 VDD.t108 VDD.t216 765.152
R77 VDD.t339 VDD.t255 765.152
R78 VDD.t457 VDD.t276 765.152
R79 VDD.t205 VDD.t233 765.152
R80 VDD.t154 VDD.t118 765.152
R81 VDD.t410 VDD.t179 765.152
R82 VDD.t242 VDD.t202 765.152
R83 VDD.t152 VDD.t115 765.152
R84 VDD.t247 VDD.t161 765.152
R85 VDD.t144 VDD.t139 765.152
R86 VDD.t298 VDD.t249 765.152
R87 VDD.t27 VDD.t220 765.152
R88 VDD.t265 VDD.t5 765.152
R89 VDD.t398 VDD.t214 765.152
R90 VDD.t392 VDD.t101 765.152
R91 VDD.t235 VDD.t432 765.152
R92 VDD.t395 VDD.t211 765.152
R93 VDD.t192 VDD.t103 765.152
R94 VDD.t181 VDD.t262 765.152
R95 VDD.t444 VDD.t159 765.152
R96 VDD.t174 VDD.t343 765.152
R97 VDD.t369 VDD.t18 765.152
R98 VDD.t441 VDD.t156 765.152
R99 VDD.t359 VDD.t341 765.152
R100 VDD.t271 VDD.t172 765.152
R101 VDD.t333 VDD.t469 765.152
R102 VDD.t131 VDD.t390 765.152
R103 VDD.t141 VDD.t351 765.152
R104 VDD.t251 VDD.t301 765.152
R105 VDD.t380 VDD.t353 765.152
R106 VDD.n292 VDD.t335 676.191
R107 VDD.t290 VDD.t274 536.798
R108 VDD.t357 VDD.t412 501.002
R109 VDD.t382 VDD.t96 501.002
R110 VDD.t331 VDD.t10 501.002
R111 VDD.n125 VDD.t401 485.714
R112 VDD.n293 VDD.t66 485.714
R113 VDD VDD.n141 451.327
R114 VDD.n188 VDD 448.709
R115 VDD VDD.n138 445.577
R116 VDD.n176 VDD 442.993
R117 VDD VDD.n134 431.3
R118 VDD VDD.n68 429.187
R119 VDD VDD.n243 429.187
R120 VDD.n408 VDD 429.187
R121 VDD VDD.n165 428.8
R122 VDD.n50 VDD 427.092
R123 VDD.n502 VDD 427.092
R124 VDD VDD.n222 426.699
R125 VDD VDD.n271 426.699
R126 VDD.t327 VDD.n125 426.44
R127 VDD.t16 VDD.n293 426.44
R128 VDD VDD.n130 425.019
R129 VDD VDD.n52 420.935
R130 VDD.n68 VDD.t459 386.365
R131 VDD.t46 VDD.n408 386.365
R132 VDD.n243 VDD.t43 386.365
R133 VDD.t59 VDD.n222 386.365
R134 VDD.t76 VDD.n271 386.365
R135 VDD.t319 VDD.t3 380.952
R136 VDD.t13 VDD.t452 380.952
R137 VDD.t169 VDD.n130 378.788
R138 VDD.t122 VDD.n134 378.788
R139 VDD.t374 VDD.n138 378.788
R140 VDD.t208 VDD.n141 378.788
R141 VDD.t87 VDD.n165 378.788
R142 VDD.t133 VDD.n176 378.788
R143 VDD.t244 VDD.n188 378.788
R144 VDD.n450 VDD.t33 362.8
R145 VDD.n452 VDD.t218 362.8
R146 VDD.n454 VDD.t36 359.49
R147 VDD.n422 VDD.t285 359.49
R148 VDD.n52 VDD.t147 322.223
R149 VDD.t308 VDD.n50 320.635
R150 VDD.t282 VDD.n502 309.341
R151 VDD.t403 VDD.t311 303.031
R152 VDD.t187 VDD.t347 303.031
R153 VDD.t324 VDD.t303 303.031
R154 VDD.t228 VDD.t339 303.031
R155 VDD.t316 VDD.t457 303.031
R156 VDD.t222 VDD.t154 303.031
R157 VDD.t79 VDD.t410 303.031
R158 VDD.t161 VDD.t377 303.031
R159 VDD.t136 VDD.t27 303.031
R160 VDD.t5 VDD.t111 303.031
R161 VDD.t432 VDD.t113 303.031
R162 VDD.t190 VDD.t395 303.031
R163 VDD.t262 VDD.t430 303.031
R164 VDD.t18 VDD.t424 303.031
R165 VDD.t90 VDD.t441 303.031
R166 VDD.t184 VDD.t333 303.031
R167 VDD.t197 VDD.t131 303.031
R168 VDD.t225 VDD.t251 303.031
R169 VDD.t125 VDD.t380 303.031
R170 VDD.n423 VDD.t287 296.538
R171 VDD.t257 VDD.n118 285.714
R172 VDD.n292 VDD.t466 285.714
R173 VDD.n104 VDD.t0 242.857
R174 VDD.n113 VDD.t105 242.857
R175 VDD.n119 VDD.t257 242.857
R176 VDD.n124 VDD.t319 242.857
R177 VDD.n274 VDD.t449 242.857
R178 VDD.n280 VDD.t268 242.857
R179 VDD.t466 VDD.n284 242.857
R180 VDD.n289 VDD.t13 242.857
R181 VDD.t367 VDD.n424 227.456
R182 VDD.n59 VDD.t461 193.183
R183 VDD.n36 VDD.t149 193.183
R184 VDD.n42 VDD.t387 193.183
R185 VDD.n43 VDD.t364 193.183
R186 VDD.n67 VDD.t311 193.183
R187 VDD.n15 VDD.t305 193.183
R188 VDD.n17 VDD.t384 193.183
R189 VDD.n20 VDD.t187 193.183
R190 VDD.n23 VDD.t324 193.183
R191 VDD.n71 VDD.t454 193.183
R192 VDD.n73 VDD.t108 193.183
R193 VDD.n76 VDD.t228 193.183
R194 VDD.n79 VDD.t316 193.183
R195 VDD.n132 VDD.t169 193.183
R196 VDD.n136 VDD.t122 193.183
R197 VDD.n140 VDD.t374 193.183
R198 VDD.n143 VDD.t208 193.183
R199 VDD.n463 VDD.t407 193.183
R200 VDD.n465 VDD.t205 193.183
R201 VDD.n468 VDD.t222 193.183
R202 VDD.n471 VDD.t79 193.183
R203 VDD.n164 VDD.t21 193.183
R204 VDD.n167 VDD.t87 193.183
R205 VDD.n182 VDD.t133 193.183
R206 VDD.n189 VDD.t244 193.183
R207 VDD.n412 VDD.t163 193.183
R208 VDD.t202 VDD.n411 193.183
R209 VDD.t115 VDD.n410 193.183
R210 VDD.t377 VDD.n409 193.183
R211 VDD.n225 VDD.t24 193.183
R212 VDD.n231 VDD.t144 193.183
R213 VDD.n235 VDD.t298 193.183
R214 VDD.n240 VDD.t136 193.183
R215 VDD.n245 VDD.t128 193.183
R216 VDD.n247 VDD.t271 193.183
R217 VDD.n250 VDD.t184 193.183
R218 VDD.n253 VDD.t197 193.183
R219 VDD.n196 VDD.t82 193.183
R220 VDD.n198 VDD.t141 193.183
R221 VDD.n201 VDD.t225 193.183
R222 VDD.n204 VDD.t125 193.183
R223 VDD.t111 VDD.n227 191.288
R224 VDD.t214 VDD.n234 191.288
R225 VDD.t101 VDD.n237 191.288
R226 VDD.n242 VDD.t8 191.288
R227 VDD.t113 VDD.n366 191.288
R228 VDD.n367 VDD.t190 191.288
R229 VDD.t103 VDD.n375 191.288
R230 VDD.n376 VDD.t419 191.288
R231 VDD.t430 VDD.n276 191.288
R232 VDD.t159 VDD.n283 191.288
R233 VDD.t343 VDD.n286 191.288
R234 VDD.n291 VDD.t260 191.288
R235 VDD.t424 VDD.n310 191.288
R236 VDD.n311 VDD.t90 191.288
R237 VDD.t341 VDD.n319 191.288
R238 VDD.n320 VDD.t195 191.288
R239 VDD.n450 VDD.n424 167.588
R240 VDD.n51 VDD.t308 142.857
R241 VDD.n104 VDD.t200 138.095
R242 VDD.n113 VDD.t337 138.095
R243 VDD.n119 VDD.t231 138.095
R244 VDD.t401 VDD.n124 138.095
R245 VDD.t253 VDD.n274 138.095
R246 VDD.t335 VDD.n280 138.095
R247 VDD.t309 VDD.n284 138.095
R248 VDD.t66 VDD.n289 138.095
R249 VDD.n503 VDD.t282 137.826
R250 VDD.n453 VDD.n452 119.706
R251 VDD.n454 VDD.n453 118.614
R252 VDD.n227 VDD.t59 111.743
R253 VDD.n234 VDD.t265 111.743
R254 VDD.n237 VDD.t398 111.743
R255 VDD.n242 VDD.t392 111.743
R256 VDD.n366 VDD.t52 111.743
R257 VDD.n367 VDD.t235 111.743
R258 VDD.n375 VDD.t211 111.743
R259 VDD.n376 VDD.t192 111.743
R260 VDD.n276 VDD.t76 111.743
R261 VDD.n283 VDD.t181 111.743
R262 VDD.n286 VDD.t444 111.743
R263 VDD.n291 VDD.t174 111.743
R264 VDD.n310 VDD.t72 111.743
R265 VDD.n311 VDD.t369 111.743
R266 VDD.n319 VDD.t156 111.743
R267 VDD.n320 VDD.t359 111.743
R268 VDD.t147 VDD.n51 111.112
R269 VDD.n59 VDD.t322 109.849
R270 VDD.n36 VDD.t345 109.849
R271 VDD.t349 VDD.n42 109.849
R272 VDD.n43 VDD.t92 109.849
R273 VDD.t459 VDD.n67 109.849
R274 VDD.t293 VDD.n15 109.849
R275 VDD.t362 VDD.n17 109.849
R276 VDD.t31 VDD.n20 109.849
R277 VDD.n23 VDD.t40 109.849
R278 VDD.t216 VDD.n71 109.849
R279 VDD.t255 VDD.n73 109.849
R280 VDD.t276 VDD.n76 109.849
R281 VDD.n79 VDD.t49 109.849
R282 VDD.t372 VDD.n132 109.849
R283 VDD.t437 VDD.n136 109.849
R284 VDD.t355 VDD.n140 109.849
R285 VDD.n143 VDD.t428 109.849
R286 VDD.t233 VDD.n463 109.849
R287 VDD.t118 VDD.n465 109.849
R288 VDD.t179 VDD.n468 109.849
R289 VDD.n471 VDD.t69 109.849
R290 VDD.t415 VDD.n164 109.849
R291 VDD.t417 VDD.n167 109.849
R292 VDD.t240 VDD.n182 109.849
R293 VDD.n189 VDD.t426 109.849
R294 VDD.n412 VDD.t242 109.849
R295 VDD.n411 VDD.t152 109.849
R296 VDD.n410 VDD.t247 109.849
R297 VDD.n409 VDD.t46 109.849
R298 VDD.t139 VDD.n225 109.849
R299 VDD.t249 VDD.n231 109.849
R300 VDD.t220 VDD.n235 109.849
R301 VDD.t43 VDD.n240 109.849
R302 VDD.t172 VDD.n245 109.849
R303 VDD.t469 VDD.n247 109.849
R304 VDD.t390 VDD.n250 109.849
R305 VDD.n253 VDD.t63 109.849
R306 VDD.t351 VDD.n196 109.849
R307 VDD.t301 VDD.n198 109.849
R308 VDD.t353 VDD.n201 109.849
R309 VDD.n204 VDD.t56 109.849
R310 VDD.n503 VDD.t405 107.198
R311 VDD.n423 VDD.n422 100.365
R312 VDD.n188 VDD.t329 65.4455
R313 VDD.n176 VDD.t280 64.6
R314 VDD.n141 VDD.t447 62.8277
R315 VDD.n165 VDD.t177 62.5005
R316 VDD.n222 VDD.t166 62.1896
R317 VDD.n271 VDD.t421 62.1896
R318 VDD.n138 VDD.t238 62.016
R319 VDD.n134 VDD.t99 60.0005
R320 VDD.n68 VDD.t314 59.702
R321 VDD.n408 VDD.t85 59.702
R322 VDD.n243 VDD.t120 59.702
R323 VDD.n50 VDD.t278 59.4064
R324 VDD.n502 VDD.t283 59.4064
R325 VDD.n130 VDD.t94 59.1138
R326 VDD.n52 VDD.t464 58.5371
R327 VDD.n453 VDD.n424 47.8826
R328 VDD.n80 VDD.t39 30.9379
R329 VDD.n474 VDD.t68 30.9379
R330 VDD.n472 VDD.t45 30.9379
R331 VDD.n356 VDD.t51 30.9379
R332 VDD.n358 VDD.t58 30.9379
R333 VDD.n300 VDD.t71 30.9379
R334 VDD.n301 VDD.t75 30.9379
R335 VDD.n254 VDD.t65 30.9379
R336 VDD.n256 VDD.t62 30.9379
R337 VDD.n205 VDD.t42 30.9379
R338 VDD.n207 VDD.t55 30.9379
R339 VDD.n85 VDD.t48 30.0062
R340 VDD.n459 VDD.t287 28.139
R341 VDD.t274 VDD.n459 28.139
R342 VDD.n460 VDD.t290 28.139
R343 VDD.n460 VDD.t439 28.139
R344 VDD.n80 VDD.t474 24.5101
R345 VDD.n474 VDD.t479 24.5101
R346 VDD.n472 VDD.t485 24.5101
R347 VDD.n356 VDD.t483 24.5101
R348 VDD.n358 VDD.t478 24.5101
R349 VDD.n300 VDD.t477 24.5101
R350 VDD.n301 VDD.t475 24.5101
R351 VDD.n254 VDD.t472 24.5101
R352 VDD.n256 VDD.t482 24.5101
R353 VDD.n205 VDD.t473 24.5101
R354 VDD.n207 VDD.t486 24.5101
R355 VDD.n84 VDD.t484 24.4392
R356 VDD.n435 VDD.t295 22.0446
R357 VDD.n436 VDD.t357 22.0446
R358 VDD.n439 VDD.t412 22.0446
R359 VDD.n440 VDD.t382 22.0446
R360 VDD.n443 VDD.t96 22.0446
R361 VDD.n444 VDD.t331 22.0446
R362 VDD.n447 VDD.t10 21.0426
R363 VDD.n448 VDD.t367 21.0426
R364 VDD.n453 VDD.n423 18.2487
R365 VDD VDD.t327 10.5649
R366 VDD VDD.t16 10.5649
R367 VDD.n432 VDD.t358 8.94586
R368 VDD.n430 VDD.t383 8.94586
R369 VDD.n428 VDD.t332 8.94586
R370 VDD.n426 VDD.t368 8.92336
R371 VDD.n82 VDD.n81 6.98838
R372 VDD.n185 VDD.t330 6.62407
R373 VDD.n54 VDD.n51 6.3005
R374 VDD.n24 VDD.n23 6.3005
R375 VDD.n27 VDD.n20 6.3005
R376 VDD.n30 VDD.n17 6.3005
R377 VDD.n33 VDD.n15 6.3005
R378 VDD.n44 VDD.n43 6.3005
R379 VDD.n42 VDD.n41 6.3005
R380 VDD.n37 VDD.n36 6.3005
R381 VDD.n60 VDD.n59 6.3005
R382 VDD.n92 VDD.n79 6.3005
R383 VDD.n95 VDD.n76 6.3005
R384 VDD.n98 VDD.n73 6.3005
R385 VDD.n101 VDD.n71 6.3005
R386 VDD.n124 VDD.n123 6.3005
R387 VDD.n120 VDD.n119 6.3005
R388 VDD.n114 VDD.n113 6.3005
R389 VDD.n105 VDD.n104 6.3005
R390 VDD.n67 VDD.n66 6.3005
R391 VDD.n144 VDD.n143 6.3005
R392 VDD.n148 VDD.n140 6.3005
R393 VDD.n153 VDD.n136 6.3005
R394 VDD.n158 VDD.n132 6.3005
R395 VDD.n435 VDD 6.3005
R396 VDD VDD.n436 6.3005
R397 VDD.n439 VDD 6.3005
R398 VDD VDD.n440 6.3005
R399 VDD.n443 VDD 6.3005
R400 VDD VDD.n444 6.3005
R401 VDD.n447 VDD 6.3005
R402 VDD VDD.n448 6.3005
R403 VDD.n452 VDD 6.3005
R404 VDD VDD.n450 6.3005
R405 VDD.n487 VDD.n463 6.3005
R406 VDD.n484 VDD.n465 6.3005
R407 VDD.n481 VDD.n468 6.3005
R408 VDD.n478 VDD.n471 6.3005
R409 VDD.n310 VDD.n309 6.3005
R410 VDD.n312 VDD.n311 6.3005
R411 VDD.n319 VDD.n318 6.3005
R412 VDD.n321 VDD.n320 6.3005
R413 VDD.n260 VDD.n253 6.3005
R414 VDD.n263 VDD.n250 6.3005
R415 VDD.n266 VDD.n247 6.3005
R416 VDD.n269 VDD.n245 6.3005
R417 VDD.n343 VDD.n276 6.3005
R418 VDD.n336 VDD.n283 6.3005
R419 VDD.n331 VDD.n286 6.3005
R420 VDD.n325 VDD.n291 6.3005
R421 VDD.n328 VDD.n289 6.3005
R422 VDD.n335 VDD.n284 6.3005
R423 VDD.n340 VDD.n280 6.3005
R424 VDD.n346 VDD.n274 6.3005
R425 VDD.n366 VDD.n365 6.3005
R426 VDD.n368 VDD.n367 6.3005
R427 VDD.n375 VDD.n374 6.3005
R428 VDD.n377 VDD.n376 6.3005
R429 VDD.n211 VDD.n204 6.3005
R430 VDD.n214 VDD.n201 6.3005
R431 VDD.n217 VDD.n198 6.3005
R432 VDD.n220 VDD.n196 6.3005
R433 VDD.n400 VDD.n227 6.3005
R434 VDD.n393 VDD.n234 6.3005
R435 VDD.n388 VDD.n237 6.3005
R436 VDD.n382 VDD.n242 6.3005
R437 VDD.n385 VDD.n240 6.3005
R438 VDD.n392 VDD.n235 6.3005
R439 VDD.n397 VDD.n231 6.3005
R440 VDD.n403 VDD.n225 6.3005
R441 VDD.n409 VDD.n193 6.3005
R442 VDD.n190 VDD.n189 6.3005
R443 VDD.n182 VDD.n181 6.3005
R444 VDD.n410 VDD.n170 6.3005
R445 VDD.n411 VDD.n169 6.3005
R446 VDD.n413 VDD.n412 6.3005
R447 VDD.n493 VDD.n167 6.3005
R448 VDD.n497 VDD.n164 6.3005
R449 VDD VDD.n161 6.3005
R450 VDD VDD.n162 6.3005
R451 VDD.n504 VDD.n503 6.3005
R452 VDD.n109 VDD.n108 6.15559
R453 VDD.n111 VDD.n110 6.1505
R454 VDD.n117 VDD.n0 6.13918
R455 VDD.n128 VDD.n127 6.13239
R456 VDD.n507 VDD.n506 6.01749
R457 VDD.n323 VDD.t17 5.85907
R458 VDD.n380 VDD.t121 5.85907
R459 VDD.n405 VDD.n223 5.85007
R460 VDD.n348 VDD.n272 5.85007
R461 VDD.n56 VDD.n55 5.50832
R462 VDD.n62 VDD.n6 5.32833
R463 VDD.n57 VDD.n56 5.32746
R464 VDD.n24 VDD.t41 5.213
R465 VDD VDD.t429 5.1878
R466 VDD.n434 VDD.n433 5.15595
R467 VDD VDD.t418 5.1508
R468 VDD.n45 VDD.t93 5.13287
R469 VDD.n11 VDD.n10 5.13287
R470 VDD.n40 VDD.t350 5.13287
R471 VDD.n39 VDD.n12 5.13287
R472 VDD.n38 VDD.t346 5.13287
R473 VDD.n35 VDD.n13 5.13287
R474 VDD.n26 VDD.t32 5.13287
R475 VDD.n29 VDD.t363 5.13287
R476 VDD.n31 VDD.n16 5.13287
R477 VDD.n32 VDD.t294 5.13287
R478 VDD.n34 VDD.n14 5.13287
R479 VDD.n94 VDD.t277 5.13287
R480 VDD.n97 VDD.t256 5.13287
R481 VDD.n99 VDD.n72 5.13287
R482 VDD.n100 VDD.t217 5.13287
R483 VDD.n102 VDD.n70 5.13287
R484 VDD.n145 VDD.n142 5.13287
R485 VDD.n147 VDD.t356 5.13287
R486 VDD.n149 VDD.n139 5.13287
R487 VDD.n152 VDD.t438 5.13287
R488 VDD.n154 VDD.n135 5.13287
R489 VDD.n157 VDD.t373 5.13287
R490 VDD.n159 VDD.n131 5.13287
R491 VDD.n477 VDD.t70 5.13287
R492 VDD.n480 VDD.t180 5.13287
R493 VDD.n483 VDD.t119 5.13287
R494 VDD.n485 VDD.n464 5.13287
R495 VDD.n486 VDD.t234 5.13287
R496 VDD.n488 VDD.n462 5.13287
R497 VDD.n414 VDD.t243 5.13287
R498 VDD.n402 VDD.n226 5.13287
R499 VDD.n395 VDD.n232 5.13287
R500 VDD.n391 VDD.t215 5.13287
R501 VDD.n389 VDD.n236 5.13287
R502 VDD.n386 VDD.t102 5.13287
R503 VDD.n384 VDD.n241 5.13287
R504 VDD.n381 VDD.t9 5.13287
R505 VDD.n345 VDD.n275 5.13287
R506 VDD.n338 VDD.n281 5.13287
R507 VDD.n334 VDD.t160 5.13287
R508 VDD.n332 VDD.n285 5.13287
R509 VDD.n329 VDD.t344 5.13287
R510 VDD.n327 VDD.n290 5.13287
R511 VDD.n324 VDD.t261 5.13287
R512 VDD.n305 VDD.n299 5.13287
R513 VDD.n298 VDD.n297 5.13287
R514 VDD.n314 VDD.n294 5.13287
R515 VDD.n317 VDD.t342 5.13287
R516 VDD.n316 VDD.n315 5.13287
R517 VDD.n322 VDD.t196 5.13287
R518 VDD.n326 VDD.t67 5.13287
R519 VDD.n333 VDD.t310 5.13287
R520 VDD.n337 VDD.n282 5.13287
R521 VDD.n339 VDD.t336 5.13287
R522 VDD.n342 VDD.n277 5.13287
R523 VDD.n344 VDD.t254 5.13287
R524 VDD.n347 VDD.n273 5.13287
R525 VDD.n259 VDD.t64 5.13287
R526 VDD.n262 VDD.t391 5.13287
R527 VDD.n265 VDD.t470 5.13287
R528 VDD.n267 VDD.n246 5.13287
R529 VDD.n268 VDD.t173 5.13287
R530 VDD.n270 VDD.n244 5.13287
R531 VDD.n361 VDD.n355 5.13287
R532 VDD.n354 VDD.n353 5.13287
R533 VDD.n370 VDD.n350 5.13287
R534 VDD.n373 VDD.t104 5.13287
R535 VDD.n372 VDD.n371 5.13287
R536 VDD.n378 VDD.t420 5.13287
R537 VDD.n383 VDD.t44 5.13287
R538 VDD.n390 VDD.t221 5.13287
R539 VDD.n394 VDD.n233 5.13287
R540 VDD.n396 VDD.t250 5.13287
R541 VDD.n399 VDD.n228 5.13287
R542 VDD.n401 VDD.t140 5.13287
R543 VDD.n404 VDD.n224 5.13287
R544 VDD.n210 VDD.t57 5.13287
R545 VDD.n213 VDD.t354 5.13287
R546 VDD.n216 VDD.t302 5.13287
R547 VDD.n218 VDD.n197 5.13287
R548 VDD.n219 VDD.t352 5.13287
R549 VDD.n221 VDD.n195 5.13287
R550 VDD.n194 VDD.t47 5.13287
R551 VDD.n174 VDD.n173 5.13287
R552 VDD.n191 VDD.t427 5.13287
R553 VDD.n175 VDD.t248 5.13287
R554 VDD.n179 VDD.n178 5.13287
R555 VDD.n183 VDD.t241 5.13287
R556 VDD.n187 VDD.n186 5.13287
R557 VDD.n184 VDD.t153 5.13287
R558 VDD.n180 VDD.n177 5.13287
R559 VDD.n494 VDD.n166 5.13287
R560 VDD.n498 VDD.n163 5.13287
R561 VDD.n496 VDD.t416 5.13287
R562 VDD VDD.t328 5.12757
R563 VDD.n61 VDD.t323 5.12339
R564 VDD.n58 VDD.n48 5.12339
R565 VDD.n126 VDD.t402 5.11708
R566 VDD.n121 VDD.t232 5.11708
R567 VDD.n116 VDD.n3 5.11708
R568 VDD.n115 VDD.t338 5.11708
R569 VDD.n112 VDD.n4 5.11708
R570 VDD.n5 VDD.t201 5.11708
R571 VDD.n106 VDD.n103 5.11708
R572 VDD.n7 VDD.t460 5.11708
R573 VDD VDD.t281 5.10366
R574 VDD VDD.t279 5.10321
R575 VDD.n446 VDD.n427 5.09836
R576 VDD.n442 VDD.n429 5.09836
R577 VDD.n438 VDD.n431 5.09836
R578 VDD.n449 VDD.n425 5.09836
R579 VDD.n451 VDD.t219 5.09836
R580 VDD.n421 VDD.n420 5.09836
R581 VDD.n456 VDD.t286 5.09836
R582 VDD.n457 VDD.n419 5.09836
R583 VDD.n458 VDD.t275 5.09836
R584 VDD.n418 VDD.n417 5.09836
R585 VDD.n461 VDD.t440 5.09836
R586 VDD.n49 VDD.t465 5.09407
R587 VDD.n69 VDD.t315 5.09407
R588 VDD.n146 VDD.t448 5.09407
R589 VDD.n150 VDD.t239 5.09407
R590 VDD.n155 VDD.t100 5.09407
R591 VDD.n160 VDD.t95 5.09407
R592 VDD.n407 VDD.t86 5.09407
R593 VDD.n495 VDD.t178 5.09407
R594 VDD.n500 VDD.t30 5.09407
R595 VDD.n499 VDD.t436 5.09407
R596 VDD.n501 VDD.t284 5.09407
R597 VDD.n448 VDD.n447 5.01052
R598 VDD.n416 VDD.n415 4.97242
R599 VDD.n489 VDD.n461 4.93241
R600 VDD.n91 VDD.t50 4.8755
R601 VDD.n437 VDD.n430 4.5905
R602 VDD.n441 VDD.n428 4.5905
R603 VDD.n445 VDD.n426 4.5905
R604 VDD.n161 VDD.t29 4.26489
R605 VDD.n162 VDD.t435 4.26489
R606 VDD.n505 VDD.t406 4.12326
R607 VDD.n53 VDD.t148 4.11379
R608 VDD.n208 VDD.n207 4.08741
R609 VDD VDD.n300 4.08362
R610 VDD.n255 VDD.n254 4.07437
R611 VDD.n475 VDD.n474 4.07346
R612 VDD.n257 VDD.n256 4.06995
R613 VDD.n206 VDD.n205 4.06354
R614 VDD VDD.n356 4.0592
R615 VDD.n473 VDD.n472 4.05141
R616 VDD.n359 VDD.n358 4.04913
R617 VDD.n436 VDD.n435 4.00852
R618 VDD.n440 VDD.n439 4.00852
R619 VDD.n444 VDD.n443 4.00852
R620 VDD.n302 VDD.n301 4.0005
R621 VDD.n86 VDD.n85 3.61662
R622 VDD.n455 VDD.n454 3.1505
R623 VDD.n455 VDD.n422 3.1505
R624 VDD.n459 VDD 3.1505
R625 VDD VDD.n460 3.1505
R626 VDD.n258 VDD.n255 3.06712
R627 VDD.n209 VDD.n206 3.0645
R628 VDD.n360 VDD.n359 3.00562
R629 VDD.n476 VDD.n473 2.95066
R630 VDD.n209 VDD.n208 2.92128
R631 VDD.n304 VDD.n303 2.91332
R632 VDD.n46 VDD.n9 2.85787
R633 VDD.n25 VDD.n22 2.85787
R634 VDD.n28 VDD.n19 2.85787
R635 VDD.n93 VDD.n78 2.85787
R636 VDD.n96 VDD.n75 2.85787
R637 VDD.n479 VDD.n470 2.85787
R638 VDD.n482 VDD.n467 2.85787
R639 VDD.n398 VDD.n230 2.85787
R640 VDD.n341 VDD.n279 2.85787
R641 VDD.n308 VDD.n307 2.85787
R642 VDD.n313 VDD.n296 2.85787
R643 VDD.n330 VDD.n288 2.85787
R644 VDD.n261 VDD.n252 2.85787
R645 VDD.n264 VDD.n249 2.85787
R646 VDD.n364 VDD.n363 2.85787
R647 VDD.n369 VDD.n352 2.85787
R648 VDD.n387 VDD.n239 2.85787
R649 VDD.n212 VDD.n203 2.85787
R650 VDD.n215 VDD.n200 2.85787
R651 VDD.n192 VDD.n172 2.85787
R652 VDD.n258 VDD.n257 2.85553
R653 VDD.n122 VDD.n2 2.84208
R654 VDD.n304 VDD 2.82101
R655 VDD.n360 VDD.n357 2.8124
R656 VDD.n476 VDD.n475 2.79396
R657 VDD.n9 VDD.t404 2.2755
R658 VDD.n9 VDD.n8 2.2755
R659 VDD.n22 VDD.t304 2.2755
R660 VDD.n22 VDD.n21 2.2755
R661 VDD.n19 VDD.t348 2.2755
R662 VDD.n19 VDD.n18 2.2755
R663 VDD.n2 VDD.t4 2.2755
R664 VDD.n2 VDD.n1 2.2755
R665 VDD.n78 VDD.t458 2.2755
R666 VDD.n78 VDD.n77 2.2755
R667 VDD.n75 VDD.t340 2.2755
R668 VDD.n75 VDD.n74 2.2755
R669 VDD.n470 VDD.t411 2.2755
R670 VDD.n470 VDD.n469 2.2755
R671 VDD.n467 VDD.t155 2.2755
R672 VDD.n467 VDD.n466 2.2755
R673 VDD.n230 VDD.t112 2.2755
R674 VDD.n230 VDD.n229 2.2755
R675 VDD.n279 VDD.t431 2.2755
R676 VDD.n279 VDD.n278 2.2755
R677 VDD.n307 VDD.t425 2.2755
R678 VDD.n307 VDD.n306 2.2755
R679 VDD.n296 VDD.t91 2.2755
R680 VDD.n296 VDD.n295 2.2755
R681 VDD.n288 VDD.t453 2.2755
R682 VDD.n288 VDD.n287 2.2755
R683 VDD.n252 VDD.t132 2.2755
R684 VDD.n252 VDD.n251 2.2755
R685 VDD.n249 VDD.t334 2.2755
R686 VDD.n249 VDD.n248 2.2755
R687 VDD.n363 VDD.t114 2.2755
R688 VDD.n363 VDD.n362 2.2755
R689 VDD.n352 VDD.t191 2.2755
R690 VDD.n352 VDD.n351 2.2755
R691 VDD.n239 VDD.t28 2.2755
R692 VDD.n239 VDD.n238 2.2755
R693 VDD.n203 VDD.t381 2.2755
R694 VDD.n203 VDD.n202 2.2755
R695 VDD.n200 VDD.t252 2.2755
R696 VDD.n200 VDD.n199 2.2755
R697 VDD.n172 VDD.t162 2.2755
R698 VDD.n172 VDD.n171 2.2755
R699 VDD.n361 VDD.n360 2.27547
R700 VDD.n305 VDD.n304 2.27315
R701 VDD.n210 VDD.n209 2.26966
R702 VDD.n259 VDD.n258 2.26502
R703 VDD.n477 VDD.n476 2.26153
R704 VDD.n81 VDD.n80 2.11318
R705 VDD VDD.n455 1.5755
R706 VDD.n83 VDD.n82 1.54785
R707 VDD.n506 VDD 1.37899
R708 VDD VDD.n322 1.21661
R709 VDD.n349 VDD.n270 1.18347
R710 VDD.n35 VDD.n34 1.16167
R711 VDD.n406 VDD.n221 1.12775
R712 VDD.n379 VDD.n378 1.12407
R713 VDD.n129 VDD.n128 1.06492
R714 VDD.n107 VDD.n102 1.01882
R715 VDD.n490 VDD.n489 0.986314
R716 VDD.n85 VDD.n84 0.840632
R717 VDD.n65 VDD.n64 0.7205
R718 VDD.n490 VDD.n416 0.559447
R719 VDD.n64 VDD.n47 0.487926
R720 VDD.n504 VDD.n501 0.388218
R721 VDD.n133 VDD.n129 0.341963
R722 VDD.n92 VDD.n91 0.337997
R723 VDD.n91 VDD.n90 0.328132
R724 VDD.n416 VDD.n414 0.279974
R725 VDD.n109 VDD.n6 0.247933
R726 VDD.n137 VDD.n133 0.247664
R727 VDD.n29 VDD.n28 0.233919
R728 VDD.n26 VDD.n25 0.233919
R729 VDD.n97 VDD.n96 0.233919
R730 VDD.n94 VDD.n93 0.233919
R731 VDD.n483 VDD.n482 0.233919
R732 VDD.n480 VDD.n479 0.233919
R733 VDD.n308 VDD.n298 0.233919
R734 VDD.n314 VDD.n313 0.233919
R735 VDD.n265 VDD.n264 0.233919
R736 VDD.n262 VDD.n261 0.233919
R737 VDD.n364 VDD.n354 0.233919
R738 VDD.n370 VDD.n369 0.233919
R739 VDD.n216 VDD.n215 0.233919
R740 VDD.n213 VDD.n212 0.233919
R741 VDD.n128 VDD.n0 0.224828
R742 VDD.n63 VDD.n62 0.215786
R743 VDD.n137 VDD 0.213007
R744 VDD.n110 VDD.n0 0.205754
R745 VDD.n110 VDD.n109 0.193664
R746 VDD.n379 VDD.n349 0.178068
R747 VDD.n56 VDD.n6 0.16653
R748 VDD.n53 VDD 0.162783
R749 VDD.n407 VDD.n406 0.162742
R750 VDD.n55 VDD 0.155173
R751 VDD.n63 VDD 0.150503
R752 VDD.n437 VDD 0.143635
R753 VDD.n441 VDD 0.143635
R754 VDD.n445 VDD 0.143635
R755 VDD.n32 VDD.n31 0.141016
R756 VDD.n39 VDD.n38 0.141016
R757 VDD.n40 VDD.n11 0.141016
R758 VDD.n100 VDD.n99 0.141016
R759 VDD.n486 VDD.n485 0.141016
R760 VDD.n317 VDD.n316 0.141016
R761 VDD.n268 VDD.n267 0.141016
R762 VDD.n373 VDD.n372 0.141016
R763 VDD.n219 VDD.n218 0.141016
R764 VDD VDD.n7 0.13207
R765 VDD.n126 VDD 0.13207
R766 VDD.n496 VDD 0.126036
R767 VDD.n500 VDD 0.125632
R768 VDD VDD.n45 0.122435
R769 VDD VDD.n302 0.121547
R770 VDD.n157 VDD.n156 0.121517
R771 VDD.n64 VDD.n63 0.120236
R772 VDD.n506 VDD.n505 0.119239
R773 VDD.n147 VDD 0.11887
R774 VDD VDD.n129 0.112318
R775 VDD.n46 VDD 0.111984
R776 VDD.n505 VDD 0.110164
R777 VDD.n34 VDD.n33 0.107339
R778 VDD.n31 VDD.n30 0.107339
R779 VDD.n37 VDD.n35 0.107339
R780 VDD.n41 VDD.n39 0.107339
R781 VDD.n44 VDD.n11 0.107339
R782 VDD.n102 VDD.n101 0.107339
R783 VDD.n99 VDD.n98 0.107339
R784 VDD.n488 VDD.n487 0.107339
R785 VDD.n485 VDD.n484 0.107339
R786 VDD.n318 VDD.n317 0.107339
R787 VDD.n322 VDD.n321 0.107339
R788 VDD.n270 VDD.n269 0.107339
R789 VDD.n267 VDD.n266 0.107339
R790 VDD.n374 VDD.n373 0.107339
R791 VDD.n378 VDD.n377 0.107339
R792 VDD.n221 VDD.n220 0.107339
R793 VDD.n218 VDD.n217 0.107339
R794 VDD.n81 VDD 0.106795
R795 VDD VDD.n308 0.106758
R796 VDD.n313 VDD 0.106758
R797 VDD VDD.n364 0.106758
R798 VDD.n369 VDD 0.106758
R799 VDD.n28 VDD 0.106177
R800 VDD.n25 VDD 0.106177
R801 VDD.n96 VDD 0.106177
R802 VDD.n93 VDD 0.106177
R803 VDD.n482 VDD 0.106177
R804 VDD.n479 VDD 0.106177
R805 VDD.n264 VDD 0.106177
R806 VDD.n261 VDD 0.106177
R807 VDD.n215 VDD 0.106177
R808 VDD.n212 VDD 0.106177
R809 VDD.n152 VDD.n151 0.105286
R810 VDD.n458 VDD.n418 0.102798
R811 VDD.n457 VDD.n456 0.102778
R812 VDD.n451 VDD.n421 0.0987707
R813 VDD.n146 VDD.n145 0.0984239
R814 VDD.n116 VDD.n115 0.0981682
R815 VDD.n150 VDD.n149 0.0962255
R816 VDD.n160 VDD.n159 0.0962255
R817 VDD.n499 VDD.n498 0.0962255
R818 VDD.n107 VDD.n106 0.0925179
R819 VDD.n60 VDD.n58 0.0925
R820 VDD.n155 VDD.n154 0.0917202
R821 VDD.n495 VDD.n494 0.0917202
R822 VDD.n491 VDD.n490 0.0908448
R823 VDD.n58 VDD.n57 0.0888696
R824 VDD VDD.n121 0.0852534
R825 VDD VDD.n458 0.0815938
R826 VDD VDD.n457 0.081125
R827 VDD.n507 VDD 0.0810263
R828 VDD VDD.n194 0.0808411
R829 VDD.n27 VDD.n26 0.080629
R830 VDD.n95 VDD.n94 0.080629
R831 VDD.n481 VDD.n480 0.080629
R832 VDD.n478 VDD.n477 0.080629
R833 VDD.n309 VDD.n305 0.080629
R834 VDD.n312 VDD.n298 0.080629
R835 VDD.n263 VDD.n262 0.080629
R836 VDD.n260 VDD.n259 0.080629
R837 VDD.n365 VDD.n361 0.080629
R838 VDD.n368 VDD.n354 0.080629
R839 VDD.n214 VDD.n213 0.080629
R840 VDD.n211 VDD.n210 0.080629
R841 VDD.n151 VDD.n137 0.0796304
R842 VDD.n156 VDD.n133 0.0796304
R843 VDD VDD.n32 0.0794677
R844 VDD VDD.n29 0.0794677
R845 VDD.n38 VDD 0.0794677
R846 VDD VDD.n40 0.0794677
R847 VDD.n45 VDD 0.0794677
R848 VDD VDD.n100 0.0794677
R849 VDD VDD.n97 0.0794677
R850 VDD VDD.n486 0.0794677
R851 VDD VDD.n483 0.0794677
R852 VDD VDD.n268 0.0794677
R853 VDD VDD.n265 0.0794677
R854 VDD VDD.n219 0.0794677
R855 VDD VDD.n216 0.0794677
R856 VDD VDD.n314 0.0788871
R857 VDD.n316 VDD 0.0788871
R858 VDD VDD.n370 0.0788871
R859 VDD.n372 VDD 0.0788871
R860 VDD.n145 VDD.n144 0.0782465
R861 VDD.n122 VDD 0.0779888
R862 VDD.n149 VDD.n148 0.0764633
R863 VDD.n159 VDD.n158 0.0764633
R864 VDD.n498 VDD.n497 0.0764633
R865 VDD.n108 VDD.n69 0.0759709
R866 VDD.n106 VDD.n105 0.0747601
R867 VDD.n114 VDD.n112 0.0747601
R868 VDD.n461 VDD 0.0742915
R869 VDD VDD.n122 0.0739529
R870 VDD.n456 VDD 0.0739434
R871 VDD VDD.n418 0.0738649
R872 VDD VDD.n421 0.0735189
R873 VDD.n89 VDD 0.0733571
R874 VDD VDD.n53 0.073
R875 VDD.n154 VDD.n153 0.0728144
R876 VDD.n494 VDD.n493 0.0728144
R877 VDD VDD.n501 0.0709717
R878 VDD.n47 VDD.n46 0.0669867
R879 VDD.n61 VDD 0.0655
R880 VDD.n111 VDD.n5 0.0610381
R881 VDD VDD.n451 0.0594773
R882 VDD VDD.n449 0.0591364
R883 VDD VDD.n438 0.0582099
R884 VDD VDD.n442 0.0582099
R885 VDD VDD.n446 0.0576483
R886 VDD VDD.n5 0.0553879
R887 VDD.n115 VDD 0.0553879
R888 VDD.n121 VDD 0.0553879
R889 VDD.n62 VDD.n61 0.055
R890 VDD VDD.n147 0.0541697
R891 VDD VDD.n157 0.0541697
R892 VDD VDD.n496 0.0541697
R893 VDD.n491 VDD 0.0523961
R894 VDD.n492 VDD.n491 0.0518793
R895 VDD VDD.n152 0.0515917
R896 VDD.n65 VDD.n7 0.0501413
R897 VDD VDD.n168 0.0493571
R898 VDD.n90 VDD.n89 0.0471071
R899 VDD.n127 VDD.n126 0.0452982
R900 VDD VDD.n192 0.0435288
R901 VDD.n489 VDD.n488 0.0434677
R902 VDD.n117 VDD.n116 0.0428767
R903 VDD VDD.n49 0.0410978
R904 VDD.n349 VDD 0.0403112
R905 VDD.n55 VDD.n54 0.0395
R906 VDD VDD.n379 0.0394651
R907 VDD.n406 VDD 0.0394564
R908 VDD VDD.n184 0.0392961
R909 VDD.n404 VDD.n403 0.038569
R910 VDD.n382 VDD.n381 0.038569
R911 VDD.n347 VDD.n346 0.0377135
R912 VDD.n325 VDD.n324 0.0377135
R913 VDD.n112 VDD.n111 0.03763
R914 VDD.n88 VDD.n87 0.0358571
R915 VDD.n449 VDD 0.0352326
R916 VDD.n194 VDD.n193 0.0350961
R917 VDD.n90 VDD.n88 0.03425
R918 VDD.n69 VDD 0.0339978
R919 VDD VDD.n146 0.0339978
R920 VDD VDD.n150 0.0332632
R921 VDD VDD.n160 0.0332632
R922 VDD VDD.n499 0.0332632
R923 VDD.n187 VDD.n170 0.0326553
R924 VDD.n120 VDD.n117 0.0323834
R925 VDD.n393 VDD.n392 0.0323621
R926 VDD VDD.n155 0.0317552
R927 VDD VDD.n495 0.0317552
R928 VDD.n190 VDD.n175 0.0313824
R929 VDD.n339 VDD.n338 0.0312416
R930 VDD.n333 VDD.n332 0.0312416
R931 VDD.n57 VDD.n49 0.0293587
R932 VDD.n396 VDD.n395 0.0282241
R933 VDD.n390 VDD.n389 0.0282241
R934 VDD.n336 VDD.n335 0.0280056
R935 VDD.n398 VDD.n397 0.0273966
R936 VDD.n388 VDD.n387 0.0273966
R937 VDD VDD.n399 0.0271897
R938 VDD.n386 VDD 0.0269828
R939 VDD.n344 VDD.n343 0.0267921
R940 VDD.n328 VDD.n327 0.0267921
R941 VDD VDD.n345 0.0263876
R942 VDD.n326 VDD 0.0261854
R943 VDD.n401 VDD.n400 0.0236724
R944 VDD.n385 VDD.n384 0.0236724
R945 VDD VDD.n402 0.0232586
R946 VDD.n341 VDD.n340 0.0231517
R947 VDD.n331 VDD.n330 0.0231517
R948 VDD.n383 VDD 0.0230517
R949 VDD VDD.n342 0.0229494
R950 VDD.n174 VDD 0.0228998
R951 VDD.n395 VDD.n394 0.0228448
R952 VDD.n391 VDD.n390 0.0228448
R953 VDD.n329 VDD 0.0227472
R954 VDD.n492 VDD 0.0222241
R955 VDD.n179 VDD.n168 0.0214709
R956 VDD VDD.n407 0.0207439
R957 VDD.n181 VDD.n180 0.0205971
R958 VDD.n338 VDD.n337 0.0187022
R959 VDD.n334 VDD.n333 0.0187022
R960 VDD.n191 VDD 0.0186765
R961 VDD.n359 VDD 0.0181958
R962 VDD.n151 VDD 0.0174737
R963 VDD VDD.n396 0.016431
R964 VDD.n389 VDD 0.0162241
R965 VDD.n192 VDD.n191 0.0162059
R966 VDD.n255 VDD 0.0157113
R967 VDD.n303 VDD 0.0152541
R968 VDD.n342 VDD.n341 0.0150618
R969 VDD.n330 VDD.n329 0.0150618
R970 VDD.n475 VDD 0.0133571
R971 VDD.n473 VDD 0.0132059
R972 VDD.n180 VDD.n179 0.0125583
R973 VDD.n184 VDD.n183 0.0125583
R974 VDD.n438 VDD.n437 0.0125512
R975 VDD.n442 VDD.n441 0.0125512
R976 VDD.n446 VDD.n445 0.0125094
R977 VDD VDD.n339 0.0124326
R978 VDD.n332 VDD 0.0122303
R979 VDD.n183 VDD 0.0122087
R980 VDD.n399 VDD.n398 0.0116724
R981 VDD.n387 VDD.n386 0.0116724
R982 VDD.n127 VDD.n123 0.0113969
R983 VDD VDD.n169 0.0111602
R984 VDD.n206 VDD 0.0110882
R985 VDD.n414 VDD.n413 0.0105519
R986 VDD.n257 VDD 0.00981034
R987 VDD VDD.n334 0.00980337
R988 VDD.n337 VDD 0.00960112
R989 VDD VDD.n500 0.00839474
R990 VDD.n108 VDD.n107 0.00816816
R991 VDD.n66 VDD.n65 0.00655381
R992 VDD.n405 VDD.n404 0.0065
R993 VDD VDD.n391 0.0062931
R994 VDD.n381 VDD.n380 0.0062931
R995 VDD.n394 VDD 0.00608621
R996 VDD.n402 VDD.n401 0.00587931
R997 VDD.n384 VDD.n383 0.00587931
R998 VDD.n357 VDD 0.00579412
R999 VDD VDD.n504 0.00579412
R1000 VDD.n156 VDD 0.00501883
R1001 VDD.n47 VDD 0.00493946
R1002 VDD.n89 VDD 0.00478571
R1003 VDD VDD.n60 0.0045
R1004 VDD.n303 VDD.n302 0.00419863
R1005 VDD VDD.n507 0.00400649
R1006 VDD.n54 VDD 0.004
R1007 VDD.n144 VDD 0.00388028
R1008 VDD.n148 VDD 0.00380275
R1009 VDD.n158 VDD 0.00380275
R1010 VDD.n497 VDD 0.00380275
R1011 VDD.n87 VDD.n86 0.00371429
R1012 VDD.n153 VDD 0.0036441
R1013 VDD.n208 VDD 0.00307143
R1014 VDD.n348 VDD.n347 0.00272472
R1015 VDD.n324 VDD.n323 0.00252247
R1016 VDD.n185 VDD 0.00242233
R1017 VDD.n318 VDD 0.00224194
R1018 VDD.n321 VDD 0.00224194
R1019 VDD.n374 VDD 0.00224194
R1020 VDD.n377 VDD 0.00224194
R1021 VDD.n345 VDD.n344 0.00211798
R1022 VDD.n327 VDD.n326 0.00211798
R1023 VDD.n86 VDD.n83 0.00210714
R1024 VDD.n175 VDD.n174 0.00208824
R1025 VDD VDD.n190 0.00191176
R1026 VDD.n181 VDD 0.00189806
R1027 VDD VDD.n187 0.0017233
R1028 VDD.n434 VDD.n432 0.00167963
R1029 VDD.n491 VDD.n168 0.00166883
R1030 VDD.n413 VDD 0.00166883
R1031 VDD.n33 VDD 0.00166129
R1032 VDD.n30 VDD 0.00166129
R1033 VDD VDD.n27 0.00166129
R1034 VDD VDD.n24 0.00166129
R1035 VDD VDD.n37 0.00166129
R1036 VDD.n41 VDD 0.00166129
R1037 VDD VDD.n44 0.00166129
R1038 VDD.n101 VDD 0.00166129
R1039 VDD.n98 VDD 0.00166129
R1040 VDD VDD.n95 0.00166129
R1041 VDD VDD.n92 0.00166129
R1042 VDD.n487 VDD 0.00166129
R1043 VDD.n484 VDD 0.00166129
R1044 VDD VDD.n481 0.00166129
R1045 VDD VDD.n478 0.00166129
R1046 VDD.n269 VDD 0.00166129
R1047 VDD.n266 VDD 0.00166129
R1048 VDD VDD.n263 0.00166129
R1049 VDD VDD.n260 0.00166129
R1050 VDD.n220 VDD 0.00166129
R1051 VDD.n217 VDD 0.00166129
R1052 VDD VDD.n214 0.00166129
R1053 VDD VDD.n211 0.00166129
R1054 VDD.n357 VDD 0.00155882
R1055 VDD VDD.n426 0.00152662
R1056 VDD.n66 VDD 0.00130718
R1057 VDD.n105 VDD 0.00130718
R1058 VDD VDD.n114 0.00130718
R1059 VDD VDD.n120 0.00130718
R1060 VDD.n123 VDD 0.00130718
R1061 VDD VDD.n432 0.00118702
R1062 VDD VDD.n430 0.00118702
R1063 VDD VDD.n430 0.00118702
R1064 VDD VDD.n428 0.00118702
R1065 VDD VDD.n428 0.00118702
R1066 VDD VDD.n426 0.00118441
R1067 VDD VDD.n393 0.00112069
R1068 VDD VDD.n388 0.00112069
R1069 VDD VDD.n382 0.00112069
R1070 VDD VDD.n336 0.00110674
R1071 VDD VDD.n331 0.00110674
R1072 VDD VDD.n325 0.00110674
R1073 VDD.n309 VDD 0.00108064
R1074 VDD VDD.n312 0.00108064
R1075 VDD.n365 VDD 0.00108064
R1076 VDD VDD.n368 0.00108064
R1077 VDD VDD.n434 0.00100731
R1078 VDD.n193 VDD 0.00100139
R1079 VDD VDD.n405 0.000913793
R1080 VDD.n403 VDD 0.000913793
R1081 VDD.n397 VDD 0.000913793
R1082 VDD.n392 VDD 0.000913793
R1083 VDD VDD.n385 0.000913793
R1084 VDD.n380 VDD 0.000913793
R1085 VDD VDD.n348 0.000904494
R1086 VDD.n346 VDD 0.000904494
R1087 VDD.n340 VDD 0.000904494
R1088 VDD.n335 VDD 0.000904494
R1089 VDD VDD.n328 0.000904494
R1090 VDD.n323 VDD 0.000904494
R1091 VDD.n493 VDD.n492 0.000893013
R1092 VDD VDD.n169 0.000849515
R1093 VDD VDD.n185 0.000849515
R1094 VDD VDD.n170 0.000849515
R1095 VDD.n400 VDD 0.000706897
R1096 VDD.n343 VDD 0.000702247
R1097 VSS.n158 VSS.n157 3.10619e+06
R1098 VSS.n158 VSS.n103 685750
R1099 VSS.n310 VSS.n309 26028.4
R1100 VSS.n276 VSS.n274 18801.2
R1101 VSS.n79 VSS.n71 16250
R1102 VSS.n156 VSS.n155 9901.08
R1103 VSS.n102 VSS.n98 9750
R1104 VSS.n51 VSS.n50 7243.74
R1105 VSS.n232 VSS.n231 5598.39
R1106 VSS.n277 VSS.n276 5365.74
R1107 VSS.n142 VSS.n129 5347.83
R1108 VSS.t120 VSS.n338 4659.04
R1109 VSS.n48 VSS.n47 4152.58
R1110 VSS.n134 VSS.t33 4024.27
R1111 VSS.n273 VSS.n217 3893.61
R1112 VSS.n308 VSS.t270 3750
R1113 VSS.n9 VSS.n8 3574.4
R1114 VSS.n120 VSS.n119 3494.13
R1115 VSS.n378 VSS.n377 3330.48
R1116 VSS.n157 VSS.n156 3205.8
R1117 VSS.n338 VSS.n44 2949.84
R1118 VSS.n309 VSS.n206 2896.63
R1119 VSS.t302 VSS.t87 2781.65
R1120 VSS.n322 VSS.n45 2502.44
R1121 VSS.n231 VSS.t265 2336.12
R1122 VSS.t86 VSS.t83 2307.56
R1123 VSS.t195 VSS.t154 2307.56
R1124 VSS.t157 VSS.t165 2307.56
R1125 VSS.t217 VSS.t304 2307.56
R1126 VSS.t2 VSS.t162 2307.56
R1127 VSS.t130 VSS.t262 2307.56
R1128 VSS.t66 VSS.t258 2307.56
R1129 VSS.t126 VSS.t149 2307.56
R1130 VSS.t72 VSS.t91 2307.56
R1131 VSS.t152 VSS.t97 2307.56
R1132 VSS.t249 VSS.t26 2307.56
R1133 VSS.t224 VSS.t255 2307.56
R1134 VSS.t227 VSS.t240 2307.56
R1135 VSS.t57 VSS.t89 2307.56
R1136 VSS.t299 VSS.t209 2307.56
R1137 VSS.t68 VSS.t123 2307.56
R1138 VSS.t159 VSS.t220 2307.56
R1139 VSS.t1 VSS.t139 2307.56
R1140 VSS.n10 VSS.n9 2206.03
R1141 VSS.n129 VSS.t75 2085.4
R1142 VSS.n13 VSS.t252 2062.12
R1143 VSS.n15 VSS.t243 2062.12
R1144 VSS.t180 VSS.n386 2062.12
R1145 VSS.t167 VSS.n385 2062.12
R1146 VSS.n14 VSS.t215 2058.2
R1147 VSS.t46 VSS.n217 1806.5
R1148 VSS.t301 VSS.n217 1802.23
R1149 VSS.t254 VSS.t188 1725.36
R1150 VSS.t197 VSS.t16 1725.36
R1151 VSS.t69 VSS.t131 1725.36
R1152 VSS.t297 VSS.t169 1725.36
R1153 VSS.n274 VSS.t0 1713.53
R1154 VSS.t3 VSS.n51 1672
R1155 VSS.n50 VSS.n46 1611.34
R1156 VSS.t171 VSS.n232 1601.22
R1157 VSS.n206 VSS.n205 1597.63
R1158 VSS.n155 VSS.t12 1577.93
R1159 VSS.n274 VSS.n273 1565.03
R1160 VSS.n129 VSS.t24 1513.35
R1161 VSS.t166 VSS.t103 1450.83
R1162 VSS.t76 VSS.t256 1450.83
R1163 VSS.t125 VSS.t141 1438.12
R1164 VSS.t109 VSS.t151 1438.12
R1165 VSS.t85 VSS.t229 1436.54
R1166 VSS.n305 VSS.n210 1405.57
R1167 VSS.n309 VSS.n308 1350.61
R1168 VSS.n388 VSS.n387 1293.73
R1169 VSS.n173 VSS.n158 1282.2
R1170 VSS.n6 VSS.t207 1272.1
R1171 VSS.n142 VSS.t272 1226.37
R1172 VSS.t48 VSS.n144 1199.47
R1173 VSS.t50 VSS.n134 1199.47
R1174 VSS.n173 VSS.t37 1199.47
R1175 VSS.n7 VSS.t266 1199.47
R1176 VSS.n377 VSS.t98 1153.78
R1177 VSS.n128 VSS.t77 1152.75
R1178 VSS.n124 VSS.n123 1119.51
R1179 VSS.t269 VSS.n105 1117.74
R1180 VSS.t40 VSS.n322 1035.69
R1181 VSS.t245 VSS.t10 1016.25
R1182 VSS.t67 VSS.t116 1015.47
R1183 VSS.n119 VSS.n26 961.587
R1184 VSS.n50 VSS.n49 960.539
R1185 VSS.n209 VSS.t18 927.717
R1186 VSS.n210 VSS.t21 919.253
R1187 VSS.n293 VSS.t4 919.253
R1188 VSS.t81 VSS.t13 913.885
R1189 VSS.t122 VSS.t296 913.885
R1190 VSS.t102 VSS.t2 913.885
R1191 VSS.t97 VSS.t251 913.885
R1192 VSS.t89 VSS.t211 913.885
R1193 VSS.t203 VSS.t1 913.885
R1194 VSS.n307 VSS.n209 879.836
R1195 VSS.n381 VSS.n380 839.716
R1196 VSS.n119 VSS.t35 808.298
R1197 VSS.n235 VSS.t198 776.83
R1198 VSS.n205 VSS.t14 771.441
R1199 VSS.n288 VSS.t175 753.193
R1200 VSS.n276 VSS.n275 749.452
R1201 VSS.n8 VSS.n7 738.636
R1202 VSS.n30 VSS.t7 728.939
R1203 VSS.n305 VSS.t182 709.049
R1204 VSS.n30 VSS.t231 707.605
R1205 VSS.n322 VSS.t279 703.503
R1206 VSS.t115 VSS.t226 683.312
R1207 VSS.t206 VSS.t197 683.312
R1208 VSS.t55 VSS.t222 683.312
R1209 VSS.t212 VSS.t297 683.312
R1210 VSS.n308 VSS.n207 676.096
R1211 VSS.n307 VSS.n306 673.139
R1212 VSS.n101 VSS.n100 629.365
R1213 VSS.n88 VSS.n87 629.365
R1214 VSS.n96 VSS.n95 626.053
R1215 VSS.n85 VSS.n84 626.053
R1216 VSS.n72 VSS.n70 616.962
R1217 VSS.n200 VSS.n199 616.962
R1218 VSS.n78 VSS.n77 615.048
R1219 VSS.n82 VSS.n81 615.048
R1220 VSS.t121 VSS.t76 574.587
R1221 VSS.t138 VSS.t90 569.552
R1222 VSS.t151 VSS.t53 569.552
R1223 VSS.t113 VSS.t156 568.928
R1224 VSS.t87 VSS.n235 554.879
R1225 VSS.t12 VSS.n154 548.331
R1226 VSS.n125 VSS.t86 548.331
R1227 VSS.n126 VSS.t195 548.331
R1228 VSS.n145 VSS.t81 548.331
R1229 VSS.t272 VSS.n141 548.331
R1230 VSS.t165 VSS.n140 548.331
R1231 VSS.t304 VSS.n139 548.331
R1232 VSS.n135 VSS.t122 548.331
R1233 VSS.n172 VSS.t102 548.331
R1234 VSS.n171 VSS.t130 548.331
R1235 VSS.n170 VSS.t66 548.331
R1236 VSS.n169 VSS.t3 548.331
R1237 VSS.t98 VSS.n376 548.331
R1238 VSS.n22 VSS.t126 548.331
R1239 VSS.n23 VSS.t72 548.331
R1240 VSS.t265 VSS.n230 548.331
R1241 VSS.t255 VSS.n229 548.331
R1242 VSS.t240 VSS.n228 548.331
R1243 VSS.t211 VSS.n227 548.331
R1244 VSS.t0 VSS.n0 548.331
R1245 VSS.n1 VSS.t68 548.331
R1246 VSS.n2 VSS.t159 548.331
R1247 VSS.n3 VSS.t203 548.331
R1248 VSS.n239 VSS.t298 546.41
R1249 VSS.t30 VSS.n310 512.745
R1250 VSS.n103 VSS.n88 491.8
R1251 VSS.n102 VSS.n101 484.921
R1252 VSS.n98 VSS.n85 472.106
R1253 VSS.n206 VSS.n70 468.62
R1254 VSS.t273 VSS.n280 455.26
R1255 VSS.n281 VSS.t61 455.26
R1256 VSS.n97 VSS.n96 455
R1257 VSS.n199 VSS.n71 448.392
R1258 VSS.n49 VSS.n48 443.99
R1259 VSS.n79 VSS.n78 430.197
R1260 VSS.n82 VSS.n79 426.837
R1261 VSS.n121 VSS.n120 420.916
R1262 VSS.n249 VSS.t196 409.988
R1263 VSS.n250 VSS.t254 409.988
R1264 VSS.n254 VSS.t115 409.988
R1265 VSS.n255 VSS.t206 409.988
R1266 VSS.n258 VSS.t301 409.988
R1267 VSS.n259 VSS.t69 409.988
R1268 VSS.n260 VSS.t55 409.988
R1269 VSS.n261 VSS.t212 409.988
R1270 VSS.n41 VSS.t8 404.618
R1271 VSS.t10 VSS.t283 402.478
R1272 VSS.t56 VSS.t291 402.478
R1273 VSS.t71 VSS.t285 402.166
R1274 VSS.t137 VSS.t261 402.166
R1275 VSS.n338 VSS.n51 378.765
R1276 VSS.n174 VSS.t99 372.873
R1277 VSS.n154 VSS.t83 365.555
R1278 VSS.t154 VSS.n125 365.555
R1279 VSS.n126 VSS.t135 365.555
R1280 VSS.n145 VSS.t48 365.555
R1281 VSS.n141 VSS.t157 365.555
R1282 VSS.n140 VSS.t217 365.555
R1283 VSS.n139 VSS.t201 365.555
R1284 VSS.n135 VSS.t50 365.555
R1285 VSS.t37 VSS.n172 365.555
R1286 VSS.t162 VSS.n171 365.555
R1287 VSS.t262 VSS.n170 365.555
R1288 VSS.t258 VSS.n169 365.555
R1289 VSS.n376 VSS.t149 365.555
R1290 VSS.t91 VSS.n22 365.555
R1291 VSS.n23 VSS.t152 365.555
R1292 VSS.t26 VSS.n24 365.555
R1293 VSS.n230 VSS.t224 365.555
R1294 VSS.n229 VSS.t227 365.555
R1295 VSS.n228 VSS.t57 365.555
R1296 VSS.n227 VSS.t299 365.555
R1297 VSS.t123 VSS.n0 365.555
R1298 VSS.t220 VSS.n1 365.555
R1299 VSS.t139 VSS.n2 365.555
R1300 VSS.t266 VSS.n3 365.555
R1301 VSS.n239 VSS.t204 364.274
R1302 VSS.n296 VSS.n209 347.168
R1303 VSS.n35 VSS.t166 344.752
R1304 VSS.n37 VSS.t114 344.752
R1305 VSS.n108 VSS.t269 341.731
R1306 VSS.n109 VSS.t125 341.731
R1307 VSS.n118 VSS.t53 341.731
R1308 VSS.n27 VSS.t54 341.358
R1309 VSS.n28 VSS.t85 341.358
R1310 VSS.n29 VSS.t113 341.358
R1311 VSS.n31 VSS.t80 341.358
R1312 VSS.n34 VSS.n33 337.57
R1313 VSS.t11 VSS.t294 337.038
R1314 VSS.t268 VSS.t213 337.038
R1315 VSS.t233 VSS.t146 335.264
R1316 VSS.t79 VSS.t173 335.264
R1317 VSS.t70 VSS.t59 330.394
R1318 VSS.t119 VSS.t286 330.394
R1319 VSS.t82 VSS.t64 329.37
R1320 VSS.t52 VSS.t107 329.37
R1321 VSS.t188 VSS.n249 273.325
R1322 VSS.n250 VSS.t241 273.325
R1323 VSS.t16 VSS.n254 273.325
R1324 VSS.n255 VSS.t46 273.325
R1325 VSS.t131 VSS.n258 273.325
R1326 VSS.n259 VSS.t160 273.325
R1327 VSS.t169 VSS.n260 273.325
R1328 VSS.n261 VSS.t28 273.325
R1329 VSS.n38 VSS.t121 272.928
R1330 VSS.n12 VSS.n11 266.587
R1331 VSS.t283 VSS.n323 241.487
R1332 VSS.n325 VSS.t56 241.487
R1333 VSS.n327 VSS.t223 241.487
R1334 VSS.n339 VSS.t120 241.487
R1335 VSS.n311 VSS.t71 241.299
R1336 VSS.n314 VSS.t137 241.299
R1337 VSS.n317 VSS.t67 241.299
R1338 VSS.t279 VSS.n321 241.299
R1339 VSS.t190 VSS.n277 237.15
R1340 VSS.t103 VSS.n34 229.834
R1341 VSS.n35 VSS.t305 229.834
R1342 VSS.t256 VSS.n37 229.834
R1343 VSS.t33 VSS.n39 229.834
R1344 VSS.t141 VSS.n108 227.821
R1345 VSS.n109 VSS.t73 227.821
R1346 VSS.n114 VSS.t109 227.821
R1347 VSS.t35 VSS.n118 227.821
R1348 VSS.t229 VSS.n27 227.571
R1349 VSS.n28 VSS.t193 227.571
R1350 VSS.t231 VSS.n29 227.571
R1351 VSS.t24 VSS.n31 227.571
R1352 VSS.n36 VSS.t219 211.879
R1353 VSS.n155 VSS.n124 204.131
R1354 VSS.n338 VSS.n45 196.673
R1355 VSS.n100 VSS.t11 196.032
R1356 VSS.n87 VSS.t268 196.032
R1357 VSS.n95 VSS.t233 195
R1358 VSS.n84 VSS.t79 195
R1359 VSS.n72 VSS.t70 192.168
R1360 VSS.n200 VSS.t119 192.168
R1361 VSS.n77 VSS.t82 191.572
R1362 VSS.n81 VSS.t52 191.572
R1363 VSS.n112 VSS.t138 181.544
R1364 VSS.n288 VSS.n207 171.989
R1365 VSS.n105 VSS.n104 167.306
R1366 VSS.t175 VSS.t178 166.059
R1367 VSS.n323 VSS.t40 160.992
R1368 VSS.n325 VSS.t245 160.992
R1369 VSS.n327 VSS.t93 160.992
R1370 VSS.n339 VSS.t237 160.992
R1371 VSS.n311 VSS.t30 160.867
R1372 VSS.n314 VSS.t143 160.867
R1373 VSS.n317 VSS.t127 160.867
R1374 VSS.n321 VSS.t116 160.867
R1375 VSS.n306 VSS.n305 154.197
R1376 VSS.n273 VSS.n272 119.948
R1377 VSS.t96 VSS.t280 112.944
R1378 VSS.n380 VSS.n379 100.334
R1379 VSS.n10 VSS.t235 86.249
R1380 VSS.t252 VSS.n12 86.249
R1381 VSS.t215 VSS.n13 86.249
R1382 VSS.t243 VSS.n14 86.249
R1383 VSS.n15 VSS.t133 86.249
R1384 VSS.n387 VSS.t180 86.249
R1385 VSS.n386 VSS.t167 86.249
R1386 VSS.n385 VSS.t289 86.249
R1387 VSS.n380 VSS.t185 74.768
R1388 VSS.t182 VSS.n304 72.8445
R1389 VSS.n379 VSS.n378 59.271
R1390 VSS.n308 VSS.n208 56.3094
R1391 VSS.n233 VSS.t171 47.5615
R1392 VSS.n7 VSS.n6 41.0359
R1393 VSS.n337 VSS.t43 40.3374
R1394 VSS.n144 VSS.n128 37.1859
R1395 VSS.n272 VSS.t209 34.2711
R1396 VSS.n236 VSS.t302 34.1511
R1397 VSS.n144 VSS.n143 29.7488
R1398 VSS.t43 VSS.t96 25.3551
R1399 VSS.n121 VSS.t249 22.8476
R1400 VSS.t54 VSS.n26 21.3353
R1401 VSS.n98 VSS.n97 20.5268
R1402 VSS.n280 VSS.t190 19.0418
R1403 VSS.n281 VSS.t273 19.0418
R1404 VSS.t61 VSS.n208 18.7705
R1405 VSS.n206 VSS.n71 16.8573
R1406 VSS.n143 VSS.n142 16.6063
R1407 VSS.n308 VSS.n307 13.8894
R1408 VSS.n134 VSS.n41 13.0527
R1409 VSS.n123 VSS.n121 11.424
R1410 VSS.n103 VSS.n102 10.318
R1411 VSS.n289 VSS.t179 10.2719
R1412 VSS.n174 VSS.n173 9.623
R1413 VSS VSS.t271 9.43705
R1414 VSS.n5 VSS.t208 9.3736
R1415 VSS.n122 VSS.t250 9.3736
R1416 VSS.n127 VSS.t78 9.3736
R1417 VSS.n271 VSS.t210 9.3736
R1418 VSS.n175 VSS.n93 9.37275
R1419 VSS.n336 VSS.n52 9.37275
R1420 VSS.n238 VSS.t303 9.36521
R1421 VSS.n73 VSS.t60 9.3533
R1422 VSS.n94 VSS.t147 9.3533
R1423 VSS.n83 VSS.t174 9.3533
R1424 VSS.n99 VSS.t295 9.35181
R1425 VSS.n86 VSS.t214 9.35181
R1426 VSS.n279 VSS.n278 9.33837
R1427 VSS.n287 VSS.n285 9.3221
R1428 VSS.n244 VSS.n234 9.3221
R1429 VSS.n242 VSS.t88 9.3221
R1430 VSS.n201 VSS.t287 9.31766
R1431 VSS.n76 VSS.t65 9.31744
R1432 VSS.n80 VSS.t108 9.31744
R1433 VSS.n341 VSS.t9 9.30652
R1434 VSS.n203 VSS.t15 9.30652
R1435 VSS.n21 VSS.n20 9.30652
R1436 VSS.n299 VSS.n211 9.30652
R1437 VSS.n297 VSS.n212 9.30652
R1438 VSS.n245 VSS.t172 9.30652
R1439 VSS.n399 VSS.t236 9.30518
R1440 VSS.n396 VSS.t253 9.30518
R1441 VSS.n394 VSS.t216 9.30518
R1442 VSS.n392 VSS.t244 9.30518
R1443 VSS.n390 VSS.t134 9.30518
R1444 VSS.n17 VSS.t181 9.30518
R1445 VSS.n300 VSS.t168 9.30518
R1446 VSS.n383 VSS.t290 9.30518
R1447 VSS.n292 VSS.n291 9.28776
R1448 VSS.n295 VSS.n213 9.26757
R1449 VSS.n283 VSS.n214 9.26488
R1450 VSS.n216 VSS.n215 9.26488
R1451 VSS VSS.t205 7.30633
R1452 VSS.n106 VSS.t142 7.19156
R1453 VSS.n111 VSS.t74 7.19156
R1454 VSS.n167 VSS.n166 7.19156
R1455 VSS.n164 VSS.n163 7.19156
R1456 VSS.n161 VSS.n160 7.19156
R1457 VSS.n59 VSS.n57 7.19156
R1458 VSS.n61 VSS.n56 7.19156
R1459 VSS.n63 VSS.n55 7.19156
R1460 VSS.n43 VSS.n42 7.19156
R1461 VSS.n329 VSS.n326 7.19156
R1462 VSS.n363 VSS.t230 7.19156
R1463 VSS.n361 VSS.t194 7.19156
R1464 VSS.n152 VSS.t84 7.19156
R1465 VSS.n150 VSS.t155 7.19156
R1466 VSS.n148 VSS.t136 7.19156
R1467 VSS.n131 VSS.t158 7.19156
R1468 VSS.n133 VSS.t218 7.19156
R1469 VSS.n137 VSS.t202 7.19156
R1470 VSS.n319 VSS.n67 7.19156
R1471 VSS.n316 VSS.n68 7.19156
R1472 VSS.n374 VSS.t150 7.19156
R1473 VSS.n372 VSS.t92 7.19156
R1474 VSS.n370 VSS.t153 7.19156
R1475 VSS.n247 VSS.t189 7.19156
R1476 VSS.n252 VSS.t242 7.19156
R1477 VSS.n221 VSS.t225 7.19156
R1478 VSS.n223 VSS.t228 7.19156
R1479 VSS.n225 VSS.t58 7.19156
R1480 VSS.n267 VSS.t132 7.19156
R1481 VSS.n265 VSS.t161 7.19156
R1482 VSS.n409 VSS.t124 7.19156
R1483 VSS.n407 VSS.t221 7.19156
R1484 VSS.n405 VSS.t140 7.19156
R1485 VSS.t75 VSS.n33 7.18282
R1486 VSS.n352 VSS.t104 7.17823
R1487 VSS.n350 VSS.t306 7.17823
R1488 VSS.n179 VSS.t278 7.14823
R1489 VSS.n178 VSS.t284 7.14823
R1490 VSS.n197 VSS.t248 7.13989
R1491 VSS.n185 VSS.t234 7.13989
R1492 VSS.n184 VSS.t148 7.13989
R1493 VSS.n196 VSS.t276 7.13989
R1494 VSS.n191 VSS.t288 7.12156
R1495 VSS.n190 VSS.t277 7.12156
R1496 VSS.n54 VSS.n45 6.85706
R1497 VSS.n302 VSS.n301 6.06679
R1498 VSS.n116 VSS.t110 5.91399
R1499 VSS.n25 VSS.t36 5.91399
R1500 VSS.n92 VSS.n91 5.91399
R1501 VSS.n65 VSS.n53 5.91399
R1502 VSS.n331 VSS.n324 5.91399
R1503 VSS.n333 VSS.n66 5.91399
R1504 VSS.n359 VSS.t232 5.91399
R1505 VSS.n356 VSS.t25 5.91399
R1506 VSS.n146 VSS.t49 5.91399
R1507 VSS.n40 VSS.t51 5.91399
R1508 VSS.n313 VSS.n69 5.91399
R1509 VSS.n90 VSS.n89 5.91399
R1510 VSS.n368 VSS.t27 5.91399
R1511 VSS.n219 VSS.t17 5.91399
R1512 VSS.n257 VSS.t47 5.91399
R1513 VSS.n218 VSS.t300 5.91399
R1514 VSS.n263 VSS.t170 5.91399
R1515 VSS.n4 VSS.t29 5.91399
R1516 VSS.n403 VSS.t267 5.91399
R1517 VSS.n347 VSS.t257 5.90065
R1518 VSS.n344 VSS.t34 5.90065
R1519 VSS.n304 VSS.n303 5.82215
R1520 VSS.n284 VSS.n208 5.40486
R1521 VSS.n389 VSS.n388 5.2005
R1522 VSS.n398 VSS.n11 5.2005
R1523 VSS.n400 VSS.n10 5.2005
R1524 VSS.n397 VSS.n12 5.2005
R1525 VSS.n395 VSS.n13 5.2005
R1526 VSS.n393 VSS.n14 5.2005
R1527 VSS.n391 VSS.n15 5.2005
R1528 VSS.n387 VSS.n16 5.2005
R1529 VSS.n385 VSS.n384 5.2005
R1530 VSS.n386 VSS.n18 5.2005
R1531 VSS.n154 VSS.n153 5.2005
R1532 VSS.n151 VSS.n125 5.2005
R1533 VSS.n149 VSS.n126 5.2005
R1534 VSS.n147 VSS.n145 5.2005
R1535 VSS.n136 VSS.n135 5.2005
R1536 VSS.n139 VSS.n138 5.2005
R1537 VSS.n140 VSS.n132 5.2005
R1538 VSS.n141 VSS.n130 5.2005
R1539 VSS.n353 VSS.n34 5.2005
R1540 VSS.n351 VSS.n35 5.2005
R1541 VSS.n348 VSS.n37 5.2005
R1542 VSS.n345 VSS.n39 5.2005
R1543 VSS.n354 VSS.n33 5.2005
R1544 VSS.n349 VSS.n36 5.2005
R1545 VSS.n346 VSS.n38 5.2005
R1546 VSS.n342 VSS.n41 5.2005
R1547 VSS.n332 VSS.n323 5.2005
R1548 VSS.n330 VSS.n325 5.2005
R1549 VSS.n328 VSS.n327 5.2005
R1550 VSS.n340 VSS.n339 5.2005
R1551 VSS.n58 VSS.n54 5.2005
R1552 VSS.n60 VSS.n54 5.2005
R1553 VSS.n62 VSS.n54 5.2005
R1554 VSS.n64 VSS.n54 5.2005
R1555 VSS.n337 VSS.n336 5.2005
R1556 VSS.n312 VSS.n311 5.2005
R1557 VSS.n315 VSS.n314 5.2005
R1558 VSS.n318 VSS.n317 5.2005
R1559 VSS.n321 VSS.n320 5.2005
R1560 VSS.n73 VSS.n72 5.2005
R1561 VSS.n201 VSS.n200 5.2005
R1562 VSS.n199 VSS.n198 5.2005
R1563 VSS.n77 VSS.n76 5.2005
R1564 VSS.n192 VSS.n82 5.2005
R1565 VSS.n81 VSS.n80 5.2005
R1566 VSS.n95 VSS.n94 5.2005
R1567 VSS.n186 VSS.n85 5.2005
R1568 VSS.n84 VSS.n83 5.2005
R1569 VSS.n100 VSS.n99 5.2005
R1570 VSS.n180 VSS.n88 5.2005
R1571 VSS.n87 VSS.n86 5.2005
R1572 VSS.n175 VSS.n174 5.2005
R1573 VSS.n169 VSS.n168 5.2005
R1574 VSS.n170 VSS.n165 5.2005
R1575 VSS.n171 VSS.n162 5.2005
R1576 VSS.n172 VSS.n159 5.2005
R1577 VSS.n128 VSS.n127 5.2005
R1578 VSS.n357 VSS.n31 5.2005
R1579 VSS.n360 VSS.n29 5.2005
R1580 VSS.n362 VSS.n28 5.2005
R1581 VSS.n364 VSS.n27 5.2005
R1582 VSS.n358 VSS.n30 5.2005
R1583 VSS.n365 VSS.n26 5.2005
R1584 VSS.n123 VSS.n122 5.2005
R1585 VSS.n376 VSS.n375 5.2005
R1586 VSS.n373 VSS.n22 5.2005
R1587 VSS.n371 VSS.n23 5.2005
R1588 VSS.n369 VSS.n24 5.2005
R1589 VSS.n118 VSS.n117 5.2005
R1590 VSS.n115 VSS.n114 5.2005
R1591 VSS.n110 VSS.n109 5.2005
R1592 VSS.n108 VSS.n107 5.2005
R1593 VSS.n113 VSS.n112 5.2005
R1594 VSS.n105 VSS.n19 5.2005
R1595 VSS.n298 VSS.n210 5.2005
R1596 VSS.n294 VSS.n293 5.2005
R1597 VSS.n286 VSS.n207 5.2005
R1598 VSS.n289 VSS.n288 5.2005
R1599 VSS.n205 VSS.n204 5.2005
R1600 VSS.n280 VSS.n279 5.2005
R1601 VSS.n282 VSS.n281 5.2005
R1602 VSS.n240 VSS.n239 5.2005
R1603 VSS.n237 VSS.n236 5.2005
R1604 VSS.n243 VSS.n235 5.2005
R1605 VSS.n246 VSS.n233 5.2005
R1606 VSS.n6 VSS.n5 5.2005
R1607 VSS.n262 VSS.n261 5.2005
R1608 VSS.n264 VSS.n260 5.2005
R1609 VSS.n266 VSS.n259 5.2005
R1610 VSS.n268 VSS.n258 5.2005
R1611 VSS.n256 VSS.n255 5.2005
R1612 VSS.n254 VSS.n253 5.2005
R1613 VSS.n251 VSS.n250 5.2005
R1614 VSS.n249 VSS.n248 5.2005
R1615 VSS.n230 VSS.n220 5.2005
R1616 VSS.n229 VSS.n222 5.2005
R1617 VSS.n228 VSS.n224 5.2005
R1618 VSS.n227 VSS.n226 5.2005
R1619 VSS.n272 VSS.n271 5.2005
R1620 VSS.n410 VSS.n0 5.2005
R1621 VSS.n408 VSS.n1 5.2005
R1622 VSS.n406 VSS.n2 5.2005
R1623 VSS.n404 VSS.n3 5.2005
R1624 VSS.n178 VSS.n177 4.93566
R1625 VSS.n338 VSS.n337 4.61043
R1626 VSS.n382 VSS 2.96937
R1627 VSS.n341 VSS 2.0829
R1628 VSS.n344 VSS.n343 0.850616
R1629 VSS.n355 VSS.n32 0.845914
R1630 VSS.n367 VSS.n366 0.845914
R1631 VSS.n270 VSS.n269 0.845914
R1632 VSS.n335 VSS.n334 0.844811
R1633 VSS.n177 VSS.n90 0.729114
R1634 VSS.n402 VSS.n401 0.637841
R1635 VSS.n164 VSS 0.343161
R1636 VSS.n167 VSS 0.343161
R1637 VSS VSS.n61 0.343161
R1638 VSS VSS.n59 0.343161
R1639 VSS.n152 VSS 0.343161
R1640 VSS.n150 VSS 0.343161
R1641 VSS VSS.n131 0.343161
R1642 VSS VSS.n133 0.343161
R1643 VSS.n374 VSS 0.343161
R1644 VSS.n372 VSS 0.343161
R1645 VSS VSS.n221 0.343161
R1646 VSS VSS.n223 0.343161
R1647 VSS.n409 VSS 0.343161
R1648 VSS.n407 VSS 0.343161
R1649 VSS.n242 VSS.n241 0.309418
R1650 VSS.n334 VSS 0.290741
R1651 VSS VSS.n159 0.289491
R1652 VSS.n64 VSS 0.289491
R1653 VSS VSS.n147 0.289491
R1654 VSS VSS.n136 0.289491
R1655 VSS VSS.n369 0.289491
R1656 VSS.n226 VSS 0.289491
R1657 VSS VSS.n404 0.289491
R1658 VSS.n241 VSS.n240 0.255008
R1659 VSS.n332 VSS.n331 0.253109
R1660 VSS.n330 VSS.n329 0.253109
R1661 VSS.n313 VSS.n312 0.251894
R1662 VSS.n316 VSS.n315 0.251894
R1663 VSS.n161 VSS 0.191234
R1664 VSS VSS.n63 0.191234
R1665 VSS.n148 VSS 0.191234
R1666 VSS.n137 VSS 0.191234
R1667 VSS.n370 VSS 0.191234
R1668 VSS VSS.n225 0.191234
R1669 VSS.n405 VSS 0.191234
R1670 VSS VSS.n43 0.180935
R1671 VSS.n319 VSS 0.180067
R1672 VSS.n245 VSS.n244 0.168119
R1673 VSS VSS.n216 0.152427
R1674 VSS.n283 VSS 0.152427
R1675 VSS.n253 VSS.n252 0.151192
R1676 VSS.n256 VSS.n219 0.151192
R1677 VSS.n265 VSS.n264 0.151192
R1678 VSS.n263 VSS.n262 0.151192
R1679 VSS.n297 VSS 0.151087
R1680 VSS.n295 VSS 0.150362
R1681 VSS.n299 VSS 0.141998
R1682 VSS.n241 VSS.n238 0.141461
R1683 VSS.n402 VSS 0.137685
R1684 VSS.n367 VSS 0.137685
R1685 VSS VSS.n32 0.137685
R1686 VSS VSS.n270 0.137685
R1687 VSS.n176 VSS 0.137136
R1688 VSS VSS.n335 0.137136
R1689 VSS.n287 VSS.n286 0.136634
R1690 VSS.n244 VSS.n243 0.136634
R1691 VSS.n343 VSS.n40 0.135964
R1692 VSS.n162 VSS.n161 0.118573
R1693 VSS.n165 VSS.n164 0.118573
R1694 VSS.n168 VSS.n167 0.118573
R1695 VSS.n63 VSS.n62 0.118573
R1696 VSS.n61 VSS.n60 0.118573
R1697 VSS.n59 VSS.n58 0.118573
R1698 VSS.n153 VSS.n152 0.118573
R1699 VSS.n151 VSS.n150 0.118573
R1700 VSS.n149 VSS.n148 0.118573
R1701 VSS.n131 VSS.n130 0.118573
R1702 VSS.n133 VSS.n132 0.118573
R1703 VSS.n138 VSS.n137 0.118573
R1704 VSS.n375 VSS.n374 0.118573
R1705 VSS.n373 VSS.n372 0.118573
R1706 VSS.n371 VSS.n370 0.118573
R1707 VSS.n221 VSS.n220 0.118573
R1708 VSS.n223 VSS.n222 0.118573
R1709 VSS.n225 VSS.n224 0.118573
R1710 VSS.n410 VSS.n409 0.118573
R1711 VSS.n408 VSS.n407 0.118573
R1712 VSS.n406 VSS.n405 0.118573
R1713 VSS VSS.n242 0.115458
R1714 VSS VSS.n92 0.115271
R1715 VSS.n65 VSS 0.115271
R1716 VSS VSS.n146 0.115271
R1717 VSS VSS.n40 0.115271
R1718 VSS VSS.n368 0.115271
R1719 VSS VSS.n218 0.115271
R1720 VSS VSS.n403 0.115271
R1721 VSS VSS.n302 0.111993
R1722 VSS.n247 VSS 0.108137
R1723 VSS.n267 VSS 0.108137
R1724 VSS.n117 VSS.n116 0.10529
R1725 VSS.n361 VSS.n360 0.10508
R1726 VSS.n194 VSS.n193 0.103269
R1727 VSS.n188 VSS.n187 0.103269
R1728 VSS.n182 VSS.n181 0.103269
R1729 VSS.n355 VSS.n354 0.102565
R1730 VSS.n176 VSS.n92 0.10206
R1731 VSS.n335 VSS.n65 0.10206
R1732 VSS.n146 VSS.n32 0.10206
R1733 VSS.n368 VSS.n367 0.10206
R1734 VSS.n270 VSS.n218 0.10206
R1735 VSS.n403 VSS.n402 0.10206
R1736 VSS.n347 VSS.n346 0.101682
R1737 VSS.n334 VSS.n333 0.0985362
R1738 VSS.n113 VSS.n111 0.0971733
R1739 VSS.n290 VSS.n287 0.0844496
R1740 VSS.n358 VSS.n357 0.08348
R1741 VSS.n352 VSS 0.0753497
R1742 VSS.n106 VSS 0.0753497
R1743 VSS.n363 VSS 0.0752
R1744 VSS.n282 VSS.n216 0.0739862
R1745 VSS.n284 VSS.n283 0.0739862
R1746 VSS.n296 VSS.n295 0.0739862
R1747 VSS VSS.n19 0.0733657
R1748 VSS.n401 VSS 0.0717187
R1749 VSS.n298 VSS.n297 0.066973
R1750 VSS.n381 VSS.n21 0.0666983
R1751 VSS.n196 VSS.n195 0.0664039
R1752 VSS.n190 VSS.n189 0.0637265
R1753 VSS.n329 VSS.n328 0.0626739
R1754 VSS.n340 VSS.n43 0.0626739
R1755 VSS.n318 VSS.n316 0.062375
R1756 VSS.n320 VSS.n319 0.062375
R1757 VSS.n303 VSS.n299 0.0618793
R1758 VSS.n75 VSS.n74 0.061873
R1759 VSS.n333 VSS 0.0609348
R1760 VSS.n331 VSS 0.0609348
R1761 VSS.n90 VSS 0.0606442
R1762 VSS VSS.n313 0.0606442
R1763 VSS.n177 VSS.n176 0.059582
R1764 VSS.n269 VSS.n257 0.0593761
R1765 VSS.n238 VSS.n237 0.0589274
R1766 VSS.n269 VSS 0.0580792
R1767 VSS.n349 VSS.n348 0.0573136
R1768 VSS.n246 VSS.n245 0.0564843
R1769 VSS.n396 VSS 0.0553671
R1770 VSS VSS.n17 0.0553671
R1771 VSS.n394 VSS 0.0552176
R1772 VSS.n292 VSS.n290 0.0540556
R1773 VSS.n366 VSS 0.0537064
R1774 VSS.n184 VSS 0.053635
R1775 VSS.n401 VSS.n4 0.0533747
R1776 VSS VSS.n365 0.0532782
R1777 VSS.n383 VSS.n382 0.0514681
R1778 VSS.n74 VSS 0.0502725
R1779 VSS.n389 VSS 0.0495365
R1780 VSS.n350 VSS.n349 0.048476
R1781 VSS.n399 VSS.n398 0.0455
R1782 VSS.n202 VSS.n74 0.0423182
R1783 VSS.n366 VSS.n25 0.0414419
R1784 VSS.n356 VSS.n355 0.04136
R1785 VSS.n248 VSS.n247 0.0375893
R1786 VSS.n252 VSS.n251 0.0375893
R1787 VSS.n268 VSS.n267 0.0375893
R1788 VSS.n266 VSS.n265 0.0375893
R1789 VSS.n301 VSS 0.0366794
R1790 VSS VSS.n219 0.0365519
R1791 VSS.n257 VSS 0.0365519
R1792 VSS VSS.n263 0.0365519
R1793 VSS VSS.n4 0.0365519
R1794 VSS.n294 VSS.n292 0.032289
R1795 VSS.n202 VSS 0.0311818
R1796 VSS.n343 VSS 0.030089
R1797 VSS.n203 VSS.n202 0.0295323
R1798 VSS VSS.n197 0.0289211
R1799 VSS VSS.n191 0.0289211
R1800 VSS VSS.n185 0.0289211
R1801 VSS VSS.n179 0.0289211
R1802 VSS.n392 VSS 0.0278588
R1803 VSS.n400 VSS.n399 0.0272608
R1804 VSS.n397 VSS.n396 0.0272608
R1805 VSS.n395 VSS.n394 0.0272608
R1806 VSS.n393 VSS.n392 0.0272608
R1807 VSS.n391 VSS.n390 0.0272608
R1808 VSS.n17 VSS.n16 0.0272608
R1809 VSS.n300 VSS.n18 0.0272608
R1810 VSS.n384 VSS.n383 0.0272608
R1811 VSS.n292 VSS 0.026922
R1812 VSS.n353 VSS.n352 0.0262916
R1813 VSS.n351 VSS.n350 0.0262916
R1814 VSS.n107 VSS.n106 0.0262916
R1815 VSS.n111 VSS.n110 0.0262916
R1816 VSS.n364 VSS.n363 0.02624
R1817 VSS.n362 VSS.n361 0.02624
R1818 VSS VSS.n347 0.0255701
R1819 VSS VSS.n344 0.0255701
R1820 VSS.n116 VSS 0.0255701
R1821 VSS VSS.n25 0.0255701
R1822 VSS.n302 VSS.n21 0.0255299
R1823 VSS VSS.n359 0.02552
R1824 VSS VSS.n356 0.02552
R1825 VSS.n342 VSS.n341 0.0248493
R1826 VSS.n359 VSS.n358 0.0221
R1827 VSS.n195 VSS 0.0205495
R1828 VSS.n194 VSS 0.0205495
R1829 VSS.n301 VSS.n300 0.0191877
R1830 VSS.n365 VSS 0.01778
R1831 VSS.n354 VSS 0.0163717
R1832 VSS VSS.n203 0.0135645
R1833 VSS.n398 VSS 0.0103671
R1834 VSS VSS.n183 0.00935583
R1835 VSS.n115 VSS.n113 0.00861623
R1836 VSS.n204 VSS 0.00654839
R1837 VSS.n390 VSS.n389 0.00633057
R1838 VSS.n382 VSS.n19 0.00627154
R1839 VSS VSS.n162 0.00545413
R1840 VSS VSS.n165 0.00545413
R1841 VSS.n168 VSS 0.00545413
R1842 VSS.n62 VSS 0.00545413
R1843 VSS.n60 VSS 0.00545413
R1844 VSS.n58 VSS 0.00545413
R1845 VSS.n153 VSS 0.00545413
R1846 VSS VSS.n151 0.00545413
R1847 VSS VSS.n149 0.00545413
R1848 VSS.n130 VSS 0.00545413
R1849 VSS.n132 VSS 0.00545413
R1850 VSS.n138 VSS 0.00545413
R1851 VSS.n375 VSS 0.00545413
R1852 VSS VSS.n373 0.00545413
R1853 VSS VSS.n371 0.00545413
R1854 VSS.n220 VSS 0.00545413
R1855 VSS.n222 VSS 0.00545413
R1856 VSS.n224 VSS 0.00545413
R1857 VSS VSS.n410 0.00545413
R1858 VSS VSS.n408 0.00545413
R1859 VSS VSS.n406 0.00545413
R1860 VSS.n290 VSS 0.00427778
R1861 VSS.n346 VSS.n345 0.00410721
R1862 VSS.n159 VSS 0.00380275
R1863 VSS VSS.n64 0.00380275
R1864 VSS.n147 VSS 0.00380275
R1865 VSS.n136 VSS 0.00380275
R1866 VSS.n369 VSS 0.00380275
R1867 VSS.n226 VSS 0.00380275
R1868 VSS.n240 VSS 0.00380275
R1869 VSS.n404 VSS 0.00380275
R1870 VSS.n286 VSS 0.00352521
R1871 VSS.n243 VSS 0.00352521
R1872 VSS.n328 VSS 0.0031087
R1873 VSS VSS.n340 0.0031087
R1874 VSS VSS.n318 0.00309615
R1875 VSS.n320 VSS 0.00309615
R1876 VSS.n189 VSS 0.00286842
R1877 VSS.n188 VSS 0.00286842
R1878 VSS.n183 VSS 0.00279299
R1879 VSS.n182 VSS 0.00279299
R1880 VSS VSS.n332 0.00223913
R1881 VSS VSS.n330 0.00223913
R1882 VSS.n312 VSS 0.00223077
R1883 VSS.n315 VSS 0.00223077
R1884 VSS.n5 VSS 0.00219811
R1885 VSS.n122 VSS 0.00219811
R1886 VSS VSS.n175 0.00219811
R1887 VSS.n127 VSS 0.00219811
R1888 VSS.n336 VSS 0.00219811
R1889 VSS.n271 VSS 0.00219811
R1890 VSS.n237 VSS 0.00219811
R1891 VSS.n248 VSS 0.0020562
R1892 VSS.n251 VSS 0.0020562
R1893 VSS VSS.n268 0.0020562
R1894 VSS VSS.n266 0.0020562
R1895 VSS VSS.n246 0.00191732
R1896 VSS VSS.n73 0.00168421
R1897 VSS.n94 VSS 0.00168421
R1898 VSS.n83 VSS 0.00168421
R1899 VSS.n99 VSS 0.0016465
R1900 VSS.n86 VSS 0.0016465
R1901 VSS VSS.n353 0.00158216
R1902 VSS VSS.n351 0.00158216
R1903 VSS.n107 VSS 0.00158216
R1904 VSS.n110 VSS 0.00158216
R1905 VSS VSS.n364 0.00158
R1906 VSS VSS.n362 0.00158
R1907 VSS.n253 VSS 0.00153746
R1908 VSS VSS.n256 0.00153746
R1909 VSS.n264 VSS 0.00153746
R1910 VSS.n262 VSS 0.00153746
R1911 VSS.n279 VSS 0.00132569
R1912 VSS VSS.n282 0.00132569
R1913 VSS VSS.n284 0.00132569
R1914 VSS VSS.n294 0.00132569
R1915 VSS VSS.n296 0.00132569
R1916 VSS VSS.n298 0.00124689
R1917 VSS VSS.n381 0.0012438
R1918 VSS.n348 VSS 0.00122144
R1919 VSS.n345 VSS 0.00122144
R1920 VSS VSS.n115 0.00122144
R1921 VSS.n117 VSS 0.00122144
R1922 VSS.n360 VSS 0.00122
R1923 VSS.n357 VSS 0.00122
R1924 VSS.n303 VSS 0.00118965
R1925 VSS.n198 VSS 0.00111785
R1926 VSS.n192 VSS 0.00111785
R1927 VSS.n186 VSS 0.00111785
R1928 VSS.n180 VSS 0.00111785
R1929 VSS VSS.n342 0.00111644
R1930 VSS.n204 VSS 0.000983871
R1931 VSS VSS.n201 0.000954545
R1932 VSS.n76 VSS 0.000945545
R1933 VSS.n80 VSS 0.000945545
R1934 VSS VSS.n289 0.000944444
R1935 VSS VSS.n400 0.000799003
R1936 VSS VSS.n397 0.000799003
R1937 VSS VSS.n395 0.000799003
R1938 VSS VSS.n393 0.000799003
R1939 VSS VSS.n391 0.000799003
R1940 VSS.n16 VSS 0.000799003
R1941 VSS.n18 VSS 0.000799003
R1942 VSS.n384 VSS 0.000799003
R1943 VSS.n198 VSS.n75 0.00070595
R1944 VSS.n197 VSS.n196 0.00070595
R1945 VSS.n195 VSS.n194 0.00070595
R1946 VSS.n193 VSS.n192 0.00070595
R1947 VSS.n191 VSS.n190 0.00070595
R1948 VSS.n189 VSS.n188 0.00070595
R1949 VSS.n187 VSS.n186 0.00070595
R1950 VSS.n185 VSS.n184 0.00070595
R1951 VSS.n183 VSS.n182 0.00070595
R1952 VSS.n181 VSS.n180 0.00070595
R1953 VSS.n179 VSS.n178 0.00070595
R1954 CLK_div_31_mag_0.Q3.n2 CLK_div_31_mag_0.Q3.t2 36.935
R1955 CLK_div_31_mag_0.Q3.n9 CLK_div_31_mag_0.Q3.t13 36.935
R1956 CLK_div_31_mag_0.Q3.n8 CLK_div_31_mag_0.Q3.t7 36.935
R1957 CLK_div_31_mag_0.Q3.n3 CLK_div_31_mag_0.Q3.t9 31.528
R1958 CLK_div_31_mag_0.Q3.n5 CLK_div_31_mag_0.Q3.t14 31.528
R1959 CLK_div_31_mag_0.Q3.n6 CLK_div_31_mag_0.Q3.t4 31.528
R1960 CLK_div_31_mag_0.Q3.n11 CLK_div_31_mag_0.Q3.t6 25.5364
R1961 CLK_div_31_mag_0.Q3.n2 CLK_div_31_mag_0.Q3.t15 18.1962
R1962 CLK_div_31_mag_0.Q3.n9 CLK_div_31_mag_0.Q3.t11 18.1962
R1963 CLK_div_31_mag_0.Q3.n8 CLK_div_31_mag_0.Q3.t3 18.1962
R1964 CLK_div_31_mag_0.Q3.n3 CLK_div_31_mag_0.Q3.t5 15.3826
R1965 CLK_div_31_mag_0.Q3.n5 CLK_div_31_mag_0.Q3.t10 15.3826
R1966 CLK_div_31_mag_0.Q3.n6 CLK_div_31_mag_0.Q3.t8 15.3826
R1967 CLK_div_31_mag_0.Q3.n11 CLK_div_31_mag_0.Q3.t12 14.0749
R1968 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q3.n6 7.63631
R1969 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q3.n3 6.86134
R1970 CLK_div_31_mag_0.Q3.n7 CLK_div_31_mag_0.Q3 6.23913
R1971 CLK_div_31_mag_0.Q3.n1 CLK_div_31_mag_0.Q3.n5 8.03067
R1972 CLK_div_31_mag_0.Q3.n4 CLK_div_31_mag_0.Q3 5.01116
R1973 CLK_div_31_mag_0.Q3.n0 CLK_div_31_mag_0.Q3 4.5005
R1974 CLK_div_31_mag_0.Q3.n10 CLK_div_31_mag_0.Q3 3.25197
R1975 CLK_div_31_mag_0.Q3.n7 CLK_div_31_mag_0.Q3 2.91397
R1976 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q3.n1 2.52047
R1977 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q3.n12 2.3025
R1978 CLK_div_31_mag_0.Q3.n10 CLK_div_31_mag_0.Q3 2.25107
R1979 CLK_div_31_mag_0.Q3.n1 CLK_div_31_mag_0.Q3 2.24713
R1980 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q3.n2 2.13398
R1981 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q3.n8 2.12175
R1982 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q3.n9 2.12075
R1983 CLK_div_31_mag_0.Q3.n0 CLK_div_31_mag_0.Q3.n7 1.69271
R1984 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q3.n11 1.42706
R1985 CLK_div_31_mag_0.Q3.n12 CLK_div_31_mag_0.Q3.n4 1.32654
R1986 CLK_div_31_mag_0.Q3.n4 CLK_div_31_mag_0.Q3 1.12056
R1987 CLK_div_31_mag_0.Q3.n0 CLK_div_31_mag_0.Q3.n10 1.02402
R1988 CLK_div_31_mag_0.Q3.n12 CLK_div_31_mag_0.Q3.n0 0.557773
R1989 CLK_div_31_mag_0.Q1.n4 CLK_div_31_mag_0.Q1.t8 36.935
R1990 CLK_div_31_mag_0.Q1.n13 CLK_div_31_mag_0.Q1.t16 36.935
R1991 CLK_div_31_mag_0.Q1.n12 CLK_div_31_mag_0.Q1.t15 36.935
R1992 CLK_div_31_mag_0.Q1.n5 CLK_div_31_mag_0.Q1.t9 31.528
R1993 CLK_div_31_mag_0.Q1.n6 CLK_div_31_mag_0.Q1.t12 31.528
R1994 CLK_div_31_mag_0.Q1.n9 CLK_div_31_mag_0.Q1.t13 31.4332
R1995 CLK_div_31_mag_0.Q1.n11 CLK_div_31_mag_0.Q1.t5 25.5364
R1996 CLK_div_31_mag_0.Q1.n4 CLK_div_31_mag_0.Q1.t7 18.1962
R1997 CLK_div_31_mag_0.Q1.n13 CLK_div_31_mag_0.Q1.t4 18.1962
R1998 CLK_div_31_mag_0.Q1.n12 CLK_div_31_mag_0.Q1.t14 18.1962
R1999 CLK_div_31_mag_0.Q1.n9 CLK_div_31_mag_0.Q1.t11 15.3826
R2000 CLK_div_31_mag_0.Q1.n5 CLK_div_31_mag_0.Q1.t3 15.3826
R2001 CLK_div_31_mag_0.Q1.n6 CLK_div_31_mag_0.Q1.t10 15.3826
R2002 CLK_div_31_mag_0.Q1.n11 CLK_div_31_mag_0.Q1.t6 14.0749
R2003 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n5 7.63417
R2004 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n6 7.62076
R2005 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.t2 7.09905
R2006 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n9 6.86029
R2007 CLK_div_31_mag_0.Q1.n8 CLK_div_31_mag_0.Q1.n7 6.65668
R2008 CLK_div_31_mag_0.Q1.n7 CLK_div_31_mag_0.Q1 5.46205
R2009 CLK_div_31_mag_0.Q1.n7 CLK_div_31_mag_0.Q1 4.73586
R2010 CLK_div_31_mag_0.Q1.n10 CLK_div_31_mag_0.Q1.n8 3.41968
R2011 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n3 3.25053
R2012 CLK_div_31_mag_0.Q1.n3 CLK_div_31_mag_0.Q1.t0 2.2755
R2013 CLK_div_31_mag_0.Q1.n3 CLK_div_31_mag_0.Q1.n2 2.2755
R2014 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n4 2.13459
R2015 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n13 2.13151
R2016 CLK_div_31_mag_0.Q1.n1 CLK_div_31_mag_0.Q1 2.63808
R2017 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n12 2.13042
R2018 CLK_div_31_mag_0.Q1.n8 CLK_div_31_mag_0.Q1 1.5916
R2019 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n10 1.49033
R2020 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n11 1.43689
R2021 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n0 1.22411
R2022 CLK_div_31_mag_0.Q1.n10 CLK_div_31_mag_0.Q1 1.12067
R2023 CLK_div_31_mag_0.Q1.n0 CLK_div_31_mag_0.Q1 1.12013
R2024 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q1.n1 1.11863
R2025 CLK_div_31_mag_0.Q1.n0 CLK_div_31_mag_0.Q1.n1 0.927577
R2026 CLK_div_31_mag_0.Q4.n3 CLK_div_31_mag_0.Q4.t4 40.2519
R2027 CLK_div_31_mag_0.Q4.n0 CLK_div_31_mag_0.Q4.t3 36.935
R2028 CLK_div_31_mag_0.Q4.n4 CLK_div_31_mag_0.Q4.t5 31.528
R2029 CLK_div_31_mag_0.Q4.n1 CLK_div_31_mag_0.Q4.t7 31.528
R2030 CLK_div_31_mag_0.Q4.n0 CLK_div_31_mag_0.Q4.t8 18.1962
R2031 CLK_div_31_mag_0.Q4.n3 CLK_div_31_mag_0.Q4.t9 15.3826
R2032 CLK_div_31_mag_0.Q4.n4 CLK_div_31_mag_0.Q4.t2 15.3826
R2033 CLK_div_31_mag_0.Q4.n1 CLK_div_31_mag_0.Q4.t6 15.3826
R2034 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Q4.n4 7.63442
R2035 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Q4.n1 6.86134
R2036 CLK_div_31_mag_0.Q4.n2 CLK_div_31_mag_0.Q4 5.01116
R2037 CLK_div_31_mag_0.Q4.n5 CLK_div_31_mag_0.Q4 3.11241
R2038 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Q4.n6 2.25871
R2039 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Q4.n0 2.13398
R2040 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Q4.n3 2.12278
R2041 CLK_div_31_mag_0.Q4.n5 CLK_div_31_mag_0.Q4 2.10026
R2042 CLK_div_31_mag_0.Q4.n6 CLK_div_31_mag_0.Q4.n2 1.37588
R2043 CLK_div_31_mag_0.Q4.n6 CLK_div_31_mag_0.Q4.n5 1.26898
R2044 CLK_div_31_mag_0.Q4.n2 CLK_div_31_mag_0.Q4 1.12056
R2045 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 37.1986
R2046 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 31.528
R2047 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 30.5184
R2048 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 24.7029
R2049 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 17.6614
R2050 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 15.3826
R2051 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 12.0843
R2052 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 9.86691
R2053 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R2054 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 2.99416
R2055 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.t1 2.2755
R2056 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2755
R2057 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 2.2505
R2058 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.24173
R2059 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.93723
R2060 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n2 1.81225
R2061 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.43709
R2062 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n1 0.281955
R2063 RST.n35 RST.t9 37.1991
R2064 RST.n30 RST.t8 36.935
R2065 RST.n21 RST.t6 36.935
R2066 RST.n26 RST.t14 36.935
R2067 RST.n0 RST.t11 36.935
R2068 RST.n12 RST.t4 36.935
R2069 RST.n39 RST.t2 36.935
R2070 RST.n30 RST.t5 18.1962
R2071 RST.n21 RST.t13 18.1962
R2072 RST.n26 RST.t12 18.1962
R2073 RST.n0 RST.t10 18.1962
R2074 RST.n12 RST.t3 18.1962
R2075 RST.n39 RST.t15 18.1962
R2076 RST.n35 RST.t7 17.66
R2077 RST.n54 RST.n45 11.4652
R2078 RST.n50 RST.n48 9.33985
R2079 RST.n55 RST.n54 6.23435
R2080 RST.n45 RST.n38 5.63145
R2081 RST.n28 RST.n27 5.42044
R2082 RST.n50 RST.n49 5.17836
R2083 RST.n57 RST.n56 4.51909
R2084 RST.n14 RST.n10 4.5005
R2085 RST.n14 RST.n13 4.5005
R2086 RST.n16 RST.n15 4.5005
R2087 RST.n44 RST.n43 4.5005
R2088 RST.n45 RST.n44 3.78663
R2089 RST.n32 RST.n31 3.49993
R2090 RST.n56 RST.n55 2.78304
R2091 RST.n51 RST 2.27453
R2092 RST.n41 RST.n40 2.25731
R2093 RST.n5 RST.n3 2.2505
R2094 RST.n17 RST.n16 2.2505
R2095 RST.n38 RST.n37 2.24157
R2096 RST.n27 RST.n26 2.15059
R2097 RST.n31 RST.n30 2.14848
R2098 RST.n41 RST.n39 2.12457
R2099 RST.n1 RST.n0 2.1224
R2100 RST.n13 RST.n12 2.12207
R2101 RST.n22 RST.n21 2.1217
R2102 RST.n55 RST.n20 2.06221
R2103 RST.n55 RST.n32 1.79221
R2104 RST.n20 RST.n7 1.78161
R2105 RST.n32 RST.n29 1.72354
R2106 RST.n20 RST.n19 1.53272
R2107 RST.n52 RST.n51 1.50509
R2108 RST.n36 RST.n35 1.41552
R2109 RST.n29 RST.n25 1.1266
R2110 RST.n7 RST.n6 0.940487
R2111 RST RST.n57 0.938927
R2112 RST.n24 RST.n23 0.898026
R2113 RST.n46 RST 0.723675
R2114 RST.n54 RST.n53 0.473577
R2115 RST RST.n50 0.109973
R2116 RST.n42 RST 0.0593097
R2117 RST.n31 RST 0.0563307
R2118 RST.n27 RST 0.0558741
R2119 RST.n23 RST 0.0553557
R2120 RST.n34 RST 0.0410354
R2121 RST.n2 RST 0.0377414
R2122 RST.n3 RST.n2 0.0361897
R2123 RST.n37 RST.n34 0.0361897
R2124 RST.n10 RST 0.0348285
R2125 RST.n44 RST 0.0293
R2126 RST.n23 RST.n22 0.0275188
R2127 RST.n53 RST.n52 0.0274231
R2128 RST.n5 RST.n4 0.0267025
R2129 RST.n14 RST.n11 0.0255
R2130 RST.n9 RST.n8 0.0235
R2131 RST.n38 RST.n33 0.0230258
R2132 RST RST.n56 0.019087
R2133 RST.n43 RST.n42 0.0187743
R2134 RST.n29 RST.n28 0.0175868
R2135 RST.n52 RST.n46 0.0140977
R2136 RST.n3 RST.n1 0.00515517
R2137 RST.n37 RST.n36 0.00515517
R2138 RST.n25 RST.n24 0.00494444
R2139 RST.n6 RST.n5 0.00372575
R2140 RST.n43 RST.n41 0.00333412
R2141 RST.n51 RST.n47 0.00217441
R2142 RST.n40 RST 0.0017
R2143 RST.n16 RST.n9 0.0015
R2144 RST.n16 RST.n14 0.0015
R2145 RST.n19 RST.n18 0.0015
R2146 RST.n18 RST.n17 0.0015
R2147 CLK_div_31_mag_0.JK_FF_mag_0.QB.n2 CLK_div_31_mag_0.JK_FF_mag_0.QB.t4 37.1981
R2148 CLK_div_31_mag_0.JK_FF_mag_0.QB.n1 CLK_div_31_mag_0.JK_FF_mag_0.QB.t3 31.528
R2149 CLK_div_31_mag_0.JK_FF_mag_0.QB.n2 CLK_div_31_mag_0.JK_FF_mag_0.QB.t6 17.6611
R2150 CLK_div_31_mag_0.JK_FF_mag_0.QB.n1 CLK_div_31_mag_0.JK_FF_mag_0.QB.t5 15.3826
R2151 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_0.QB.n1 7.62751
R2152 CLK_div_31_mag_0.JK_FF_mag_0.QB.n3 CLK_div_31_mag_0.JK_FF_mag_0.QB 6.09789
R2153 CLK_div_31_mag_0.JK_FF_mag_0.QB.n0 CLK_div_31_mag_0.JK_FF_mag_0.QB.n5 2.99416
R2154 CLK_div_31_mag_0.JK_FF_mag_0.QB.n3 CLK_div_31_mag_0.JK_FF_mag_0.QB 2.67866
R2155 CLK_div_31_mag_0.JK_FF_mag_0.QB.n5 CLK_div_31_mag_0.JK_FF_mag_0.QB.t0 2.2755
R2156 CLK_div_31_mag_0.JK_FF_mag_0.QB.n5 CLK_div_31_mag_0.JK_FF_mag_0.QB.n4 2.2755
R2157 CLK_div_31_mag_0.JK_FF_mag_0.QB.n0 CLK_div_31_mag_0.JK_FF_mag_0.QB.n3 2.2505
R2158 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_0.QB.n2 1.43706
R2159 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_0.QB.n0 0.281955
R2160 CLK.n8 CLK.t3 36.935
R2161 CLK.n12 CLK.t7 36.935
R2162 CLK.n0 CLK.t4 31.528
R2163 CLK.n20 CLK.t0 25.4744
R2164 CLK.n8 CLK.t5 18.1962
R2165 CLK.n12 CLK.t6 18.1962
R2166 CLK.n0 CLK.t1 15.3826
R2167 CLK.n20 CLK.t2 14.1417
R2168 CLK.n1 CLK.n0 7.62171
R2169 CLK.n32 CLK.n31 6.57848
R2170 CLK.n3 CLK.n2 6.33303
R2171 CLK.n2 CLK.n1 5.0581
R2172 CLK.n33 CLK.n32 4.53391
R2173 CLK.n28 CLK.n7 2.26042
R2174 CLK.n19 CLK.n11 2.25107
R2175 CLK.n7 CLK.n6 2.2505
R2176 CLK.n23 CLK.n22 2.24319
R2177 CLK.n27 CLK.n26 2.24244
R2178 CLK.n15 CLK.n12 2.12464
R2179 CLK.n9 CLK.n8 2.12188
R2180 CLK.n18 CLK.n17 1.71671
R2181 CLK.n16 CLK.n15 1.50503
R2182 CLK.n21 CLK.n20 1.42118
R2183 CLK.n31 CLK.n30 1.32117
R2184 CLK.n23 CLK.n19 0.964895
R2185 CLK CLK.n33 0.916495
R2186 CLK.n31 CLK.n3 0.158593
R2187 CLK.n6 CLK.n5 0.09875
R2188 CLK.n6 CLK 0.04775
R2189 CLK.n10 CLK 0.0457995
R2190 CLK.n13 CLK 0.0457995
R2191 CLK.n26 CLK.n25 0.0403734
R2192 CLK.n17 CLK.n16 0.0386356
R2193 CLK.n11 CLK.n10 0.0377414
R2194 CLK.n14 CLK.n13 0.0377414
R2195 CLK.n25 CLK.n24 0.03466
R2196 CLK CLK.n32 0.0339132
R2197 CLK.n30 CLK.n29 0.0328596
R2198 CLK.n1 CLK 0.0316785
R2199 CLK.n24 CLK.n23 0.0207183
R2200 CLK.n28 CLK.n27 0.0181256
R2201 CLK.n19 CLK.n18 0.0122182
R2202 CLK.n2 CLK 0.0095
R2203 CLK.n3 CLK 0.00469786
R2204 CLK.n11 CLK.n9 0.00360345
R2205 CLK.n29 CLK.n4 0.00286842
R2206 CLK.n15 CLK.n14 0.00203726
R2207 CLK.n22 CLK.n21 0.00175
R2208 CLK.n29 CLK.n28 0.00151124
R2209 Vdiv93.n2 Vdiv93.n1 9.33985
R2210 Vdiv93.n2 Vdiv93.n0 5.17836
R2211 Vdiv93 Vdiv93.n2 0.0749828
C0 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.CLK 0.298f
C1 a_15342_208# CLK_div_3_mag_0.Q1 0.00789f
C2 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 7.03e-21
C3 a_18199_208# CLK_div_3_mag_0.CLK 0.00117f
C4 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q3 0.983f
C5 VDD CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.744f
C6 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 0.111f
C7 a_7506_3203# CLK_div_31_mag_0.Q2 0.00692f
C8 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00112f
C9 CLK_div_31_mag_0.JK_FF_mag_1.QB a_7095_1457# 1.72e-20
C10 VDD CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.471f
C11 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00169f
C12 CLK_div_3_mag_0.JK_FF_mag_1.K VDD 2.63f
C13 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_2528_4227# 0.0202f
C14 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.16f
C15 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.or_2_mag_0.IN2 5.32e-19
C16 CLK a_5428_4226# 0.00539f
C17 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.Q0 0.00335f
C18 a_1699_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C19 CLK_div_31_mag_0.Q0 a_5422_3129# 4.21e-19
C20 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_8383_1501# 0.011f
C21 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_20057_1349# 0.00118f
C22 a_7095_1457# RST 0.00185f
C23 a_2833_1493# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.21e-19
C24 a_4140_4226# RST 8.06e-19
C25 a_17194_252# RST 0.00114f
C26 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C27 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.00668f
C28 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C29 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2362_3130# 3.87e-20
C30 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C31 a_19647_252# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C32 a_1141_1449# RST 7.68e-19
C33 a_15182_208# CLK_div_3_mag_0.Q1 0.00335f
C34 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.17e-19
C35 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.0357f
C36 a_7973_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 2.88e-20
C37 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C38 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C39 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C40 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN RST 0.015f
C41 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.16f
C42 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.75e-19
C43 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 3.58e-19
C44 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00103f
C45 CLK CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00254f
C46 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q2 0.0264f
C47 CLK_div_3_mag_0.JK_FF_mag_1.QB a_15912_1349# 3.33e-19
C48 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.01f
C49 a_4017_361# RST 0.00189f
C50 a_7249_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 1.5e-20
C51 a_2833_1493# VDD 3.56e-19
C52 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 4.21e-20
C53 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_2368_4227# 0.0731f
C54 CLK a_4864_4226# 0.00148f
C55 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C56 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN Vdiv93 0.129f
C57 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_31_mag_0.Q2 3.91e-20
C58 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_19493_1349# 0.011f
C59 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C60 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_7819_1501# 1.43e-19
C61 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_0.QB 0.199f
C62 a_3576_4226# RST 8.24e-19
C63 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.Q2 2.39f
C64 a_16630_252# RST 0.00164f
C65 a_7813_360# CLK_div_31_mag_0.Q4 0.0102f
C66 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.127f
C67 VDD CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.655f
C68 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD 0.802f
C69 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q1 2.08f
C70 a_2522_3130# RST 0.00264f
C71 VDD CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C72 a_2423_396# CLK_div_31_mag_0.JK_FF_mag_0.QB 0.00964f
C73 a_10367_3208# RST 9.29e-19
C74 CLK a_10368_3965# 0.00479f
C75 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_17040_1349# 4.52e-20
C76 CLK_div_3_mag_0.JK_FF_mag_1.QB a_15348_1305# 0.00392f
C77 CLK_div_31_mag_0.Q4 a_7255_1457# 2.79e-20
C78 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.23e-19
C79 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_1804_4227# 9.1e-19
C80 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VDD 0.519f
C81 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_0.QB 3.48e-19
C82 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C83 CLK_div_31_mag_0.Q0 a_4294_3129# 6.14e-21
C84 VDD CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.749f
C85 CLK a_4704_4226# 0.00145f
C86 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_18929_1349# 1.43e-19
C87 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_7255_1457# 0.00119f
C88 a_16066_208# RST 0.00228f
C89 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0877f
C90 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00103f
C91 a_670_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C92 a_4183_1458# CLK_div_31_mag_0.JK_FF_mag_0.QB 1.07e-20
C93 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0725f
C94 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_3.QB 0.0592f
C95 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN RST 0.0388f
C96 a_4017_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C97 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C98 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C99 a_9403_3219# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 8.97e-21
C100 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_3.QB 0.103f
C101 a_2987_396# CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C102 a_2269_1493# CLK_div_31_mag_0.JK_FF_mag_0.QB 2.96e-19
C103 a_2362_3130# RST 0.00204f
C104 VDD a_11989_2561# 0.165f
C105 a_7973_360# CLK_div_31_mag_0.JK_FF_mag_4.QB 0.00696f
C106 a_16630_252# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C107 CLK a_9404_3954# 7.37e-19
C108 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C109 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 RST 0.0188f
C110 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN a_10368_3965# 0.069f
C111 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.11e-19
C112 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT RST 0.0981f
C113 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.61e-20
C114 CLK_div_3_mag_0.Q0 RST 0.0447f
C115 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_3.QB 9.89e-20
C116 a_4177_361# CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C117 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 6.04e-20
C118 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_1644_4227# 2.88e-20
C119 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD 0.746f
C120 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_31_mag_0.or_2_mag_0.IN1 2.97e-19
C121 CLK a_4140_4226# 0.00178f
C122 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_31_mag_0.Q2 2.93e-20
C123 CLK_div_31_mag_0.Q0 a_3730_3129# 0.069f
C124 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.CLK 0.235f
C125 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_18365_1305# 0.00119f
C126 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN RST 0.00968f
C127 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.Q0 0.149f
C128 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 RST 0.00252f
C129 a_15906_208# RST 0.00187f
C130 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q2 0.892f
C131 a_4023_1458# CLK_div_31_mag_0.JK_FF_mag_0.QB 1.4e-20
C132 a_5875_1502# CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C133 a_2423_396# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C134 VDD CLK_div_3_mag_0.Q1 2.52f
C135 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN RST 0.00661f
C136 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.CLK 0.0215f
C137 a_975_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C138 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00579f
C139 a_1705_1493# CLK_div_31_mag_0.JK_FF_mag_0.QB 3.33e-19
C140 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q2 0.671f
C141 a_1798_3130# RST 6.28e-19
C142 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK 8.46e-19
C143 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C144 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C145 a_16066_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C146 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.12f
C147 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 0.519f
C148 CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 3.21e-19
C149 a_4741_361# CLK_div_31_mag_0.JK_FF_mag_1.QB 0.00695f
C150 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0016f
C151 CLK a_3576_4226# 0.00178f
C152 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN RST 0.0227f
C153 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.Q3 0.102f
C154 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.128f
C155 a_2269_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C156 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C157 a_4741_361# RST 0.00171f
C158 a_7973_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.0733f
C159 a_15342_208# RST 0.00218f
C160 a_18205_1305# a_18365_1305# 0.0504f
C161 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C162 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.298f
C163 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q1 0.363f
C164 a_8452_3208# RST 3.66e-19
C165 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_5588_4226# 1.17e-20
C166 a_1141_1449# CLK_div_31_mag_0.JK_FF_mag_0.QB 0.00392f
C167 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.305f
C168 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT RST 0.0231f
C169 a_15342_208# CLK_div_3_mag_0.CLK 0.00164f
C170 a_10367_3208# CLK 2.43e-19
C171 a_1234_3130# RST 6.04e-19
C172 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C173 CLK_div_31_mag_0.JK_FF_mag_3.QB VDD 0.915f
C174 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C175 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00113f
C176 a_8537_404# CLK_div_31_mag_0.Q4 0.00859f
C177 CLK_div_31_mag_0.and_5_mag_0.VOUT VDD 1.03f
C178 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0957f
C179 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 4.92e-19
C180 a_3730_3129# CLK_div_31_mag_0.Q2 5.1e-19
C181 CLK_div_3_mag_0.Q0 Vdiv93 0.00953f
C182 a_15906_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C183 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.314f
C184 a_8537_404# CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.0036f
C185 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_31_mag_0.Q4 2.35e-19
C186 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0822f
C187 a_1705_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C188 a_7813_360# a_7973_360# 0.0504f
C189 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.0123f
C190 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.652f
C191 a_5422_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00119f
C192 a_15182_208# RST 0.00218f
C193 a_981_1449# a_1141_1449# 0.0504f
C194 a_4858_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0697f
C195 a_11989_2561# CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C196 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.Q1 0.0177f
C197 a_15182_208# CLK_div_3_mag_0.CLK 0.00117f
C198 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_1.QB 3.09e-19
C199 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 4.92e-21
C200 a_4741_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C201 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_2.QB 0.198f
C202 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.28e-19
C203 a_7507_3970# VDD 3.14e-19
C204 a_15342_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C205 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_31_mag_0.and_5_mag_0.VOUT 0.0974f
C206 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C207 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 RST 0.02f
C208 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C209 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 0.0275f
C210 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.28f
C211 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 7.98e-19
C212 a_4747_1502# CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.61e-20
C213 CLK_div_31_mag_0.JK_FF_mag_2.QB a_1804_4227# 0.00695f
C214 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT RST 0.0508f
C215 a_9101_404# CLK_div_31_mag_0.JK_FF_mag_4.QB 0.0811f
C216 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.9e-21
C217 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_5428_4226# 1.5e-20
C218 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.0104f
C219 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 0.338f
C220 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN VDD 0.418f
C221 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.02e-20
C222 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 0.00846f
C223 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0385f
C224 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00237f
C225 a_4858_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.43e-19
C226 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00335f
C227 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0126f
C228 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C229 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C230 a_4294_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0059f
C231 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 RST 0.2f
C232 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 2.62e-19
C233 CLK_div_31_mag_0.Q1 a_975_352# 0.00117f
C234 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 5.32e-19
C235 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 8.18e-19
C236 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.Q3 0.0124f
C237 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C238 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_1644_4227# 8.64e-19
C239 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 2.02e-19
C240 a_15182_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C241 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00119f
C242 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.and_5_mag_0.VOUT 0.00384f
C243 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_5875_1502# 0.00372f
C244 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.129f
C245 a_1699_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C246 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.00832f
C247 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.00382f
C248 CLK_div_31_mag_0.Q1 a_2528_4227# 0.0122f
C249 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 6.85e-19
C250 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_0.QB 0.0592f
C251 CLK_div_31_mag_0.JK_FF_mag_2.QB a_1644_4227# 0.00696f
C252 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_4864_4226# 0.0203f
C253 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_4140_4226# 0.069f
C254 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_670_3130# 0.00372f
C255 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0218f
C256 CLK_div_31_mag_0.Q4 a_8452_3208# 3.11e-21
C257 CLK_div_31_mag_0.Q0 a_2528_4227# 0.00144f
C258 a_5465_405# CLK_div_31_mag_0.JK_FF_mag_1.QB 0.00964f
C259 a_4294_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.011f
C260 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.00183f
C261 RST CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.061f
C262 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.768f
C263 a_8452_3208# CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 3.66e-20
C264 CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4e-20
C265 CLK a_1234_3130# 3.7e-19
C266 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.Q3 0.235f
C267 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.112f
C268 a_5465_405# RST 9.62e-19
C269 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_2.QB 0.25f
C270 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.Q3 0.0246f
C271 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.128f
C272 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C273 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_5311_1502# 0.069f
C274 CLK_div_31_mag_0.JK_FF_mag_1.QB VDD 0.915f
C275 CLK_div_31_mag_0.Q1 a_2368_4227# 0.0151f
C276 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00314f
C277 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_4704_4226# 0.0733f
C278 CLK_div_31_mag_0.JK_FF_mag_2.QB a_1080_4227# 0.00964f
C279 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.Q0 0.0635f
C280 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2833_1493# 0.00118f
C281 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_3576_4226# 0.00372f
C282 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 RST 0.00889f
C283 VDD a_516_4227# 3.14e-19
C284 a_5422_3129# CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.42e-20
C285 VDD RST 5.36f
C286 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0124f
C287 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.Q2 0.00542f
C288 CLK_div_31_mag_0.Q0 a_2368_4227# 0.00169f
C289 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 RST 8.23e-19
C290 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C291 a_3730_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C292 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 0.00617f
C293 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q0 7.24e-19
C294 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 0.107f
C295 VDD CLK_div_3_mag_0.CLK 2.94f
C296 a_975_352# CLK_div_31_mag_0.Q2 0.00335f
C297 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C298 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C299 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C300 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_0.QB 3.01e-20
C301 a_5875_1502# CLK_div_31_mag_0.Q3 0.069f
C302 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK 3.92e-20
C303 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C304 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C305 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.101f
C306 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 4.29e-20
C307 CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.79e-20
C308 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.or_2_mag_0.IN2 4.52e-20
C309 a_1234_3130# CLK_div_31_mag_0.JK_FF_mag_0.QB 5e-20
C310 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 8.36e-19
C311 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK 0.263f
C312 a_7089_360# CLK_div_31_mag_0.Q3 0.00182f
C313 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_31_mag_0.Q2 0.28f
C314 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VDD 0.39f
C315 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 2.08e-19
C316 CLK_div_31_mag_0.Q1 a_1804_4227# 0.0102f
C317 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT RST 0.0118f
C318 a_5465_405# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C319 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_4140_4226# 0.00378f
C320 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 2.06e-19
C321 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 6.95e-19
C322 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.00102f
C323 CLK_div_3_mag_0.JK_FF_mag_1.K RST 0.254f
C324 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.Q3 0.00525f
C325 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.129f
C326 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.00168f
C327 a_1798_3130# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 5e-20
C328 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C329 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.343f
C330 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0983f
C331 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.CLK 2.12f
C332 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD 0.998f
C333 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD 1f
C334 CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 1.56e-19
C335 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.Q3 0.308f
C336 a_5311_1502# CLK_div_31_mag_0.Q3 6.03e-21
C337 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.Q1 6.7e-19
C338 a_4017_361# a_4177_361# 0.0504f
C339 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_19493_1349# 4.52e-20
C340 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 a_10368_3965# 0.00347f
C341 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN a_11989_2561# 4.15e-20
C342 CLK_div_31_mag_0.Q1 a_1644_4227# 0.0101f
C343 VDD Vdiv93 0.156f
C344 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00122f
C345 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_10367_3208# 8.67e-20
C346 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 RST 0.156f
C347 a_2833_1493# RST 0.00221f
C348 CLK CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C349 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 1.01e-20
C350 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.109f
C351 a_17194_252# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0811f
C352 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK 1.31f
C353 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_16476_1349# 0.0059f
C354 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.QB 0.0592f
C355 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0346f
C356 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 6.2e-19
C357 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.Q2 1.05e-20
C358 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C359 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_18929_1349# 0.0202f
C360 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 a_9404_3954# 8.97e-21
C361 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.116f
C362 CLK_div_31_mag_0.Q4 VDD 3.43f
C363 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 RST 0.206f
C364 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD 0.744f
C365 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT RST 0.0843f
C366 CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN RST 0.0148f
C367 CLK_div_31_mag_0.Q1 a_1080_4227# 0.00859f
C368 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 6.64e-19
C369 CLK VDD 2.59f
C370 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VDD 0.519f
C371 a_2269_1493# CLK_div_31_mag_0.JK_FF_mag_2.QB 5e-20
C372 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN Vdiv93 1e-19
C373 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C374 CLK_div_3_mag_0.JK_FF_mag_1.K Vdiv93 4.46e-19
C375 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.36f
C376 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_31_mag_0.Q4 0.0638f
C377 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 4.73e-19
C378 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.CLK 0.235f
C379 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 VDD 1.22f
C380 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.0622f
C381 CLK_div_3_mag_0.CLK CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.13f
C382 CLK_div_31_mag_0.Q1 a_5588_4226# 0.00613f
C383 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.Q3 8.94e-19
C384 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT RST 0.0859f
C385 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN RST 0.0275f
C386 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.321f
C387 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0502f
C388 a_16630_252# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00964f
C389 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.0388f
C390 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.233f
C391 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_7819_1501# 0.00378f
C392 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_3_mag_0.CLK 1.34e-20
C393 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.75e-19
C394 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_15912_1349# 0.0697f
C395 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00541f
C396 CLK_div_31_mag_0.Q3 a_7819_1501# 6.43e-21
C397 CLK_div_31_mag_0.Q0 a_5588_4226# 0.0117f
C398 a_19647_252# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C399 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C400 a_4183_1458# CLK_div_31_mag_0.Q3 2.79e-20
C401 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_4.QB 9.12e-20
C402 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C403 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 4.09e-19
C404 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.Q2 0.66f
C405 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.23e-19
C406 a_1699_352# CLK_div_31_mag_0.Q2 0.0102f
C407 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.119f
C408 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.VOUT 1.26e-19
C409 a_11989_2561# RST 0.00703f
C410 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_4.QB 6.38e-19
C411 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD 0.427f
C412 VDD CLK_div_31_mag_0.JK_FF_mag_0.QB 0.915f
C413 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.Q2 0.0782f
C414 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT RST 0.0206f
C415 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q0 0.107f
C416 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C417 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_8383_1501# 0.0059f
C418 a_16066_208# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00696f
C419 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_7255_1457# 0.0732f
C420 CLK_div_31_mag_0.Q3 a_7255_1457# 0.00939f
C421 CLK_div_3_mag_0.Q1 RST 0.135f
C422 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C423 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C424 a_5875_1502# CLK_div_31_mag_0.Q2 4.6e-19
C425 CLK_div_31_mag_0.Q1 a_5428_4226# 0.006f
C426 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C427 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_9403_3219# 1.05e-20
C428 a_8452_3208# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 4.18e-21
C429 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.517f
C430 a_20057_1349# CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C431 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.Q1 1.03f
C432 a_9101_404# CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 5.06e-20
C433 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C434 a_1859_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C435 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN RST 0.0185f
C436 a_981_1449# VDD 0.00533f
C437 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_9404_3954# 1.05e-20
C438 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.768f
C439 CLK_div_31_mag_0.Q0 a_5428_4226# 0.016f
C440 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 5.53e-19
C441 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C442 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.77e-19
C443 VDD a_18641_2448# 5.95e-19
C444 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C445 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 2.59e-20
C446 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VDD 0.514f
C447 a_17194_252# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00372f
C448 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.34e-21
C449 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.Q2 0.102f
C450 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_7819_1501# 0.0697f
C451 a_15906_208# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00695f
C452 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_7095_1457# 0.0203f
C453 CLK_div_31_mag_0.Q3 a_9404_3954# 9.22e-21
C454 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.11f
C455 a_2368_4227# a_2528_4227# 0.0504f
C456 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD 0.649f
C457 CLK_div_31_mag_0.Q3 a_7095_1457# 0.0101f
C458 a_2987_396# VDD 3.14e-19
C459 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0495f
C460 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.Q2 2.42e-20
C461 CLK_div_31_mag_0.Q1 a_4864_4226# 9.09e-19
C462 CLK_div_3_mag_0.or_2_mag_0.IN2 a_19614_2684# 8.64e-19
C463 a_981_1449# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C464 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 1.48e-20
C465 CLK_div_31_mag_0.JK_FF_mag_3.QB RST 0.186f
C466 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 6.4e-20
C467 VDD CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.998f
C468 CLK_div_31_mag_0.and_5_mag_0.VOUT RST 0.0374f
C469 a_1135_352# CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C470 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.Q1 0.0343f
C471 CLK_div_31_mag_0.Q0 a_4864_4226# 0.0102f
C472 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 2.91e-19
C473 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.112f
C474 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_8453_3965# 0.069f
C475 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.0836f
C476 CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_3_mag_0.CLK 0.248f
C477 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q3 0.00164f
C478 a_16630_252# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.069f
C479 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 8.93e-21
C480 a_15188_1305# a_15348_1305# 0.0504f
C481 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.198f
C482 a_4017_361# CLK_div_31_mag_0.Q3 0.00335f
C483 a_2833_1493# CLK_div_31_mag_0.JK_FF_mag_0.QB 0.0114f
C484 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_18641_2448# 0.069f
C485 CLK_div_3_mag_0.Q1 Vdiv93 2.53e-19
C486 CLK_div_31_mag_0.Q3 a_8453_3965# 0.00943f
C487 CLK_div_31_mag_0.Q1 a_10368_3965# 2.43e-19
C488 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.64e-19
C489 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 RST 0.143f
C490 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C491 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00975f
C492 CLK_div_31_mag_0.Q4 a_11989_2561# 8.64e-19
C493 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C494 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C495 a_18359_208# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C496 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C497 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.CLK 0.00254f
C498 a_4747_1502# CLK_div_31_mag_0.Q2 6.43e-21
C499 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C500 CLK_div_31_mag_0.Q1 a_4704_4226# 9.09e-19
C501 CLK_div_31_mag_0.Q1 a_1705_1493# 6.43e-21
C502 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.392f
C503 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.038f
C504 CLK_div_31_mag_0.Q0 a_4704_4226# 0.0101f
C505 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 7.87e-19
C506 CLK CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 1.56e-21
C507 a_2423_396# CLK_div_31_mag_0.Q2 0.00859f
C508 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 5.06e-21
C509 a_2362_3130# CLK_div_31_mag_0.JK_FF_mag_2.QB 0.00392f
C510 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 RST 0.129f
C511 a_10367_3208# CLK_div_31_mag_0.Q3 4.35e-19
C512 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.09e-19
C513 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 8.64e-20
C514 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.Q2 5.76e-22
C515 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN RST 0.147f
C516 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.QB 3.48e-19
C517 a_7506_3203# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.91e-21
C518 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_8452_3208# 3.85e-20
C519 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C520 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.CLK 1e-20
C521 CLK_div_31_mag_0.Q1 a_4140_4226# 0.00108f
C522 a_4183_1458# CLK_div_31_mag_0.Q2 0.00939f
C523 a_5465_405# CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.069f
C524 a_1798_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0697f
C525 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.00527f
C526 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.0829f
C527 CLK_div_31_mag_0.Q1 a_1141_1449# 0.00939f
C528 a_2269_1493# CLK_div_31_mag_0.Q2 1.46e-21
C529 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C530 CLK_div_31_mag_0.Q0 a_4140_4226# 0.00859f
C531 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.11f
C532 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_10368_3965# 8.67e-20
C533 a_1798_3130# CLK_div_31_mag_0.JK_FF_mag_2.QB 3.33e-19
C534 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0016f
C535 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.3f
C536 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C537 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_2528_4227# 1.17e-20
C538 a_4741_361# a_4901_361# 0.0504f
C539 VDD CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.391f
C540 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.Q0 0.0655f
C541 a_20057_1349# CLK_div_3_mag_0.Q0 0.069f
C542 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.429f
C543 CLK_div_31_mag_0.Q2 a_10368_3965# 4.35e-19
C544 CLK_div_31_mag_0.Q1 a_8453_3965# 3.11e-21
C545 a_670_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C546 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00113f
C547 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.QB 0.343f
C548 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_19614_2684# 1.4e-19
C549 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C550 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.and_5_mag_0.VOUT 5.03e-20
C551 CLK CLK_div_31_mag_0.JK_FF_mag_3.QB 0.414f
C552 a_4023_1458# CLK_div_31_mag_0.Q2 0.0101f
C553 CLK_div_31_mag_0.Q1 a_3576_4226# 0.00108f
C554 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.75f
C555 CLK CLK_div_31_mag_0.and_5_mag_0.VOUT 0.0102f
C556 CLK_div_31_mag_0.Q0 a_8453_3965# 6.36e-20
C557 a_1234_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0059f
C558 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD 0.998f
C559 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q3 0.0264f
C560 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN a_8947_1501# 6.6e-20
C561 CLK_div_31_mag_0.Q1 a_2522_3130# 4.47e-19
C562 CLK_div_31_mag_0.Q0 a_3576_4226# 0.0157f
C563 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.00185f
C564 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_9404_3954# 0.069f
C565 CLK_div_31_mag_0.JK_FF_mag_1.QB RST 0.221f
C566 a_1234_3130# CLK_div_31_mag_0.JK_FF_mag_2.QB 2.96e-19
C567 CLK_div_31_mag_0.Q1 a_10367_3208# 0.00479f
C568 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_2368_4227# 1.5e-20
C569 a_670_3130# VDD 3.56e-19
C570 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 8.99e-19
C571 CLK_div_31_mag_0.Q0 a_2522_3130# 0.0101f
C572 a_9403_3219# VDD 3.14e-19
C573 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C574 CLK_div_31_mag_0.Q2 a_9404_3954# 0.0193f
C575 a_1644_4227# a_1804_4227# 0.0504f
C576 CLK_div_3_mag_0.CLK RST 0.0548f
C577 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.112f
C578 a_4741_361# CLK_div_31_mag_0.Q3 0.0102f
C579 CLK_div_3_mag_0.Q1 a_18641_2448# 0.01f
C580 CLK a_7507_3970# 2.25e-19
C581 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.VOUT 0.122f
C582 a_8452_3208# CLK_div_31_mag_0.Q3 0.0114f
C583 a_1141_1449# CLK_div_31_mag_0.Q2 2.79e-20
C584 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.122f
C585 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.Q3 8.36e-19
C586 a_9101_404# VDD 3.14e-19
C587 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 0.101f
C588 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.31e-19
C589 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN a_8383_1501# 2.72e-20
C590 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 RST 0.00628f
C591 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 0.00872f
C592 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C593 CLK_div_31_mag_0.Q1 a_2362_3130# 3.43e-19
C594 a_9101_404# CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.00372f
C595 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_8453_3965# 4.56e-21
C596 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_1804_4227# 0.0203f
C597 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD 0.877f
C598 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_1080_4227# 0.069f
C599 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.48e-20
C600 a_4017_361# CLK_div_31_mag_0.Q2 0.00185f
C601 CLK_div_31_mag_0.Q0 a_2362_3130# 0.00939f
C602 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C603 CLK_div_31_mag_0.Q2 a_8453_3965# 0.0114f
C604 a_4901_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C605 CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.00174f
C606 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C607 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.28e-19
C608 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST 0.289f
C609 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST 0.335f
C610 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 VDD 0.386f
C611 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0477f
C612 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.111f
C613 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.CLK 0.00481f
C614 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5875_1502# 0.00118f
C615 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.431f
C616 a_7089_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.0202f
C617 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C618 a_4183_1458# CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.42e-20
C619 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.QB 0.28f
C620 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_1644_4227# 0.0733f
C621 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.Q0 0.0175f
C622 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 5.52e-20
C623 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C624 a_4704_4226# CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 8.64e-19
C625 CLK_div_31_mag_0.Q0 a_1798_3130# 6.43e-21
C626 a_18365_1305# CLK_div_3_mag_0.Q0 2.79e-20
C627 a_1859_352# RST 0.00186f
C628 a_8453_3965# CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.85e-20
C629 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C630 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.402f
C631 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_15912_1349# 0.00378f
C632 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_1.QB 1.34e-19
C633 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C634 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.QB 0.28f
C635 VDD CLK_div_31_mag_0.or_2_mag_0.IN1 0.729f
C636 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VDD 0.515f
C637 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_4.QB 0.103f
C638 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.Q3 0.00381f
C639 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C640 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK 2.15e-19
C641 a_4177_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C642 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 6.23e-20
C643 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT RST 0.012f
C644 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5311_1502# 0.011f
C645 CLK_div_31_mag_0.Q4 RST 1.1f
C646 a_7506_3203# VDD 3.14e-19
C647 CLK a_516_4227# 0.00207f
C648 CLK RST 0.662f
C649 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN RST 0.0239f
C650 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_1080_4227# 0.00378f
C651 a_19647_252# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C652 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C653 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 RST 0.0432f
C654 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.Q2 0.11f
C655 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_3_mag_0.CLK 2.47e-20
C656 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.655f
C657 a_7249_360# RST 0.00189f
C658 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_3.QB 0.199f
C659 VDD CLK_div_31_mag_0.JK_FF_mag_2.QB 0.911f
C660 VDD CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.752f
C661 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.00173f
C662 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_15348_1305# 0.0732f
C663 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C664 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C665 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C666 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q2 0.318f
C667 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 0.103f
C668 a_5465_405# CLK_div_31_mag_0.Q3 0.00859f
C669 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 1.59e-19
C670 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_4747_1502# 1.43e-19
C671 a_5582_3129# VDD 0.00503f
C672 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.394f
C673 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 6.28e-19
C674 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.431f
C675 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_0.QB 2e-21
C676 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_4140_4226# 0.0036f
C677 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN RST 5.63e-20
C678 a_19083_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C679 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 3.27e-20
C680 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 a_8453_3965# 0.00347f
C681 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C682 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD 0.745f
C683 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00542f
C684 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.77e-19
C685 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_31_mag_0.Q3 1.48e-20
C686 CLK_div_31_mag_0.JK_FF_mag_0.QB RST 0.169f
C687 VDD CLK_div_3_mag_0.or_2_mag_0.IN2 0.491f
C688 CLK_div_31_mag_0.Q3 VDD 3.04f
C689 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.121f
C690 VDD a_20057_1349# 3.56e-19
C691 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.516f
C692 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.107f
C693 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_17040_1349# 0.00372f
C694 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_15188_1305# 0.0203f
C695 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.365f
C696 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_4294_3129# 0.069f
C697 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1 1.12e-19
C698 a_1135_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C699 a_8452_3208# CLK_div_31_mag_0.Q2 0.00952f
C700 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN RST 0.0116f
C701 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.Q2 0.274f
C702 CLK_div_31_mag_0.JK_FF_mag_4.QB a_8947_1501# 0.0114f
C703 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_4183_1458# 0.00119f
C704 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_3_mag_0.CLK 3.46e-19
C705 a_18923_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C706 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VDD 0.517f
C707 a_981_1449# RST 9.22e-19
C708 a_7813_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 9.1e-19
C709 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 RST 0.00239f
C710 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN RST 0.00861f
C711 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_3.QB 0.25f
C712 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_31_mag_0.or_2_mag_0.IN1 1.18e-19
C713 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 4.02e-20
C714 VDD a_19493_1349# 3.14e-19
C715 CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.208f
C716 a_5428_4226# a_5588_4226# 0.0504f
C717 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.IN2 0.124f
C718 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 1.94f
C719 CLK_div_3_mag_0.CLK a_18641_2448# 0.0103f
C720 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.or_2_mag_0.IN2 0.00761f
C721 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 a_8383_1501# 3.59e-20
C722 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_16476_1349# 0.069f
C723 CLK_div_3_mag_0.JK_FF_mag_1.K a_20057_1349# 0.012f
C724 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT RST 0.00412f
C725 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 8.46e-19
C726 a_2987_396# RST 9.7e-19
C727 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_3730_3129# 0.00372f
C728 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00975f
C729 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0295f
C730 a_7089_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 1.17e-20
C731 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK 0.274f
C732 a_16066_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C733 CLK_div_31_mag_0.Q4 CLK 0.00641f
C734 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.CLK 0.272f
C735 CLK_div_31_mag_0.JK_FF_mag_4.QB a_8383_1501# 2.96e-19
C736 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.118f
C737 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.244f
C738 a_4858_3129# VDD 3.14e-19
C739 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST 0.27f
C740 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.41f
C741 a_18359_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C742 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C743 a_18923_208# a_19083_208# 0.0504f
C744 a_7249_360# CLK_div_31_mag_0.Q4 0.00789f
C745 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.Q2 0.00733f
C746 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.109f
C747 a_4901_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C748 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VDD 0.655f
C749 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0016f
C750 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.QB 1.14e-19
C751 a_6029_405# VDD 3.15e-19
C752 a_7249_360# CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 1.46e-19
C753 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 3.86e-20
C754 CLK_div_31_mag_0.Q1 VDD 3.87f
C755 a_1859_352# CLK_div_31_mag_0.JK_FF_mag_0.QB 0.00696f
C756 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.118f
C757 VDD a_18929_1349# 3.14e-19
C758 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 5.82e-21
C759 CLK_div_31_mag_0.or_2_mag_0.IN1 a_11989_2561# 0.0144f
C760 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.25f
C761 CLK_div_3_mag_0.JK_FF_mag_1.K a_19493_1349# 2.96e-19
C762 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.0012f
C763 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C764 a_7973_360# RST 0.00147f
C765 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C766 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.Q2 0.00281f
C767 CLK_div_31_mag_0.Q0 VDD 2.57f
C768 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.and_5_mag_0.VOUT 1.53e-22
C769 CLK_div_31_mag_0.JK_FF_mag_4.QB a_7819_1501# 3.33e-19
C770 CLK CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.3f
C771 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.11f
C772 a_4294_3129# VDD 3.14e-19
C773 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 RST 0.0212f
C774 a_18199_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C775 a_1705_1493# CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 5e-20
C776 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_670_3130# 2.21e-19
C777 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.269f
C778 CLK_div_3_mag_0.Q1 CLK_div_31_mag_0.or_2_mag_0.IN1 1.71e-20
C779 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_3_mag_0.Q1 5.66e-20
C780 a_2423_396# CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C781 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.08f
C782 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 a_9404_3954# 0.00347f
C783 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C784 a_7813_360# CLK_div_31_mag_0.JK_FF_mag_4.QB 0.00695f
C785 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 6.95e-19
C786 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 a_10367_3208# 0.00347f
C787 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_8383_1501# 4.52e-20
C788 CLK_div_3_mag_0.JK_FF_mag_1.K a_18929_1349# 1.75e-19
C789 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C790 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 7e-19
C791 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.QB 0.343f
C792 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.0405f
C793 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00127f
C794 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 3.59e-20
C795 CLK_div_31_mag_0.JK_FF_mag_4.QB a_7255_1457# 0.00392f
C796 a_3730_3129# VDD 3.56e-19
C797 a_1859_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C798 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.43f
C799 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.199f
C800 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_31_mag_0.Q4 0.00279f
C801 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 0.112f
C802 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_3.QB 3.09e-19
C803 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.01e-19
C804 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 RST 0.0196f
C805 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C806 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_31_mag_0.Q2 4.94e-20
C807 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C808 VDD a_18205_1305# 2.27e-19
C809 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 1.15e-19
C810 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.Q1 0.0636f
C811 CLK_div_31_mag_0.Q2 VDD 4.61f
C812 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN RST 0.00738f
C813 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_7819_1501# 0.0202f
C814 CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.or_2_mag_0.IN1 0.0103f
C815 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_31_mag_0.and_5_mag_0.VOUT 0.00527f
C816 CLK_div_3_mag_0.JK_FF_mag_1.K a_18365_1305# 0.00392f
C817 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.109f
C818 RST CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0865f
C819 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.or_2_mag_0.IN2 0.0138f
C820 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00166f
C821 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT RST 0.273f
C822 a_4177_361# RST 0.00189f
C823 a_7813_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.0203f
C824 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.119f
C825 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 1.97e-19
C826 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 3.81e-19
C827 CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.JK_FF_mag_2.QB 2.46e-21
C828 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.97e-19
C829 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 6.26e-20
C830 a_670_3130# RST 6.04e-19
C831 a_7973_360# CLK_div_31_mag_0.Q4 0.0101f
C832 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 7.4e-22
C833 a_9403_3219# RST 2.96e-19
C834 VDD a_17040_1349# 3.6e-19
C835 VDD CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.429f
C836 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.36f
C837 a_2987_396# CLK_div_31_mag_0.JK_FF_mag_0.QB 0.0811f
C838 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C839 CLK CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0108f
C840 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.CLK 7.81e-19
C841 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C842 a_20211_252# CLK_div_3_mag_0.Q0 0.0157f
C843 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.4e-21
C844 a_4023_1458# a_4183_1458# 0.0504f
C845 a_4704_4226# a_4864_4226# 0.0504f
C846 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.00517f
C847 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C848 a_18199_208# a_18359_208# 0.0504f
C849 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 a_9403_3219# 0.00347f
C850 CLK_div_31_mag_0.Q1 a_11989_2561# 1.78e-19
C851 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00103f
C852 CLK_div_3_mag_0.JK_FF_mag_1.QB RST 0.684f
C853 CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.106f
C854 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.98e-19
C855 a_4177_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C856 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 8.93e-21
C857 VDD a_16476_1349# 3.18e-19
C858 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C859 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.QB 0.00541f
C860 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.CLK 0.362f
C861 a_2833_1493# CLK_div_31_mag_0.Q2 0.069f
C862 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00107f
C863 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C864 a_5422_3129# CLK_div_31_mag_0.JK_FF_mag_3.QB 0.00392f
C865 a_8537_404# CLK_div_31_mag_0.JK_FF_mag_4.QB 0.00964f
C866 a_19647_252# CLK_div_3_mag_0.Q0 0.00859f
C867 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.Q0 0.0343f
C868 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.or_2_mag_0.IN2 1.82e-19
C869 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 1.03e-19
C870 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_7507_3970# 4.6e-21
C871 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.108f
C872 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.267f
C873 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 RST 1.08e-19
C874 VDD CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.655f
C875 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN RST 0.00657f
C876 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00392f
C877 CLK_div_31_mag_0.Q3 a_7507_3970# 0.00665f
C878 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0886f
C879 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00229f
C880 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00196f
C881 a_1798_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0202f
C882 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK 8.09e-19
C883 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 VDD 0.388f
C884 VDD a_15912_1349# 3.18e-19
C885 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_17040_1349# 0.00118f
C886 a_1135_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C887 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C888 CLK CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.013f
C889 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q3 3.08e-19
C890 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.657f
C891 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C892 a_4858_3129# CLK_div_31_mag_0.JK_FF_mag_3.QB 3.29e-19
C893 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C894 a_975_352# VDD 0.00108f
C895 a_19083_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C896 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.Q1 0.104f
C897 CLK CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0219f
C898 a_19083_208# CLK_div_3_mag_0.Q0 0.0101f
C899 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 4.17e-19
C900 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C901 a_7095_1457# a_7255_1457# 0.0504f
C902 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 RST 0.0132f
C903 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_19493_1349# 0.0059f
C904 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 2.63e-20
C905 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.12f
C906 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 8.53e-19
C907 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.515f
C908 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 3.34e-21
C909 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.2f
C910 a_4901_361# CLK_div_31_mag_0.JK_FF_mag_1.QB 0.00696f
C911 CLK_div_31_mag_0.or_2_mag_0.IN1 RST 0.226f
C912 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN RST 0.0233f
C913 a_19614_2684# CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C914 VDD a_2528_4227# 0.00108f
C915 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_8947_1501# 3.59e-20
C916 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_3.QB 0.00585f
C917 a_7506_3203# RST 3.99e-19
C918 CLK a_670_3130# 3.7e-19
C919 CLK_div_3_mag_0.CLK CLK_div_31_mag_0.or_2_mag_0.IN1 0.00923f
C920 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_3_mag_0.CLK 0.00153f
C921 a_4901_361# RST 0.00187f
C922 a_1234_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 4.52e-20
C923 a_8537_404# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.00378f
C924 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_2368_4227# 8.66e-20
C925 VDD a_15348_1305# 2.65e-19
C926 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C927 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 RST 0.163f
C928 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.QB 1.97f
C929 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_16476_1349# 0.011f
C930 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.04e-20
C931 a_4294_3129# CLK_div_31_mag_0.JK_FF_mag_3.QB 2.96e-19
C932 CLK_div_31_mag_0.JK_FF_mag_2.QB a_516_4227# 0.0811f
C933 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT RST 0.051f
C934 a_18923_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C935 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C936 RST CLK_div_31_mag_0.JK_FF_mag_2.QB 0.117f
C937 a_9101_404# CLK_div_31_mag_0.Q4 0.0157f
C938 a_18923_208# CLK_div_3_mag_0.Q0 0.0102f
C939 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_18929_1349# 0.0697f
C940 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 a_8452_3208# 0.00347f
C941 a_18205_1305# CLK_div_3_mag_0.Q1 0.00149f
C942 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C943 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 2.74e-20
C944 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C945 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C946 a_5582_3129# RST 8.67e-19
C947 CLK_div_31_mag_0.Q1 a_7507_3970# 0.00353f
C948 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 RST 0.0606f
C949 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.Q3 1.97f
C950 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.431f
C951 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT RST 0.0173f
C952 VDD a_15188_1305# 6.05e-19
C953 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.CLK 5.57e-19
C954 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_15912_1349# 1.43e-19
C955 CLK_div_31_mag_0.Q0 a_7507_3970# 0.00389f
C956 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 0.0103f
C957 a_4901_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C958 a_3730_3129# CLK_div_31_mag_0.JK_FF_mag_3.QB 0.0114f
C959 CLK_div_31_mag_0.Q3 RST 0.328f
C960 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C961 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C962 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN RST 0.00749f
C963 a_18359_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C964 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00133f
C965 a_18359_208# CLK_div_3_mag_0.Q0 0.00789f
C966 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.392f
C967 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 5.96e-22
C968 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VDD 0.385f
C969 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.or_2_mag_0.IN2 6.62e-20
C970 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_2269_1493# 0.069f
C971 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.VOUT 5.82e-21
C972 CLK CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.101f
C973 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.3f
C974 a_17040_1349# CLK_div_3_mag_0.Q1 0.069f
C975 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN CLK_div_3_mag_0.CLK 0.00347f
C976 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK 0.00127f
C977 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VDD 0.519f
C978 VDD a_1804_4227# 2.21e-19
C979 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 2.36e-20
C980 a_5422_3129# RST 7.2e-19
C981 CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.Q2 0.0154f
C982 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_4747_1502# 0.00378f
C983 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.and_5_mag_0.VOUT 3.56e-19
C984 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_5588_4226# 0.0202f
C985 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.Q3 0.0781f
C986 a_5465_405# CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C987 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN RST 0.0163f
C988 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00166f
C989 CLK_div_31_mag_0.Q1 a_1135_352# 0.00164f
C990 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_15348_1305# 0.00119f
C991 CLK_div_3_mag_0.JK_FF_mag_1.K a_15188_1305# 8.64e-19
C992 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C993 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK 1.44e-19
C994 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C995 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.or_2_mag_0.IN1 0.091f
C996 a_18199_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C997 a_18199_208# CLK_div_3_mag_0.Q0 0.00335f
C998 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD 0.75f
C999 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C1000 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.112f
C1001 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.108f
C1002 a_1859_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C1003 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.118f
C1004 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VDD 0.512f
C1005 CLK_div_31_mag_0.Q4 a_7506_3203# 0.00353f
C1006 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.24f
C1007 a_1699_352# VDD 2.21e-19
C1008 a_20211_252# VDD 3.14e-19
C1009 a_7506_3203# CLK 2.26e-19
C1010 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.16f
C1011 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.Q3 0.0345f
C1012 a_10367_3208# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.069f
C1013 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_1234_3130# 0.069f
C1014 a_4858_3129# RST 3.98e-19
C1015 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_5311_1502# 0.0059f
C1016 CLK_div_31_mag_0.Q2 a_7507_3970# 0.0108f
C1017 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_4183_1458# 0.0732f
C1018 CLK CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00955f
C1019 a_6029_405# CLK_div_31_mag_0.JK_FF_mag_1.QB 0.0811f
C1020 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_1080_4227# 0.0036f
C1021 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 VDD 0.389f
C1022 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.Q2 0.0262f
C1023 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 RST 0.162f
C1024 a_6029_405# RST 9.82e-19
C1025 CLK CLK_div_31_mag_0.JK_FF_mag_2.QB 0.106f
C1026 CLK_div_31_mag_0.Q1 a_516_4227# 0.0157f
C1027 CLK_div_31_mag_0.Q1 RST 0.23f
C1028 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_5428_4226# 0.0731f
C1029 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C1030 a_18929_1349# RST 1.9e-19
C1031 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.122f
C1032 CLK_div_3_mag_0.Q0 a_19614_2684# 0.0134f
C1033 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.998f
C1034 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.517f
C1035 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_5582_3129# 0.0203f
C1036 a_5875_1502# VDD 3.56e-19
C1037 a_4294_3129# CLK_div_31_mag_0.JK_FF_mag_1.QB 4.61e-20
C1038 a_19647_252# VDD 3.14e-19
C1039 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.995f
C1040 a_18929_1349# CLK_div_3_mag_0.CLK 6.43e-21
C1041 a_5582_3129# CLK 0.0118f
C1042 CLK_div_31_mag_0.Q0 RST 0.274f
C1043 a_7089_360# VDD 0.00108f
C1044 a_20211_252# CLK_div_3_mag_0.JK_FF_mag_1.K 0.0811f
C1045 VDD a_1080_4227# 3.14e-19
C1046 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 1.73e-20
C1047 CLK CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0477f
C1048 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.Q1 0.00335f
C1049 a_4294_3129# RST 0.00173f
C1050 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_4747_1502# 0.0697f
C1051 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.00669f
C1052 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_4023_1458# 0.0203f
C1053 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Q3 0.29f
C1054 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0512f
C1055 a_7507_3970# CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C1056 a_5588_4226# VDD 0.00108f
C1057 CLK CLK_div_31_mag_0.Q3 0.198f
C1058 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 2.66e-19
C1059 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.0886f
C1060 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 4.31e-19
C1061 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VDD 0.39f
C1062 a_4858_3129# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.61e-20
C1063 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 RST 0.00941f
C1064 a_1135_352# CLK_div_31_mag_0.Q2 0.00789f
C1065 CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 1.14e-19
C1066 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.0181f
C1067 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.Q3 0.438f
C1068 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.00527f
C1069 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK 0.471f
C1070 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_4864_4226# 9.1e-19
C1071 a_18365_1305# RST 6.43e-19
C1072 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 a_8947_1501# 0.00372f
C1073 a_2362_3130# a_2522_3130# 0.0504f
C1074 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.0592f
C1075 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_0.QB 0.103f
C1076 CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0386f
C1077 VDD a_8947_1501# 3.56e-19
C1078 a_7249_360# CLK_div_31_mag_0.Q3 0.00214f
C1079 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_5422_3129# 0.0732f
C1080 a_5311_1502# VDD 3.14e-19
C1081 CLK_div_31_mag_0.JK_FF_mag_4.QB VDD 0.912f
C1082 a_15348_1305# CLK_div_3_mag_0.Q1 2.79e-20
C1083 a_18365_1305# CLK_div_3_mag_0.CLK 0.00939f
C1084 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 a_8947_1501# 4.52e-20
C1085 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_4.QB 0.199f
C1086 a_5422_3129# CLK 0.0106f
C1087 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C1088 a_19647_252# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00964f
C1089 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C1090 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_31_mag_0.Q4 0.00141f
C1091 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.00162f
C1092 a_3730_3129# RST 0.00252f
C1093 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN RST 3.56e-20
C1094 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.Q2 0.321f
C1095 a_8537_404# CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.76e-20
C1096 a_18205_1305# RST 7.78e-19
C1097 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.QB 0.28f
C1098 CLK_div_31_mag_0.Q2 RST 1.03f
C1099 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_4704_4226# 2.88e-20
C1100 VDD CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C1101 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 a_8383_1501# 0.069f
C1102 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.JK_FF_mag_0.QB 2.1e-19
C1103 a_9403_3219# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C1104 VDD a_8383_1501# 3.14e-19
C1105 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_4858_3129# 0.00378f
C1106 a_4747_1502# VDD 3.14e-19
C1107 a_18205_1305# CLK_div_3_mag_0.CLK 0.0101f
C1108 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.36f
C1109 a_18923_208# VDD 2.21e-19
C1110 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C1111 a_4858_3129# CLK 3.01e-19
C1112 a_19083_208# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00696f
C1113 a_15906_208# a_16066_208# 0.0504f
C1114 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.00662f
C1115 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 3.48e-19
C1116 a_2423_396# VDD 3.14e-19
C1117 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.112f
C1118 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.33e-20
C1119 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.Q2 0.0127f
C1120 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 0.338f
C1121 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q4 0.79f
C1122 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.233f
C1123 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.00975f
C1124 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C1125 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 3.48e-19
C1126 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VDD 0.998f
C1127 CLK_div_31_mag_0.Q1 CLK 1.26f
C1128 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.122f
C1129 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 6.25e-19
C1130 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD 0.401f
C1131 a_17040_1349# RST 7.24e-19
C1132 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 9.41e-19
C1133 CLK_div_3_mag_0.or_2_mag_0.IN2 a_18641_2448# 7.48e-20
C1134 VDD a_7819_1501# 3.14e-19
C1135 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_20057_1349# 4.52e-20
C1136 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.Q4 0.197f
C1137 a_4864_4226# VDD 2.21e-19
C1138 CLK_div_31_mag_0.Q0 CLK 0.636f
C1139 a_17040_1349# CLK_div_3_mag_0.CLK 9.45e-19
C1140 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 7.44e-19
C1141 a_18359_208# VDD 0.00305f
C1142 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.00376f
C1143 a_18923_208# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00695f
C1144 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.Q2 0.00182f
C1145 a_2269_1493# VDD 3.14e-19
C1146 a_7813_360# VDD 2.21e-19
C1147 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1.9e-21
C1148 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 8.4e-19
C1149 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.112f
C1150 a_10368_3965# VDD 5.2e-19
C1151 a_16476_1349# RST 8.63e-19
C1152 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 8.03e-20
C1153 a_975_352# a_1135_352# 0.0504f
C1154 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_0.QB 0.308f
C1155 a_2833_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C1156 a_4023_1458# VDD 0.00519f
C1157 a_1859_352# CLK_div_31_mag_0.Q2 0.0101f
C1158 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C1159 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.664f
C1160 VDD CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.426f
C1161 a_18199_208# VDD 0.00743f
C1162 a_16476_1349# CLK_div_3_mag_0.CLK 6.06e-21
C1163 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C1164 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 5.09e-24
C1165 a_1705_1493# VDD 3.14e-19
C1166 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 9.89e-20
C1167 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_0.QB 0.00258f
C1168 CLK CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.046f
C1169 RST CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.204f
C1170 a_1141_1449# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 3.87e-20
C1171 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.Q1 4.33e-19
C1172 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.Q2 0.00739f
C1173 a_8452_3208# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C1174 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Q2 0.197f
C1175 CLK CLK_div_31_mag_0.Q2 0.327f
C1176 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 RST 2.65e-20
C1177 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_3.QB 6.46e-19
C1178 CLK_div_31_mag_0.Q1 a_981_1449# 0.0101f
C1179 a_15912_1349# RST 2.23e-19
C1180 a_9404_3954# VDD 3.14e-19
C1181 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.Q2 7.84e-19
C1182 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 1.56e-21
C1183 a_1705_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C1184 VDD a_7095_1457# 0.00554f
C1185 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 RST 0.21f
C1186 a_15912_1349# CLK_div_3_mag_0.CLK 6.43e-21
C1187 a_4140_4226# VDD 3.14e-19
C1188 a_17194_252# VDD 0.00149f
C1189 VDD a_19614_2684# 0.172f
C1190 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 6.46e-19
C1191 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C1192 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00161f
C1193 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C1194 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.CLK 0.013f
C1195 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN RST 0.0149f
C1196 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_18929_1349# 0.00378f
C1197 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C1198 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_16476_1349# 4.52e-20
C1199 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 2.8e-19
C1200 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 RST 0.0968f
C1201 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_2.QB 0.103f
C1202 RST a_2528_4227# 9.7e-19
C1203 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.4e-19
C1204 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD 0.431f
C1205 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 9.67e-20
C1206 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00164f
C1207 CLK CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0454f
C1208 a_4017_361# VDD 0.00108f
C1209 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C1210 a_8453_3965# VDD 3.14e-19
C1211 a_15348_1305# RST 6.43e-19
C1212 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 3.09e-19
C1213 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C1214 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.QB 2f
C1215 a_1141_1449# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C1216 a_2269_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C1217 a_670_3130# CLK_div_31_mag_0.JK_FF_mag_2.QB 0.0114f
C1218 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C1219 a_15348_1305# CLK_div_3_mag_0.CLK 0.00939f
C1220 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q3 0.314f
C1221 a_3576_4226# VDD 3.15e-19
C1222 a_7973_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 8.64e-19
C1223 a_16630_252# VDD 0.00149f
C1224 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C1225 CLK_div_3_mag_0.JK_FF_mag_1.K a_19614_2684# 0.00168f
C1226 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 4.48e-19
C1227 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_19614_2684# 3.25e-19
C1228 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_18365_1305# 0.0732f
C1229 a_15182_208# a_15342_208# 0.0504f
C1230 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_15912_1349# 0.0202f
C1231 a_2522_3130# VDD 0.00523f
C1232 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C1233 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C1234 RST a_2368_4227# 9.7e-19
C1235 a_4177_361# CLK_div_31_mag_0.Q3 0.00789f
C1236 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00288f
C1237 a_10367_3208# VDD 5.19e-19
C1238 a_18923_208# CLK_div_3_mag_0.Q1 3.6e-22
C1239 a_2362_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00119f
C1240 a_5311_1502# CLK_div_31_mag_0.JK_FF_mag_3.QB 4.61e-20
C1241 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.61e-20
C1242 a_8537_404# VDD 3.14e-19
C1243 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C1244 a_15188_1305# RST 7.78e-19
C1245 a_1705_1493# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C1246 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C1247 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 5.53e-19
C1248 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00279f
C1249 a_8537_404# CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.069f
C1250 a_9403_3219# CLK_div_31_mag_0.Q3 0.0193f
C1251 a_15188_1305# CLK_div_3_mag_0.CLK 0.0101f
C1252 a_16066_208# VDD 9.82e-19
C1253 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VDD 0.519f
C1254 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.or_2_mag_0.IN2 3.81e-19
C1255 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_516_4227# 0.00372f
C1256 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C1257 RST CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 8.38e-19
C1258 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_20057_1349# 0.00372f
C1259 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 RST 0.00927f
C1260 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_18205_1305# 0.0203f
C1261 a_7506_3203# CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C1262 CLK CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00418f
C1263 a_2987_396# CLK_div_31_mag_0.Q2 0.0157f
C1264 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN RST 0.0417f
C1265 a_19083_208# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C1266 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.175f
C1267 RST a_1804_4227# 0.00155f
C1268 a_18359_208# CLK_div_3_mag_0.Q1 1.86e-20
C1269 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C1270 CLK CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0502f
C1271 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C1272 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.401f
C1273 a_1798_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.43e-19
C1274 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD 0.739f
C1275 VDD CLK_div_3_mag_0.Q0 1.29f
C1276 a_6029_405# CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00372f
C1277 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.207f
C1278 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 4.92e-21
C1279 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VDD 0.769f
C1280 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.0169f
C1281 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C1282 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.403f
C1283 a_4858_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0202f
C1284 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 7.75e-19
C1285 a_3730_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C1286 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.089f
C1287 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.046f
C1288 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT RST 0.0826f
C1289 a_15906_208# VDD 0.0012f
C1290 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 3e-20
C1291 CLK CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.417f
C1292 a_16630_252# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C1293 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 5.47e-20
C1294 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 1.97e-19
C1295 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_19493_1349# 0.069f
C1296 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 3.68e-19
C1297 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 RST 0.126f
C1298 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.432f
C1299 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN RST 0.0411f
C1300 CLK a_2528_4227# 0.00165f
C1301 a_1699_352# RST 8.64e-19
C1302 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.349f
C1303 a_1798_3130# VDD 3.14e-19
C1304 RST a_1644_4227# 0.00127f
C1305 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 7.24e-19
C1306 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00139f
C1307 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0048f
C1308 a_18199_208# CLK_div_3_mag_0.Q1 2.55e-20
C1309 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 6.2e-20
C1310 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_31_mag_0.Q2 2.84e-19
C1311 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 1.05e-20
C1312 a_1234_3130# CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C1313 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q3 0.0129f
C1314 CLK_div_31_mag_0.JK_FF_mag_3.QB a_4864_4226# 0.00695f
C1315 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.235f
C1316 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.0881f
C1317 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 RST 4.4e-20
C1318 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C1319 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q0 8.04e-19
C1320 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0 2.37f
C1321 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0343f
C1322 a_4017_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C1323 VDD CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.517f
C1324 CLK_div_31_mag_0.Q1 a_670_3130# 0.069f
C1325 CLK_div_31_mag_0.JK_FF_mag_1.QB a_5875_1502# 0.0114f
C1326 a_4294_3129# CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.52e-20
C1327 a_4741_361# VDD 2.21e-19
C1328 a_15342_208# VDD 0.00888f
C1329 CLK_div_31_mag_0.Q1 a_9403_3219# 7.37e-19
C1330 RST CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.263f
C1331 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_31_mag_0.JK_FF_mag_2.QB 0.0381f
C1332 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C1333 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN RST 0.022f
C1334 a_5875_1502# RST 0.00126f
C1335 a_8452_3208# VDD 3.14e-19
C1336 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST 0.276f
C1337 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.745f
C1338 CLK a_2368_4227# 0.00165f
C1339 a_2423_396# CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C1340 a_1234_3130# VDD 3.14e-19
C1341 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_31_mag_0.Q3 0.109f
C1342 a_7089_360# RST 0.00189f
C1343 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.00165f
C1344 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.CLK 0.00302f
C1345 a_17194_252# CLK_div_3_mag_0.Q1 0.0157f
C1346 CLK_div_3_mag_0.Q1 a_19614_2684# 6.83e-19
C1347 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C1348 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.012f
C1349 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 7e-19
C1350 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00116f
C1351 CLK_div_31_mag_0.JK_FF_mag_3.QB a_4704_4226# 0.00696f
C1352 a_7506_3203# CLK_div_31_mag_0.Q3 0.0108f
C1353 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_2833_1493# 0.00372f
C1354 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00279f
C1355 a_4901_361# CLK_div_31_mag_0.Q3 0.0101f
C1356 a_16066_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C1357 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.93e-19
C1358 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 RST 0.00589f
C1359 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.and_5_mag_0.VOUT 2.17e-20
C1360 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 2.44e-21
C1361 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.00203f
C1362 CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_31_mag_0.JK_FF_mag_4.QB 2.42e-21
C1363 CLK_div_31_mag_0.JK_FF_mag_1.QB a_5311_1502# 2.96e-19
C1364 CLK CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0132f
C1365 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.4e-19
C1366 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C1367 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK 0.0014f
C1368 a_15182_208# VDD 0.0132f
C1369 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C1370 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q2 8.87e-19
C1371 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_31_mag_0.Q4 0.00138f
C1372 CLK_div_31_mag_0.JK_FF_mag_4.QB RST 0.11f
C1373 a_8947_1501# RST 6.56e-19
C1374 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2269_1493# 0.011f
C1375 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_31_mag_0.or_2_mag_0.IN1 0.0042f
C1376 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 0.112f
C1377 a_5311_1502# RST 0.00126f
C1378 CLK a_1804_4227# 0.00133f
C1379 a_19083_208# RST 0.00103f
C1380 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C1381 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.00102f
C1382 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_2522_3130# 0.0203f
C1383 a_1699_352# a_1859_352# 0.0504f
C1384 a_16630_252# CLK_div_3_mag_0.Q1 0.00859f
C1385 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 4.3e-20
C1386 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 5.06e-21
C1387 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_31_mag_0.Q2 0.00147f
C1388 a_4177_361# CLK_div_31_mag_0.Q2 0.00216f
C1389 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.402f
C1390 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0014f
C1391 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD 0.756f
C1392 CLK_div_31_mag_0.JK_FF_mag_3.QB a_4140_4226# 0.00964f
C1393 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C1394 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0443f
C1395 a_975_352# CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C1396 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.Q4 0.338f
C1397 CLK_div_31_mag_0.Q3 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.318f
C1398 a_15906_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C1399 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_31_mag_0.JK_FF_mag_4.QB 3.95e-19
C1400 CLK_div_3_mag_0.JK_FF_mag_1.QB a_18365_1305# 1.41e-20
C1401 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01e-19
C1402 CLK_div_31_mag_0.JK_FF_mag_1.QB a_4747_1502# 3.25e-19
C1403 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 0.00956f
C1404 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_31_mag_0.Q3 0.269f
C1405 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.00118f
C1406 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK 6.68e-19
C1407 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 RST 0.0205f
C1408 a_9403_3219# CLK_div_31_mag_0.Q2 9.22e-21
C1409 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0943f
C1410 a_15342_208# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C1411 a_8383_1501# RST 6.56e-19
C1412 a_4747_1502# RST 6.86e-19
C1413 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_1705_1493# 1.43e-19
C1414 a_5422_3129# a_5582_3129# 0.0504f
C1415 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.655f
C1416 CLK a_1644_4227# 0.00133f
C1417 a_7249_360# CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.0731f
C1418 a_18923_208# RST 0.00119f
C1419 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_2362_3130# 0.0732f
C1420 a_16066_208# CLK_div_3_mag_0.Q1 0.0101f
C1421 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.or_2_mag_0.IN1 1.64e-19
C1422 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_5311_1502# 4.52e-20
C1423 CLK CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0512f
C1424 a_2423_396# RST 9.46e-19
C1425 CLK_div_31_mag_0.JK_FF_mag_3.QB a_3576_4226# 0.0811f
C1426 a_15342_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C1427 CLK_div_31_mag_0.Q1 a_7506_3203# 2.95e-21
C1428 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT RST 0.259f
C1429 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.00907f
C1430 CLK_div_3_mag_0.JK_FF_mag_1.QB a_18205_1305# 1.86e-20
C1431 CLK CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.019f
C1432 CLK_div_31_mag_0.JK_FF_mag_1.QB a_4183_1458# 0.00392f
C1433 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 RST 0.00822f
C1434 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 0.00529f
C1435 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00396f
C1436 a_7089_360# CLK_div_31_mag_0.Q4 0.00335f
C1437 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.321f
C1438 CLK_div_31_mag_0.Q0 a_7506_3203# 0.00347f
C1439 CLK_div_31_mag_0.JK_FF_mag_3.QB a_2522_3130# 1.76e-20
C1440 a_7819_1501# RST 5.43e-19
C1441 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 9.98e-19
C1442 VDD CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.32f
C1443 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q0 0.0285f
C1444 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_1141_1449# 0.00119f
C1445 a_4741_361# CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C1446 a_19493_1349# CLK_div_3_mag_0.or_2_mag_0.IN2 4.9e-20
C1447 a_4183_1458# RST 0.00229f
C1448 a_4864_4226# RST 8.64e-19
C1449 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.127f
C1450 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C1451 CLK a_1080_4227# 0.00194f
C1452 a_5465_405# VDD 3.14e-19
C1453 a_18359_208# RST 0.00218f
C1454 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_31_mag_0.JK_FF_mag_0.QB 7.57e-20
C1455 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_2.QB 1.99f
C1456 a_1699_352# CLK_div_31_mag_0.JK_FF_mag_0.QB 0.00695f
C1457 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C1458 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 9.71e-20
C1459 a_2269_1493# RST 0.00165f
C1460 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1 0.109f
C1461 a_18359_208# CLK_div_3_mag_0.CLK 0.00164f
C1462 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_1798_3130# 0.00378f
C1463 a_15906_208# CLK_div_3_mag_0.Q1 0.0102f
C1464 a_7089_360# a_7249_360# 0.0504f
C1465 CLK a_5588_4226# 0.00544f
C1466 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4747_1502# 0.0202f
C1467 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0107f
C1468 CLK_div_31_mag_0.Q2 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0127f
C1469 a_7813_360# RST 0.0017f
C1470 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_2.QB 0.307f
C1471 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 0.128f
C1472 a_15182_208# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C1473 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_31_mag_0.Q2 0.0728f
C1474 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 1.29e-20
C1475 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.88e-19
C1476 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.122f
C1477 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VDD 0.4f
C1478 CLK_div_31_mag_0.Q4 a_8947_1501# 0.0695f
C1479 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00122f
C1480 CLK_div_3_mag_0.JK_FF_mag_1.QB a_17040_1349# 0.0112f
C1481 CLK_div_31_mag_0.JK_FF_mag_1.QB a_7255_1457# 1.33e-20
C1482 CLK_div_31_mag_0.Q4 CLK_div_31_mag_0.JK_FF_mag_4.QB 1.98f
C1483 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_31_mag_0.Q3 3.38e-19
C1484 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 8.16e-20
C1485 a_10368_3965# RST 6.53e-20
C1486 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VDD 0.391f
C1487 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 8.48e-20
C1488 CLK_div_31_mag_0.JK_FF_mag_3.QB a_2362_3130# 1.35e-20
C1489 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_8947_1501# 0.00118f
C1490 CLK_div_31_mag_0.Q0 a_5582_3129# 5.54e-19
C1491 a_6029_405# CLK_div_31_mag_0.Q3 0.0157f
C1492 CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.28f
C1493 a_7255_1457# RST 0.00154f
C1494 CLK_div_31_mag_0.Q1 CLK_div_31_mag_0.Q3 0.812f
C1495 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 6.3e-20
C1496 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C1497 a_4023_1458# RST 0.003f
C1498 a_4704_4226# RST 0.00173f
C1499 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT RST 0.0042f
C1500 a_18199_208# RST 0.00218f
C1501 a_20211_252# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C1502 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_31_mag_0.Q2 0.0064f
C1503 CLK_div_31_mag_0.Q0 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 2.86e-19
C1504 a_1705_1493# RST 3.21e-19
C1505 a_20211_252# VSS 0.0675f
C1506 a_19647_252# VSS 0.0676f
C1507 a_19083_208# VSS 0.0343f
C1508 a_18923_208# VSS 0.0881f
C1509 a_18359_208# VSS 0.0343f
C1510 a_18199_208# VSS 0.0881f
C1511 a_17194_252# VSS 0.0675f
C1512 a_16630_252# VSS 0.0676f
C1513 a_16066_208# VSS 0.0343f
C1514 a_15906_208# VSS 0.0881f
C1515 a_15342_208# VSS 0.0343f
C1516 a_15182_208# VSS 0.0881f
C1517 a_9101_404# VSS 0.0675f
C1518 a_8537_404# VSS 0.0676f
C1519 a_7973_360# VSS 0.0343f
C1520 a_7813_360# VSS 0.0881f
C1521 a_7249_360# VSS 0.0343f
C1522 a_7089_360# VSS 0.0881f
C1523 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C1524 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.541f
C1525 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C1526 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C1527 a_6029_405# VSS 0.0675f
C1528 a_5465_405# VSS 0.0676f
C1529 a_4901_361# VSS 0.0343f
C1530 a_4741_361# VSS 0.0881f
C1531 a_4177_361# VSS 0.0343f
C1532 a_4017_361# VSS 0.0881f
C1533 a_2987_396# VSS 0.0686f
C1534 a_2423_396# VSS 0.0687f
C1535 a_1859_352# VSS 0.036f
C1536 a_1699_352# VSS 0.0898f
C1537 a_1135_352# VSS 0.036f
C1538 a_975_352# VSS 0.0899f
C1539 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VSS 0.677f
C1540 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VSS 0.662f
C1541 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VSS 0.662f
C1542 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VSS 0.662f
C1543 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VSS 0.666f
C1544 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VSS 0.677f
C1545 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VSS 0.762f
C1546 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VSS 0.417f
C1547 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VSS 0.541f
C1548 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C1549 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.541f
C1550 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.419f
C1551 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.546f
C1552 a_20057_1349# VSS 0.0676f
C1553 a_19493_1349# VSS 0.0676f
C1554 a_18929_1349# VSS 0.0676f
C1555 a_18365_1305# VSS 0.0343f
C1556 a_18205_1305# VSS 0.0881f
C1557 a_17040_1349# VSS 0.0676f
C1558 a_16476_1349# VSS 0.0676f
C1559 a_15912_1349# VSS 0.0676f
C1560 a_15348_1305# VSS 0.0343f
C1561 a_15188_1305# VSS 0.0881f
C1562 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VSS 0.707f
C1563 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VSS 0.698f
C1564 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VSS 0.698f
C1565 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VSS 0.708f
C1566 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VSS 0.681f
C1567 a_8947_1501# VSS 0.0676f
C1568 a_8383_1501# VSS 0.0676f
C1569 a_7819_1501# VSS 0.0676f
C1570 a_7255_1457# VSS 0.0343f
C1571 a_7095_1457# VSS 0.0881f
C1572 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VSS 0.761f
C1573 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS 1.68f
C1574 CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VSS 0.703f
C1575 a_5875_1502# VSS 0.0676f
C1576 a_5311_1502# VSS 0.0676f
C1577 a_4747_1502# VSS 0.0676f
C1578 a_4183_1458# VSS 0.0343f
C1579 a_4023_1458# VSS 0.0881f
C1580 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1581 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.692f
C1582 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C1583 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C1584 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1585 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1586 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.695f
C1587 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C1588 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C1589 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C1590 CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.859f
C1591 CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.56f
C1592 a_2833_1493# VSS 0.0676f
C1593 a_2269_1493# VSS 0.0676f
C1594 a_1705_1493# VSS 0.0676f
C1595 a_1141_1449# VSS 0.0343f
C1596 a_981_1449# VSS 0.0881f
C1597 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VSS 0.413f
C1598 CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 VSS 0.706f
C1599 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VSS 0.724f
C1600 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VSS 0.809f
C1601 CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VSS 0.507f
C1602 CLK_div_31_mag_0.JK_FF_mag_4.QB VSS 0.929f
C1603 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C1604 CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.691f
C1605 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.724f
C1606 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.809f
C1607 CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.507f
C1608 CLK_div_31_mag_0.JK_FF_mag_1.QB VSS 0.886f
C1609 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.413f
C1610 CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.739f
C1611 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C1612 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.814f
C1613 CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.507f
C1614 CLK_div_31_mag_0.JK_FF_mag_0.QB VSS 1.61f
C1615 a_18641_2448# VSS 0.0676f
C1616 Vdiv93 VSS 0.425f
C1617 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C1618 a_19614_2684# VSS 0.0247f
C1619 CLK_div_3_mag_0.Q0 VSS 1.99f
C1620 CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.418f
C1621 CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.602f
C1622 a_11989_2561# VSS 0.0247f
C1623 CLK_div_31_mag_0.or_2_mag_0.IN1 VSS 1.34f
C1624 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C1625 CLK_div_3_mag_0.Q1 VSS 1.77f
C1626 CLK_div_3_mag_0.CLK VSS 3.53f
C1627 CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN VSS 0.413f
C1628 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.446f
C1629 a_10367_3208# VSS 0.073f
C1630 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS 0.4f
C1631 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.451f
C1632 a_9403_3219# VSS 0.0757f
C1633 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS 0.397f
C1634 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.443f
C1635 a_8452_3208# VSS 0.073f
C1636 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS 0.393f
C1637 CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.445f
C1638 a_7506_3203# VSS 0.072f
C1639 a_5582_3129# VSS 0.0881f
C1640 a_5422_3129# VSS 0.0343f
C1641 a_4858_3129# VSS 0.0676f
C1642 a_4294_3129# VSS 0.0676f
C1643 a_3730_3129# VSS 0.0676f
C1644 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.507f
C1645 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.412f
C1646 CLK_div_31_mag_0.Q4 VSS 3.96f
C1647 a_2522_3130# VSS 0.0881f
C1648 a_2362_3130# VSS 0.0343f
C1649 a_1798_3130# VSS 0.0676f
C1650 a_1234_3130# VSS 0.0676f
C1651 a_670_3130# VSS 0.0676f
C1652 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C1653 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.413f
C1654 a_10368_3965# VSS 0.073f
C1655 a_9404_3954# VSS 0.0757f
C1656 a_8453_3965# VSS 0.073f
C1657 CLK_div_31_mag_0.and_5_mag_0.VOUT VSS 2.97f
C1658 a_7507_3970# VSS 0.0717f
C1659 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.465f
C1660 CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS 0.4f
C1661 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.451f
C1662 CLK_div_31_mag_0.Q2 VSS 4.42f
C1663 CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS 0.398f
C1664 a_5588_4226# VSS 0.0881f
C1665 a_5428_4226# VSS 0.0343f
C1666 a_4864_4226# VSS 0.0881f
C1667 a_4704_4226# VSS 0.0343f
C1668 a_4140_4226# VSS 0.0676f
C1669 a_3576_4226# VSS 0.0675f
C1670 CLK_div_31_mag_0.JK_FF_mag_3.QB VSS 0.885f
C1671 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.807f
C1672 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.699f
C1673 CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.416f
C1674 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.445f
C1675 CLK_div_31_mag_0.Q3 VSS 6.07f
C1676 CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS 0.395f
C1677 CLK VSS 4.43f
C1678 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.537f
C1679 CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.723f
C1680 a_2528_4227# VSS 0.0881f
C1681 a_2368_4227# VSS 0.0343f
C1682 a_1804_4227# VSS 0.0881f
C1683 a_1644_4227# VSS 0.0343f
C1684 a_1080_4227# VSS 0.0676f
C1685 a_516_4227# VSS 0.0675f
C1686 CLK_div_31_mag_0.JK_FF_mag_2.QB VSS 0.923f
C1687 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.807f
C1688 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.716f
C1689 CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.416f
C1690 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.54f
C1691 RST VSS 9.08f
C1692 CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.723f
C1693 CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.448f
C1694 CLK_div_31_mag_0.Q1 VSS 7.39f
C1695 CLK_div_31_mag_0.Q0 VSS 3.73f
C1696 VDD VSS 0.148p
C1697 CLK.t1 VSS 0.00895f
C1698 CLK.t4 VSS 0.0112f
C1699 CLK.n0 VSS 0.0265f
C1700 CLK.n1 VSS 0.193f
C1701 CLK.n2 VSS 0.359f
C1702 CLK.n3 VSS 0.136f
C1703 CLK.n4 VSS 0.00274f
C1704 CLK.n5 VSS 0.00708f
C1705 CLK.n6 VSS 0.00868f
C1706 CLK.n7 VSS 0.00722f
C1707 CLK.t3 VSS 0.0156f
C1708 CLK.t5 VSS 0.0103f
C1709 CLK.n8 VSS 0.0276f
C1710 CLK.n9 VSS 0.0036f
C1711 CLK.n10 VSS 0.00259f
C1712 CLK.n11 VSS 0.00128f
C1713 CLK.t7 VSS 0.0156f
C1714 CLK.t6 VSS 0.0103f
C1715 CLK.n12 VSS 0.0276f
C1716 CLK.n13 VSS 0.00259f
C1717 CLK.n14 VSS 0.00129f
C1718 CLK.n15 VSS 0.0036f
C1719 CLK.n16 VSS 0.00509f
C1720 CLK.n17 VSS 0.0517f
C1721 CLK.n18 VSS 0.0509f
C1722 CLK.n19 VSS 0.0325f
C1723 CLK.t0 VSS 0.0129f
C1724 CLK.t2 VSS 0.00333f
C1725 CLK.n20 VSS 0.0213f
C1726 CLK.n21 VSS 0.00453f
C1727 CLK.n22 VSS 0.00158f
C1728 CLK.n23 VSS 0.0328f
C1729 CLK.n24 VSS 0.00656f
C1730 CLK.n25 VSS 0.00516f
C1731 CLK.n26 VSS 0.00332f
C1732 CLK.n27 VSS 0.00348f
C1733 CLK.n28 VSS 0.00266f
C1734 CLK.n29 VSS 0.00493f
C1735 CLK.n30 VSS 0.1f
C1736 CLK.n31 VSS 0.604f
C1737 CLK.n32 VSS 0.517f
C1738 CLK.n33 VSS 0.175f
C1739 CLK_div_31_mag_0.JK_FF_mag_0.QB.n0 VSS 0.123f
C1740 CLK_div_31_mag_0.JK_FF_mag_0.QB.t5 VSS 0.0265f
C1741 CLK_div_31_mag_0.JK_FF_mag_0.QB.t3 VSS 0.0332f
C1742 CLK_div_31_mag_0.JK_FF_mag_0.QB.n1 VSS 0.0786f
C1743 CLK_div_31_mag_0.JK_FF_mag_0.QB.t6 VSS 0.0297f
C1744 CLK_div_31_mag_0.JK_FF_mag_0.QB.t4 VSS 0.0466f
C1745 CLK_div_31_mag_0.JK_FF_mag_0.QB.n2 VSS 0.0825f
C1746 CLK_div_31_mag_0.JK_FF_mag_0.QB.n3 VSS 0.763f
C1747 CLK_div_31_mag_0.JK_FF_mag_0.QB.t0 VSS 0.0207f
C1748 CLK_div_31_mag_0.JK_FF_mag_0.QB.n4 VSS 0.0207f
C1749 CLK_div_31_mag_0.JK_FF_mag_0.QB.n5 VSS 0.0489f
C1750 RST.t11 VSS 0.0129f
C1751 RST.t10 VSS 0.00851f
C1752 RST.n0 VSS 0.0228f
C1753 RST.n1 VSS 0.0031f
C1754 RST.n2 VSS 0.0019f
C1755 RST.n3 VSS 0.00105f
C1756 RST.n4 VSS 0.00233f
C1757 RST.n5 VSS 0.00143f
C1758 RST.n6 VSS 0.00582f
C1759 RST.n7 VSS 0.0993f
C1760 RST.n8 VSS 0.00422f
C1761 RST.n9 VSS 0.0015f
C1762 RST.n10 VSS 0.00182f
C1763 RST.n11 VSS 0.00397f
C1764 RST.t4 VSS 0.0129f
C1765 RST.t3 VSS 0.00851f
C1766 RST.n12 VSS 0.0228f
C1767 RST.n13 VSS 0.00314f
C1768 RST.n14 VSS 0.00163f
C1769 RST.n15 VSS 0.00117f
C1770 RST.n16 VSS 1.25e-19
C1771 RST.n17 VSS 0.00568f
C1772 RST.n18 VSS 1.25e-19
C1773 RST.n19 VSS 0.0834f
C1774 RST.n20 VSS 0.265f
C1775 RST.t13 VSS 0.00851f
C1776 RST.t6 VSS 0.0129f
C1777 RST.n21 VSS 0.0228f
C1778 RST.n22 VSS 0.004f
C1779 RST.n23 VSS 0.00152f
C1780 RST.n24 VSS 0.0047f
C1781 RST.n25 VSS 0.0056f
C1782 RST.t12 VSS 0.00851f
C1783 RST.t14 VSS 0.0129f
C1784 RST.n26 VSS 0.0229f
C1785 RST.n27 VSS 0.126f
C1786 RST.n28 VSS 0.221f
C1787 RST.n29 VSS 0.0778f
C1788 RST.t5 VSS 0.00851f
C1789 RST.t8 VSS 0.0129f
C1790 RST.n30 VSS 0.0229f
C1791 RST.n31 VSS 0.0609f
C1792 RST.n32 VSS 0.284f
C1793 RST.n33 VSS 0.00383f
C1794 RST.n34 VSS 0.00198f
C1795 RST.t9 VSS 0.013f
C1796 RST.t7 VSS 0.0083f
C1797 RST.n35 VSS 0.0229f
C1798 RST.n36 VSS 0.00294f
C1799 RST.n37 VSS 0.00105f
C1800 RST.n38 VSS 0.0695f
C1801 RST.t15 VSS 0.00851f
C1802 RST.t2 VSS 0.0129f
C1803 RST.n39 VSS 0.0228f
C1804 RST.n40 VSS 0.004f
C1805 RST.n41 VSS 0.00294f
C1806 RST.n42 VSS 0.00137f
C1807 RST.n43 VSS 0.00107f
C1808 RST.n44 VSS 0.0742f
C1809 RST.n45 VSS 0.417f
C1810 RST.n46 VSS 0.0857f
C1811 RST.n47 VSS 0.00876f
C1812 RST.n48 VSS 0.00435f
C1813 RST.n49 VSS 0.0145f
C1814 RST.n50 VSS 0.0501f
C1815 RST.n51 VSS 0.00929f
C1816 RST.n52 VSS 0.00434f
C1817 RST.n53 VSS 0.0532f
C1818 RST.n54 VSS 1.01f
C1819 RST.n55 VSS 1.13f
C1820 RST.n56 VSS 0.32f
C1821 RST.n57 VSS 0.175f
C1822 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.15f
C1823 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.208f
C1824 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.0724f
C1825 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0562f
C1826 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.143f
C1827 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.0449f
C1828 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0563f
C1829 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.145f
C1830 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.079f
C1831 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS 0.0503f
C1832 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.14f
C1833 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 1.2f
C1834 CLK_div_3_mag_0.JK_FF_mag_1.K.t1 VSS 0.0351f
C1835 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 0.0351f
C1836 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.0828f
C1837 CLK_div_31_mag_0.Q4.t8 VSS 0.0156f
C1838 CLK_div_31_mag_0.Q4.t3 VSS 0.0237f
C1839 CLK_div_31_mag_0.Q4.n0 VSS 0.0421f
C1840 CLK_div_31_mag_0.Q4.t6 VSS 0.0136f
C1841 CLK_div_31_mag_0.Q4.t7 VSS 0.0171f
C1842 CLK_div_31_mag_0.Q4.n1 VSS 0.0395f
C1843 CLK_div_31_mag_0.Q4.n2 VSS 0.308f
C1844 CLK_div_31_mag_0.Q4.t4 VSS 0.0389f
C1845 CLK_div_31_mag_0.Q4.t9 VSS 0.00562f
C1846 CLK_div_31_mag_0.Q4.n3 VSS 0.0323f
C1847 CLK_div_31_mag_0.Q4.t2 VSS 0.0136f
C1848 CLK_div_31_mag_0.Q4.t5 VSS 0.0171f
C1849 CLK_div_31_mag_0.Q4.n4 VSS 0.0404f
C1850 CLK_div_31_mag_0.Q4.n5 VSS 1.36f
C1851 CLK_div_31_mag_0.Q4.n6 VSS 0.186f
C1852 CLK_div_31_mag_0.Q1.n0 VSS 0.353f
C1853 CLK_div_31_mag_0.Q1.n1 VSS 0.227f
C1854 CLK_div_31_mag_0.Q1.t2 VSS 0.0191f
C1855 CLK_div_31_mag_0.Q1.t0 VSS 0.0157f
C1856 CLK_div_31_mag_0.Q1.n2 VSS 0.0157f
C1857 CLK_div_31_mag_0.Q1.n3 VSS 0.0378f
C1858 CLK_div_31_mag_0.Q1.t8 VSS 0.035f
C1859 CLK_div_31_mag_0.Q1.t7 VSS 0.0231f
C1860 CLK_div_31_mag_0.Q1.n4 VSS 0.0622f
C1861 CLK_div_31_mag_0.Q1.t3 VSS 0.0201f
C1862 CLK_div_31_mag_0.Q1.t9 VSS 0.0252f
C1863 CLK_div_31_mag_0.Q1.n5 VSS 0.0596f
C1864 CLK_div_31_mag_0.Q1.t10 VSS 0.0201f
C1865 CLK_div_31_mag_0.Q1.t12 VSS 0.0252f
C1866 CLK_div_31_mag_0.Q1.n6 VSS 0.0596f
C1867 CLK_div_31_mag_0.Q1.n7 VSS 1.06f
C1868 CLK_div_31_mag_0.Q1.n8 VSS 0.789f
C1869 CLK_div_31_mag_0.Q1.t13 VSS 0.0251f
C1870 CLK_div_31_mag_0.Q1.t11 VSS 0.0201f
C1871 CLK_div_31_mag_0.Q1.n9 VSS 0.0584f
C1872 CLK_div_31_mag_0.Q1.n10 VSS 0.362f
C1873 CLK_div_31_mag_0.Q1.t5 VSS 0.029f
C1874 CLK_div_31_mag_0.Q1.t6 VSS 0.0074f
C1875 CLK_div_31_mag_0.Q1.n11 VSS 0.048f
C1876 CLK_div_31_mag_0.Q1.t14 VSS 0.0231f
C1877 CLK_div_31_mag_0.Q1.t15 VSS 0.035f
C1878 CLK_div_31_mag_0.Q1.n12 VSS 0.0619f
C1879 CLK_div_31_mag_0.Q1.t4 VSS 0.0231f
C1880 CLK_div_31_mag_0.Q1.t16 VSS 0.035f
C1881 CLK_div_31_mag_0.Q1.n13 VSS 0.0619f
C1882 CLK_div_31_mag_0.Q3.n0 VSS 0.651f
C1883 CLK_div_31_mag_0.Q3.n1 VSS 0.242f
C1884 CLK_div_31_mag_0.Q3.t15 VSS 0.0256f
C1885 CLK_div_31_mag_0.Q3.t2 VSS 0.0388f
C1886 CLK_div_31_mag_0.Q3.n2 VSS 0.0689f
C1887 CLK_div_31_mag_0.Q3.t5 VSS 0.0223f
C1888 CLK_div_31_mag_0.Q3.t9 VSS 0.0279f
C1889 CLK_div_31_mag_0.Q3.n3 VSS 0.0646f
C1890 CLK_div_31_mag_0.Q3.n4 VSS 0.499f
C1891 CLK_div_31_mag_0.Q3.t10 VSS 0.0223f
C1892 CLK_div_31_mag_0.Q3.t14 VSS 0.0279f
C1893 CLK_div_31_mag_0.Q3.n5 VSS 0.0726f
C1894 CLK_div_31_mag_0.Q3.t8 VSS 0.0223f
C1895 CLK_div_31_mag_0.Q3.t4 VSS 0.0279f
C1896 CLK_div_31_mag_0.Q3.n6 VSS 0.0661f
C1897 CLK_div_31_mag_0.Q3.n7 VSS 0.67f
C1898 CLK_div_31_mag_0.Q3.t3 VSS 0.0256f
C1899 CLK_div_31_mag_0.Q3.t7 VSS 0.0388f
C1900 CLK_div_31_mag_0.Q3.n8 VSS 0.0686f
C1901 CLK_div_31_mag_0.Q3.t11 VSS 0.0256f
C1902 CLK_div_31_mag_0.Q3.t13 VSS 0.0388f
C1903 CLK_div_31_mag_0.Q3.n9 VSS 0.0686f
C1904 CLK_div_31_mag_0.Q3.n10 VSS 0.276f
C1905 CLK_div_31_mag_0.Q3.t6 VSS 0.0321f
C1906 CLK_div_31_mag_0.Q3.t12 VSS 0.0082f
C1907 CLK_div_31_mag_0.Q3.n11 VSS 0.0531f
C1908 CLK_div_31_mag_0.Q3.n12 VSS 0.204f
C1909 VDD.n0 VSS 0.275f
C1910 VDD.t4 VSS 0.00226f
C1911 VDD.n1 VSS 0.00226f
C1912 VDD.n2 VSS 0.0049f
C1913 VDD.t232 VSS 0.00547f
C1914 VDD.n3 VSS 0.00546f
C1915 VDD.t338 VSS 0.00547f
C1916 VDD.n4 VSS 0.00546f
C1917 VDD.t201 VSS 0.00547f
C1918 VDD.n5 VSS 0.0264f
C1919 VDD.n6 VSS 0.254f
C1920 VDD.t315 VSS 0.00547f
C1921 VDD.t460 VSS 0.00547f
C1922 VDD.n7 VSS 0.0363f
C1923 VDD.t314 VSS 0.0485f
C1924 VDD.t311 VSS 0.0376f
C1925 VDD.t404 VSS 0.00226f
C1926 VDD.n8 VSS 0.00226f
C1927 VDD.n9 VSS 0.00493f
C1928 VDD.t93 VSS 0.0055f
C1929 VDD.n10 VSS 0.00549f
C1930 VDD.n11 VSS 0.0272f
C1931 VDD.t387 VSS 0.0725f
C1932 VDD.n12 VSS 0.00549f
C1933 VDD.t346 VSS 0.0055f
C1934 VDD.n13 VSS 0.00549f
C1935 VDD.n14 VSS 0.00549f
C1936 VDD.t305 VSS 0.0715f
C1937 VDD.n15 VSS 0.0341f
C1938 VDD.t294 VSS 0.0055f
C1939 VDD.n16 VSS 0.00549f
C1940 VDD.t293 VSS 0.0662f
C1941 VDD.t384 VSS 0.0725f
C1942 VDD.n17 VSS 0.0341f
C1943 VDD.t363 VSS 0.0055f
C1944 VDD.t348 VSS 0.00226f
C1945 VDD.n18 VSS 0.00226f
C1946 VDD.n19 VSS 0.00493f
C1947 VDD.t362 VSS 0.0662f
C1948 VDD.t347 VSS 0.0809f
C1949 VDD.t187 VSS 0.0376f
C1950 VDD.n20 VSS 0.0341f
C1951 VDD.t32 VSS 0.0055f
C1952 VDD.t304 VSS 0.00226f
C1953 VDD.n21 VSS 0.00226f
C1954 VDD.n22 VSS 0.00493f
C1955 VDD.t31 VSS 0.0662f
C1956 VDD.t303 VSS 0.0809f
C1957 VDD.t324 VSS 0.0376f
C1958 VDD.t40 VSS 0.066f
C1959 VDD.n23 VSS 0.0341f
C1960 VDD.t41 VSS 0.00589f
C1961 VDD.n24 VSS 0.0423f
C1962 VDD.n25 VSS 0.0313f
C1963 VDD.n26 VSS 0.0321f
C1964 VDD.n27 VSS 0.017f
C1965 VDD.n28 VSS 0.0313f
C1966 VDD.n29 VSS 0.032f
C1967 VDD.n30 VSS 0.019f
C1968 VDD.n31 VSS 0.0272f
C1969 VDD.n32 VSS 0.0253f
C1970 VDD.n33 VSS 0.019f
C1971 VDD.n34 VSS 0.0518f
C1972 VDD.n35 VSS 0.0589f
C1973 VDD.t149 VSS 0.0715f
C1974 VDD.t345 VSS 0.0662f
C1975 VDD.n36 VSS 0.0341f
C1976 VDD.n37 VSS 0.019f
C1977 VDD.n38 VSS 0.0253f
C1978 VDD.n39 VSS 0.0272f
C1979 VDD.t350 VSS 0.0055f
C1980 VDD.n40 VSS 0.0253f
C1981 VDD.n41 VSS 0.019f
C1982 VDD.n42 VSS 0.0341f
C1983 VDD.t349 VSS 0.0662f
C1984 VDD.t364 VSS 0.0725f
C1985 VDD.t403 VSS 0.0809f
C1986 VDD.t92 VSS 0.0662f
C1987 VDD.n43 VSS 0.0341f
C1988 VDD.n44 VSS 0.019f
C1989 VDD.n45 VSS 0.024f
C1990 VDD.n46 VSS 0.0208f
C1991 VDD.n47 VSS 0.0213f
C1992 VDD.t323 VSS 0.00548f
C1993 VDD.n48 VSS 0.00547f
C1994 VDD.t465 VSS 0.00547f
C1995 VDD.n49 VSS 0.0172f
C1996 VDD.t279 VSS 0.0055f
C1997 VDD.t278 VSS 0.0487f
C1998 VDD.n50 VSS 0.0564f
C1999 VDD.t308 VSS 0.0492f
C2000 VDD.n51 VSS 0.0332f
C2001 VDD.t148 VSS 0.0131f
C2002 VDD.t464 VSS 0.0494f
C2003 VDD.t147 VSS 0.0467f
C2004 VDD.n52 VSS 0.0856f
C2005 VDD.n53 VSS 0.0377f
C2006 VDD.n54 VSS 0.0162f
C2007 VDD.n55 VSS 0.162f
C2008 VDD.n56 VSS 0.775f
C2009 VDD.n57 VSS 0.125f
C2010 VDD.n58 VSS 0.0268f
C2011 VDD.t461 VSS 0.0433f
C2012 VDD.t322 VSS 0.066f
C2013 VDD.n59 VSS 0.0341f
C2014 VDD.n60 VSS 0.0205f
C2015 VDD.n61 VSS 0.0209f
C2016 VDD.n62 VSS 0.146f
C2017 VDD.n63 VSS 0.00887f
C2018 VDD.n64 VSS 0.0372f
C2019 VDD.n65 VSS 0.0149f
C2020 VDD.n66 VSS 0.0122f
C2021 VDD.n67 VSS 0.0341f
C2022 VDD.t459 VSS 0.0376f
C2023 VDD.n68 VSS 0.051f
C2024 VDD.n69 VSS 0.0265f
C2025 VDD.n70 VSS 0.00549f
C2026 VDD.t454 VSS 0.0715f
C2027 VDD.n71 VSS 0.0341f
C2028 VDD.t217 VSS 0.0055f
C2029 VDD.n72 VSS 0.00549f
C2030 VDD.t216 VSS 0.0662f
C2031 VDD.t108 VSS 0.0725f
C2032 VDD.n73 VSS 0.0341f
C2033 VDD.t256 VSS 0.0055f
C2034 VDD.t340 VSS 0.00226f
C2035 VDD.n74 VSS 0.00226f
C2036 VDD.n75 VSS 0.00493f
C2037 VDD.t255 VSS 0.0662f
C2038 VDD.t339 VSS 0.0809f
C2039 VDD.t228 VSS 0.0376f
C2040 VDD.n76 VSS 0.0341f
C2041 VDD.t277 VSS 0.0055f
C2042 VDD.t458 VSS 0.00226f
C2043 VDD.n77 VSS 0.00226f
C2044 VDD.n78 VSS 0.00493f
C2045 VDD.t276 VSS 0.0662f
C2046 VDD.t457 VSS 0.0809f
C2047 VDD.t316 VSS 0.0376f
C2048 VDD.t49 VSS 0.066f
C2049 VDD.n79 VSS 0.0341f
C2050 VDD.t50 VSS 0.00513f
C2051 VDD.t39 VSS 0.00471f
C2052 VDD.t474 VSS 0.00357f
C2053 VDD.n80 VSS 0.0092f
C2054 VDD.n81 VSS 0.0516f
C2055 VDD.n82 VSS 0.0675f
C2056 VDD.n83 VSS 0.0012f
C2057 VDD.t484 VSS 0.00356f
C2058 VDD.n84 VSS 0.00483f
C2059 VDD.t48 VSS 0.00458f
C2060 VDD.n85 VSS 0.00452f
C2061 VDD.n86 VSS 4.56e-20
C2062 VDD.n87 VSS 0.00142f
C2063 VDD.n88 VSS 6.54e-19
C2064 VDD.n89 VSS 5.43e-19
C2065 VDD.n90 VSS 0.00409f
C2066 VDD.n91 VSS 0.0128f
C2067 VDD.n92 VSS 0.0314f
C2068 VDD.n93 VSS 0.0313f
C2069 VDD.n94 VSS 0.0321f
C2070 VDD.n95 VSS 0.017f
C2071 VDD.n96 VSS 0.0313f
C2072 VDD.n97 VSS 0.032f
C2073 VDD.n98 VSS 0.019f
C2074 VDD.n99 VSS 0.0272f
C2075 VDD.n100 VSS 0.0253f
C2076 VDD.n101 VSS 0.019f
C2077 VDD.n102 VSS 0.0474f
C2078 VDD.n103 VSS 0.00546f
C2079 VDD.t0 VSS 0.0577f
C2080 VDD.t200 VSS 0.0527f
C2081 VDD.n104 VSS 0.0294f
C2082 VDD.n105 VSS 0.0224f
C2083 VDD.n106 VSS 0.0339f
C2084 VDD.n107 VSS 0.0379f
C2085 VDD.n108 VSS 0.143f
C2086 VDD.n109 VSS 0.28f
C2087 VDD.n110 VSS 0.265f
C2088 VDD.n111 VSS 0.144f
C2089 VDD.n112 VSS 0.0257f
C2090 VDD.t105 VSS 0.0577f
C2091 VDD.t337 VSS 0.039f
C2092 VDD.n113 VSS 0.0294f
C2093 VDD.n114 VSS 0.0224f
C2094 VDD.n115 VSS 0.032f
C2095 VDD.n116 VSS 0.03f
C2096 VDD.n117 VSS 0.14f
C2097 VDD.n118 VSS 0.151f
C2098 VDD.t257 VSS 0.0253f
C2099 VDD.t231 VSS 0.0527f
C2100 VDD.n119 VSS 0.0294f
C2101 VDD.n120 VSS 0.0161f
C2102 VDD.n121 VSS 0.0301f
C2103 VDD.n122 VSS 0.0291f
C2104 VDD.n123 VSS 0.0129f
C2105 VDD.t402 VSS 0.00547f
C2106 VDD.t3 VSS 0.0643f
C2107 VDD.t319 VSS 0.0299f
C2108 VDD.n124 VSS 0.0294f
C2109 VDD.t401 VSS 0.0299f
C2110 VDD.n125 VSS 0.0841f
C2111 VDD.t327 VSS 0.0605f
C2112 VDD.t328 VSS 0.00566f
C2113 VDD.n126 VSS 0.0356f
C2114 VDD.n127 VSS 0.136f
C2115 VDD.n128 VSS 0.564f
C2116 VDD.n129 VSS 0.494f
C2117 VDD.t94 VSS 0.049f
C2118 VDD.n130 VSS 0.0507f
C2119 VDD.t95 VSS 0.00547f
C2120 VDD.n131 VSS 0.00549f
C2121 VDD.t169 VSS 0.0433f
C2122 VDD.n132 VSS 0.0341f
C2123 VDD.t373 VSS 0.0055f
C2124 VDD.n133 VSS 0.21f
C2125 VDD.t372 VSS 0.0645f
C2126 VDD.t99 VSS 0.0482f
C2127 VDD.n134 VSS 0.0527f
C2128 VDD.t100 VSS 0.00547f
C2129 VDD.n135 VSS 0.00549f
C2130 VDD.t122 VSS 0.0433f
C2131 VDD.n136 VSS 0.0341f
C2132 VDD.t438 VSS 0.0055f
C2133 VDD.n137 VSS 0.166f
C2134 VDD.t437 VSS 0.0656f
C2135 VDD.t238 VSS 0.0467f
C2136 VDD.n138 VSS 0.0508f
C2137 VDD.t239 VSS 0.00547f
C2138 VDD.n139 VSS 0.00549f
C2139 VDD.t374 VSS 0.0433f
C2140 VDD.n140 VSS 0.0341f
C2141 VDD.t356 VSS 0.0055f
C2142 VDD.t355 VSS 0.0657f
C2143 VDD.t447 VSS 0.0461f
C2144 VDD.n141 VSS 0.0504f
C2145 VDD.t448 VSS 0.00547f
C2146 VDD.n142 VSS 0.00549f
C2147 VDD.t208 VSS 0.0433f
C2148 VDD.t428 VSS 0.066f
C2149 VDD.n143 VSS 0.0341f
C2150 VDD.t429 VSS 0.00582f
C2151 VDD.n144 VSS 0.0223f
C2152 VDD.n145 VSS 0.0336f
C2153 VDD.n146 VSS 0.0295f
C2154 VDD.n147 VSS 0.0344f
C2155 VDD.n148 VSS 0.0225f
C2156 VDD.n149 VSS 0.0342f
C2157 VDD.n150 VSS 0.03f
C2158 VDD.n151 VSS 0.0294f
C2159 VDD.n152 VSS 0.034f
C2160 VDD.n153 VSS 0.0231f
C2161 VDD.n154 VSS 0.0355f
C2162 VDD.n155 VSS 0.0309f
C2163 VDD.n156 VSS 0.0313f
C2164 VDD.n157 VSS 0.0357f
C2165 VDD.n158 VSS 0.0225f
C2166 VDD.n159 VSS 0.0342f
C2167 VDD.n160 VSS 0.03f
C2168 VDD.t29 VSS 0.0517f
C2169 VDD.n161 VSS 0.0581f
C2170 VDD.t30 VSS 0.00547f
C2171 VDD.t435 VSS 0.0509f
C2172 VDD.n162 VSS 0.0586f
C2173 VDD.t436 VSS 0.00547f
C2174 VDD.n163 VSS 0.00549f
C2175 VDD.t21 VSS 0.0722f
C2176 VDD.n164 VSS 0.0341f
C2177 VDD.t416 VSS 0.0055f
C2178 VDD.t415 VSS 0.0645f
C2179 VDD.t177 VSS 0.0483f
C2180 VDD.n165 VSS 0.0527f
C2181 VDD.t178 VSS 0.00547f
C2182 VDD.n166 VSS 0.00549f
C2183 VDD.t87 VSS 0.0433f
C2184 VDD.n167 VSS 0.0341f
C2185 VDD.t418 VSS 0.00554f
C2186 VDD.t281 VSS 0.0055f
C2187 VDD.n168 VSS 0.0392f
C2188 VDD.t243 VSS 0.0055f
C2189 VDD.t163 VSS 0.0715f
C2190 VDD.n169 VSS 0.02f
C2191 VDD.n170 VSS 0.0372f
C2192 VDD.t162 VSS 0.00226f
C2193 VDD.n171 VSS 0.00226f
C2194 VDD.n172 VSS 0.00493f
C2195 VDD.t427 VSS 0.0055f
C2196 VDD.t248 VSS 0.0055f
C2197 VDD.n173 VSS 0.00549f
C2198 VDD.n174 VSS 0.0281f
C2199 VDD.n175 VSS 0.0349f
C2200 VDD.t417 VSS 0.0656f
C2201 VDD.t280 VSS 0.0468f
C2202 VDD.n176 VSS 0.0508f
C2203 VDD.t133 VSS 0.0433f
C2204 VDD.n177 VSS 0.00549f
C2205 VDD.n178 VSS 0.00549f
C2206 VDD.n179 VSS 0.0357f
C2207 VDD.n180 VSS 0.035f
C2208 VDD.n181 VSS 0.0284f
C2209 VDD.n182 VSS 0.0341f
C2210 VDD.t240 VSS 0.0657f
C2211 VDD.t329 VSS 0.0462f
C2212 VDD.t330 VSS 0.00791f
C2213 VDD.t153 VSS 0.0055f
C2214 VDD.t241 VSS 0.0055f
C2215 VDD.n183 VSS 0.0284f
C2216 VDD.n184 VSS 0.0501f
C2217 VDD.n185 VSS 0.0106f
C2218 VDD.n186 VSS 0.00549f
C2219 VDD.n187 VSS 0.036f
C2220 VDD.n188 VSS 0.0504f
C2221 VDD.t244 VSS 0.0433f
C2222 VDD.t426 VSS 0.066f
C2223 VDD.n189 VSS 0.0341f
C2224 VDD.n190 VSS 0.0365f
C2225 VDD.n191 VSS 0.036f
C2226 VDD.n192 VSS 0.0403f
C2227 VDD.n193 VSS 0.0248f
C2228 VDD.t47 VSS 0.0055f
C2229 VDD.n194 VSS 0.0548f
C2230 VDD.t86 VSS 0.00547f
C2231 VDD.n195 VSS 0.00549f
C2232 VDD.t82 VSS 0.0715f
C2233 VDD.n196 VSS 0.0341f
C2234 VDD.t352 VSS 0.0055f
C2235 VDD.n197 VSS 0.00549f
C2236 VDD.t351 VSS 0.0662f
C2237 VDD.t141 VSS 0.0725f
C2238 VDD.n198 VSS 0.0341f
C2239 VDD.t302 VSS 0.0055f
C2240 VDD.t252 VSS 0.00226f
C2241 VDD.n199 VSS 0.00226f
C2242 VDD.n200 VSS 0.00493f
C2243 VDD.t301 VSS 0.0662f
C2244 VDD.t251 VSS 0.0809f
C2245 VDD.t225 VSS 0.0376f
C2246 VDD.n201 VSS 0.0341f
C2247 VDD.t354 VSS 0.0055f
C2248 VDD.t381 VSS 0.00226f
C2249 VDD.n202 VSS 0.00226f
C2250 VDD.n203 VSS 0.00493f
C2251 VDD.t353 VSS 0.0662f
C2252 VDD.t380 VSS 0.0809f
C2253 VDD.t125 VSS 0.0376f
C2254 VDD.t56 VSS 0.066f
C2255 VDD.n204 VSS 0.0341f
C2256 VDD.t57 VSS 0.0055f
C2257 VDD.t42 VSS 0.00471f
C2258 VDD.t473 VSS 0.00357f
C2259 VDD.n205 VSS 0.00925f
C2260 VDD.n206 VSS 0.00867f
C2261 VDD.t55 VSS 0.00471f
C2262 VDD.t486 VSS 0.00357f
C2263 VDD.n207 VSS 0.00927f
C2264 VDD.n208 VSS 0.00696f
C2265 VDD.n209 VSS 0.0362f
C2266 VDD.n210 VSS 0.0256f
C2267 VDD.n211 VSS 0.017f
C2268 VDD.n212 VSS 0.0313f
C2269 VDD.n213 VSS 0.0321f
C2270 VDD.n214 VSS 0.017f
C2271 VDD.n215 VSS 0.0313f
C2272 VDD.n216 VSS 0.032f
C2273 VDD.n217 VSS 0.019f
C2274 VDD.n218 VSS 0.0272f
C2275 VDD.n219 VSS 0.0253f
C2276 VDD.n220 VSS 0.019f
C2277 VDD.n221 VSS 0.0489f
C2278 VDD.t166 VSS 0.0486f
C2279 VDD.n222 VSS 0.051f
C2280 VDD.n223 VSS 0.00689f
C2281 VDD.n224 VSS 0.00549f
C2282 VDD.t24 VSS 0.0715f
C2283 VDD.n225 VSS 0.0341f
C2284 VDD.n226 VSS 0.0055f
C2285 VDD.t140 VSS 0.0055f
C2286 VDD.t59 VSS 0.0377f
C2287 VDD.n227 VSS 0.0341f
C2288 VDD.n228 VSS 0.00549f
C2289 VDD.t112 VSS 0.00226f
C2290 VDD.n229 VSS 0.00226f
C2291 VDD.n230 VSS 0.00493f
C2292 VDD.t139 VSS 0.0662f
C2293 VDD.t144 VSS 0.0725f
C2294 VDD.n231 VSS 0.0341f
C2295 VDD.t250 VSS 0.0055f
C2296 VDD.n232 VSS 0.0055f
C2297 VDD.n233 VSS 0.00549f
C2298 VDD.t111 VSS 0.0374f
C2299 VDD.t5 VSS 0.0809f
C2300 VDD.t265 VSS 0.0664f
C2301 VDD.n234 VSS 0.0341f
C2302 VDD.t249 VSS 0.0662f
C2303 VDD.t298 VSS 0.0725f
C2304 VDD.n235 VSS 0.0341f
C2305 VDD.t215 VSS 0.00549f
C2306 VDD.t221 VSS 0.0055f
C2307 VDD.n236 VSS 0.0055f
C2308 VDD.t214 VSS 0.0724f
C2309 VDD.t398 VSS 0.0664f
C2310 VDD.n237 VSS 0.0341f
C2311 VDD.t28 VSS 0.00226f
C2312 VDD.n238 VSS 0.00226f
C2313 VDD.n239 VSS 0.00493f
C2314 VDD.t102 VSS 0.00549f
C2315 VDD.t220 VSS 0.0662f
C2316 VDD.t27 VSS 0.0809f
C2317 VDD.t136 VSS 0.0376f
C2318 VDD.n240 VSS 0.0341f
C2319 VDD.n241 VSS 0.0055f
C2320 VDD.t44 VSS 0.0055f
C2321 VDD.t101 VSS 0.0724f
C2322 VDD.t392 VSS 0.0664f
C2323 VDD.t8 VSS 0.0714f
C2324 VDD.n242 VSS 0.0341f
C2325 VDD.t9 VSS 0.00549f
C2326 VDD.t121 VSS 0.00691f
C2327 VDD.t120 VSS 0.0485f
C2328 VDD.t43 VSS 0.0376f
C2329 VDD.n243 VSS 0.051f
C2330 VDD.n244 VSS 0.00549f
C2331 VDD.t128 VSS 0.0715f
C2332 VDD.n245 VSS 0.0341f
C2333 VDD.t173 VSS 0.0055f
C2334 VDD.n246 VSS 0.00549f
C2335 VDD.t172 VSS 0.0662f
C2336 VDD.t271 VSS 0.0725f
C2337 VDD.n247 VSS 0.0341f
C2338 VDD.t470 VSS 0.0055f
C2339 VDD.t334 VSS 0.00226f
C2340 VDD.n248 VSS 0.00226f
C2341 VDD.n249 VSS 0.00493f
C2342 VDD.t469 VSS 0.0662f
C2343 VDD.t333 VSS 0.0809f
C2344 VDD.t184 VSS 0.0376f
C2345 VDD.n250 VSS 0.0341f
C2346 VDD.t391 VSS 0.0055f
C2347 VDD.t132 VSS 0.00226f
C2348 VDD.n251 VSS 0.00226f
C2349 VDD.n252 VSS 0.00493f
C2350 VDD.t390 VSS 0.0662f
C2351 VDD.t131 VSS 0.0809f
C2352 VDD.t197 VSS 0.0376f
C2353 VDD.t63 VSS 0.066f
C2354 VDD.n253 VSS 0.0341f
C2355 VDD.t64 VSS 0.0055f
C2356 VDD.t65 VSS 0.00471f
C2357 VDD.t472 VSS 0.00357f
C2358 VDD.n254 VSS 0.00926f
C2359 VDD.n255 VSS 0.00765f
C2360 VDD.t62 VSS 0.00471f
C2361 VDD.t482 VSS 0.00357f
C2362 VDD.n256 VSS 0.00926f
C2363 VDD.n257 VSS 0.00736f
C2364 VDD.n258 VSS 0.0377f
C2365 VDD.n259 VSS 0.0256f
C2366 VDD.n260 VSS 0.017f
C2367 VDD.n261 VSS 0.0313f
C2368 VDD.n262 VSS 0.0321f
C2369 VDD.n263 VSS 0.017f
C2370 VDD.n264 VSS 0.0313f
C2371 VDD.n265 VSS 0.032f
C2372 VDD.n266 VSS 0.019f
C2373 VDD.n267 VSS 0.0272f
C2374 VDD.n268 VSS 0.0253f
C2375 VDD.n269 VSS 0.019f
C2376 VDD.n270 VSS 0.0496f
C2377 VDD.t421 VSS 0.0486f
C2378 VDD.n271 VSS 0.051f
C2379 VDD.n272 VSS 0.00689f
C2380 VDD.n273 VSS 0.00549f
C2381 VDD.t449 VSS 0.0577f
C2382 VDD.n274 VSS 0.0294f
C2383 VDD.n275 VSS 0.0055f
C2384 VDD.t254 VSS 0.0055f
C2385 VDD.t76 VSS 0.0377f
C2386 VDD.n276 VSS 0.0341f
C2387 VDD.n277 VSS 0.00549f
C2388 VDD.t431 VSS 0.00226f
C2389 VDD.n278 VSS 0.00226f
C2390 VDD.n279 VSS 0.00493f
C2391 VDD.t253 VSS 0.0527f
C2392 VDD.t268 VSS 0.0577f
C2393 VDD.n280 VSS 0.0294f
C2394 VDD.t336 VSS 0.0055f
C2395 VDD.n281 VSS 0.0055f
C2396 VDD.n282 VSS 0.00549f
C2397 VDD.t430 VSS 0.0374f
C2398 VDD.t262 VSS 0.0809f
C2399 VDD.t181 VSS 0.0664f
C2400 VDD.n283 VSS 0.0341f
C2401 VDD.n284 VSS 0.0294f
C2402 VDD.t160 VSS 0.00549f
C2403 VDD.t310 VSS 0.0055f
C2404 VDD.n285 VSS 0.0055f
C2405 VDD.t159 VSS 0.0724f
C2406 VDD.t444 VSS 0.0664f
C2407 VDD.n286 VSS 0.0341f
C2408 VDD.t453 VSS 0.00226f
C2409 VDD.n287 VSS 0.00226f
C2410 VDD.n288 VSS 0.00493f
C2411 VDD.t344 VSS 0.00549f
C2412 VDD.t309 VSS 0.0527f
C2413 VDD.t452 VSS 0.0643f
C2414 VDD.t13 VSS 0.0299f
C2415 VDD.n289 VSS 0.0294f
C2416 VDD.n290 VSS 0.0055f
C2417 VDD.t67 VSS 0.0055f
C2418 VDD.t343 VSS 0.0724f
C2419 VDD.t174 VSS 0.0664f
C2420 VDD.t260 VSS 0.0714f
C2421 VDD.n291 VSS 0.0341f
C2422 VDD.t261 VSS 0.00549f
C2423 VDD.t17 VSS 0.00691f
C2424 VDD.t66 VSS 0.0299f
C2425 VDD.t335 VSS 0.039f
C2426 VDD.t466 VSS 0.0253f
C2427 VDD.n292 VSS 0.152f
C2428 VDD.n293 VSS 0.0842f
C2429 VDD.t16 VSS 0.0605f
C2430 VDD.t196 VSS 0.00549f
C2431 VDD.t156 VSS 0.0664f
C2432 VDD.n294 VSS 0.0055f
C2433 VDD.t91 VSS 0.00226f
C2434 VDD.n295 VSS 0.00226f
C2435 VDD.n296 VSS 0.00493f
C2436 VDD.n297 VSS 0.0055f
C2437 VDD.n298 VSS 0.0321f
C2438 VDD.t72 VSS 0.0662f
C2439 VDD.n299 VSS 0.0055f
C2440 VDD.t477 VSS 0.00357f
C2441 VDD.t71 VSS 0.00471f
C2442 VDD.n300 VSS 0.00927f
C2443 VDD.t475 VSS 0.00357f
C2444 VDD.t75 VSS 0.00471f
C2445 VDD.n301 VSS 0.0092f
C2446 VDD.n302 VSS 0.0014f
C2447 VDD.n303 VSS 0.00834f
C2448 VDD.n304 VSS 0.0455f
C2449 VDD.n305 VSS 0.0256f
C2450 VDD.t425 VSS 0.00226f
C2451 VDD.n306 VSS 0.00226f
C2452 VDD.n307 VSS 0.00493f
C2453 VDD.n308 VSS 0.0313f
C2454 VDD.n309 VSS 0.017f
C2455 VDD.n310 VSS 0.0341f
C2456 VDD.t424 VSS 0.0374f
C2457 VDD.t18 VSS 0.0809f
C2458 VDD.t369 VSS 0.0664f
C2459 VDD.t441 VSS 0.0809f
C2460 VDD.t90 VSS 0.0374f
C2461 VDD.n311 VSS 0.0341f
C2462 VDD.n312 VSS 0.017f
C2463 VDD.n313 VSS 0.0313f
C2464 VDD.n314 VSS 0.032f
C2465 VDD.t342 VSS 0.00549f
C2466 VDD.n315 VSS 0.0055f
C2467 VDD.n316 VSS 0.0253f
C2468 VDD.n317 VSS 0.0272f
C2469 VDD.n318 VSS 0.019f
C2470 VDD.n319 VSS 0.0341f
C2471 VDD.t341 VSS 0.0724f
C2472 VDD.t359 VSS 0.0664f
C2473 VDD.t195 VSS 0.0714f
C2474 VDD.n320 VSS 0.0341f
C2475 VDD.n321 VSS 0.019f
C2476 VDD.n322 VSS 0.0513f
C2477 VDD.n323 VSS 0.0124f
C2478 VDD.n324 VSS 0.0327f
C2479 VDD.n325 VSS 0.0337f
C2480 VDD.n326 VSS 0.0257f
C2481 VDD.n327 VSS 0.0261f
C2482 VDD.n328 VSS 0.0271f
C2483 VDD.n329 VSS 0.0313f
C2484 VDD.n330 VSS 0.0289f
C2485 VDD.n331 VSS 0.025f
C2486 VDD.n332 VSS 0.0348f
C2487 VDD.n333 VSS 0.0386f
C2488 VDD.n334 VSS 0.0257f
C2489 VDD.n335 VSS 0.0278f
C2490 VDD.n336 VSS 0.0279f
C2491 VDD.n337 VSS 0.0256f
C2492 VDD.n338 VSS 0.0386f
C2493 VDD.n339 VSS 0.0349f
C2494 VDD.n340 VSS 0.0249f
C2495 VDD.n341 VSS 0.0289f
C2496 VDD.n342 VSS 0.0314f
C2497 VDD.n343 VSS 0.027f
C2498 VDD.n344 VSS 0.0261f
C2499 VDD.n345 VSS 0.0258f
C2500 VDD.n346 VSS 0.0336f
C2501 VDD.n347 VSS 0.0328f
C2502 VDD.n348 VSS 0.0125f
C2503 VDD.n349 VSS 0.0593f
C2504 VDD.t420 VSS 0.00549f
C2505 VDD.t211 VSS 0.0664f
C2506 VDD.n350 VSS 0.0055f
C2507 VDD.t191 VSS 0.00226f
C2508 VDD.n351 VSS 0.00226f
C2509 VDD.n352 VSS 0.00493f
C2510 VDD.n353 VSS 0.0055f
C2511 VDD.n354 VSS 0.0321f
C2512 VDD.t52 VSS 0.0662f
C2513 VDD.n355 VSS 0.0055f
C2514 VDD.t483 VSS 0.00357f
C2515 VDD.t51 VSS 0.00471f
C2516 VDD.n356 VSS 0.00925f
C2517 VDD.n357 VSS 0.00258f
C2518 VDD.t478 VSS 0.00357f
C2519 VDD.t58 VSS 0.00471f
C2520 VDD.n358 VSS 0.00923f
C2521 VDD.n359 VSS 0.00753f
C2522 VDD.n360 VSS 0.041f
C2523 VDD.n361 VSS 0.0256f
C2524 VDD.t114 VSS 0.00226f
C2525 VDD.n362 VSS 0.00226f
C2526 VDD.n363 VSS 0.00493f
C2527 VDD.n364 VSS 0.0313f
C2528 VDD.n365 VSS 0.017f
C2529 VDD.n366 VSS 0.0341f
C2530 VDD.t113 VSS 0.0374f
C2531 VDD.t432 VSS 0.0809f
C2532 VDD.t235 VSS 0.0664f
C2533 VDD.t395 VSS 0.0809f
C2534 VDD.t190 VSS 0.0374f
C2535 VDD.n367 VSS 0.0341f
C2536 VDD.n368 VSS 0.017f
C2537 VDD.n369 VSS 0.0313f
C2538 VDD.n370 VSS 0.032f
C2539 VDD.t104 VSS 0.00549f
C2540 VDD.n371 VSS 0.0055f
C2541 VDD.n372 VSS 0.0253f
C2542 VDD.n373 VSS 0.0272f
C2543 VDD.n374 VSS 0.019f
C2544 VDD.n375 VSS 0.0341f
C2545 VDD.t103 VSS 0.0724f
C2546 VDD.t192 VSS 0.0664f
C2547 VDD.t419 VSS 0.0714f
C2548 VDD.n376 VSS 0.0341f
C2549 VDD.n377 VSS 0.019f
C2550 VDD.n378 VSS 0.0488f
C2551 VDD.n379 VSS 0.0565f
C2552 VDD.n380 VSS 0.0144f
C2553 VDD.n381 VSS 0.0343f
C2554 VDD.n382 VSS 0.0332f
C2555 VDD.n383 VSS 0.0253f
C2556 VDD.n384 VSS 0.0257f
C2557 VDD.n385 VSS 0.0246f
C2558 VDD.n386 VSS 0.0308f
C2559 VDD.n387 VSS 0.0284f
C2560 VDD.n388 VSS 0.0269f
C2561 VDD.n389 VSS 0.0342f
C2562 VDD.n390 VSS 0.038f
C2563 VDD.n391 VSS 0.0253f
C2564 VDD.n392 VSS 0.0296f
C2565 VDD.n393 VSS 0.0297f
C2566 VDD.n394 VSS 0.0252f
C2567 VDD.n395 VSS 0.038f
C2568 VDD.n396 VSS 0.0343f
C2569 VDD.n397 VSS 0.0267f
C2570 VDD.n398 VSS 0.0284f
C2571 VDD.n399 VSS 0.0309f
C2572 VDD.n400 VSS 0.0245f
C2573 VDD.n401 VSS 0.0257f
C2574 VDD.n402 VSS 0.0255f
C2575 VDD.n403 VSS 0.0331f
C2576 VDD.n404 VSS 0.0344f
C2577 VDD.n405 VSS 0.0146f
C2578 VDD.n406 VSS 0.0582f
C2579 VDD.n407 VSS 0.0529f
C2580 VDD.t85 VSS 0.0485f
C2581 VDD.n408 VSS 0.051f
C2582 VDD.t46 VSS 0.0376f
C2583 VDD.n409 VSS 0.0341f
C2584 VDD.t377 VSS 0.0376f
C2585 VDD.t161 VSS 0.0809f
C2586 VDD.t247 VSS 0.0662f
C2587 VDD.n410 VSS 0.0341f
C2588 VDD.t115 VSS 0.0725f
C2589 VDD.t152 VSS 0.0662f
C2590 VDD.n411 VSS 0.0341f
C2591 VDD.t202 VSS 0.0725f
C2592 VDD.t242 VSS 0.0662f
C2593 VDD.n412 VSS 0.0341f
C2594 VDD.n413 VSS 0.0162f
C2595 VDD.n414 VSS 0.0151f
C2596 VDD.n415 VSS 0.00523f
C2597 VDD.n416 VSS 0.00802f
C2598 VDD.t440 VSS 0.00547f
C2599 VDD.n417 VSS 0.00547f
C2600 VDD.n418 VSS 0.0301f
C2601 VDD.t287 VSS 0.0753f
C2602 VDD.n419 VSS 0.00547f
C2603 VDD.t286 VSS 0.00547f
C2604 VDD.n420 VSS 0.00547f
C2605 VDD.n421 VSS 0.03f
C2606 VDD.t285 VSS 0.0918f
C2607 VDD.n422 VSS 0.0375f
C2608 VDD.t36 VSS 0.0918f
C2609 VDD.n423 VSS 0.0784f
C2610 VDD.n424 VSS 0.0788f
C2611 VDD.n425 VSS 0.00547f
C2612 VDD.t368 VSS 0.00992f
C2613 VDD.n426 VSS 0.00669f
C2614 VDD.t10 VSS 0.141f
C2615 VDD.n427 VSS 0.00547f
C2616 VDD.t332 VSS 0.00993f
C2617 VDD.n428 VSS 0.0066f
C2618 VDD.t96 VSS 0.141f
C2619 VDD.n429 VSS 0.00547f
C2620 VDD.t383 VSS 0.00993f
C2621 VDD.n430 VSS 0.0066f
C2622 VDD.t412 VSS 0.141f
C2623 VDD.n431 VSS 0.00547f
C2624 VDD.t358 VSS 0.00993f
C2625 VDD.n432 VSS 0.00668f
C2626 VDD.t295 VSS 0.115f
C2627 VDD.n433 VSS 0.00578f
C2628 VDD.n434 VSS 0.0274f
C2629 VDD.n435 VSS 0.0142f
C2630 VDD.t357 VSS 0.141f
C2631 VDD.n436 VSS 0.0142f
C2632 VDD.n437 VSS 0.0191f
C2633 VDD.n438 VSS 0.0246f
C2634 VDD.n439 VSS 0.0142f
C2635 VDD.t382 VSS 0.141f
C2636 VDD.n440 VSS 0.0142f
C2637 VDD.n441 VSS 0.0191f
C2638 VDD.n442 VSS 0.0246f
C2639 VDD.n443 VSS 0.0142f
C2640 VDD.t331 VSS 0.141f
C2641 VDD.n444 VSS 0.0142f
C2642 VDD.n445 VSS 0.0191f
C2643 VDD.n446 VSS 0.0245f
C2644 VDD.n447 VSS 0.0142f
C2645 VDD.t367 VSS 0.0672f
C2646 VDD.n448 VSS 0.0142f
C2647 VDD.n449 VSS 0.0277f
C2648 VDD.t33 VSS 0.091f
C2649 VDD.n450 VSS 0.0497f
C2650 VDD.t219 VSS 0.00547f
C2651 VDD.n451 VSS 0.0336f
C2652 VDD.t218 VSS 0.091f
C2653 VDD.n452 VSS 0.0458f
C2654 VDD.n453 VSS 0.0246f
C2655 VDD.n454 VSS 0.039f
C2656 VDD.n455 VSS 0.037f
C2657 VDD.n456 VSS 0.0302f
C2658 VDD.n457 VSS 0.0288f
C2659 VDD.t275 VSS 0.00547f
C2660 VDD.n458 VSS 0.0288f
C2661 VDD.n459 VSS 0.0298f
C2662 VDD.t274 VSS 0.131f
C2663 VDD.t290 VSS 0.125f
C2664 VDD.t439 VSS 0.104f
C2665 VDD.n460 VSS 0.0314f
C2666 VDD.n461 VSS 0.0443f
C2667 VDD.n462 VSS 0.00549f
C2668 VDD.t407 VSS 0.0715f
C2669 VDD.n463 VSS 0.0341f
C2670 VDD.t234 VSS 0.0055f
C2671 VDD.n464 VSS 0.00549f
C2672 VDD.t233 VSS 0.0662f
C2673 VDD.t205 VSS 0.0725f
C2674 VDD.n465 VSS 0.0341f
C2675 VDD.t119 VSS 0.0055f
C2676 VDD.t155 VSS 0.00226f
C2677 VDD.n466 VSS 0.00226f
C2678 VDD.n467 VSS 0.00493f
C2679 VDD.t118 VSS 0.0662f
C2680 VDD.t154 VSS 0.0809f
C2681 VDD.t222 VSS 0.0376f
C2682 VDD.n468 VSS 0.0341f
C2683 VDD.t180 VSS 0.0055f
C2684 VDD.t411 VSS 0.00226f
C2685 VDD.n469 VSS 0.00226f
C2686 VDD.n470 VSS 0.00493f
C2687 VDD.t179 VSS 0.0662f
C2688 VDD.t410 VSS 0.0809f
C2689 VDD.t79 VSS 0.0376f
C2690 VDD.t69 VSS 0.066f
C2691 VDD.n471 VSS 0.0341f
C2692 VDD.t70 VSS 0.0055f
C2693 VDD.t45 VSS 0.00471f
C2694 VDD.t485 VSS 0.00357f
C2695 VDD.n472 VSS 0.00924f
C2696 VDD.n473 VSS 0.00852f
C2697 VDD.t68 VSS 0.00471f
C2698 VDD.t479 VSS 0.00357f
C2699 VDD.n474 VSS 0.00926f
C2700 VDD.n475 VSS 0.00691f
C2701 VDD.n476 VSS 0.0441f
C2702 VDD.n477 VSS 0.0256f
C2703 VDD.n478 VSS 0.017f
C2704 VDD.n479 VSS 0.0313f
C2705 VDD.n480 VSS 0.0321f
C2706 VDD.n481 VSS 0.017f
C2707 VDD.n482 VSS 0.0313f
C2708 VDD.n483 VSS 0.032f
C2709 VDD.n484 VSS 0.019f
C2710 VDD.n485 VSS 0.0272f
C2711 VDD.n486 VSS 0.0253f
C2712 VDD.n487 VSS 0.019f
C2713 VDD.n488 VSS 0.0201f
C2714 VDD.n489 VSS 0.0449f
C2715 VDD.n490 VSS 0.0412f
C2716 VDD.n491 VSS 0.0529f
C2717 VDD.n492 VSS 0.0151f
C2718 VDD.n493 VSS 0.0227f
C2719 VDD.n494 VSS 0.0355f
C2720 VDD.n495 VSS 0.0309f
C2721 VDD.n496 VSS 0.0364f
C2722 VDD.n497 VSS 0.0225f
C2723 VDD.n498 VSS 0.0342f
C2724 VDD.n499 VSS 0.03f
C2725 VDD.n500 VSS 0.031f
C2726 VDD.t406 VSS 0.0131f
C2727 VDD.t284 VSS 0.00547f
C2728 VDD.n501 VSS 0.0294f
C2729 VDD.t283 VSS 0.0487f
C2730 VDD.n502 VSS 0.0577f
C2731 VDD.t282 VSS 0.0518f
C2732 VDD.t405 VSS 0.084f
C2733 VDD.n503 VSS 0.0404f
C2734 VDD.n504 VSS 0.0292f
C2735 VDD.n505 VSS 0.0244f
C2736 VDD.n506 VSS 0.0956f
C2737 VDD.n507 VSS 0.139f
C2738 CLK_div_31_mag_0.Q0.n0 VSS 0.109f
C2739 CLK_div_31_mag_0.Q0.n1 VSS 0.0183f
C2740 CLK_div_31_mag_0.Q0.t0 VSS 0.0256f
C2741 CLK_div_31_mag_0.Q0.t2 VSS 0.0211f
C2742 CLK_div_31_mag_0.Q0.n2 VSS 0.0211f
C2743 CLK_div_31_mag_0.Q0.n3 VSS 0.0508f
C2744 CLK_div_31_mag_0.Q0.n4 VSS 0.158f
C2745 CLK_div_31_mag_0.Q0.n5 VSS 0.0296f
C2746 CLK_div_31_mag_0.Q0.t12 VSS 0.0388f
C2747 CLK_div_31_mag_0.Q0.t14 VSS 0.0101f
C2748 CLK_div_31_mag_0.Q0.n6 VSS 0.0644f
C2749 CLK_div_31_mag_0.Q0.n7 VSS 0.00386f
C2750 CLK_div_31_mag_0.Q0.n8 VSS 0.0154f
C2751 CLK_div_31_mag_0.Q0.t11 VSS 0.0471f
C2752 CLK_div_31_mag_0.Q0.t9 VSS 0.031f
C2753 CLK_div_31_mag_0.Q0.n9 VSS 0.0832f
C2754 CLK_div_31_mag_0.Q0.n10 VSS 0.0109f
C2755 CLK_div_31_mag_0.Q0.n11 VSS 0.00782f
C2756 CLK_div_31_mag_0.Q0.n12 VSS 0.0039f
C2757 CLK_div_31_mag_0.Q0.n13 VSS 0.156f
C2758 CLK_div_31_mag_0.Q0.t8 VSS 0.0471f
C2759 CLK_div_31_mag_0.Q0.t5 VSS 0.031f
C2760 CLK_div_31_mag_0.Q0.n14 VSS 0.0832f
C2761 CLK_div_31_mag_0.Q0.n15 VSS 0.0109f
C2762 CLK_div_31_mag_0.Q0.n16 VSS 0.00782f
C2763 CLK_div_31_mag_0.Q0.n17 VSS 0.154f
C2764 CLK_div_31_mag_0.Q0.n18 VSS 0.0951f
C2765 CLK_div_31_mag_0.Q0.n19 VSS 0.1f
C2766 CLK_div_31_mag_0.Q0.t4 VSS 0.0471f
C2767 CLK_div_31_mag_0.Q0.t3 VSS 0.031f
C2768 CLK_div_31_mag_0.Q0.n20 VSS 0.0836f
C2769 CLK_div_31_mag_0.Q0.n21 VSS 0.0283f
C2770 CLK_div_31_mag_0.Q0.t6 VSS 0.0441f
C2771 CLK_div_31_mag_0.Q0.t16 VSS 0.0241f
C2772 CLK_div_31_mag_0.Q0.n22 VSS 0.0838f
C2773 CLK_div_31_mag_0.Q0.t10 VSS 0.0241f
C2774 CLK_div_31_mag_0.Q0.t7 VSS 0.0441f
C2775 CLK_div_31_mag_0.Q0.n23 VSS 0.0838f
C2776 CLK_div_31_mag_0.Q0.n24 VSS 0.479f
C2777 CLK_div_31_mag_0.Q0.n25 VSS 0.725f
C2778 CLK_div_31_mag_0.Q0.t15 VSS 0.0338f
C2779 CLK_div_31_mag_0.Q0.t13 VSS 0.027f
C2780 CLK_div_31_mag_0.Q0.n26 VSS 0.0785f
C2781 CLK_div_31_mag_0.Q0.n27 VSS 0.0487f
C2782 CLK_div_31_mag_0.Q0.n28 VSS 0.5f
C2783 CLK_div_31_mag_0.Q0.n29 VSS 0.02f
.ends

