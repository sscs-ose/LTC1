magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -9345 -2095 9345 2095
<< psubdiff >>
rect -7345 70 7345 95
rect -7345 -70 -7308 70
rect 7308 -70 7345 70
rect -7345 -95 7345 -70
<< psubdiffcont >>
rect -7308 -70 7308 70
<< metal1 >>
rect -7334 70 7334 84
rect -7334 -70 -7308 70
rect 7308 -70 7334 70
rect -7334 -84 7334 -70
<< end >>
