magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1071 1045 1071
<< metal1 >>
rect -45 65 45 71
rect -45 -65 -39 65
rect 39 -65 45 65
rect -45 -71 45 -65
<< via1 >>
rect -39 -65 39 65
<< metal2 >>
rect -45 65 45 71
rect -45 -65 -39 65
rect 39 -65 45 65
rect -45 -71 45 -65
<< end >>
