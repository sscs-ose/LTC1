magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2083 -2083 4795 4575
<< isosubstrate >>
rect 1197 -83 2795 2575
<< nwell >>
rect -83 1281 857 2439
rect 1197 1281 2795 2575
<< polysilicon >>
rect 316 698 456 1442
rect 1561 1202 1701 1578
rect 1805 1202 1945 1578
rect 1561 991 1945 1202
rect 1561 698 1701 991
rect 1805 698 1945 991
rect 2049 1202 2189 1578
rect 2293 1202 2433 1578
rect 2049 991 2433 1202
rect 2049 698 2189 991
rect 2293 698 2433 991
<< metal1 >>
rect 79 2413 165 2481
rect 226 1486 302 2468
rect 609 2413 695 2481
rect 1359 2413 1445 2481
rect 470 1186 546 2086
rect 1471 1622 1547 2451
rect 1715 1186 1791 2222
rect 1959 1622 2035 2451
rect 470 1008 1655 1186
rect 1715 1008 2143 1186
rect 79 11 165 79
rect 226 42 302 654
rect 470 354 546 1008
rect 609 11 695 79
rect 1359 11 1445 79
rect 1471 39 1547 654
rect 1715 354 1791 1008
rect 1959 39 2035 654
rect 2203 354 2279 2222
rect 2447 1622 2523 2451
rect 2547 2413 2633 2481
rect 2447 39 2523 654
rect 2547 11 2633 79
use M1_NWELL_CDNS_40661953145273  M1_NWELL_CDNS_40661953145273_0
timestamp 1713338890
transform 1 0 387 0 1 2447
box -316 -128 316 128
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_0
timestamp 1713338890
transform 1 0 1325 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_1
timestamp 1713338890
transform 1 0 729 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_2
timestamp 1713338890
transform 1 0 45 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_3
timestamp 1713338890
transform 1 0 2667 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145322  M1_NWELL_CDNS_40661953145322_0
timestamp 1713338890
transform 1 0 1996 0 1 2447
box -645 -128 645 128
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform 1 0 376 0 1 1097
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform 1 0 1621 0 1 1097
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_2
timestamp 1713338890
transform 1 0 2109 0 1 1097
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 1 0 45 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 1 0 2667 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165611  M1_PSUB_CDNS_69033583165611_0
timestamp 1713338890
transform 1 0 729 0 -1 468
box -45 -468 45 468
use M1_PSUB_CDNS_69033583165611  M1_PSUB_CDNS_69033583165611_1
timestamp 1713338890
transform 1 0 1325 0 -1 468
box -45 -468 45 468
use M1_PSUB_CDNS_69033583165620  M1_PSUB_CDNS_69033583165620_0
timestamp 1713338890
transform 1 0 1996 0 -1 45
box -562 -45 562 45
use M1_PSUB_CDNS_69033583165621  M1_PSUB_CDNS_69033583165621_0
timestamp 1713338890
transform 1 0 387 0 -1 45
box -233 -45 233 45
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_0
timestamp 1713338890
transform 1 0 316 0 1 354
box -88 -44 228 344
use nmos_6p0_CDNS_4066195314531  nmos_6p0_CDNS_4066195314531_0
timestamp 1713338890
transform 1 0 1561 0 1 354
box -88 -44 472 344
use nmos_6p0_CDNS_4066195314531  nmos_6p0_CDNS_4066195314531_1
timestamp 1713338890
transform 1 0 2049 0 1 354
box -88 -44 472 344
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1713338890
transform 1 0 316 0 1 1486
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314529  pmos_6p0_CDNS_4066195314529_0
timestamp 1713338890
transform 1 0 1561 0 1 1622
box -208 -120 592 720
use pmos_6p0_CDNS_4066195314529  pmos_6p0_CDNS_4066195314529_1
timestamp 1713338890
transform 1 0 2049 0 1 1622
box -208 -120 592 720
<< labels >>
rlabel metal1 s 2242 1098 2242 1098 4 ZB
port 1 nsew
rlabel metal1 s 29 2452 29 2452 4 VDD
port 2 nsew
rlabel metal1 s 376 1098 376 1098 4 A
port 3 nsew
rlabel metal1 s 2348 2452 2348 2452 4 DVDD
port 4 nsew
rlabel metal1 s 2339 45 2339 45 4 DVSS
port 5 nsew
rlabel metal1 s 263 45 263 45 4 VSS
port 6 nsew
rlabel metal1 s 1987 1098 1987 1098 4 Z
port 7 nsew
<< end >>
