magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1319 -2540 1319 2540
<< metal4 >>
rect -316 1532 316 1537
rect -316 1504 -311 1532
rect -283 1504 -245 1532
rect -217 1504 -179 1532
rect -151 1504 -113 1532
rect -85 1504 -47 1532
rect -19 1504 19 1532
rect 47 1504 85 1532
rect 113 1504 151 1532
rect 179 1504 217 1532
rect 245 1504 283 1532
rect 311 1504 316 1532
rect -316 1466 316 1504
rect -316 1438 -311 1466
rect -283 1438 -245 1466
rect -217 1438 -179 1466
rect -151 1438 -113 1466
rect -85 1438 -47 1466
rect -19 1438 19 1466
rect 47 1438 85 1466
rect 113 1438 151 1466
rect 179 1438 217 1466
rect 245 1438 283 1466
rect 311 1438 316 1466
rect -316 1400 316 1438
rect -316 1372 -311 1400
rect -283 1372 -245 1400
rect -217 1372 -179 1400
rect -151 1372 -113 1400
rect -85 1372 -47 1400
rect -19 1372 19 1400
rect 47 1372 85 1400
rect 113 1372 151 1400
rect 179 1372 217 1400
rect 245 1372 283 1400
rect 311 1372 316 1400
rect -316 1334 316 1372
rect -316 1306 -311 1334
rect -283 1306 -245 1334
rect -217 1306 -179 1334
rect -151 1306 -113 1334
rect -85 1306 -47 1334
rect -19 1306 19 1334
rect 47 1306 85 1334
rect 113 1306 151 1334
rect 179 1306 217 1334
rect 245 1306 283 1334
rect 311 1306 316 1334
rect -316 1268 316 1306
rect -316 1240 -311 1268
rect -283 1240 -245 1268
rect -217 1240 -179 1268
rect -151 1240 -113 1268
rect -85 1240 -47 1268
rect -19 1240 19 1268
rect 47 1240 85 1268
rect 113 1240 151 1268
rect 179 1240 217 1268
rect 245 1240 283 1268
rect 311 1240 316 1268
rect -316 1202 316 1240
rect -316 1174 -311 1202
rect -283 1174 -245 1202
rect -217 1174 -179 1202
rect -151 1174 -113 1202
rect -85 1174 -47 1202
rect -19 1174 19 1202
rect 47 1174 85 1202
rect 113 1174 151 1202
rect 179 1174 217 1202
rect 245 1174 283 1202
rect 311 1174 316 1202
rect -316 1136 316 1174
rect -316 1108 -311 1136
rect -283 1108 -245 1136
rect -217 1108 -179 1136
rect -151 1108 -113 1136
rect -85 1108 -47 1136
rect -19 1108 19 1136
rect 47 1108 85 1136
rect 113 1108 151 1136
rect 179 1108 217 1136
rect 245 1108 283 1136
rect 311 1108 316 1136
rect -316 1070 316 1108
rect -316 1042 -311 1070
rect -283 1042 -245 1070
rect -217 1042 -179 1070
rect -151 1042 -113 1070
rect -85 1042 -47 1070
rect -19 1042 19 1070
rect 47 1042 85 1070
rect 113 1042 151 1070
rect 179 1042 217 1070
rect 245 1042 283 1070
rect 311 1042 316 1070
rect -316 1004 316 1042
rect -316 976 -311 1004
rect -283 976 -245 1004
rect -217 976 -179 1004
rect -151 976 -113 1004
rect -85 976 -47 1004
rect -19 976 19 1004
rect 47 976 85 1004
rect 113 976 151 1004
rect 179 976 217 1004
rect 245 976 283 1004
rect 311 976 316 1004
rect -316 938 316 976
rect -316 910 -311 938
rect -283 910 -245 938
rect -217 910 -179 938
rect -151 910 -113 938
rect -85 910 -47 938
rect -19 910 19 938
rect 47 910 85 938
rect 113 910 151 938
rect 179 910 217 938
rect 245 910 283 938
rect 311 910 316 938
rect -316 872 316 910
rect -316 844 -311 872
rect -283 844 -245 872
rect -217 844 -179 872
rect -151 844 -113 872
rect -85 844 -47 872
rect -19 844 19 872
rect 47 844 85 872
rect 113 844 151 872
rect 179 844 217 872
rect 245 844 283 872
rect 311 844 316 872
rect -316 806 316 844
rect -316 778 -311 806
rect -283 778 -245 806
rect -217 778 -179 806
rect -151 778 -113 806
rect -85 778 -47 806
rect -19 778 19 806
rect 47 778 85 806
rect 113 778 151 806
rect 179 778 217 806
rect 245 778 283 806
rect 311 778 316 806
rect -316 740 316 778
rect -316 712 -311 740
rect -283 712 -245 740
rect -217 712 -179 740
rect -151 712 -113 740
rect -85 712 -47 740
rect -19 712 19 740
rect 47 712 85 740
rect 113 712 151 740
rect 179 712 217 740
rect 245 712 283 740
rect 311 712 316 740
rect -316 674 316 712
rect -316 646 -311 674
rect -283 646 -245 674
rect -217 646 -179 674
rect -151 646 -113 674
rect -85 646 -47 674
rect -19 646 19 674
rect 47 646 85 674
rect 113 646 151 674
rect 179 646 217 674
rect 245 646 283 674
rect 311 646 316 674
rect -316 608 316 646
rect -316 580 -311 608
rect -283 580 -245 608
rect -217 580 -179 608
rect -151 580 -113 608
rect -85 580 -47 608
rect -19 580 19 608
rect 47 580 85 608
rect 113 580 151 608
rect 179 580 217 608
rect 245 580 283 608
rect 311 580 316 608
rect -316 542 316 580
rect -316 514 -311 542
rect -283 514 -245 542
rect -217 514 -179 542
rect -151 514 -113 542
rect -85 514 -47 542
rect -19 514 19 542
rect 47 514 85 542
rect 113 514 151 542
rect 179 514 217 542
rect 245 514 283 542
rect 311 514 316 542
rect -316 476 316 514
rect -316 448 -311 476
rect -283 448 -245 476
rect -217 448 -179 476
rect -151 448 -113 476
rect -85 448 -47 476
rect -19 448 19 476
rect 47 448 85 476
rect 113 448 151 476
rect 179 448 217 476
rect 245 448 283 476
rect 311 448 316 476
rect -316 410 316 448
rect -316 382 -311 410
rect -283 382 -245 410
rect -217 382 -179 410
rect -151 382 -113 410
rect -85 382 -47 410
rect -19 382 19 410
rect 47 382 85 410
rect 113 382 151 410
rect 179 382 217 410
rect 245 382 283 410
rect 311 382 316 410
rect -316 344 316 382
rect -316 316 -311 344
rect -283 316 -245 344
rect -217 316 -179 344
rect -151 316 -113 344
rect -85 316 -47 344
rect -19 316 19 344
rect 47 316 85 344
rect 113 316 151 344
rect 179 316 217 344
rect 245 316 283 344
rect 311 316 316 344
rect -316 278 316 316
rect -316 250 -311 278
rect -283 250 -245 278
rect -217 250 -179 278
rect -151 250 -113 278
rect -85 250 -47 278
rect -19 250 19 278
rect 47 250 85 278
rect 113 250 151 278
rect 179 250 217 278
rect 245 250 283 278
rect 311 250 316 278
rect -316 212 316 250
rect -316 184 -311 212
rect -283 184 -245 212
rect -217 184 -179 212
rect -151 184 -113 212
rect -85 184 -47 212
rect -19 184 19 212
rect 47 184 85 212
rect 113 184 151 212
rect 179 184 217 212
rect 245 184 283 212
rect 311 184 316 212
rect -316 146 316 184
rect -316 118 -311 146
rect -283 118 -245 146
rect -217 118 -179 146
rect -151 118 -113 146
rect -85 118 -47 146
rect -19 118 19 146
rect 47 118 85 146
rect 113 118 151 146
rect 179 118 217 146
rect 245 118 283 146
rect 311 118 316 146
rect -316 80 316 118
rect -316 52 -311 80
rect -283 52 -245 80
rect -217 52 -179 80
rect -151 52 -113 80
rect -85 52 -47 80
rect -19 52 19 80
rect 47 52 85 80
rect 113 52 151 80
rect 179 52 217 80
rect 245 52 283 80
rect 311 52 316 80
rect -316 14 316 52
rect -316 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 19 14
rect 47 -14 85 14
rect 113 -14 151 14
rect 179 -14 217 14
rect 245 -14 283 14
rect 311 -14 316 14
rect -316 -52 316 -14
rect -316 -80 -311 -52
rect -283 -80 -245 -52
rect -217 -80 -179 -52
rect -151 -80 -113 -52
rect -85 -80 -47 -52
rect -19 -80 19 -52
rect 47 -80 85 -52
rect 113 -80 151 -52
rect 179 -80 217 -52
rect 245 -80 283 -52
rect 311 -80 316 -52
rect -316 -118 316 -80
rect -316 -146 -311 -118
rect -283 -146 -245 -118
rect -217 -146 -179 -118
rect -151 -146 -113 -118
rect -85 -146 -47 -118
rect -19 -146 19 -118
rect 47 -146 85 -118
rect 113 -146 151 -118
rect 179 -146 217 -118
rect 245 -146 283 -118
rect 311 -146 316 -118
rect -316 -184 316 -146
rect -316 -212 -311 -184
rect -283 -212 -245 -184
rect -217 -212 -179 -184
rect -151 -212 -113 -184
rect -85 -212 -47 -184
rect -19 -212 19 -184
rect 47 -212 85 -184
rect 113 -212 151 -184
rect 179 -212 217 -184
rect 245 -212 283 -184
rect 311 -212 316 -184
rect -316 -250 316 -212
rect -316 -278 -311 -250
rect -283 -278 -245 -250
rect -217 -278 -179 -250
rect -151 -278 -113 -250
rect -85 -278 -47 -250
rect -19 -278 19 -250
rect 47 -278 85 -250
rect 113 -278 151 -250
rect 179 -278 217 -250
rect 245 -278 283 -250
rect 311 -278 316 -250
rect -316 -316 316 -278
rect -316 -344 -311 -316
rect -283 -344 -245 -316
rect -217 -344 -179 -316
rect -151 -344 -113 -316
rect -85 -344 -47 -316
rect -19 -344 19 -316
rect 47 -344 85 -316
rect 113 -344 151 -316
rect 179 -344 217 -316
rect 245 -344 283 -316
rect 311 -344 316 -316
rect -316 -382 316 -344
rect -316 -410 -311 -382
rect -283 -410 -245 -382
rect -217 -410 -179 -382
rect -151 -410 -113 -382
rect -85 -410 -47 -382
rect -19 -410 19 -382
rect 47 -410 85 -382
rect 113 -410 151 -382
rect 179 -410 217 -382
rect 245 -410 283 -382
rect 311 -410 316 -382
rect -316 -448 316 -410
rect -316 -476 -311 -448
rect -283 -476 -245 -448
rect -217 -476 -179 -448
rect -151 -476 -113 -448
rect -85 -476 -47 -448
rect -19 -476 19 -448
rect 47 -476 85 -448
rect 113 -476 151 -448
rect 179 -476 217 -448
rect 245 -476 283 -448
rect 311 -476 316 -448
rect -316 -514 316 -476
rect -316 -542 -311 -514
rect -283 -542 -245 -514
rect -217 -542 -179 -514
rect -151 -542 -113 -514
rect -85 -542 -47 -514
rect -19 -542 19 -514
rect 47 -542 85 -514
rect 113 -542 151 -514
rect 179 -542 217 -514
rect 245 -542 283 -514
rect 311 -542 316 -514
rect -316 -580 316 -542
rect -316 -608 -311 -580
rect -283 -608 -245 -580
rect -217 -608 -179 -580
rect -151 -608 -113 -580
rect -85 -608 -47 -580
rect -19 -608 19 -580
rect 47 -608 85 -580
rect 113 -608 151 -580
rect 179 -608 217 -580
rect 245 -608 283 -580
rect 311 -608 316 -580
rect -316 -646 316 -608
rect -316 -674 -311 -646
rect -283 -674 -245 -646
rect -217 -674 -179 -646
rect -151 -674 -113 -646
rect -85 -674 -47 -646
rect -19 -674 19 -646
rect 47 -674 85 -646
rect 113 -674 151 -646
rect 179 -674 217 -646
rect 245 -674 283 -646
rect 311 -674 316 -646
rect -316 -712 316 -674
rect -316 -740 -311 -712
rect -283 -740 -245 -712
rect -217 -740 -179 -712
rect -151 -740 -113 -712
rect -85 -740 -47 -712
rect -19 -740 19 -712
rect 47 -740 85 -712
rect 113 -740 151 -712
rect 179 -740 217 -712
rect 245 -740 283 -712
rect 311 -740 316 -712
rect -316 -778 316 -740
rect -316 -806 -311 -778
rect -283 -806 -245 -778
rect -217 -806 -179 -778
rect -151 -806 -113 -778
rect -85 -806 -47 -778
rect -19 -806 19 -778
rect 47 -806 85 -778
rect 113 -806 151 -778
rect 179 -806 217 -778
rect 245 -806 283 -778
rect 311 -806 316 -778
rect -316 -844 316 -806
rect -316 -872 -311 -844
rect -283 -872 -245 -844
rect -217 -872 -179 -844
rect -151 -872 -113 -844
rect -85 -872 -47 -844
rect -19 -872 19 -844
rect 47 -872 85 -844
rect 113 -872 151 -844
rect 179 -872 217 -844
rect 245 -872 283 -844
rect 311 -872 316 -844
rect -316 -910 316 -872
rect -316 -938 -311 -910
rect -283 -938 -245 -910
rect -217 -938 -179 -910
rect -151 -938 -113 -910
rect -85 -938 -47 -910
rect -19 -938 19 -910
rect 47 -938 85 -910
rect 113 -938 151 -910
rect 179 -938 217 -910
rect 245 -938 283 -910
rect 311 -938 316 -910
rect -316 -976 316 -938
rect -316 -1004 -311 -976
rect -283 -1004 -245 -976
rect -217 -1004 -179 -976
rect -151 -1004 -113 -976
rect -85 -1004 -47 -976
rect -19 -1004 19 -976
rect 47 -1004 85 -976
rect 113 -1004 151 -976
rect 179 -1004 217 -976
rect 245 -1004 283 -976
rect 311 -1004 316 -976
rect -316 -1042 316 -1004
rect -316 -1070 -311 -1042
rect -283 -1070 -245 -1042
rect -217 -1070 -179 -1042
rect -151 -1070 -113 -1042
rect -85 -1070 -47 -1042
rect -19 -1070 19 -1042
rect 47 -1070 85 -1042
rect 113 -1070 151 -1042
rect 179 -1070 217 -1042
rect 245 -1070 283 -1042
rect 311 -1070 316 -1042
rect -316 -1108 316 -1070
rect -316 -1136 -311 -1108
rect -283 -1136 -245 -1108
rect -217 -1136 -179 -1108
rect -151 -1136 -113 -1108
rect -85 -1136 -47 -1108
rect -19 -1136 19 -1108
rect 47 -1136 85 -1108
rect 113 -1136 151 -1108
rect 179 -1136 217 -1108
rect 245 -1136 283 -1108
rect 311 -1136 316 -1108
rect -316 -1174 316 -1136
rect -316 -1202 -311 -1174
rect -283 -1202 -245 -1174
rect -217 -1202 -179 -1174
rect -151 -1202 -113 -1174
rect -85 -1202 -47 -1174
rect -19 -1202 19 -1174
rect 47 -1202 85 -1174
rect 113 -1202 151 -1174
rect 179 -1202 217 -1174
rect 245 -1202 283 -1174
rect 311 -1202 316 -1174
rect -316 -1240 316 -1202
rect -316 -1268 -311 -1240
rect -283 -1268 -245 -1240
rect -217 -1268 -179 -1240
rect -151 -1268 -113 -1240
rect -85 -1268 -47 -1240
rect -19 -1268 19 -1240
rect 47 -1268 85 -1240
rect 113 -1268 151 -1240
rect 179 -1268 217 -1240
rect 245 -1268 283 -1240
rect 311 -1268 316 -1240
rect -316 -1306 316 -1268
rect -316 -1334 -311 -1306
rect -283 -1334 -245 -1306
rect -217 -1334 -179 -1306
rect -151 -1334 -113 -1306
rect -85 -1334 -47 -1306
rect -19 -1334 19 -1306
rect 47 -1334 85 -1306
rect 113 -1334 151 -1306
rect 179 -1334 217 -1306
rect 245 -1334 283 -1306
rect 311 -1334 316 -1306
rect -316 -1372 316 -1334
rect -316 -1400 -311 -1372
rect -283 -1400 -245 -1372
rect -217 -1400 -179 -1372
rect -151 -1400 -113 -1372
rect -85 -1400 -47 -1372
rect -19 -1400 19 -1372
rect 47 -1400 85 -1372
rect 113 -1400 151 -1372
rect 179 -1400 217 -1372
rect 245 -1400 283 -1372
rect 311 -1400 316 -1372
rect -316 -1438 316 -1400
rect -316 -1466 -311 -1438
rect -283 -1466 -245 -1438
rect -217 -1466 -179 -1438
rect -151 -1466 -113 -1438
rect -85 -1466 -47 -1438
rect -19 -1466 19 -1438
rect 47 -1466 85 -1438
rect 113 -1466 151 -1438
rect 179 -1466 217 -1438
rect 245 -1466 283 -1438
rect 311 -1466 316 -1438
rect -316 -1504 316 -1466
rect -316 -1532 -311 -1504
rect -283 -1532 -245 -1504
rect -217 -1532 -179 -1504
rect -151 -1532 -113 -1504
rect -85 -1532 -47 -1504
rect -19 -1532 19 -1504
rect 47 -1532 85 -1504
rect 113 -1532 151 -1504
rect 179 -1532 217 -1504
rect 245 -1532 283 -1504
rect 311 -1532 316 -1504
rect -316 -1537 316 -1532
<< via4 >>
rect -311 1504 -283 1532
rect -245 1504 -217 1532
rect -179 1504 -151 1532
rect -113 1504 -85 1532
rect -47 1504 -19 1532
rect 19 1504 47 1532
rect 85 1504 113 1532
rect 151 1504 179 1532
rect 217 1504 245 1532
rect 283 1504 311 1532
rect -311 1438 -283 1466
rect -245 1438 -217 1466
rect -179 1438 -151 1466
rect -113 1438 -85 1466
rect -47 1438 -19 1466
rect 19 1438 47 1466
rect 85 1438 113 1466
rect 151 1438 179 1466
rect 217 1438 245 1466
rect 283 1438 311 1466
rect -311 1372 -283 1400
rect -245 1372 -217 1400
rect -179 1372 -151 1400
rect -113 1372 -85 1400
rect -47 1372 -19 1400
rect 19 1372 47 1400
rect 85 1372 113 1400
rect 151 1372 179 1400
rect 217 1372 245 1400
rect 283 1372 311 1400
rect -311 1306 -283 1334
rect -245 1306 -217 1334
rect -179 1306 -151 1334
rect -113 1306 -85 1334
rect -47 1306 -19 1334
rect 19 1306 47 1334
rect 85 1306 113 1334
rect 151 1306 179 1334
rect 217 1306 245 1334
rect 283 1306 311 1334
rect -311 1240 -283 1268
rect -245 1240 -217 1268
rect -179 1240 -151 1268
rect -113 1240 -85 1268
rect -47 1240 -19 1268
rect 19 1240 47 1268
rect 85 1240 113 1268
rect 151 1240 179 1268
rect 217 1240 245 1268
rect 283 1240 311 1268
rect -311 1174 -283 1202
rect -245 1174 -217 1202
rect -179 1174 -151 1202
rect -113 1174 -85 1202
rect -47 1174 -19 1202
rect 19 1174 47 1202
rect 85 1174 113 1202
rect 151 1174 179 1202
rect 217 1174 245 1202
rect 283 1174 311 1202
rect -311 1108 -283 1136
rect -245 1108 -217 1136
rect -179 1108 -151 1136
rect -113 1108 -85 1136
rect -47 1108 -19 1136
rect 19 1108 47 1136
rect 85 1108 113 1136
rect 151 1108 179 1136
rect 217 1108 245 1136
rect 283 1108 311 1136
rect -311 1042 -283 1070
rect -245 1042 -217 1070
rect -179 1042 -151 1070
rect -113 1042 -85 1070
rect -47 1042 -19 1070
rect 19 1042 47 1070
rect 85 1042 113 1070
rect 151 1042 179 1070
rect 217 1042 245 1070
rect 283 1042 311 1070
rect -311 976 -283 1004
rect -245 976 -217 1004
rect -179 976 -151 1004
rect -113 976 -85 1004
rect -47 976 -19 1004
rect 19 976 47 1004
rect 85 976 113 1004
rect 151 976 179 1004
rect 217 976 245 1004
rect 283 976 311 1004
rect -311 910 -283 938
rect -245 910 -217 938
rect -179 910 -151 938
rect -113 910 -85 938
rect -47 910 -19 938
rect 19 910 47 938
rect 85 910 113 938
rect 151 910 179 938
rect 217 910 245 938
rect 283 910 311 938
rect -311 844 -283 872
rect -245 844 -217 872
rect -179 844 -151 872
rect -113 844 -85 872
rect -47 844 -19 872
rect 19 844 47 872
rect 85 844 113 872
rect 151 844 179 872
rect 217 844 245 872
rect 283 844 311 872
rect -311 778 -283 806
rect -245 778 -217 806
rect -179 778 -151 806
rect -113 778 -85 806
rect -47 778 -19 806
rect 19 778 47 806
rect 85 778 113 806
rect 151 778 179 806
rect 217 778 245 806
rect 283 778 311 806
rect -311 712 -283 740
rect -245 712 -217 740
rect -179 712 -151 740
rect -113 712 -85 740
rect -47 712 -19 740
rect 19 712 47 740
rect 85 712 113 740
rect 151 712 179 740
rect 217 712 245 740
rect 283 712 311 740
rect -311 646 -283 674
rect -245 646 -217 674
rect -179 646 -151 674
rect -113 646 -85 674
rect -47 646 -19 674
rect 19 646 47 674
rect 85 646 113 674
rect 151 646 179 674
rect 217 646 245 674
rect 283 646 311 674
rect -311 580 -283 608
rect -245 580 -217 608
rect -179 580 -151 608
rect -113 580 -85 608
rect -47 580 -19 608
rect 19 580 47 608
rect 85 580 113 608
rect 151 580 179 608
rect 217 580 245 608
rect 283 580 311 608
rect -311 514 -283 542
rect -245 514 -217 542
rect -179 514 -151 542
rect -113 514 -85 542
rect -47 514 -19 542
rect 19 514 47 542
rect 85 514 113 542
rect 151 514 179 542
rect 217 514 245 542
rect 283 514 311 542
rect -311 448 -283 476
rect -245 448 -217 476
rect -179 448 -151 476
rect -113 448 -85 476
rect -47 448 -19 476
rect 19 448 47 476
rect 85 448 113 476
rect 151 448 179 476
rect 217 448 245 476
rect 283 448 311 476
rect -311 382 -283 410
rect -245 382 -217 410
rect -179 382 -151 410
rect -113 382 -85 410
rect -47 382 -19 410
rect 19 382 47 410
rect 85 382 113 410
rect 151 382 179 410
rect 217 382 245 410
rect 283 382 311 410
rect -311 316 -283 344
rect -245 316 -217 344
rect -179 316 -151 344
rect -113 316 -85 344
rect -47 316 -19 344
rect 19 316 47 344
rect 85 316 113 344
rect 151 316 179 344
rect 217 316 245 344
rect 283 316 311 344
rect -311 250 -283 278
rect -245 250 -217 278
rect -179 250 -151 278
rect -113 250 -85 278
rect -47 250 -19 278
rect 19 250 47 278
rect 85 250 113 278
rect 151 250 179 278
rect 217 250 245 278
rect 283 250 311 278
rect -311 184 -283 212
rect -245 184 -217 212
rect -179 184 -151 212
rect -113 184 -85 212
rect -47 184 -19 212
rect 19 184 47 212
rect 85 184 113 212
rect 151 184 179 212
rect 217 184 245 212
rect 283 184 311 212
rect -311 118 -283 146
rect -245 118 -217 146
rect -179 118 -151 146
rect -113 118 -85 146
rect -47 118 -19 146
rect 19 118 47 146
rect 85 118 113 146
rect 151 118 179 146
rect 217 118 245 146
rect 283 118 311 146
rect -311 52 -283 80
rect -245 52 -217 80
rect -179 52 -151 80
rect -113 52 -85 80
rect -47 52 -19 80
rect 19 52 47 80
rect 85 52 113 80
rect 151 52 179 80
rect 217 52 245 80
rect 283 52 311 80
rect -311 -14 -283 14
rect -245 -14 -217 14
rect -179 -14 -151 14
rect -113 -14 -85 14
rect -47 -14 -19 14
rect 19 -14 47 14
rect 85 -14 113 14
rect 151 -14 179 14
rect 217 -14 245 14
rect 283 -14 311 14
rect -311 -80 -283 -52
rect -245 -80 -217 -52
rect -179 -80 -151 -52
rect -113 -80 -85 -52
rect -47 -80 -19 -52
rect 19 -80 47 -52
rect 85 -80 113 -52
rect 151 -80 179 -52
rect 217 -80 245 -52
rect 283 -80 311 -52
rect -311 -146 -283 -118
rect -245 -146 -217 -118
rect -179 -146 -151 -118
rect -113 -146 -85 -118
rect -47 -146 -19 -118
rect 19 -146 47 -118
rect 85 -146 113 -118
rect 151 -146 179 -118
rect 217 -146 245 -118
rect 283 -146 311 -118
rect -311 -212 -283 -184
rect -245 -212 -217 -184
rect -179 -212 -151 -184
rect -113 -212 -85 -184
rect -47 -212 -19 -184
rect 19 -212 47 -184
rect 85 -212 113 -184
rect 151 -212 179 -184
rect 217 -212 245 -184
rect 283 -212 311 -184
rect -311 -278 -283 -250
rect -245 -278 -217 -250
rect -179 -278 -151 -250
rect -113 -278 -85 -250
rect -47 -278 -19 -250
rect 19 -278 47 -250
rect 85 -278 113 -250
rect 151 -278 179 -250
rect 217 -278 245 -250
rect 283 -278 311 -250
rect -311 -344 -283 -316
rect -245 -344 -217 -316
rect -179 -344 -151 -316
rect -113 -344 -85 -316
rect -47 -344 -19 -316
rect 19 -344 47 -316
rect 85 -344 113 -316
rect 151 -344 179 -316
rect 217 -344 245 -316
rect 283 -344 311 -316
rect -311 -410 -283 -382
rect -245 -410 -217 -382
rect -179 -410 -151 -382
rect -113 -410 -85 -382
rect -47 -410 -19 -382
rect 19 -410 47 -382
rect 85 -410 113 -382
rect 151 -410 179 -382
rect 217 -410 245 -382
rect 283 -410 311 -382
rect -311 -476 -283 -448
rect -245 -476 -217 -448
rect -179 -476 -151 -448
rect -113 -476 -85 -448
rect -47 -476 -19 -448
rect 19 -476 47 -448
rect 85 -476 113 -448
rect 151 -476 179 -448
rect 217 -476 245 -448
rect 283 -476 311 -448
rect -311 -542 -283 -514
rect -245 -542 -217 -514
rect -179 -542 -151 -514
rect -113 -542 -85 -514
rect -47 -542 -19 -514
rect 19 -542 47 -514
rect 85 -542 113 -514
rect 151 -542 179 -514
rect 217 -542 245 -514
rect 283 -542 311 -514
rect -311 -608 -283 -580
rect -245 -608 -217 -580
rect -179 -608 -151 -580
rect -113 -608 -85 -580
rect -47 -608 -19 -580
rect 19 -608 47 -580
rect 85 -608 113 -580
rect 151 -608 179 -580
rect 217 -608 245 -580
rect 283 -608 311 -580
rect -311 -674 -283 -646
rect -245 -674 -217 -646
rect -179 -674 -151 -646
rect -113 -674 -85 -646
rect -47 -674 -19 -646
rect 19 -674 47 -646
rect 85 -674 113 -646
rect 151 -674 179 -646
rect 217 -674 245 -646
rect 283 -674 311 -646
rect -311 -740 -283 -712
rect -245 -740 -217 -712
rect -179 -740 -151 -712
rect -113 -740 -85 -712
rect -47 -740 -19 -712
rect 19 -740 47 -712
rect 85 -740 113 -712
rect 151 -740 179 -712
rect 217 -740 245 -712
rect 283 -740 311 -712
rect -311 -806 -283 -778
rect -245 -806 -217 -778
rect -179 -806 -151 -778
rect -113 -806 -85 -778
rect -47 -806 -19 -778
rect 19 -806 47 -778
rect 85 -806 113 -778
rect 151 -806 179 -778
rect 217 -806 245 -778
rect 283 -806 311 -778
rect -311 -872 -283 -844
rect -245 -872 -217 -844
rect -179 -872 -151 -844
rect -113 -872 -85 -844
rect -47 -872 -19 -844
rect 19 -872 47 -844
rect 85 -872 113 -844
rect 151 -872 179 -844
rect 217 -872 245 -844
rect 283 -872 311 -844
rect -311 -938 -283 -910
rect -245 -938 -217 -910
rect -179 -938 -151 -910
rect -113 -938 -85 -910
rect -47 -938 -19 -910
rect 19 -938 47 -910
rect 85 -938 113 -910
rect 151 -938 179 -910
rect 217 -938 245 -910
rect 283 -938 311 -910
rect -311 -1004 -283 -976
rect -245 -1004 -217 -976
rect -179 -1004 -151 -976
rect -113 -1004 -85 -976
rect -47 -1004 -19 -976
rect 19 -1004 47 -976
rect 85 -1004 113 -976
rect 151 -1004 179 -976
rect 217 -1004 245 -976
rect 283 -1004 311 -976
rect -311 -1070 -283 -1042
rect -245 -1070 -217 -1042
rect -179 -1070 -151 -1042
rect -113 -1070 -85 -1042
rect -47 -1070 -19 -1042
rect 19 -1070 47 -1042
rect 85 -1070 113 -1042
rect 151 -1070 179 -1042
rect 217 -1070 245 -1042
rect 283 -1070 311 -1042
rect -311 -1136 -283 -1108
rect -245 -1136 -217 -1108
rect -179 -1136 -151 -1108
rect -113 -1136 -85 -1108
rect -47 -1136 -19 -1108
rect 19 -1136 47 -1108
rect 85 -1136 113 -1108
rect 151 -1136 179 -1108
rect 217 -1136 245 -1108
rect 283 -1136 311 -1108
rect -311 -1202 -283 -1174
rect -245 -1202 -217 -1174
rect -179 -1202 -151 -1174
rect -113 -1202 -85 -1174
rect -47 -1202 -19 -1174
rect 19 -1202 47 -1174
rect 85 -1202 113 -1174
rect 151 -1202 179 -1174
rect 217 -1202 245 -1174
rect 283 -1202 311 -1174
rect -311 -1268 -283 -1240
rect -245 -1268 -217 -1240
rect -179 -1268 -151 -1240
rect -113 -1268 -85 -1240
rect -47 -1268 -19 -1240
rect 19 -1268 47 -1240
rect 85 -1268 113 -1240
rect 151 -1268 179 -1240
rect 217 -1268 245 -1240
rect 283 -1268 311 -1240
rect -311 -1334 -283 -1306
rect -245 -1334 -217 -1306
rect -179 -1334 -151 -1306
rect -113 -1334 -85 -1306
rect -47 -1334 -19 -1306
rect 19 -1334 47 -1306
rect 85 -1334 113 -1306
rect 151 -1334 179 -1306
rect 217 -1334 245 -1306
rect 283 -1334 311 -1306
rect -311 -1400 -283 -1372
rect -245 -1400 -217 -1372
rect -179 -1400 -151 -1372
rect -113 -1400 -85 -1372
rect -47 -1400 -19 -1372
rect 19 -1400 47 -1372
rect 85 -1400 113 -1372
rect 151 -1400 179 -1372
rect 217 -1400 245 -1372
rect 283 -1400 311 -1372
rect -311 -1466 -283 -1438
rect -245 -1466 -217 -1438
rect -179 -1466 -151 -1438
rect -113 -1466 -85 -1438
rect -47 -1466 -19 -1438
rect 19 -1466 47 -1438
rect 85 -1466 113 -1438
rect 151 -1466 179 -1438
rect 217 -1466 245 -1438
rect 283 -1466 311 -1438
rect -311 -1532 -283 -1504
rect -245 -1532 -217 -1504
rect -179 -1532 -151 -1504
rect -113 -1532 -85 -1504
rect -47 -1532 -19 -1504
rect 19 -1532 47 -1504
rect 85 -1532 113 -1504
rect 151 -1532 179 -1504
rect 217 -1532 245 -1504
rect 283 -1532 311 -1504
<< metal5 >>
rect -319 1532 319 1540
rect -319 1504 -311 1532
rect -283 1504 -245 1532
rect -217 1504 -179 1532
rect -151 1504 -113 1532
rect -85 1504 -47 1532
rect -19 1504 19 1532
rect 47 1504 85 1532
rect 113 1504 151 1532
rect 179 1504 217 1532
rect 245 1504 283 1532
rect 311 1504 319 1532
rect -319 1466 319 1504
rect -319 1438 -311 1466
rect -283 1438 -245 1466
rect -217 1438 -179 1466
rect -151 1438 -113 1466
rect -85 1438 -47 1466
rect -19 1438 19 1466
rect 47 1438 85 1466
rect 113 1438 151 1466
rect 179 1438 217 1466
rect 245 1438 283 1466
rect 311 1438 319 1466
rect -319 1400 319 1438
rect -319 1372 -311 1400
rect -283 1372 -245 1400
rect -217 1372 -179 1400
rect -151 1372 -113 1400
rect -85 1372 -47 1400
rect -19 1372 19 1400
rect 47 1372 85 1400
rect 113 1372 151 1400
rect 179 1372 217 1400
rect 245 1372 283 1400
rect 311 1372 319 1400
rect -319 1334 319 1372
rect -319 1306 -311 1334
rect -283 1306 -245 1334
rect -217 1306 -179 1334
rect -151 1306 -113 1334
rect -85 1306 -47 1334
rect -19 1306 19 1334
rect 47 1306 85 1334
rect 113 1306 151 1334
rect 179 1306 217 1334
rect 245 1306 283 1334
rect 311 1306 319 1334
rect -319 1268 319 1306
rect -319 1240 -311 1268
rect -283 1240 -245 1268
rect -217 1240 -179 1268
rect -151 1240 -113 1268
rect -85 1240 -47 1268
rect -19 1240 19 1268
rect 47 1240 85 1268
rect 113 1240 151 1268
rect 179 1240 217 1268
rect 245 1240 283 1268
rect 311 1240 319 1268
rect -319 1202 319 1240
rect -319 1174 -311 1202
rect -283 1174 -245 1202
rect -217 1174 -179 1202
rect -151 1174 -113 1202
rect -85 1174 -47 1202
rect -19 1174 19 1202
rect 47 1174 85 1202
rect 113 1174 151 1202
rect 179 1174 217 1202
rect 245 1174 283 1202
rect 311 1174 319 1202
rect -319 1136 319 1174
rect -319 1108 -311 1136
rect -283 1108 -245 1136
rect -217 1108 -179 1136
rect -151 1108 -113 1136
rect -85 1108 -47 1136
rect -19 1108 19 1136
rect 47 1108 85 1136
rect 113 1108 151 1136
rect 179 1108 217 1136
rect 245 1108 283 1136
rect 311 1108 319 1136
rect -319 1070 319 1108
rect -319 1042 -311 1070
rect -283 1042 -245 1070
rect -217 1042 -179 1070
rect -151 1042 -113 1070
rect -85 1042 -47 1070
rect -19 1042 19 1070
rect 47 1042 85 1070
rect 113 1042 151 1070
rect 179 1042 217 1070
rect 245 1042 283 1070
rect 311 1042 319 1070
rect -319 1004 319 1042
rect -319 976 -311 1004
rect -283 976 -245 1004
rect -217 976 -179 1004
rect -151 976 -113 1004
rect -85 976 -47 1004
rect -19 976 19 1004
rect 47 976 85 1004
rect 113 976 151 1004
rect 179 976 217 1004
rect 245 976 283 1004
rect 311 976 319 1004
rect -319 938 319 976
rect -319 910 -311 938
rect -283 910 -245 938
rect -217 910 -179 938
rect -151 910 -113 938
rect -85 910 -47 938
rect -19 910 19 938
rect 47 910 85 938
rect 113 910 151 938
rect 179 910 217 938
rect 245 910 283 938
rect 311 910 319 938
rect -319 872 319 910
rect -319 844 -311 872
rect -283 844 -245 872
rect -217 844 -179 872
rect -151 844 -113 872
rect -85 844 -47 872
rect -19 844 19 872
rect 47 844 85 872
rect 113 844 151 872
rect 179 844 217 872
rect 245 844 283 872
rect 311 844 319 872
rect -319 806 319 844
rect -319 778 -311 806
rect -283 778 -245 806
rect -217 778 -179 806
rect -151 778 -113 806
rect -85 778 -47 806
rect -19 778 19 806
rect 47 778 85 806
rect 113 778 151 806
rect 179 778 217 806
rect 245 778 283 806
rect 311 778 319 806
rect -319 740 319 778
rect -319 712 -311 740
rect -283 712 -245 740
rect -217 712 -179 740
rect -151 712 -113 740
rect -85 712 -47 740
rect -19 712 19 740
rect 47 712 85 740
rect 113 712 151 740
rect 179 712 217 740
rect 245 712 283 740
rect 311 712 319 740
rect -319 674 319 712
rect -319 646 -311 674
rect -283 646 -245 674
rect -217 646 -179 674
rect -151 646 -113 674
rect -85 646 -47 674
rect -19 646 19 674
rect 47 646 85 674
rect 113 646 151 674
rect 179 646 217 674
rect 245 646 283 674
rect 311 646 319 674
rect -319 608 319 646
rect -319 580 -311 608
rect -283 580 -245 608
rect -217 580 -179 608
rect -151 580 -113 608
rect -85 580 -47 608
rect -19 580 19 608
rect 47 580 85 608
rect 113 580 151 608
rect 179 580 217 608
rect 245 580 283 608
rect 311 580 319 608
rect -319 542 319 580
rect -319 514 -311 542
rect -283 514 -245 542
rect -217 514 -179 542
rect -151 514 -113 542
rect -85 514 -47 542
rect -19 514 19 542
rect 47 514 85 542
rect 113 514 151 542
rect 179 514 217 542
rect 245 514 283 542
rect 311 514 319 542
rect -319 476 319 514
rect -319 448 -311 476
rect -283 448 -245 476
rect -217 448 -179 476
rect -151 448 -113 476
rect -85 448 -47 476
rect -19 448 19 476
rect 47 448 85 476
rect 113 448 151 476
rect 179 448 217 476
rect 245 448 283 476
rect 311 448 319 476
rect -319 410 319 448
rect -319 382 -311 410
rect -283 382 -245 410
rect -217 382 -179 410
rect -151 382 -113 410
rect -85 382 -47 410
rect -19 382 19 410
rect 47 382 85 410
rect 113 382 151 410
rect 179 382 217 410
rect 245 382 283 410
rect 311 382 319 410
rect -319 344 319 382
rect -319 316 -311 344
rect -283 316 -245 344
rect -217 316 -179 344
rect -151 316 -113 344
rect -85 316 -47 344
rect -19 316 19 344
rect 47 316 85 344
rect 113 316 151 344
rect 179 316 217 344
rect 245 316 283 344
rect 311 316 319 344
rect -319 278 319 316
rect -319 250 -311 278
rect -283 250 -245 278
rect -217 250 -179 278
rect -151 250 -113 278
rect -85 250 -47 278
rect -19 250 19 278
rect 47 250 85 278
rect 113 250 151 278
rect 179 250 217 278
rect 245 250 283 278
rect 311 250 319 278
rect -319 212 319 250
rect -319 184 -311 212
rect -283 184 -245 212
rect -217 184 -179 212
rect -151 184 -113 212
rect -85 184 -47 212
rect -19 184 19 212
rect 47 184 85 212
rect 113 184 151 212
rect 179 184 217 212
rect 245 184 283 212
rect 311 184 319 212
rect -319 146 319 184
rect -319 118 -311 146
rect -283 118 -245 146
rect -217 118 -179 146
rect -151 118 -113 146
rect -85 118 -47 146
rect -19 118 19 146
rect 47 118 85 146
rect 113 118 151 146
rect 179 118 217 146
rect 245 118 283 146
rect 311 118 319 146
rect -319 80 319 118
rect -319 52 -311 80
rect -283 52 -245 80
rect -217 52 -179 80
rect -151 52 -113 80
rect -85 52 -47 80
rect -19 52 19 80
rect 47 52 85 80
rect 113 52 151 80
rect 179 52 217 80
rect 245 52 283 80
rect 311 52 319 80
rect -319 14 319 52
rect -319 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 19 14
rect 47 -14 85 14
rect 113 -14 151 14
rect 179 -14 217 14
rect 245 -14 283 14
rect 311 -14 319 14
rect -319 -52 319 -14
rect -319 -80 -311 -52
rect -283 -80 -245 -52
rect -217 -80 -179 -52
rect -151 -80 -113 -52
rect -85 -80 -47 -52
rect -19 -80 19 -52
rect 47 -80 85 -52
rect 113 -80 151 -52
rect 179 -80 217 -52
rect 245 -80 283 -52
rect 311 -80 319 -52
rect -319 -118 319 -80
rect -319 -146 -311 -118
rect -283 -146 -245 -118
rect -217 -146 -179 -118
rect -151 -146 -113 -118
rect -85 -146 -47 -118
rect -19 -146 19 -118
rect 47 -146 85 -118
rect 113 -146 151 -118
rect 179 -146 217 -118
rect 245 -146 283 -118
rect 311 -146 319 -118
rect -319 -184 319 -146
rect -319 -212 -311 -184
rect -283 -212 -245 -184
rect -217 -212 -179 -184
rect -151 -212 -113 -184
rect -85 -212 -47 -184
rect -19 -212 19 -184
rect 47 -212 85 -184
rect 113 -212 151 -184
rect 179 -212 217 -184
rect 245 -212 283 -184
rect 311 -212 319 -184
rect -319 -250 319 -212
rect -319 -278 -311 -250
rect -283 -278 -245 -250
rect -217 -278 -179 -250
rect -151 -278 -113 -250
rect -85 -278 -47 -250
rect -19 -278 19 -250
rect 47 -278 85 -250
rect 113 -278 151 -250
rect 179 -278 217 -250
rect 245 -278 283 -250
rect 311 -278 319 -250
rect -319 -316 319 -278
rect -319 -344 -311 -316
rect -283 -344 -245 -316
rect -217 -344 -179 -316
rect -151 -344 -113 -316
rect -85 -344 -47 -316
rect -19 -344 19 -316
rect 47 -344 85 -316
rect 113 -344 151 -316
rect 179 -344 217 -316
rect 245 -344 283 -316
rect 311 -344 319 -316
rect -319 -382 319 -344
rect -319 -410 -311 -382
rect -283 -410 -245 -382
rect -217 -410 -179 -382
rect -151 -410 -113 -382
rect -85 -410 -47 -382
rect -19 -410 19 -382
rect 47 -410 85 -382
rect 113 -410 151 -382
rect 179 -410 217 -382
rect 245 -410 283 -382
rect 311 -410 319 -382
rect -319 -448 319 -410
rect -319 -476 -311 -448
rect -283 -476 -245 -448
rect -217 -476 -179 -448
rect -151 -476 -113 -448
rect -85 -476 -47 -448
rect -19 -476 19 -448
rect 47 -476 85 -448
rect 113 -476 151 -448
rect 179 -476 217 -448
rect 245 -476 283 -448
rect 311 -476 319 -448
rect -319 -514 319 -476
rect -319 -542 -311 -514
rect -283 -542 -245 -514
rect -217 -542 -179 -514
rect -151 -542 -113 -514
rect -85 -542 -47 -514
rect -19 -542 19 -514
rect 47 -542 85 -514
rect 113 -542 151 -514
rect 179 -542 217 -514
rect 245 -542 283 -514
rect 311 -542 319 -514
rect -319 -580 319 -542
rect -319 -608 -311 -580
rect -283 -608 -245 -580
rect -217 -608 -179 -580
rect -151 -608 -113 -580
rect -85 -608 -47 -580
rect -19 -608 19 -580
rect 47 -608 85 -580
rect 113 -608 151 -580
rect 179 -608 217 -580
rect 245 -608 283 -580
rect 311 -608 319 -580
rect -319 -646 319 -608
rect -319 -674 -311 -646
rect -283 -674 -245 -646
rect -217 -674 -179 -646
rect -151 -674 -113 -646
rect -85 -674 -47 -646
rect -19 -674 19 -646
rect 47 -674 85 -646
rect 113 -674 151 -646
rect 179 -674 217 -646
rect 245 -674 283 -646
rect 311 -674 319 -646
rect -319 -712 319 -674
rect -319 -740 -311 -712
rect -283 -740 -245 -712
rect -217 -740 -179 -712
rect -151 -740 -113 -712
rect -85 -740 -47 -712
rect -19 -740 19 -712
rect 47 -740 85 -712
rect 113 -740 151 -712
rect 179 -740 217 -712
rect 245 -740 283 -712
rect 311 -740 319 -712
rect -319 -778 319 -740
rect -319 -806 -311 -778
rect -283 -806 -245 -778
rect -217 -806 -179 -778
rect -151 -806 -113 -778
rect -85 -806 -47 -778
rect -19 -806 19 -778
rect 47 -806 85 -778
rect 113 -806 151 -778
rect 179 -806 217 -778
rect 245 -806 283 -778
rect 311 -806 319 -778
rect -319 -844 319 -806
rect -319 -872 -311 -844
rect -283 -872 -245 -844
rect -217 -872 -179 -844
rect -151 -872 -113 -844
rect -85 -872 -47 -844
rect -19 -872 19 -844
rect 47 -872 85 -844
rect 113 -872 151 -844
rect 179 -872 217 -844
rect 245 -872 283 -844
rect 311 -872 319 -844
rect -319 -910 319 -872
rect -319 -938 -311 -910
rect -283 -938 -245 -910
rect -217 -938 -179 -910
rect -151 -938 -113 -910
rect -85 -938 -47 -910
rect -19 -938 19 -910
rect 47 -938 85 -910
rect 113 -938 151 -910
rect 179 -938 217 -910
rect 245 -938 283 -910
rect 311 -938 319 -910
rect -319 -976 319 -938
rect -319 -1004 -311 -976
rect -283 -1004 -245 -976
rect -217 -1004 -179 -976
rect -151 -1004 -113 -976
rect -85 -1004 -47 -976
rect -19 -1004 19 -976
rect 47 -1004 85 -976
rect 113 -1004 151 -976
rect 179 -1004 217 -976
rect 245 -1004 283 -976
rect 311 -1004 319 -976
rect -319 -1042 319 -1004
rect -319 -1070 -311 -1042
rect -283 -1070 -245 -1042
rect -217 -1070 -179 -1042
rect -151 -1070 -113 -1042
rect -85 -1070 -47 -1042
rect -19 -1070 19 -1042
rect 47 -1070 85 -1042
rect 113 -1070 151 -1042
rect 179 -1070 217 -1042
rect 245 -1070 283 -1042
rect 311 -1070 319 -1042
rect -319 -1108 319 -1070
rect -319 -1136 -311 -1108
rect -283 -1136 -245 -1108
rect -217 -1136 -179 -1108
rect -151 -1136 -113 -1108
rect -85 -1136 -47 -1108
rect -19 -1136 19 -1108
rect 47 -1136 85 -1108
rect 113 -1136 151 -1108
rect 179 -1136 217 -1108
rect 245 -1136 283 -1108
rect 311 -1136 319 -1108
rect -319 -1174 319 -1136
rect -319 -1202 -311 -1174
rect -283 -1202 -245 -1174
rect -217 -1202 -179 -1174
rect -151 -1202 -113 -1174
rect -85 -1202 -47 -1174
rect -19 -1202 19 -1174
rect 47 -1202 85 -1174
rect 113 -1202 151 -1174
rect 179 -1202 217 -1174
rect 245 -1202 283 -1174
rect 311 -1202 319 -1174
rect -319 -1240 319 -1202
rect -319 -1268 -311 -1240
rect -283 -1268 -245 -1240
rect -217 -1268 -179 -1240
rect -151 -1268 -113 -1240
rect -85 -1268 -47 -1240
rect -19 -1268 19 -1240
rect 47 -1268 85 -1240
rect 113 -1268 151 -1240
rect 179 -1268 217 -1240
rect 245 -1268 283 -1240
rect 311 -1268 319 -1240
rect -319 -1306 319 -1268
rect -319 -1334 -311 -1306
rect -283 -1334 -245 -1306
rect -217 -1334 -179 -1306
rect -151 -1334 -113 -1306
rect -85 -1334 -47 -1306
rect -19 -1334 19 -1306
rect 47 -1334 85 -1306
rect 113 -1334 151 -1306
rect 179 -1334 217 -1306
rect 245 -1334 283 -1306
rect 311 -1334 319 -1306
rect -319 -1372 319 -1334
rect -319 -1400 -311 -1372
rect -283 -1400 -245 -1372
rect -217 -1400 -179 -1372
rect -151 -1400 -113 -1372
rect -85 -1400 -47 -1372
rect -19 -1400 19 -1372
rect 47 -1400 85 -1372
rect 113 -1400 151 -1372
rect 179 -1400 217 -1372
rect 245 -1400 283 -1372
rect 311 -1400 319 -1372
rect -319 -1438 319 -1400
rect -319 -1466 -311 -1438
rect -283 -1466 -245 -1438
rect -217 -1466 -179 -1438
rect -151 -1466 -113 -1438
rect -85 -1466 -47 -1438
rect -19 -1466 19 -1438
rect 47 -1466 85 -1438
rect 113 -1466 151 -1438
rect 179 -1466 217 -1438
rect 245 -1466 283 -1438
rect 311 -1466 319 -1438
rect -319 -1504 319 -1466
rect -319 -1532 -311 -1504
rect -283 -1532 -245 -1504
rect -217 -1532 -179 -1504
rect -151 -1532 -113 -1504
rect -85 -1532 -47 -1504
rect -19 -1532 19 -1504
rect 47 -1532 85 -1504
rect 113 -1532 151 -1504
rect 179 -1532 217 -1504
rect 245 -1532 283 -1504
rect 311 -1532 319 -1504
rect -319 -1540 319 -1532
<< end >>
