* NGSPICE file created from dec_3x8_ibr_mag_flat.ext - technology: gf180mcuC

.subckt pex_dec_3x8_ibr_mag IN1 VSS VDD D0 D1 D2 D3 D4 D5 D6 D7 IN3 IN2
X0 and_3_ibr_5.nand3_mag_ibr_0.OUT IN3.t0 a_1516_n344# VSS.t5 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1 D5 and_3_ibr_6.nand3_mag_ibr_0.OUT VSS.t8 VSS.t7 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2 and_3_ibr_5.nand3_mag_ibr_0.OUT IN3.t1 VDD.t9 VDD.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 and_3_ibr_0.nand3_mag_ibr_0.OUT and_3_ibr_5.IN3 VDD.t38 VDD.t37 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 VDD IN2.t0 and_3_ibr_3.nand3_mag_ibr_0.OUT VDD.t72 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X5 D1 and_3_ibr_4.nand3_mag_ibr_0.OUT VDD.t69 VDD.t68 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 D0 and_3_ibr_0.nand3_mag_ibr_0.OUT VDD.t19 VDD.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 a_230_n344# and_3_ibr_6.IN3 VSS.t32 VSS.t2 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X8 a_230_212# and_3_ibr_5.IN3 VSS.t22 VSS.t21 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X9 a_3768_212# IN2.t1 a_3608_212# VSS.t6 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X10 and_3_ibr_3.IN1 IN3.t2 VDD.t7 VDD.t6 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 and_3_ibr_4.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 VDD.t64 VDD.t63 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X12 and_3_ibr_1.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 VDD.t55 VDD.t54 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 and_3_ibr_3.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 VDD.t53 VDD.t52 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X14 D3 and_3_ibr_5.nand3_mag_ibr_0.OUT VSS.t35 VSS.t27 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X15 and_3_ibr_5.IN3 IN1.t0 VSS.t10 VSS.t9 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X16 and_3_ibr_2.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 VDD.t51 VDD.t50 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X17 a_1516_n344# IN2.t2 a_1356_n344# VSS.t13 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X18 and_3_ibr_1.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 a_1516_212# VSS.t5 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X19 and_3_ibr_3.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 a_3768_212# VSS.t4 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X20 a_1356_n344# and_3_ibr_5.IN3 VSS.t20 VSS.t18 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X21 and_3_ibr_7.nand3_mag_ibr_0.OUT IN3.t3 a_3768_n344# VSS.t4 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X22 and_3_ibr_2.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 a_2642_212# VSS.t3 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X23 a_3768_n344# IN2.t3 a_3608_n344# VSS.t6 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X24 VDD IN2.t4 and_3_ibr_5.nand3_mag_ibr_0.OUT VDD.t39 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 D5 and_3_ibr_6.nand3_mag_ibr_0.OUT VDD.t11 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X26 and_3_ibr_5.nand3_mag_ibr_0.OUT and_3_ibr_5.IN3 VDD.t36 VDD.t35 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X27 and_3_ibr_7.nand3_mag_ibr_0.OUT IN3.t4 VDD.t5 VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X28 D4 and_3_ibr_2.nand3_mag_ibr_0.OUT VDD.t26 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X29 D6 and_3_ibr_3.nand3_mag_ibr_0.OUT VDD.t21 VDD.t20 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X30 VDD IN2.t5 and_3_ibr_7.nand3_mag_ibr_0.OUT VDD.t75 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X31 D2 and_3_ibr_1.nand3_mag_ibr_0.OUT VDD.t47 VDD.t46 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X32 D0 and_3_ibr_0.nand3_mag_ibr_0.OUT VSS.t15 VSS.t14 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X33 and_3_ibr_6.IN3 IN2.t6 VSS.t26 VSS.t25 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X34 VDD and_3_ibr_6.IN3 and_3_ibr_0.nand3_mag_ibr_0.OUT VDD.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 and_3_ibr_6.nand3_mag_ibr_0.OUT IN3.t5 a_2642_n344# VSS.t3 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X36 D3 and_3_ibr_5.nand3_mag_ibr_0.OUT VDD.t71 VDD.t70 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 D7 and_3_ibr_7.nand3_mag_ibr_0.OUT VSS.t12 VSS.t11 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X38 and_3_ibr_6.nand3_mag_ibr_0.OUT IN3.t6 VDD.t3 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X39 a_390_212# and_3_ibr_6.IN3 a_230_212# VSS.t21 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X40 and_3_ibr_1.nand3_mag_ibr_0.OUT and_3_ibr_5.IN3 VDD.t34 VDD.t33 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X41 and_3_ibr_3.nand3_mag_ibr_0.OUT IN1.t1 VDD.t13 VDD.t12 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X42 a_3608_n344# IN1.t2 VSS.t24 VSS.t23 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X43 and_3_ibr_0.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 VDD.t49 VDD.t48 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X44 and_3_ibr_2.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 VDD.t59 VDD.t58 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X45 and_3_ibr_7.nand3_mag_ibr_0.OUT IN1.t3 VDD.t17 VDD.t16 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X46 a_1356_212# and_3_ibr_5.IN3 VSS.t19 VSS.t18 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X47 D4 and_3_ibr_2.nand3_mag_ibr_0.OUT VSS.t17 VSS.t7 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X48 a_3608_212# IN1.t4 VSS.t36 VSS.t23 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X49 D1 and_3_ibr_4.nand3_mag_ibr_0.OUT VSS.t34 VSS.t14 nfet_03v3 ad=0.157p pd=1.68u as=0.152p ps=1.64u w=0.22u l=0.28u
X50 and_3_ibr_0.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 a_390_212# VSS.t21 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X51 D2 and_3_ibr_1.nand3_mag_ibr_0.OUT VSS.t28 VSS.t27 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X52 a_2482_212# and_3_ibr_6.IN3 VSS.t31 VSS.t29 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X53 D6 and_3_ibr_3.nand3_mag_ibr_0.OUT VSS.t16 VSS.t11 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X54 and_3_ibr_6.IN3 IN2.t7 VDD.t43 VDD.t42 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X55 VDD IN2.t8 and_3_ibr_1.nand3_mag_ibr_0.OUT VDD.t65 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X56 VDD IN1.t5 and_3_ibr_2.nand3_mag_ibr_0.OUT VDD.t27 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X57 and_3_ibr_4.nand3_mag_ibr_0.OUT IN3.t7 a_390_n344# VSS.t2 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X58 a_2642_n344# IN1.t6 a_2482_n344# VSS.t33 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X59 and_3_ibr_3.IN1 IN3.t8 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X60 a_390_n344# and_3_ibr_5.IN3 a_230_n344# VSS.t2 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X61 a_2482_n344# and_3_ibr_6.IN3 VSS.t30 VSS.t29 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X62 and_3_ibr_4.nand3_mag_ibr_0.OUT IN3.t9 VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X63 VDD IN1.t7 and_3_ibr_6.nand3_mag_ibr_0.OUT VDD.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X64 D7 and_3_ibr_7.nand3_mag_ibr_0.OUT VDD.t15 VDD.t14 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X65 and_3_ibr_5.IN3 IN1.t8 VDD.t45 VDD.t44 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 a_1516_212# IN2.t9 a_1356_212# VSS.t13 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X67 a_2642_212# IN1.t9 a_2482_212# VSS.t33 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X68 VDD and_3_ibr_5.IN3 and_3_ibr_4.nand3_mag_ibr_0.OUT VDD.t30 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X69 and_3_ibr_6.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 VDD.t57 VDD.t56 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 IN3.n5 IN3.t3 36.935
R1 IN3.n12 IN3.t5 36.935
R2 IN3.n19 IN3.t7 36.935
R3 IN3.n16 IN3.t0 36.7829
R4 IN3.n0 IN3.t2 25.432
R5 IN3.n5 IN3.t4 18.1962
R6 IN3.n12 IN3.t6 18.1962
R7 IN3.n19 IN3.t9 18.1962
R8 IN3.n15 IN3.t1 17.5436
R9 IN3.n1 IN3.t8 12.4441
R10 IN3.n17 IN3.n16 4.5005
R11 IN3.n22 IN3.n21 4.5005
R12 IN3.n26 IN3.n4 4.5005
R13 IN3.n20 IN3.n19 2.88176
R14 IN3.n15 IN3 2.31681
R15 IN3.n28 IN3.n27 2.24831
R16 IN3 IN3.n1 2.20644
R17 IN3.n6 IN3.n5 2.12014
R18 IN3.n13 IN3.n12 2.11861
R19 IN3.n23 IN3.n22 1.79371
R20 IN3.n25 IN3.n24 1.60479
R21 IN3.n24 IN3.n23 1.59764
R22 IN3.n10 IN3.n9 1.49986
R23 IN3.n26 IN3.n25 1.3167
R24 IN3.n24 IN3.n14 1.27535
R25 IN3.n23 IN3.n18 1.2731
R26 IN3.n22 IN3.n20 1.1306
R27 IN3.n1 IN3.n0 0.802693
R28 IN3.n16 IN3.n15 0.582843
R29 IN3.n25 IN3.n11 0.128961
R30 IN3.n18 IN3 0.0537005
R31 IN3.n21 IN3 0.0534349
R32 IN3.n14 IN3 0.0533296
R33 IN3.n9 IN3 0.0532041
R34 IN3.n21 IN3 0.0371102
R35 IN3.n11 IN3.n10 0.0273966
R36 IN3.n14 IN3.n13 0.0222526
R37 IN3 IN3.n26 0.0183125
R38 IN3.n18 IN3.n17 0.0173852
R39 IN3.n4 IN3.n3 0.0161522
R40 IN3.n8 IN3.n7 0.0122391
R41 IN3.n9 IN3.n8 0.00925458
R42 IN3.n27 IN3 0.008
R43 IN3 IN3.n29 0.00734783
R44 IN3.n17 IN3 0.00692857
R45 IN3.n29 IN3.n28 0.00637401
R46 IN3.n28 IN3.n4 0.00637401
R47 IN3.n13 IN3 0.00468281
R48 IN3.n3 IN3.n2 0.00343478
R49 IN3.n7 IN3.n6 0.00306851
R50 IN3.n6 IN3 0.00284273
R51 IN3 IN3.n20 0.00176228
R52 VSS.t4 VSS.t11 1310.38
R53 VSS.t3 VSS.t7 1310.38
R54 VSS.t5 VSS.t27 1310.38
R55 VSS.t7 VSS.t23 1303.89
R56 VSS.t27 VSS.t29 1303.89
R57 VSS.t14 VSS.t18 1303.89
R58 VSS.n33 VSS.t14 655.191
R59 VSS.t6 VSS.t4 518.962
R60 VSS.t33 VSS.t3 518.962
R61 VSS.t13 VSS.t5 518.962
R62 VSS.n32 VSS.n31 412.745
R63 VSS.n35 VSS.n34 412.745
R64 VSS.n9 VSS.t6 311.377
R65 VSS.n17 VSS.t33 311.377
R66 VSS.n26 VSS.t13 311.377
R67 VSS.t21 VSS.t9 294.406
R68 VSS.t2 VSS.t25 291.519
R69 VSS.n31 VSS.t21 216.475
R70 VSS.n35 VSS.t2 216.475
R71 VSS.n9 VSS.t23 207.585
R72 VSS.n17 VSS.t29 207.585
R73 VSS.t18 VSS.n26 207.585
R74 VSS.n33 VSS.n32 173.179
R75 VSS.n34 VSS.n33 173.179
R76 VSS.n8 VSS.n4 35.7094
R77 VSS VSS.t10 9.40995
R78 VSS VSS.t26 9.40995
R79 VSS.n24 VSS.t28 9.34566
R80 VSS.n15 VSS.t17 9.34566
R81 VSS.n3 VSS.t16 9.34566
R82 VSS.n28 VSS.t15 9.34566
R83 VSS.n41 VSS.t34 9.34566
R84 VSS.n6 VSS.t12 9.34566
R85 VSS.n5 VSS.t1 9.34566
R86 VSS.n13 VSS.t8 9.34566
R87 VSS.n22 VSS.t35 9.34566
R88 VSS.n19 VSS.t31 8.70232
R89 VSS.n19 VSS.t30 8.70232
R90 VSS.n38 VSS.t22 5.91399
R91 VSS.n38 VSS.t32 5.91399
R92 VSS.n11 VSS.t36 5.91399
R93 VSS.n11 VSS.t24 5.91399
R94 VSS.n44 VSS.t19 5.91399
R95 VSS.n44 VSS.t20 5.91399
R96 VSS.t11 VSS 5.20126
R97 VSS.n31 VSS.n30 5.2005
R98 VSS.n36 VSS.n35 5.2005
R99 VSS.t7 VSS.n16 5.2005
R100 VSS.t27 VSS.n25 5.2005
R101 VSS.n27 VSS.t14 5.2005
R102 VSS.n42 VSS.t14 5.2005
R103 VSS.t7 VSS.n14 5.2005
R104 VSS.t27 VSS.n21 5.2005
R105 VSS.n34 VSS.n29 3.36413
R106 VSS.n10 VSS.n9 2.6035
R107 VSS.n18 VSS.n17 2.6035
R108 VSS.n26 VSS.n0 2.6035
R109 VSS VSS.n4 2.60126
R110 VSS.n8 VSS.n7 2.6005
R111 VSS.t11 VSS.n8 2.6005
R112 VSS.n4 VSS.t0 2.6005
R113 VSS.n39 VSS.n29 0.919774
R114 VSS.n14 VSS.n12 0.273398
R115 VSS.n21 VSS.n20 0.262705
R116 VSS.n43 VSS.n42 0.249789
R117 VSS.n7 VSS.n5 0.240248
R118 VSS.n37 VSS.n36 0.234244
R119 VSS.n15 VSS 0.154224
R120 VSS.n3 VSS 0.154224
R121 VSS VSS.n28 0.154224
R122 VSS.n41 VSS 0.154224
R123 VSS.n6 VSS 0.154224
R124 VSS.n13 VSS 0.154224
R125 VSS VSS.n22 0.154224
R126 VSS.n24 VSS 0.1528
R127 VSS.n40 VSS.n39 0.119812
R128 VSS.n10 VSS.n2 0.119812
R129 VSS.n18 VSS.n1 0.119812
R130 VSS.n23 VSS.n0 0.119812
R131 VSS.n19 VSS 0.0706835
R132 VSS VSS.n24 0.0647857
R133 VSS VSS.n15 0.0647857
R134 VSS VSS.n3 0.0647857
R135 VSS.n28 VSS 0.0647857
R136 VSS VSS.n41 0.0647857
R137 VSS.n5 VSS 0.0647857
R138 VSS VSS.n6 0.0647857
R139 VSS VSS.n13 0.0647857
R140 VSS.n22 VSS 0.0647857
R141 VSS VSS.n38 0.0578853
R142 VSS.n11 VSS 0.0578853
R143 VSS VSS.n44 0.0549954
R144 VSS.n38 VSS.n37 0.0372431
R145 VSS.n12 VSS.n11 0.0372431
R146 VSS.n44 VSS.n43 0.0372431
R147 VSS.n20 VSS.n19 0.0242273
R148 VSS.n40 VSS 0.021555
R149 VSS VSS.n40 0.021555
R150 VSS VSS.n2 0.021555
R151 VSS VSS.n2 0.021555
R152 VSS VSS.n1 0.021555
R153 VSS VSS.n1 0.021555
R154 VSS VSS.n23 0.021555
R155 VSS.n23 VSS 0.021555
R156 VSS.n39 VSS 0.00215138
R157 VSS VSS.n10 0.00215138
R158 VSS VSS.n18 0.00215138
R159 VSS VSS.n0 0.00215138
R160 VSS.n25 VSS 0.0012563
R161 VSS.n16 VSS 0.0012563
R162 VSS.n36 VSS 0.0012563
R163 VSS VSS.n27 0.0012563
R164 VSS.n42 VSS 0.0012563
R165 VSS.n30 VSS 0.0012563
R166 VSS.n7 VSS 0.0012563
R167 VSS.n14 VSS 0.0012563
R168 VSS VSS.n21 0.0012563
R169 D5.n1 D5.n0 6.74465
R170 D5 D5.n2 5.13104
R171 D5.n1 D5 4.65319
R172 D5 D5.n1 0.150788
R173 VDD.t52 VDD.n50 765.153
R174 VDD.t50 VDD.t25 765.152
R175 VDD.t54 VDD.t46 765.152
R176 VDD.t48 VDD.t18 765.152
R177 VDD.t10 VDD.t2 765.152
R178 VDD.t70 VDD.t8 765.152
R179 VDD.t68 VDD.t0 765.152
R180 VDD.n59 VDD.t12 759.471
R181 VDD.n65 VDD.t58 759.471
R182 VDD.n67 VDD.t33 759.471
R183 VDD.t37 VDD.n72 759.471
R184 VDD.t16 VDD.n40 759.471
R185 VDD.t56 VDD.n38 759.471
R186 VDD.t35 VDD.n36 759.471
R187 VDD.t63 VDD.n34 759.471
R188 VDD.t14 VDD.t4 749.85
R189 VDD.t6 VDD.n42 730.909
R190 VDD.t72 VDD.t52 303.031
R191 VDD.t27 VDD.t50 303.031
R192 VDD.t65 VDD.t54 303.031
R193 VDD.t60 VDD.t48 303.031
R194 VDD.t4 VDD.t75 303.031
R195 VDD.t2 VDD.t22 303.031
R196 VDD.t8 VDD.t39 303.031
R197 VDD.t0 VDD.t30 303.031
R198 VDD.n51 VDD.t72 193.183
R199 VDD.n60 VDD.t27 193.183
R200 VDD.n66 VDD.t65 193.183
R201 VDD.n73 VDD.t60 193.183
R202 VDD.t75 VDD.n41 193.183
R203 VDD.t22 VDD.n39 193.183
R204 VDD.t39 VDD.n37 193.183
R205 VDD.t30 VDD.n35 193.183
R206 VDD.n51 VDD.t12 109.849
R207 VDD.n60 VDD.t58 109.849
R208 VDD.t33 VDD.n66 109.849
R209 VDD.n73 VDD.t37 109.849
R210 VDD.n41 VDD.t16 109.849
R211 VDD.n39 VDD.t56 109.849
R212 VDD.n37 VDD.t35 109.849
R213 VDD.n35 VDD.t63 109.849
R214 VDD.n43 VDD.n4 35.263
R215 VDD.n50 VDD.n49 8.19491
R216 VDD.n74 VDD.n73 6.3005
R217 VDD.n77 VDD.n67 6.3005
R218 VDD.n72 VDD.n71 6.3005
R219 VDD.n34 VDD.n33 6.3005
R220 VDD.n35 VDD.n31 6.3005
R221 VDD.n36 VDD.n26 6.3005
R222 VDD.n37 VDD.n24 6.3005
R223 VDD.n38 VDD.n19 6.3005
R224 VDD.n39 VDD.n17 6.3005
R225 VDD.n40 VDD.n12 6.3005
R226 VDD.n41 VDD.n10 6.3005
R227 VDD.n52 VDD.n51 6.3005
R228 VDD.n59 VDD.n58 6.3005
R229 VDD.n61 VDD.n60 6.3005
R230 VDD.n65 VDD.n64 6.3005
R231 VDD.n79 VDD.n66 6.3005
R232 VDD.n71 VDD.t45 5.19258
R233 VDD.n33 VDD.t43 5.19258
R234 VDD.n29 VDD.t69 5.14703
R235 VDD.n22 VDD.t71 5.14703
R236 VDD.n15 VDD.t11 5.14703
R237 VDD.n3 VDD.t7 5.14703
R238 VDD.n8 VDD.t15 5.14703
R239 VDD.n57 VDD.t26 5.14703
R240 VDD.n63 VDD.t47 5.14491
R241 VDD.n76 VDD.t19 5.14046
R242 VDD.n48 VDD.t21 5.13792
R243 VDD.n70 VDD.t38 5.13287
R244 VDD.n32 VDD.t64 5.13287
R245 VDD.n25 VDD.t36 5.13287
R246 VDD.n18 VDD.t57 5.13287
R247 VDD.n11 VDD.t17 5.13287
R248 VDD.n53 VDD.t13 5.13287
R249 VDD.n78 VDD.t34 5.13287
R250 VDD.n62 VDD.t59 5.12141
R251 VDD.n43 VDD.t6 4.96868
R252 VDD.n7 VDD.n4 3.1505
R253 VDD.n42 VDD.n4 3.1505
R254 VDD.n44 VDD.n43 3.1505
R255 VDD.n75 VDD.n69 2.85787
R256 VDD.n30 VDD.n28 2.85787
R257 VDD.n23 VDD.n21 2.85787
R258 VDD.n16 VDD.n14 2.85787
R259 VDD.n9 VDD.n6 2.85787
R260 VDD.n2 VDD.n1 2.85561
R261 VDD.n47 VDD.n46 2.84433
R262 VDD.n56 VDD.n55 2.84433
R263 VDD.n69 VDD.t49 2.2755
R264 VDD.n69 VDD.n68 2.2755
R265 VDD.n28 VDD.t1 2.2755
R266 VDD.n28 VDD.n27 2.2755
R267 VDD.n21 VDD.t9 2.2755
R268 VDD.n21 VDD.n20 2.2755
R269 VDD.n14 VDD.t3 2.2755
R270 VDD.n14 VDD.n13 2.2755
R271 VDD.n6 VDD.t5 2.2755
R272 VDD.n6 VDD.n5 2.2755
R273 VDD.n46 VDD.t53 2.2755
R274 VDD.n46 VDD.n45 2.2755
R275 VDD.n55 VDD.t51 2.2755
R276 VDD.n55 VDD.n54 2.2755
R277 VDD.n1 VDD.t55 2.2755
R278 VDD.n1 VDD.n0 2.2755
R279 VDD.t25 VDD.n59 1.89444
R280 VDD.t46 VDD.n65 1.89444
R281 VDD.t18 VDD.n67 1.89444
R282 VDD.n72 VDD.t44 1.89444
R283 VDD.n40 VDD.t10 1.89444
R284 VDD.n38 VDD.t70 1.89444
R285 VDD.n36 VDD.t68 1.89444
R286 VDD.n34 VDD.t42 1.89444
R287 VDD.n42 VDD.t14 1.81868
R288 VDD VDD.n70 0.181314
R289 VDD.n78 VDD 0.181314
R290 VDD VDD.n32 0.181314
R291 VDD VDD.n25 0.181314
R292 VDD VDD.n18 0.181314
R293 VDD VDD.n11 0.181314
R294 VDD VDD.n53 0.181314
R295 VDD VDD.n62 0.181314
R296 VDD VDD.n3 0.178278
R297 VDD VDD.n75 0.163383
R298 VDD VDD.n47 0.163383
R299 VDD VDD.n56 0.163383
R300 VDD VDD.n2 0.163383
R301 VDD.n30 VDD 0.163383
R302 VDD.n23 VDD 0.163383
R303 VDD.n16 VDD 0.163383
R304 VDD.n9 VDD 0.163383
R305 VDD.n75 VDD 0.106177
R306 VDD VDD.n30 0.106177
R307 VDD VDD.n23 0.106177
R308 VDD VDD.n16 0.106177
R309 VDD VDD.n9 0.106177
R310 VDD.n47 VDD 0.106177
R311 VDD.n56 VDD 0.106177
R312 VDD VDD.n2 0.106177
R313 VDD.n74 VDD.n70 0.080629
R314 VDD.n32 VDD.n31 0.080629
R315 VDD.n25 VDD.n24 0.080629
R316 VDD.n18 VDD.n17 0.080629
R317 VDD.n11 VDD.n10 0.080629
R318 VDD.n53 VDD.n52 0.080629
R319 VDD.n62 VDD.n61 0.080629
R320 VDD VDD.n78 0.0788871
R321 VDD.n76 VDD 0.0671667
R322 VDD VDD.n29 0.0671667
R323 VDD VDD.n22 0.0671667
R324 VDD VDD.n15 0.0671667
R325 VDD VDD.n8 0.0671667
R326 VDD.n48 VDD 0.0671667
R327 VDD.n57 VDD 0.0671667
R328 VDD.n63 VDD 0.0671667
R329 VDD.n77 VDD.n76 0.0460556
R330 VDD.n29 VDD.n26 0.0460556
R331 VDD.n22 VDD.n19 0.0460556
R332 VDD.n15 VDD.n12 0.0460556
R333 VDD.n44 VDD.n3 0.0460556
R334 VDD.n8 VDD.n7 0.0460556
R335 VDD.n49 VDD.n48 0.0460556
R336 VDD.n58 VDD.n57 0.0460556
R337 VDD.n64 VDD.n63 0.0460556
R338 VDD.n79 VDD 0.00224194
R339 VDD VDD.n74 0.00166129
R340 VDD.n31 VDD 0.00166129
R341 VDD.n24 VDD 0.00166129
R342 VDD.n17 VDD 0.00166129
R343 VDD.n10 VDD 0.00166129
R344 VDD.n52 VDD 0.00166129
R345 VDD.n61 VDD 0.00166129
R346 VDD VDD.n79 0.00166129
R347 VDD.n71 VDD 0.00105556
R348 VDD VDD.n77 0.00105556
R349 VDD.n33 VDD 0.00105556
R350 VDD.n26 VDD 0.00105556
R351 VDD.n19 VDD 0.00105556
R352 VDD.n12 VDD 0.00105556
R353 VDD VDD.n44 0.00105556
R354 VDD.n7 VDD 0.00105556
R355 VDD.n49 VDD 0.00105556
R356 VDD.n58 VDD 0.00105556
R357 VDD.n64 VDD 0.00105556
R358 VDD.n50 VDD.t20 0.00101274
R359 IN2.n22 IN2.t9 36.935
R360 IN2.n10 IN2.t3 36.935
R361 IN2.n5 IN2.t1 36.859
R362 IN2.n31 IN2.t2 36.8284
R363 IN2.n39 IN2.t7 25.515
R364 IN2.n22 IN2.t8 18.1962
R365 IN2.n10 IN2.t5 18.1962
R366 IN2.n4 IN2.t0 17.5837
R367 IN2.n30 IN2.t4 17.2177
R368 IN2.n37 IN2.t6 11.0572
R369 IN2 IN2.n5 8.02236
R370 IN2.n10 IN2 8.0192
R371 IN2.n31 IN2 8.01903
R372 IN2.n35 IN2.n15 5.77472
R373 IN2.n15 IN2.n14 4.55209
R374 IN2.n26 IN2.n25 4.53206
R375 IN2.n34 IN2.n33 4.52972
R376 IN2.n27 IN2.n21 4.5005
R377 IN2.n20 IN2.n19 4.5005
R378 IN2.n33 IN2.n18 4.5005
R379 IN2.n33 IN2.n32 4.5005
R380 IN2.n32 IN2.n31 4.5005
R381 IN2.n28 IN2.n27 4.5005
R382 IN2.n17 IN2.n16 4.5005
R383 IN2.n3 IN2.n2 4.5005
R384 IN2.n6 IN2.n2 4.5005
R385 IN2.n13 IN2.n12 4.5005
R386 IN2.n30 IN2.n29 3.61051
R387 IN2.n25 IN2.n24 2.99669
R388 IN2.n36 IN2.n35 2.96291
R389 IN2.n11 IN2.n10 2.88073
R390 IN2.n40 IN2.n39 2.8805
R391 IN2.n35 IN2.n34 2.64379
R392 IN2.n15 IN2.n1 2.25429
R393 IN2.n40 IN2 2.25188
R394 IN2.n27 IN2.n26 2.2505
R395 IN2.n36 IN2.n0 2.24638
R396 IN2.n8 IN2.n7 2.24478
R397 IN2.n38 IN2.n37 2.24027
R398 IN2.n23 IN2.n22 2.11839
R399 IN2.n6 IN2.n4 1.81009
R400 IN2.n14 IN2.n8 1.63145
R401 IN2.n9 IN2.n1 1.12663
R402 IN2.n31 IN2.n30 0.857233
R403 IN2.n5 IN2.n4 0.435263
R404 IN2.n39 IN2.n38 0.249364
R405 IN2.n3 IN2 0.0768393
R406 IN2.n24 IN2 0.0752567
R407 IN2.n21 IN2 0.0719706
R408 IN2.n9 IN2 0.0464863
R409 IN2.n34 IN2.n16 0.0320584
R410 IN2.n7 IN2.n3 0.0300714
R411 IN2.n27 IN2.n20 0.0273831
R412 IN2.n19 IN2.n18 0.0269706
R413 IN2 IN2.n36 0.0237421
R414 IN2.n12 IN2.n9 0.0215918
R415 IN2.n8 IN2.n2 0.0177728
R416 IN2.n24 IN2.n23 0.016845
R417 IN2.n11 IN2 0.0099298
R418 IN2 IN2.n29 0.00976471
R419 IN2.n6 IN2 0.0095
R420 IN2.n23 IN2 0.00885048
R421 IN2.n7 IN2.n6 0.00692857
R422 IN2.n21 IN2.n18 0.00579412
R423 IN2.n32 IN2.n28 0.00579412
R424 IN2.n25 IN2.n20 0.00517532
R425 IN2.n13 IN2.n1 0.00484133
R426 IN2.n32 IN2.n29 0.00447059
R427 IN2.n28 IN2.n19 0.00314706
R428 IN2.n33 IN2.n17 0.00283766
R429 IN2.n41 IN2.n40 0.00194385
R430 IN2.n27 IN2.n17 0.00166883
R431 IN2.n26 IN2.n16 0.00166883
R432 IN2.n14 IN2.n13 0.00159756
R433 IN2.n12 IN2.n11 0.00142074
R434 IN2 IN2.n41 0.000981283
R435 IN2.n40 IN2.n0 0.000981283
R436 D1.n1 D1.n0 6.57033
R437 D1.n1 D1 5.38904
R438 D1 D1.n2 5.13104
R439 D1 D1.n1 0.18262
R440 D0.n2 D0.n1 8.64529
R441 D0 D0.n0 5.13104
R442 D0.n2 D0 2.59619
R443 D0 D0.n2 0.17112
R444 D3.n1 D3.n0 8.64364
R445 D3 D3.n2 5.13104
R446 D3.n1 D3 4.3719
R447 D3 D3.n1 0.179746
R448 IN1.n11 IN1.t6 36.7069
R449 IN1.n25 IN1.t9 36.5548
R450 IN1.n16 IN1.t3 30.9379
R451 IN1.n2 IN1.t1 30.4206
R452 IN1.n2 IN1.t4 24.7698
R453 IN1.n16 IN1.t2 24.5101
R454 IN1.n31 IN1.t8 23.4411
R455 IN1.n24 IN1.t5 17.4145
R456 IN1.n10 IN1.t7 17.3258
R457 IN1.n32 IN1.t0 10.8912
R458 IN1.n20 IN1.n14 10.468
R459 IN1 IN1.n30 8.62191
R460 IN1.n31 IN1.n0 8.02876
R461 IN1.n11 IN1 8.02168
R462 IN1.n25 IN1 8.01896
R463 IN1.n8 IN1.n7 4.5005
R464 IN1.n12 IN1.n7 4.5005
R465 IN1.n12 IN1.n11 4.5005
R466 IN1.n3 IN1.n1 4.5005
R467 IN1.n4 IN1.n1 4.5005
R468 IN1.n18 IN1.n15 4.5005
R469 IN1.n29 IN1.n28 4.5005
R470 IN1.n29 IN1.n26 4.5005
R471 IN1.n26 IN1.n25 4.5005
R472 IN1.n24 IN1.n23 3.66972
R473 IN1.n10 IN1.n9 3.63801
R474 IN1.n17 IN1.n16 2.88138
R475 IN1.n33 IN1.n32 2.40618
R476 IN1.n33 IN1.n31 2.32323
R477 IN1.n19 IN1 2.251
R478 IN1.n14 IN1.n13 2.24496
R479 IN1.n6 IN1.n5 2.2444
R480 IN1.n34 IN1.n33 2.11815
R481 IN1.n22 IN1.n21 1.66028
R482 IN1.n18 IN1.n17 1.50386
R483 IN1.n34 IN1 1.50158
R484 IN1.n27 IN1.n22 1.49405
R485 IN1.n3 IN1.n2 1.42163
R486 IN1.n25 IN1.n24 1.04377
R487 IN1.n11 IN1.n10 0.955106
R488 IN1.n21 IN1.n20 0.575955
R489 IN1.n28 IN1 0.484751
R490 IN1.n21 IN1.n6 0.381035
R491 IN1.n20 IN1.n19 0.296719
R492 IN1.n4 IN1 0.192359
R493 IN1.n15 IN1 0.0793218
R494 IN1.n8 IN1 0.041692
R495 IN1.n13 IN1.n8 0.0309412
R496 IN1.n15 IN1 0.028625
R497 IN1.n5 IN1.n4 0.0275
R498 IN1.n28 IN1.n27 0.0270385
R499 IN1.n30 IN1.n22 0.0255368
R500 IN1.n14 IN1.n7 0.0200059
R501 IN1.n6 IN1.n1 0.017373
R502 IN1.n19 IN1.n18 0.0152683
R503 IN1 IN1.n9 0.00976471
R504 IN1 IN1.n23 0.00857692
R505 IN1.n27 IN1.n26 0.00626923
R506 IN1.n5 IN1 0.006125
R507 IN1.n13 IN1.n12 0.00447059
R508 IN1.n30 IN1.n29 0.00284618
R509 IN1.n12 IN1.n9 0.00182353
R510 IN1.n17 IN1 0.0017491
R511 IN1.n26 IN1.n23 0.00165385
R512 IN1 IN1.n3 0.001625
R513 IN1.n34 IN1.n0 0.00154651
R514 IN1 IN1.n34 0.00154651
R515 D4.n2 D4.n1 8.64671
R516 D4 D4.n0 5.1189
R517 D4.n2 D4 3.99616
R518 D4 D4.n2 0.17421
R519 D6.n2 D6.n1 7.02949
R520 D6 D6.n0 5.11937
R521 D6.n2 D6 3.85641
R522 D6 D6.n2 0.164487
R523 D2.n2 D2.n1 9.16414
R524 D2.n2 D2 5.233
R525 D2 D2.n0 5.118
R526 D2 D2.n2 0.152915
R527 D7 D7.n8 5.13104
R528 D7.n2 D7.n1 4.9917
R529 D7.n3 D7 3.92264
R530 D7.n4 D7.n2 2.21368
R531 D7.n2 D7.n0 0.707829
R532 D7.n4 D7.n3 0.654546
R533 D7 D7.n7 0.161084
R534 D7.n6 D7.n5 0.0177727
R535 D7.n5 D7.n4 0.00231818
R536 D7.n7 D7.n6 0.00231818
C0 IN2 D3 0.0249f
C1 a_1356_212# and_3_ibr_6.IN3 0.00182f
C2 VDD a_1356_212# 2.21e-19
C3 IN2 a_1516_212# 0.00993f
C4 a_3608_212# IN3 5.62e-19
C5 D5 and_3_ibr_6.nand3_mag_ibr_0.OUT 0.147f
C6 D5 and_3_ibr_7.nand3_mag_ibr_0.OUT 0.0241f
C7 IN1 a_3608_212# 0.00692f
C8 a_390_n344# and_3_ibr_6.IN3 0.00216f
C9 D5 a_2642_n344# 0.00174f
C10 and_3_ibr_0.nand3_mag_ibr_0.OUT IN2 4.8e-19
C11 IN2 and_3_ibr_4.nand3_mag_ibr_0.OUT 0.0355f
C12 D5 a_2482_n344# 0.00139f
C13 D5 D3 0.0576f
C14 a_3768_n344# and_3_ibr_6.nand3_mag_ibr_0.OUT 3.58e-20
C15 D4 and_3_ibr_2.nand3_mag_ibr_0.OUT 0.142f
C16 a_390_212# and_3_ibr_5.IN3 0.00903f
C17 a_3768_n344# and_3_ibr_7.nand3_mag_ibr_0.OUT 0.0779f
C18 and_3_ibr_5.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 0.00136f
C19 a_3608_n344# and_3_ibr_6.nand3_mag_ibr_0.OUT 6.08e-20
C20 a_390_212# IN1 3.45e-20
C21 D7 D6 0.184f
C22 a_3608_n344# and_3_ibr_7.nand3_mag_ibr_0.OUT 0.0249f
C23 and_3_ibr_3.nand3_mag_ibr_0.OUT D6 0.151f
C24 and_3_ibr_5.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 0.0184f
C25 VDD and_3_ibr_5.nand3_mag_ibr_0.OUT 0.671f
C26 D1 and_3_ibr_5.IN3 0.284f
C27 D1 IN3 0.0475f
C28 D2 IN3 0.00388f
C29 D1 IN1 0.0329f
C30 a_230_212# and_3_ibr_0.nand3_mag_ibr_0.OUT 0.0249f
C31 D1 a_1356_212# 0.00123f
C32 D2 IN1 0.112f
C33 and_3_ibr_5.IN3 D0 0.118f
C34 and_3_ibr_3.IN1 and_3_ibr_6.IN3 0.779f
C35 D7 and_3_ibr_2.nand3_mag_ibr_0.OUT 1.51e-19
C36 VDD and_3_ibr_3.IN1 1.68f
C37 D6 IN3 0.00169f
C38 and_3_ibr_2.nand3_mag_ibr_0.OUT and_3_ibr_3.nand3_mag_ibr_0.OUT 6.97e-19
C39 D7 a_3768_212# 0.00156f
C40 and_3_ibr_3.nand3_mag_ibr_0.OUT a_3768_212# 0.0779f
C41 a_1516_n344# IN3 0.00193f
C42 D0 IN1 0.0354f
C43 VDD and_3_ibr_6.IN3 1.04f
C44 D5 IN2 0.0131f
C45 D1 a_390_n344# 0.00167f
C46 a_1356_212# D0 8.75e-20
C47 a_1356_n344# and_3_ibr_5.IN3 0.00657f
C48 a_1356_n344# IN3 0.00181f
C49 and_3_ibr_3.IN1 a_3608_212# 0.00175f
C50 and_3_ibr_2.nand3_mag_ibr_0.OUT IN3 3.87e-19
C51 and_3_ibr_6.nand3_mag_ibr_0.OUT D7 9.08e-20
C52 a_3768_212# IN3 2.63e-19
C53 a_230_212# IN2 4.46e-19
C54 and_3_ibr_7.nand3_mag_ibr_0.OUT D7 0.154f
C55 VDD a_3608_212# 2.21e-19
C56 and_3_ibr_2.nand3_mag_ibr_0.OUT IN1 0.351f
C57 and_3_ibr_5.IN3 and_3_ibr_1.nand3_mag_ibr_0.OUT 0.119f
C58 and_3_ibr_2.nand3_mag_ibr_0.OUT a_2642_212# 0.0779f
C59 and_3_ibr_1.nand3_mag_ibr_0.OUT IN3 0.00222f
C60 and_3_ibr_7.nand3_mag_ibr_0.OUT and_3_ibr_3.nand3_mag_ibr_0.OUT 0.00141f
C61 a_2482_212# IN3 5.62e-19
C62 a_3768_n344# IN2 0.0112f
C63 and_3_ibr_1.nand3_mag_ibr_0.OUT a_2642_212# 3.58e-20
C64 and_3_ibr_1.nand3_mag_ibr_0.OUT IN1 0.0189f
C65 a_2482_212# a_2642_212# 0.0504f
C66 IN1 a_2482_212# 0.00241f
C67 a_3608_n344# IN2 0.00741f
C68 D1 and_3_ibr_5.nand3_mag_ibr_0.OUT 0.0206f
C69 and_3_ibr_6.nand3_mag_ibr_0.OUT IN3 0.327f
C70 a_1356_212# and_3_ibr_1.nand3_mag_ibr_0.OUT 0.0249f
C71 a_390_212# and_3_ibr_3.IN1 8.64e-19
C72 and_3_ibr_7.nand3_mag_ibr_0.OUT IN3 0.35f
C73 and_3_ibr_6.nand3_mag_ibr_0.OUT IN1 0.298f
C74 and_3_ibr_5.IN3 a_230_n344# 0.00321f
C75 a_2642_n344# IN3 8.64e-19
C76 a_390_212# and_3_ibr_6.IN3 0.00418f
C77 D4 IN2 0.00535f
C78 and_3_ibr_7.nand3_mag_ibr_0.OUT IN1 0.108f
C79 D5 a_3768_n344# 7.87e-19
C80 a_2642_n344# IN1 0.00981f
C81 D1 and_3_ibr_3.IN1 0.0341f
C82 a_2482_n344# IN3 0.00181f
C83 D3 and_3_ibr_5.IN3 0.00663f
C84 D3 IN3 0.0471f
C85 a_1516_n344# and_3_ibr_5.nand3_mag_ibr_0.OUT 0.0779f
C86 a_1516_212# IN3 3.14e-19
C87 D5 a_3608_n344# 0.00132f
C88 D2 and_3_ibr_3.IN1 0.0621f
C89 a_2482_n344# IN1 0.00237f
C90 D1 and_3_ibr_6.IN3 0.0619f
C91 D1 VDD 0.218f
C92 D3 a_2642_212# 0.00126f
C93 D3 IN1 0.0422f
C94 a_1356_n344# and_3_ibr_5.nand3_mag_ibr_0.OUT 0.0249f
C95 D2 and_3_ibr_6.IN3 0.169f
C96 and_3_ibr_3.IN1 D0 0.0578f
C97 D3 a_1356_212# 0.00118f
C98 and_3_ibr_0.nand3_mag_ibr_0.OUT and_3_ibr_5.IN3 0.245f
C99 and_3_ibr_3.IN1 D6 0.157f
C100 VDD D2 0.245f
C101 and_3_ibr_0.nand3_mag_ibr_0.OUT IN3 5.81e-20
C102 a_1356_212# a_1516_212# 0.0504f
C103 and_3_ibr_5.IN3 and_3_ibr_4.nand3_mag_ibr_0.OUT 0.288f
C104 and_3_ibr_4.nand3_mag_ibr_0.OUT IN3 0.283f
C105 a_230_n344# a_390_n344# 0.0504f
C106 D5 D4 0.206f
C107 a_1516_n344# and_3_ibr_3.IN1 3.18e-19
C108 D0 and_3_ibr_6.IN3 0.106f
C109 and_3_ibr_0.nand3_mag_ibr_0.OUT IN1 0.0275f
C110 VDD D0 0.204f
C111 VDD D6 0.579f
C112 and_3_ibr_5.nand3_mag_ibr_0.OUT and_3_ibr_1.nand3_mag_ibr_0.OUT 0.00141f
C113 IN2 D7 0.0384f
C114 a_3608_n344# a_3768_n344# 0.0504f
C115 a_1516_n344# and_3_ibr_6.IN3 0.00103f
C116 a_1356_n344# and_3_ibr_3.IN1 5.51e-19
C117 IN2 and_3_ibr_3.nand3_mag_ibr_0.OUT 0.24f
C118 and_3_ibr_0.nand3_mag_ibr_0.OUT a_1356_212# 6.08e-20
C119 and_3_ibr_2.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 0.321f
C120 a_1356_n344# and_3_ibr_6.IN3 8.19e-19
C121 and_3_ibr_3.IN1 a_3768_212# 0.00244f
C122 a_1356_n344# VDD 2.21e-19
C123 and_3_ibr_6.nand3_mag_ibr_0.OUT and_3_ibr_5.nand3_mag_ibr_0.OUT 6.66e-19
C124 and_3_ibr_2.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 0.127f
C125 and_3_ibr_3.IN1 and_3_ibr_1.nand3_mag_ibr_0.OUT 0.317f
C126 VDD and_3_ibr_2.nand3_mag_ibr_0.OUT 0.729f
C127 and_3_ibr_3.IN1 a_2482_212# 0.00175f
C128 a_390_n344# and_3_ibr_4.nand3_mag_ibr_0.OUT 0.0779f
C129 a_2642_n344# and_3_ibr_5.nand3_mag_ibr_0.OUT 3.58e-20
C130 IN2 and_3_ibr_5.IN3 0.379f
C131 IN2 IN3 1.72f
C132 D1 a_390_212# 0.00167f
C133 and_3_ibr_1.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 0.0785f
C134 D5 D7 0.0512f
C135 and_3_ibr_6.IN3 a_2482_212# 0.00699f
C136 VDD and_3_ibr_1.nand3_mag_ibr_0.OUT 0.714f
C137 D5 and_3_ibr_3.nand3_mag_ibr_0.OUT 6.71e-19
C138 VDD a_2482_212# 2.21e-19
C139 IN2 IN1 0.353f
C140 and_3_ibr_6.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 3.53e-19
C141 a_2482_n344# and_3_ibr_5.nand3_mag_ibr_0.OUT 6.08e-20
C142 and_3_ibr_5.nand3_mag_ibr_0.OUT D3 0.144f
C143 IN2 a_1356_212# 0.00731f
C144 and_3_ibr_2.nand3_mag_ibr_0.OUT a_3608_212# 6.08e-20
C145 and_3_ibr_7.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 0.00275f
C146 and_3_ibr_6.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 0.11f
C147 a_3608_212# a_3768_212# 0.0504f
C148 and_3_ibr_6.nand3_mag_ibr_0.OUT VDD 0.671f
C149 a_230_n344# and_3_ibr_6.IN3 0.00284f
C150 a_2642_n344# and_3_ibr_6.IN3 0.00297f
C151 a_2482_n344# and_3_ibr_3.IN1 5.51e-19
C152 VDD and_3_ibr_7.nand3_mag_ibr_0.OUT 0.67f
C153 D5 IN3 0.0491f
C154 a_3768_n344# D7 0.00172f
C155 VDD a_230_n344# 2.21e-19
C156 IN2 a_390_n344# 3.58e-20
C157 and_3_ibr_5.nand3_mag_ibr_0.OUT and_3_ibr_4.nand3_mag_ibr_0.OUT 6.66e-19
C158 D3 and_3_ibr_3.IN1 0.0448f
C159 and_3_ibr_3.IN1 a_1516_212# 0.00193f
C160 D1 D0 0.318f
C161 a_2482_n344# and_3_ibr_6.IN3 0.00699f
C162 D5 IN1 0.323f
C163 D5 a_2642_212# 0.00174f
C164 a_3608_n344# D7 0.00153f
C165 a_2482_n344# VDD 2.21e-19
C166 D3 and_3_ibr_6.IN3 0.153f
C167 VDD D3 0.21f
C168 a_1516_212# and_3_ibr_6.IN3 0.00194f
C169 D1 a_1516_n344# 8.68e-19
C170 and_3_ibr_0.nand3_mag_ibr_0.OUT and_3_ibr_3.IN1 0.271f
C171 a_230_212# and_3_ibr_5.IN3 0.0079f
C172 and_3_ibr_3.IN1 and_3_ibr_4.nand3_mag_ibr_0.OUT 5.81e-20
C173 a_3768_n344# IN3 0.00168f
C174 D4 D7 0.0503f
C175 D1 a_1356_n344# 0.00148f
C176 a_230_212# IN1 5.87e-20
C177 and_3_ibr_0.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 0.263f
C178 D4 and_3_ibr_3.nand3_mag_ibr_0.OUT 0.0295f
C179 and_3_ibr_0.nand3_mag_ibr_0.OUT VDD 0.712f
C180 and_3_ibr_4.nand3_mag_ibr_0.OUT and_3_ibr_6.IN3 0.133f
C181 VDD and_3_ibr_4.nand3_mag_ibr_0.OUT 0.671f
C182 a_3608_n344# IN3 0.00181f
C183 IN2 and_3_ibr_5.nand3_mag_ibr_0.OUT 0.259f
C184 D2 and_3_ibr_2.nand3_mag_ibr_0.OUT 0.031f
C185 D1 and_3_ibr_1.nand3_mag_ibr_0.OUT 6.58e-19
C186 a_3608_n344# IN1 0.00692f
C187 D4 IN3 1.44e-21
C188 D2 and_3_ibr_1.nand3_mag_ibr_0.OUT 0.139f
C189 a_1356_n344# a_1516_n344# 0.0504f
C190 D6 a_3768_212# 2.34e-19
C191 IN2 and_3_ibr_3.IN1 0.428f
C192 D4 IN1 0.0946f
C193 D0 and_3_ibr_1.nand3_mag_ibr_0.OUT 0.0266f
C194 IN2 and_3_ibr_6.IN3 0.294f
C195 D5 and_3_ibr_5.nand3_mag_ibr_0.OUT 2.54e-21
C196 D7 and_3_ibr_3.nand3_mag_ibr_0.OUT 0.0334f
C197 D1 a_230_n344# 0.00132f
C198 IN2 VDD 2.02f
C199 and_3_ibr_2.nand3_mag_ibr_0.OUT a_3768_212# 3.58e-20
C200 a_390_212# and_3_ibr_0.nand3_mag_ibr_0.OUT 0.0779f
C201 D1 D3 0.0415f
C202 D1 a_1516_212# 7.02e-19
C203 and_3_ibr_7.nand3_mag_ibr_0.OUT D6 3.42e-19
C204 D5 and_3_ibr_3.IN1 0.0593f
C205 and_3_ibr_2.nand3_mag_ibr_0.OUT and_3_ibr_1.nand3_mag_ibr_0.OUT 6.94e-19
C206 and_3_ibr_2.nand3_mag_ibr_0.OUT a_2482_212# 0.0249f
C207 IN2 a_3608_212# 0.00741f
C208 D3 D2 0.208f
C209 D7 IN3 0.0922f
C210 and_3_ibr_3.nand3_mag_ibr_0.OUT IN3 0.00223f
C211 D5 and_3_ibr_6.IN3 0.00791f
C212 D5 VDD 0.219f
C213 D1 and_3_ibr_0.nand3_mag_ibr_0.OUT 0.0179f
C214 and_3_ibr_1.nand3_mag_ibr_0.OUT a_2482_212# 6.08e-20
C215 D3 D0 0.0371f
C216 D7 IN1 0.011f
C217 D1 and_3_ibr_4.nand3_mag_ibr_0.OUT 0.147f
C218 and_3_ibr_3.nand3_mag_ibr_0.OUT IN1 0.111f
C219 and_3_ibr_6.nand3_mag_ibr_0.OUT and_3_ibr_2.nand3_mag_ibr_0.OUT 0.00141f
C220 a_1516_212# D0 5.38e-20
C221 a_1516_n344# D3 0.0011f
C222 a_3768_n344# and_3_ibr_3.IN1 6.46e-19
C223 and_3_ibr_5.IN3 IN3 0.293f
C224 a_230_212# and_3_ibr_6.IN3 0.00284f
C225 and_3_ibr_0.nand3_mag_ibr_0.OUT D0 0.146f
C226 a_1356_n344# D3 0.00101f
C227 a_230_212# VDD 2.09e-19
C228 D5 a_3608_212# 0.00124f
C229 a_3608_n344# and_3_ibr_3.IN1 5.51e-19
C230 and_3_ibr_5.IN3 IN1 0.168f
C231 IN1 IN3 0.353f
C232 D3 and_3_ibr_2.nand3_mag_ibr_0.OUT 8.8e-19
C233 a_1516_n344# and_3_ibr_4.nand3_mag_ibr_0.OUT 3.58e-20
C234 and_3_ibr_5.IN3 a_1356_212# 0.00657f
C235 a_1356_212# IN3 5.62e-19
C236 IN1 a_2642_212# 0.0115f
C237 a_3608_n344# VDD 2.21e-19
C238 D3 and_3_ibr_1.nand3_mag_ibr_0.OUT 0.0244f
C239 and_3_ibr_6.nand3_mag_ibr_0.OUT and_3_ibr_7.nand3_mag_ibr_0.OUT 6.66e-19
C240 a_1356_n344# and_3_ibr_4.nand3_mag_ibr_0.OUT 6.08e-20
C241 D3 a_2482_212# 0.0016f
C242 D1 IN2 0.0127f
C243 a_2642_n344# and_3_ibr_6.nand3_mag_ibr_0.OUT 0.0779f
C244 a_1516_212# and_3_ibr_1.nand3_mag_ibr_0.OUT 0.0779f
C245 D4 and_3_ibr_3.IN1 0.0858f
C246 IN2 D2 0.00708f
C247 and_3_ibr_5.IN3 a_390_n344# 0.0104f
C248 a_2482_n344# and_3_ibr_6.nand3_mag_ibr_0.OUT 0.0249f
C249 a_390_n344# IN3 8.64e-19
C250 D4 VDD 0.223f
C251 and_3_ibr_6.nand3_mag_ibr_0.OUT D3 0.0244f
C252 and_3_ibr_0.nand3_mag_ibr_0.OUT and_3_ibr_1.nand3_mag_ibr_0.OUT 6.9e-19
C253 IN2 D0 0.00364f
C254 a_2482_n344# a_2642_n344# 0.0504f
C255 IN2 D6 0.00936f
C256 a_2642_n344# D3 0.00137f
C257 a_1516_n344# IN2 0.0102f
C258 a_230_212# a_390_212# 0.0504f
C259 a_2482_n344# D3 0.00174f
C260 a_1356_n344# IN2 0.00731f
C261 D5 D2 0.0233f
C262 D3 a_1516_212# 0.00116f
C263 D7 and_3_ibr_3.IN1 0.117f
C264 and_3_ibr_3.IN1 and_3_ibr_3.nand3_mag_ibr_0.OUT 0.336f
C265 a_230_n344# and_3_ibr_4.nand3_mag_ibr_0.OUT 0.0249f
C266 IN2 and_3_ibr_2.nand3_mag_ibr_0.OUT 7.8e-19
C267 and_3_ibr_5.nand3_mag_ibr_0.OUT and_3_ibr_5.IN3 0.117f
C268 and_3_ibr_5.nand3_mag_ibr_0.OUT IN3 0.344f
C269 IN2 a_3768_212# 0.0103f
C270 D1 a_230_212# 0.00132f
C271 VDD D7 0.25f
C272 and_3_ibr_0.nand3_mag_ibr_0.OUT D3 8.06e-20
C273 IN2 and_3_ibr_1.nand3_mag_ibr_0.OUT 0.216f
C274 VDD and_3_ibr_3.nand3_mag_ibr_0.OUT 0.717f
C275 and_3_ibr_5.nand3_mag_ibr_0.OUT IN1 6.84e-19
C276 and_3_ibr_0.nand3_mag_ibr_0.OUT a_1516_212# 3.58e-20
C277 and_3_ibr_3.IN1 and_3_ibr_5.IN3 0.0986f
C278 and_3_ibr_3.IN1 IN3 0.221f
C279 and_3_ibr_6.nand3_mag_ibr_0.OUT IN2 0.025f
C280 and_3_ibr_0.nand3_mag_ibr_0.OUT and_3_ibr_4.nand3_mag_ibr_0.OUT 0.00141f
C281 D7 a_3608_212# 0.00153f
C282 D5 and_3_ibr_2.nand3_mag_ibr_0.OUT 0.0249f
C283 and_3_ibr_5.IN3 and_3_ibr_6.IN3 0.546f
C284 and_3_ibr_3.IN1 a_2642_212# 8.64e-19
C285 and_3_ibr_3.IN1 IN1 1.23f
C286 and_3_ibr_3.nand3_mag_ibr_0.OUT a_3608_212# 0.0249f
C287 and_3_ibr_6.IN3 IN3 0.0547f
C288 D5 a_3768_212# 7.36e-19
C289 IN2 and_3_ibr_7.nand3_mag_ibr_0.OUT 0.273f
C290 VDD and_3_ibr_5.IN3 0.915f
C291 VDD IN3 1.35f
C292 IN2 a_230_n344# 0.00132f
C293 and_3_ibr_3.IN1 a_1356_212# 0.00175f
C294 D5 and_3_ibr_1.nand3_mag_ibr_0.OUT 1.25e-20
C295 and_3_ibr_6.IN3 IN1 0.442f
C296 and_3_ibr_6.IN3 a_2642_212# 0.00297f
C297 D5 a_2482_212# 0.00139f
C298 VDD IN1 1.69f
C299 D7 VSS 0.484f
C300 and_3_ibr_7.nand3_mag_ibr_0.OUT VSS 0.506f
C301 a_3768_n344# VSS 0.034f
C302 a_3608_n344# VSS 0.0878f
C303 D5 VSS 0.313f
C304 and_3_ibr_6.nand3_mag_ibr_0.OUT VSS 0.507f
C305 a_2642_n344# VSS 0.034f
C306 a_2482_n344# VSS 0.0878f
C307 D3 VSS 0.355f
C308 and_3_ibr_5.nand3_mag_ibr_0.OUT VSS 0.505f
C309 a_1516_n344# VSS 0.034f
C310 a_1356_n344# VSS 0.0878f
C311 D1 VSS 0.414f
C312 and_3_ibr_4.nand3_mag_ibr_0.OUT VSS 0.507f
C313 a_390_n344# VSS 0.034f
C314 a_230_n344# VSS 0.0878f
C315 IN3 VSS 1.42f
C316 a_3768_212# VSS 0.034f
C317 a_3608_212# VSS 0.0878f
C318 a_2642_212# VSS 0.034f
C319 a_2482_212# VSS 0.0878f
C320 D6 VSS 0.305f
C321 a_1516_212# VSS 0.034f
C322 a_1356_212# VSS 0.0878f
C323 and_3_ibr_3.nand3_mag_ibr_0.OUT VSS 0.517f
C324 D4 VSS 0.134f
C325 a_390_212# VSS 0.034f
C326 a_230_212# VSS 0.0878f
C327 and_3_ibr_2.nand3_mag_ibr_0.OUT VSS 0.501f
C328 D2 VSS 0.204f
C329 and_3_ibr_1.nand3_mag_ibr_0.OUT VSS 0.501f
C330 D0 VSS 0.153f
C331 IN2 VSS 2.29f
C332 and_3_ibr_0.nand3_mag_ibr_0.OUT VSS 0.501f
C333 and_3_ibr_3.IN1 VSS 1.67f
C334 and_3_ibr_6.IN3 VSS 2.11f
C335 and_3_ibr_5.IN3 VSS 1.93f
C336 IN1 VSS 2.39f
C337 VDD VSS 19.8f
C338 IN2.n0 VSS 0.023f
C339 IN2.n1 VSS 0.00613f
C340 IN2.n2 VSS 0.0107f
C341 IN2.n3 VSS 0.00696f
C342 IN2.t0 VSS 0.0178f
C343 IN2.n4 VSS 0.0157f
C344 IN2.t1 VSS 0.0277f
C345 IN2.n5 VSS 0.0339f
C346 IN2.n6 VSS 0.00126f
C347 IN2.n7 VSS 0.00294f
C348 IN2.n8 VSS 0.101f
C349 IN2.n9 VSS 0.00458f
C350 IN2.t3 VSS 0.0278f
C351 IN2.t5 VSS 0.0183f
C352 IN2.n10 VSS 0.049f
C353 IN2.n11 VSS 7.98e-19
C354 IN2.n12 VSS 0.00328f
C355 IN2.n13 VSS 6.1e-19
C356 IN2.n14 VSS 0.106f
C357 IN2.n15 VSS 0.193f
C358 IN2.n16 VSS 0.00323f
C359 IN2.n17 VSS 3.44e-19
C360 IN2.n18 VSS 0.00244f
C361 IN2.n19 VSS 0.00224f
C362 IN2.n20 VSS 0.00302f
C363 IN2.n21 VSS 0.00413f
C364 IN2.t8 VSS 0.0183f
C365 IN2.t9 VSS 0.0278f
C366 IN2.n22 VSS 0.049f
C367 IN2.n23 VSS 0.00205f
C368 IN2.n24 VSS 0.079f
C369 IN2.n25 VSS 0.136f
C370 IN2.n26 VSS 0.00935f
C371 IN2.n27 VSS 0.00183f
C372 IN2.n28 VSS 6.11e-19
C373 IN2.n29 VSS 0.00102f
C374 IN2.t2 VSS 0.0277f
C375 IN2.t4 VSS 0.0175f
C376 IN2.n30 VSS 0.0161f
C377 IN2.n31 VSS 0.0339f
C378 IN2.n32 VSS 7.13e-19
C379 IN2.n33 VSS 0.00735f
C380 IN2.n34 VSS 0.0534f
C381 IN2.n35 VSS 0.519f
C382 IN2.n36 VSS 0.193f
C383 IN2.t6 VSS 0.00359f
C384 IN2.n37 VSS 0.0132f
C385 IN2.n38 VSS 0.00395f
C386 IN2.t7 VSS 0.0229f
C387 IN2.n39 VSS 0.0229f
C388 IN2.n40 VSS 0.00112f
C389 IN2.n41 VSS 0.00112f
C390 VDD.t55 VSS 9.68e-19
C391 VDD.n0 VSS 9.68e-19
C392 VDD.n1 VSS 0.00212f
C393 VDD.n2 VSS 0.0113f
C394 VDD.t58 VSS 0.0282f
C395 VDD.t59 VSS 0.00236f
C396 VDD.t12 VSS 0.0282f
C397 VDD.t13 VSS 0.00236f
C398 VDD.t7 VSS 0.00236f
C399 VDD.n3 VSS 0.0117f
C400 VDD.n4 VSS 0.00638f
C401 VDD.t5 VSS 9.68e-19
C402 VDD.n5 VSS 9.68e-19
C403 VDD.n6 VSS 0.00211f
C404 VDD.t15 VSS 0.00236f
C405 VDD.n7 VSS 0.00157f
C406 VDD.n8 VSS 0.00795f
C407 VDD.n9 VSS 0.0112f
C408 VDD.n10 VSS 0.00731f
C409 VDD.t17 VSS 0.00236f
C410 VDD.n11 VSS 0.0123f
C411 VDD.n12 VSS 0.00455f
C412 VDD.t3 VSS 9.68e-19
C413 VDD.n13 VSS 9.68e-19
C414 VDD.n14 VSS 0.00211f
C415 VDD.t11 VSS 0.00236f
C416 VDD.n15 VSS 0.00795f
C417 VDD.n16 VSS 0.0112f
C418 VDD.n17 VSS 0.00731f
C419 VDD.t57 VSS 0.00236f
C420 VDD.n18 VSS 0.0123f
C421 VDD.n19 VSS 0.00455f
C422 VDD.t9 VSS 9.68e-19
C423 VDD.n20 VSS 9.68e-19
C424 VDD.n21 VSS 0.00211f
C425 VDD.t71 VSS 0.00236f
C426 VDD.n22 VSS 0.00795f
C427 VDD.n23 VSS 0.0112f
C428 VDD.n24 VSS 0.00731f
C429 VDD.t36 VSS 0.00236f
C430 VDD.n25 VSS 0.0123f
C431 VDD.n26 VSS 0.00455f
C432 VDD.t1 VSS 9.68e-19
C433 VDD.n27 VSS 9.68e-19
C434 VDD.n28 VSS 0.00211f
C435 VDD.t69 VSS 0.00236f
C436 VDD.n29 VSS 0.00795f
C437 VDD.n30 VSS 0.0112f
C438 VDD.n31 VSS 0.00731f
C439 VDD.t42 VSS 0.0228f
C440 VDD.t64 VSS 0.00236f
C441 VDD.n32 VSS 0.0123f
C442 VDD.t43 VSS 0.00245f
C443 VDD.n33 VSS 0.0147f
C444 VDD.n34 VSS 0.0277f
C445 VDD.t63 VSS 0.0282f
C446 VDD.n35 VSS 0.0146f
C447 VDD.t30 VSS 0.0161f
C448 VDD.t0 VSS 0.0347f
C449 VDD.t68 VSS 0.0228f
C450 VDD.n36 VSS 0.0277f
C451 VDD.t35 VSS 0.0282f
C452 VDD.n37 VSS 0.0146f
C453 VDD.t39 VSS 0.0161f
C454 VDD.t8 VSS 0.0347f
C455 VDD.t70 VSS 0.0228f
C456 VDD.n38 VSS 0.0277f
C457 VDD.t56 VSS 0.0282f
C458 VDD.n39 VSS 0.0146f
C459 VDD.t22 VSS 0.0161f
C460 VDD.t2 VSS 0.0347f
C461 VDD.t10 VSS 0.0228f
C462 VDD.n40 VSS 0.0277f
C463 VDD.t16 VSS 0.0282f
C464 VDD.n41 VSS 0.0146f
C465 VDD.t75 VSS 0.0161f
C466 VDD.t4 VSS 0.0347f
C467 VDD.t14 VSS 0.0259f
C468 VDD.n42 VSS 0.0258f
C469 VDD.t6 VSS 0.042f
C470 VDD.n43 VSS 0.0157f
C471 VDD.n44 VSS 0.00157f
C472 VDD.t21 VSS 0.00237f
C473 VDD.t53 VSS 9.68e-19
C474 VDD.n45 VSS 9.68e-19
C475 VDD.n46 VSS 0.00213f
C476 VDD.n47 VSS 0.0115f
C477 VDD.n48 VSS 0.00824f
C478 VDD.n49 VSS 0.011f
C479 VDD.t20 VSS 1.23e-19
C480 VDD.n50 VSS 0.0482f
C481 VDD.t52 VSS 0.0347f
C482 VDD.t72 VSS 0.0161f
C483 VDD.n51 VSS 0.0146f
C484 VDD.n52 VSS 0.00731f
C485 VDD.n53 VSS 0.0123f
C486 VDD.t26 VSS 0.00236f
C487 VDD.t51 VSS 9.68e-19
C488 VDD.n54 VSS 9.68e-19
C489 VDD.n55 VSS 0.00213f
C490 VDD.n56 VSS 0.0115f
C491 VDD.n57 VSS 0.00795f
C492 VDD.n58 VSS 0.00455f
C493 VDD.n59 VSS 0.0277f
C494 VDD.t25 VSS 0.0249f
C495 VDD.t50 VSS 0.0347f
C496 VDD.t27 VSS 0.0161f
C497 VDD.n60 VSS 0.0146f
C498 VDD.n61 VSS 0.00731f
C499 VDD.n62 VSS 0.0126f
C500 VDD.t47 VSS 0.00238f
C501 VDD.n63 VSS 0.00821f
C502 VDD.n64 VSS 0.00455f
C503 VDD.n65 VSS 0.0277f
C504 VDD.t46 VSS 0.0249f
C505 VDD.t54 VSS 0.0347f
C506 VDD.t65 VSS 0.0161f
C507 VDD.n66 VSS 0.0146f
C508 VDD.t34 VSS 0.00236f
C509 VDD.t33 VSS 0.0282f
C510 VDD.n67 VSS 0.0277f
C511 VDD.t19 VSS 0.00237f
C512 VDD.t49 VSS 9.68e-19
C513 VDD.n68 VSS 9.68e-19
C514 VDD.n69 VSS 0.00211f
C515 VDD.t38 VSS 0.00236f
C516 VDD.n70 VSS 0.0123f
C517 VDD.t18 VSS 0.0249f
C518 VDD.t48 VSS 0.0347f
C519 VDD.t60 VSS 0.0161f
C520 VDD.t45 VSS 0.00245f
C521 VDD.n71 VSS 0.0147f
C522 VDD.t44 VSS 0.0248f
C523 VDD.n72 VSS 0.0277f
C524 VDD.t37 VSS 0.0282f
C525 VDD.n73 VSS 0.0146f
C526 VDD.n74 VSS 0.00731f
C527 VDD.n75 VSS 0.0112f
C528 VDD.n76 VSS 0.00814f
C529 VDD.n77 VSS 0.00455f
C530 VDD.n78 VSS 0.0123f
C531 VDD.n79 VSS 0.00487f
.ends

