magic
tech gf180mcuC
magscale 1 10
timestamp 1694514513
<< metal1 >>
rect 6149 15237 6160 15283
rect 6218 14976 6318 15386
rect 6374 15237 6385 15283
rect 6535 15141 6635 15416
rect 9419 15380 10475 15480
rect 6789 15237 6800 15283
rect 6851 15221 7294 15309
rect 7438 15301 7657 15313
rect 7438 15283 7451 15301
rect 7334 15237 7345 15283
rect 7429 15237 7451 15283
rect 7515 15237 7581 15301
rect 7645 15283 7657 15301
rect 7645 15237 7665 15283
rect 7749 15237 7760 15283
rect 7438 15225 7657 15237
rect 7831 15219 8223 15307
rect 8397 15301 8616 15313
rect 8397 15283 8409 15301
rect 8294 15237 8305 15283
rect 8389 15237 8409 15283
rect 8473 15237 8539 15301
rect 8603 15283 8616 15301
rect 8603 15237 8625 15283
rect 8709 15237 8720 15283
rect 8397 15225 8616 15237
rect 8760 15221 9203 15309
rect 9254 15237 9265 15283
rect 9349 15237 9360 15283
rect 9419 15241 9519 15380
rect 9574 15237 9585 15283
rect 9669 15237 9680 15283
rect 9749 15222 10147 15310
rect 10214 15237 10225 15283
rect 10309 15237 10320 15283
rect 10375 15241 10475 15380
rect 10534 15237 10545 15283
rect 10629 15237 10640 15283
rect 10691 15221 11134 15309
rect 11278 15301 11497 15313
rect 11278 15283 11291 15301
rect 11174 15237 11185 15283
rect 11269 15237 11291 15283
rect 11355 15237 11421 15301
rect 11485 15283 11497 15301
rect 11485 15237 11505 15283
rect 11589 15237 11600 15283
rect 11278 15225 11497 15237
rect 11671 15219 12063 15307
rect 12237 15301 12456 15313
rect 12237 15283 12249 15301
rect 12134 15237 12145 15283
rect 12229 15237 12249 15283
rect 12313 15237 12379 15301
rect 12443 15283 12456 15301
rect 12443 15237 12465 15283
rect 12549 15237 12560 15283
rect 12237 15225 12456 15237
rect 12600 15221 13043 15309
rect 13414 15304 13504 15453
rect 13094 15237 13105 15283
rect 13189 15237 13200 15283
rect 13264 15214 13676 15304
rect 13734 15237 13745 15283
rect 6535 15041 6950 15141
rect 6158 14964 6377 14976
rect 6158 14951 6171 14964
rect 5667 14920 5755 14932
rect 5667 14856 5679 14920
rect 5743 14856 5755 14920
rect 6149 14905 6171 14951
rect 6158 14900 6171 14905
rect 6235 14900 6301 14964
rect 6365 14951 6377 14964
rect 6475 14962 6694 14974
rect 6475 14951 6488 14962
rect 6365 14905 6385 14951
rect 6469 14905 6488 14951
rect 6365 14900 6377 14905
rect 6158 14888 6377 14900
rect 6475 14898 6488 14905
rect 6552 14898 6618 14962
rect 6682 14951 6694 14962
rect 6682 14905 6705 14951
rect 6850 14917 6950 15041
rect 7109 14905 7120 14951
rect 6682 14898 6694 14905
rect 6475 14886 6694 14898
rect 5667 14813 5755 14856
rect 7177 14824 7277 14949
rect 7334 14905 7345 14951
rect 7429 14905 7440 14951
rect 7486 14886 7929 14974
rect 8125 14886 8568 14974
rect 9037 14965 9256 14977
rect 9037 14951 9049 14965
rect 8614 14905 8625 14951
rect 8709 14905 8720 14951
rect 8777 14824 8877 14949
rect 8934 14905 8945 14951
rect 9029 14905 9049 14951
rect 9037 14901 9049 14905
rect 9113 14901 9179 14965
rect 9243 14951 9256 14965
rect 9360 14962 9579 14974
rect 9360 14951 9372 14962
rect 9243 14905 9265 14951
rect 9349 14905 9372 14951
rect 9243 14901 9256 14905
rect 9037 14889 9256 14901
rect 9360 14898 9372 14905
rect 9436 14898 9502 14962
rect 9566 14951 9579 14962
rect 9677 14964 9896 14976
rect 9677 14951 9689 14964
rect 9566 14905 9585 14951
rect 9669 14905 9689 14951
rect 9566 14898 9579 14905
rect 9360 14886 9579 14898
rect 9677 14900 9689 14905
rect 9753 14900 9819 14964
rect 9883 14951 9896 14964
rect 9998 14964 10217 14976
rect 9998 14951 10011 14964
rect 9883 14905 9905 14951
rect 9989 14905 10011 14951
rect 9883 14900 9896 14905
rect 9677 14888 9896 14900
rect 9998 14900 10011 14905
rect 10075 14900 10141 14964
rect 10205 14951 10217 14964
rect 10315 14962 10534 14974
rect 10315 14951 10328 14962
rect 10205 14905 10225 14951
rect 10309 14905 10328 14951
rect 10205 14900 10217 14905
rect 9998 14888 10217 14900
rect 10315 14898 10328 14905
rect 10392 14898 10458 14962
rect 10522 14951 10534 14962
rect 10638 14965 10857 14977
rect 10638 14951 10651 14965
rect 10522 14905 10545 14951
rect 10629 14905 10651 14951
rect 10522 14898 10534 14905
rect 10315 14886 10534 14898
rect 10638 14901 10651 14905
rect 10715 14901 10781 14965
rect 10845 14951 10857 14965
rect 10845 14905 10865 14951
rect 10949 14905 10960 14951
rect 10845 14901 10857 14905
rect 10638 14889 10857 14901
rect 5667 14790 6638 14813
rect 5667 14726 5679 14790
rect 5743 14726 6638 14790
rect 5667 14713 6638 14726
rect 7177 14724 7600 14824
rect 6171 14615 6306 14650
rect 6171 14562 6313 14615
rect 6374 14585 6385 14631
rect 6469 14585 6480 14631
rect 6538 14593 6638 14713
rect 6694 14585 6705 14631
rect 6789 14585 6800 14631
rect 6847 14566 7290 14654
rect 7334 14585 7345 14631
rect 7429 14585 7440 14631
rect 7500 14591 7600 14724
rect 8454 14724 8877 14824
rect 11017 14824 11117 14949
rect 11174 14905 11185 14951
rect 11269 14905 11280 14951
rect 11326 14886 11769 14974
rect 11965 14886 12408 14974
rect 12877 14965 13096 14977
rect 13576 14976 13676 15214
rect 12877 14951 12889 14965
rect 12454 14905 12465 14951
rect 12549 14905 12560 14951
rect 12617 14824 12717 14949
rect 12774 14905 12785 14951
rect 12869 14905 12889 14951
rect 12877 14901 12889 14905
rect 12953 14901 13019 14965
rect 13083 14951 13096 14965
rect 13200 14962 13419 14974
rect 13200 14951 13212 14962
rect 13083 14905 13105 14951
rect 13189 14905 13212 14951
rect 13083 14901 13096 14905
rect 12877 14889 13096 14901
rect 13200 14898 13212 14905
rect 13276 14898 13342 14962
rect 13406 14951 13419 14962
rect 13517 14964 13736 14976
rect 13517 14951 13529 14964
rect 13406 14905 13425 14951
rect 13509 14905 13529 14951
rect 13406 14898 13419 14905
rect 13200 14886 13419 14898
rect 13517 14900 13529 14905
rect 13593 14900 13659 14964
rect 13723 14951 13736 14964
rect 13723 14905 13745 14951
rect 13723 14900 13736 14905
rect 13517 14888 13736 14900
rect 7654 14585 7665 14631
rect 7749 14585 7760 14631
rect 7800 14578 8240 14666
rect 8294 14585 8305 14631
rect 8389 14585 8400 14631
rect 8454 14591 8554 14724
rect 9416 14713 10478 14813
rect 11017 14724 11440 14824
rect 8614 14585 8625 14631
rect 8709 14585 8720 14631
rect 8764 14566 9207 14654
rect 9254 14585 9265 14631
rect 9349 14585 9360 14631
rect 9416 14593 9516 14713
rect 9574 14585 9585 14631
rect 9669 14585 9680 14631
rect 9748 14562 10146 14650
rect 10214 14585 10225 14631
rect 10309 14585 10320 14631
rect 10378 14593 10478 14713
rect 10534 14585 10545 14631
rect 10629 14585 10640 14631
rect 10687 14566 11130 14654
rect 11174 14585 11185 14631
rect 11269 14585 11280 14631
rect 11340 14591 11440 14724
rect 12294 14724 12717 14824
rect 11494 14585 11505 14631
rect 11589 14585 11600 14631
rect 11643 14576 12083 14664
rect 12134 14585 12145 14631
rect 12229 14585 12240 14631
rect 12294 14591 12394 14724
rect 13256 14713 14227 14813
rect 12454 14585 12465 14631
rect 12549 14585 12560 14631
rect 12604 14566 13047 14654
rect 13094 14585 13105 14631
rect 13189 14585 13200 14631
rect 13256 14593 13356 14713
rect 13414 14585 13425 14631
rect 6213 14497 6313 14562
rect 5667 14397 6313 14497
rect 13574 14495 13674 14617
rect 5667 13847 5767 14397
rect 6213 14321 6313 14397
rect 7496 14395 8558 14495
rect 6155 14309 6374 14321
rect 6155 14299 6168 14309
rect 6149 14253 6168 14299
rect 6155 14245 6168 14253
rect 6232 14245 6298 14309
rect 6362 14299 6374 14309
rect 6477 14308 6696 14320
rect 6477 14299 6490 14308
rect 6362 14253 6385 14299
rect 6469 14253 6490 14299
rect 6362 14245 6374 14253
rect 6155 14233 6374 14245
rect 6477 14244 6490 14253
rect 6554 14244 6620 14308
rect 6684 14299 6696 14308
rect 7119 14304 7338 14316
rect 7119 14299 7132 14304
rect 6684 14253 6705 14299
rect 6789 14253 6800 14299
rect 6684 14244 6696 14253
rect 6477 14232 6696 14244
rect 6831 14150 6931 14290
rect 7014 14253 7025 14299
rect 7109 14253 7132 14299
rect 7119 14240 7132 14253
rect 7196 14240 7262 14304
rect 7326 14299 7338 14304
rect 7326 14253 7345 14299
rect 7429 14253 7440 14299
rect 7496 14258 7596 14395
rect 7759 14312 7978 14324
rect 7759 14299 7772 14312
rect 7654 14253 7665 14299
rect 7749 14253 7772 14299
rect 7326 14240 7338 14253
rect 7119 14228 7338 14240
rect 7759 14248 7772 14253
rect 7836 14248 7902 14312
rect 7966 14299 7978 14312
rect 8076 14312 8295 14324
rect 8076 14299 8088 14312
rect 7966 14253 7985 14299
rect 8069 14253 8088 14299
rect 7966 14248 7978 14253
rect 7759 14236 7978 14248
rect 8076 14248 8088 14253
rect 8152 14248 8218 14312
rect 8282 14299 8295 14312
rect 8282 14253 8305 14299
rect 8389 14253 8400 14299
rect 8458 14258 8558 14395
rect 11336 14395 12398 14495
rect 13574 14475 14060 14495
rect 13574 14411 13853 14475
rect 13917 14411 13983 14475
rect 14047 14411 14060 14475
rect 13574 14395 14060 14411
rect 8716 14304 8935 14316
rect 8716 14299 8728 14304
rect 8614 14253 8625 14299
rect 8709 14253 8728 14299
rect 8282 14248 8295 14253
rect 8076 14236 8295 14248
rect 8716 14240 8728 14253
rect 8792 14240 8858 14304
rect 8922 14299 8935 14304
rect 9358 14308 9577 14320
rect 9358 14299 9370 14308
rect 8922 14253 8945 14299
rect 9029 14253 9040 14299
rect 8922 14240 8935 14253
rect 8716 14228 8935 14240
rect 6216 14050 6931 14150
rect 7502 14052 8552 14151
rect 6149 13933 6160 13979
rect 6216 13967 6316 14050
rect 7502 14041 7601 14052
rect 6475 13989 6694 14001
rect 7118 13991 7337 14003
rect 6475 13979 6488 13989
rect 6216 13939 6317 13967
rect 6217 13847 6317 13939
rect 6374 13933 6385 13979
rect 6469 13933 6488 13979
rect 6475 13925 6488 13933
rect 6552 13925 6618 13989
rect 6682 13979 6694 13989
rect 6796 13979 7015 13990
rect 7118 13979 7131 13991
rect 6682 13933 6705 13979
rect 6789 13978 7025 13979
rect 6789 13933 6809 13978
rect 6682 13925 6694 13933
rect 6475 13913 6694 13925
rect 6796 13914 6809 13933
rect 6873 13914 6939 13978
rect 7003 13933 7025 13978
rect 7109 13933 7131 13979
rect 7003 13914 7015 13933
rect 7118 13927 7131 13933
rect 7195 13927 7261 13991
rect 7325 13979 7337 13991
rect 7325 13933 7345 13979
rect 7429 13933 7440 13979
rect 7501 13944 7601 14041
rect 8453 14041 8552 14052
rect 9123 14150 9223 14290
rect 9254 14253 9265 14299
rect 9349 14253 9370 14299
rect 9358 14244 9370 14253
rect 9434 14244 9500 14308
rect 9564 14299 9577 14308
rect 9680 14309 9899 14321
rect 9680 14299 9692 14309
rect 9564 14253 9585 14299
rect 9669 14253 9692 14299
rect 9564 14244 9577 14253
rect 9358 14232 9577 14244
rect 9680 14245 9692 14253
rect 9756 14245 9822 14309
rect 9886 14299 9899 14309
rect 9995 14309 10214 14321
rect 9995 14299 10008 14309
rect 9886 14253 9905 14299
rect 9989 14253 10008 14299
rect 9886 14245 9899 14253
rect 9680 14233 9899 14245
rect 9995 14245 10008 14253
rect 10072 14245 10138 14309
rect 10202 14299 10214 14309
rect 10317 14308 10536 14320
rect 10317 14299 10330 14308
rect 10202 14253 10225 14299
rect 10309 14253 10330 14299
rect 10202 14245 10214 14253
rect 9995 14233 10214 14245
rect 10317 14244 10330 14253
rect 10394 14244 10460 14308
rect 10524 14299 10536 14308
rect 10959 14304 11178 14316
rect 10959 14299 10972 14304
rect 10524 14253 10545 14299
rect 10629 14253 10640 14299
rect 10524 14244 10536 14253
rect 10317 14232 10536 14244
rect 10671 14150 10771 14290
rect 10854 14253 10865 14299
rect 10949 14253 10972 14299
rect 10959 14240 10972 14253
rect 11036 14240 11102 14304
rect 11166 14299 11178 14304
rect 11166 14253 11185 14299
rect 11269 14253 11280 14299
rect 11336 14258 11436 14395
rect 11599 14312 11818 14324
rect 11599 14299 11612 14312
rect 11494 14253 11505 14299
rect 11589 14253 11612 14299
rect 11166 14240 11178 14253
rect 10959 14228 11178 14240
rect 11599 14248 11612 14253
rect 11676 14248 11742 14312
rect 11806 14299 11818 14312
rect 11916 14312 12135 14324
rect 11916 14299 11928 14312
rect 11806 14253 11825 14299
rect 11909 14253 11928 14299
rect 11806 14248 11818 14253
rect 11599 14236 11818 14248
rect 11916 14248 11928 14253
rect 11992 14248 12058 14312
rect 12122 14299 12135 14312
rect 12122 14253 12145 14299
rect 12229 14253 12240 14299
rect 12298 14258 12398 14395
rect 12556 14304 12775 14316
rect 12556 14299 12568 14304
rect 12454 14253 12465 14299
rect 12549 14253 12568 14299
rect 12122 14248 12135 14253
rect 11916 14236 12135 14248
rect 12556 14240 12568 14253
rect 12632 14240 12698 14304
rect 12762 14299 12775 14304
rect 13198 14308 13417 14320
rect 13198 14299 13210 14308
rect 12762 14253 12785 14299
rect 12869 14253 12880 14299
rect 12762 14240 12775 14253
rect 12556 14228 12775 14240
rect 9123 14050 9838 14150
rect 7758 13987 7977 13999
rect 7758 13979 7771 13987
rect 7654 13933 7665 13979
rect 7749 13933 7771 13979
rect 7325 13927 7337 13933
rect 7118 13915 7337 13927
rect 7758 13923 7771 13933
rect 7835 13923 7901 13987
rect 7965 13979 7977 13987
rect 8077 13987 8296 13999
rect 8077 13979 8089 13987
rect 7965 13933 7985 13979
rect 8069 13933 8089 13979
rect 7965 13923 7977 13933
rect 6796 13902 7015 13914
rect 7758 13911 7977 13923
rect 8077 13923 8089 13933
rect 8153 13923 8219 13987
rect 8283 13979 8296 13987
rect 8283 13933 8305 13979
rect 8389 13933 8400 13979
rect 8453 13944 8553 14041
rect 8717 13991 8936 14003
rect 8717 13979 8729 13991
rect 8614 13933 8625 13979
rect 8709 13933 8729 13979
rect 8283 13923 8296 13933
rect 8077 13911 8296 13923
rect 8717 13927 8729 13933
rect 8793 13927 8859 13991
rect 8923 13979 8936 13991
rect 9039 13979 9258 13990
rect 9360 13989 9579 14001
rect 9360 13979 9372 13989
rect 8923 13933 8945 13979
rect 9029 13978 9265 13979
rect 9029 13933 9051 13978
rect 8923 13927 8936 13933
rect 8717 13915 8936 13927
rect 9039 13914 9051 13933
rect 9115 13914 9181 13978
rect 9245 13933 9265 13978
rect 9349 13933 9372 13979
rect 9245 13914 9258 13933
rect 9039 13902 9258 13914
rect 9360 13925 9372 13933
rect 9436 13925 9502 13989
rect 9566 13979 9579 13989
rect 9566 13933 9585 13979
rect 9669 13933 9680 13979
rect 9738 13939 9838 14050
rect 10056 14050 10771 14150
rect 11342 14052 12392 14151
rect 10056 13939 10156 14050
rect 11342 14041 11441 14052
rect 10315 13989 10534 14001
rect 10958 13991 11177 14003
rect 10315 13979 10328 13989
rect 10214 13933 10225 13979
rect 10309 13933 10328 13979
rect 9566 13925 9579 13933
rect 9360 13913 9579 13925
rect 10315 13925 10328 13933
rect 10392 13925 10458 13989
rect 10522 13979 10534 13989
rect 10636 13979 10855 13990
rect 10958 13979 10971 13991
rect 10522 13933 10545 13979
rect 10629 13978 10865 13979
rect 10629 13933 10649 13978
rect 10522 13925 10534 13933
rect 10315 13913 10534 13925
rect 10636 13914 10649 13933
rect 10713 13914 10779 13978
rect 10843 13933 10865 13978
rect 10949 13933 10971 13979
rect 10843 13914 10855 13933
rect 10958 13927 10971 13933
rect 11035 13927 11101 13991
rect 11165 13979 11177 13991
rect 11165 13933 11185 13979
rect 11269 13933 11280 13979
rect 11341 13944 11441 14041
rect 12293 14041 12392 14052
rect 12963 14150 13063 14290
rect 13094 14253 13105 14299
rect 13189 14253 13210 14299
rect 13198 14244 13210 14253
rect 13274 14244 13340 14308
rect 13404 14299 13417 14308
rect 13520 14309 13739 14321
rect 13520 14299 13532 14309
rect 13404 14253 13425 14299
rect 13509 14253 13532 14299
rect 13404 14244 13417 14253
rect 13198 14232 13417 14244
rect 13520 14245 13532 14253
rect 13596 14245 13662 14309
rect 13726 14299 13739 14309
rect 13726 14253 13745 14299
rect 13726 14245 13739 14253
rect 13520 14233 13739 14245
rect 12963 14050 13678 14150
rect 11598 13987 11817 13999
rect 11598 13979 11611 13987
rect 11494 13933 11505 13979
rect 11589 13933 11611 13979
rect 11165 13927 11177 13933
rect 10958 13915 11177 13927
rect 11598 13923 11611 13933
rect 11675 13923 11741 13987
rect 11805 13979 11817 13987
rect 11917 13987 12136 13999
rect 11917 13979 11929 13987
rect 11805 13933 11825 13979
rect 11909 13933 11929 13979
rect 11805 13923 11817 13933
rect 10636 13902 10855 13914
rect 11598 13911 11817 13923
rect 11917 13923 11929 13933
rect 11993 13923 12059 13987
rect 12123 13979 12136 13987
rect 12123 13933 12145 13979
rect 12229 13933 12240 13979
rect 12293 13944 12393 14041
rect 12557 13991 12776 14003
rect 12557 13979 12569 13991
rect 12454 13933 12465 13979
rect 12549 13933 12569 13979
rect 12123 13923 12136 13933
rect 11917 13911 12136 13923
rect 12557 13927 12569 13933
rect 12633 13927 12699 13991
rect 12763 13979 12776 13991
rect 12879 13979 13098 13990
rect 13200 13989 13419 14001
rect 13200 13979 13212 13989
rect 12763 13933 12785 13979
rect 12869 13978 13105 13979
rect 12869 13933 12891 13978
rect 12763 13927 12776 13933
rect 12557 13915 12776 13927
rect 12879 13914 12891 13933
rect 12955 13914 13021 13978
rect 13085 13933 13105 13978
rect 13189 13933 13212 13979
rect 13085 13914 13098 13933
rect 12879 13902 13098 13914
rect 13200 13925 13212 13933
rect 13276 13925 13342 13989
rect 13406 13979 13419 13989
rect 13406 13933 13425 13979
rect 13509 13933 13520 13979
rect 13578 13939 13678 14050
rect 13734 13933 13745 13979
rect 13406 13925 13419 13933
rect 13200 13913 13419 13925
rect 5667 13747 6317 13847
rect 6217 13579 6317 13747
rect 6534 13732 7599 13832
rect 6374 13601 6385 13647
rect 6469 13601 6480 13647
rect 6534 13606 6634 13732
rect 6694 13601 6705 13647
rect 6789 13601 6800 13647
rect 6854 13576 7297 13664
rect 7334 13601 7345 13647
rect 7429 13601 7440 13647
rect 7499 13602 7599 13732
rect 8455 13732 9520 13832
rect 7654 13601 7665 13647
rect 7749 13601 7760 13647
rect 7807 13578 8247 13666
rect 8294 13601 8305 13647
rect 8389 13601 8400 13647
rect 8455 13602 8555 13732
rect 8614 13601 8625 13647
rect 8709 13601 8720 13647
rect 8757 13576 9200 13664
rect 9254 13601 9265 13647
rect 9349 13601 9360 13647
rect 9420 13606 9520 13732
rect 10374 13732 11439 13832
rect 9574 13601 9585 13647
rect 9669 13601 9680 13647
rect 9770 13579 10124 13667
rect 10214 13601 10225 13647
rect 10309 13601 10320 13647
rect 10374 13606 10474 13732
rect 10534 13601 10545 13647
rect 10629 13601 10640 13647
rect 10694 13576 11137 13664
rect 11174 13601 11185 13647
rect 11269 13601 11280 13647
rect 11339 13602 11439 13732
rect 12295 13732 13360 13832
rect 14127 13830 14227 14713
rect 16308 14317 16396 14329
rect 16308 14253 16320 14317
rect 16384 14253 16396 14317
rect 16308 14187 16396 14253
rect 16308 14123 16320 14187
rect 16384 14123 16396 14187
rect 16308 14110 16396 14123
rect 11494 13601 11505 13647
rect 11589 13601 11600 13647
rect 11647 13578 12087 13666
rect 12134 13601 12145 13647
rect 12229 13601 12240 13647
rect 12295 13602 12395 13732
rect 12454 13601 12465 13647
rect 12549 13601 12560 13647
rect 12597 13576 13040 13664
rect 13094 13601 13105 13647
rect 13189 13601 13200 13647
rect 13260 13606 13360 13732
rect 13575 13730 14227 13830
rect 13414 13601 13425 13647
rect 13575 13604 13675 13730
rect 15908 13612 16127 13624
rect 15908 13548 15921 13612
rect 15985 13548 16051 13612
rect 16115 13548 16127 13612
rect 15908 13536 16127 13548
rect 7179 13403 8875 13503
rect 5667 13293 5755 13305
rect 5667 13229 5679 13293
rect 5743 13229 5755 13293
rect 6149 13281 6160 13327
rect 6211 13269 6654 13357
rect 6797 13339 7016 13351
rect 6797 13327 6810 13339
rect 6694 13281 6705 13327
rect 6789 13281 6810 13327
rect 6797 13275 6810 13281
rect 6874 13275 6940 13339
rect 7004 13327 7016 13339
rect 7004 13281 7025 13327
rect 7109 13281 7120 13327
rect 7179 13291 7279 13403
rect 7438 13332 7657 13344
rect 7438 13327 7451 13332
rect 7334 13281 7345 13327
rect 7429 13281 7451 13327
rect 7004 13275 7016 13281
rect 5667 13181 5755 13229
rect 6222 13181 6317 13269
rect 6797 13263 7016 13275
rect 7438 13268 7451 13281
rect 7515 13268 7581 13332
rect 7645 13327 7657 13332
rect 7758 13343 7977 13355
rect 7758 13327 7771 13343
rect 7645 13281 7665 13327
rect 7749 13281 7771 13327
rect 7645 13268 7657 13281
rect 7438 13256 7657 13268
rect 7758 13279 7771 13281
rect 7835 13279 7901 13343
rect 7965 13327 7977 13343
rect 8077 13343 8296 13355
rect 8077 13327 8089 13343
rect 7965 13281 7985 13327
rect 8069 13281 8089 13327
rect 7965 13279 7977 13281
rect 7758 13267 7977 13279
rect 8077 13279 8089 13281
rect 8153 13279 8219 13343
rect 8283 13327 8296 13343
rect 8397 13332 8616 13344
rect 8397 13327 8409 13332
rect 8283 13281 8305 13327
rect 8389 13281 8409 13327
rect 8283 13279 8296 13281
rect 8077 13267 8296 13279
rect 8397 13268 8409 13281
rect 8473 13268 8539 13332
rect 8603 13327 8616 13332
rect 8603 13281 8625 13327
rect 8709 13281 8720 13327
rect 8775 13291 8875 13403
rect 11019 13403 12715 13503
rect 9038 13339 9257 13351
rect 9038 13327 9050 13339
rect 8934 13281 8945 13327
rect 9029 13281 9050 13327
rect 8603 13268 8616 13281
rect 8397 13256 8616 13268
rect 9038 13275 9050 13281
rect 9114 13275 9180 13339
rect 9244 13327 9257 13339
rect 9244 13281 9265 13327
rect 9349 13281 9360 13327
rect 9244 13275 9257 13281
rect 9038 13263 9257 13275
rect 9400 13269 9843 13357
rect 10051 13269 10494 13357
rect 10637 13339 10856 13351
rect 10637 13327 10650 13339
rect 10534 13281 10545 13327
rect 10629 13281 10650 13327
rect 10637 13275 10650 13281
rect 10714 13275 10780 13339
rect 10844 13327 10856 13339
rect 10844 13281 10865 13327
rect 10949 13281 10960 13327
rect 11019 13291 11119 13403
rect 11278 13332 11497 13344
rect 11278 13327 11291 13332
rect 11174 13281 11185 13327
rect 11269 13281 11291 13327
rect 10844 13275 10856 13281
rect 10637 13263 10856 13275
rect 11278 13268 11291 13281
rect 11355 13268 11421 13332
rect 11485 13327 11497 13332
rect 11598 13343 11817 13355
rect 11598 13327 11611 13343
rect 11485 13281 11505 13327
rect 11589 13281 11611 13327
rect 11485 13268 11497 13281
rect 11278 13256 11497 13268
rect 11598 13279 11611 13281
rect 11675 13279 11741 13343
rect 11805 13327 11817 13343
rect 11917 13343 12136 13355
rect 11917 13327 11929 13343
rect 11805 13281 11825 13327
rect 11909 13281 11929 13327
rect 11805 13279 11817 13281
rect 11598 13267 11817 13279
rect 11917 13279 11929 13281
rect 11993 13279 12059 13343
rect 12123 13327 12136 13343
rect 12237 13332 12456 13344
rect 12237 13327 12249 13332
rect 12123 13281 12145 13327
rect 12229 13281 12249 13327
rect 12123 13279 12136 13281
rect 11917 13267 12136 13279
rect 12237 13268 12249 13281
rect 12313 13268 12379 13332
rect 12443 13327 12456 13332
rect 12443 13281 12465 13327
rect 12549 13281 12560 13327
rect 12615 13291 12715 13403
rect 15913 13369 16132 13381
rect 12878 13339 13097 13351
rect 12878 13327 12890 13339
rect 12774 13281 12785 13327
rect 12869 13281 12890 13327
rect 12443 13268 12456 13281
rect 12237 13256 12456 13268
rect 12878 13275 12890 13281
rect 12954 13275 13020 13339
rect 13084 13327 13097 13339
rect 13084 13281 13105 13327
rect 13189 13281 13200 13327
rect 13084 13275 13097 13281
rect 12878 13263 13097 13275
rect 13240 13269 13683 13357
rect 13734 13281 13745 13327
rect 15913 13305 15926 13369
rect 15990 13305 16056 13369
rect 16120 13305 16132 13369
rect 15913 13293 16132 13305
rect 5667 13163 6317 13181
rect 5667 13099 5679 13163
rect 5743 13099 6317 13163
rect 5667 13086 6317 13099
rect 6222 12925 6317 13086
rect 13581 13182 13676 13269
rect 13581 13087 14227 13182
rect 6374 12949 6385 12995
rect 6469 12949 6480 12995
rect 6538 12872 6638 12994
rect 6694 12949 6705 12995
rect 6789 12949 6800 12995
rect 6855 12928 7298 13016
rect 7334 12949 7345 12995
rect 7429 12949 7440 12995
rect 7491 12872 7591 12987
rect 7654 12949 7665 12995
rect 7749 12949 7760 12995
rect 7811 12924 8243 13012
rect 8294 12949 8305 12995
rect 8389 12949 8400 12995
rect 6538 12772 7591 12872
rect 8463 12872 8563 12987
rect 8614 12949 8625 12995
rect 8709 12949 8720 12995
rect 8756 12928 9199 13016
rect 9254 12949 9265 12995
rect 9349 12949 9360 12995
rect 9416 12872 9516 12994
rect 9574 12949 9585 12995
rect 9669 12949 9680 12995
rect 9731 12925 10134 13013
rect 10214 12949 10225 12995
rect 10309 12949 10320 12995
rect 8463 12772 9516 12872
rect 10378 12872 10478 12994
rect 10534 12949 10545 12995
rect 10629 12949 10640 12995
rect 10695 12928 11138 13016
rect 11174 12949 11185 12995
rect 11269 12949 11280 12995
rect 11331 12872 11431 12987
rect 11494 12949 11505 12995
rect 11589 12949 11600 12995
rect 11651 12924 12083 13012
rect 12134 12949 12145 12995
rect 12229 12949 12240 12995
rect 10378 12772 11431 12872
rect 12303 12872 12403 12987
rect 12454 12949 12465 12995
rect 12549 12949 12560 12995
rect 12596 12928 13039 13016
rect 13581 13013 13676 13087
rect 13094 12949 13105 12995
rect 13189 12949 13200 12995
rect 13256 12872 13356 12994
rect 13414 12949 13425 12995
rect 13509 12949 13520 12995
rect 13572 12925 13676 13013
rect 12303 12772 13356 12872
rect 6435 10417 6535 10827
rect 6752 10682 6852 10826
rect 9804 10821 11028 10921
rect 7068 10662 7511 10750
rect 7655 10742 7874 10754
rect 7655 10678 7668 10742
rect 7732 10678 7798 10742
rect 7862 10678 7874 10742
rect 7655 10666 7874 10678
rect 8048 10660 8608 10748
rect 8782 10742 9001 10754
rect 8782 10678 8794 10742
rect 8858 10678 8924 10742
rect 8988 10678 9001 10742
rect 8782 10666 9001 10678
rect 9145 10662 9588 10750
rect 9804 10682 9904 10821
rect 10134 10663 10700 10751
rect 10928 10682 11028 10821
rect 11244 10662 11687 10750
rect 11831 10742 12050 10754
rect 11831 10678 11844 10742
rect 11908 10678 11974 10742
rect 12038 10678 12050 10742
rect 11831 10666 12050 10678
rect 12224 10660 12784 10748
rect 12958 10742 13177 10754
rect 12958 10678 12970 10742
rect 13034 10678 13100 10742
rect 13164 10678 13177 10742
rect 12958 10666 13177 10678
rect 13321 10662 13764 10750
rect 13980 10682 14080 10826
rect 6375 10405 6594 10417
rect 6375 10341 6388 10405
rect 6452 10341 6518 10405
rect 6582 10341 6594 10405
rect 6375 10329 6594 10341
rect 6692 10403 6911 10415
rect 6692 10339 6705 10403
rect 6769 10339 6835 10403
rect 6899 10339 6911 10403
rect 6692 10327 6911 10339
rect 7015 10406 7234 10418
rect 7015 10342 7028 10406
rect 7092 10342 7158 10406
rect 7222 10342 7234 10406
rect 7015 10330 7234 10342
rect 7394 10265 7494 10390
rect 7703 10327 8146 10415
rect 8510 10327 8953 10415
rect 9422 10406 9641 10418
rect 9162 10265 9262 10390
rect 9422 10342 9434 10406
rect 9498 10342 9564 10406
rect 9628 10342 9641 10406
rect 9422 10330 9641 10342
rect 9745 10403 9964 10415
rect 9745 10339 9757 10403
rect 9821 10339 9887 10403
rect 9951 10339 9964 10403
rect 9745 10327 9964 10339
rect 10062 10405 10281 10417
rect 10062 10341 10074 10405
rect 10138 10341 10204 10405
rect 10268 10341 10281 10405
rect 10062 10329 10281 10341
rect 10551 10405 10770 10417
rect 10551 10341 10564 10405
rect 10628 10341 10694 10405
rect 10758 10341 10770 10405
rect 10551 10329 10770 10341
rect 10868 10403 11087 10415
rect 10868 10339 10881 10403
rect 10945 10339 11011 10403
rect 11075 10339 11087 10403
rect 10868 10327 11087 10339
rect 11191 10406 11410 10418
rect 11191 10342 11204 10406
rect 11268 10342 11334 10406
rect 11398 10342 11410 10406
rect 11191 10330 11410 10342
rect 6210 10154 6855 10254
rect 7394 10165 7817 10265
rect 6210 10056 6523 10091
rect 6210 10003 6530 10056
rect 6755 10034 6855 10154
rect 7064 10007 7507 10095
rect 7717 10032 7817 10165
rect 8839 10165 9262 10265
rect 11570 10265 11670 10390
rect 11879 10327 12322 10415
rect 12686 10327 13129 10415
rect 13598 10406 13817 10418
rect 14297 10417 14397 10827
rect 13338 10265 13438 10390
rect 13598 10342 13610 10406
rect 13674 10342 13740 10406
rect 13804 10342 13817 10406
rect 13598 10330 13817 10342
rect 13921 10403 14140 10415
rect 13921 10339 13933 10403
rect 13997 10339 14063 10403
rect 14127 10339 14140 10403
rect 13921 10327 14140 10339
rect 14238 10405 14457 10417
rect 14238 10341 14250 10405
rect 14314 10341 14380 10405
rect 14444 10341 14457 10405
rect 14238 10329 14457 10341
rect 8017 10019 8625 10107
rect 8839 10032 8939 10165
rect 9801 10154 11031 10254
rect 11570 10165 11993 10265
rect 9149 10007 9592 10095
rect 9801 10034 9901 10154
rect 10133 10003 10699 10091
rect 10931 10034 11031 10154
rect 11240 10007 11683 10095
rect 11893 10032 11993 10165
rect 13015 10165 13438 10265
rect 12196 10017 12804 10105
rect 13015 10032 13115 10165
rect 13977 10154 14630 10254
rect 13325 10007 13768 10095
rect 13977 10034 14077 10154
rect 14309 10003 14630 10091
rect 6430 9762 6530 10003
rect 7713 9836 8943 9936
rect 6372 9750 6591 9762
rect 6372 9686 6385 9750
rect 6449 9686 6515 9750
rect 6579 9686 6591 9750
rect 6372 9674 6591 9686
rect 6694 9749 6913 9761
rect 6694 9685 6707 9749
rect 6771 9685 6837 9749
rect 6901 9685 6913 9749
rect 7336 9745 7555 9757
rect 6694 9673 6913 9685
rect 7048 9591 7148 9731
rect 7336 9681 7349 9745
rect 7413 9681 7479 9745
rect 7543 9681 7555 9745
rect 7713 9699 7813 9836
rect 7976 9753 8195 9765
rect 7336 9669 7555 9681
rect 7976 9689 7989 9753
rect 8053 9689 8119 9753
rect 8183 9689 8195 9753
rect 7976 9677 8195 9689
rect 8461 9753 8680 9765
rect 8461 9689 8473 9753
rect 8537 9689 8603 9753
rect 8667 9689 8680 9753
rect 8843 9699 8943 9836
rect 11889 9836 13119 9936
rect 9101 9745 9320 9757
rect 8461 9677 8680 9689
rect 9101 9681 9113 9745
rect 9177 9681 9243 9745
rect 9307 9681 9320 9745
rect 9743 9749 9962 9761
rect 9101 9669 9320 9681
rect 6433 9491 7148 9591
rect 7719 9493 8937 9592
rect 6433 9408 6533 9491
rect 7719 9482 7818 9493
rect 6692 9430 6911 9442
rect 7335 9432 7554 9444
rect 6433 9380 6534 9408
rect 6434 9108 6534 9380
rect 6692 9366 6705 9430
rect 6769 9366 6835 9430
rect 6899 9366 6911 9430
rect 6692 9354 6911 9366
rect 7013 9419 7232 9431
rect 7013 9355 7026 9419
rect 7090 9355 7156 9419
rect 7220 9355 7232 9419
rect 7335 9368 7348 9432
rect 7412 9368 7478 9432
rect 7542 9368 7554 9432
rect 7718 9385 7818 9482
rect 8838 9482 8937 9493
rect 9508 9591 9608 9731
rect 9743 9685 9755 9749
rect 9819 9685 9885 9749
rect 9949 9685 9962 9749
rect 9743 9673 9962 9685
rect 10065 9750 10284 9762
rect 10065 9686 10077 9750
rect 10141 9686 10207 9750
rect 10271 9686 10284 9750
rect 10065 9674 10284 9686
rect 10548 9750 10767 9762
rect 10548 9686 10561 9750
rect 10625 9686 10691 9750
rect 10755 9686 10767 9750
rect 10548 9674 10767 9686
rect 10870 9749 11089 9761
rect 10870 9685 10883 9749
rect 10947 9685 11013 9749
rect 11077 9685 11089 9749
rect 11512 9745 11731 9757
rect 10870 9673 11089 9685
rect 11224 9591 11324 9731
rect 11512 9681 11525 9745
rect 11589 9681 11655 9745
rect 11719 9681 11731 9745
rect 11889 9699 11989 9836
rect 12152 9753 12371 9765
rect 11512 9669 11731 9681
rect 12152 9689 12165 9753
rect 12229 9689 12295 9753
rect 12359 9689 12371 9753
rect 12152 9677 12371 9689
rect 12637 9753 12856 9765
rect 12637 9689 12649 9753
rect 12713 9689 12779 9753
rect 12843 9689 12856 9753
rect 13019 9699 13119 9836
rect 13277 9745 13496 9757
rect 12637 9677 12856 9689
rect 13277 9681 13289 9745
rect 13353 9681 13419 9745
rect 13483 9681 13496 9745
rect 13919 9749 14138 9761
rect 13277 9669 13496 9681
rect 9508 9491 10223 9591
rect 7975 9428 8194 9440
rect 7335 9356 7554 9368
rect 7975 9364 7988 9428
rect 8052 9364 8118 9428
rect 8182 9364 8194 9428
rect 7013 9343 7232 9355
rect 7975 9352 8194 9364
rect 8462 9428 8681 9440
rect 8462 9364 8474 9428
rect 8538 9364 8604 9428
rect 8668 9364 8681 9428
rect 8838 9385 8938 9482
rect 9102 9432 9321 9444
rect 8462 9352 8681 9364
rect 9102 9368 9114 9432
rect 9178 9368 9244 9432
rect 9308 9368 9321 9432
rect 9102 9356 9321 9368
rect 9424 9419 9643 9431
rect 9424 9355 9436 9419
rect 9500 9355 9566 9419
rect 9630 9355 9643 9419
rect 9424 9343 9643 9355
rect 9745 9430 9964 9442
rect 9745 9366 9757 9430
rect 9821 9366 9887 9430
rect 9951 9366 9964 9430
rect 10123 9380 10223 9491
rect 10609 9491 11324 9591
rect 11895 9493 13113 9592
rect 10609 9380 10709 9491
rect 11895 9482 11994 9493
rect 10868 9430 11087 9442
rect 11511 9432 11730 9444
rect 9745 9354 9964 9366
rect 10868 9366 10881 9430
rect 10945 9366 11011 9430
rect 11075 9366 11087 9430
rect 10868 9354 11087 9366
rect 11189 9419 11408 9431
rect 11189 9355 11202 9419
rect 11266 9355 11332 9419
rect 11396 9355 11408 9419
rect 11511 9368 11524 9432
rect 11588 9368 11654 9432
rect 11718 9368 11730 9432
rect 11894 9385 11994 9482
rect 13014 9482 13113 9493
rect 13684 9591 13784 9731
rect 13919 9685 13931 9749
rect 13995 9685 14061 9749
rect 14125 9685 14138 9749
rect 13919 9673 14138 9685
rect 14241 9750 14460 9762
rect 14241 9686 14253 9750
rect 14317 9686 14383 9750
rect 14447 9686 14460 9750
rect 14241 9674 14460 9686
rect 13684 9491 14399 9591
rect 12151 9428 12370 9440
rect 11511 9356 11730 9368
rect 12151 9364 12164 9428
rect 12228 9364 12294 9428
rect 12358 9364 12370 9428
rect 11189 9343 11408 9355
rect 12151 9352 12370 9364
rect 12638 9428 12857 9440
rect 12638 9364 12650 9428
rect 12714 9364 12780 9428
rect 12844 9364 12857 9428
rect 13014 9385 13114 9482
rect 13278 9432 13497 9444
rect 12638 9352 12857 9364
rect 13278 9368 13290 9432
rect 13354 9368 13420 9432
rect 13484 9368 13497 9432
rect 13278 9356 13497 9368
rect 13600 9419 13819 9431
rect 13600 9355 13612 9419
rect 13676 9355 13742 9419
rect 13806 9355 13819 9419
rect 13600 9343 13819 9355
rect 13921 9430 14140 9442
rect 13921 9366 13933 9430
rect 13997 9366 14063 9430
rect 14127 9366 14140 9430
rect 14299 9380 14399 9491
rect 13921 9354 14140 9366
rect 6210 9050 6534 9108
rect 6751 9173 7816 9273
rect 6210 9020 6501 9050
rect 6751 9047 6851 9173
rect 7071 9017 7514 9105
rect 7716 9043 7816 9173
rect 8840 9173 9905 9273
rect 8024 9019 8632 9107
rect 8840 9043 8940 9173
rect 9142 9017 9585 9105
rect 9805 9047 9905 9173
rect 10927 9173 11992 9273
rect 10155 9020 10677 9108
rect 10927 9047 11027 9173
rect 11247 9017 11690 9105
rect 11892 9043 11992 9173
rect 13016 9173 14081 9273
rect 12200 9019 12808 9107
rect 13016 9043 13116 9173
rect 13318 9017 13761 9105
rect 13981 9047 14081 9173
rect 14331 9020 14560 9108
rect 7396 8844 9260 8944
rect 6428 8710 6871 8798
rect 7014 8780 7233 8792
rect 7014 8716 7027 8780
rect 7091 8716 7157 8780
rect 7221 8716 7233 8780
rect 7396 8732 7496 8844
rect 7655 8773 7874 8785
rect 6439 8454 6534 8710
rect 7014 8704 7233 8716
rect 7655 8709 7668 8773
rect 7732 8709 7798 8773
rect 7862 8709 7874 8773
rect 7655 8697 7874 8709
rect 7975 8784 8194 8796
rect 7975 8720 7988 8784
rect 8052 8720 8118 8784
rect 8182 8720 8194 8784
rect 7975 8708 8194 8720
rect 8462 8784 8681 8796
rect 8462 8720 8474 8784
rect 8538 8720 8604 8784
rect 8668 8720 8681 8784
rect 8462 8708 8681 8720
rect 8782 8773 9001 8785
rect 8782 8709 8794 8773
rect 8858 8709 8924 8773
rect 8988 8709 9001 8773
rect 9160 8732 9260 8844
rect 11572 8844 13436 8944
rect 9423 8780 9642 8792
rect 8782 8697 9001 8709
rect 9423 8716 9435 8780
rect 9499 8716 9565 8780
rect 9629 8716 9642 8780
rect 9423 8704 9642 8716
rect 9785 8710 10228 8798
rect 10604 8710 11047 8798
rect 11190 8780 11409 8792
rect 11190 8716 11203 8780
rect 11267 8716 11333 8780
rect 11397 8716 11409 8780
rect 11572 8732 11672 8844
rect 11831 8773 12050 8785
rect 11190 8704 11409 8716
rect 11831 8709 11844 8773
rect 11908 8709 11974 8773
rect 12038 8709 12050 8773
rect 11831 8697 12050 8709
rect 12151 8784 12370 8796
rect 12151 8720 12164 8784
rect 12228 8720 12294 8784
rect 12358 8720 12370 8784
rect 12151 8708 12370 8720
rect 12638 8784 12857 8796
rect 12638 8720 12650 8784
rect 12714 8720 12780 8784
rect 12844 8720 12857 8784
rect 12638 8708 12857 8720
rect 12958 8773 13177 8785
rect 12958 8709 12970 8773
rect 13034 8709 13100 8773
rect 13164 8709 13177 8773
rect 13336 8732 13436 8844
rect 13599 8780 13818 8792
rect 12958 8697 13177 8709
rect 13599 8716 13611 8780
rect 13675 8716 13741 8780
rect 13805 8716 13818 8780
rect 13599 8704 13818 8716
rect 13961 8710 14404 8798
rect 6210 8407 6534 8454
rect 6210 8366 6511 8407
rect 6755 8313 6855 8435
rect 7072 8369 7515 8457
rect 7708 8313 7808 8428
rect 8028 8365 8628 8453
rect 6755 8213 7808 8313
rect 8848 8313 8948 8428
rect 9141 8369 9584 8457
rect 9801 8313 9901 8435
rect 10116 8366 10687 8454
rect 8848 8213 9901 8313
rect 10931 8313 11031 8435
rect 11248 8369 11691 8457
rect 11884 8313 11984 8428
rect 12204 8365 12804 8453
rect 10931 8213 11984 8313
rect 13024 8313 13124 8428
rect 13317 8369 13760 8457
rect 14302 8454 14397 8710
rect 13977 8313 14077 8435
rect 14293 8366 14630 8454
rect 13024 8213 14077 8313
rect 5587 1473 5687 1617
rect 5904 1472 6004 1616
rect 6220 1452 6663 1540
rect 6807 1532 7026 1544
rect 6807 1468 6820 1532
rect 6884 1468 6950 1532
rect 7014 1468 7026 1532
rect 6807 1456 7026 1468
rect 7200 1450 7643 1538
rect 4448 1269 4667 1281
rect 4448 1205 4461 1269
rect 4525 1205 4591 1269
rect 4655 1205 4667 1269
rect 4448 1193 4667 1205
rect 5527 1195 5746 1207
rect 5527 1131 5540 1195
rect 5604 1131 5670 1195
rect 5734 1131 5746 1195
rect 5527 1119 5746 1131
rect 5844 1193 6063 1205
rect 5844 1129 5857 1193
rect 5921 1129 5987 1193
rect 6051 1129 6063 1193
rect 5844 1117 6063 1129
rect 6167 1196 6386 1208
rect 6167 1132 6180 1196
rect 6244 1132 6310 1196
rect 6374 1132 6386 1196
rect 6167 1120 6386 1132
rect 6546 1055 6646 1180
rect 6855 1117 7298 1205
rect 4453 1026 4672 1038
rect 4453 962 4466 1026
rect 4530 962 4596 1026
rect 4660 962 4672 1026
rect 4453 950 4672 962
rect 5233 944 6007 1044
rect 6546 955 6969 1055
rect 5232 785 5675 873
rect 5907 816 6007 944
rect 6216 789 6659 877
rect 6869 814 6969 955
rect 7192 933 7642 1033
rect 7192 810 7292 933
rect 6865 618 7626 718
rect 5524 532 5743 544
rect 5524 468 5537 532
rect 5601 468 5667 532
rect 5731 468 5743 532
rect 5524 456 5743 468
rect 5846 531 6065 543
rect 5846 467 5859 531
rect 5923 467 5989 531
rect 6053 467 6065 531
rect 6488 527 6707 539
rect 5846 455 6065 467
rect 6200 373 6300 513
rect 6488 463 6501 527
rect 6565 463 6631 527
rect 6695 463 6707 527
rect 6865 481 6965 618
rect 7128 535 7347 547
rect 6488 451 6707 463
rect 7128 471 7141 535
rect 7205 471 7271 535
rect 7335 471 7347 535
rect 7128 459 7347 471
rect 4347 141 4447 285
rect 5585 273 6300 373
rect 6871 275 7601 374
rect 5585 154 5685 273
rect 6871 258 6970 275
rect 5844 204 6063 216
rect 6487 206 6706 218
rect 5844 140 5857 204
rect 5921 140 5987 204
rect 6051 140 6063 204
rect 5844 128 6063 140
rect 6165 193 6384 205
rect 6165 129 6178 193
rect 6242 129 6308 193
rect 6372 129 6384 193
rect 6487 142 6500 206
rect 6564 142 6630 206
rect 6694 142 6706 206
rect 6870 159 6970 258
rect 7127 202 7346 214
rect 6487 130 6706 142
rect 7127 138 7140 202
rect 7204 138 7270 202
rect 7334 138 7346 202
rect 6165 117 6384 129
rect 7127 126 7346 138
rect 5903 -53 6968 47
rect 5210 -206 5653 -118
rect 5903 -179 6003 -53
rect 6223 -209 6666 -121
rect 6868 -183 6968 -53
rect 7176 -207 7619 -119
rect 6548 -382 7619 -282
rect 5580 -524 6023 -436
rect 6166 -454 6385 -442
rect 6166 -518 6179 -454
rect 6243 -518 6309 -454
rect 6373 -518 6385 -454
rect 6548 -502 6648 -382
rect 6807 -461 7026 -449
rect 6166 -530 6385 -518
rect 6807 -525 6820 -461
rect 6884 -525 6950 -461
rect 7014 -525 7026 -461
rect 6807 -537 7026 -525
rect 7127 -450 7346 -438
rect 7127 -514 7140 -450
rect 7204 -514 7270 -450
rect 7334 -514 7346 -450
rect 7127 -526 7346 -514
rect 5220 -868 5663 -780
rect 5907 -921 6007 -799
rect 6224 -865 6667 -777
rect 6860 -921 6960 -806
rect 7180 -869 7623 -781
rect 5907 -1021 6960 -921
<< via1 >>
rect 7451 15237 7515 15301
rect 7581 15237 7645 15301
rect 8409 15237 8473 15301
rect 8539 15237 8603 15301
rect 11291 15237 11355 15301
rect 11421 15237 11485 15301
rect 12249 15237 12313 15301
rect 12379 15237 12443 15301
rect 5679 14856 5743 14920
rect 6171 14900 6235 14964
rect 6301 14900 6365 14964
rect 6488 14898 6552 14962
rect 6618 14898 6682 14962
rect 9049 14901 9113 14965
rect 9179 14901 9243 14965
rect 9372 14898 9436 14962
rect 9502 14898 9566 14962
rect 9689 14900 9753 14964
rect 9819 14900 9883 14964
rect 10011 14900 10075 14964
rect 10141 14900 10205 14964
rect 10328 14898 10392 14962
rect 10458 14898 10522 14962
rect 10651 14901 10715 14965
rect 10781 14901 10845 14965
rect 5679 14726 5743 14790
rect 12889 14901 12953 14965
rect 13019 14901 13083 14965
rect 13212 14898 13276 14962
rect 13342 14898 13406 14962
rect 13529 14900 13593 14964
rect 13659 14900 13723 14964
rect 6168 14245 6232 14309
rect 6298 14245 6362 14309
rect 6490 14244 6554 14308
rect 6620 14244 6684 14308
rect 7132 14240 7196 14304
rect 7262 14240 7326 14304
rect 7772 14248 7836 14312
rect 7902 14248 7966 14312
rect 8088 14248 8152 14312
rect 8218 14248 8282 14312
rect 13853 14411 13917 14475
rect 13983 14411 14047 14475
rect 8728 14240 8792 14304
rect 8858 14240 8922 14304
rect 6488 13925 6552 13989
rect 6618 13925 6682 13989
rect 6809 13914 6873 13978
rect 6939 13914 7003 13978
rect 7131 13927 7195 13991
rect 7261 13927 7325 13991
rect 9370 14244 9434 14308
rect 9500 14244 9564 14308
rect 9692 14245 9756 14309
rect 9822 14245 9886 14309
rect 10008 14245 10072 14309
rect 10138 14245 10202 14309
rect 10330 14244 10394 14308
rect 10460 14244 10524 14308
rect 10972 14240 11036 14304
rect 11102 14240 11166 14304
rect 11612 14248 11676 14312
rect 11742 14248 11806 14312
rect 11928 14248 11992 14312
rect 12058 14248 12122 14312
rect 12568 14240 12632 14304
rect 12698 14240 12762 14304
rect 7771 13923 7835 13987
rect 7901 13923 7965 13987
rect 8089 13923 8153 13987
rect 8219 13923 8283 13987
rect 8729 13927 8793 13991
rect 8859 13927 8923 13991
rect 9051 13914 9115 13978
rect 9181 13914 9245 13978
rect 9372 13925 9436 13989
rect 9502 13925 9566 13989
rect 10328 13925 10392 13989
rect 10458 13925 10522 13989
rect 10649 13914 10713 13978
rect 10779 13914 10843 13978
rect 10971 13927 11035 13991
rect 11101 13927 11165 13991
rect 13210 14244 13274 14308
rect 13340 14244 13404 14308
rect 13532 14245 13596 14309
rect 13662 14245 13726 14309
rect 11611 13923 11675 13987
rect 11741 13923 11805 13987
rect 11929 13923 11993 13987
rect 12059 13923 12123 13987
rect 12569 13927 12633 13991
rect 12699 13927 12763 13991
rect 12891 13914 12955 13978
rect 13021 13914 13085 13978
rect 13212 13925 13276 13989
rect 13342 13925 13406 13989
rect 16320 14253 16384 14317
rect 16320 14123 16384 14187
rect 15921 13548 15985 13612
rect 16051 13548 16115 13612
rect 5679 13229 5743 13293
rect 6810 13275 6874 13339
rect 6940 13275 7004 13339
rect 7451 13268 7515 13332
rect 7581 13268 7645 13332
rect 7771 13279 7835 13343
rect 7901 13279 7965 13343
rect 8089 13279 8153 13343
rect 8219 13279 8283 13343
rect 8409 13268 8473 13332
rect 8539 13268 8603 13332
rect 9050 13275 9114 13339
rect 9180 13275 9244 13339
rect 10650 13275 10714 13339
rect 10780 13275 10844 13339
rect 11291 13268 11355 13332
rect 11421 13268 11485 13332
rect 11611 13279 11675 13343
rect 11741 13279 11805 13343
rect 11929 13279 11993 13343
rect 12059 13279 12123 13343
rect 12249 13268 12313 13332
rect 12379 13268 12443 13332
rect 12890 13275 12954 13339
rect 13020 13275 13084 13339
rect 15926 13305 15990 13369
rect 16056 13305 16120 13369
rect 5679 13099 5743 13163
rect 7668 10678 7732 10742
rect 7798 10678 7862 10742
rect 8794 10678 8858 10742
rect 8924 10678 8988 10742
rect 11844 10678 11908 10742
rect 11974 10678 12038 10742
rect 12970 10678 13034 10742
rect 13100 10678 13164 10742
rect 6388 10341 6452 10405
rect 6518 10341 6582 10405
rect 6705 10339 6769 10403
rect 6835 10339 6899 10403
rect 7028 10342 7092 10406
rect 7158 10342 7222 10406
rect 9434 10342 9498 10406
rect 9564 10342 9628 10406
rect 9757 10339 9821 10403
rect 9887 10339 9951 10403
rect 10074 10341 10138 10405
rect 10204 10341 10268 10405
rect 10564 10341 10628 10405
rect 10694 10341 10758 10405
rect 10881 10339 10945 10403
rect 11011 10339 11075 10403
rect 11204 10342 11268 10406
rect 11334 10342 11398 10406
rect 13610 10342 13674 10406
rect 13740 10342 13804 10406
rect 13933 10339 13997 10403
rect 14063 10339 14127 10403
rect 14250 10341 14314 10405
rect 14380 10341 14444 10405
rect 6385 9686 6449 9750
rect 6515 9686 6579 9750
rect 6707 9685 6771 9749
rect 6837 9685 6901 9749
rect 7349 9681 7413 9745
rect 7479 9681 7543 9745
rect 7989 9689 8053 9753
rect 8119 9689 8183 9753
rect 8473 9689 8537 9753
rect 8603 9689 8667 9753
rect 9113 9681 9177 9745
rect 9243 9681 9307 9745
rect 6705 9366 6769 9430
rect 6835 9366 6899 9430
rect 7026 9355 7090 9419
rect 7156 9355 7220 9419
rect 7348 9368 7412 9432
rect 7478 9368 7542 9432
rect 9755 9685 9819 9749
rect 9885 9685 9949 9749
rect 10077 9686 10141 9750
rect 10207 9686 10271 9750
rect 10561 9686 10625 9750
rect 10691 9686 10755 9750
rect 10883 9685 10947 9749
rect 11013 9685 11077 9749
rect 11525 9681 11589 9745
rect 11655 9681 11719 9745
rect 12165 9689 12229 9753
rect 12295 9689 12359 9753
rect 12649 9689 12713 9753
rect 12779 9689 12843 9753
rect 13289 9681 13353 9745
rect 13419 9681 13483 9745
rect 7988 9364 8052 9428
rect 8118 9364 8182 9428
rect 8474 9364 8538 9428
rect 8604 9364 8668 9428
rect 9114 9368 9178 9432
rect 9244 9368 9308 9432
rect 9436 9355 9500 9419
rect 9566 9355 9630 9419
rect 9757 9366 9821 9430
rect 9887 9366 9951 9430
rect 10881 9366 10945 9430
rect 11011 9366 11075 9430
rect 11202 9355 11266 9419
rect 11332 9355 11396 9419
rect 11524 9368 11588 9432
rect 11654 9368 11718 9432
rect 13931 9685 13995 9749
rect 14061 9685 14125 9749
rect 14253 9686 14317 9750
rect 14383 9686 14447 9750
rect 12164 9364 12228 9428
rect 12294 9364 12358 9428
rect 12650 9364 12714 9428
rect 12780 9364 12844 9428
rect 13290 9368 13354 9432
rect 13420 9368 13484 9432
rect 13612 9355 13676 9419
rect 13742 9355 13806 9419
rect 13933 9366 13997 9430
rect 14063 9366 14127 9430
rect 7027 8716 7091 8780
rect 7157 8716 7221 8780
rect 7668 8709 7732 8773
rect 7798 8709 7862 8773
rect 7988 8720 8052 8784
rect 8118 8720 8182 8784
rect 8474 8720 8538 8784
rect 8604 8720 8668 8784
rect 8794 8709 8858 8773
rect 8924 8709 8988 8773
rect 9435 8716 9499 8780
rect 9565 8716 9629 8780
rect 11203 8716 11267 8780
rect 11333 8716 11397 8780
rect 11844 8709 11908 8773
rect 11974 8709 12038 8773
rect 12164 8720 12228 8784
rect 12294 8720 12358 8784
rect 12650 8720 12714 8784
rect 12780 8720 12844 8784
rect 12970 8709 13034 8773
rect 13100 8709 13164 8773
rect 13611 8716 13675 8780
rect 13741 8716 13805 8780
rect 6820 1468 6884 1532
rect 6950 1468 7014 1532
rect 4461 1205 4525 1269
rect 4591 1205 4655 1269
rect 5540 1131 5604 1195
rect 5670 1131 5734 1195
rect 5857 1129 5921 1193
rect 5987 1129 6051 1193
rect 6180 1132 6244 1196
rect 6310 1132 6374 1196
rect 4466 962 4530 1026
rect 4596 962 4660 1026
rect 5537 468 5601 532
rect 5667 468 5731 532
rect 5859 467 5923 531
rect 5989 467 6053 531
rect 6501 463 6565 527
rect 6631 463 6695 527
rect 7141 471 7205 535
rect 7271 471 7335 535
rect 5857 140 5921 204
rect 5987 140 6051 204
rect 6178 129 6242 193
rect 6308 129 6372 193
rect 6500 142 6564 206
rect 6630 142 6694 206
rect 7140 138 7204 202
rect 7270 138 7334 202
rect 6179 -518 6243 -454
rect 6309 -518 6373 -454
rect 6820 -525 6884 -461
rect 6950 -525 7014 -461
rect 7140 -514 7204 -450
rect 7270 -514 7334 -450
<< metal2 >>
rect 9098 15380 10796 15480
rect 7438 15301 7657 15313
rect 7438 15237 7451 15301
rect 7515 15237 7581 15301
rect 7645 15237 7657 15301
rect 7438 15225 7657 15237
rect 8397 15301 8616 15313
rect 8397 15237 8409 15301
rect 8473 15237 8539 15301
rect 8603 15237 8616 15301
rect 8397 15225 8616 15237
rect 9098 14977 9198 15380
rect 10696 14977 10796 15380
rect 11278 15301 11497 15313
rect 11278 15237 11291 15301
rect 11355 15237 11421 15301
rect 11485 15237 11497 15301
rect 11278 15225 11497 15237
rect 12237 15301 12456 15313
rect 12237 15237 12249 15301
rect 12313 15237 12379 15301
rect 12443 15237 12456 15301
rect 12237 15225 12456 15237
rect 12938 15148 13038 15480
rect 12938 15048 14003 15148
rect 12938 14977 13038 15048
rect 6158 14964 6377 14976
rect 5667 14920 5755 14932
rect 5667 14856 5679 14920
rect 5743 14856 5755 14920
rect 6158 14900 6171 14964
rect 6235 14900 6301 14964
rect 6365 14900 6377 14964
rect 6158 14888 6377 14900
rect 6475 14962 6694 14974
rect 6475 14898 6488 14962
rect 6552 14898 6618 14962
rect 6682 14898 6694 14962
rect 5667 14790 5755 14856
rect 5667 14726 5679 14790
rect 5743 14726 5755 14790
rect 5667 13293 5755 14726
rect 6202 14490 6302 14888
rect 6475 14886 6694 14898
rect 9037 14965 9256 14977
rect 9037 14901 9049 14965
rect 9113 14901 9179 14965
rect 9243 14901 9256 14965
rect 9037 14889 9256 14901
rect 9360 14962 9579 14974
rect 9360 14898 9372 14962
rect 9436 14898 9502 14962
rect 9566 14898 9579 14962
rect 9360 14886 9579 14898
rect 9677 14964 9896 14976
rect 9677 14900 9689 14964
rect 9753 14900 9819 14964
rect 9883 14900 9896 14964
rect 9677 14888 9896 14900
rect 9998 14964 10217 14976
rect 9998 14900 10011 14964
rect 10075 14900 10141 14964
rect 10205 14900 10217 14964
rect 9998 14888 10217 14900
rect 10315 14962 10534 14974
rect 10315 14898 10328 14962
rect 10392 14898 10458 14962
rect 10522 14898 10534 14962
rect 6202 14390 6934 14490
rect 6155 14309 6374 14321
rect 6155 14245 6168 14309
rect 6232 14245 6298 14309
rect 6362 14245 6374 14309
rect 6155 14233 6374 14245
rect 6477 14308 6696 14320
rect 6477 14244 6490 14308
rect 6554 14244 6620 14308
rect 6684 14244 6696 14308
rect 6216 13839 6316 14233
rect 6477 14232 6696 14244
rect 6834 14150 6934 14390
rect 7173 14395 7586 14495
rect 7173 14316 7273 14395
rect 7119 14304 7338 14316
rect 7119 14240 7132 14304
rect 7196 14240 7262 14304
rect 7326 14240 7338 14304
rect 7119 14228 7338 14240
rect 6533 14050 6934 14150
rect 7486 14154 7586 14395
rect 8468 14395 8881 14495
rect 9752 14490 9852 14888
rect 7759 14312 7978 14324
rect 7759 14248 7772 14312
rect 7836 14248 7902 14312
rect 7966 14248 7978 14312
rect 7759 14236 7978 14248
rect 8076 14312 8295 14324
rect 8076 14248 8088 14312
rect 8152 14248 8218 14312
rect 8282 14248 8295 14312
rect 8076 14236 8295 14248
rect 8468 14154 8568 14395
rect 8781 14316 8881 14395
rect 9120 14390 9852 14490
rect 10042 14490 10142 14888
rect 10315 14886 10534 14898
rect 10638 14965 10857 14977
rect 10638 14901 10651 14965
rect 10715 14901 10781 14965
rect 10845 14901 10857 14965
rect 10638 14889 10857 14901
rect 12877 14965 13096 14977
rect 12877 14901 12889 14965
rect 12953 14901 13019 14965
rect 13083 14901 13096 14965
rect 12877 14889 13096 14901
rect 13200 14962 13419 14974
rect 13200 14898 13212 14962
rect 13276 14898 13342 14962
rect 13406 14898 13419 14962
rect 13200 14886 13419 14898
rect 13517 14964 13736 14976
rect 13517 14900 13529 14964
rect 13593 14900 13659 14964
rect 13723 14900 13736 14964
rect 13517 14888 13736 14900
rect 10042 14390 10774 14490
rect 8716 14304 8935 14316
rect 8716 14240 8728 14304
rect 8792 14240 8858 14304
rect 8922 14240 8935 14304
rect 8716 14228 8935 14240
rect 7486 14054 7913 14154
rect 6533 14001 6694 14050
rect 6475 13989 6694 14001
rect 7118 13991 7337 14003
rect 6475 13925 6488 13989
rect 6552 13925 6618 13989
rect 6682 13925 6694 13989
rect 6475 13913 6694 13925
rect 6796 13978 7015 13990
rect 6796 13914 6809 13978
rect 6873 13914 6939 13978
rect 7003 13914 7015 13978
rect 7118 13927 7131 13991
rect 7195 13927 7261 13991
rect 7325 13927 7337 13991
rect 7118 13915 7337 13927
rect 7758 13999 7913 14054
rect 8141 14054 8568 14154
rect 9120 14150 9220 14390
rect 9358 14308 9577 14320
rect 9358 14244 9370 14308
rect 9434 14244 9500 14308
rect 9564 14244 9577 14308
rect 9358 14232 9577 14244
rect 9680 14309 9899 14321
rect 9680 14245 9692 14309
rect 9756 14245 9822 14309
rect 9886 14245 9899 14309
rect 9680 14233 9899 14245
rect 9995 14309 10214 14321
rect 9995 14245 10008 14309
rect 10072 14245 10138 14309
rect 10202 14245 10214 14309
rect 9995 14233 10214 14245
rect 10317 14308 10536 14320
rect 10317 14244 10330 14308
rect 10394 14244 10460 14308
rect 10524 14244 10536 14308
rect 8141 13999 8296 14054
rect 9120 14050 9521 14150
rect 7758 13987 7977 13999
rect 7758 13923 7771 13987
rect 7835 13923 7901 13987
rect 7965 13923 7977 13987
rect 6796 13902 7015 13914
rect 6858 13839 6958 13902
rect 6216 13739 6958 13839
rect 7173 13836 7273 13915
rect 7758 13911 7977 13923
rect 8077 13987 8296 13999
rect 8077 13923 8089 13987
rect 8153 13923 8219 13987
rect 8283 13923 8296 13987
rect 8077 13911 8296 13923
rect 8717 13991 8936 14003
rect 8717 13927 8729 13991
rect 8793 13927 8859 13991
rect 8923 13927 8936 13991
rect 9360 14001 9521 14050
rect 8717 13915 8936 13927
rect 9039 13978 9258 13990
rect 8781 13836 8881 13915
rect 9039 13914 9051 13978
rect 9115 13914 9181 13978
rect 9245 13914 9258 13978
rect 9039 13902 9258 13914
rect 9360 13989 9579 14001
rect 9360 13925 9372 13989
rect 9436 13925 9502 13989
rect 9566 13925 9579 13989
rect 9360 13913 9579 13925
rect 7173 13818 7958 13836
rect 7173 13754 7762 13818
rect 7826 13754 7882 13818
rect 7946 13754 7958 13818
rect 7173 13736 7958 13754
rect 8096 13818 8881 13836
rect 8096 13754 8108 13818
rect 8172 13754 8228 13818
rect 8292 13754 8881 13818
rect 8096 13736 8881 13754
rect 9096 13839 9196 13902
rect 9738 13839 9838 14233
rect 9096 13739 9838 13839
rect 10056 13839 10156 14233
rect 10317 14232 10536 14244
rect 10674 14150 10774 14390
rect 11013 14395 11426 14495
rect 11013 14316 11113 14395
rect 10959 14304 11178 14316
rect 10959 14240 10972 14304
rect 11036 14240 11102 14304
rect 11166 14240 11178 14304
rect 10959 14228 11178 14240
rect 10373 14050 10774 14150
rect 11326 14154 11426 14395
rect 12308 14395 12721 14495
rect 13592 14490 13692 14888
rect 11599 14312 11818 14324
rect 11599 14248 11612 14312
rect 11676 14248 11742 14312
rect 11806 14248 11818 14312
rect 11599 14236 11818 14248
rect 11916 14312 12135 14324
rect 11916 14248 11928 14312
rect 11992 14248 12058 14312
rect 12122 14248 12135 14312
rect 11916 14236 12135 14248
rect 12308 14154 12408 14395
rect 12621 14316 12721 14395
rect 12960 14390 13692 14490
rect 13903 14487 14003 15048
rect 13840 14475 14059 14487
rect 13840 14411 13853 14475
rect 13917 14411 13983 14475
rect 14047 14411 14059 14475
rect 13840 14399 14059 14411
rect 12556 14304 12775 14316
rect 12556 14240 12568 14304
rect 12632 14240 12698 14304
rect 12762 14240 12775 14304
rect 12556 14228 12775 14240
rect 11326 14054 11753 14154
rect 10373 14001 10534 14050
rect 10315 13989 10534 14001
rect 10958 13991 11177 14003
rect 10315 13925 10328 13989
rect 10392 13925 10458 13989
rect 10522 13925 10534 13989
rect 10315 13913 10534 13925
rect 10636 13978 10855 13990
rect 10636 13914 10649 13978
rect 10713 13914 10779 13978
rect 10843 13914 10855 13978
rect 10958 13927 10971 13991
rect 11035 13927 11101 13991
rect 11165 13927 11177 13991
rect 10958 13915 11177 13927
rect 11598 13999 11753 14054
rect 11981 14054 12408 14154
rect 12960 14150 13060 14390
rect 13198 14308 13417 14320
rect 13198 14244 13210 14308
rect 13274 14244 13340 14308
rect 13404 14244 13417 14308
rect 13198 14232 13417 14244
rect 13520 14309 13739 14321
rect 13520 14245 13532 14309
rect 13596 14245 13662 14309
rect 13726 14245 13739 14309
rect 13520 14233 13739 14245
rect 16308 14317 16396 14329
rect 16308 14253 16320 14317
rect 16384 14253 16396 14317
rect 11981 13999 12136 14054
rect 12960 14050 13361 14150
rect 11598 13987 11817 13999
rect 11598 13923 11611 13987
rect 11675 13923 11741 13987
rect 11805 13923 11817 13987
rect 10636 13902 10855 13914
rect 10698 13839 10798 13902
rect 10056 13739 10798 13839
rect 11013 13836 11113 13915
rect 11598 13911 11817 13923
rect 11917 13987 12136 13999
rect 11917 13923 11929 13987
rect 11993 13923 12059 13987
rect 12123 13923 12136 13987
rect 11917 13911 12136 13923
rect 12557 13991 12776 14003
rect 12557 13927 12569 13991
rect 12633 13927 12699 13991
rect 12763 13927 12776 13991
rect 13200 14001 13361 14050
rect 12557 13915 12776 13927
rect 12879 13978 13098 13990
rect 12621 13836 12721 13915
rect 12879 13914 12891 13978
rect 12955 13914 13021 13978
rect 13085 13914 13098 13978
rect 12879 13902 13098 13914
rect 13200 13989 13419 14001
rect 13200 13925 13212 13989
rect 13276 13925 13342 13989
rect 13406 13925 13419 13989
rect 13200 13913 13419 13925
rect 11013 13818 11798 13836
rect 11013 13754 11602 13818
rect 11666 13754 11722 13818
rect 11786 13754 11798 13818
rect 11013 13736 11798 13754
rect 11936 13818 12721 13836
rect 11936 13754 11948 13818
rect 12012 13754 12068 13818
rect 12132 13754 12721 13818
rect 11936 13736 12721 13754
rect 12936 13839 13036 13902
rect 13578 13839 13678 14233
rect 16308 14187 16396 14253
rect 16308 14123 16320 14187
rect 16384 14123 16396 14187
rect 16308 14110 16396 14123
rect 12936 13739 13678 13839
rect 15908 13612 16127 13624
rect 15908 13548 15921 13612
rect 15985 13548 16051 13612
rect 16115 13548 16127 13612
rect 15908 13536 16127 13548
rect 15913 13369 16132 13381
rect 5667 13229 5679 13293
rect 5743 13229 5755 13293
rect 6797 13339 7016 13351
rect 6797 13275 6810 13339
rect 6874 13275 6940 13339
rect 7004 13275 7016 13339
rect 6797 13263 7016 13275
rect 7438 13332 7657 13344
rect 7438 13268 7451 13332
rect 7515 13268 7581 13332
rect 7645 13268 7657 13332
rect 7438 13256 7657 13268
rect 7758 13343 7977 13355
rect 7758 13279 7771 13343
rect 7835 13279 7901 13343
rect 7965 13279 7977 13343
rect 7758 13267 7977 13279
rect 8077 13343 8296 13355
rect 8077 13279 8089 13343
rect 8153 13279 8219 13343
rect 8283 13279 8296 13343
rect 8077 13267 8296 13279
rect 8397 13332 8616 13344
rect 8397 13268 8409 13332
rect 8473 13268 8539 13332
rect 8603 13268 8616 13332
rect 8397 13256 8616 13268
rect 9038 13339 9257 13351
rect 9038 13275 9050 13339
rect 9114 13275 9180 13339
rect 9244 13275 9257 13339
rect 9038 13263 9257 13275
rect 10637 13339 10856 13351
rect 10637 13275 10650 13339
rect 10714 13275 10780 13339
rect 10844 13275 10856 13339
rect 10637 13263 10856 13275
rect 11278 13332 11497 13344
rect 11278 13268 11291 13332
rect 11355 13268 11421 13332
rect 11485 13268 11497 13332
rect 11278 13256 11497 13268
rect 11598 13343 11817 13355
rect 11598 13279 11611 13343
rect 11675 13279 11741 13343
rect 11805 13279 11817 13343
rect 11598 13267 11817 13279
rect 11917 13343 12136 13355
rect 11917 13279 11929 13343
rect 11993 13279 12059 13343
rect 12123 13279 12136 13343
rect 11917 13267 12136 13279
rect 12237 13332 12456 13344
rect 12237 13268 12249 13332
rect 12313 13268 12379 13332
rect 12443 13268 12456 13332
rect 12237 13256 12456 13268
rect 12878 13339 13097 13351
rect 12878 13275 12890 13339
rect 12954 13275 13020 13339
rect 13084 13275 13097 13339
rect 15913 13305 15926 13369
rect 15990 13305 16056 13369
rect 16120 13305 16132 13369
rect 15913 13293 16132 13305
rect 12878 13263 13097 13275
rect 5667 13163 5755 13229
rect 5667 13099 5679 13163
rect 5743 13099 5755 13163
rect 5667 13086 5755 13099
rect 7073 10418 7173 10921
rect 9483 10821 11349 10921
rect 7655 10742 7874 10754
rect 7655 10678 7668 10742
rect 7732 10678 7798 10742
rect 7862 10678 7874 10742
rect 7655 10666 7874 10678
rect 8782 10742 9001 10754
rect 8782 10678 8794 10742
rect 8858 10678 8924 10742
rect 8988 10678 9001 10742
rect 8782 10666 9001 10678
rect 9483 10418 9583 10821
rect 11249 10418 11349 10821
rect 11831 10742 12050 10754
rect 11831 10678 11844 10742
rect 11908 10678 11974 10742
rect 12038 10678 12050 10742
rect 11831 10666 12050 10678
rect 12958 10742 13177 10754
rect 12958 10678 12970 10742
rect 13034 10678 13100 10742
rect 13164 10678 13177 10742
rect 12958 10666 13177 10678
rect 13659 10418 13759 10921
rect 6375 10405 6594 10417
rect 6375 10341 6388 10405
rect 6452 10341 6518 10405
rect 6582 10341 6594 10405
rect 6375 10329 6594 10341
rect 6692 10403 6911 10415
rect 6692 10339 6705 10403
rect 6769 10339 6835 10403
rect 6899 10339 6911 10403
rect 6419 9931 6519 10329
rect 6692 10327 6911 10339
rect 7015 10406 7234 10418
rect 7015 10342 7028 10406
rect 7092 10342 7158 10406
rect 7222 10342 7234 10406
rect 7015 10330 7234 10342
rect 9422 10406 9641 10418
rect 9422 10342 9434 10406
rect 9498 10342 9564 10406
rect 9628 10342 9641 10406
rect 9422 10330 9641 10342
rect 9745 10403 9964 10415
rect 9745 10339 9757 10403
rect 9821 10339 9887 10403
rect 9951 10339 9964 10403
rect 9745 10327 9964 10339
rect 10062 10405 10281 10417
rect 10062 10341 10074 10405
rect 10138 10341 10204 10405
rect 10268 10341 10281 10405
rect 10062 10329 10281 10341
rect 10551 10405 10770 10417
rect 10551 10341 10564 10405
rect 10628 10341 10694 10405
rect 10758 10341 10770 10405
rect 10551 10329 10770 10341
rect 10868 10403 11087 10415
rect 10868 10339 10881 10403
rect 10945 10339 11011 10403
rect 11075 10339 11087 10403
rect 6419 9831 7151 9931
rect 6372 9750 6591 9762
rect 6372 9686 6385 9750
rect 6449 9686 6515 9750
rect 6579 9686 6591 9750
rect 6372 9674 6591 9686
rect 6694 9749 6913 9761
rect 6694 9685 6707 9749
rect 6771 9685 6837 9749
rect 6901 9685 6913 9749
rect 6433 9280 6533 9674
rect 6694 9673 6913 9685
rect 7051 9591 7151 9831
rect 7390 9836 7803 9936
rect 7390 9757 7490 9836
rect 7336 9745 7555 9757
rect 7336 9681 7349 9745
rect 7413 9681 7479 9745
rect 7543 9681 7555 9745
rect 7336 9669 7555 9681
rect 6750 9491 7151 9591
rect 7703 9595 7803 9836
rect 8853 9836 9266 9936
rect 10137 9931 10237 10329
rect 7976 9753 8195 9765
rect 7976 9689 7989 9753
rect 8053 9689 8119 9753
rect 8183 9689 8195 9753
rect 7976 9677 8195 9689
rect 8461 9753 8680 9765
rect 8461 9689 8473 9753
rect 8537 9689 8603 9753
rect 8667 9689 8680 9753
rect 8461 9677 8680 9689
rect 8853 9595 8953 9836
rect 9166 9757 9266 9836
rect 9505 9831 10237 9931
rect 10595 9931 10695 10329
rect 10868 10327 11087 10339
rect 11191 10406 11410 10418
rect 11191 10342 11204 10406
rect 11268 10342 11334 10406
rect 11398 10342 11410 10406
rect 11191 10330 11410 10342
rect 13598 10406 13817 10418
rect 13598 10342 13610 10406
rect 13674 10342 13740 10406
rect 13804 10342 13817 10406
rect 13598 10330 13817 10342
rect 13921 10403 14140 10415
rect 13921 10339 13933 10403
rect 13997 10339 14063 10403
rect 14127 10339 14140 10403
rect 13921 10327 14140 10339
rect 14238 10405 14457 10417
rect 14238 10341 14250 10405
rect 14314 10341 14380 10405
rect 14444 10341 14457 10405
rect 14238 10329 14457 10341
rect 10595 9831 11327 9931
rect 9101 9745 9320 9757
rect 9101 9681 9113 9745
rect 9177 9681 9243 9745
rect 9307 9681 9320 9745
rect 9101 9669 9320 9681
rect 7703 9495 8130 9595
rect 6750 9442 6911 9491
rect 6692 9430 6911 9442
rect 7335 9432 7554 9444
rect 6692 9366 6705 9430
rect 6769 9366 6835 9430
rect 6899 9366 6911 9430
rect 6692 9354 6911 9366
rect 7013 9419 7232 9431
rect 7013 9355 7026 9419
rect 7090 9355 7156 9419
rect 7220 9355 7232 9419
rect 7335 9368 7348 9432
rect 7412 9368 7478 9432
rect 7542 9368 7554 9432
rect 7335 9356 7554 9368
rect 7975 9440 8130 9495
rect 8526 9495 8953 9595
rect 9505 9591 9605 9831
rect 9743 9749 9962 9761
rect 9743 9685 9755 9749
rect 9819 9685 9885 9749
rect 9949 9685 9962 9749
rect 9743 9673 9962 9685
rect 10065 9750 10284 9762
rect 10065 9686 10077 9750
rect 10141 9686 10207 9750
rect 10271 9686 10284 9750
rect 10065 9674 10284 9686
rect 10548 9750 10767 9762
rect 10548 9686 10561 9750
rect 10625 9686 10691 9750
rect 10755 9686 10767 9750
rect 10548 9674 10767 9686
rect 10870 9749 11089 9761
rect 10870 9685 10883 9749
rect 10947 9685 11013 9749
rect 11077 9685 11089 9749
rect 8526 9440 8681 9495
rect 9505 9491 9906 9591
rect 7975 9428 8194 9440
rect 7975 9364 7988 9428
rect 8052 9364 8118 9428
rect 8182 9364 8194 9428
rect 7013 9343 7232 9355
rect 7075 9280 7175 9343
rect 6433 9180 7175 9280
rect 7390 9277 7490 9356
rect 7975 9352 8194 9364
rect 8462 9428 8681 9440
rect 8462 9364 8474 9428
rect 8538 9364 8604 9428
rect 8668 9364 8681 9428
rect 8462 9352 8681 9364
rect 9102 9432 9321 9444
rect 9102 9368 9114 9432
rect 9178 9368 9244 9432
rect 9308 9368 9321 9432
rect 9745 9442 9906 9491
rect 9102 9356 9321 9368
rect 9424 9419 9643 9431
rect 9166 9277 9266 9356
rect 9424 9355 9436 9419
rect 9500 9355 9566 9419
rect 9630 9355 9643 9419
rect 9424 9343 9643 9355
rect 9745 9430 9964 9442
rect 9745 9366 9757 9430
rect 9821 9366 9887 9430
rect 9951 9366 9964 9430
rect 9745 9354 9964 9366
rect 7390 9259 8175 9277
rect 7390 9195 7979 9259
rect 8043 9195 8099 9259
rect 8163 9195 8175 9259
rect 7390 9177 8175 9195
rect 8481 9259 9266 9277
rect 8481 9195 8493 9259
rect 8557 9195 8613 9259
rect 8677 9195 9266 9259
rect 8481 9177 9266 9195
rect 9481 9280 9581 9343
rect 10123 9280 10223 9674
rect 9481 9180 10223 9280
rect 10609 9280 10709 9674
rect 10870 9673 11089 9685
rect 11227 9591 11327 9831
rect 11566 9836 11979 9936
rect 11566 9757 11666 9836
rect 11512 9745 11731 9757
rect 11512 9681 11525 9745
rect 11589 9681 11655 9745
rect 11719 9681 11731 9745
rect 11512 9669 11731 9681
rect 10926 9491 11327 9591
rect 11879 9595 11979 9836
rect 13029 9836 13442 9936
rect 14313 9931 14413 10329
rect 12152 9753 12371 9765
rect 12152 9689 12165 9753
rect 12229 9689 12295 9753
rect 12359 9689 12371 9753
rect 12152 9677 12371 9689
rect 12637 9753 12856 9765
rect 12637 9689 12649 9753
rect 12713 9689 12779 9753
rect 12843 9689 12856 9753
rect 12637 9677 12856 9689
rect 13029 9595 13129 9836
rect 13342 9757 13442 9836
rect 13681 9831 14413 9931
rect 13277 9745 13496 9757
rect 13277 9681 13289 9745
rect 13353 9681 13419 9745
rect 13483 9681 13496 9745
rect 13277 9669 13496 9681
rect 11879 9495 12306 9595
rect 10926 9442 11087 9491
rect 10868 9430 11087 9442
rect 11511 9432 11730 9444
rect 10868 9366 10881 9430
rect 10945 9366 11011 9430
rect 11075 9366 11087 9430
rect 10868 9354 11087 9366
rect 11189 9419 11408 9431
rect 11189 9355 11202 9419
rect 11266 9355 11332 9419
rect 11396 9355 11408 9419
rect 11511 9368 11524 9432
rect 11588 9368 11654 9432
rect 11718 9368 11730 9432
rect 11511 9356 11730 9368
rect 12151 9440 12306 9495
rect 12702 9495 13129 9595
rect 13681 9591 13781 9831
rect 13919 9749 14138 9761
rect 13919 9685 13931 9749
rect 13995 9685 14061 9749
rect 14125 9685 14138 9749
rect 13919 9673 14138 9685
rect 14241 9750 14460 9762
rect 14241 9686 14253 9750
rect 14317 9686 14383 9750
rect 14447 9686 14460 9750
rect 14241 9674 14460 9686
rect 12702 9440 12857 9495
rect 13681 9491 14082 9591
rect 12151 9428 12370 9440
rect 12151 9364 12164 9428
rect 12228 9364 12294 9428
rect 12358 9364 12370 9428
rect 11189 9343 11408 9355
rect 11251 9280 11351 9343
rect 10609 9180 11351 9280
rect 11566 9277 11666 9356
rect 12151 9352 12370 9364
rect 12638 9428 12857 9440
rect 12638 9364 12650 9428
rect 12714 9364 12780 9428
rect 12844 9364 12857 9428
rect 12638 9352 12857 9364
rect 13278 9432 13497 9444
rect 13278 9368 13290 9432
rect 13354 9368 13420 9432
rect 13484 9368 13497 9432
rect 13921 9442 14082 9491
rect 13278 9356 13497 9368
rect 13600 9419 13819 9431
rect 13342 9277 13442 9356
rect 13600 9355 13612 9419
rect 13676 9355 13742 9419
rect 13806 9355 13819 9419
rect 13600 9343 13819 9355
rect 13921 9430 14140 9442
rect 13921 9366 13933 9430
rect 13997 9366 14063 9430
rect 14127 9366 14140 9430
rect 13921 9354 14140 9366
rect 11566 9259 12351 9277
rect 11566 9195 12155 9259
rect 12219 9195 12275 9259
rect 12339 9195 12351 9259
rect 11566 9177 12351 9195
rect 12657 9259 13442 9277
rect 12657 9195 12669 9259
rect 12733 9195 12789 9259
rect 12853 9195 13442 9259
rect 12657 9177 13442 9195
rect 13657 9280 13757 9343
rect 14299 9280 14399 9674
rect 13657 9180 14399 9280
rect 7014 8780 7233 8792
rect 7014 8716 7027 8780
rect 7091 8716 7157 8780
rect 7221 8716 7233 8780
rect 7014 8704 7233 8716
rect 7655 8773 7874 8785
rect 7655 8709 7668 8773
rect 7732 8709 7798 8773
rect 7862 8709 7874 8773
rect 7655 8697 7874 8709
rect 7975 8784 8194 8796
rect 7975 8720 7988 8784
rect 8052 8720 8118 8784
rect 8182 8720 8194 8784
rect 7975 8708 8194 8720
rect 8462 8784 8681 8796
rect 8462 8720 8474 8784
rect 8538 8720 8604 8784
rect 8668 8720 8681 8784
rect 8462 8708 8681 8720
rect 8782 8773 9001 8785
rect 8782 8709 8794 8773
rect 8858 8709 8924 8773
rect 8988 8709 9001 8773
rect 8782 8697 9001 8709
rect 9423 8780 9642 8792
rect 9423 8716 9435 8780
rect 9499 8716 9565 8780
rect 9629 8716 9642 8780
rect 9423 8704 9642 8716
rect 11190 8780 11409 8792
rect 11190 8716 11203 8780
rect 11267 8716 11333 8780
rect 11397 8716 11409 8780
rect 11190 8704 11409 8716
rect 11831 8773 12050 8785
rect 11831 8709 11844 8773
rect 11908 8709 11974 8773
rect 12038 8709 12050 8773
rect 11831 8697 12050 8709
rect 12151 8784 12370 8796
rect 12151 8720 12164 8784
rect 12228 8720 12294 8784
rect 12358 8720 12370 8784
rect 12151 8708 12370 8720
rect 12638 8784 12857 8796
rect 12638 8720 12650 8784
rect 12714 8720 12780 8784
rect 12844 8720 12857 8784
rect 12638 8708 12857 8720
rect 12958 8773 13177 8785
rect 12958 8709 12970 8773
rect 13034 8709 13100 8773
rect 13164 8709 13177 8773
rect 12958 8697 13177 8709
rect 13599 8780 13818 8792
rect 13599 8716 13611 8780
rect 13675 8716 13741 8780
rect 13805 8716 13818 8780
rect 13599 8704 13818 8716
rect 4448 1269 4667 1281
rect 4448 1205 4461 1269
rect 4525 1205 4591 1269
rect 4655 1205 4667 1269
rect 6225 1208 6325 1711
rect 6807 1532 7026 1544
rect 6807 1468 6820 1532
rect 6884 1468 6950 1532
rect 7014 1468 7026 1532
rect 6807 1456 7026 1468
rect 4448 1193 4667 1205
rect 5527 1195 5746 1207
rect 5527 1131 5540 1195
rect 5604 1131 5670 1195
rect 5734 1131 5746 1195
rect 5527 1119 5746 1131
rect 5844 1193 6063 1205
rect 5844 1129 5857 1193
rect 5921 1129 5987 1193
rect 6051 1129 6063 1193
rect 4453 1026 4672 1038
rect 4453 962 4466 1026
rect 4530 962 4596 1026
rect 4660 962 4672 1026
rect 4453 950 4672 962
rect 5571 713 5671 1119
rect 5844 1117 6063 1129
rect 6167 1196 6386 1208
rect 6167 1132 6180 1196
rect 6244 1132 6310 1196
rect 6374 1132 6386 1196
rect 6167 1120 6386 1132
rect 5571 613 6303 713
rect 5524 532 5743 544
rect 5524 468 5537 532
rect 5601 468 5667 532
rect 5731 468 5743 532
rect 5524 456 5743 468
rect 5846 531 6065 543
rect 5846 467 5859 531
rect 5923 467 5989 531
rect 6053 467 6065 531
rect 5585 54 5685 456
rect 5846 455 6065 467
rect 6203 373 6303 613
rect 6542 618 6955 718
rect 6542 539 6642 618
rect 6488 527 6707 539
rect 6488 463 6501 527
rect 6565 463 6631 527
rect 6695 463 6707 527
rect 6488 451 6707 463
rect 5902 273 6303 373
rect 6855 377 6955 618
rect 7128 535 7347 547
rect 7128 471 7141 535
rect 7205 471 7271 535
rect 7335 471 7347 535
rect 7128 459 7347 471
rect 6855 277 7282 377
rect 5902 216 6002 273
rect 5844 204 6063 216
rect 6487 206 6706 218
rect 7182 214 7282 277
rect 5844 140 5857 204
rect 5921 140 5987 204
rect 6051 140 6063 204
rect 5844 128 6063 140
rect 6165 193 6384 205
rect 6165 129 6178 193
rect 6242 129 6308 193
rect 6372 129 6384 193
rect 6487 142 6500 206
rect 6564 142 6630 206
rect 6694 142 6706 206
rect 6487 130 6706 142
rect 7127 202 7346 214
rect 7127 138 7140 202
rect 7204 138 7270 202
rect 7334 138 7346 202
rect 6165 117 6384 129
rect 6227 54 6327 117
rect 5585 -46 6327 54
rect 6542 51 6642 130
rect 7127 126 7346 138
rect 6542 33 7327 51
rect 6542 -31 7131 33
rect 7195 -31 7251 33
rect 7315 -31 7327 33
rect 6542 -49 7327 -31
rect 6166 -454 6385 -442
rect 6166 -518 6179 -454
rect 6243 -518 6309 -454
rect 6373 -518 6385 -454
rect 6166 -530 6385 -518
rect 6807 -461 7026 -449
rect 6807 -525 6820 -461
rect 6884 -525 6950 -461
rect 7014 -525 7026 -461
rect 6807 -537 7026 -525
rect 7127 -450 7346 -438
rect 7127 -514 7140 -450
rect 7204 -514 7270 -450
rect 7334 -514 7346 -450
rect 7127 -526 7346 -514
<< via2 >>
rect 7451 15237 7515 15301
rect 7581 15237 7645 15301
rect 8409 15237 8473 15301
rect 8539 15237 8603 15301
rect 11291 15237 11355 15301
rect 11421 15237 11485 15301
rect 12249 15237 12313 15301
rect 12379 15237 12443 15301
rect 6488 14898 6552 14962
rect 6618 14898 6682 14962
rect 9372 14898 9436 14962
rect 9502 14898 9566 14962
rect 10328 14898 10392 14962
rect 10458 14898 10522 14962
rect 6490 14244 6554 14308
rect 6620 14244 6684 14308
rect 7772 14248 7836 14312
rect 7902 14248 7966 14312
rect 8088 14248 8152 14312
rect 8218 14248 8282 14312
rect 13212 14898 13276 14962
rect 13342 14898 13406 14962
rect 9370 14244 9434 14308
rect 9500 14244 9564 14308
rect 10330 14244 10394 14308
rect 10460 14244 10524 14308
rect 7762 13754 7826 13818
rect 7882 13754 7946 13818
rect 8108 13754 8172 13818
rect 8228 13754 8292 13818
rect 11612 14248 11676 14312
rect 11742 14248 11806 14312
rect 11928 14248 11992 14312
rect 12058 14248 12122 14312
rect 13210 14244 13274 14308
rect 13340 14244 13404 14308
rect 11602 13754 11666 13818
rect 11722 13754 11786 13818
rect 11948 13754 12012 13818
rect 12068 13754 12132 13818
rect 6810 13275 6874 13339
rect 6940 13275 7004 13339
rect 7451 13268 7515 13332
rect 7581 13268 7645 13332
rect 7771 13279 7835 13343
rect 7901 13279 7965 13343
rect 8089 13279 8153 13343
rect 8219 13279 8283 13343
rect 8409 13268 8473 13332
rect 8539 13268 8603 13332
rect 9050 13275 9114 13339
rect 9180 13275 9244 13339
rect 10650 13275 10714 13339
rect 10780 13275 10844 13339
rect 11291 13268 11355 13332
rect 11421 13268 11485 13332
rect 11611 13279 11675 13343
rect 11741 13279 11805 13343
rect 11929 13279 11993 13343
rect 12059 13279 12123 13343
rect 12249 13268 12313 13332
rect 12379 13268 12443 13332
rect 12890 13275 12954 13339
rect 13020 13275 13084 13339
rect 15926 13305 15990 13369
rect 16056 13305 16120 13369
rect 7668 10678 7732 10742
rect 7798 10678 7862 10742
rect 8794 10678 8858 10742
rect 8924 10678 8988 10742
rect 11844 10678 11908 10742
rect 11974 10678 12038 10742
rect 12970 10678 13034 10742
rect 13100 10678 13164 10742
rect 6705 10339 6769 10403
rect 6835 10339 6899 10403
rect 9757 10339 9821 10403
rect 9887 10339 9951 10403
rect 10881 10339 10945 10403
rect 11011 10339 11075 10403
rect 6707 9685 6771 9749
rect 6837 9685 6901 9749
rect 7989 9689 8053 9753
rect 8119 9689 8183 9753
rect 8473 9689 8537 9753
rect 8603 9689 8667 9753
rect 13933 10339 13997 10403
rect 14063 10339 14127 10403
rect 9755 9685 9819 9749
rect 9885 9685 9949 9749
rect 10883 9685 10947 9749
rect 11013 9685 11077 9749
rect 7979 9195 8043 9259
rect 8099 9195 8163 9259
rect 8493 9195 8557 9259
rect 8613 9195 8677 9259
rect 12165 9689 12229 9753
rect 12295 9689 12359 9753
rect 12649 9689 12713 9753
rect 12779 9689 12843 9753
rect 13931 9685 13995 9749
rect 14061 9685 14125 9749
rect 12155 9195 12219 9259
rect 12275 9195 12339 9259
rect 12669 9195 12733 9259
rect 12789 9195 12853 9259
rect 7027 8716 7091 8780
rect 7157 8716 7221 8780
rect 7668 8709 7732 8773
rect 7798 8709 7862 8773
rect 7988 8720 8052 8784
rect 8118 8720 8182 8784
rect 8474 8720 8538 8784
rect 8604 8720 8668 8784
rect 8794 8709 8858 8773
rect 8924 8709 8988 8773
rect 9435 8716 9499 8780
rect 9565 8716 9629 8780
rect 11203 8716 11267 8780
rect 11333 8716 11397 8780
rect 11844 8709 11908 8773
rect 11974 8709 12038 8773
rect 12164 8720 12228 8784
rect 12294 8720 12358 8784
rect 12650 8720 12714 8784
rect 12780 8720 12844 8784
rect 12970 8709 13034 8773
rect 13100 8709 13164 8773
rect 13611 8716 13675 8780
rect 13741 8716 13805 8780
rect 6820 1468 6884 1532
rect 6950 1468 7014 1532
rect 5857 1129 5921 1193
rect 5987 1129 6051 1193
rect 4466 962 4530 1026
rect 4596 962 4660 1026
rect 5859 467 5923 531
rect 5989 467 6053 531
rect 7141 471 7205 535
rect 7271 471 7335 535
rect 7131 -31 7195 33
rect 7251 -31 7315 33
rect 6179 -518 6243 -454
rect 6309 -518 6373 -454
rect 6820 -525 6884 -461
rect 6950 -525 7014 -461
rect 7140 -514 7204 -450
rect 7270 -514 7334 -450
<< metal3 >>
rect 7438 15301 7657 15313
rect 7438 15237 7451 15301
rect 7515 15237 7581 15301
rect 7645 15237 7657 15301
rect 7438 15225 7657 15237
rect 8397 15301 8616 15313
rect 8397 15237 8409 15301
rect 8473 15237 8539 15301
rect 8603 15237 8616 15301
rect 8397 15225 8616 15237
rect 11278 15301 11497 15313
rect 11278 15237 11291 15301
rect 11355 15237 11421 15301
rect 11485 15237 11497 15301
rect 11278 15225 11497 15237
rect 12237 15301 12456 15313
rect 12237 15237 12249 15301
rect 12313 15237 12379 15301
rect 12443 15237 12456 15301
rect 12237 15225 12456 15237
rect 6475 14962 6694 14974
rect 6475 14898 6488 14962
rect 6552 14898 6618 14962
rect 6682 14898 6694 14962
rect 6475 14886 6694 14898
rect 6515 14806 6615 14886
rect 6515 14706 7275 14806
rect 6477 14308 6696 14320
rect 6477 14244 6490 14308
rect 6554 14244 6620 14308
rect 6684 14244 6696 14308
rect 6477 14232 6696 14244
rect 6533 14171 6633 14232
rect 6533 14071 6956 14171
rect 6856 13351 6956 14071
rect 6797 13339 7016 13351
rect 6797 13275 6810 13339
rect 6874 13275 6940 13339
rect 7004 13275 7016 13339
rect 6797 13263 7016 13275
rect 7175 13199 7275 14706
rect 7494 13344 7594 15225
rect 7759 14312 7978 14324
rect 7759 14248 7772 14312
rect 7836 14248 7902 14312
rect 7966 14248 7978 14312
rect 7759 14236 7978 14248
rect 8076 14312 8295 14324
rect 8076 14248 8088 14312
rect 8152 14248 8218 14312
rect 8282 14248 8295 14312
rect 8076 14236 8295 14248
rect 7808 13836 7908 14236
rect 8146 13836 8246 14236
rect 7749 13818 7958 13836
rect 7749 13754 7762 13818
rect 7826 13754 7882 13818
rect 7946 13754 7958 13818
rect 7749 13736 7958 13754
rect 8096 13818 8305 13836
rect 8096 13754 8108 13818
rect 8172 13754 8228 13818
rect 8292 13754 8305 13818
rect 8096 13736 8305 13754
rect 7438 13332 7657 13344
rect 7438 13268 7451 13332
rect 7515 13268 7581 13332
rect 7645 13268 7657 13332
rect 7438 13256 7657 13268
rect 7758 13343 7977 13355
rect 7758 13279 7771 13343
rect 7835 13279 7901 13343
rect 7965 13279 7977 13343
rect 7758 13267 7977 13279
rect 8077 13343 8296 13355
rect 8460 13344 8560 15225
rect 9360 14962 9579 14974
rect 9360 14898 9372 14962
rect 9436 14898 9502 14962
rect 9566 14898 9579 14962
rect 9360 14886 9579 14898
rect 10315 14962 10534 14974
rect 10315 14898 10328 14962
rect 10392 14898 10458 14962
rect 10522 14898 10534 14962
rect 10315 14886 10534 14898
rect 9439 14806 9539 14886
rect 8779 14706 9539 14806
rect 10355 14806 10455 14886
rect 10355 14706 11115 14806
rect 8077 13279 8089 13343
rect 8153 13279 8219 13343
rect 8283 13279 8296 13343
rect 8077 13267 8296 13279
rect 8397 13332 8616 13344
rect 8397 13268 8409 13332
rect 8473 13268 8539 13332
rect 8603 13268 8616 13332
rect 7806 13199 7906 13267
rect 7175 13099 7906 13199
rect 8148 13199 8248 13267
rect 8397 13256 8616 13268
rect 8779 13199 8879 14706
rect 9358 14308 9577 14320
rect 9358 14244 9370 14308
rect 9434 14244 9500 14308
rect 9564 14244 9577 14308
rect 9358 14232 9577 14244
rect 10317 14308 10536 14320
rect 10317 14244 10330 14308
rect 10394 14244 10460 14308
rect 10524 14244 10536 14308
rect 10317 14232 10536 14244
rect 9421 14171 9521 14232
rect 9098 14071 9521 14171
rect 10373 14171 10473 14232
rect 10373 14071 10796 14171
rect 9098 13351 9198 14071
rect 10696 13351 10796 14071
rect 9038 13339 9257 13351
rect 9038 13275 9050 13339
rect 9114 13275 9180 13339
rect 9244 13275 9257 13339
rect 9038 13263 9257 13275
rect 10637 13339 10856 13351
rect 10637 13275 10650 13339
rect 10714 13275 10780 13339
rect 10844 13275 10856 13339
rect 10637 13263 10856 13275
rect 8148 13099 8879 13199
rect 11015 13199 11115 14706
rect 11334 13344 11434 15225
rect 11599 14312 11818 14324
rect 11599 14248 11612 14312
rect 11676 14248 11742 14312
rect 11806 14248 11818 14312
rect 11599 14236 11818 14248
rect 11916 14312 12135 14324
rect 11916 14248 11928 14312
rect 11992 14248 12058 14312
rect 12122 14248 12135 14312
rect 11916 14236 12135 14248
rect 11648 13836 11748 14236
rect 11986 13836 12086 14236
rect 11589 13818 11798 13836
rect 11589 13754 11602 13818
rect 11666 13754 11722 13818
rect 11786 13754 11798 13818
rect 11589 13736 11798 13754
rect 11936 13818 12145 13836
rect 11936 13754 11948 13818
rect 12012 13754 12068 13818
rect 12132 13754 12145 13818
rect 11936 13736 12145 13754
rect 11278 13332 11497 13344
rect 11278 13268 11291 13332
rect 11355 13268 11421 13332
rect 11485 13268 11497 13332
rect 11278 13256 11497 13268
rect 11598 13343 11817 13355
rect 11598 13279 11611 13343
rect 11675 13279 11741 13343
rect 11805 13279 11817 13343
rect 11598 13267 11817 13279
rect 11917 13343 12136 13355
rect 12300 13344 12400 15225
rect 13200 14962 13419 14974
rect 13200 14898 13212 14962
rect 13276 14898 13342 14962
rect 13406 14898 13419 14962
rect 13200 14886 13419 14898
rect 13279 14806 13379 14886
rect 12619 14706 13379 14806
rect 11917 13279 11929 13343
rect 11993 13279 12059 13343
rect 12123 13279 12136 13343
rect 11917 13267 12136 13279
rect 12237 13332 12456 13344
rect 12237 13268 12249 13332
rect 12313 13268 12379 13332
rect 12443 13268 12456 13332
rect 11646 13199 11746 13267
rect 11015 13099 11746 13199
rect 11988 13199 12088 13267
rect 12237 13256 12456 13268
rect 12619 13199 12719 14706
rect 13198 14308 13417 14320
rect 13198 14244 13210 14308
rect 13274 14244 13340 14308
rect 13404 14244 13417 14308
rect 13198 14232 13417 14244
rect 13261 14171 13361 14232
rect 12938 14071 13361 14171
rect 12938 13351 13038 14071
rect 15913 13369 16132 13381
rect 12878 13339 13097 13351
rect 12878 13275 12890 13339
rect 12954 13275 13020 13339
rect 13084 13275 13097 13339
rect 15913 13305 15926 13369
rect 15990 13305 16056 13369
rect 16120 13305 16132 13369
rect 15913 13293 16132 13305
rect 12878 13263 13097 13275
rect 11988 13099 12719 13199
rect 7655 10742 7874 10754
rect 7655 10678 7668 10742
rect 7732 10678 7798 10742
rect 7862 10678 7874 10742
rect 7655 10666 7874 10678
rect 8782 10742 9001 10754
rect 8782 10678 8794 10742
rect 8858 10678 8924 10742
rect 8988 10678 9001 10742
rect 8782 10666 9001 10678
rect 11831 10742 12050 10754
rect 11831 10678 11844 10742
rect 11908 10678 11974 10742
rect 12038 10678 12050 10742
rect 11831 10666 12050 10678
rect 12958 10742 13177 10754
rect 12958 10678 12970 10742
rect 13034 10678 13100 10742
rect 13164 10678 13177 10742
rect 12958 10666 13177 10678
rect 6692 10403 6911 10415
rect 6692 10339 6705 10403
rect 6769 10339 6835 10403
rect 6899 10339 6911 10403
rect 6692 10327 6911 10339
rect 6732 10247 6832 10327
rect 6732 10147 7492 10247
rect 6694 9749 6913 9761
rect 6694 9685 6707 9749
rect 6771 9685 6837 9749
rect 6901 9685 6913 9749
rect 6694 9673 6913 9685
rect 6750 9612 6850 9673
rect 6750 9512 7173 9612
rect 7073 8792 7173 9512
rect 7014 8780 7233 8792
rect 7014 8716 7027 8780
rect 7091 8716 7157 8780
rect 7221 8716 7233 8780
rect 7014 8704 7233 8716
rect 7392 8640 7492 10147
rect 7711 8785 7811 10666
rect 7976 9753 8195 9765
rect 7976 9689 7989 9753
rect 8053 9689 8119 9753
rect 8183 9689 8195 9753
rect 7976 9677 8195 9689
rect 8461 9753 8680 9765
rect 8461 9689 8473 9753
rect 8537 9689 8603 9753
rect 8667 9689 8680 9753
rect 8461 9677 8680 9689
rect 8025 9277 8125 9677
rect 8531 9277 8631 9677
rect 7966 9259 8175 9277
rect 7966 9195 7979 9259
rect 8043 9195 8099 9259
rect 8163 9195 8175 9259
rect 7966 9177 8175 9195
rect 8481 9259 8690 9277
rect 8481 9195 8493 9259
rect 8557 9195 8613 9259
rect 8677 9195 8690 9259
rect 8481 9177 8690 9195
rect 7655 8773 7874 8785
rect 7655 8709 7668 8773
rect 7732 8709 7798 8773
rect 7862 8709 7874 8773
rect 7655 8697 7874 8709
rect 7975 8784 8194 8796
rect 7975 8720 7988 8784
rect 8052 8720 8118 8784
rect 8182 8720 8194 8784
rect 7975 8708 8194 8720
rect 8462 8784 8681 8796
rect 8845 8785 8945 10666
rect 9745 10403 9964 10415
rect 9745 10339 9757 10403
rect 9821 10339 9887 10403
rect 9951 10339 9964 10403
rect 9745 10327 9964 10339
rect 10868 10403 11087 10415
rect 10868 10339 10881 10403
rect 10945 10339 11011 10403
rect 11075 10339 11087 10403
rect 10868 10327 11087 10339
rect 9824 10247 9924 10327
rect 9164 10147 9924 10247
rect 10908 10247 11008 10327
rect 10908 10147 11668 10247
rect 8462 8720 8474 8784
rect 8538 8720 8604 8784
rect 8668 8720 8681 8784
rect 8462 8708 8681 8720
rect 8782 8773 9001 8785
rect 8782 8709 8794 8773
rect 8858 8709 8924 8773
rect 8988 8709 9001 8773
rect 8023 8640 8123 8708
rect 7392 8540 8123 8640
rect 8533 8640 8633 8708
rect 8782 8697 9001 8709
rect 9164 8640 9264 10147
rect 9743 9749 9962 9761
rect 9743 9685 9755 9749
rect 9819 9685 9885 9749
rect 9949 9685 9962 9749
rect 9743 9673 9962 9685
rect 10870 9749 11089 9761
rect 10870 9685 10883 9749
rect 10947 9685 11013 9749
rect 11077 9685 11089 9749
rect 10870 9673 11089 9685
rect 9806 9612 9906 9673
rect 9483 9512 9906 9612
rect 10926 9612 11026 9673
rect 10926 9512 11349 9612
rect 9483 8792 9583 9512
rect 11249 8792 11349 9512
rect 9423 8780 9642 8792
rect 9423 8716 9435 8780
rect 9499 8716 9565 8780
rect 9629 8716 9642 8780
rect 9423 8704 9642 8716
rect 11190 8780 11409 8792
rect 11190 8716 11203 8780
rect 11267 8716 11333 8780
rect 11397 8716 11409 8780
rect 11190 8704 11409 8716
rect 8533 8540 9264 8640
rect 11568 8640 11668 10147
rect 11887 8785 11987 10666
rect 12152 9753 12371 9765
rect 12152 9689 12165 9753
rect 12229 9689 12295 9753
rect 12359 9689 12371 9753
rect 12152 9677 12371 9689
rect 12637 9753 12856 9765
rect 12637 9689 12649 9753
rect 12713 9689 12779 9753
rect 12843 9689 12856 9753
rect 12637 9677 12856 9689
rect 12201 9277 12301 9677
rect 12707 9277 12807 9677
rect 12142 9259 12351 9277
rect 12142 9195 12155 9259
rect 12219 9195 12275 9259
rect 12339 9195 12351 9259
rect 12142 9177 12351 9195
rect 12657 9259 12866 9277
rect 12657 9195 12669 9259
rect 12733 9195 12789 9259
rect 12853 9195 12866 9259
rect 12657 9177 12866 9195
rect 11831 8773 12050 8785
rect 11831 8709 11844 8773
rect 11908 8709 11974 8773
rect 12038 8709 12050 8773
rect 11831 8697 12050 8709
rect 12151 8784 12370 8796
rect 12151 8720 12164 8784
rect 12228 8720 12294 8784
rect 12358 8720 12370 8784
rect 12151 8708 12370 8720
rect 12638 8784 12857 8796
rect 13021 8785 13121 10666
rect 13921 10403 14140 10415
rect 13921 10339 13933 10403
rect 13997 10339 14063 10403
rect 14127 10339 14140 10403
rect 13921 10327 14140 10339
rect 14000 10247 14100 10327
rect 13340 10147 14100 10247
rect 12638 8720 12650 8784
rect 12714 8720 12780 8784
rect 12844 8720 12857 8784
rect 12638 8708 12857 8720
rect 12958 8773 13177 8785
rect 12958 8709 12970 8773
rect 13034 8709 13100 8773
rect 13164 8709 13177 8773
rect 12199 8640 12299 8708
rect 11568 8540 12299 8640
rect 12709 8640 12809 8708
rect 12958 8697 13177 8709
rect 13340 8640 13440 10147
rect 13919 9749 14138 9761
rect 13919 9685 13931 9749
rect 13995 9685 14061 9749
rect 14125 9685 14138 9749
rect 13919 9673 14138 9685
rect 13982 9612 14082 9673
rect 13659 9512 14082 9612
rect 13659 8792 13759 9512
rect 13599 8780 13818 8792
rect 13599 8716 13611 8780
rect 13675 8716 13741 8780
rect 13805 8716 13818 8780
rect 13599 8704 13818 8716
rect 12709 8540 13440 8640
rect 6807 1532 7026 1544
rect 6807 1468 6820 1532
rect 6884 1468 6950 1532
rect 7014 1468 7026 1532
rect 6807 1456 7026 1468
rect 5844 1193 6063 1205
rect 5844 1129 5857 1193
rect 5921 1129 5987 1193
rect 6051 1129 6063 1193
rect 5844 1117 6063 1129
rect 4453 1026 4672 1038
rect 4453 962 4466 1026
rect 4530 962 4596 1026
rect 4660 962 4672 1026
rect 4453 950 4672 962
rect 5884 1037 5984 1117
rect 5884 937 6644 1037
rect 5846 531 6065 543
rect 5846 467 5859 531
rect 5923 467 5989 531
rect 6053 467 6065 531
rect 5846 455 6065 467
rect 5902 394 6002 455
rect 5902 294 6325 394
rect 6225 -442 6325 294
rect 6166 -454 6385 -442
rect 6166 -518 6179 -454
rect 6243 -518 6309 -454
rect 6373 -518 6385 -454
rect 6166 -530 6385 -518
rect 6544 -594 6644 937
rect 6863 -449 6963 1456
rect 7128 535 7347 547
rect 7128 471 7141 535
rect 7205 471 7271 535
rect 7335 471 7347 535
rect 7128 459 7347 471
rect 7177 51 7277 459
rect 7118 33 7327 51
rect 7118 -31 7131 33
rect 7195 -31 7251 33
rect 7315 -31 7327 33
rect 7118 -49 7327 -31
rect 6807 -461 7026 -449
rect 6807 -525 6820 -461
rect 6884 -525 6950 -461
rect 7014 -525 7026 -461
rect 6807 -537 7026 -525
rect 7127 -450 7346 -438
rect 7127 -514 7140 -450
rect 7204 -514 7270 -450
rect 7334 -514 7346 -450
rect 7127 -526 7346 -514
rect 7175 -594 7275 -526
rect 6544 -694 7275 -594
use ppolyf_u_GQDF3M  ppolyf_u_GQDF3M_0
timestamp 1694501647
transform 1 0 5996 0 1 8579
box -304 -386 304 386
use ppolyf_u_GQDF3M  ppolyf_u_GQDF3M_1
timestamp 1694501647
transform 1 0 14836 0 1 10535
box -304 -386 304 386
use ppolyf_u_GQDF3M  ppolyf_u_GQDF3M_2
timestamp 1694501647
transform 1 0 14836 0 1 9883
box -304 -386 304 386
use ppolyf_u_GQDF3M  ppolyf_u_GQDF3M_3
timestamp 1694501647
transform 1 0 14836 0 1 9231
box -304 -386 304 386
use ppolyf_u_GQDF3M  ppolyf_u_GQDF3M_4
timestamp 1694501647
transform 1 0 14836 0 1 8579
box -304 -386 304 386
use ppolyf_u_GQDF3M  ppolyf_u_GQDF3M_5
timestamp 1694501647
transform 1 0 5996 0 1 10535
box -304 -386 304 386
use ppolyf_u_GQDF3M  ppolyf_u_GQDF3M_6
timestamp 1694501647
transform 1 0 5996 0 1 9883
box -304 -386 304 386
use ppolyf_u_GQDF3M  ppolyf_u_GQDF3M_7
timestamp 1694501647
transform 1 0 5996 0 1 9231
box -304 -386 304 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_0
timestamp 1694501647
transform 1 0 7284 0 1 9231
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_1
timestamp 1694501647
transform 1 0 7284 0 1 9883
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_2
timestamp 1694501647
transform 1 0 7284 0 1 8579
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_3
timestamp 1694501647
transform -1 0 9372 0 1 9231
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_4
timestamp 1694501647
transform 1 0 6436 0 1 5
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_5
timestamp 1694501647
transform 1 0 6436 0 1 665
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_6
timestamp 1694501647
transform 1 0 6436 0 1 1325
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_7
timestamp 1694501647
transform 1 0 6436 0 1 -655
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_8
timestamp 1694501647
transform -1 0 9372 0 1 9883
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_9
timestamp 1694501647
transform -1 0 9372 0 1 8579
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_10
timestamp 1694501647
transform 1 0 7284 0 1 10535
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_11
timestamp 1694501647
transform -1 0 9372 0 1 10535
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_12
timestamp 1694501647
transform 1 0 11460 0 1 9231
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_13
timestamp 1694501647
transform 1 0 11460 0 1 9883
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_14
timestamp 1694501647
transform 1 0 11460 0 1 8579
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_15
timestamp 1694501647
transform -1 0 13548 0 1 9231
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_16
timestamp 1694501647
transform -1 0 13548 0 1 9883
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_17
timestamp 1694501647
transform -1 0 13548 0 1 8579
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_18
timestamp 1694501647
transform 1 0 11460 0 1 10535
box -1104 -386 1104 386
use ppolyf_u_GQDP2M  ppolyf_u_GQDP2M_19
timestamp 1694501647
transform -1 0 13548 0 1 10535
box -1104 -386 1104 386
use ppolyf_u_W5AMT6  ppolyf_u_W5AMT6_0
timestamp 1694513024
transform 1 0 9947 0 1 13138
box -4304 -386 4304 386
use ppolyf_u_W5AMT6  ppolyf_u_W5AMT6_1
timestamp 1694513024
transform 1 0 9947 0 1 15094
box -4304 -386 4304 386
use ppolyf_u_W5AMT6  ppolyf_u_W5AMT6_2
timestamp 1694513024
transform 1 0 9947 0 1 14442
box -4304 -386 4304 386
use ppolyf_u_W5AMT6  ppolyf_u_W5AMT6_3
timestamp 1694513024
transform 1 0 9947 0 1 13790
box -4304 -386 4304 386
<< labels >>
flabel metal1 6263 15330 6263 15330 0 FreeSans 1600 0 0 0 A
port 1 nsew
flabel metal1 13459 15339 13459 15339 0 FreeSans 1600 0 0 0 B
port 3 nsew
flabel metal1 6588 15339 6588 15339 0 FreeSans 1600 0 0 0 C
port 5 nsew
flabel metal2 12986 15349 12986 15349 0 FreeSans 1600 0 0 0 D
port 7 nsew
flabel metal1 5746 14447 5746 14447 0 FreeSans 1600 0 0 0 E
port 9 nsew
flabel metal1 14122 14758 14122 14758 0 FreeSans 1600 0 0 0 F
port 10 nsew
flabel metal1 5794 14766 5794 14766 0 FreeSans 1600 0 0 0 G
port 14 nsew
flabel metal1 14151 13143 14151 13143 0 FreeSans 1600 0 0 0 H
port 15 nsew
<< end >>
