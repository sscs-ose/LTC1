magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2208 -2120 2592 2550
<< nwell >>
rect -208 -120 592 550
<< mvpmos >>
rect 0 0 140 430
rect 244 0 384 430
<< mvpdiff >>
rect -88 417 0 430
rect -88 371 -75 417
rect -29 371 0 417
rect -88 298 0 371
rect -88 252 -75 298
rect -29 252 0 298
rect -88 179 0 252
rect -88 133 -75 179
rect -29 133 0 179
rect -88 59 0 133
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 417 244 430
rect 140 371 169 417
rect 215 371 244 417
rect 140 298 244 371
rect 140 252 169 298
rect 215 252 244 298
rect 140 179 244 252
rect 140 133 169 179
rect 215 133 244 179
rect 140 59 244 133
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 417 472 430
rect 384 371 413 417
rect 459 371 472 417
rect 384 298 472 371
rect 384 252 413 298
rect 459 252 472 298
rect 384 179 472 252
rect 384 133 413 179
rect 459 133 472 179
rect 384 59 472 133
rect 384 13 413 59
rect 459 13 472 59
rect 384 0 472 13
<< mvpdiffc >>
rect -75 371 -29 417
rect -75 252 -29 298
rect -75 133 -29 179
rect -75 13 -29 59
rect 169 371 215 417
rect 169 252 215 298
rect 169 133 215 179
rect 169 13 215 59
rect 413 371 459 417
rect 413 252 459 298
rect 413 133 459 179
rect 413 13 459 59
<< polysilicon >>
rect 0 430 140 474
rect 244 430 384 474
rect 0 -44 140 0
rect 244 -44 384 0
<< metal1 >>
rect -75 417 -29 430
rect -75 298 -29 371
rect -75 179 -29 252
rect -75 59 -29 133
rect -75 0 -29 13
rect 169 417 215 430
rect 169 298 215 371
rect 169 179 215 252
rect 169 59 215 133
rect 169 0 215 13
rect 413 417 459 430
rect 413 298 459 371
rect 413 179 459 252
rect 413 59 459 133
rect 413 0 459 13
<< labels >>
rlabel metal1 192 215 192 215 4 D
rlabel metal1 436 215 436 215 4 S
rlabel metal1 -52 215 -52 215 4 S
<< end >>
