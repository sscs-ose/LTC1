magic
tech gf180mcuC
magscale 1 10
timestamp 1693483456
<< error_p >>
rect -2154 -23 -2143 23
rect -1942 -23 -1931 23
rect -1730 -23 -1719 23
rect -1518 -23 -1507 23
rect -1306 -23 -1295 23
rect -1094 -23 -1083 23
rect -882 -23 -871 23
rect -670 -23 -659 23
rect -458 -23 -447 23
rect -246 -23 -235 23
rect -34 -23 -23 23
rect 178 -23 189 23
rect 390 -23 401 23
rect 602 -23 613 23
rect 814 -23 825 23
rect 1026 -23 1037 23
rect 1238 -23 1249 23
rect 1450 -23 1461 23
rect 1662 -23 1673 23
rect 1874 -23 1885 23
rect 2086 -23 2097 23
<< pwell >>
rect -2180 -97 2180 97
<< nmos >>
rect -2064 -22 -1964 22
rect -1852 -22 -1752 22
rect -1640 -22 -1540 22
rect -1428 -22 -1328 22
rect -1216 -22 -1116 22
rect -1004 -22 -904 22
rect -792 -22 -692 22
rect -580 -22 -480 22
rect -368 -22 -268 22
rect -156 -22 -56 22
rect 56 -22 156 22
rect 268 -22 368 22
rect 480 -22 580 22
rect 692 -22 792 22
rect 904 -22 1004 22
rect 1116 -22 1216 22
rect 1328 -22 1428 22
rect 1540 -22 1640 22
rect 1752 -22 1852 22
rect 1964 -22 2064 22
<< ndiff >>
rect -2156 23 -2084 36
rect -2156 -23 -2143 23
rect -2097 22 -2084 23
rect -1944 23 -1872 36
rect -1944 22 -1931 23
rect -2097 -22 -2064 22
rect -1964 -22 -1931 22
rect -2097 -23 -2084 -22
rect -2156 -36 -2084 -23
rect -1944 -23 -1931 -22
rect -1885 22 -1872 23
rect -1732 23 -1660 36
rect -1732 22 -1719 23
rect -1885 -22 -1852 22
rect -1752 -22 -1719 22
rect -1885 -23 -1872 -22
rect -1944 -36 -1872 -23
rect -1732 -23 -1719 -22
rect -1673 22 -1660 23
rect -1520 23 -1448 36
rect -1520 22 -1507 23
rect -1673 -22 -1640 22
rect -1540 -22 -1507 22
rect -1673 -23 -1660 -22
rect -1732 -36 -1660 -23
rect -1520 -23 -1507 -22
rect -1461 22 -1448 23
rect -1308 23 -1236 36
rect -1308 22 -1295 23
rect -1461 -22 -1428 22
rect -1328 -22 -1295 22
rect -1461 -23 -1448 -22
rect -1520 -36 -1448 -23
rect -1308 -23 -1295 -22
rect -1249 22 -1236 23
rect -1096 23 -1024 36
rect -1096 22 -1083 23
rect -1249 -22 -1216 22
rect -1116 -22 -1083 22
rect -1249 -23 -1236 -22
rect -1308 -36 -1236 -23
rect -1096 -23 -1083 -22
rect -1037 22 -1024 23
rect -884 23 -812 36
rect -884 22 -871 23
rect -1037 -22 -1004 22
rect -904 -22 -871 22
rect -1037 -23 -1024 -22
rect -1096 -36 -1024 -23
rect -884 -23 -871 -22
rect -825 22 -812 23
rect -672 23 -600 36
rect -672 22 -659 23
rect -825 -22 -792 22
rect -692 -22 -659 22
rect -825 -23 -812 -22
rect -884 -36 -812 -23
rect -672 -23 -659 -22
rect -613 22 -600 23
rect -460 23 -388 36
rect -460 22 -447 23
rect -613 -22 -580 22
rect -480 -22 -447 22
rect -613 -23 -600 -22
rect -672 -36 -600 -23
rect -460 -23 -447 -22
rect -401 22 -388 23
rect -248 23 -176 36
rect -248 22 -235 23
rect -401 -22 -368 22
rect -268 -22 -235 22
rect -401 -23 -388 -22
rect -460 -36 -388 -23
rect -248 -23 -235 -22
rect -189 22 -176 23
rect -36 23 36 36
rect -36 22 -23 23
rect -189 -22 -156 22
rect -56 -22 -23 22
rect -189 -23 -176 -22
rect -248 -36 -176 -23
rect -36 -23 -23 -22
rect 23 22 36 23
rect 176 23 248 36
rect 176 22 189 23
rect 23 -22 56 22
rect 156 -22 189 22
rect 23 -23 36 -22
rect -36 -36 36 -23
rect 176 -23 189 -22
rect 235 22 248 23
rect 388 23 460 36
rect 388 22 401 23
rect 235 -22 268 22
rect 368 -22 401 22
rect 235 -23 248 -22
rect 176 -36 248 -23
rect 388 -23 401 -22
rect 447 22 460 23
rect 600 23 672 36
rect 600 22 613 23
rect 447 -22 480 22
rect 580 -22 613 22
rect 447 -23 460 -22
rect 388 -36 460 -23
rect 600 -23 613 -22
rect 659 22 672 23
rect 812 23 884 36
rect 812 22 825 23
rect 659 -22 692 22
rect 792 -22 825 22
rect 659 -23 672 -22
rect 600 -36 672 -23
rect 812 -23 825 -22
rect 871 22 884 23
rect 1024 23 1096 36
rect 1024 22 1037 23
rect 871 -22 904 22
rect 1004 -22 1037 22
rect 871 -23 884 -22
rect 812 -36 884 -23
rect 1024 -23 1037 -22
rect 1083 22 1096 23
rect 1236 23 1308 36
rect 1236 22 1249 23
rect 1083 -22 1116 22
rect 1216 -22 1249 22
rect 1083 -23 1096 -22
rect 1024 -36 1096 -23
rect 1236 -23 1249 -22
rect 1295 22 1308 23
rect 1448 23 1520 36
rect 1448 22 1461 23
rect 1295 -22 1328 22
rect 1428 -22 1461 22
rect 1295 -23 1308 -22
rect 1236 -36 1308 -23
rect 1448 -23 1461 -22
rect 1507 22 1520 23
rect 1660 23 1732 36
rect 1660 22 1673 23
rect 1507 -22 1540 22
rect 1640 -22 1673 22
rect 1507 -23 1520 -22
rect 1448 -36 1520 -23
rect 1660 -23 1673 -22
rect 1719 22 1732 23
rect 1872 23 1944 36
rect 1872 22 1885 23
rect 1719 -22 1752 22
rect 1852 -22 1885 22
rect 1719 -23 1732 -22
rect 1660 -36 1732 -23
rect 1872 -23 1885 -22
rect 1931 22 1944 23
rect 2084 23 2156 36
rect 2084 22 2097 23
rect 1931 -22 1964 22
rect 2064 -22 2097 22
rect 1931 -23 1944 -22
rect 1872 -36 1944 -23
rect 2084 -23 2097 -22
rect 2143 -23 2156 23
rect 2084 -36 2156 -23
<< ndiffc >>
rect -2143 -23 -2097 23
rect -1931 -23 -1885 23
rect -1719 -23 -1673 23
rect -1507 -23 -1461 23
rect -1295 -23 -1249 23
rect -1083 -23 -1037 23
rect -871 -23 -825 23
rect -659 -23 -613 23
rect -447 -23 -401 23
rect -235 -23 -189 23
rect -23 -23 23 23
rect 189 -23 235 23
rect 401 -23 447 23
rect 613 -23 659 23
rect 825 -23 871 23
rect 1037 -23 1083 23
rect 1249 -23 1295 23
rect 1461 -23 1507 23
rect 1673 -23 1719 23
rect 1885 -23 1931 23
rect 2097 -23 2143 23
<< polysilicon >>
rect -2064 22 -1964 66
rect -2064 -66 -1964 -22
rect -1852 22 -1752 66
rect -1852 -66 -1752 -22
rect -1640 22 -1540 66
rect -1640 -66 -1540 -22
rect -1428 22 -1328 66
rect -1428 -66 -1328 -22
rect -1216 22 -1116 66
rect -1216 -66 -1116 -22
rect -1004 22 -904 66
rect -1004 -66 -904 -22
rect -792 22 -692 66
rect -792 -66 -692 -22
rect -580 22 -480 66
rect -580 -66 -480 -22
rect -368 22 -268 66
rect -368 -66 -268 -22
rect -156 22 -56 66
rect -156 -66 -56 -22
rect 56 22 156 66
rect 56 -66 156 -22
rect 268 22 368 66
rect 268 -66 368 -22
rect 480 22 580 66
rect 480 -66 580 -22
rect 692 22 792 66
rect 692 -66 792 -22
rect 904 22 1004 66
rect 904 -66 1004 -22
rect 1116 22 1216 66
rect 1116 -66 1216 -22
rect 1328 22 1428 66
rect 1328 -66 1428 -22
rect 1540 22 1640 66
rect 1540 -66 1640 -22
rect 1752 22 1852 66
rect 1752 -66 1852 -22
rect 1964 22 2064 66
rect 1964 -66 2064 -22
<< metal1 >>
rect -2154 -23 -2143 23
rect -2097 -23 -2086 23
rect -1942 -23 -1931 23
rect -1885 -23 -1874 23
rect -1730 -23 -1719 23
rect -1673 -23 -1662 23
rect -1518 -23 -1507 23
rect -1461 -23 -1450 23
rect -1306 -23 -1295 23
rect -1249 -23 -1238 23
rect -1094 -23 -1083 23
rect -1037 -23 -1026 23
rect -882 -23 -871 23
rect -825 -23 -814 23
rect -670 -23 -659 23
rect -613 -23 -602 23
rect -458 -23 -447 23
rect -401 -23 -390 23
rect -246 -23 -235 23
rect -189 -23 -178 23
rect -34 -23 -23 23
rect 23 -23 34 23
rect 178 -23 189 23
rect 235 -23 246 23
rect 390 -23 401 23
rect 447 -23 458 23
rect 602 -23 613 23
rect 659 -23 670 23
rect 814 -23 825 23
rect 871 -23 882 23
rect 1026 -23 1037 23
rect 1083 -23 1094 23
rect 1238 -23 1249 23
rect 1295 -23 1306 23
rect 1450 -23 1461 23
rect 1507 -23 1518 23
rect 1662 -23 1673 23
rect 1719 -23 1730 23
rect 1874 -23 1885 23
rect 1931 -23 1942 23
rect 2086 -23 2097 23
rect 2143 -23 2154 23
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.22 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
