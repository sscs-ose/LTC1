magic
tech gf180mcuC
magscale 1 10
timestamp 1693911244
<< nwell >>
rect -442 -1902 442 1902
<< pmos >>
rect -268 1172 -212 1772
rect -108 1172 -52 1772
rect 52 1172 108 1772
rect 212 1172 268 1772
rect -268 436 -212 1036
rect -108 436 -52 1036
rect 52 436 108 1036
rect 212 436 268 1036
rect -268 -300 -212 300
rect -108 -300 -52 300
rect 52 -300 108 300
rect 212 -300 268 300
rect -268 -1036 -212 -436
rect -108 -1036 -52 -436
rect 52 -1036 108 -436
rect 212 -1036 268 -436
rect -268 -1772 -212 -1172
rect -108 -1772 -52 -1172
rect 52 -1772 108 -1172
rect 212 -1772 268 -1172
<< pdiff >>
rect -356 1759 -268 1772
rect -356 1185 -343 1759
rect -297 1185 -268 1759
rect -356 1172 -268 1185
rect -212 1759 -108 1772
rect -212 1185 -183 1759
rect -137 1185 -108 1759
rect -212 1172 -108 1185
rect -52 1759 52 1772
rect -52 1185 -23 1759
rect 23 1185 52 1759
rect -52 1172 52 1185
rect 108 1759 212 1772
rect 108 1185 137 1759
rect 183 1185 212 1759
rect 108 1172 212 1185
rect 268 1759 356 1772
rect 268 1185 297 1759
rect 343 1185 356 1759
rect 268 1172 356 1185
rect -356 1023 -268 1036
rect -356 449 -343 1023
rect -297 449 -268 1023
rect -356 436 -268 449
rect -212 1023 -108 1036
rect -212 449 -183 1023
rect -137 449 -108 1023
rect -212 436 -108 449
rect -52 1023 52 1036
rect -52 449 -23 1023
rect 23 449 52 1023
rect -52 436 52 449
rect 108 1023 212 1036
rect 108 449 137 1023
rect 183 449 212 1023
rect 108 436 212 449
rect 268 1023 356 1036
rect 268 449 297 1023
rect 343 449 356 1023
rect 268 436 356 449
rect -356 287 -268 300
rect -356 -287 -343 287
rect -297 -287 -268 287
rect -356 -300 -268 -287
rect -212 287 -108 300
rect -212 -287 -183 287
rect -137 -287 -108 287
rect -212 -300 -108 -287
rect -52 287 52 300
rect -52 -287 -23 287
rect 23 -287 52 287
rect -52 -300 52 -287
rect 108 287 212 300
rect 108 -287 137 287
rect 183 -287 212 287
rect 108 -300 212 -287
rect 268 287 356 300
rect 268 -287 297 287
rect 343 -287 356 287
rect 268 -300 356 -287
rect -356 -449 -268 -436
rect -356 -1023 -343 -449
rect -297 -1023 -268 -449
rect -356 -1036 -268 -1023
rect -212 -449 -108 -436
rect -212 -1023 -183 -449
rect -137 -1023 -108 -449
rect -212 -1036 -108 -1023
rect -52 -449 52 -436
rect -52 -1023 -23 -449
rect 23 -1023 52 -449
rect -52 -1036 52 -1023
rect 108 -449 212 -436
rect 108 -1023 137 -449
rect 183 -1023 212 -449
rect 108 -1036 212 -1023
rect 268 -449 356 -436
rect 268 -1023 297 -449
rect 343 -1023 356 -449
rect 268 -1036 356 -1023
rect -356 -1185 -268 -1172
rect -356 -1759 -343 -1185
rect -297 -1759 -268 -1185
rect -356 -1772 -268 -1759
rect -212 -1185 -108 -1172
rect -212 -1759 -183 -1185
rect -137 -1759 -108 -1185
rect -212 -1772 -108 -1759
rect -52 -1185 52 -1172
rect -52 -1759 -23 -1185
rect 23 -1759 52 -1185
rect -52 -1772 52 -1759
rect 108 -1185 212 -1172
rect 108 -1759 137 -1185
rect 183 -1759 212 -1185
rect 108 -1772 212 -1759
rect 268 -1185 356 -1172
rect 268 -1759 297 -1185
rect 343 -1759 356 -1185
rect 268 -1772 356 -1759
<< pdiffc >>
rect -343 1185 -297 1759
rect -183 1185 -137 1759
rect -23 1185 23 1759
rect 137 1185 183 1759
rect 297 1185 343 1759
rect -343 449 -297 1023
rect -183 449 -137 1023
rect -23 449 23 1023
rect 137 449 183 1023
rect 297 449 343 1023
rect -343 -287 -297 287
rect -183 -287 -137 287
rect -23 -287 23 287
rect 137 -287 183 287
rect 297 -287 343 287
rect -343 -1023 -297 -449
rect -183 -1023 -137 -449
rect -23 -1023 23 -449
rect 137 -1023 183 -449
rect 297 -1023 343 -449
rect -343 -1759 -297 -1185
rect -183 -1759 -137 -1185
rect -23 -1759 23 -1185
rect 137 -1759 183 -1185
rect 297 -1759 343 -1185
<< polysilicon >>
rect -268 1772 -212 1816
rect -108 1772 -52 1816
rect 52 1772 108 1816
rect 212 1772 268 1816
rect -268 1128 -212 1172
rect -108 1128 -52 1172
rect 52 1128 108 1172
rect 212 1128 268 1172
rect -268 1036 -212 1080
rect -108 1036 -52 1080
rect 52 1036 108 1080
rect 212 1036 268 1080
rect -268 392 -212 436
rect -108 392 -52 436
rect 52 392 108 436
rect 212 392 268 436
rect -268 300 -212 344
rect -108 300 -52 344
rect 52 300 108 344
rect 212 300 268 344
rect -268 -344 -212 -300
rect -108 -344 -52 -300
rect 52 -344 108 -300
rect 212 -344 268 -300
rect -268 -436 -212 -392
rect -108 -436 -52 -392
rect 52 -436 108 -392
rect 212 -436 268 -392
rect -268 -1080 -212 -1036
rect -108 -1080 -52 -1036
rect 52 -1080 108 -1036
rect 212 -1080 268 -1036
rect -268 -1172 -212 -1128
rect -108 -1172 -52 -1128
rect 52 -1172 108 -1128
rect 212 -1172 268 -1128
rect -268 -1816 -212 -1772
rect -108 -1816 -52 -1772
rect 52 -1816 108 -1772
rect 212 -1816 268 -1772
<< metal1 >>
rect -343 1759 -297 1770
rect -343 1174 -297 1185
rect -183 1759 -137 1770
rect -183 1174 -137 1185
rect -23 1759 23 1770
rect -23 1174 23 1185
rect 137 1759 183 1770
rect 137 1174 183 1185
rect 297 1759 343 1770
rect 297 1174 343 1185
rect -343 1023 -297 1034
rect -343 438 -297 449
rect -183 1023 -137 1034
rect -183 438 -137 449
rect -23 1023 23 1034
rect -23 438 23 449
rect 137 1023 183 1034
rect 137 438 183 449
rect 297 1023 343 1034
rect 297 438 343 449
rect -343 287 -297 298
rect -343 -298 -297 -287
rect -183 287 -137 298
rect -183 -298 -137 -287
rect -23 287 23 298
rect -23 -298 23 -287
rect 137 287 183 298
rect 137 -298 183 -287
rect 297 287 343 298
rect 297 -298 343 -287
rect -343 -449 -297 -438
rect -343 -1034 -297 -1023
rect -183 -449 -137 -438
rect -183 -1034 -137 -1023
rect -23 -449 23 -438
rect -23 -1034 23 -1023
rect 137 -449 183 -438
rect 137 -1034 183 -1023
rect 297 -449 343 -438
rect 297 -1034 343 -1023
rect -343 -1185 -297 -1174
rect -343 -1770 -297 -1759
rect -183 -1185 -137 -1174
rect -183 -1770 -137 -1759
rect -23 -1185 23 -1174
rect -23 -1770 23 -1759
rect 137 -1185 183 -1174
rect 137 -1770 183 -1759
rect 297 -1185 343 -1174
rect 297 -1770 343 -1759
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 5 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
