** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/pex_4x1_mux_TB_ibr..sym
**.subckt pex_4x1_mux_TB_ibr.
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V4 S0 VSS pulse(3.3 0 0 100p 100p 200n 400n)
.save i(v4)
V6 I0 VSS pulse(0 3.3 0 100p 100p 100n 200n)3.3
.save i(v6)
V7 I1 VSS pulse(0 3.3 0 100p 100p 200n 400n)
.save i(v7)
V5 S1 VSS pulse(3.3 0 0 100p 100p 400n 800n)
.save i(v5)
V3 I2 VSS pulse(0 3.3 0 100p 100p 400n 800n)3.3
.save i(v3)
V8 I3 VSS pulse(0 3.3 0 100p 100p 800n 1600n)3.3
.save i(v8)
x1 VDD S1 VSS I2 I3 S0 I0 I1 OUT pex_mux_4x1_ibr
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_mux_4x1_ibr.spice
.control
save all
tran 50p 800n
plot v(S0) v(S1)+4  v(I0)+8 v(I1)+12 I2+16 I3+20  v(OUT)+24


*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
