* NGSPICE file created from inv_flat.ext - technology: gf180mcuC

.subckt inv_flat VDD VSS IN OUT
X0 OUT IN.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 OUT IN.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
R0 IN.n0 IN.t0 25.4398
R1 IN.n0 IN.t1 17.6975
R2 IN IN.n0 4.24656
R3 VDD.n0 VDD.t0 547.89
R4 VDD VDD.n0 6.3005
R5 VDD VDD.n0 6.3005
R6 VDD VDD.t1 5.2211
R7 OUT.n2 OUT.n1 9.40108
R8 OUT.n2 OUT.n0 5.21162
R9 OUT OUT.n2 0.143142
R10 VSS.n1 VSS.t0 1603.59
R11 VSS.n2 VSS.t1 9.44211
R12 VSS.n2 VSS.n1 2.6005
R13 VSS.n1 VSS.n0 0.0926053
R14 VSS VSS.n2 0.00128947
C0 OUT IN 0.111f
C1 VDD IN 0.184f
C2 OUT VDD 0.131f
.ends

