** sch_path: /home/shahid/OSPDKs/gf180mcuC/libs.tech/xschem/gf180mcu_tests/test_cap_mim_2p0fF.sch
**.subckt test_cap_mim_2p0fF
XC1 P GND cap_mim_2f0fF c_width=10e-6 c_length=10e-6 m=10
V1 IN GND pwl 0 0 200n 3.3
.save i(v1)
R2 P IN 100k m=1
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
* .lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_statistical



.control
save all
tran 0.1n 200n
write test_cap_mim_2p0fF.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
