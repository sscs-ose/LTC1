* NGSPICE file created from nmos_3p3_GGGST2_flat.ext - technology: gf180mcuC

.subckt nmos_3p3_GGGST2_flat A B C OUT VDD VSS
X0 OUT a_24_68.t6 VDD.t6 VDD.t5 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1 OUT a_24_68.t7 VSS.t9 VSS.t8 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 VSS C.t0 a_648_68.t0 VSS.t1 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X3 VDD C.t2 a_24_68.t0 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 VSS C.t3 a_648_68.t5 VSS.t13 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 VDD A.t3 a_24_68.t3 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
R0 a_24_68.n0 a_24_68.t7 63.282
R1 a_24_68.n0 a_24_68.t6 43.207
R2 a_24_68.n3 a_24_68.t1 7.2365
R3 a_24_68.n5 a_24_68.n0 4.89072
R4 a_24_68.n4 a_24_68.t3 4.72376
R5 a_24_68.n3 a_24_68.n2 3.33441
R6 a_24_68.n2 a_24_68.t5 3.2765
R7 a_24_68.n2 a_24_68.n1 3.2765
R8 a_24_68.n7 a_24_68.n5 2.90376
R9 a_24_68.t0 a_24_68.n7 1.8205
R10 a_24_68.n7 a_24_68.n6 1.8205
R11 a_24_68.n5 a_24_68.n4 0.626587
R12 a_24_68.n4 a_24_68.n3 0.472022
R13 VDD.n9 VDD.t0 154.44
R14 VDD.n4 VDD.t5 85.6379
R15 VDD.n15 VDD.t7 85.6365
R16 VDD.t0 VDD.n8 27.0275
R17 VDD.n17 VDD.t3 27.0275
R18 VDD.n10 VDD.n7 8.2255
R19 VDD.n18 VDD.n10 8.2255
R20 VDD VDD.n10 6.3005
R21 VDD VDD.n10 6.3005
R22 VDD.n3 VDD.n2 3.1505
R23 VDD.n7 VDD.n6 3.1505
R24 VDD.n8 VDD.n7 3.1505
R25 VDD.n10 VDD.n9 3.1505
R26 VDD.n19 VDD.n18 3.1505
R27 VDD.n18 VDD.n17 3.1505
R28 VDD.n14 VDD.n13 3.1505
R29 VDD.n5 VDD.n1 2.91941
R30 VDD.n16 VDD.n12 2.91705
R31 VDD.n4 VDD.n3 1.87098
R32 VDD.n15 VDD.n14 1.8708
R33 VDD.n12 VDD.t4 1.8205
R34 VDD.n12 VDD.n11 1.8205
R35 VDD.n1 VDD.t6 1.8205
R36 VDD.n1 VDD.n0 1.8205
R37 VDD.n5 VDD.n4 0.58998
R38 VDD.n16 VDD.n15 0.588573
R39 VDD VDD.n6 0.0760357
R40 VDD VDD.n19 0.0760357
R41 VDD.n19 VDD.n16 0.0551429
R42 VDD.n6 VDD.n5 0.0535357
R43 OUT.n2 OUT.n0 7.06041
R44 OUT.n2 OUT.n1 5.46137
R45 OUT OUT.n2 0.196152
R46 A.n1 A.t3 39.6291
R47 A.n0 A.t1 29.9826
R48 A.t2 A.n0 29.9826
R49 A.n1 A.t2 28.9398
R50 A A.n1 21.7803
R51 A.n0 A.t0 9.1255
R52 a_168_68.n4 a_168_68.n3 3.9605
R53 a_168_68.n5 a_168_68.n4 3.9605
R54 a_168_68.n4 a_168_68.n1 3.33441
R55 a_168_68.n3 a_168_68.t0 3.2765
R56 a_168_68.n3 a_168_68.n2 3.2765
R57 a_168_68.n1 a_168_68.t2 3.2765
R58 a_168_68.n1 a_168_68.n0 3.2765
R59 a_168_68.n5 a_168_68.t5 3.2765
R60 a_168_68.n6 a_168_68.n5 3.2765
R61 VSS.n13 VSS.t1 231.768
R62 VSS.n36 VSS.t12 221.232
R63 VSS.n0 VSS.t0 179.093
R64 VSS.n52 VSS.t6 168.559
R65 VSS.n39 VSS.t10 126.418
R66 VSS.n16 VSS.t4 115.883
R67 VSS.n6 VSS.t8 84.2793
R68 VSS.n30 VSS.t11 73.7444
R69 VSS.n23 VSS.t13 31.605
R70 VSS.n45 VSS.t7 21.0702
R71 VSS VSS.n1 4.66717
R72 VSS VSS.n53 4.47272
R73 VSS.n9 VSS.n5 3.76289
R74 VSS.n22 VSS.n3 3.76289
R75 VSS.n5 VSS.t9 3.2765
R76 VSS.n5 VSS.n4 3.2765
R77 VSS.n3 VSS.t5 3.2765
R78 VSS.n3 VSS.n2 3.2765
R79 VSS.n7 VSS.n6 2.6005
R80 VSS.n12 VSS.n11 2.6005
R81 VSS.n11 VSS.n10 2.6005
R82 VSS.n15 VSS.n14 2.6005
R83 VSS.n14 VSS.n13 2.6005
R84 VSS.n18 VSS.n17 2.6005
R85 VSS.n17 VSS.n16 2.6005
R86 VSS.n21 VSS.n20 2.6005
R87 VSS.n20 VSS.n19 2.6005
R88 VSS.n25 VSS.n24 2.6005
R89 VSS.n24 VSS.n23 2.6005
R90 VSS.n28 VSS.n27 2.6005
R91 VSS.n27 VSS.n26 2.6005
R92 VSS.n1 VSS.n0 2.6005
R93 VSS.n53 VSS.n51 2.6005
R94 VSS.n53 VSS.n52 2.6005
R95 VSS.n50 VSS.n49 2.6005
R96 VSS.n49 VSS.n48 2.6005
R97 VSS.n47 VSS.n46 2.6005
R98 VSS.n46 VSS.n45 2.6005
R99 VSS.n44 VSS.n43 2.6005
R100 VSS.n43 VSS.n42 2.6005
R101 VSS.n41 VSS.n40 2.6005
R102 VSS.n40 VSS.n39 2.6005
R103 VSS.n38 VSS.n37 2.6005
R104 VSS.n37 VSS.n36 2.6005
R105 VSS.n35 VSS.n34 2.6005
R106 VSS.n34 VSS.n33 2.6005
R107 VSS.n31 VSS.n30 2.6005
R108 VSS.n8 VSS.n7 1.64943
R109 VSS.n32 VSS.n31 1.64943
R110 VSS.n35 VSS.n32 0.559135
R111 VSS.n9 VSS.n8 0.535028
R112 VSS.n15 VSS.n12 0.0760357
R113 VSS.n18 VSS.n15 0.0760357
R114 VSS.n21 VSS.n18 0.0760357
R115 VSS.n28 VSS.n25 0.0760357
R116 VSS.n29 VSS.n28 0.0760357
R117 VSS.n51 VSS.n29 0.0760357
R118 VSS.n51 VSS.n50 0.0760357
R119 VSS.n50 VSS.n47 0.0760357
R120 VSS.n47 VSS.n44 0.0760357
R121 VSS.n44 VSS.n41 0.0760357
R122 VSS.n41 VSS.n38 0.0760357
R123 VSS.n38 VSS.n35 0.0760357
R124 VSS.n25 VSS.n22 0.0696071
R125 VSS.n12 VSS.n9 0.0246071
R126 VSS.n22 VSS.n21 0.00692857
R127 B.t2 B.t1 55.0112
R128 B.n0 B.t0 29.9826
R129 B B.n1 27.1952
R130 B.n1 B.t3 22.5523
R131 B.n0 B.t2 9.1255
R132 B.n1 B.n0 7.43086
R133 a_648_68.n4 a_648_68.n3 3.9605
R134 a_648_68.n4 a_648_68.n1 3.9605
R135 a_648_68.n5 a_648_68.n4 3.33441
R136 a_648_68.n3 a_648_68.t3 3.2765
R137 a_648_68.n3 a_648_68.n2 3.2765
R138 a_648_68.n1 a_648_68.t0 3.2765
R139 a_648_68.n1 a_648_68.n0 3.2765
R140 a_648_68.n5 a_648_68.t5 3.2765
R141 a_648_68.n6 a_648_68.n5 3.2765
R142 C.t3 C.t2 68.5684
R143 C C.n1 37.2709
R144 C.n0 C.t3 29.9826
R145 C.n1 C.n0 20.8576
R146 C.n1 C.t0 9.1255
R147 C.n0 C.t1 9.1255
C0 B C 0.061f
C1 A B 0.0428f
C2 B OUT 1.47e-19
C3 VDD C 0.136f
C4 A VDD 0.17f
C5 VDD OUT 0.147f
C6 VDD B 0.109f
C7 C OUT 0.0364f
.ends

