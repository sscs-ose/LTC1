magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1247 -1133 1247 1133
<< metal1 >>
rect -247 127 247 133
rect -247 101 -241 127
rect -215 101 -165 127
rect -139 101 -89 127
rect -63 101 -13 127
rect 13 101 63 127
rect 89 101 139 127
rect 165 101 215 127
rect 241 101 247 127
rect -247 51 247 101
rect -247 25 -241 51
rect -215 25 -165 51
rect -139 25 -89 51
rect -63 25 -13 51
rect 13 25 63 51
rect 89 25 139 51
rect 165 25 215 51
rect 241 25 247 51
rect -247 -25 247 25
rect -247 -51 -241 -25
rect -215 -51 -165 -25
rect -139 -51 -89 -25
rect -63 -51 -13 -25
rect 13 -51 63 -25
rect 89 -51 139 -25
rect 165 -51 215 -25
rect 241 -51 247 -25
rect -247 -101 247 -51
rect -247 -127 -241 -101
rect -215 -127 -165 -101
rect -139 -127 -89 -101
rect -63 -127 -13 -101
rect 13 -127 63 -101
rect 89 -127 139 -101
rect 165 -127 215 -101
rect 241 -127 247 -101
rect -247 -133 247 -127
<< via1 >>
rect -241 101 -215 127
rect -165 101 -139 127
rect -89 101 -63 127
rect -13 101 13 127
rect 63 101 89 127
rect 139 101 165 127
rect 215 101 241 127
rect -241 25 -215 51
rect -165 25 -139 51
rect -89 25 -63 51
rect -13 25 13 51
rect 63 25 89 51
rect 139 25 165 51
rect 215 25 241 51
rect -241 -51 -215 -25
rect -165 -51 -139 -25
rect -89 -51 -63 -25
rect -13 -51 13 -25
rect 63 -51 89 -25
rect 139 -51 165 -25
rect 215 -51 241 -25
rect -241 -127 -215 -101
rect -165 -127 -139 -101
rect -89 -127 -63 -101
rect -13 -127 13 -101
rect 63 -127 89 -101
rect 139 -127 165 -101
rect 215 -127 241 -101
<< metal2 >>
rect -247 127 247 133
rect -247 101 -241 127
rect -215 101 -165 127
rect -139 101 -89 127
rect -63 101 -13 127
rect 13 101 63 127
rect 89 101 139 127
rect 165 101 215 127
rect 241 101 247 127
rect -247 51 247 101
rect -247 25 -241 51
rect -215 25 -165 51
rect -139 25 -89 51
rect -63 25 -13 51
rect 13 25 63 51
rect 89 25 139 51
rect 165 25 215 51
rect 241 25 247 51
rect -247 -25 247 25
rect -247 -51 -241 -25
rect -215 -51 -165 -25
rect -139 -51 -89 -25
rect -63 -51 -13 -25
rect 13 -51 63 -25
rect 89 -51 139 -25
rect 165 -51 215 -25
rect 241 -51 247 -25
rect -247 -101 247 -51
rect -247 -127 -241 -101
rect -215 -127 -165 -101
rect -139 -127 -89 -101
rect -63 -127 -13 -101
rect 13 -127 63 -101
rect 89 -127 139 -101
rect 165 -127 215 -101
rect 241 -127 247 -101
rect -247 -133 247 -127
<< end >>
