magic
tech gf180mcuC
magscale 1 10
timestamp 1691428809
<< error_p >>
rect -343 70 -297 166
rect -183 70 -137 166
rect -23 70 23 166
rect 137 70 183 166
rect 297 70 343 166
rect -343 -166 -297 -70
rect -183 -166 -137 -70
rect -23 -166 23 -70
rect 137 -166 183 -70
rect 297 -166 343 -70
<< pwell >>
rect -380 -236 380 236
<< nmos >>
rect -268 68 -212 168
rect -108 68 -52 168
rect 52 68 108 168
rect 212 68 268 168
rect -268 -168 -212 -68
rect -108 -168 -52 -68
rect 52 -168 108 -68
rect 212 -168 268 -68
<< ndiff >>
rect -356 155 -268 168
rect -356 81 -343 155
rect -297 81 -268 155
rect -356 68 -268 81
rect -212 155 -108 168
rect -212 81 -183 155
rect -137 81 -108 155
rect -212 68 -108 81
rect -52 155 52 168
rect -52 81 -23 155
rect 23 81 52 155
rect -52 68 52 81
rect 108 155 212 168
rect 108 81 137 155
rect 183 81 212 155
rect 108 68 212 81
rect 268 155 356 168
rect 268 81 297 155
rect 343 81 356 155
rect 268 68 356 81
rect -356 -81 -268 -68
rect -356 -155 -343 -81
rect -297 -155 -268 -81
rect -356 -168 -268 -155
rect -212 -81 -108 -68
rect -212 -155 -183 -81
rect -137 -155 -108 -81
rect -212 -168 -108 -155
rect -52 -81 52 -68
rect -52 -155 -23 -81
rect 23 -155 52 -81
rect -52 -168 52 -155
rect 108 -81 212 -68
rect 108 -155 137 -81
rect 183 -155 212 -81
rect 108 -168 212 -155
rect 268 -81 356 -68
rect 268 -155 297 -81
rect 343 -155 356 -81
rect 268 -168 356 -155
<< ndiffc >>
rect -343 81 -297 155
rect -183 81 -137 155
rect -23 81 23 155
rect 137 81 183 155
rect 297 81 343 155
rect -343 -155 -297 -81
rect -183 -155 -137 -81
rect -23 -155 23 -81
rect 137 -155 183 -81
rect 297 -155 343 -81
<< polysilicon >>
rect -268 168 -212 212
rect -108 168 -52 212
rect 52 168 108 212
rect 212 168 268 212
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect -268 -212 -212 -168
rect -108 -212 -52 -168
rect 52 -212 108 -168
rect 212 -212 268 -168
<< metal1 >>
rect -343 155 -297 166
rect -343 70 -297 81
rect -183 155 -137 166
rect -183 70 -137 81
rect -23 155 23 166
rect -23 70 23 81
rect 137 155 183 166
rect 137 70 183 81
rect 297 155 343 166
rect 297 70 343 81
rect -343 -81 -297 -70
rect -343 -166 -297 -155
rect -183 -81 -137 -70
rect -183 -166 -137 -155
rect -23 -81 23 -70
rect -23 -166 23 -155
rect 137 -81 183 -70
rect 137 -166 183 -155
rect 297 -81 343 -70
rect 297 -166 343 -155
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.5 l 0.280 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
