magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1285 -1285 1285 1285
<< metal1 >>
rect -285 279 285 285
rect -285 253 -279 279
rect -253 253 -203 279
rect -177 253 -127 279
rect -101 253 -51 279
rect -25 253 25 279
rect 51 253 101 279
rect 127 253 177 279
rect 203 253 253 279
rect 279 253 285 279
rect -285 203 285 253
rect -285 177 -279 203
rect -253 177 -203 203
rect -177 177 -127 203
rect -101 177 -51 203
rect -25 177 25 203
rect 51 177 101 203
rect 127 177 177 203
rect 203 177 253 203
rect 279 177 285 203
rect -285 127 285 177
rect -285 101 -279 127
rect -253 101 -203 127
rect -177 101 -127 127
rect -101 101 -51 127
rect -25 101 25 127
rect 51 101 101 127
rect 127 101 177 127
rect 203 101 253 127
rect 279 101 285 127
rect -285 51 285 101
rect -285 25 -279 51
rect -253 25 -203 51
rect -177 25 -127 51
rect -101 25 -51 51
rect -25 25 25 51
rect 51 25 101 51
rect 127 25 177 51
rect 203 25 253 51
rect 279 25 285 51
rect -285 -25 285 25
rect -285 -51 -279 -25
rect -253 -51 -203 -25
rect -177 -51 -127 -25
rect -101 -51 -51 -25
rect -25 -51 25 -25
rect 51 -51 101 -25
rect 127 -51 177 -25
rect 203 -51 253 -25
rect 279 -51 285 -25
rect -285 -101 285 -51
rect -285 -127 -279 -101
rect -253 -127 -203 -101
rect -177 -127 -127 -101
rect -101 -127 -51 -101
rect -25 -127 25 -101
rect 51 -127 101 -101
rect 127 -127 177 -101
rect 203 -127 253 -101
rect 279 -127 285 -101
rect -285 -177 285 -127
rect -285 -203 -279 -177
rect -253 -203 -203 -177
rect -177 -203 -127 -177
rect -101 -203 -51 -177
rect -25 -203 25 -177
rect 51 -203 101 -177
rect 127 -203 177 -177
rect 203 -203 253 -177
rect 279 -203 285 -177
rect -285 -253 285 -203
rect -285 -279 -279 -253
rect -253 -279 -203 -253
rect -177 -279 -127 -253
rect -101 -279 -51 -253
rect -25 -279 25 -253
rect 51 -279 101 -253
rect 127 -279 177 -253
rect 203 -279 253 -253
rect 279 -279 285 -253
rect -285 -285 285 -279
<< via1 >>
rect -279 253 -253 279
rect -203 253 -177 279
rect -127 253 -101 279
rect -51 253 -25 279
rect 25 253 51 279
rect 101 253 127 279
rect 177 253 203 279
rect 253 253 279 279
rect -279 177 -253 203
rect -203 177 -177 203
rect -127 177 -101 203
rect -51 177 -25 203
rect 25 177 51 203
rect 101 177 127 203
rect 177 177 203 203
rect 253 177 279 203
rect -279 101 -253 127
rect -203 101 -177 127
rect -127 101 -101 127
rect -51 101 -25 127
rect 25 101 51 127
rect 101 101 127 127
rect 177 101 203 127
rect 253 101 279 127
rect -279 25 -253 51
rect -203 25 -177 51
rect -127 25 -101 51
rect -51 25 -25 51
rect 25 25 51 51
rect 101 25 127 51
rect 177 25 203 51
rect 253 25 279 51
rect -279 -51 -253 -25
rect -203 -51 -177 -25
rect -127 -51 -101 -25
rect -51 -51 -25 -25
rect 25 -51 51 -25
rect 101 -51 127 -25
rect 177 -51 203 -25
rect 253 -51 279 -25
rect -279 -127 -253 -101
rect -203 -127 -177 -101
rect -127 -127 -101 -101
rect -51 -127 -25 -101
rect 25 -127 51 -101
rect 101 -127 127 -101
rect 177 -127 203 -101
rect 253 -127 279 -101
rect -279 -203 -253 -177
rect -203 -203 -177 -177
rect -127 -203 -101 -177
rect -51 -203 -25 -177
rect 25 -203 51 -177
rect 101 -203 127 -177
rect 177 -203 203 -177
rect 253 -203 279 -177
rect -279 -279 -253 -253
rect -203 -279 -177 -253
rect -127 -279 -101 -253
rect -51 -279 -25 -253
rect 25 -279 51 -253
rect 101 -279 127 -253
rect 177 -279 203 -253
rect 253 -279 279 -253
<< metal2 >>
rect -285 279 285 285
rect -285 253 -279 279
rect -253 253 -203 279
rect -177 253 -127 279
rect -101 253 -51 279
rect -25 253 25 279
rect 51 253 101 279
rect 127 253 177 279
rect 203 253 253 279
rect 279 253 285 279
rect -285 203 285 253
rect -285 177 -279 203
rect -253 177 -203 203
rect -177 177 -127 203
rect -101 177 -51 203
rect -25 177 25 203
rect 51 177 101 203
rect 127 177 177 203
rect 203 177 253 203
rect 279 177 285 203
rect -285 127 285 177
rect -285 101 -279 127
rect -253 101 -203 127
rect -177 101 -127 127
rect -101 101 -51 127
rect -25 101 25 127
rect 51 101 101 127
rect 127 101 177 127
rect 203 101 253 127
rect 279 101 285 127
rect -285 51 285 101
rect -285 25 -279 51
rect -253 25 -203 51
rect -177 25 -127 51
rect -101 25 -51 51
rect -25 25 25 51
rect 51 25 101 51
rect 127 25 177 51
rect 203 25 253 51
rect 279 25 285 51
rect -285 -25 285 25
rect -285 -51 -279 -25
rect -253 -51 -203 -25
rect -177 -51 -127 -25
rect -101 -51 -51 -25
rect -25 -51 25 -25
rect 51 -51 101 -25
rect 127 -51 177 -25
rect 203 -51 253 -25
rect 279 -51 285 -25
rect -285 -101 285 -51
rect -285 -127 -279 -101
rect -253 -127 -203 -101
rect -177 -127 -127 -101
rect -101 -127 -51 -101
rect -25 -127 25 -101
rect 51 -127 101 -101
rect 127 -127 177 -101
rect 203 -127 253 -101
rect 279 -127 285 -101
rect -285 -177 285 -127
rect -285 -203 -279 -177
rect -253 -203 -203 -177
rect -177 -203 -127 -177
rect -101 -203 -51 -177
rect -25 -203 25 -177
rect 51 -203 101 -177
rect 127 -203 177 -177
rect 203 -203 253 -177
rect 279 -203 285 -177
rect -285 -253 285 -203
rect -285 -279 -279 -253
rect -253 -279 -203 -253
rect -177 -279 -127 -253
rect -101 -279 -51 -253
rect -25 -279 25 -253
rect 51 -279 101 -253
rect 127 -279 177 -253
rect 203 -279 253 -253
rect 279 -279 285 -253
rect -285 -285 285 -279
<< end >>
