magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1391 -2879 1391 2879
<< metal1 >>
rect -391 1873 391 1879
rect -391 1847 -385 1873
rect -359 1847 -323 1873
rect -297 1847 -261 1873
rect -235 1847 -199 1873
rect -173 1847 -137 1873
rect -111 1847 -75 1873
rect -49 1847 -13 1873
rect 13 1847 49 1873
rect 75 1847 111 1873
rect 137 1847 173 1873
rect 199 1847 235 1873
rect 261 1847 297 1873
rect 323 1847 359 1873
rect 385 1847 391 1873
rect -391 1811 391 1847
rect -391 1785 -385 1811
rect -359 1785 -323 1811
rect -297 1785 -261 1811
rect -235 1785 -199 1811
rect -173 1785 -137 1811
rect -111 1785 -75 1811
rect -49 1785 -13 1811
rect 13 1785 49 1811
rect 75 1785 111 1811
rect 137 1785 173 1811
rect 199 1785 235 1811
rect 261 1785 297 1811
rect 323 1785 359 1811
rect 385 1785 391 1811
rect -391 1749 391 1785
rect -391 1723 -385 1749
rect -359 1723 -323 1749
rect -297 1723 -261 1749
rect -235 1723 -199 1749
rect -173 1723 -137 1749
rect -111 1723 -75 1749
rect -49 1723 -13 1749
rect 13 1723 49 1749
rect 75 1723 111 1749
rect 137 1723 173 1749
rect 199 1723 235 1749
rect 261 1723 297 1749
rect 323 1723 359 1749
rect 385 1723 391 1749
rect -391 1687 391 1723
rect -391 1661 -385 1687
rect -359 1661 -323 1687
rect -297 1661 -261 1687
rect -235 1661 -199 1687
rect -173 1661 -137 1687
rect -111 1661 -75 1687
rect -49 1661 -13 1687
rect 13 1661 49 1687
rect 75 1661 111 1687
rect 137 1661 173 1687
rect 199 1661 235 1687
rect 261 1661 297 1687
rect 323 1661 359 1687
rect 385 1661 391 1687
rect -391 1625 391 1661
rect -391 1599 -385 1625
rect -359 1599 -323 1625
rect -297 1599 -261 1625
rect -235 1599 -199 1625
rect -173 1599 -137 1625
rect -111 1599 -75 1625
rect -49 1599 -13 1625
rect 13 1599 49 1625
rect 75 1599 111 1625
rect 137 1599 173 1625
rect 199 1599 235 1625
rect 261 1599 297 1625
rect 323 1599 359 1625
rect 385 1599 391 1625
rect -391 1563 391 1599
rect -391 1537 -385 1563
rect -359 1537 -323 1563
rect -297 1537 -261 1563
rect -235 1537 -199 1563
rect -173 1537 -137 1563
rect -111 1537 -75 1563
rect -49 1537 -13 1563
rect 13 1537 49 1563
rect 75 1537 111 1563
rect 137 1537 173 1563
rect 199 1537 235 1563
rect 261 1537 297 1563
rect 323 1537 359 1563
rect 385 1537 391 1563
rect -391 1501 391 1537
rect -391 1475 -385 1501
rect -359 1475 -323 1501
rect -297 1475 -261 1501
rect -235 1475 -199 1501
rect -173 1475 -137 1501
rect -111 1475 -75 1501
rect -49 1475 -13 1501
rect 13 1475 49 1501
rect 75 1475 111 1501
rect 137 1475 173 1501
rect 199 1475 235 1501
rect 261 1475 297 1501
rect 323 1475 359 1501
rect 385 1475 391 1501
rect -391 1439 391 1475
rect -391 1413 -385 1439
rect -359 1413 -323 1439
rect -297 1413 -261 1439
rect -235 1413 -199 1439
rect -173 1413 -137 1439
rect -111 1413 -75 1439
rect -49 1413 -13 1439
rect 13 1413 49 1439
rect 75 1413 111 1439
rect 137 1413 173 1439
rect 199 1413 235 1439
rect 261 1413 297 1439
rect 323 1413 359 1439
rect 385 1413 391 1439
rect -391 1377 391 1413
rect -391 1351 -385 1377
rect -359 1351 -323 1377
rect -297 1351 -261 1377
rect -235 1351 -199 1377
rect -173 1351 -137 1377
rect -111 1351 -75 1377
rect -49 1351 -13 1377
rect 13 1351 49 1377
rect 75 1351 111 1377
rect 137 1351 173 1377
rect 199 1351 235 1377
rect 261 1351 297 1377
rect 323 1351 359 1377
rect 385 1351 391 1377
rect -391 1315 391 1351
rect -391 1289 -385 1315
rect -359 1289 -323 1315
rect -297 1289 -261 1315
rect -235 1289 -199 1315
rect -173 1289 -137 1315
rect -111 1289 -75 1315
rect -49 1289 -13 1315
rect 13 1289 49 1315
rect 75 1289 111 1315
rect 137 1289 173 1315
rect 199 1289 235 1315
rect 261 1289 297 1315
rect 323 1289 359 1315
rect 385 1289 391 1315
rect -391 1253 391 1289
rect -391 1227 -385 1253
rect -359 1227 -323 1253
rect -297 1227 -261 1253
rect -235 1227 -199 1253
rect -173 1227 -137 1253
rect -111 1227 -75 1253
rect -49 1227 -13 1253
rect 13 1227 49 1253
rect 75 1227 111 1253
rect 137 1227 173 1253
rect 199 1227 235 1253
rect 261 1227 297 1253
rect 323 1227 359 1253
rect 385 1227 391 1253
rect -391 1191 391 1227
rect -391 1165 -385 1191
rect -359 1165 -323 1191
rect -297 1165 -261 1191
rect -235 1165 -199 1191
rect -173 1165 -137 1191
rect -111 1165 -75 1191
rect -49 1165 -13 1191
rect 13 1165 49 1191
rect 75 1165 111 1191
rect 137 1165 173 1191
rect 199 1165 235 1191
rect 261 1165 297 1191
rect 323 1165 359 1191
rect 385 1165 391 1191
rect -391 1129 391 1165
rect -391 1103 -385 1129
rect -359 1103 -323 1129
rect -297 1103 -261 1129
rect -235 1103 -199 1129
rect -173 1103 -137 1129
rect -111 1103 -75 1129
rect -49 1103 -13 1129
rect 13 1103 49 1129
rect 75 1103 111 1129
rect 137 1103 173 1129
rect 199 1103 235 1129
rect 261 1103 297 1129
rect 323 1103 359 1129
rect 385 1103 391 1129
rect -391 1067 391 1103
rect -391 1041 -385 1067
rect -359 1041 -323 1067
rect -297 1041 -261 1067
rect -235 1041 -199 1067
rect -173 1041 -137 1067
rect -111 1041 -75 1067
rect -49 1041 -13 1067
rect 13 1041 49 1067
rect 75 1041 111 1067
rect 137 1041 173 1067
rect 199 1041 235 1067
rect 261 1041 297 1067
rect 323 1041 359 1067
rect 385 1041 391 1067
rect -391 1005 391 1041
rect -391 979 -385 1005
rect -359 979 -323 1005
rect -297 979 -261 1005
rect -235 979 -199 1005
rect -173 979 -137 1005
rect -111 979 -75 1005
rect -49 979 -13 1005
rect 13 979 49 1005
rect 75 979 111 1005
rect 137 979 173 1005
rect 199 979 235 1005
rect 261 979 297 1005
rect 323 979 359 1005
rect 385 979 391 1005
rect -391 943 391 979
rect -391 917 -385 943
rect -359 917 -323 943
rect -297 917 -261 943
rect -235 917 -199 943
rect -173 917 -137 943
rect -111 917 -75 943
rect -49 917 -13 943
rect 13 917 49 943
rect 75 917 111 943
rect 137 917 173 943
rect 199 917 235 943
rect 261 917 297 943
rect 323 917 359 943
rect 385 917 391 943
rect -391 881 391 917
rect -391 855 -385 881
rect -359 855 -323 881
rect -297 855 -261 881
rect -235 855 -199 881
rect -173 855 -137 881
rect -111 855 -75 881
rect -49 855 -13 881
rect 13 855 49 881
rect 75 855 111 881
rect 137 855 173 881
rect 199 855 235 881
rect 261 855 297 881
rect 323 855 359 881
rect 385 855 391 881
rect -391 819 391 855
rect -391 793 -385 819
rect -359 793 -323 819
rect -297 793 -261 819
rect -235 793 -199 819
rect -173 793 -137 819
rect -111 793 -75 819
rect -49 793 -13 819
rect 13 793 49 819
rect 75 793 111 819
rect 137 793 173 819
rect 199 793 235 819
rect 261 793 297 819
rect 323 793 359 819
rect 385 793 391 819
rect -391 757 391 793
rect -391 731 -385 757
rect -359 731 -323 757
rect -297 731 -261 757
rect -235 731 -199 757
rect -173 731 -137 757
rect -111 731 -75 757
rect -49 731 -13 757
rect 13 731 49 757
rect 75 731 111 757
rect 137 731 173 757
rect 199 731 235 757
rect 261 731 297 757
rect 323 731 359 757
rect 385 731 391 757
rect -391 695 391 731
rect -391 669 -385 695
rect -359 669 -323 695
rect -297 669 -261 695
rect -235 669 -199 695
rect -173 669 -137 695
rect -111 669 -75 695
rect -49 669 -13 695
rect 13 669 49 695
rect 75 669 111 695
rect 137 669 173 695
rect 199 669 235 695
rect 261 669 297 695
rect 323 669 359 695
rect 385 669 391 695
rect -391 633 391 669
rect -391 607 -385 633
rect -359 607 -323 633
rect -297 607 -261 633
rect -235 607 -199 633
rect -173 607 -137 633
rect -111 607 -75 633
rect -49 607 -13 633
rect 13 607 49 633
rect 75 607 111 633
rect 137 607 173 633
rect 199 607 235 633
rect 261 607 297 633
rect 323 607 359 633
rect 385 607 391 633
rect -391 571 391 607
rect -391 545 -385 571
rect -359 545 -323 571
rect -297 545 -261 571
rect -235 545 -199 571
rect -173 545 -137 571
rect -111 545 -75 571
rect -49 545 -13 571
rect 13 545 49 571
rect 75 545 111 571
rect 137 545 173 571
rect 199 545 235 571
rect 261 545 297 571
rect 323 545 359 571
rect 385 545 391 571
rect -391 509 391 545
rect -391 483 -385 509
rect -359 483 -323 509
rect -297 483 -261 509
rect -235 483 -199 509
rect -173 483 -137 509
rect -111 483 -75 509
rect -49 483 -13 509
rect 13 483 49 509
rect 75 483 111 509
rect 137 483 173 509
rect 199 483 235 509
rect 261 483 297 509
rect 323 483 359 509
rect 385 483 391 509
rect -391 447 391 483
rect -391 421 -385 447
rect -359 421 -323 447
rect -297 421 -261 447
rect -235 421 -199 447
rect -173 421 -137 447
rect -111 421 -75 447
rect -49 421 -13 447
rect 13 421 49 447
rect 75 421 111 447
rect 137 421 173 447
rect 199 421 235 447
rect 261 421 297 447
rect 323 421 359 447
rect 385 421 391 447
rect -391 385 391 421
rect -391 359 -385 385
rect -359 359 -323 385
rect -297 359 -261 385
rect -235 359 -199 385
rect -173 359 -137 385
rect -111 359 -75 385
rect -49 359 -13 385
rect 13 359 49 385
rect 75 359 111 385
rect 137 359 173 385
rect 199 359 235 385
rect 261 359 297 385
rect 323 359 359 385
rect 385 359 391 385
rect -391 323 391 359
rect -391 297 -385 323
rect -359 297 -323 323
rect -297 297 -261 323
rect -235 297 -199 323
rect -173 297 -137 323
rect -111 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 111 323
rect 137 297 173 323
rect 199 297 235 323
rect 261 297 297 323
rect 323 297 359 323
rect 385 297 391 323
rect -391 261 391 297
rect -391 235 -385 261
rect -359 235 -323 261
rect -297 235 -261 261
rect -235 235 -199 261
rect -173 235 -137 261
rect -111 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 111 261
rect 137 235 173 261
rect 199 235 235 261
rect 261 235 297 261
rect 323 235 359 261
rect 385 235 391 261
rect -391 199 391 235
rect -391 173 -385 199
rect -359 173 -323 199
rect -297 173 -261 199
rect -235 173 -199 199
rect -173 173 -137 199
rect -111 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 111 199
rect 137 173 173 199
rect 199 173 235 199
rect 261 173 297 199
rect 323 173 359 199
rect 385 173 391 199
rect -391 137 391 173
rect -391 111 -385 137
rect -359 111 -323 137
rect -297 111 -261 137
rect -235 111 -199 137
rect -173 111 -137 137
rect -111 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 111 137
rect 137 111 173 137
rect 199 111 235 137
rect 261 111 297 137
rect 323 111 359 137
rect 385 111 391 137
rect -391 75 391 111
rect -391 49 -385 75
rect -359 49 -323 75
rect -297 49 -261 75
rect -235 49 -199 75
rect -173 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 173 75
rect 199 49 235 75
rect 261 49 297 75
rect 323 49 359 75
rect 385 49 391 75
rect -391 13 391 49
rect -391 -13 -385 13
rect -359 -13 -323 13
rect -297 -13 -261 13
rect -235 -13 -199 13
rect -173 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 173 13
rect 199 -13 235 13
rect 261 -13 297 13
rect 323 -13 359 13
rect 385 -13 391 13
rect -391 -49 391 -13
rect -391 -75 -385 -49
rect -359 -75 -323 -49
rect -297 -75 -261 -49
rect -235 -75 -199 -49
rect -173 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 173 -49
rect 199 -75 235 -49
rect 261 -75 297 -49
rect 323 -75 359 -49
rect 385 -75 391 -49
rect -391 -111 391 -75
rect -391 -137 -385 -111
rect -359 -137 -323 -111
rect -297 -137 -261 -111
rect -235 -137 -199 -111
rect -173 -137 -137 -111
rect -111 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 111 -111
rect 137 -137 173 -111
rect 199 -137 235 -111
rect 261 -137 297 -111
rect 323 -137 359 -111
rect 385 -137 391 -111
rect -391 -173 391 -137
rect -391 -199 -385 -173
rect -359 -199 -323 -173
rect -297 -199 -261 -173
rect -235 -199 -199 -173
rect -173 -199 -137 -173
rect -111 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 111 -173
rect 137 -199 173 -173
rect 199 -199 235 -173
rect 261 -199 297 -173
rect 323 -199 359 -173
rect 385 -199 391 -173
rect -391 -235 391 -199
rect -391 -261 -385 -235
rect -359 -261 -323 -235
rect -297 -261 -261 -235
rect -235 -261 -199 -235
rect -173 -261 -137 -235
rect -111 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 111 -235
rect 137 -261 173 -235
rect 199 -261 235 -235
rect 261 -261 297 -235
rect 323 -261 359 -235
rect 385 -261 391 -235
rect -391 -297 391 -261
rect -391 -323 -385 -297
rect -359 -323 -323 -297
rect -297 -323 -261 -297
rect -235 -323 -199 -297
rect -173 -323 -137 -297
rect -111 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 111 -297
rect 137 -323 173 -297
rect 199 -323 235 -297
rect 261 -323 297 -297
rect 323 -323 359 -297
rect 385 -323 391 -297
rect -391 -359 391 -323
rect -391 -385 -385 -359
rect -359 -385 -323 -359
rect -297 -385 -261 -359
rect -235 -385 -199 -359
rect -173 -385 -137 -359
rect -111 -385 -75 -359
rect -49 -385 -13 -359
rect 13 -385 49 -359
rect 75 -385 111 -359
rect 137 -385 173 -359
rect 199 -385 235 -359
rect 261 -385 297 -359
rect 323 -385 359 -359
rect 385 -385 391 -359
rect -391 -421 391 -385
rect -391 -447 -385 -421
rect -359 -447 -323 -421
rect -297 -447 -261 -421
rect -235 -447 -199 -421
rect -173 -447 -137 -421
rect -111 -447 -75 -421
rect -49 -447 -13 -421
rect 13 -447 49 -421
rect 75 -447 111 -421
rect 137 -447 173 -421
rect 199 -447 235 -421
rect 261 -447 297 -421
rect 323 -447 359 -421
rect 385 -447 391 -421
rect -391 -483 391 -447
rect -391 -509 -385 -483
rect -359 -509 -323 -483
rect -297 -509 -261 -483
rect -235 -509 -199 -483
rect -173 -509 -137 -483
rect -111 -509 -75 -483
rect -49 -509 -13 -483
rect 13 -509 49 -483
rect 75 -509 111 -483
rect 137 -509 173 -483
rect 199 -509 235 -483
rect 261 -509 297 -483
rect 323 -509 359 -483
rect 385 -509 391 -483
rect -391 -545 391 -509
rect -391 -571 -385 -545
rect -359 -571 -323 -545
rect -297 -571 -261 -545
rect -235 -571 -199 -545
rect -173 -571 -137 -545
rect -111 -571 -75 -545
rect -49 -571 -13 -545
rect 13 -571 49 -545
rect 75 -571 111 -545
rect 137 -571 173 -545
rect 199 -571 235 -545
rect 261 -571 297 -545
rect 323 -571 359 -545
rect 385 -571 391 -545
rect -391 -607 391 -571
rect -391 -633 -385 -607
rect -359 -633 -323 -607
rect -297 -633 -261 -607
rect -235 -633 -199 -607
rect -173 -633 -137 -607
rect -111 -633 -75 -607
rect -49 -633 -13 -607
rect 13 -633 49 -607
rect 75 -633 111 -607
rect 137 -633 173 -607
rect 199 -633 235 -607
rect 261 -633 297 -607
rect 323 -633 359 -607
rect 385 -633 391 -607
rect -391 -669 391 -633
rect -391 -695 -385 -669
rect -359 -695 -323 -669
rect -297 -695 -261 -669
rect -235 -695 -199 -669
rect -173 -695 -137 -669
rect -111 -695 -75 -669
rect -49 -695 -13 -669
rect 13 -695 49 -669
rect 75 -695 111 -669
rect 137 -695 173 -669
rect 199 -695 235 -669
rect 261 -695 297 -669
rect 323 -695 359 -669
rect 385 -695 391 -669
rect -391 -731 391 -695
rect -391 -757 -385 -731
rect -359 -757 -323 -731
rect -297 -757 -261 -731
rect -235 -757 -199 -731
rect -173 -757 -137 -731
rect -111 -757 -75 -731
rect -49 -757 -13 -731
rect 13 -757 49 -731
rect 75 -757 111 -731
rect 137 -757 173 -731
rect 199 -757 235 -731
rect 261 -757 297 -731
rect 323 -757 359 -731
rect 385 -757 391 -731
rect -391 -793 391 -757
rect -391 -819 -385 -793
rect -359 -819 -323 -793
rect -297 -819 -261 -793
rect -235 -819 -199 -793
rect -173 -819 -137 -793
rect -111 -819 -75 -793
rect -49 -819 -13 -793
rect 13 -819 49 -793
rect 75 -819 111 -793
rect 137 -819 173 -793
rect 199 -819 235 -793
rect 261 -819 297 -793
rect 323 -819 359 -793
rect 385 -819 391 -793
rect -391 -855 391 -819
rect -391 -881 -385 -855
rect -359 -881 -323 -855
rect -297 -881 -261 -855
rect -235 -881 -199 -855
rect -173 -881 -137 -855
rect -111 -881 -75 -855
rect -49 -881 -13 -855
rect 13 -881 49 -855
rect 75 -881 111 -855
rect 137 -881 173 -855
rect 199 -881 235 -855
rect 261 -881 297 -855
rect 323 -881 359 -855
rect 385 -881 391 -855
rect -391 -917 391 -881
rect -391 -943 -385 -917
rect -359 -943 -323 -917
rect -297 -943 -261 -917
rect -235 -943 -199 -917
rect -173 -943 -137 -917
rect -111 -943 -75 -917
rect -49 -943 -13 -917
rect 13 -943 49 -917
rect 75 -943 111 -917
rect 137 -943 173 -917
rect 199 -943 235 -917
rect 261 -943 297 -917
rect 323 -943 359 -917
rect 385 -943 391 -917
rect -391 -979 391 -943
rect -391 -1005 -385 -979
rect -359 -1005 -323 -979
rect -297 -1005 -261 -979
rect -235 -1005 -199 -979
rect -173 -1005 -137 -979
rect -111 -1005 -75 -979
rect -49 -1005 -13 -979
rect 13 -1005 49 -979
rect 75 -1005 111 -979
rect 137 -1005 173 -979
rect 199 -1005 235 -979
rect 261 -1005 297 -979
rect 323 -1005 359 -979
rect 385 -1005 391 -979
rect -391 -1041 391 -1005
rect -391 -1067 -385 -1041
rect -359 -1067 -323 -1041
rect -297 -1067 -261 -1041
rect -235 -1067 -199 -1041
rect -173 -1067 -137 -1041
rect -111 -1067 -75 -1041
rect -49 -1067 -13 -1041
rect 13 -1067 49 -1041
rect 75 -1067 111 -1041
rect 137 -1067 173 -1041
rect 199 -1067 235 -1041
rect 261 -1067 297 -1041
rect 323 -1067 359 -1041
rect 385 -1067 391 -1041
rect -391 -1103 391 -1067
rect -391 -1129 -385 -1103
rect -359 -1129 -323 -1103
rect -297 -1129 -261 -1103
rect -235 -1129 -199 -1103
rect -173 -1129 -137 -1103
rect -111 -1129 -75 -1103
rect -49 -1129 -13 -1103
rect 13 -1129 49 -1103
rect 75 -1129 111 -1103
rect 137 -1129 173 -1103
rect 199 -1129 235 -1103
rect 261 -1129 297 -1103
rect 323 -1129 359 -1103
rect 385 -1129 391 -1103
rect -391 -1165 391 -1129
rect -391 -1191 -385 -1165
rect -359 -1191 -323 -1165
rect -297 -1191 -261 -1165
rect -235 -1191 -199 -1165
rect -173 -1191 -137 -1165
rect -111 -1191 -75 -1165
rect -49 -1191 -13 -1165
rect 13 -1191 49 -1165
rect 75 -1191 111 -1165
rect 137 -1191 173 -1165
rect 199 -1191 235 -1165
rect 261 -1191 297 -1165
rect 323 -1191 359 -1165
rect 385 -1191 391 -1165
rect -391 -1227 391 -1191
rect -391 -1253 -385 -1227
rect -359 -1253 -323 -1227
rect -297 -1253 -261 -1227
rect -235 -1253 -199 -1227
rect -173 -1253 -137 -1227
rect -111 -1253 -75 -1227
rect -49 -1253 -13 -1227
rect 13 -1253 49 -1227
rect 75 -1253 111 -1227
rect 137 -1253 173 -1227
rect 199 -1253 235 -1227
rect 261 -1253 297 -1227
rect 323 -1253 359 -1227
rect 385 -1253 391 -1227
rect -391 -1289 391 -1253
rect -391 -1315 -385 -1289
rect -359 -1315 -323 -1289
rect -297 -1315 -261 -1289
rect -235 -1315 -199 -1289
rect -173 -1315 -137 -1289
rect -111 -1315 -75 -1289
rect -49 -1315 -13 -1289
rect 13 -1315 49 -1289
rect 75 -1315 111 -1289
rect 137 -1315 173 -1289
rect 199 -1315 235 -1289
rect 261 -1315 297 -1289
rect 323 -1315 359 -1289
rect 385 -1315 391 -1289
rect -391 -1351 391 -1315
rect -391 -1377 -385 -1351
rect -359 -1377 -323 -1351
rect -297 -1377 -261 -1351
rect -235 -1377 -199 -1351
rect -173 -1377 -137 -1351
rect -111 -1377 -75 -1351
rect -49 -1377 -13 -1351
rect 13 -1377 49 -1351
rect 75 -1377 111 -1351
rect 137 -1377 173 -1351
rect 199 -1377 235 -1351
rect 261 -1377 297 -1351
rect 323 -1377 359 -1351
rect 385 -1377 391 -1351
rect -391 -1413 391 -1377
rect -391 -1439 -385 -1413
rect -359 -1439 -323 -1413
rect -297 -1439 -261 -1413
rect -235 -1439 -199 -1413
rect -173 -1439 -137 -1413
rect -111 -1439 -75 -1413
rect -49 -1439 -13 -1413
rect 13 -1439 49 -1413
rect 75 -1439 111 -1413
rect 137 -1439 173 -1413
rect 199 -1439 235 -1413
rect 261 -1439 297 -1413
rect 323 -1439 359 -1413
rect 385 -1439 391 -1413
rect -391 -1475 391 -1439
rect -391 -1501 -385 -1475
rect -359 -1501 -323 -1475
rect -297 -1501 -261 -1475
rect -235 -1501 -199 -1475
rect -173 -1501 -137 -1475
rect -111 -1501 -75 -1475
rect -49 -1501 -13 -1475
rect 13 -1501 49 -1475
rect 75 -1501 111 -1475
rect 137 -1501 173 -1475
rect 199 -1501 235 -1475
rect 261 -1501 297 -1475
rect 323 -1501 359 -1475
rect 385 -1501 391 -1475
rect -391 -1537 391 -1501
rect -391 -1563 -385 -1537
rect -359 -1563 -323 -1537
rect -297 -1563 -261 -1537
rect -235 -1563 -199 -1537
rect -173 -1563 -137 -1537
rect -111 -1563 -75 -1537
rect -49 -1563 -13 -1537
rect 13 -1563 49 -1537
rect 75 -1563 111 -1537
rect 137 -1563 173 -1537
rect 199 -1563 235 -1537
rect 261 -1563 297 -1537
rect 323 -1563 359 -1537
rect 385 -1563 391 -1537
rect -391 -1599 391 -1563
rect -391 -1625 -385 -1599
rect -359 -1625 -323 -1599
rect -297 -1625 -261 -1599
rect -235 -1625 -199 -1599
rect -173 -1625 -137 -1599
rect -111 -1625 -75 -1599
rect -49 -1625 -13 -1599
rect 13 -1625 49 -1599
rect 75 -1625 111 -1599
rect 137 -1625 173 -1599
rect 199 -1625 235 -1599
rect 261 -1625 297 -1599
rect 323 -1625 359 -1599
rect 385 -1625 391 -1599
rect -391 -1661 391 -1625
rect -391 -1687 -385 -1661
rect -359 -1687 -323 -1661
rect -297 -1687 -261 -1661
rect -235 -1687 -199 -1661
rect -173 -1687 -137 -1661
rect -111 -1687 -75 -1661
rect -49 -1687 -13 -1661
rect 13 -1687 49 -1661
rect 75 -1687 111 -1661
rect 137 -1687 173 -1661
rect 199 -1687 235 -1661
rect 261 -1687 297 -1661
rect 323 -1687 359 -1661
rect 385 -1687 391 -1661
rect -391 -1723 391 -1687
rect -391 -1749 -385 -1723
rect -359 -1749 -323 -1723
rect -297 -1749 -261 -1723
rect -235 -1749 -199 -1723
rect -173 -1749 -137 -1723
rect -111 -1749 -75 -1723
rect -49 -1749 -13 -1723
rect 13 -1749 49 -1723
rect 75 -1749 111 -1723
rect 137 -1749 173 -1723
rect 199 -1749 235 -1723
rect 261 -1749 297 -1723
rect 323 -1749 359 -1723
rect 385 -1749 391 -1723
rect -391 -1785 391 -1749
rect -391 -1811 -385 -1785
rect -359 -1811 -323 -1785
rect -297 -1811 -261 -1785
rect -235 -1811 -199 -1785
rect -173 -1811 -137 -1785
rect -111 -1811 -75 -1785
rect -49 -1811 -13 -1785
rect 13 -1811 49 -1785
rect 75 -1811 111 -1785
rect 137 -1811 173 -1785
rect 199 -1811 235 -1785
rect 261 -1811 297 -1785
rect 323 -1811 359 -1785
rect 385 -1811 391 -1785
rect -391 -1847 391 -1811
rect -391 -1873 -385 -1847
rect -359 -1873 -323 -1847
rect -297 -1873 -261 -1847
rect -235 -1873 -199 -1847
rect -173 -1873 -137 -1847
rect -111 -1873 -75 -1847
rect -49 -1873 -13 -1847
rect 13 -1873 49 -1847
rect 75 -1873 111 -1847
rect 137 -1873 173 -1847
rect 199 -1873 235 -1847
rect 261 -1873 297 -1847
rect 323 -1873 359 -1847
rect 385 -1873 391 -1847
rect -391 -1879 391 -1873
<< via1 >>
rect -385 1847 -359 1873
rect -323 1847 -297 1873
rect -261 1847 -235 1873
rect -199 1847 -173 1873
rect -137 1847 -111 1873
rect -75 1847 -49 1873
rect -13 1847 13 1873
rect 49 1847 75 1873
rect 111 1847 137 1873
rect 173 1847 199 1873
rect 235 1847 261 1873
rect 297 1847 323 1873
rect 359 1847 385 1873
rect -385 1785 -359 1811
rect -323 1785 -297 1811
rect -261 1785 -235 1811
rect -199 1785 -173 1811
rect -137 1785 -111 1811
rect -75 1785 -49 1811
rect -13 1785 13 1811
rect 49 1785 75 1811
rect 111 1785 137 1811
rect 173 1785 199 1811
rect 235 1785 261 1811
rect 297 1785 323 1811
rect 359 1785 385 1811
rect -385 1723 -359 1749
rect -323 1723 -297 1749
rect -261 1723 -235 1749
rect -199 1723 -173 1749
rect -137 1723 -111 1749
rect -75 1723 -49 1749
rect -13 1723 13 1749
rect 49 1723 75 1749
rect 111 1723 137 1749
rect 173 1723 199 1749
rect 235 1723 261 1749
rect 297 1723 323 1749
rect 359 1723 385 1749
rect -385 1661 -359 1687
rect -323 1661 -297 1687
rect -261 1661 -235 1687
rect -199 1661 -173 1687
rect -137 1661 -111 1687
rect -75 1661 -49 1687
rect -13 1661 13 1687
rect 49 1661 75 1687
rect 111 1661 137 1687
rect 173 1661 199 1687
rect 235 1661 261 1687
rect 297 1661 323 1687
rect 359 1661 385 1687
rect -385 1599 -359 1625
rect -323 1599 -297 1625
rect -261 1599 -235 1625
rect -199 1599 -173 1625
rect -137 1599 -111 1625
rect -75 1599 -49 1625
rect -13 1599 13 1625
rect 49 1599 75 1625
rect 111 1599 137 1625
rect 173 1599 199 1625
rect 235 1599 261 1625
rect 297 1599 323 1625
rect 359 1599 385 1625
rect -385 1537 -359 1563
rect -323 1537 -297 1563
rect -261 1537 -235 1563
rect -199 1537 -173 1563
rect -137 1537 -111 1563
rect -75 1537 -49 1563
rect -13 1537 13 1563
rect 49 1537 75 1563
rect 111 1537 137 1563
rect 173 1537 199 1563
rect 235 1537 261 1563
rect 297 1537 323 1563
rect 359 1537 385 1563
rect -385 1475 -359 1501
rect -323 1475 -297 1501
rect -261 1475 -235 1501
rect -199 1475 -173 1501
rect -137 1475 -111 1501
rect -75 1475 -49 1501
rect -13 1475 13 1501
rect 49 1475 75 1501
rect 111 1475 137 1501
rect 173 1475 199 1501
rect 235 1475 261 1501
rect 297 1475 323 1501
rect 359 1475 385 1501
rect -385 1413 -359 1439
rect -323 1413 -297 1439
rect -261 1413 -235 1439
rect -199 1413 -173 1439
rect -137 1413 -111 1439
rect -75 1413 -49 1439
rect -13 1413 13 1439
rect 49 1413 75 1439
rect 111 1413 137 1439
rect 173 1413 199 1439
rect 235 1413 261 1439
rect 297 1413 323 1439
rect 359 1413 385 1439
rect -385 1351 -359 1377
rect -323 1351 -297 1377
rect -261 1351 -235 1377
rect -199 1351 -173 1377
rect -137 1351 -111 1377
rect -75 1351 -49 1377
rect -13 1351 13 1377
rect 49 1351 75 1377
rect 111 1351 137 1377
rect 173 1351 199 1377
rect 235 1351 261 1377
rect 297 1351 323 1377
rect 359 1351 385 1377
rect -385 1289 -359 1315
rect -323 1289 -297 1315
rect -261 1289 -235 1315
rect -199 1289 -173 1315
rect -137 1289 -111 1315
rect -75 1289 -49 1315
rect -13 1289 13 1315
rect 49 1289 75 1315
rect 111 1289 137 1315
rect 173 1289 199 1315
rect 235 1289 261 1315
rect 297 1289 323 1315
rect 359 1289 385 1315
rect -385 1227 -359 1253
rect -323 1227 -297 1253
rect -261 1227 -235 1253
rect -199 1227 -173 1253
rect -137 1227 -111 1253
rect -75 1227 -49 1253
rect -13 1227 13 1253
rect 49 1227 75 1253
rect 111 1227 137 1253
rect 173 1227 199 1253
rect 235 1227 261 1253
rect 297 1227 323 1253
rect 359 1227 385 1253
rect -385 1165 -359 1191
rect -323 1165 -297 1191
rect -261 1165 -235 1191
rect -199 1165 -173 1191
rect -137 1165 -111 1191
rect -75 1165 -49 1191
rect -13 1165 13 1191
rect 49 1165 75 1191
rect 111 1165 137 1191
rect 173 1165 199 1191
rect 235 1165 261 1191
rect 297 1165 323 1191
rect 359 1165 385 1191
rect -385 1103 -359 1129
rect -323 1103 -297 1129
rect -261 1103 -235 1129
rect -199 1103 -173 1129
rect -137 1103 -111 1129
rect -75 1103 -49 1129
rect -13 1103 13 1129
rect 49 1103 75 1129
rect 111 1103 137 1129
rect 173 1103 199 1129
rect 235 1103 261 1129
rect 297 1103 323 1129
rect 359 1103 385 1129
rect -385 1041 -359 1067
rect -323 1041 -297 1067
rect -261 1041 -235 1067
rect -199 1041 -173 1067
rect -137 1041 -111 1067
rect -75 1041 -49 1067
rect -13 1041 13 1067
rect 49 1041 75 1067
rect 111 1041 137 1067
rect 173 1041 199 1067
rect 235 1041 261 1067
rect 297 1041 323 1067
rect 359 1041 385 1067
rect -385 979 -359 1005
rect -323 979 -297 1005
rect -261 979 -235 1005
rect -199 979 -173 1005
rect -137 979 -111 1005
rect -75 979 -49 1005
rect -13 979 13 1005
rect 49 979 75 1005
rect 111 979 137 1005
rect 173 979 199 1005
rect 235 979 261 1005
rect 297 979 323 1005
rect 359 979 385 1005
rect -385 917 -359 943
rect -323 917 -297 943
rect -261 917 -235 943
rect -199 917 -173 943
rect -137 917 -111 943
rect -75 917 -49 943
rect -13 917 13 943
rect 49 917 75 943
rect 111 917 137 943
rect 173 917 199 943
rect 235 917 261 943
rect 297 917 323 943
rect 359 917 385 943
rect -385 855 -359 881
rect -323 855 -297 881
rect -261 855 -235 881
rect -199 855 -173 881
rect -137 855 -111 881
rect -75 855 -49 881
rect -13 855 13 881
rect 49 855 75 881
rect 111 855 137 881
rect 173 855 199 881
rect 235 855 261 881
rect 297 855 323 881
rect 359 855 385 881
rect -385 793 -359 819
rect -323 793 -297 819
rect -261 793 -235 819
rect -199 793 -173 819
rect -137 793 -111 819
rect -75 793 -49 819
rect -13 793 13 819
rect 49 793 75 819
rect 111 793 137 819
rect 173 793 199 819
rect 235 793 261 819
rect 297 793 323 819
rect 359 793 385 819
rect -385 731 -359 757
rect -323 731 -297 757
rect -261 731 -235 757
rect -199 731 -173 757
rect -137 731 -111 757
rect -75 731 -49 757
rect -13 731 13 757
rect 49 731 75 757
rect 111 731 137 757
rect 173 731 199 757
rect 235 731 261 757
rect 297 731 323 757
rect 359 731 385 757
rect -385 669 -359 695
rect -323 669 -297 695
rect -261 669 -235 695
rect -199 669 -173 695
rect -137 669 -111 695
rect -75 669 -49 695
rect -13 669 13 695
rect 49 669 75 695
rect 111 669 137 695
rect 173 669 199 695
rect 235 669 261 695
rect 297 669 323 695
rect 359 669 385 695
rect -385 607 -359 633
rect -323 607 -297 633
rect -261 607 -235 633
rect -199 607 -173 633
rect -137 607 -111 633
rect -75 607 -49 633
rect -13 607 13 633
rect 49 607 75 633
rect 111 607 137 633
rect 173 607 199 633
rect 235 607 261 633
rect 297 607 323 633
rect 359 607 385 633
rect -385 545 -359 571
rect -323 545 -297 571
rect -261 545 -235 571
rect -199 545 -173 571
rect -137 545 -111 571
rect -75 545 -49 571
rect -13 545 13 571
rect 49 545 75 571
rect 111 545 137 571
rect 173 545 199 571
rect 235 545 261 571
rect 297 545 323 571
rect 359 545 385 571
rect -385 483 -359 509
rect -323 483 -297 509
rect -261 483 -235 509
rect -199 483 -173 509
rect -137 483 -111 509
rect -75 483 -49 509
rect -13 483 13 509
rect 49 483 75 509
rect 111 483 137 509
rect 173 483 199 509
rect 235 483 261 509
rect 297 483 323 509
rect 359 483 385 509
rect -385 421 -359 447
rect -323 421 -297 447
rect -261 421 -235 447
rect -199 421 -173 447
rect -137 421 -111 447
rect -75 421 -49 447
rect -13 421 13 447
rect 49 421 75 447
rect 111 421 137 447
rect 173 421 199 447
rect 235 421 261 447
rect 297 421 323 447
rect 359 421 385 447
rect -385 359 -359 385
rect -323 359 -297 385
rect -261 359 -235 385
rect -199 359 -173 385
rect -137 359 -111 385
rect -75 359 -49 385
rect -13 359 13 385
rect 49 359 75 385
rect 111 359 137 385
rect 173 359 199 385
rect 235 359 261 385
rect 297 359 323 385
rect 359 359 385 385
rect -385 297 -359 323
rect -323 297 -297 323
rect -261 297 -235 323
rect -199 297 -173 323
rect -137 297 -111 323
rect -75 297 -49 323
rect -13 297 13 323
rect 49 297 75 323
rect 111 297 137 323
rect 173 297 199 323
rect 235 297 261 323
rect 297 297 323 323
rect 359 297 385 323
rect -385 235 -359 261
rect -323 235 -297 261
rect -261 235 -235 261
rect -199 235 -173 261
rect -137 235 -111 261
rect -75 235 -49 261
rect -13 235 13 261
rect 49 235 75 261
rect 111 235 137 261
rect 173 235 199 261
rect 235 235 261 261
rect 297 235 323 261
rect 359 235 385 261
rect -385 173 -359 199
rect -323 173 -297 199
rect -261 173 -235 199
rect -199 173 -173 199
rect -137 173 -111 199
rect -75 173 -49 199
rect -13 173 13 199
rect 49 173 75 199
rect 111 173 137 199
rect 173 173 199 199
rect 235 173 261 199
rect 297 173 323 199
rect 359 173 385 199
rect -385 111 -359 137
rect -323 111 -297 137
rect -261 111 -235 137
rect -199 111 -173 137
rect -137 111 -111 137
rect -75 111 -49 137
rect -13 111 13 137
rect 49 111 75 137
rect 111 111 137 137
rect 173 111 199 137
rect 235 111 261 137
rect 297 111 323 137
rect 359 111 385 137
rect -385 49 -359 75
rect -323 49 -297 75
rect -261 49 -235 75
rect -199 49 -173 75
rect -137 49 -111 75
rect -75 49 -49 75
rect -13 49 13 75
rect 49 49 75 75
rect 111 49 137 75
rect 173 49 199 75
rect 235 49 261 75
rect 297 49 323 75
rect 359 49 385 75
rect -385 -13 -359 13
rect -323 -13 -297 13
rect -261 -13 -235 13
rect -199 -13 -173 13
rect -137 -13 -111 13
rect -75 -13 -49 13
rect -13 -13 13 13
rect 49 -13 75 13
rect 111 -13 137 13
rect 173 -13 199 13
rect 235 -13 261 13
rect 297 -13 323 13
rect 359 -13 385 13
rect -385 -75 -359 -49
rect -323 -75 -297 -49
rect -261 -75 -235 -49
rect -199 -75 -173 -49
rect -137 -75 -111 -49
rect -75 -75 -49 -49
rect -13 -75 13 -49
rect 49 -75 75 -49
rect 111 -75 137 -49
rect 173 -75 199 -49
rect 235 -75 261 -49
rect 297 -75 323 -49
rect 359 -75 385 -49
rect -385 -137 -359 -111
rect -323 -137 -297 -111
rect -261 -137 -235 -111
rect -199 -137 -173 -111
rect -137 -137 -111 -111
rect -75 -137 -49 -111
rect -13 -137 13 -111
rect 49 -137 75 -111
rect 111 -137 137 -111
rect 173 -137 199 -111
rect 235 -137 261 -111
rect 297 -137 323 -111
rect 359 -137 385 -111
rect -385 -199 -359 -173
rect -323 -199 -297 -173
rect -261 -199 -235 -173
rect -199 -199 -173 -173
rect -137 -199 -111 -173
rect -75 -199 -49 -173
rect -13 -199 13 -173
rect 49 -199 75 -173
rect 111 -199 137 -173
rect 173 -199 199 -173
rect 235 -199 261 -173
rect 297 -199 323 -173
rect 359 -199 385 -173
rect -385 -261 -359 -235
rect -323 -261 -297 -235
rect -261 -261 -235 -235
rect -199 -261 -173 -235
rect -137 -261 -111 -235
rect -75 -261 -49 -235
rect -13 -261 13 -235
rect 49 -261 75 -235
rect 111 -261 137 -235
rect 173 -261 199 -235
rect 235 -261 261 -235
rect 297 -261 323 -235
rect 359 -261 385 -235
rect -385 -323 -359 -297
rect -323 -323 -297 -297
rect -261 -323 -235 -297
rect -199 -323 -173 -297
rect -137 -323 -111 -297
rect -75 -323 -49 -297
rect -13 -323 13 -297
rect 49 -323 75 -297
rect 111 -323 137 -297
rect 173 -323 199 -297
rect 235 -323 261 -297
rect 297 -323 323 -297
rect 359 -323 385 -297
rect -385 -385 -359 -359
rect -323 -385 -297 -359
rect -261 -385 -235 -359
rect -199 -385 -173 -359
rect -137 -385 -111 -359
rect -75 -385 -49 -359
rect -13 -385 13 -359
rect 49 -385 75 -359
rect 111 -385 137 -359
rect 173 -385 199 -359
rect 235 -385 261 -359
rect 297 -385 323 -359
rect 359 -385 385 -359
rect -385 -447 -359 -421
rect -323 -447 -297 -421
rect -261 -447 -235 -421
rect -199 -447 -173 -421
rect -137 -447 -111 -421
rect -75 -447 -49 -421
rect -13 -447 13 -421
rect 49 -447 75 -421
rect 111 -447 137 -421
rect 173 -447 199 -421
rect 235 -447 261 -421
rect 297 -447 323 -421
rect 359 -447 385 -421
rect -385 -509 -359 -483
rect -323 -509 -297 -483
rect -261 -509 -235 -483
rect -199 -509 -173 -483
rect -137 -509 -111 -483
rect -75 -509 -49 -483
rect -13 -509 13 -483
rect 49 -509 75 -483
rect 111 -509 137 -483
rect 173 -509 199 -483
rect 235 -509 261 -483
rect 297 -509 323 -483
rect 359 -509 385 -483
rect -385 -571 -359 -545
rect -323 -571 -297 -545
rect -261 -571 -235 -545
rect -199 -571 -173 -545
rect -137 -571 -111 -545
rect -75 -571 -49 -545
rect -13 -571 13 -545
rect 49 -571 75 -545
rect 111 -571 137 -545
rect 173 -571 199 -545
rect 235 -571 261 -545
rect 297 -571 323 -545
rect 359 -571 385 -545
rect -385 -633 -359 -607
rect -323 -633 -297 -607
rect -261 -633 -235 -607
rect -199 -633 -173 -607
rect -137 -633 -111 -607
rect -75 -633 -49 -607
rect -13 -633 13 -607
rect 49 -633 75 -607
rect 111 -633 137 -607
rect 173 -633 199 -607
rect 235 -633 261 -607
rect 297 -633 323 -607
rect 359 -633 385 -607
rect -385 -695 -359 -669
rect -323 -695 -297 -669
rect -261 -695 -235 -669
rect -199 -695 -173 -669
rect -137 -695 -111 -669
rect -75 -695 -49 -669
rect -13 -695 13 -669
rect 49 -695 75 -669
rect 111 -695 137 -669
rect 173 -695 199 -669
rect 235 -695 261 -669
rect 297 -695 323 -669
rect 359 -695 385 -669
rect -385 -757 -359 -731
rect -323 -757 -297 -731
rect -261 -757 -235 -731
rect -199 -757 -173 -731
rect -137 -757 -111 -731
rect -75 -757 -49 -731
rect -13 -757 13 -731
rect 49 -757 75 -731
rect 111 -757 137 -731
rect 173 -757 199 -731
rect 235 -757 261 -731
rect 297 -757 323 -731
rect 359 -757 385 -731
rect -385 -819 -359 -793
rect -323 -819 -297 -793
rect -261 -819 -235 -793
rect -199 -819 -173 -793
rect -137 -819 -111 -793
rect -75 -819 -49 -793
rect -13 -819 13 -793
rect 49 -819 75 -793
rect 111 -819 137 -793
rect 173 -819 199 -793
rect 235 -819 261 -793
rect 297 -819 323 -793
rect 359 -819 385 -793
rect -385 -881 -359 -855
rect -323 -881 -297 -855
rect -261 -881 -235 -855
rect -199 -881 -173 -855
rect -137 -881 -111 -855
rect -75 -881 -49 -855
rect -13 -881 13 -855
rect 49 -881 75 -855
rect 111 -881 137 -855
rect 173 -881 199 -855
rect 235 -881 261 -855
rect 297 -881 323 -855
rect 359 -881 385 -855
rect -385 -943 -359 -917
rect -323 -943 -297 -917
rect -261 -943 -235 -917
rect -199 -943 -173 -917
rect -137 -943 -111 -917
rect -75 -943 -49 -917
rect -13 -943 13 -917
rect 49 -943 75 -917
rect 111 -943 137 -917
rect 173 -943 199 -917
rect 235 -943 261 -917
rect 297 -943 323 -917
rect 359 -943 385 -917
rect -385 -1005 -359 -979
rect -323 -1005 -297 -979
rect -261 -1005 -235 -979
rect -199 -1005 -173 -979
rect -137 -1005 -111 -979
rect -75 -1005 -49 -979
rect -13 -1005 13 -979
rect 49 -1005 75 -979
rect 111 -1005 137 -979
rect 173 -1005 199 -979
rect 235 -1005 261 -979
rect 297 -1005 323 -979
rect 359 -1005 385 -979
rect -385 -1067 -359 -1041
rect -323 -1067 -297 -1041
rect -261 -1067 -235 -1041
rect -199 -1067 -173 -1041
rect -137 -1067 -111 -1041
rect -75 -1067 -49 -1041
rect -13 -1067 13 -1041
rect 49 -1067 75 -1041
rect 111 -1067 137 -1041
rect 173 -1067 199 -1041
rect 235 -1067 261 -1041
rect 297 -1067 323 -1041
rect 359 -1067 385 -1041
rect -385 -1129 -359 -1103
rect -323 -1129 -297 -1103
rect -261 -1129 -235 -1103
rect -199 -1129 -173 -1103
rect -137 -1129 -111 -1103
rect -75 -1129 -49 -1103
rect -13 -1129 13 -1103
rect 49 -1129 75 -1103
rect 111 -1129 137 -1103
rect 173 -1129 199 -1103
rect 235 -1129 261 -1103
rect 297 -1129 323 -1103
rect 359 -1129 385 -1103
rect -385 -1191 -359 -1165
rect -323 -1191 -297 -1165
rect -261 -1191 -235 -1165
rect -199 -1191 -173 -1165
rect -137 -1191 -111 -1165
rect -75 -1191 -49 -1165
rect -13 -1191 13 -1165
rect 49 -1191 75 -1165
rect 111 -1191 137 -1165
rect 173 -1191 199 -1165
rect 235 -1191 261 -1165
rect 297 -1191 323 -1165
rect 359 -1191 385 -1165
rect -385 -1253 -359 -1227
rect -323 -1253 -297 -1227
rect -261 -1253 -235 -1227
rect -199 -1253 -173 -1227
rect -137 -1253 -111 -1227
rect -75 -1253 -49 -1227
rect -13 -1253 13 -1227
rect 49 -1253 75 -1227
rect 111 -1253 137 -1227
rect 173 -1253 199 -1227
rect 235 -1253 261 -1227
rect 297 -1253 323 -1227
rect 359 -1253 385 -1227
rect -385 -1315 -359 -1289
rect -323 -1315 -297 -1289
rect -261 -1315 -235 -1289
rect -199 -1315 -173 -1289
rect -137 -1315 -111 -1289
rect -75 -1315 -49 -1289
rect -13 -1315 13 -1289
rect 49 -1315 75 -1289
rect 111 -1315 137 -1289
rect 173 -1315 199 -1289
rect 235 -1315 261 -1289
rect 297 -1315 323 -1289
rect 359 -1315 385 -1289
rect -385 -1377 -359 -1351
rect -323 -1377 -297 -1351
rect -261 -1377 -235 -1351
rect -199 -1377 -173 -1351
rect -137 -1377 -111 -1351
rect -75 -1377 -49 -1351
rect -13 -1377 13 -1351
rect 49 -1377 75 -1351
rect 111 -1377 137 -1351
rect 173 -1377 199 -1351
rect 235 -1377 261 -1351
rect 297 -1377 323 -1351
rect 359 -1377 385 -1351
rect -385 -1439 -359 -1413
rect -323 -1439 -297 -1413
rect -261 -1439 -235 -1413
rect -199 -1439 -173 -1413
rect -137 -1439 -111 -1413
rect -75 -1439 -49 -1413
rect -13 -1439 13 -1413
rect 49 -1439 75 -1413
rect 111 -1439 137 -1413
rect 173 -1439 199 -1413
rect 235 -1439 261 -1413
rect 297 -1439 323 -1413
rect 359 -1439 385 -1413
rect -385 -1501 -359 -1475
rect -323 -1501 -297 -1475
rect -261 -1501 -235 -1475
rect -199 -1501 -173 -1475
rect -137 -1501 -111 -1475
rect -75 -1501 -49 -1475
rect -13 -1501 13 -1475
rect 49 -1501 75 -1475
rect 111 -1501 137 -1475
rect 173 -1501 199 -1475
rect 235 -1501 261 -1475
rect 297 -1501 323 -1475
rect 359 -1501 385 -1475
rect -385 -1563 -359 -1537
rect -323 -1563 -297 -1537
rect -261 -1563 -235 -1537
rect -199 -1563 -173 -1537
rect -137 -1563 -111 -1537
rect -75 -1563 -49 -1537
rect -13 -1563 13 -1537
rect 49 -1563 75 -1537
rect 111 -1563 137 -1537
rect 173 -1563 199 -1537
rect 235 -1563 261 -1537
rect 297 -1563 323 -1537
rect 359 -1563 385 -1537
rect -385 -1625 -359 -1599
rect -323 -1625 -297 -1599
rect -261 -1625 -235 -1599
rect -199 -1625 -173 -1599
rect -137 -1625 -111 -1599
rect -75 -1625 -49 -1599
rect -13 -1625 13 -1599
rect 49 -1625 75 -1599
rect 111 -1625 137 -1599
rect 173 -1625 199 -1599
rect 235 -1625 261 -1599
rect 297 -1625 323 -1599
rect 359 -1625 385 -1599
rect -385 -1687 -359 -1661
rect -323 -1687 -297 -1661
rect -261 -1687 -235 -1661
rect -199 -1687 -173 -1661
rect -137 -1687 -111 -1661
rect -75 -1687 -49 -1661
rect -13 -1687 13 -1661
rect 49 -1687 75 -1661
rect 111 -1687 137 -1661
rect 173 -1687 199 -1661
rect 235 -1687 261 -1661
rect 297 -1687 323 -1661
rect 359 -1687 385 -1661
rect -385 -1749 -359 -1723
rect -323 -1749 -297 -1723
rect -261 -1749 -235 -1723
rect -199 -1749 -173 -1723
rect -137 -1749 -111 -1723
rect -75 -1749 -49 -1723
rect -13 -1749 13 -1723
rect 49 -1749 75 -1723
rect 111 -1749 137 -1723
rect 173 -1749 199 -1723
rect 235 -1749 261 -1723
rect 297 -1749 323 -1723
rect 359 -1749 385 -1723
rect -385 -1811 -359 -1785
rect -323 -1811 -297 -1785
rect -261 -1811 -235 -1785
rect -199 -1811 -173 -1785
rect -137 -1811 -111 -1785
rect -75 -1811 -49 -1785
rect -13 -1811 13 -1785
rect 49 -1811 75 -1785
rect 111 -1811 137 -1785
rect 173 -1811 199 -1785
rect 235 -1811 261 -1785
rect 297 -1811 323 -1785
rect 359 -1811 385 -1785
rect -385 -1873 -359 -1847
rect -323 -1873 -297 -1847
rect -261 -1873 -235 -1847
rect -199 -1873 -173 -1847
rect -137 -1873 -111 -1847
rect -75 -1873 -49 -1847
rect -13 -1873 13 -1847
rect 49 -1873 75 -1847
rect 111 -1873 137 -1847
rect 173 -1873 199 -1847
rect 235 -1873 261 -1847
rect 297 -1873 323 -1847
rect 359 -1873 385 -1847
<< metal2 >>
rect -391 1873 391 1879
rect -391 1847 -385 1873
rect -359 1847 -323 1873
rect -297 1847 -261 1873
rect -235 1847 -199 1873
rect -173 1847 -137 1873
rect -111 1847 -75 1873
rect -49 1847 -13 1873
rect 13 1847 49 1873
rect 75 1847 111 1873
rect 137 1847 173 1873
rect 199 1847 235 1873
rect 261 1847 297 1873
rect 323 1847 359 1873
rect 385 1847 391 1873
rect -391 1811 391 1847
rect -391 1785 -385 1811
rect -359 1785 -323 1811
rect -297 1785 -261 1811
rect -235 1785 -199 1811
rect -173 1785 -137 1811
rect -111 1785 -75 1811
rect -49 1785 -13 1811
rect 13 1785 49 1811
rect 75 1785 111 1811
rect 137 1785 173 1811
rect 199 1785 235 1811
rect 261 1785 297 1811
rect 323 1785 359 1811
rect 385 1785 391 1811
rect -391 1749 391 1785
rect -391 1723 -385 1749
rect -359 1723 -323 1749
rect -297 1723 -261 1749
rect -235 1723 -199 1749
rect -173 1723 -137 1749
rect -111 1723 -75 1749
rect -49 1723 -13 1749
rect 13 1723 49 1749
rect 75 1723 111 1749
rect 137 1723 173 1749
rect 199 1723 235 1749
rect 261 1723 297 1749
rect 323 1723 359 1749
rect 385 1723 391 1749
rect -391 1687 391 1723
rect -391 1661 -385 1687
rect -359 1661 -323 1687
rect -297 1661 -261 1687
rect -235 1661 -199 1687
rect -173 1661 -137 1687
rect -111 1661 -75 1687
rect -49 1661 -13 1687
rect 13 1661 49 1687
rect 75 1661 111 1687
rect 137 1661 173 1687
rect 199 1661 235 1687
rect 261 1661 297 1687
rect 323 1661 359 1687
rect 385 1661 391 1687
rect -391 1625 391 1661
rect -391 1599 -385 1625
rect -359 1599 -323 1625
rect -297 1599 -261 1625
rect -235 1599 -199 1625
rect -173 1599 -137 1625
rect -111 1599 -75 1625
rect -49 1599 -13 1625
rect 13 1599 49 1625
rect 75 1599 111 1625
rect 137 1599 173 1625
rect 199 1599 235 1625
rect 261 1599 297 1625
rect 323 1599 359 1625
rect 385 1599 391 1625
rect -391 1563 391 1599
rect -391 1537 -385 1563
rect -359 1537 -323 1563
rect -297 1537 -261 1563
rect -235 1537 -199 1563
rect -173 1537 -137 1563
rect -111 1537 -75 1563
rect -49 1537 -13 1563
rect 13 1537 49 1563
rect 75 1537 111 1563
rect 137 1537 173 1563
rect 199 1537 235 1563
rect 261 1537 297 1563
rect 323 1537 359 1563
rect 385 1537 391 1563
rect -391 1501 391 1537
rect -391 1475 -385 1501
rect -359 1475 -323 1501
rect -297 1475 -261 1501
rect -235 1475 -199 1501
rect -173 1475 -137 1501
rect -111 1475 -75 1501
rect -49 1475 -13 1501
rect 13 1475 49 1501
rect 75 1475 111 1501
rect 137 1475 173 1501
rect 199 1475 235 1501
rect 261 1475 297 1501
rect 323 1475 359 1501
rect 385 1475 391 1501
rect -391 1439 391 1475
rect -391 1413 -385 1439
rect -359 1413 -323 1439
rect -297 1413 -261 1439
rect -235 1413 -199 1439
rect -173 1413 -137 1439
rect -111 1413 -75 1439
rect -49 1413 -13 1439
rect 13 1413 49 1439
rect 75 1413 111 1439
rect 137 1413 173 1439
rect 199 1413 235 1439
rect 261 1413 297 1439
rect 323 1413 359 1439
rect 385 1413 391 1439
rect -391 1377 391 1413
rect -391 1351 -385 1377
rect -359 1351 -323 1377
rect -297 1351 -261 1377
rect -235 1351 -199 1377
rect -173 1351 -137 1377
rect -111 1351 -75 1377
rect -49 1351 -13 1377
rect 13 1351 49 1377
rect 75 1351 111 1377
rect 137 1351 173 1377
rect 199 1351 235 1377
rect 261 1351 297 1377
rect 323 1351 359 1377
rect 385 1351 391 1377
rect -391 1315 391 1351
rect -391 1289 -385 1315
rect -359 1289 -323 1315
rect -297 1289 -261 1315
rect -235 1289 -199 1315
rect -173 1289 -137 1315
rect -111 1289 -75 1315
rect -49 1289 -13 1315
rect 13 1289 49 1315
rect 75 1289 111 1315
rect 137 1289 173 1315
rect 199 1289 235 1315
rect 261 1289 297 1315
rect 323 1289 359 1315
rect 385 1289 391 1315
rect -391 1253 391 1289
rect -391 1227 -385 1253
rect -359 1227 -323 1253
rect -297 1227 -261 1253
rect -235 1227 -199 1253
rect -173 1227 -137 1253
rect -111 1227 -75 1253
rect -49 1227 -13 1253
rect 13 1227 49 1253
rect 75 1227 111 1253
rect 137 1227 173 1253
rect 199 1227 235 1253
rect 261 1227 297 1253
rect 323 1227 359 1253
rect 385 1227 391 1253
rect -391 1191 391 1227
rect -391 1165 -385 1191
rect -359 1165 -323 1191
rect -297 1165 -261 1191
rect -235 1165 -199 1191
rect -173 1165 -137 1191
rect -111 1165 -75 1191
rect -49 1165 -13 1191
rect 13 1165 49 1191
rect 75 1165 111 1191
rect 137 1165 173 1191
rect 199 1165 235 1191
rect 261 1165 297 1191
rect 323 1165 359 1191
rect 385 1165 391 1191
rect -391 1129 391 1165
rect -391 1103 -385 1129
rect -359 1103 -323 1129
rect -297 1103 -261 1129
rect -235 1103 -199 1129
rect -173 1103 -137 1129
rect -111 1103 -75 1129
rect -49 1103 -13 1129
rect 13 1103 49 1129
rect 75 1103 111 1129
rect 137 1103 173 1129
rect 199 1103 235 1129
rect 261 1103 297 1129
rect 323 1103 359 1129
rect 385 1103 391 1129
rect -391 1067 391 1103
rect -391 1041 -385 1067
rect -359 1041 -323 1067
rect -297 1041 -261 1067
rect -235 1041 -199 1067
rect -173 1041 -137 1067
rect -111 1041 -75 1067
rect -49 1041 -13 1067
rect 13 1041 49 1067
rect 75 1041 111 1067
rect 137 1041 173 1067
rect 199 1041 235 1067
rect 261 1041 297 1067
rect 323 1041 359 1067
rect 385 1041 391 1067
rect -391 1005 391 1041
rect -391 979 -385 1005
rect -359 979 -323 1005
rect -297 979 -261 1005
rect -235 979 -199 1005
rect -173 979 -137 1005
rect -111 979 -75 1005
rect -49 979 -13 1005
rect 13 979 49 1005
rect 75 979 111 1005
rect 137 979 173 1005
rect 199 979 235 1005
rect 261 979 297 1005
rect 323 979 359 1005
rect 385 979 391 1005
rect -391 943 391 979
rect -391 917 -385 943
rect -359 917 -323 943
rect -297 917 -261 943
rect -235 917 -199 943
rect -173 917 -137 943
rect -111 917 -75 943
rect -49 917 -13 943
rect 13 917 49 943
rect 75 917 111 943
rect 137 917 173 943
rect 199 917 235 943
rect 261 917 297 943
rect 323 917 359 943
rect 385 917 391 943
rect -391 881 391 917
rect -391 855 -385 881
rect -359 855 -323 881
rect -297 855 -261 881
rect -235 855 -199 881
rect -173 855 -137 881
rect -111 855 -75 881
rect -49 855 -13 881
rect 13 855 49 881
rect 75 855 111 881
rect 137 855 173 881
rect 199 855 235 881
rect 261 855 297 881
rect 323 855 359 881
rect 385 855 391 881
rect -391 819 391 855
rect -391 793 -385 819
rect -359 793 -323 819
rect -297 793 -261 819
rect -235 793 -199 819
rect -173 793 -137 819
rect -111 793 -75 819
rect -49 793 -13 819
rect 13 793 49 819
rect 75 793 111 819
rect 137 793 173 819
rect 199 793 235 819
rect 261 793 297 819
rect 323 793 359 819
rect 385 793 391 819
rect -391 757 391 793
rect -391 731 -385 757
rect -359 731 -323 757
rect -297 731 -261 757
rect -235 731 -199 757
rect -173 731 -137 757
rect -111 731 -75 757
rect -49 731 -13 757
rect 13 731 49 757
rect 75 731 111 757
rect 137 731 173 757
rect 199 731 235 757
rect 261 731 297 757
rect 323 731 359 757
rect 385 731 391 757
rect -391 695 391 731
rect -391 669 -385 695
rect -359 669 -323 695
rect -297 669 -261 695
rect -235 669 -199 695
rect -173 669 -137 695
rect -111 669 -75 695
rect -49 669 -13 695
rect 13 669 49 695
rect 75 669 111 695
rect 137 669 173 695
rect 199 669 235 695
rect 261 669 297 695
rect 323 669 359 695
rect 385 669 391 695
rect -391 633 391 669
rect -391 607 -385 633
rect -359 607 -323 633
rect -297 607 -261 633
rect -235 607 -199 633
rect -173 607 -137 633
rect -111 607 -75 633
rect -49 607 -13 633
rect 13 607 49 633
rect 75 607 111 633
rect 137 607 173 633
rect 199 607 235 633
rect 261 607 297 633
rect 323 607 359 633
rect 385 607 391 633
rect -391 571 391 607
rect -391 545 -385 571
rect -359 545 -323 571
rect -297 545 -261 571
rect -235 545 -199 571
rect -173 545 -137 571
rect -111 545 -75 571
rect -49 545 -13 571
rect 13 545 49 571
rect 75 545 111 571
rect 137 545 173 571
rect 199 545 235 571
rect 261 545 297 571
rect 323 545 359 571
rect 385 545 391 571
rect -391 509 391 545
rect -391 483 -385 509
rect -359 483 -323 509
rect -297 483 -261 509
rect -235 483 -199 509
rect -173 483 -137 509
rect -111 483 -75 509
rect -49 483 -13 509
rect 13 483 49 509
rect 75 483 111 509
rect 137 483 173 509
rect 199 483 235 509
rect 261 483 297 509
rect 323 483 359 509
rect 385 483 391 509
rect -391 447 391 483
rect -391 421 -385 447
rect -359 421 -323 447
rect -297 421 -261 447
rect -235 421 -199 447
rect -173 421 -137 447
rect -111 421 -75 447
rect -49 421 -13 447
rect 13 421 49 447
rect 75 421 111 447
rect 137 421 173 447
rect 199 421 235 447
rect 261 421 297 447
rect 323 421 359 447
rect 385 421 391 447
rect -391 385 391 421
rect -391 359 -385 385
rect -359 359 -323 385
rect -297 359 -261 385
rect -235 359 -199 385
rect -173 359 -137 385
rect -111 359 -75 385
rect -49 359 -13 385
rect 13 359 49 385
rect 75 359 111 385
rect 137 359 173 385
rect 199 359 235 385
rect 261 359 297 385
rect 323 359 359 385
rect 385 359 391 385
rect -391 323 391 359
rect -391 297 -385 323
rect -359 297 -323 323
rect -297 297 -261 323
rect -235 297 -199 323
rect -173 297 -137 323
rect -111 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 111 323
rect 137 297 173 323
rect 199 297 235 323
rect 261 297 297 323
rect 323 297 359 323
rect 385 297 391 323
rect -391 261 391 297
rect -391 235 -385 261
rect -359 235 -323 261
rect -297 235 -261 261
rect -235 235 -199 261
rect -173 235 -137 261
rect -111 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 111 261
rect 137 235 173 261
rect 199 235 235 261
rect 261 235 297 261
rect 323 235 359 261
rect 385 235 391 261
rect -391 199 391 235
rect -391 173 -385 199
rect -359 173 -323 199
rect -297 173 -261 199
rect -235 173 -199 199
rect -173 173 -137 199
rect -111 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 111 199
rect 137 173 173 199
rect 199 173 235 199
rect 261 173 297 199
rect 323 173 359 199
rect 385 173 391 199
rect -391 137 391 173
rect -391 111 -385 137
rect -359 111 -323 137
rect -297 111 -261 137
rect -235 111 -199 137
rect -173 111 -137 137
rect -111 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 111 137
rect 137 111 173 137
rect 199 111 235 137
rect 261 111 297 137
rect 323 111 359 137
rect 385 111 391 137
rect -391 75 391 111
rect -391 49 -385 75
rect -359 49 -323 75
rect -297 49 -261 75
rect -235 49 -199 75
rect -173 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 173 75
rect 199 49 235 75
rect 261 49 297 75
rect 323 49 359 75
rect 385 49 391 75
rect -391 13 391 49
rect -391 -13 -385 13
rect -359 -13 -323 13
rect -297 -13 -261 13
rect -235 -13 -199 13
rect -173 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 173 13
rect 199 -13 235 13
rect 261 -13 297 13
rect 323 -13 359 13
rect 385 -13 391 13
rect -391 -49 391 -13
rect -391 -75 -385 -49
rect -359 -75 -323 -49
rect -297 -75 -261 -49
rect -235 -75 -199 -49
rect -173 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 173 -49
rect 199 -75 235 -49
rect 261 -75 297 -49
rect 323 -75 359 -49
rect 385 -75 391 -49
rect -391 -111 391 -75
rect -391 -137 -385 -111
rect -359 -137 -323 -111
rect -297 -137 -261 -111
rect -235 -137 -199 -111
rect -173 -137 -137 -111
rect -111 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 111 -111
rect 137 -137 173 -111
rect 199 -137 235 -111
rect 261 -137 297 -111
rect 323 -137 359 -111
rect 385 -137 391 -111
rect -391 -173 391 -137
rect -391 -199 -385 -173
rect -359 -199 -323 -173
rect -297 -199 -261 -173
rect -235 -199 -199 -173
rect -173 -199 -137 -173
rect -111 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 111 -173
rect 137 -199 173 -173
rect 199 -199 235 -173
rect 261 -199 297 -173
rect 323 -199 359 -173
rect 385 -199 391 -173
rect -391 -235 391 -199
rect -391 -261 -385 -235
rect -359 -261 -323 -235
rect -297 -261 -261 -235
rect -235 -261 -199 -235
rect -173 -261 -137 -235
rect -111 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 111 -235
rect 137 -261 173 -235
rect 199 -261 235 -235
rect 261 -261 297 -235
rect 323 -261 359 -235
rect 385 -261 391 -235
rect -391 -297 391 -261
rect -391 -323 -385 -297
rect -359 -323 -323 -297
rect -297 -323 -261 -297
rect -235 -323 -199 -297
rect -173 -323 -137 -297
rect -111 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 111 -297
rect 137 -323 173 -297
rect 199 -323 235 -297
rect 261 -323 297 -297
rect 323 -323 359 -297
rect 385 -323 391 -297
rect -391 -359 391 -323
rect -391 -385 -385 -359
rect -359 -385 -323 -359
rect -297 -385 -261 -359
rect -235 -385 -199 -359
rect -173 -385 -137 -359
rect -111 -385 -75 -359
rect -49 -385 -13 -359
rect 13 -385 49 -359
rect 75 -385 111 -359
rect 137 -385 173 -359
rect 199 -385 235 -359
rect 261 -385 297 -359
rect 323 -385 359 -359
rect 385 -385 391 -359
rect -391 -421 391 -385
rect -391 -447 -385 -421
rect -359 -447 -323 -421
rect -297 -447 -261 -421
rect -235 -447 -199 -421
rect -173 -447 -137 -421
rect -111 -447 -75 -421
rect -49 -447 -13 -421
rect 13 -447 49 -421
rect 75 -447 111 -421
rect 137 -447 173 -421
rect 199 -447 235 -421
rect 261 -447 297 -421
rect 323 -447 359 -421
rect 385 -447 391 -421
rect -391 -483 391 -447
rect -391 -509 -385 -483
rect -359 -509 -323 -483
rect -297 -509 -261 -483
rect -235 -509 -199 -483
rect -173 -509 -137 -483
rect -111 -509 -75 -483
rect -49 -509 -13 -483
rect 13 -509 49 -483
rect 75 -509 111 -483
rect 137 -509 173 -483
rect 199 -509 235 -483
rect 261 -509 297 -483
rect 323 -509 359 -483
rect 385 -509 391 -483
rect -391 -545 391 -509
rect -391 -571 -385 -545
rect -359 -571 -323 -545
rect -297 -571 -261 -545
rect -235 -571 -199 -545
rect -173 -571 -137 -545
rect -111 -571 -75 -545
rect -49 -571 -13 -545
rect 13 -571 49 -545
rect 75 -571 111 -545
rect 137 -571 173 -545
rect 199 -571 235 -545
rect 261 -571 297 -545
rect 323 -571 359 -545
rect 385 -571 391 -545
rect -391 -607 391 -571
rect -391 -633 -385 -607
rect -359 -633 -323 -607
rect -297 -633 -261 -607
rect -235 -633 -199 -607
rect -173 -633 -137 -607
rect -111 -633 -75 -607
rect -49 -633 -13 -607
rect 13 -633 49 -607
rect 75 -633 111 -607
rect 137 -633 173 -607
rect 199 -633 235 -607
rect 261 -633 297 -607
rect 323 -633 359 -607
rect 385 -633 391 -607
rect -391 -669 391 -633
rect -391 -695 -385 -669
rect -359 -695 -323 -669
rect -297 -695 -261 -669
rect -235 -695 -199 -669
rect -173 -695 -137 -669
rect -111 -695 -75 -669
rect -49 -695 -13 -669
rect 13 -695 49 -669
rect 75 -695 111 -669
rect 137 -695 173 -669
rect 199 -695 235 -669
rect 261 -695 297 -669
rect 323 -695 359 -669
rect 385 -695 391 -669
rect -391 -731 391 -695
rect -391 -757 -385 -731
rect -359 -757 -323 -731
rect -297 -757 -261 -731
rect -235 -757 -199 -731
rect -173 -757 -137 -731
rect -111 -757 -75 -731
rect -49 -757 -13 -731
rect 13 -757 49 -731
rect 75 -757 111 -731
rect 137 -757 173 -731
rect 199 -757 235 -731
rect 261 -757 297 -731
rect 323 -757 359 -731
rect 385 -757 391 -731
rect -391 -793 391 -757
rect -391 -819 -385 -793
rect -359 -819 -323 -793
rect -297 -819 -261 -793
rect -235 -819 -199 -793
rect -173 -819 -137 -793
rect -111 -819 -75 -793
rect -49 -819 -13 -793
rect 13 -819 49 -793
rect 75 -819 111 -793
rect 137 -819 173 -793
rect 199 -819 235 -793
rect 261 -819 297 -793
rect 323 -819 359 -793
rect 385 -819 391 -793
rect -391 -855 391 -819
rect -391 -881 -385 -855
rect -359 -881 -323 -855
rect -297 -881 -261 -855
rect -235 -881 -199 -855
rect -173 -881 -137 -855
rect -111 -881 -75 -855
rect -49 -881 -13 -855
rect 13 -881 49 -855
rect 75 -881 111 -855
rect 137 -881 173 -855
rect 199 -881 235 -855
rect 261 -881 297 -855
rect 323 -881 359 -855
rect 385 -881 391 -855
rect -391 -917 391 -881
rect -391 -943 -385 -917
rect -359 -943 -323 -917
rect -297 -943 -261 -917
rect -235 -943 -199 -917
rect -173 -943 -137 -917
rect -111 -943 -75 -917
rect -49 -943 -13 -917
rect 13 -943 49 -917
rect 75 -943 111 -917
rect 137 -943 173 -917
rect 199 -943 235 -917
rect 261 -943 297 -917
rect 323 -943 359 -917
rect 385 -943 391 -917
rect -391 -979 391 -943
rect -391 -1005 -385 -979
rect -359 -1005 -323 -979
rect -297 -1005 -261 -979
rect -235 -1005 -199 -979
rect -173 -1005 -137 -979
rect -111 -1005 -75 -979
rect -49 -1005 -13 -979
rect 13 -1005 49 -979
rect 75 -1005 111 -979
rect 137 -1005 173 -979
rect 199 -1005 235 -979
rect 261 -1005 297 -979
rect 323 -1005 359 -979
rect 385 -1005 391 -979
rect -391 -1041 391 -1005
rect -391 -1067 -385 -1041
rect -359 -1067 -323 -1041
rect -297 -1067 -261 -1041
rect -235 -1067 -199 -1041
rect -173 -1067 -137 -1041
rect -111 -1067 -75 -1041
rect -49 -1067 -13 -1041
rect 13 -1067 49 -1041
rect 75 -1067 111 -1041
rect 137 -1067 173 -1041
rect 199 -1067 235 -1041
rect 261 -1067 297 -1041
rect 323 -1067 359 -1041
rect 385 -1067 391 -1041
rect -391 -1103 391 -1067
rect -391 -1129 -385 -1103
rect -359 -1129 -323 -1103
rect -297 -1129 -261 -1103
rect -235 -1129 -199 -1103
rect -173 -1129 -137 -1103
rect -111 -1129 -75 -1103
rect -49 -1129 -13 -1103
rect 13 -1129 49 -1103
rect 75 -1129 111 -1103
rect 137 -1129 173 -1103
rect 199 -1129 235 -1103
rect 261 -1129 297 -1103
rect 323 -1129 359 -1103
rect 385 -1129 391 -1103
rect -391 -1165 391 -1129
rect -391 -1191 -385 -1165
rect -359 -1191 -323 -1165
rect -297 -1191 -261 -1165
rect -235 -1191 -199 -1165
rect -173 -1191 -137 -1165
rect -111 -1191 -75 -1165
rect -49 -1191 -13 -1165
rect 13 -1191 49 -1165
rect 75 -1191 111 -1165
rect 137 -1191 173 -1165
rect 199 -1191 235 -1165
rect 261 -1191 297 -1165
rect 323 -1191 359 -1165
rect 385 -1191 391 -1165
rect -391 -1227 391 -1191
rect -391 -1253 -385 -1227
rect -359 -1253 -323 -1227
rect -297 -1253 -261 -1227
rect -235 -1253 -199 -1227
rect -173 -1253 -137 -1227
rect -111 -1253 -75 -1227
rect -49 -1253 -13 -1227
rect 13 -1253 49 -1227
rect 75 -1253 111 -1227
rect 137 -1253 173 -1227
rect 199 -1253 235 -1227
rect 261 -1253 297 -1227
rect 323 -1253 359 -1227
rect 385 -1253 391 -1227
rect -391 -1289 391 -1253
rect -391 -1315 -385 -1289
rect -359 -1315 -323 -1289
rect -297 -1315 -261 -1289
rect -235 -1315 -199 -1289
rect -173 -1315 -137 -1289
rect -111 -1315 -75 -1289
rect -49 -1315 -13 -1289
rect 13 -1315 49 -1289
rect 75 -1315 111 -1289
rect 137 -1315 173 -1289
rect 199 -1315 235 -1289
rect 261 -1315 297 -1289
rect 323 -1315 359 -1289
rect 385 -1315 391 -1289
rect -391 -1351 391 -1315
rect -391 -1377 -385 -1351
rect -359 -1377 -323 -1351
rect -297 -1377 -261 -1351
rect -235 -1377 -199 -1351
rect -173 -1377 -137 -1351
rect -111 -1377 -75 -1351
rect -49 -1377 -13 -1351
rect 13 -1377 49 -1351
rect 75 -1377 111 -1351
rect 137 -1377 173 -1351
rect 199 -1377 235 -1351
rect 261 -1377 297 -1351
rect 323 -1377 359 -1351
rect 385 -1377 391 -1351
rect -391 -1413 391 -1377
rect -391 -1439 -385 -1413
rect -359 -1439 -323 -1413
rect -297 -1439 -261 -1413
rect -235 -1439 -199 -1413
rect -173 -1439 -137 -1413
rect -111 -1439 -75 -1413
rect -49 -1439 -13 -1413
rect 13 -1439 49 -1413
rect 75 -1439 111 -1413
rect 137 -1439 173 -1413
rect 199 -1439 235 -1413
rect 261 -1439 297 -1413
rect 323 -1439 359 -1413
rect 385 -1439 391 -1413
rect -391 -1475 391 -1439
rect -391 -1501 -385 -1475
rect -359 -1501 -323 -1475
rect -297 -1501 -261 -1475
rect -235 -1501 -199 -1475
rect -173 -1501 -137 -1475
rect -111 -1501 -75 -1475
rect -49 -1501 -13 -1475
rect 13 -1501 49 -1475
rect 75 -1501 111 -1475
rect 137 -1501 173 -1475
rect 199 -1501 235 -1475
rect 261 -1501 297 -1475
rect 323 -1501 359 -1475
rect 385 -1501 391 -1475
rect -391 -1537 391 -1501
rect -391 -1563 -385 -1537
rect -359 -1563 -323 -1537
rect -297 -1563 -261 -1537
rect -235 -1563 -199 -1537
rect -173 -1563 -137 -1537
rect -111 -1563 -75 -1537
rect -49 -1563 -13 -1537
rect 13 -1563 49 -1537
rect 75 -1563 111 -1537
rect 137 -1563 173 -1537
rect 199 -1563 235 -1537
rect 261 -1563 297 -1537
rect 323 -1563 359 -1537
rect 385 -1563 391 -1537
rect -391 -1599 391 -1563
rect -391 -1625 -385 -1599
rect -359 -1625 -323 -1599
rect -297 -1625 -261 -1599
rect -235 -1625 -199 -1599
rect -173 -1625 -137 -1599
rect -111 -1625 -75 -1599
rect -49 -1625 -13 -1599
rect 13 -1625 49 -1599
rect 75 -1625 111 -1599
rect 137 -1625 173 -1599
rect 199 -1625 235 -1599
rect 261 -1625 297 -1599
rect 323 -1625 359 -1599
rect 385 -1625 391 -1599
rect -391 -1661 391 -1625
rect -391 -1687 -385 -1661
rect -359 -1687 -323 -1661
rect -297 -1687 -261 -1661
rect -235 -1687 -199 -1661
rect -173 -1687 -137 -1661
rect -111 -1687 -75 -1661
rect -49 -1687 -13 -1661
rect 13 -1687 49 -1661
rect 75 -1687 111 -1661
rect 137 -1687 173 -1661
rect 199 -1687 235 -1661
rect 261 -1687 297 -1661
rect 323 -1687 359 -1661
rect 385 -1687 391 -1661
rect -391 -1723 391 -1687
rect -391 -1749 -385 -1723
rect -359 -1749 -323 -1723
rect -297 -1749 -261 -1723
rect -235 -1749 -199 -1723
rect -173 -1749 -137 -1723
rect -111 -1749 -75 -1723
rect -49 -1749 -13 -1723
rect 13 -1749 49 -1723
rect 75 -1749 111 -1723
rect 137 -1749 173 -1723
rect 199 -1749 235 -1723
rect 261 -1749 297 -1723
rect 323 -1749 359 -1723
rect 385 -1749 391 -1723
rect -391 -1785 391 -1749
rect -391 -1811 -385 -1785
rect -359 -1811 -323 -1785
rect -297 -1811 -261 -1785
rect -235 -1811 -199 -1785
rect -173 -1811 -137 -1785
rect -111 -1811 -75 -1785
rect -49 -1811 -13 -1785
rect 13 -1811 49 -1785
rect 75 -1811 111 -1785
rect 137 -1811 173 -1785
rect 199 -1811 235 -1785
rect 261 -1811 297 -1785
rect 323 -1811 359 -1785
rect 385 -1811 391 -1785
rect -391 -1847 391 -1811
rect -391 -1873 -385 -1847
rect -359 -1873 -323 -1847
rect -297 -1873 -261 -1847
rect -235 -1873 -199 -1847
rect -173 -1873 -137 -1847
rect -111 -1873 -75 -1847
rect -49 -1873 -13 -1847
rect 13 -1873 49 -1847
rect 75 -1873 111 -1847
rect 137 -1873 173 -1847
rect 199 -1873 235 -1847
rect 261 -1873 297 -1847
rect 323 -1873 359 -1847
rect 385 -1873 391 -1847
rect -391 -1879 391 -1873
<< end >>
