magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6416 -2045 6416 2045
<< psubdiff >>
rect -4416 23 4416 45
rect -4416 -23 -4394 23
rect 4394 -23 4416 23
rect -4416 -45 4416 -23
<< psubdiffcont >>
rect -4394 -23 4394 23
<< metal1 >>
rect -4405 23 4405 34
rect -4405 -23 -4394 23
rect 4394 -23 4405 23
rect -4405 -34 4405 -23
<< end >>
