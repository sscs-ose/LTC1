magic
tech gf180mcuD
magscale 1 10
timestamp 1713358893
<< checkpaint >>
rect 1672 -3154 11606 6970
<< polysilicon >>
rect 8586 3098 8806 3202
rect 4386 2270 4606 2374
rect 8586 1442 8806 1546
rect 4386 614 4606 718
<< metal1 >>
rect 4010 4887 9182 4933
rect 4427 4741 4574 4887
rect 4088 4695 9104 4741
rect 4184 4089 4233 4695
rect 8990 4089 9039 4695
rect 4088 4043 9104 4089
rect 3766 3930 3845 3944
rect 3766 3926 3782 3930
rect 3672 3878 3782 3926
rect 3834 3878 3845 3930
rect 3672 3873 3845 3878
rect 3766 3865 3845 3873
rect 4184 -227 4233 4043
rect 4475 3930 4565 3944
rect 4475 3878 4490 3930
rect 4542 3878 4565 3930
rect 4475 3851 4565 3878
rect 4688 3867 5204 3913
rect 5288 3867 5804 3913
rect 5888 3867 6404 3913
rect 6488 3867 7004 3913
rect 7088 3867 7604 3913
rect 7688 3867 8204 3913
rect 8288 3867 8804 3913
rect 4388 3215 4904 3261
rect 4988 3215 5504 3261
rect 5588 3215 6104 3261
rect 6188 3215 6704 3261
rect 6788 3215 7304 3261
rect 7388 3215 7904 3261
rect 7988 3215 8504 3261
rect 4388 3039 4904 3085
rect 4988 3039 5504 3085
rect 5588 3039 6104 3085
rect 6188 3039 6704 3085
rect 6788 3039 7304 3085
rect 7388 3039 7904 3085
rect 7988 3039 8504 3085
rect 4688 2387 5204 2433
rect 5288 2387 5804 2433
rect 5888 2387 6404 2433
rect 6488 2387 7004 2433
rect 7088 2387 7604 2433
rect 7688 2387 8204 2433
rect 8288 2387 8804 2433
rect 4688 2211 5204 2257
rect 5288 2211 5804 2257
rect 5888 2211 6404 2257
rect 6488 2211 7004 2257
rect 7088 2211 7604 2257
rect 7688 2211 8204 2257
rect 8288 2211 8804 2257
rect 4388 1559 4904 1605
rect 4988 1559 5504 1605
rect 5588 1559 6104 1605
rect 6188 1559 6704 1605
rect 6788 1559 7304 1605
rect 7388 1559 7904 1605
rect 7988 1559 8504 1605
rect 4388 1383 4904 1429
rect 4988 1383 5504 1429
rect 5588 1383 6104 1429
rect 6188 1383 6704 1429
rect 6788 1383 7304 1429
rect 7388 1383 7904 1429
rect 7988 1383 8504 1429
rect 4688 731 5204 777
rect 5288 731 5804 777
rect 5888 731 6404 777
rect 6488 731 7004 777
rect 7088 731 7604 777
rect 7688 731 8204 777
rect 8288 731 8804 777
rect 4688 555 5204 601
rect 5288 555 5804 601
rect 5888 555 6404 601
rect 6488 555 7004 601
rect 7088 555 7604 601
rect 7688 555 8204 601
rect 8288 555 8804 601
rect 4388 -97 4904 -51
rect 4988 -97 5504 -51
rect 5588 -97 6104 -51
rect 6188 -97 6704 -51
rect 6788 -97 7304 -51
rect 7388 -97 7904 -51
rect 7988 -97 8504 -51
rect 8645 -52 8753 -33
rect 8645 -104 8663 -52
rect 8715 -104 8753 -52
rect 8645 -120 8753 -104
rect 8990 -227 9039 4043
rect 9417 -50 9499 -31
rect 9417 -102 9432 -50
rect 9484 -102 9606 -50
rect 9417 -104 9606 -102
rect 9417 -120 9499 -104
rect 4088 -273 9104 -227
rect 4184 -879 4233 -273
rect 8990 -879 9039 -273
rect 4088 -925 9104 -879
<< via1 >>
rect 3782 3878 3834 3930
rect 4490 3878 4542 3930
rect 8663 -104 8715 -52
rect 9432 -102 9484 -50
<< metal2 >>
rect 3766 3930 4610 3944
rect 3766 3878 3782 3930
rect 3834 3878 4490 3930
rect 4542 3878 4610 3930
rect 3766 3865 4610 3878
rect 8571 -31 9482 -30
rect 8571 -50 9499 -31
rect 8571 -52 9432 -50
rect 8571 -104 8663 -52
rect 8715 -102 9432 -52
rect 9484 -102 9499 -50
rect 8715 -104 9499 -102
rect 8571 -120 9499 -104
rect 8571 -121 9482 -120
use ppolyf_u_DTYK2C  ppolyf_u_DTYK2C_0
timestamp 1713274346
transform 1 0 6596 0 1 1908
box -2726 -3062 2726 3062
<< labels >>
flabel metal1 s 3714 3911 3714 3911 0 FreeSans 2500 0 0 0 M
port 1 nsew
flabel metal1 s 9563 -72 9563 -72 0 FreeSans 2500 0 0 0 P
port 2 nsew
flabel metal1 s 6495 4911 6495 4911 0 FreeSans 2500 0 0 0 VDD
port 3 nsew
<< end >>
