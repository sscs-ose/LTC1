magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1112 -1112 1112 1112
<< metal1 >>
rect -112 106 112 112
rect -112 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 112 106
rect -112 44 112 80
rect -112 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 112 44
rect -112 -18 112 18
rect -112 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 112 -18
rect -112 -80 112 -44
rect -112 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 112 -80
rect -112 -112 112 -106
<< via1 >>
rect -106 80 -80 106
rect -44 80 -18 106
rect 18 80 44 106
rect 80 80 106 106
rect -106 18 -80 44
rect -44 18 -18 44
rect 18 18 44 44
rect 80 18 106 44
rect -106 -44 -80 -18
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect 80 -44 106 -18
rect -106 -106 -80 -80
rect -44 -106 -18 -80
rect 18 -106 44 -80
rect 80 -106 106 -80
<< metal2 >>
rect -112 106 112 112
rect -112 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 112 106
rect -112 44 112 80
rect -112 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 112 44
rect -112 -18 112 18
rect -112 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 112 -18
rect -112 -80 112 -44
rect -112 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 112 -80
rect -112 -112 112 -106
<< end >>
