magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2195 -14045 2195 14045
<< psubdiff >>
rect -195 12023 195 12045
rect -195 -12023 -173 12023
rect 173 -12023 195 12023
rect -195 -12045 195 -12023
<< psubdiffcont >>
rect -173 -12023 173 12023
<< metal1 >>
rect -184 12023 184 12034
rect -184 -12023 -173 12023
rect 173 -12023 184 12023
rect -184 -12034 184 -12023
<< end >>
