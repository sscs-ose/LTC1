magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -2833 2128 2833
<< nwell >>
rect -128 -833 128 833
<< nsubdiff >>
rect -45 728 45 750
rect -45 -728 -23 728
rect 23 -728 45 728
rect -45 -750 45 -728
<< nsubdiffcont >>
rect -23 -728 23 728
<< metal1 >>
rect -34 728 34 739
rect -34 -728 -23 728
rect 23 -728 34 728
rect -34 -739 34 -728
<< end >>
