magic
tech gf180mcuC
magscale 1 10
timestamp 1699956126
<< pwell >>
rect -1182 -368 1182 368
<< nmos >>
rect -1070 -300 -970 300
rect -866 -300 -766 300
rect -662 -300 -562 300
rect -458 -300 -358 300
rect -254 -300 -154 300
rect -50 -300 50 300
rect 154 -300 254 300
rect 358 -300 458 300
rect 562 -300 662 300
rect 766 -300 866 300
rect 970 -300 1070 300
<< ndiff >>
rect -1158 287 -1070 300
rect -1158 -287 -1145 287
rect -1099 -287 -1070 287
rect -1158 -300 -1070 -287
rect -970 287 -866 300
rect -970 -287 -941 287
rect -895 -287 -866 287
rect -970 -300 -866 -287
rect -766 287 -662 300
rect -766 -287 -737 287
rect -691 -287 -662 287
rect -766 -300 -662 -287
rect -562 287 -458 300
rect -562 -287 -533 287
rect -487 -287 -458 287
rect -562 -300 -458 -287
rect -358 287 -254 300
rect -358 -287 -329 287
rect -283 -287 -254 287
rect -358 -300 -254 -287
rect -154 287 -50 300
rect -154 -287 -125 287
rect -79 -287 -50 287
rect -154 -300 -50 -287
rect 50 287 154 300
rect 50 -287 79 287
rect 125 -287 154 287
rect 50 -300 154 -287
rect 254 287 358 300
rect 254 -287 283 287
rect 329 -287 358 287
rect 254 -300 358 -287
rect 458 287 562 300
rect 458 -287 487 287
rect 533 -287 562 287
rect 458 -300 562 -287
rect 662 287 766 300
rect 662 -287 691 287
rect 737 -287 766 287
rect 662 -300 766 -287
rect 866 287 970 300
rect 866 -287 895 287
rect 941 -287 970 287
rect 866 -300 970 -287
rect 1070 287 1158 300
rect 1070 -287 1099 287
rect 1145 -287 1158 287
rect 1070 -300 1158 -287
<< ndiffc >>
rect -1145 -287 -1099 287
rect -941 -287 -895 287
rect -737 -287 -691 287
rect -533 -287 -487 287
rect -329 -287 -283 287
rect -125 -287 -79 287
rect 79 -287 125 287
rect 283 -287 329 287
rect 487 -287 533 287
rect 691 -287 737 287
rect 895 -287 941 287
rect 1099 -287 1145 287
<< polysilicon >>
rect -1070 300 -970 344
rect -866 300 -766 344
rect -662 300 -562 344
rect -458 300 -358 344
rect -254 300 -154 344
rect -50 300 50 344
rect 154 300 254 344
rect 358 300 458 344
rect 562 300 662 344
rect 766 300 866 344
rect 970 300 1070 344
rect -1070 -344 -970 -300
rect -866 -344 -766 -300
rect -662 -344 -562 -300
rect -458 -344 -358 -300
rect -254 -344 -154 -300
rect -50 -344 50 -300
rect 154 -344 254 -300
rect 358 -344 458 -300
rect 562 -344 662 -300
rect 766 -344 866 -300
rect 970 -344 1070 -300
<< metal1 >>
rect -1145 287 -1099 298
rect -1145 -298 -1099 -287
rect -941 287 -895 298
rect -941 -298 -895 -287
rect -737 287 -691 298
rect -737 -298 -691 -287
rect -533 287 -487 298
rect -533 -298 -487 -287
rect -329 287 -283 298
rect -329 -298 -283 -287
rect -125 287 -79 298
rect -125 -298 -79 -287
rect 79 287 125 298
rect 79 -298 125 -287
rect 283 287 329 298
rect 283 -298 329 -287
rect 487 287 533 298
rect 487 -298 533 -287
rect 691 287 737 298
rect 691 -298 737 -287
rect 895 287 941 298
rect 895 -298 941 -287
rect 1099 287 1145 298
rect 1099 -298 1145 -287
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 3 l 0.5 m 1 nf 11 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
