* NGSPICE file created from nmos_3p3_Z2JHD6_flat.ext - technology: gf180mcuC

.subckt nmos_3p3_Z2JHD6_flat
X0 a_0_n209# a_n181_1498.t38 a_n181_1498.t39 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_0_n209# a_n181_1498.t61 a_212_1351.t18 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X2 a_0_n209# a_n181_1498.t63 a_212_1351.t16 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X3 a_0_n209# a_n181_1498.t36 a_n181_1498.t37 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X4 a_0_n209# a_n181_1498.t64 a_212_1351.t15 a_0_n209# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X5 a_0_n209# a_n181_1498.t34 a_n181_1498.t35 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X6 a_0_n209# a_n181_1498.t65 a_212_1351.t14 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X7 a_0_n209# a_n181_1498.t30 a_n181_1498.t31 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X8 a_0_n209# a_n181_1498.t26 a_n181_1498.t27 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X9 a_0_n209# a_n181_1498.t20 a_n181_1498.t21 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X10 a_0_n209# a_n181_1498.t74 a_212_1351.t10 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X11 a_2048_1351# a_24_587.t54 a_212_1351.t39 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X12 a_0_n209# a_n181_1498.t14 a_n181_1498.t15 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X13 a_0_n209# a_n181_1498.t76 a_212_1351.t9 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X14 a_0_n209# a_n181_1498.t12 a_n181_1498.t13 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X15 a_0_n209# a_n181_1498.t78 a_212_1351.t7 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X16 a_0_n209# a_n181_1498.t80 a_212_1351.t6 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X17 a_0_n209# a_n181_1498.t6 a_n181_1498.t7 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X18 a_0_n209# a_n181_1498.t83 a_212_1351.t5 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X19 a_0_n209# a_n181_1498.t87 a_212_1351.t2 a_0_n209# nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X20 a_0_n209# a_n181_1498.t0 a_n181_1498.t1 a_0_n209# nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
R0 a_24_587.n74 a_24_587.t52 120.174
R1 a_24_587.n81 a_24_587.t60 120.174
R2 a_24_587.n16 a_24_587.n15 106.159
R3 a_24_587.n110 a_24_587.n109 106.159
R4 a_24_587.n60 a_24_587.n59 103.823
R5 a_24_587.n115 a_24_587.n114 103.823
R6 a_24_587.n76 a_24_587.n75 103.823
R7 a_24_587.n83 a_24_587.n82 103.823
R8 a_24_587.n89 a_24_587.n88 103.823
R9 a_24_587.n29 a_24_587.n28 103.823
R10 a_24_587.n42 a_24_587.n41 103.823
R11 a_24_587.n21 a_24_587.n20 103.823
R12 a_24_587.n88 a_24_587.t67 37.2224
R13 a_24_587.n28 a_24_587.t59 37.2224
R14 a_24_587.n75 a_24_587.n74 21.0894
R15 a_24_587.n77 a_24_587.n76 21.0894
R16 a_24_587.n82 a_24_587.n81 21.0894
R17 a_24_587.n84 a_24_587.n83 21.0894
R18 a_24_587.n30 a_24_587.n29 21.0894
R19 a_24_587.n97 a_24_587.n96 21.0894
R20 a_24_587.n90 a_24_587.n89 21.0894
R21 a_24_587.n74 a_24_587.t62 16.3525
R22 a_24_587.n75 a_24_587.t44 16.3525
R23 a_24_587.n76 a_24_587.t42 16.3525
R24 a_24_587.n81 a_24_587.t49 16.3525
R25 a_24_587.n82 a_24_587.t68 16.3525
R26 a_24_587.n83 a_24_587.t66 16.3525
R27 a_24_587.n88 a_24_587.t57 16.1335
R28 a_24_587.n89 a_24_587.t45 16.1335
R29 a_24_587.n28 a_24_587.t43 16.1335
R30 a_24_587.n29 a_24_587.t65 16.1335
R31 a_24_587.n96 a_24_587.t54 16.1335
R32 a_24_587.n15 a_24_587.t10 14.0165
R33 a_24_587.n17 a_24_587.t32 14.0165
R34 a_24_587.n19 a_24_587.t16 14.0165
R35 a_24_587.n109 a_24_587.t38 14.0165
R36 a_24_587.n113 a_24_587.t28 14.0165
R37 a_24_587.n105 a_24_587.t20 14.0165
R38 a_24_587.n22 a_24_587.t36 14.0165
R39 a_24_587.n111 a_24_587.t14 13.9435
R40 a_24_587.n38 a_24_587.t22 13.7975
R41 a_24_587.n40 a_24_587.t4 13.7975
R42 a_24_587.n56 a_24_587.t8 13.7975
R43 a_24_587.n58 a_24_587.t26 13.7975
R44 a_24_587.n51 a_24_587.t34 13.7975
R45 a_24_587.n70 a_24_587.t30 13.7975
R46 a_24_587.n43 a_24_587.t24 13.7975
R47 a_24_587.n85 a_24_587.t48 13.3985
R48 a_24_587.n78 a_24_587.t50 13.3702
R49 a_24_587.n25 a_24_587.t0 12.7453
R50 a_24_587.n53 a_24_587.t18 12.5263
R51 a_24_587.n92 a_24_587.t64 12.5263
R52 a_24_587.n32 a_24_587.t47 12.4812
R53 a_24_587.n99 a_24_587.t58 12.4812
R54 a_24_587.n65 a_24_587.t12 12.4795
R55 a_24_587.n45 a_24_587.t6 12.4359
R56 a_24_587.n117 a_24_587.t2 11.6805
R57 a_24_587.n15 a_24_587.n14 9.23263
R58 a_24_587.n109 a_24_587.t39 9.23263
R59 a_24_587.n18 a_24_587.n17 4.15465
R60 a_24_587.n19 a_24_587.n18 4.15465
R61 a_24_587.n39 a_24_587.n38 4.15465
R62 a_24_587.n40 a_24_587.n39 4.15465
R63 a_24_587.n57 a_24_587.n56 4.15465
R64 a_24_587.n58 a_24_587.n57 4.15465
R65 a_24_587.n52 a_24_587.n51 4.15465
R66 a_24_587.n112 a_24_587.n111 4.15465
R67 a_24_587.n113 a_24_587.n112 4.15465
R68 a_24_587.n106 a_24_587.n105 4.15465
R69 a_24_587.n71 a_24_587.n70 4.15465
R70 a_24_587.n44 a_24_587.n43 4.15465
R71 a_24_587.n120 a_24_587.n22 4.15465
R72 a_24_587.n86 a_24_587.n85 3.75668
R73 a_24_587.n79 a_24_587.n78 3.75431
R74 a_24_587.n9 a_24_587.n31 3.549
R75 a_24_587.n11 a_24_587.n91 3.51322
R76 a_24_587.n7 a_24_587.n64 3.50928
R77 a_24_587.n3 a_24_587.n53 3.50535
R78 a_24_587.n1 a_24_587.n116 3.50535
R79 a_24_587.n11 a_24_587.n92 3.50535
R80 a_24_587.n10 a_24_587.n98 3.49926
R81 a_24_587.n7 a_24_587.n65 3.49877
R82 a_24_587.n9 a_24_587.n32 3.4914
R83 a_24_587.n10 a_24_587.n99 3.4914
R84 a_24_587.n0 a_24_587.n45 3.47756
R85 a_24_587.n18 a_24_587.n13 3.43811
R86 a_24_587.n106 a_24_587.n103 3.43811
R87 a_24_587.n122 a_24_587.n120 3.43811
R88 a_24_587.n112 a_24_587.n108 3.43615
R89 a_24_587.n39 a_24_587.n37 3.43224
R90 a_24_587.n57 a_24_587.n55 3.43224
R91 a_24_587.n52 a_24_587.n49 3.43224
R92 a_24_587.n71 a_24_587.n68 3.43224
R93 a_24_587.n44 a_24_587.n35 3.43224
R94 a_24_587.n119 a_24_587.n1 3.26782
R95 a_24_587.n73 a_24_587.n0 2.90675
R96 a_24_587.n11 a_24_587.n93 2.88464
R97 a_24_587.n9 a_24_587.n33 2.88464
R98 a_24_587.n10 a_24_587.n100 2.88464
R99 a_24_587.n0 a_24_587.n47 2.88464
R100 a_24_587.n1 a_24_587.n118 2.88451
R101 a_24_587.n3 a_24_587.n61 2.88438
R102 a_24_587.n62 a_24_587.n3 2.87461
R103 a_24_587.n7 a_24_587.n66 2.8741
R104 a_24_587.n111 a_24_587.n110 2.4095
R105 a_24_587.n17 a_24_587.n16 2.3365
R106 a_24_587.n20 a_24_587.n19 2.3365
R107 a_24_587.n41 a_24_587.n40 2.3365
R108 a_24_587.n59 a_24_587.n58 2.3365
R109 a_24_587.n51 a_24_587.n50 2.3365
R110 a_24_587.n114 a_24_587.n113 2.3365
R111 a_24_587.n105 a_24_587.n104 2.3365
R112 a_24_587.n70 a_24_587.n69 2.3365
R113 a_24_587.n47 a_24_587.n46 2.3365
R114 a_24_587.n43 a_24_587.n42 2.3365
R115 a_24_587.n22 a_24_587.n21 2.3365
R116 a_24_587.n61 a_24_587.n60 2.2635
R117 a_24_587.n118 a_24_587.n117 2.2635
R118 a_24_587.n2 a_24_587.n9 2.2525
R119 a_24_587.n95 a_24_587.n11 2.2515
R120 a_24_587.n101 a_24_587.n10 2.2515
R121 a_24_587.n72 a_24_587.n7 2.2505
R122 a_24_587.n8 a_24_587.n6 2.2505
R123 a_24_587.n26 a_24_587.n24 2.1905
R124 a_24_587.n8 a_24_587.n26 2.11497
R125 a_24_587.n78 a_24_587.n77 1.92893
R126 a_24_587.n85 a_24_587.n84 1.9031
R127 a_24_587.n13 a_24_587.t33 1.6385
R128 a_24_587.n13 a_24_587.n12 1.6385
R129 a_24_587.n37 a_24_587.t23 1.6385
R130 a_24_587.n37 a_24_587.n36 1.6385
R131 a_24_587.n55 a_24_587.t27 1.6385
R132 a_24_587.n55 a_24_587.n54 1.6385
R133 a_24_587.n49 a_24_587.t35 1.6385
R134 a_24_587.n49 a_24_587.n48 1.6385
R135 a_24_587.n108 a_24_587.t29 1.6385
R136 a_24_587.n108 a_24_587.n107 1.6385
R137 a_24_587.n103 a_24_587.t21 1.6385
R138 a_24_587.n103 a_24_587.n102 1.6385
R139 a_24_587.n68 a_24_587.t31 1.6385
R140 a_24_587.n68 a_24_587.n67 1.6385
R141 a_24_587.n35 a_24_587.t25 1.6385
R142 a_24_587.n35 a_24_587.n34 1.6385
R143 a_24_587.t37 a_24_587.n122 1.6385
R144 a_24_587.n122 a_24_587.n121 1.6385
R145 a_24_587.n101 a_24_587.n95 1.26753
R146 a_24_587.n6 a_24_587.n73 1.22996
R147 a_24_587.n6 a_24_587.n2 1.18491
R148 a_24_587.n2 a_24_587.n27 1.16205
R149 a_24_587.n80 a_24_587.n79 1.16042
R150 a_24_587.n101 a_24_587.n5 1.12556
R151 a_24_587.n87 a_24_587.n86 1.12469
R152 a_24_587.n116 a_24_587.n115 1.06529
R153 a_24_587.n26 a_24_587.n25 1.06529
R154 a_24_587.n64 a_24_587.n63 1.02542
R155 a_24_587.n98 a_24_587.n97 1.01842
R156 a_24_587.n31 a_24_587.n30 1.00064
R157 a_24_587.n91 a_24_587.n90 0.99056
R158 a_24_587.n95 a_24_587.n94 0.933875
R159 a_24_587.n72 a_24_587.n62 0.652981
R160 a_24_587.n73 a_24_587.n72 0.604805
R161 a_24_587.n119 a_24_587.n101 0.545453
R162 a_24_587.n5 a_24_587.n87 0.543697
R163 a_24_587.n6 a_24_587.n119 0.266683
R164 a_24_587.n4 a_24_587.n80 0.249615
R165 a_24_587.n3 a_24_587.n52 0.156649
R166 a_24_587.n1 a_24_587.n106 0.156649
R167 a_24_587.n120 a_24_587.n8 0.15656
R168 a_24_587.n0 a_24_587.n44 0.155649
R169 a_24_587.n7 a_24_587.n71 0.155577
R170 a_24_587.n24 a_24_587.n23 0.0735
R171 a_24_587.n5 a_24_587.n4 0.0595
R172 a_n181_1498.n0 a_n181_1498.n91 74.2622
R173 a_n181_1498.n1 a_n181_1498.n23 71.202
R174 a_n181_1498.n26 a_n181_1498.t0 37.4414
R175 a_n181_1498.n92 a_n181_1498.t18 37.4414
R176 a_n181_1498.n91 a_n181_1498.n90 21.0894
R177 a_n181_1498.n90 a_n181_1498.n89 21.0894
R178 a_n181_1498.n89 a_n181_1498.n88 21.0894
R179 a_n181_1498.n88 a_n181_1498.n87 21.0894
R180 a_n181_1498.n87 a_n181_1498.n86 21.0894
R181 a_n181_1498.n86 a_n181_1498.n85 21.0894
R182 a_n181_1498.n85 a_n181_1498.n84 21.0894
R183 a_n181_1498.n84 a_n181_1498.n83 21.0894
R184 a_n181_1498.n83 a_n181_1498.n82 21.0894
R185 a_n181_1498.n15 a_n181_1498.n14 21.0894
R186 a_n181_1498.n16 a_n181_1498.n15 21.0894
R187 a_n181_1498.n17 a_n181_1498.n16 21.0894
R188 a_n181_1498.n18 a_n181_1498.n17 21.0894
R189 a_n181_1498.n19 a_n181_1498.n18 21.0894
R190 a_n181_1498.n20 a_n181_1498.n19 21.0894
R191 a_n181_1498.n21 a_n181_1498.n20 21.0894
R192 a_n181_1498.n22 a_n181_1498.n21 21.0894
R193 a_n181_1498.n23 a_n181_1498.n22 21.0894
R194 a_n181_1498.n90 a_n181_1498.t65 16.5715
R195 a_n181_1498.n89 a_n181_1498.t86 16.5715
R196 a_n181_1498.n86 a_n181_1498.t78 16.5715
R197 a_n181_1498.n85 a_n181_1498.t62 16.5715
R198 a_n181_1498.n82 a_n181_1498.t83 16.5715
R199 a_n181_1498.n14 a_n181_1498.t88 16.5715
R200 a_n181_1498.n17 a_n181_1498.t80 16.5715
R201 a_n181_1498.n18 a_n181_1498.t66 16.5715
R202 a_n181_1498.n21 a_n181_1498.t74 16.5715
R203 a_n181_1498.n22 a_n181_1498.t89 16.5715
R204 a_n181_1498.n91 a_n181_1498.t70 16.3525
R205 a_n181_1498.n88 a_n181_1498.t61 16.3525
R206 a_n181_1498.n87 a_n181_1498.t77 16.3525
R207 a_n181_1498.n84 a_n181_1498.t76 16.3525
R208 a_n181_1498.n83 a_n181_1498.t60 16.3525
R209 a_n181_1498.n15 a_n181_1498.t63 16.3525
R210 a_n181_1498.n16 a_n181_1498.t84 16.3525
R211 a_n181_1498.n19 a_n181_1498.t87 16.3525
R212 a_n181_1498.n20 a_n181_1498.t72 16.3525
R213 a_n181_1498.n23 a_n181_1498.t64 16.3525
R214 a_n181_1498.n27 a_n181_1498.t22 14.0165
R215 a_n181_1498.n30 a_n181_1498.t26 14.0165
R216 a_n181_1498.n39 a_n181_1498.t10 14.0165
R217 a_n181_1498.n42 a_n181_1498.t14 14.0165
R218 a_n181_1498.n47 a_n181_1498.t28 14.0165
R219 a_n181_1498.n50 a_n181_1498.t34 14.0165
R220 a_n181_1498.n57 a_n181_1498.t16 14.0165
R221 a_n181_1498.n60 a_n181_1498.t20 14.0165
R222 a_n181_1498.n65 a_n181_1498.t4 14.0165
R223 a_n181_1498.n68 a_n181_1498.t38 14.0165
R224 a_n181_1498.n93 a_n181_1498.t36 14.0165
R225 a_n181_1498.n96 a_n181_1498.t32 14.0165
R226 a_n181_1498.n105 a_n181_1498.t6 14.0165
R227 a_n181_1498.n108 a_n181_1498.t2 14.0165
R228 a_n181_1498.n115 a_n181_1498.t12 14.0165
R229 a_n181_1498.n118 a_n181_1498.t8 14.0165
R230 a_n181_1498.n125 a_n181_1498.t30 14.0165
R231 a_n181_1498.n73 a_n181_1498.t24 14.0165
R232 a_n181_1498.n127 a_n181_1498.n73 4.0005
R233 a_n181_1498.n126 a_n181_1498.n125 4.0005
R234 a_n181_1498.n119 a_n181_1498.n118 4.0005
R235 a_n181_1498.n116 a_n181_1498.n115 4.0005
R236 a_n181_1498.n109 a_n181_1498.n108 4.0005
R237 a_n181_1498.n106 a_n181_1498.n105 4.0005
R238 a_n181_1498.n97 a_n181_1498.n96 4.0005
R239 a_n181_1498.n94 a_n181_1498.n93 4.0005
R240 a_n181_1498.n28 a_n181_1498.n27 4.0005
R241 a_n181_1498.n31 a_n181_1498.n30 4.0005
R242 a_n181_1498.n40 a_n181_1498.n39 4.0005
R243 a_n181_1498.n43 a_n181_1498.n42 4.0005
R244 a_n181_1498.n48 a_n181_1498.n47 4.0005
R245 a_n181_1498.n51 a_n181_1498.n50 4.0005
R246 a_n181_1498.n58 a_n181_1498.n57 4.0005
R247 a_n181_1498.n61 a_n181_1498.n60 4.0005
R248 a_n181_1498.n66 a_n181_1498.n65 4.0005
R249 a_n181_1498.n69 a_n181_1498.n68 4.0005
R250 a_n181_1498.n1 a_n181_1498.n25 3.58493
R251 a_n181_1498.n103 a_n181_1498.n102 3.57898
R252 a_n181_1498.n123 a_n181_1498.n122 3.57507
R253 a_n181_1498.n0 a_n181_1498.n81 3.5665
R254 a_n181_1498.n44 a_n181_1498.n11 3.53988
R255 a_n181_1498.n112 a_n181_1498.n111 3.53861
R256 a_n181_1498.n128 a_n181_1498.n71 3.53721
R257 a_n181_1498.n113 a_n181_1498.n77 3.53202
R258 a_n181_1498.n131 a_n181_1498.n129 3.53202
R259 a_n181_1498.n120 a_n181_1498.n75 3.52224
R260 a_n181_1498.n63 a_n181_1498.n3 3.51637
R261 a_n181_1498.n45 a_n181_1498.n9 3.51246
R262 a_n181_1498.n55 a_n181_1498.n54 3.51057
R263 a_n181_1498.n34 a_n181_1498.n33 3.50854
R264 a_n181_1498.n100 a_n181_1498.n99 3.50645
R265 a_n181_1498.n37 a_n181_1498.n36 3.49699
R266 a_n181_1498.n62 a_n181_1498.n5 3.49116
R267 a_n181_1498.n52 a_n181_1498.n7 3.4806
R268 a_n181_1498.n0 a_n181_1498.n79 3.46399
R269 a_n181_1498.n1 a_n181_1498.n13 3.45496
R270 a_n181_1498.n27 a_n181_1498.n26 2.3365
R271 a_n181_1498.n30 a_n181_1498.n29 2.3365
R272 a_n181_1498.n39 a_n181_1498.n38 2.3365
R273 a_n181_1498.n42 a_n181_1498.n41 2.3365
R274 a_n181_1498.n47 a_n181_1498.n46 2.3365
R275 a_n181_1498.n50 a_n181_1498.n49 2.3365
R276 a_n181_1498.n57 a_n181_1498.n56 2.3365
R277 a_n181_1498.n60 a_n181_1498.n59 2.3365
R278 a_n181_1498.n65 a_n181_1498.n64 2.3365
R279 a_n181_1498.n68 a_n181_1498.n67 2.3365
R280 a_n181_1498.n93 a_n181_1498.n92 2.3365
R281 a_n181_1498.n96 a_n181_1498.n95 2.3365
R282 a_n181_1498.n105 a_n181_1498.n104 2.3365
R283 a_n181_1498.n108 a_n181_1498.n107 2.3365
R284 a_n181_1498.n115 a_n181_1498.n114 2.3365
R285 a_n181_1498.n118 a_n181_1498.n117 2.3365
R286 a_n181_1498.n125 a_n181_1498.n124 2.3365
R287 a_n181_1498.n73 a_n181_1498.n72 2.3365
R288 a_n181_1498.n71 a_n181_1498.t50 1.6385
R289 a_n181_1498.n71 a_n181_1498.n70 1.6385
R290 a_n181_1498.n5 a_n181_1498.t21 1.6385
R291 a_n181_1498.n5 a_n181_1498.n4 1.6385
R292 a_n181_1498.n3 a_n181_1498.t40 1.6385
R293 a_n181_1498.n3 a_n181_1498.n2 1.6385
R294 a_n181_1498.n7 a_n181_1498.t35 1.6385
R295 a_n181_1498.n7 a_n181_1498.n6 1.6385
R296 a_n181_1498.n54 a_n181_1498.t47 1.6385
R297 a_n181_1498.n54 a_n181_1498.n53 1.6385
R298 a_n181_1498.n11 a_n181_1498.t15 1.6385
R299 a_n181_1498.n11 a_n181_1498.n10 1.6385
R300 a_n181_1498.n9 a_n181_1498.t56 1.6385
R301 a_n181_1498.n9 a_n181_1498.n8 1.6385
R302 a_n181_1498.n33 a_n181_1498.t27 1.6385
R303 a_n181_1498.n33 a_n181_1498.n32 1.6385
R304 a_n181_1498.n36 a_n181_1498.t44 1.6385
R305 a_n181_1498.n36 a_n181_1498.n35 1.6385
R306 a_n181_1498.n102 a_n181_1498.t7 1.6385
R307 a_n181_1498.n102 a_n181_1498.n101 1.6385
R308 a_n181_1498.n99 a_n181_1498.t52 1.6385
R309 a_n181_1498.n99 a_n181_1498.n98 1.6385
R310 a_n181_1498.n77 a_n181_1498.t13 1.6385
R311 a_n181_1498.n77 a_n181_1498.n76 1.6385
R312 a_n181_1498.n111 a_n181_1498.t57 1.6385
R313 a_n181_1498.n111 a_n181_1498.n110 1.6385
R314 a_n181_1498.n122 a_n181_1498.t31 1.6385
R315 a_n181_1498.n122 a_n181_1498.n121 1.6385
R316 a_n181_1498.n75 a_n181_1498.t43 1.6385
R317 a_n181_1498.n75 a_n181_1498.n74 1.6385
R318 a_n181_1498.n79 a_n181_1498.t37 1.6385
R319 a_n181_1498.n79 a_n181_1498.n78 1.6385
R320 a_n181_1498.n81 a_n181_1498.t48 1.6385
R321 a_n181_1498.n81 a_n181_1498.n80 1.6385
R322 a_n181_1498.n13 a_n181_1498.t49 1.6385
R323 a_n181_1498.n13 a_n181_1498.n12 1.6385
R324 a_n181_1498.n25 a_n181_1498.t1 1.6385
R325 a_n181_1498.n25 a_n181_1498.n24 1.6385
R326 a_n181_1498.t39 a_n181_1498.n131 1.6385
R327 a_n181_1498.n131 a_n181_1498.n130 1.6385
R328 a_n181_1498.n94 a_n181_1498.n0 0.373787
R329 a_n181_1498.n127 a_n181_1498.n126 0.253351
R330 a_n181_1498.n119 a_n181_1498.n116 0.197599
R331 a_n181_1498.n97 a_n181_1498.n94 0.197599
R332 a_n181_1498.n31 a_n181_1498.n28 0.197599
R333 a_n181_1498.n51 a_n181_1498.n48 0.197599
R334 a_n181_1498.n69 a_n181_1498.n66 0.197599
R335 a_n181_1498.n109 a_n181_1498.n106 0.172031
R336 a_n181_1498.n43 a_n181_1498.n40 0.172031
R337 a_n181_1498.n61 a_n181_1498.n58 0.172031
R338 a_n181_1498.n37 a_n181_1498.n34 0.100499
R339 a_n181_1498.n45 a_n181_1498.n44 0.093148
R340 a_n181_1498.n63 a_n181_1498.n62 0.0926899
R341 a_n181_1498.n55 a_n181_1498.n52 0.0817532
R342 a_n181_1498.n123 a_n181_1498.n120 0.0807174
R343 a_n181_1498.n129 a_n181_1498.n128 0.0742956
R344 a_n181_1498.n113 a_n181_1498.n112 0.0727632
R345 a_n181_1498.n129 a_n181_1498.n69 0.0708476
R346 a_n181_1498.n116 a_n181_1498.n113 0.0705535
R347 a_n181_1498.n103 a_n181_1498.n100 0.0688207
R348 a_n181_1498.n100 a_n181_1498.n97 0.0665096
R349 a_n181_1498.n120 a_n181_1498.n119 0.0655603
R350 a_n181_1498.n66 a_n181_1498.n63 0.0636092
R351 a_n181_1498.n52 a_n181_1498.n51 0.061636
R352 a_n181_1498.n48 a_n181_1498.n45 0.0606109
R353 a_n181_1498.n34 a_n181_1498.n31 0.0579026
R354 a_n181_1498.n106 a_n181_1498.n103 0.049875
R355 a_n181_1498.n126 a_n181_1498.n123 0.0488673
R356 a_n181_1498.n112 a_n181_1498.n109 0.0443624
R357 a_n181_1498.n44 a_n181_1498.n43 0.0432184
R358 a_n181_1498.n128 a_n181_1498.n127 0.0423084
R359 a_n181_1498.n58 a_n181_1498.n55 0.0409019
R360 a_n181_1498.n62 a_n181_1498.n61 0.0397098
R361 a_n181_1498.n40 a_n181_1498.n37 0.0396398
R362 a_n181_1498.n28 a_n181_1498.n1 0.0267736
R363 a_212_1351.n43 a_212_1351.n42 3.5788
R364 a_212_1351.n23 a_212_1351.n22 3.18472
R365 a_212_1351.n0 a_212_1351.n14 3.17597
R366 a_212_1351.n5 a_212_1351.n12 3.17588
R367 a_212_1351.n4 a_212_1351.n10 3.17454
R368 a_212_1351.n2 a_212_1351.n36 3.1741
R369 a_212_1351.n24 a_212_1351.n18 3.17375
R370 a_212_1351.n57 a_212_1351.n1 3.17351
R371 a_212_1351.n3 a_212_1351.n34 3.17318
R372 a_212_1351.n6 a_212_1351.n38 3.17219
R373 a_212_1351.n4 a_212_1351.n8 2.93559
R374 a_212_1351.n43 a_212_1351.n40 2.57385
R375 a_212_1351.n23 a_212_1351.n20 2.56337
R376 a_212_1351.n25 a_212_1351.n16 2.56302
R377 a_212_1351.n6 a_212_1351.n47 2.24989
R378 a_212_1351.n5 a_212_1351.n31 2.24988
R379 a_212_1351.n0 a_212_1351.n28 2.24511
R380 a_212_1351.n2 a_212_1351.n50 2.24483
R381 a_212_1351.n1 a_212_1351.n56 2.24483
R382 a_212_1351.n3 a_212_1351.n53 2.24455
R383 a_212_1351.n46 a_212_1351.n45 1.74882
R384 a_212_1351.n55 a_212_1351.n54 1.74881
R385 a_212_1351.n49 a_212_1351.n48 1.74881
R386 a_212_1351.n30 a_212_1351.n29 1.74881
R387 a_212_1351.n16 a_212_1351.n15 1.74881
R388 a_212_1351.n40 a_212_1351.n39 1.73463
R389 a_212_1351.n27 a_212_1351.n26 1.73459
R390 a_212_1351.n52 a_212_1351.t21 1.6385
R391 a_212_1351.n52 a_212_1351.n51 1.6385
R392 a_212_1351.n42 a_212_1351.t20 1.6385
R393 a_212_1351.n42 a_212_1351.n41 1.6385
R394 a_212_1351.n38 a_212_1351.t18 1.6385
R395 a_212_1351.n38 a_212_1351.n37 1.6385
R396 a_212_1351.n36 a_212_1351.t26 1.6385
R397 a_212_1351.n36 a_212_1351.n35 1.6385
R398 a_212_1351.n34 a_212_1351.t9 1.6385
R399 a_212_1351.n34 a_212_1351.n33 1.6385
R400 a_212_1351.n8 a_212_1351.t23 1.6385
R401 a_212_1351.n8 a_212_1351.n7 1.6385
R402 a_212_1351.n20 a_212_1351.t22 1.6385
R403 a_212_1351.n20 a_212_1351.n19 1.6385
R404 a_212_1351.n22 a_212_1351.t15 1.6385
R405 a_212_1351.n22 a_212_1351.n21 1.6385
R406 a_212_1351.n18 a_212_1351.t28 1.6385
R407 a_212_1351.n18 a_212_1351.n17 1.6385
R408 a_212_1351.n14 a_212_1351.t2 1.6385
R409 a_212_1351.n14 a_212_1351.n13 1.6385
R410 a_212_1351.n12 a_212_1351.t25 1.6385
R411 a_212_1351.n12 a_212_1351.n11 1.6385
R412 a_212_1351.n10 a_212_1351.t16 1.6385
R413 a_212_1351.n10 a_212_1351.n9 1.6385
R414 a_212_1351.n57 a_212_1351.t39 1.6385
R415 a_212_1351.n58 a_212_1351.n57 1.6385
R416 a_212_1351.n27 a_212_1351.t27 1.48949
R417 a_212_1351.n40 a_212_1351.t14 1.48945
R418 a_212_1351.n55 a_212_1351.t5 1.47237
R419 a_212_1351.n49 a_212_1351.t7 1.47237
R420 a_212_1351.n30 a_212_1351.t6 1.47237
R421 a_212_1351.n16 a_212_1351.t10 1.47237
R422 a_212_1351.n46 a_212_1351.t24 1.47236
R423 a_212_1351.n53 a_212_1351.n52 1.44171
R424 a_212_1351.n47 a_212_1351.n46 1.07211
R425 a_212_1351.n50 a_212_1351.n49 1.07199
R426 a_212_1351.n31 a_212_1351.n30 1.07199
R427 a_212_1351.n56 a_212_1351.n55 1.07199
R428 a_212_1351.n28 a_212_1351.n27 1.07053
R429 a_212_1351.n1 a_212_1351.n4 0.631039
R430 a_212_1351.n0 a_212_1351.n25 0.626751
R431 a_212_1351.n2 a_212_1351.n6 0.623731
R432 a_212_1351.n24 a_212_1351.n23 0.622777
R433 a_212_1351.n5 a_212_1351.n0 0.622133
R434 a_212_1351.n1 a_212_1351.n3 0.619295
R435 a_212_1351.n3 a_212_1351.n2 0.606132
R436 a_212_1351.n4 a_212_1351.n32 0.601448
R437 a_212_1351.n44 a_212_1351.n43 0.597765
R438 a_212_1351.n32 a_212_1351.n5 0.0291239
R439 a_212_1351.n6 a_212_1351.n44 0.0287767
R440 a_212_1351.n25 a_212_1351.n24 0.0264198
R441 a_24_1802.n22 a_24_1802.n0 5.71342
R442 a_24_1802.n15 a_24_1802.t6 5.71342
R443 a_24_1802.n15 a_24_1802.n14 3.54572
R444 a_24_1802.n17 a_24_1802.n10 3.54572
R445 a_24_1802.n20 a_24_1802.n4 3.54572
R446 a_24_1802.n23 a_24_1802.n22 3.54572
R447 a_24_1802.n21 a_24_1802.n2 3.5105
R448 a_24_1802.n19 a_24_1802.n6 3.5105
R449 a_24_1802.n18 a_24_1802.n8 3.5105
R450 a_24_1802.n16 a_24_1802.n12 3.5105
R451 a_24_1802.n2 a_24_1802.t5 1.6385
R452 a_24_1802.n2 a_24_1802.n1 1.6385
R453 a_24_1802.n6 a_24_1802.t17 1.6385
R454 a_24_1802.n6 a_24_1802.n5 1.6385
R455 a_24_1802.n8 a_24_1802.t12 1.6385
R456 a_24_1802.n8 a_24_1802.n7 1.6385
R457 a_24_1802.n12 a_24_1802.t0 1.6385
R458 a_24_1802.n12 a_24_1802.n11 1.6385
R459 a_24_1802.n14 a_24_1802.t8 1.6385
R460 a_24_1802.n14 a_24_1802.n13 1.6385
R461 a_24_1802.n10 a_24_1802.t4 1.6385
R462 a_24_1802.n10 a_24_1802.n9 1.6385
R463 a_24_1802.n4 a_24_1802.t3 1.6385
R464 a_24_1802.n4 a_24_1802.n3 1.6385
R465 a_24_1802.n23 a_24_1802.t7 1.6385
R466 a_24_1802.n24 a_24_1802.n23 1.6385
R467 a_24_1802.n19 a_24_1802.n18 1.13035
R468 a_24_1802.n22 a_24_1802.n21 0.565423
R469 a_24_1802.n21 a_24_1802.n20 0.565423
R470 a_24_1802.n20 a_24_1802.n19 0.565423
R471 a_24_1802.n18 a_24_1802.n17 0.565423
R472 a_24_1802.n17 a_24_1802.n16 0.565423
R473 a_24_1802.n16 a_24_1802.n15 0.565423
C0 m1_n442_2771# a_0_n209# 0.115f $ **FLOATING
C1 a_2048_1351# a_0_n209# 0.0434f
C2 a_24_1802.t7 a_0_n209# 0.0198f
C3 a_24_1802.n0 a_0_n209# 0.0661f
C4 a_24_1802.t5 a_0_n209# 0.0198f
C5 a_24_1802.n1 a_0_n209# 0.0198f
C6 a_24_1802.n2 a_0_n209# 0.0431f
C7 a_24_1802.t3 a_0_n209# 0.0198f
C8 a_24_1802.n3 a_0_n209# 0.0198f
C9 a_24_1802.n4 a_0_n209# 0.0436f
C10 a_24_1802.t17 a_0_n209# 0.0198f
C11 a_24_1802.n5 a_0_n209# 0.0198f
C12 a_24_1802.n6 a_0_n209# 0.0431f
C13 a_24_1802.t12 a_0_n209# 0.0198f
C14 a_24_1802.n7 a_0_n209# 0.0198f
C15 a_24_1802.n8 a_0_n209# 0.0431f
C16 a_24_1802.t4 a_0_n209# 0.0198f
C17 a_24_1802.n9 a_0_n209# 0.0198f
C18 a_24_1802.n10 a_0_n209# 0.0436f
C19 a_24_1802.t0 a_0_n209# 0.0198f
C20 a_24_1802.n11 a_0_n209# 0.0198f
C21 a_24_1802.n12 a_0_n209# 0.0431f
C22 a_24_1802.t8 a_0_n209# 0.0198f
C23 a_24_1802.n13 a_0_n209# 0.0198f
C24 a_24_1802.n14 a_0_n209# 0.0436f
C25 a_24_1802.t6 a_0_n209# 0.0661f
C26 a_24_1802.n15 a_0_n209# 0.257f
C27 a_24_1802.n16 a_0_n209# 0.147f
C28 a_24_1802.n17 a_0_n209# 0.15f
C29 a_24_1802.n18 a_0_n209# 0.198f
C30 a_24_1802.n19 a_0_n209# 0.198f
C31 a_24_1802.n20 a_0_n209# 0.15f
C32 a_24_1802.n21 a_0_n209# 0.147f
C33 a_24_1802.n22 a_0_n209# 0.257f
C34 a_24_1802.n23 a_0_n209# 0.0436f
C35 a_24_1802.n24 a_0_n209# 0.0198f
C36 a_212_1351.n0 a_0_n209# 0.109f
C37 a_212_1351.n1 a_0_n209# 0.109f
C38 a_212_1351.n2 a_0_n209# 0.109f
C39 a_212_1351.n3 a_0_n209# 0.108f
C40 a_212_1351.n4 a_0_n209# 0.119f
C41 a_212_1351.n5 a_0_n209# 0.0849f
C42 a_212_1351.n6 a_0_n209# 0.0849f
C43 a_212_1351.t39 a_0_n209# 0.0106f
C44 a_212_1351.t23 a_0_n209# 0.0106f
C45 a_212_1351.n7 a_0_n209# 0.0106f
C46 a_212_1351.n8 a_0_n209# 0.0328f
C47 a_212_1351.t16 a_0_n209# 0.0106f
C48 a_212_1351.n9 a_0_n209# 0.0106f
C49 a_212_1351.n10 a_0_n209# 0.04f
C50 a_212_1351.t25 a_0_n209# 0.0106f
C51 a_212_1351.n11 a_0_n209# 0.0106f
C52 a_212_1351.n12 a_0_n209# 0.04f
C53 a_212_1351.t2 a_0_n209# 0.0106f
C54 a_212_1351.n13 a_0_n209# 0.0106f
C55 a_212_1351.n14 a_0_n209# 0.04f
C56 a_212_1351.t10 a_0_n209# 0.00993f
C57 a_212_1351.n15 a_0_n209# 0.0116f
C58 a_212_1351.n16 a_0_n209# 0.0342f
C59 a_212_1351.t28 a_0_n209# 0.0106f
C60 a_212_1351.n17 a_0_n209# 0.0106f
C61 a_212_1351.n18 a_0_n209# 0.0399f
C62 a_212_1351.t22 a_0_n209# 0.0106f
C63 a_212_1351.n19 a_0_n209# 0.0106f
C64 a_212_1351.n20 a_0_n209# 0.0312f
C65 a_212_1351.t15 a_0_n209# 0.0106f
C66 a_212_1351.n21 a_0_n209# 0.0106f
C67 a_212_1351.n22 a_0_n209# 0.0402f
C68 a_212_1351.n23 a_0_n209# 0.101f
C69 a_212_1351.n24 a_0_n209# 0.0802f
C70 a_212_1351.n25 a_0_n209# 0.0302f
C71 a_212_1351.t27 a_0_n209# 0.01f
C72 a_212_1351.n26 a_0_n209# 0.0115f
C73 a_212_1351.n27 a_0_n209# 0.0211f
C74 a_212_1351.n28 a_0_n209# 0.0225f
C75 a_212_1351.t6 a_0_n209# 0.00993f
C76 a_212_1351.n29 a_0_n209# 0.0116f
C77 a_212_1351.n30 a_0_n209# 0.021f
C78 a_212_1351.n31 a_0_n209# 0.0225f
C79 a_212_1351.n32 a_0_n209# 0.0236f
C80 a_212_1351.t9 a_0_n209# 0.0106f
C81 a_212_1351.n33 a_0_n209# 0.0106f
C82 a_212_1351.n34 a_0_n209# 0.04f
C83 a_212_1351.t26 a_0_n209# 0.0106f
C84 a_212_1351.n35 a_0_n209# 0.0106f
C85 a_212_1351.n36 a_0_n209# 0.0399f
C86 a_212_1351.t18 a_0_n209# 0.0106f
C87 a_212_1351.n37 a_0_n209# 0.0106f
C88 a_212_1351.n38 a_0_n209# 0.0399f
C89 a_212_1351.n39 a_0_n209# 0.0115f
C90 a_212_1351.t14 a_0_n209# 0.01f
C91 a_212_1351.n40 a_0_n209# 0.0342f
C92 a_212_1351.t20 a_0_n209# 0.0106f
C93 a_212_1351.n41 a_0_n209# 0.0106f
C94 a_212_1351.n42 a_0_n209# 0.0403f
C95 a_212_1351.n43 a_0_n209# 0.0964f
C96 a_212_1351.n44 a_0_n209# 0.0242f
C97 a_212_1351.t24 a_0_n209# 0.00993f
C98 a_212_1351.n45 a_0_n209# 0.0116f
C99 a_212_1351.n46 a_0_n209# 0.0211f
C100 a_212_1351.n47 a_0_n209# 0.0225f
C101 a_212_1351.t7 a_0_n209# 0.00993f
C102 a_212_1351.n48 a_0_n209# 0.0116f
C103 a_212_1351.n49 a_0_n209# 0.021f
C104 a_212_1351.n50 a_0_n209# 0.0225f
C105 a_212_1351.t21 a_0_n209# 0.0106f
C106 a_212_1351.n51 a_0_n209# 0.0106f
C107 a_212_1351.n52 a_0_n209# 0.0214f
C108 a_212_1351.n53 a_0_n209# 0.0225f
C109 a_212_1351.t5 a_0_n209# 0.00993f
C110 a_212_1351.n54 a_0_n209# 0.0116f
C111 a_212_1351.n55 a_0_n209# 0.021f
C112 a_212_1351.n56 a_0_n209# 0.0225f
C113 a_212_1351.n57 a_0_n209# 0.04f
C114 a_212_1351.n58 a_0_n209# 0.0106f
C115 a_n181_1498.n0 a_0_n209# 0.359f
C116 a_n181_1498.n1 a_0_n209# 0.362f
C117 a_n181_1498.t40 a_0_n209# 0.0105f
C118 a_n181_1498.n2 a_0_n209# 0.0105f
C119 a_n181_1498.n3 a_0_n209# 0.0228f
C120 a_n181_1498.t21 a_0_n209# 0.0105f
C121 a_n181_1498.n4 a_0_n209# 0.0105f
C122 a_n181_1498.n5 a_0_n209# 0.0227f
C123 a_n181_1498.t35 a_0_n209# 0.0105f
C124 a_n181_1498.n6 a_0_n209# 0.0105f
C125 a_n181_1498.n7 a_0_n209# 0.0226f
C126 a_n181_1498.t56 a_0_n209# 0.0105f
C127 a_n181_1498.n8 a_0_n209# 0.0105f
C128 a_n181_1498.n9 a_0_n209# 0.0228f
C129 a_n181_1498.t15 a_0_n209# 0.0105f
C130 a_n181_1498.n10 a_0_n209# 0.0105f
C131 a_n181_1498.n11 a_0_n209# 0.0231f
C132 a_n181_1498.t49 a_0_n209# 0.0105f
C133 a_n181_1498.n12 a_0_n209# 0.0105f
C134 a_n181_1498.n13 a_0_n209# 0.0226f
C135 a_n181_1498.t88 a_0_n209# 0.0342f
C136 a_n181_1498.n14 a_0_n209# 0.0341f
C137 a_n181_1498.t63 a_0_n209# 0.0339f
C138 a_n181_1498.n15 a_0_n209# 0.0338f
C139 a_n181_1498.t84 a_0_n209# 0.0339f
C140 a_n181_1498.n16 a_0_n209# 0.0338f
C141 a_n181_1498.t80 a_0_n209# 0.0342f
C142 a_n181_1498.n17 a_0_n209# 0.0341f
C143 a_n181_1498.t66 a_0_n209# 0.0342f
C144 a_n181_1498.n18 a_0_n209# 0.0341f
C145 a_n181_1498.t87 a_0_n209# 0.0339f
C146 a_n181_1498.n19 a_0_n209# 0.0338f
C147 a_n181_1498.t72 a_0_n209# 0.0339f
C148 a_n181_1498.n20 a_0_n209# 0.0338f
C149 a_n181_1498.t74 a_0_n209# 0.0342f
C150 a_n181_1498.n21 a_0_n209# 0.0341f
C151 a_n181_1498.t89 a_0_n209# 0.0342f
C152 a_n181_1498.n22 a_0_n209# 0.0341f
C153 a_n181_1498.t64 a_0_n209# 0.0339f
C154 a_n181_1498.n23 a_0_n209# 0.047f
C155 a_n181_1498.t1 a_0_n209# 0.0105f
C156 a_n181_1498.n24 a_0_n209# 0.0105f
C157 a_n181_1498.n25 a_0_n209# 0.0234f
C158 a_n181_1498.t22 a_0_n209# 0.0307f
C159 a_n181_1498.t0 a_0_n209# 0.0508f
C160 a_n181_1498.n26 a_0_n209# 0.0275f
C161 a_n181_1498.n27 a_0_n209# 0.0226f
C162 a_n181_1498.n28 a_0_n209# 0.0216f
C163 a_n181_1498.t26 a_0_n209# 0.0307f
C164 a_n181_1498.n29 a_0_n209# 0.0144f
C165 a_n181_1498.n30 a_0_n209# 0.0226f
C166 a_n181_1498.n31 a_0_n209# 0.0289f
C167 a_n181_1498.t27 a_0_n209# 0.0105f
C168 a_n181_1498.n32 a_0_n209# 0.0105f
C169 a_n181_1498.n33 a_0_n209# 0.0228f
C170 a_n181_1498.n34 a_0_n209# 0.0377f
C171 a_n181_1498.t44 a_0_n209# 0.0105f
C172 a_n181_1498.n35 a_0_n209# 0.0105f
C173 a_n181_1498.n36 a_0_n209# 0.0228f
C174 a_n181_1498.n37 a_0_n209# 0.0439f
C175 a_n181_1498.n38 a_0_n209# 0.0144f
C176 a_n181_1498.t10 a_0_n209# 0.0307f
C177 a_n181_1498.n39 a_0_n209# 0.0226f
C178 a_n181_1498.n40 a_0_n209# 0.0335f
C179 a_n181_1498.n41 a_0_n209# 0.0144f
C180 a_n181_1498.t14 a_0_n209# 0.0307f
C181 a_n181_1498.n42 a_0_n209# 0.0226f
C182 a_n181_1498.n43 a_0_n209# 0.0345f
C183 a_n181_1498.n44 a_0_n209# 0.0418f
C184 a_n181_1498.n45 a_0_n209# 0.0374f
C185 a_n181_1498.t28 a_0_n209# 0.0307f
C186 a_n181_1498.n46 a_0_n209# 0.0144f
C187 a_n181_1498.n47 a_0_n209# 0.0226f
C188 a_n181_1498.n48 a_0_n209# 0.0282f
C189 a_n181_1498.t34 a_0_n209# 0.0307f
C190 a_n181_1498.n49 a_0_n209# 0.0144f
C191 a_n181_1498.n50 a_0_n209# 0.0226f
C192 a_n181_1498.n51 a_0_n209# 0.0264f
C193 a_n181_1498.n52 a_0_n209# 0.0377f
C194 a_n181_1498.t47 a_0_n209# 0.0105f
C195 a_n181_1498.n53 a_0_n209# 0.0105f
C196 a_n181_1498.n54 a_0_n209# 0.0229f
C197 a_n181_1498.n55 a_0_n209# 0.0432f
C198 a_n181_1498.n56 a_0_n209# 0.0144f
C199 a_n181_1498.t16 a_0_n209# 0.0307f
C200 a_n181_1498.n57 a_0_n209# 0.0226f
C201 a_n181_1498.n58 a_0_n209# 0.0338f
C202 a_n181_1498.n59 a_0_n209# 0.0144f
C203 a_n181_1498.t20 a_0_n209# 0.0307f
C204 a_n181_1498.n60 a_0_n209# 0.0226f
C205 a_n181_1498.n61 a_0_n209# 0.0334f
C206 a_n181_1498.n62 a_0_n209# 0.0438f
C207 a_n181_1498.n63 a_0_n209# 0.0374f
C208 a_n181_1498.t4 a_0_n209# 0.0307f
C209 a_n181_1498.n64 a_0_n209# 0.0144f
C210 a_n181_1498.n65 a_0_n209# 0.0226f
C211 a_n181_1498.n66 a_0_n209# 0.0276f
C212 a_n181_1498.t38 a_0_n209# 0.0307f
C213 a_n181_1498.n67 a_0_n209# 0.0144f
C214 a_n181_1498.n68 a_0_n209# 0.0226f
C215 a_n181_1498.n69 a_0_n209# 0.0272f
C216 a_n181_1498.t50 a_0_n209# 0.0105f
C217 a_n181_1498.n70 a_0_n209# 0.0105f
C218 a_n181_1498.n71 a_0_n209# 0.023f
C219 a_n181_1498.n72 a_0_n209# 0.0144f
C220 a_n181_1498.t24 a_0_n209# 0.0307f
C221 a_n181_1498.n73 a_0_n209# 0.0226f
C222 a_n181_1498.t43 a_0_n209# 0.0105f
C223 a_n181_1498.n74 a_0_n209# 0.0105f
C224 a_n181_1498.n75 a_0_n209# 0.0229f
C225 a_n181_1498.t13 a_0_n209# 0.0105f
C226 a_n181_1498.n76 a_0_n209# 0.0105f
C227 a_n181_1498.n77 a_0_n209# 0.023f
C228 a_n181_1498.t37 a_0_n209# 0.0105f
C229 a_n181_1498.n78 a_0_n209# 0.0105f
C230 a_n181_1498.n79 a_0_n209# 0.0226f
C231 a_n181_1498.t48 a_0_n209# 0.0105f
C232 a_n181_1498.n80 a_0_n209# 0.0105f
C233 a_n181_1498.n81 a_0_n209# 0.0233f
C234 a_n181_1498.t70 a_0_n209# 0.0339f
C235 a_n181_1498.t65 a_0_n209# 0.0342f
C236 a_n181_1498.t86 a_0_n209# 0.0342f
C237 a_n181_1498.t61 a_0_n209# 0.0339f
C238 a_n181_1498.t77 a_0_n209# 0.0339f
C239 a_n181_1498.t78 a_0_n209# 0.0342f
C240 a_n181_1498.t62 a_0_n209# 0.0342f
C241 a_n181_1498.t76 a_0_n209# 0.0339f
C242 a_n181_1498.t60 a_0_n209# 0.0339f
C243 a_n181_1498.t83 a_0_n209# 0.0342f
C244 a_n181_1498.n82 a_0_n209# 0.0341f
C245 a_n181_1498.n83 a_0_n209# 0.0338f
C246 a_n181_1498.n84 a_0_n209# 0.0338f
C247 a_n181_1498.n85 a_0_n209# 0.0341f
C248 a_n181_1498.n86 a_0_n209# 0.0341f
C249 a_n181_1498.n87 a_0_n209# 0.0338f
C250 a_n181_1498.n88 a_0_n209# 0.0338f
C251 a_n181_1498.n89 a_0_n209# 0.0341f
C252 a_n181_1498.n90 a_0_n209# 0.0341f
C253 a_n181_1498.n91 a_0_n209# 0.0473f
C254 a_n181_1498.t36 a_0_n209# 0.0307f
C255 a_n181_1498.t18 a_0_n209# 0.0508f
C256 a_n181_1498.n92 a_0_n209# 0.0275f
C257 a_n181_1498.n93 a_0_n209# 0.0226f
C258 a_n181_1498.n94 a_0_n209# 0.0207f
C259 a_n181_1498.t32 a_0_n209# 0.0307f
C260 a_n181_1498.n95 a_0_n209# 0.0144f
C261 a_n181_1498.n96 a_0_n209# 0.0226f
C262 a_n181_1498.n97 a_0_n209# 0.0268f
C263 a_n181_1498.t52 a_0_n209# 0.0105f
C264 a_n181_1498.n98 a_0_n209# 0.0105f
C265 a_n181_1498.n99 a_0_n209# 0.0228f
C266 a_n181_1498.n100 a_0_n209# 0.0355f
C267 a_n181_1498.t7 a_0_n209# 0.0105f
C268 a_n181_1498.n101 a_0_n209# 0.0105f
C269 a_n181_1498.n102 a_0_n209# 0.0233f
C270 a_n181_1498.n103 a_0_n209# 0.0406f
C271 a_n181_1498.n104 a_0_n209# 0.0144f
C272 a_n181_1498.t6 a_0_n209# 0.0307f
C273 a_n181_1498.n105 a_0_n209# 0.0226f
C274 a_n181_1498.n106 a_0_n209# 0.0348f
C275 a_n181_1498.n107 a_0_n209# 0.0144f
C276 a_n181_1498.t2 a_0_n209# 0.0307f
C277 a_n181_1498.n108 a_0_n209# 0.0226f
C278 a_n181_1498.n109 a_0_n209# 0.0343f
C279 a_n181_1498.t57 a_0_n209# 0.0105f
C280 a_n181_1498.n110 a_0_n209# 0.0105f
C281 a_n181_1498.n111 a_0_n209# 0.023f
C282 a_n181_1498.n112 a_0_n209# 0.0412f
C283 a_n181_1498.n113 a_0_n209# 0.0358f
C284 a_n181_1498.t12 a_0_n209# 0.0307f
C285 a_n181_1498.n114 a_0_n209# 0.0144f
C286 a_n181_1498.n115 a_0_n209# 0.0226f
C287 a_n181_1498.n116 a_0_n209# 0.0273f
C288 a_n181_1498.t8 a_0_n209# 0.0307f
C289 a_n181_1498.n117 a_0_n209# 0.0144f
C290 a_n181_1498.n118 a_0_n209# 0.0226f
C291 a_n181_1498.n119 a_0_n209# 0.0276f
C292 a_n181_1498.n120 a_0_n209# 0.0359f
C293 a_n181_1498.t31 a_0_n209# 0.0105f
C294 a_n181_1498.n121 a_0_n209# 0.0105f
C295 a_n181_1498.n122 a_0_n209# 0.0233f
C296 a_n181_1498.n123 a_0_n209# 0.0406f
C297 a_n181_1498.n124 a_0_n209# 0.0144f
C298 a_n181_1498.t30 a_0_n209# 0.0307f
C299 a_n181_1498.n125 a_0_n209# 0.0226f
C300 a_n181_1498.n126 a_0_n209# 0.031f
C301 a_n181_1498.n127 a_0_n209# 0.0388f
C302 a_n181_1498.n128 a_0_n209# 0.0412f
C303 a_n181_1498.n129 a_0_n209# 0.0362f
C304 a_n181_1498.n130 a_0_n209# 0.0105f
C305 a_n181_1498.n131 a_0_n209# 0.023f
C306 a_n181_1498.t39 a_0_n209# 0.0105f
C307 a_24_587.n0 a_0_n209# 0.025f
C308 a_24_587.n1 a_0_n209# 0.0521f
C309 a_24_587.n2 a_0_n209# 0.0842f
C310 a_24_587.n3 a_0_n209# 0.0244f
C311 a_24_587.n4 a_0_n209# 0.0139f
C312 a_24_587.n5 a_0_n209# 0.0305f
C313 a_24_587.n6 a_0_n209# 0.0915f
C314 a_24_587.n7 a_0_n209# 0.0168f
C315 a_24_587.n8 a_0_n209# 0.0165f
C316 a_24_587.n9 a_0_n209# 0.0156f
C317 a_24_587.n10 a_0_n209# 0.0155f
C318 a_24_587.n11 a_0_n209# 0.0155f
C319 a_24_587.t33 a_0_n209# 0.00998f
C320 a_24_587.n12 a_0_n209# 0.00998f
C321 a_24_587.n13 a_0_n209# 0.0212f
C322 a_24_587.n14 a_0_n209# 0.0497f
C323 a_24_587.t10 a_0_n209# 0.0292f
C324 a_24_587.n15 a_0_n209# 0.0735f
C325 a_24_587.n16 a_0_n209# 0.0283f
C326 a_24_587.t32 a_0_n209# 0.0292f
C327 a_24_587.n17 a_0_n209# 0.0221f
C328 a_24_587.n18 a_0_n209# 0.0605f
C329 a_24_587.t16 a_0_n209# 0.0292f
C330 a_24_587.n19 a_0_n209# 0.0221f
C331 a_24_587.n20 a_0_n209# 0.0278f
C332 a_24_587.n21 a_0_n209# 0.0278f
C333 a_24_587.t36 a_0_n209# 0.0292f
C334 a_24_587.n22 a_0_n209# 0.0221f
C335 a_24_587.n23 a_0_n209# 0.0248f
C336 a_24_587.n24 a_0_n209# 0.00297f
C337 a_24_587.t0 a_0_n209# 0.0276f
C338 a_24_587.n25 a_0_n209# 0.0172f
C339 a_24_587.n26 a_0_n209# 0.00585f
C340 a_24_587.n27 a_0_n209# 0.035f
C341 a_24_587.t59 a_0_n209# 0.048f
C342 a_24_587.t43 a_0_n209# 0.0319f
C343 a_24_587.n28 a_0_n209# 0.0582f
C344 a_24_587.t65 a_0_n209# 0.0319f
C345 a_24_587.n29 a_0_n209# 0.0459f
C346 a_24_587.n30 a_0_n209# 0.0276f
C347 a_24_587.t47 a_0_n209# 0.0273f
C348 a_24_587.n32 a_0_n209# 0.0169f
C349 a_24_587.n33 a_0_n209# 0.00606f
C350 a_24_587.t25 a_0_n209# 0.00998f
C351 a_24_587.n34 a_0_n209# 0.00998f
C352 a_24_587.n35 a_0_n209# 0.0212f
C353 a_24_587.t24 a_0_n209# 0.0289f
C354 a_24_587.t4 a_0_n209# 0.0289f
C355 a_24_587.t23 a_0_n209# 0.00998f
C356 a_24_587.n36 a_0_n209# 0.00998f
C357 a_24_587.n37 a_0_n209# 0.0212f
C358 a_24_587.t22 a_0_n209# 0.0289f
C359 a_24_587.n38 a_0_n209# 0.0309f
C360 a_24_587.n39 a_0_n209# 0.0603f
C361 a_24_587.n40 a_0_n209# 0.0218f
C362 a_24_587.n41 a_0_n209# 0.0288f
C363 a_24_587.n42 a_0_n209# 0.0278f
C364 a_24_587.n43 a_0_n209# 0.0218f
C365 a_24_587.n44 a_0_n209# 0.0432f
C366 a_24_587.t6 a_0_n209# 0.0272f
C367 a_24_587.n45 a_0_n209# 0.0166f
C368 a_24_587.n46 a_0_n209# 0.0278f
C369 a_24_587.n47 a_0_n209# 0.00626f
C370 a_24_587.t35 a_0_n209# 0.00998f
C371 a_24_587.n48 a_0_n209# 0.00998f
C372 a_24_587.n49 a_0_n209# 0.0212f
C373 a_24_587.t34 a_0_n209# 0.0289f
C374 a_24_587.n50 a_0_n209# 0.0278f
C375 a_24_587.n51 a_0_n209# 0.0218f
C376 a_24_587.n52 a_0_n209# 0.0432f
C377 a_24_587.t18 a_0_n209# 0.0273f
C378 a_24_587.n53 a_0_n209# 0.0169f
C379 a_24_587.t26 a_0_n209# 0.0289f
C380 a_24_587.t27 a_0_n209# 0.00998f
C381 a_24_587.n54 a_0_n209# 0.00998f
C382 a_24_587.n55 a_0_n209# 0.0212f
C383 a_24_587.t8 a_0_n209# 0.0289f
C384 a_24_587.n56 a_0_n209# 0.0309f
C385 a_24_587.n57 a_0_n209# 0.0603f
C386 a_24_587.n58 a_0_n209# 0.0218f
C387 a_24_587.n59 a_0_n209# 0.0288f
C388 a_24_587.n60 a_0_n209# 0.0277f
C389 a_24_587.n61 a_0_n209# 0.00595f
C390 a_24_587.n62 a_0_n209# 0.108f
C391 a_24_587.n63 a_0_n209# 0.0278f
C392 a_24_587.t12 a_0_n209# 0.0273f
C393 a_24_587.n65 a_0_n209# 0.0167f
C394 a_24_587.n66 a_0_n209# 0.00616f
C395 a_24_587.t31 a_0_n209# 0.00998f
C396 a_24_587.n67 a_0_n209# 0.00998f
C397 a_24_587.n68 a_0_n209# 0.0212f
C398 a_24_587.t30 a_0_n209# 0.0289f
C399 a_24_587.n69 a_0_n209# 0.0278f
C400 a_24_587.n70 a_0_n209# 0.0218f
C401 a_24_587.n71 a_0_n209# 0.0441f
C402 a_24_587.n72 a_0_n209# 0.049f
C403 a_24_587.n73 a_0_n209# 0.108f
C404 a_24_587.t50 a_0_n209# 0.0285f
C405 a_24_587.t52 a_0_n209# 0.0691f
C406 a_24_587.t62 a_0_n209# 0.0322f
C407 a_24_587.n74 a_0_n209# 0.052f
C408 a_24_587.t44 a_0_n209# 0.0322f
C409 a_24_587.n75 a_0_n209# 0.0462f
C410 a_24_587.t42 a_0_n209# 0.0322f
C411 a_24_587.n76 a_0_n209# 0.0462f
C412 a_24_587.n77 a_0_n209# 0.0286f
C413 a_24_587.n78 a_0_n209# 0.0369f
C414 a_24_587.n79 a_0_n209# 0.105f
C415 a_24_587.n80 a_0_n209# 0.0792f
C416 a_24_587.t60 a_0_n209# 0.0691f
C417 a_24_587.t49 a_0_n209# 0.0322f
C418 a_24_587.n81 a_0_n209# 0.052f
C419 a_24_587.t68 a_0_n209# 0.0322f
C420 a_24_587.n82 a_0_n209# 0.0462f
C421 a_24_587.t66 a_0_n209# 0.0322f
C422 a_24_587.n83 a_0_n209# 0.0462f
C423 a_24_587.n84 a_0_n209# 0.0286f
C424 a_24_587.t48 a_0_n209# 0.0285f
C425 a_24_587.n85 a_0_n209# 0.0368f
C426 a_24_587.n86 a_0_n209# 0.105f
C427 a_24_587.n87 a_0_n209# 0.0884f
C428 a_24_587.t67 a_0_n209# 0.048f
C429 a_24_587.t57 a_0_n209# 0.0319f
C430 a_24_587.n88 a_0_n209# 0.0582f
C431 a_24_587.t45 a_0_n209# 0.0319f
C432 a_24_587.n89 a_0_n209# 0.0459f
C433 a_24_587.n90 a_0_n209# 0.0277f
C434 a_24_587.t64 a_0_n209# 0.0273f
C435 a_24_587.n92 a_0_n209# 0.0169f
C436 a_24_587.n93 a_0_n209# 0.00597f
C437 a_24_587.n94 a_0_n209# 0.0362f
C438 a_24_587.n95 a_0_n209# 0.0823f
C439 a_24_587.t54 a_0_n209# 0.0319f
C440 a_24_587.n96 a_0_n209# 0.0459f
C441 a_24_587.n97 a_0_n209# 0.0278f
C442 a_24_587.t58 a_0_n209# 0.0273f
C443 a_24_587.n99 a_0_n209# 0.0167f
C444 a_24_587.n100 a_0_n209# 0.00618f
C445 a_24_587.n101 a_0_n209# 0.0959f
C446 a_24_587.t21 a_0_n209# 0.00998f
C447 a_24_587.n102 a_0_n209# 0.00998f
C448 a_24_587.n103 a_0_n209# 0.0212f
C449 a_24_587.n104 a_0_n209# 0.0278f
C450 a_24_587.t20 a_0_n209# 0.0292f
C451 a_24_587.n105 a_0_n209# 0.0221f
C452 a_24_587.n106 a_0_n209# 0.0434f
C453 a_24_587.t29 a_0_n209# 0.00998f
C454 a_24_587.n107 a_0_n209# 0.00998f
C455 a_24_587.n108 a_0_n209# 0.0212f
C456 a_24_587.t39 a_0_n209# 0.0497f
C457 a_24_587.t38 a_0_n209# 0.0292f
C458 a_24_587.n109 a_0_n209# 0.0735f
C459 a_24_587.n110 a_0_n209# 0.0284f
C460 a_24_587.t14 a_0_n209# 0.0291f
C461 a_24_587.n111 a_0_n209# 0.0221f
C462 a_24_587.n112 a_0_n209# 0.0604f
C463 a_24_587.t28 a_0_n209# 0.0292f
C464 a_24_587.n113 a_0_n209# 0.0221f
C465 a_24_587.n114 a_0_n209# 0.0278f
C466 a_24_587.n115 a_0_n209# 0.0277f
C467 a_24_587.n116 a_0_n209# 4.21e-19
C468 a_24_587.t2 a_0_n209# 0.0261f
C469 a_24_587.n117 a_0_n209# 0.0183f
C470 a_24_587.n118 a_0_n209# 0.00595f
C471 a_24_587.n119 a_0_n209# 0.139f
C472 a_24_587.n120 a_0_n209# 0.0446f
C473 a_24_587.n121 a_0_n209# 0.00998f
C474 a_24_587.n122 a_0_n209# 0.0212f
C475 a_24_587.t37 a_0_n209# 0.00998f
.ends

