magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7578 -2284 7578 2284
<< nwell >>
rect -5578 -284 5578 284
<< nsubdiff >>
rect -5495 179 5495 201
rect -5495 133 -5428 179
rect 5428 133 5495 179
rect -5495 75 5495 133
rect -5495 29 -5428 75
rect 5428 29 5495 75
rect -5495 -29 5495 29
rect -5495 -75 -5428 -29
rect 5428 -75 5495 -29
rect -5495 -133 5495 -75
rect -5495 -179 -5428 -133
rect 5428 -179 5495 -133
rect -5495 -201 5495 -179
<< nsubdiffcont >>
rect -5428 133 5428 179
rect -5428 29 5428 75
rect -5428 -75 5428 -29
rect -5428 -179 5428 -133
<< metal1 >>
rect -5484 179 5484 190
rect -5484 133 -5428 179
rect 5428 133 5484 179
rect -5484 75 5484 133
rect -5484 29 -5428 75
rect 5428 29 5484 75
rect -5484 -29 5484 29
rect -5484 -75 -5428 -29
rect 5428 -75 5484 -29
rect -5484 -133 5484 -75
rect -5484 -179 -5428 -133
rect 5428 -179 5484 -133
rect -5484 -190 5484 -179
<< end >>
