magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2042 -2042 2042 2042
<< polysilicon >>
rect -42 23 42 42
rect -42 -23 -23 23
rect 23 -23 42 23
rect -42 -42 42 -23
<< polycontact >>
rect -23 -23 23 23
<< metal1 >>
rect -34 23 34 34
rect -34 -23 -23 23
rect 23 -23 34 23
rect -34 -34 34 -23
<< end >>
