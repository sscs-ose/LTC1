magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2139 -2045 2139 2045
<< psubdiff >>
rect -139 23 139 45
rect -139 -23 -117 23
rect 117 -23 139 23
rect -139 -45 139 -23
<< psubdiffcont >>
rect -117 -23 117 23
<< metal1 >>
rect -128 23 128 34
rect -128 -23 -117 23
rect 117 -23 128 23
rect -128 -34 128 -23
<< end >>
