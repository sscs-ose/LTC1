magic
tech gf180mcuC
magscale 1 10
timestamp 1697518002
<< nwell >>
rect -2978 -758 2978 758
<< pmos >>
rect -2804 68 -2704 628
rect -2600 68 -2500 628
rect -2396 68 -2296 628
rect -2192 68 -2092 628
rect -1988 68 -1888 628
rect -1784 68 -1684 628
rect -1580 68 -1480 628
rect -1376 68 -1276 628
rect -1172 68 -1072 628
rect -968 68 -868 628
rect -764 68 -664 628
rect -560 68 -460 628
rect -356 68 -256 628
rect -152 68 -52 628
rect 52 68 152 628
rect 256 68 356 628
rect 460 68 560 628
rect 664 68 764 628
rect 868 68 968 628
rect 1072 68 1172 628
rect 1276 68 1376 628
rect 1480 68 1580 628
rect 1684 68 1784 628
rect 1888 68 1988 628
rect 2092 68 2192 628
rect 2296 68 2396 628
rect 2500 68 2600 628
rect 2704 68 2804 628
rect -2804 -628 -2704 -68
rect -2600 -628 -2500 -68
rect -2396 -628 -2296 -68
rect -2192 -628 -2092 -68
rect -1988 -628 -1888 -68
rect -1784 -628 -1684 -68
rect -1580 -628 -1480 -68
rect -1376 -628 -1276 -68
rect -1172 -628 -1072 -68
rect -968 -628 -868 -68
rect -764 -628 -664 -68
rect -560 -628 -460 -68
rect -356 -628 -256 -68
rect -152 -628 -52 -68
rect 52 -628 152 -68
rect 256 -628 356 -68
rect 460 -628 560 -68
rect 664 -628 764 -68
rect 868 -628 968 -68
rect 1072 -628 1172 -68
rect 1276 -628 1376 -68
rect 1480 -628 1580 -68
rect 1684 -628 1784 -68
rect 1888 -628 1988 -68
rect 2092 -628 2192 -68
rect 2296 -628 2396 -68
rect 2500 -628 2600 -68
rect 2704 -628 2804 -68
<< pdiff >>
rect -2892 615 -2804 628
rect -2892 81 -2879 615
rect -2833 81 -2804 615
rect -2892 68 -2804 81
rect -2704 615 -2600 628
rect -2704 81 -2675 615
rect -2629 81 -2600 615
rect -2704 68 -2600 81
rect -2500 615 -2396 628
rect -2500 81 -2471 615
rect -2425 81 -2396 615
rect -2500 68 -2396 81
rect -2296 615 -2192 628
rect -2296 81 -2267 615
rect -2221 81 -2192 615
rect -2296 68 -2192 81
rect -2092 615 -1988 628
rect -2092 81 -2063 615
rect -2017 81 -1988 615
rect -2092 68 -1988 81
rect -1888 615 -1784 628
rect -1888 81 -1859 615
rect -1813 81 -1784 615
rect -1888 68 -1784 81
rect -1684 615 -1580 628
rect -1684 81 -1655 615
rect -1609 81 -1580 615
rect -1684 68 -1580 81
rect -1480 615 -1376 628
rect -1480 81 -1451 615
rect -1405 81 -1376 615
rect -1480 68 -1376 81
rect -1276 615 -1172 628
rect -1276 81 -1247 615
rect -1201 81 -1172 615
rect -1276 68 -1172 81
rect -1072 615 -968 628
rect -1072 81 -1043 615
rect -997 81 -968 615
rect -1072 68 -968 81
rect -868 615 -764 628
rect -868 81 -839 615
rect -793 81 -764 615
rect -868 68 -764 81
rect -664 615 -560 628
rect -664 81 -635 615
rect -589 81 -560 615
rect -664 68 -560 81
rect -460 615 -356 628
rect -460 81 -431 615
rect -385 81 -356 615
rect -460 68 -356 81
rect -256 615 -152 628
rect -256 81 -227 615
rect -181 81 -152 615
rect -256 68 -152 81
rect -52 615 52 628
rect -52 81 -23 615
rect 23 81 52 615
rect -52 68 52 81
rect 152 615 256 628
rect 152 81 181 615
rect 227 81 256 615
rect 152 68 256 81
rect 356 615 460 628
rect 356 81 385 615
rect 431 81 460 615
rect 356 68 460 81
rect 560 615 664 628
rect 560 81 589 615
rect 635 81 664 615
rect 560 68 664 81
rect 764 615 868 628
rect 764 81 793 615
rect 839 81 868 615
rect 764 68 868 81
rect 968 615 1072 628
rect 968 81 997 615
rect 1043 81 1072 615
rect 968 68 1072 81
rect 1172 615 1276 628
rect 1172 81 1201 615
rect 1247 81 1276 615
rect 1172 68 1276 81
rect 1376 615 1480 628
rect 1376 81 1405 615
rect 1451 81 1480 615
rect 1376 68 1480 81
rect 1580 615 1684 628
rect 1580 81 1609 615
rect 1655 81 1684 615
rect 1580 68 1684 81
rect 1784 615 1888 628
rect 1784 81 1813 615
rect 1859 81 1888 615
rect 1784 68 1888 81
rect 1988 615 2092 628
rect 1988 81 2017 615
rect 2063 81 2092 615
rect 1988 68 2092 81
rect 2192 615 2296 628
rect 2192 81 2221 615
rect 2267 81 2296 615
rect 2192 68 2296 81
rect 2396 615 2500 628
rect 2396 81 2425 615
rect 2471 81 2500 615
rect 2396 68 2500 81
rect 2600 615 2704 628
rect 2600 81 2629 615
rect 2675 81 2704 615
rect 2600 68 2704 81
rect 2804 615 2892 628
rect 2804 81 2833 615
rect 2879 81 2892 615
rect 2804 68 2892 81
rect -2892 -81 -2804 -68
rect -2892 -615 -2879 -81
rect -2833 -615 -2804 -81
rect -2892 -628 -2804 -615
rect -2704 -81 -2600 -68
rect -2704 -615 -2675 -81
rect -2629 -615 -2600 -81
rect -2704 -628 -2600 -615
rect -2500 -81 -2396 -68
rect -2500 -615 -2471 -81
rect -2425 -615 -2396 -81
rect -2500 -628 -2396 -615
rect -2296 -81 -2192 -68
rect -2296 -615 -2267 -81
rect -2221 -615 -2192 -81
rect -2296 -628 -2192 -615
rect -2092 -81 -1988 -68
rect -2092 -615 -2063 -81
rect -2017 -615 -1988 -81
rect -2092 -628 -1988 -615
rect -1888 -81 -1784 -68
rect -1888 -615 -1859 -81
rect -1813 -615 -1784 -81
rect -1888 -628 -1784 -615
rect -1684 -81 -1580 -68
rect -1684 -615 -1655 -81
rect -1609 -615 -1580 -81
rect -1684 -628 -1580 -615
rect -1480 -81 -1376 -68
rect -1480 -615 -1451 -81
rect -1405 -615 -1376 -81
rect -1480 -628 -1376 -615
rect -1276 -81 -1172 -68
rect -1276 -615 -1247 -81
rect -1201 -615 -1172 -81
rect -1276 -628 -1172 -615
rect -1072 -81 -968 -68
rect -1072 -615 -1043 -81
rect -997 -615 -968 -81
rect -1072 -628 -968 -615
rect -868 -81 -764 -68
rect -868 -615 -839 -81
rect -793 -615 -764 -81
rect -868 -628 -764 -615
rect -664 -81 -560 -68
rect -664 -615 -635 -81
rect -589 -615 -560 -81
rect -664 -628 -560 -615
rect -460 -81 -356 -68
rect -460 -615 -431 -81
rect -385 -615 -356 -81
rect -460 -628 -356 -615
rect -256 -81 -152 -68
rect -256 -615 -227 -81
rect -181 -615 -152 -81
rect -256 -628 -152 -615
rect -52 -81 52 -68
rect -52 -615 -23 -81
rect 23 -615 52 -81
rect -52 -628 52 -615
rect 152 -81 256 -68
rect 152 -615 181 -81
rect 227 -615 256 -81
rect 152 -628 256 -615
rect 356 -81 460 -68
rect 356 -615 385 -81
rect 431 -615 460 -81
rect 356 -628 460 -615
rect 560 -81 664 -68
rect 560 -615 589 -81
rect 635 -615 664 -81
rect 560 -628 664 -615
rect 764 -81 868 -68
rect 764 -615 793 -81
rect 839 -615 868 -81
rect 764 -628 868 -615
rect 968 -81 1072 -68
rect 968 -615 997 -81
rect 1043 -615 1072 -81
rect 968 -628 1072 -615
rect 1172 -81 1276 -68
rect 1172 -615 1201 -81
rect 1247 -615 1276 -81
rect 1172 -628 1276 -615
rect 1376 -81 1480 -68
rect 1376 -615 1405 -81
rect 1451 -615 1480 -81
rect 1376 -628 1480 -615
rect 1580 -81 1684 -68
rect 1580 -615 1609 -81
rect 1655 -615 1684 -81
rect 1580 -628 1684 -615
rect 1784 -81 1888 -68
rect 1784 -615 1813 -81
rect 1859 -615 1888 -81
rect 1784 -628 1888 -615
rect 1988 -81 2092 -68
rect 1988 -615 2017 -81
rect 2063 -615 2092 -81
rect 1988 -628 2092 -615
rect 2192 -81 2296 -68
rect 2192 -615 2221 -81
rect 2267 -615 2296 -81
rect 2192 -628 2296 -615
rect 2396 -81 2500 -68
rect 2396 -615 2425 -81
rect 2471 -615 2500 -81
rect 2396 -628 2500 -615
rect 2600 -81 2704 -68
rect 2600 -615 2629 -81
rect 2675 -615 2704 -81
rect 2600 -628 2704 -615
rect 2804 -81 2892 -68
rect 2804 -615 2833 -81
rect 2879 -615 2892 -81
rect 2804 -628 2892 -615
<< pdiffc >>
rect -2879 81 -2833 615
rect -2675 81 -2629 615
rect -2471 81 -2425 615
rect -2267 81 -2221 615
rect -2063 81 -2017 615
rect -1859 81 -1813 615
rect -1655 81 -1609 615
rect -1451 81 -1405 615
rect -1247 81 -1201 615
rect -1043 81 -997 615
rect -839 81 -793 615
rect -635 81 -589 615
rect -431 81 -385 615
rect -227 81 -181 615
rect -23 81 23 615
rect 181 81 227 615
rect 385 81 431 615
rect 589 81 635 615
rect 793 81 839 615
rect 997 81 1043 615
rect 1201 81 1247 615
rect 1405 81 1451 615
rect 1609 81 1655 615
rect 1813 81 1859 615
rect 2017 81 2063 615
rect 2221 81 2267 615
rect 2425 81 2471 615
rect 2629 81 2675 615
rect 2833 81 2879 615
rect -2879 -615 -2833 -81
rect -2675 -615 -2629 -81
rect -2471 -615 -2425 -81
rect -2267 -615 -2221 -81
rect -2063 -615 -2017 -81
rect -1859 -615 -1813 -81
rect -1655 -615 -1609 -81
rect -1451 -615 -1405 -81
rect -1247 -615 -1201 -81
rect -1043 -615 -997 -81
rect -839 -615 -793 -81
rect -635 -615 -589 -81
rect -431 -615 -385 -81
rect -227 -615 -181 -81
rect -23 -615 23 -81
rect 181 -615 227 -81
rect 385 -615 431 -81
rect 589 -615 635 -81
rect 793 -615 839 -81
rect 997 -615 1043 -81
rect 1201 -615 1247 -81
rect 1405 -615 1451 -81
rect 1609 -615 1655 -81
rect 1813 -615 1859 -81
rect 2017 -615 2063 -81
rect 2221 -615 2267 -81
rect 2425 -615 2471 -81
rect 2629 -615 2675 -81
rect 2833 -615 2879 -81
<< polysilicon >>
rect -2804 628 -2704 672
rect -2600 628 -2500 672
rect -2396 628 -2296 672
rect -2192 628 -2092 672
rect -1988 628 -1888 672
rect -1784 628 -1684 672
rect -1580 628 -1480 672
rect -1376 628 -1276 672
rect -1172 628 -1072 672
rect -968 628 -868 672
rect -764 628 -664 672
rect -560 628 -460 672
rect -356 628 -256 672
rect -152 628 -52 672
rect 52 628 152 672
rect 256 628 356 672
rect 460 628 560 672
rect 664 628 764 672
rect 868 628 968 672
rect 1072 628 1172 672
rect 1276 628 1376 672
rect 1480 628 1580 672
rect 1684 628 1784 672
rect 1888 628 1988 672
rect 2092 628 2192 672
rect 2296 628 2396 672
rect 2500 628 2600 672
rect 2704 628 2804 672
rect -2804 24 -2704 68
rect -2600 24 -2500 68
rect -2396 24 -2296 68
rect -2192 24 -2092 68
rect -1988 24 -1888 68
rect -1784 24 -1684 68
rect -1580 24 -1480 68
rect -1376 24 -1276 68
rect -1172 24 -1072 68
rect -968 24 -868 68
rect -764 24 -664 68
rect -560 24 -460 68
rect -356 24 -256 68
rect -152 24 -52 68
rect 52 24 152 68
rect 256 24 356 68
rect 460 24 560 68
rect 664 24 764 68
rect 868 24 968 68
rect 1072 24 1172 68
rect 1276 24 1376 68
rect 1480 24 1580 68
rect 1684 24 1784 68
rect 1888 24 1988 68
rect 2092 24 2192 68
rect 2296 24 2396 68
rect 2500 24 2600 68
rect 2704 24 2804 68
rect -2804 -68 -2704 -24
rect -2600 -68 -2500 -24
rect -2396 -68 -2296 -24
rect -2192 -68 -2092 -24
rect -1988 -68 -1888 -24
rect -1784 -68 -1684 -24
rect -1580 -68 -1480 -24
rect -1376 -68 -1276 -24
rect -1172 -68 -1072 -24
rect -968 -68 -868 -24
rect -764 -68 -664 -24
rect -560 -68 -460 -24
rect -356 -68 -256 -24
rect -152 -68 -52 -24
rect 52 -68 152 -24
rect 256 -68 356 -24
rect 460 -68 560 -24
rect 664 -68 764 -24
rect 868 -68 968 -24
rect 1072 -68 1172 -24
rect 1276 -68 1376 -24
rect 1480 -68 1580 -24
rect 1684 -68 1784 -24
rect 1888 -68 1988 -24
rect 2092 -68 2192 -24
rect 2296 -68 2396 -24
rect 2500 -68 2600 -24
rect 2704 -68 2804 -24
rect -2804 -672 -2704 -628
rect -2600 -672 -2500 -628
rect -2396 -672 -2296 -628
rect -2192 -672 -2092 -628
rect -1988 -672 -1888 -628
rect -1784 -672 -1684 -628
rect -1580 -672 -1480 -628
rect -1376 -672 -1276 -628
rect -1172 -672 -1072 -628
rect -968 -672 -868 -628
rect -764 -672 -664 -628
rect -560 -672 -460 -628
rect -356 -672 -256 -628
rect -152 -672 -52 -628
rect 52 -672 152 -628
rect 256 -672 356 -628
rect 460 -672 560 -628
rect 664 -672 764 -628
rect 868 -672 968 -628
rect 1072 -672 1172 -628
rect 1276 -672 1376 -628
rect 1480 -672 1580 -628
rect 1684 -672 1784 -628
rect 1888 -672 1988 -628
rect 2092 -672 2192 -628
rect 2296 -672 2396 -628
rect 2500 -672 2600 -628
rect 2704 -672 2804 -628
<< metal1 >>
rect -2879 615 -2833 626
rect -2879 70 -2833 81
rect -2675 615 -2629 626
rect -2675 70 -2629 81
rect -2471 615 -2425 626
rect -2471 70 -2425 81
rect -2267 615 -2221 626
rect -2267 70 -2221 81
rect -2063 615 -2017 626
rect -2063 70 -2017 81
rect -1859 615 -1813 626
rect -1859 70 -1813 81
rect -1655 615 -1609 626
rect -1655 70 -1609 81
rect -1451 615 -1405 626
rect -1451 70 -1405 81
rect -1247 615 -1201 626
rect -1247 70 -1201 81
rect -1043 615 -997 626
rect -1043 70 -997 81
rect -839 615 -793 626
rect -839 70 -793 81
rect -635 615 -589 626
rect -635 70 -589 81
rect -431 615 -385 626
rect -431 70 -385 81
rect -227 615 -181 626
rect -227 70 -181 81
rect -23 615 23 626
rect -23 70 23 81
rect 181 615 227 626
rect 181 70 227 81
rect 385 615 431 626
rect 385 70 431 81
rect 589 615 635 626
rect 589 70 635 81
rect 793 615 839 626
rect 793 70 839 81
rect 997 615 1043 626
rect 997 70 1043 81
rect 1201 615 1247 626
rect 1201 70 1247 81
rect 1405 615 1451 626
rect 1405 70 1451 81
rect 1609 615 1655 626
rect 1609 70 1655 81
rect 1813 615 1859 626
rect 1813 70 1859 81
rect 2017 615 2063 626
rect 2017 70 2063 81
rect 2221 615 2267 626
rect 2221 70 2267 81
rect 2425 615 2471 626
rect 2425 70 2471 81
rect 2629 615 2675 626
rect 2629 70 2675 81
rect 2833 615 2879 626
rect 2833 70 2879 81
rect -2879 -81 -2833 -70
rect -2879 -626 -2833 -615
rect -2675 -81 -2629 -70
rect -2675 -626 -2629 -615
rect -2471 -81 -2425 -70
rect -2471 -626 -2425 -615
rect -2267 -81 -2221 -70
rect -2267 -626 -2221 -615
rect -2063 -81 -2017 -70
rect -2063 -626 -2017 -615
rect -1859 -81 -1813 -70
rect -1859 -626 -1813 -615
rect -1655 -81 -1609 -70
rect -1655 -626 -1609 -615
rect -1451 -81 -1405 -70
rect -1451 -626 -1405 -615
rect -1247 -81 -1201 -70
rect -1247 -626 -1201 -615
rect -1043 -81 -997 -70
rect -1043 -626 -997 -615
rect -839 -81 -793 -70
rect -839 -626 -793 -615
rect -635 -81 -589 -70
rect -635 -626 -589 -615
rect -431 -81 -385 -70
rect -431 -626 -385 -615
rect -227 -81 -181 -70
rect -227 -626 -181 -615
rect -23 -81 23 -70
rect -23 -626 23 -615
rect 181 -81 227 -70
rect 181 -626 227 -615
rect 385 -81 431 -70
rect 385 -626 431 -615
rect 589 -81 635 -70
rect 589 -626 635 -615
rect 793 -81 839 -70
rect 793 -626 839 -615
rect 997 -81 1043 -70
rect 997 -626 1043 -615
rect 1201 -81 1247 -70
rect 1201 -626 1247 -615
rect 1405 -81 1451 -70
rect 1405 -626 1451 -615
rect 1609 -81 1655 -70
rect 1609 -626 1655 -615
rect 1813 -81 1859 -70
rect 1813 -626 1859 -615
rect 2017 -81 2063 -70
rect 2017 -626 2063 -615
rect 2221 -81 2267 -70
rect 2221 -626 2267 -615
rect 2425 -81 2471 -70
rect 2425 -626 2471 -615
rect 2629 -81 2675 -70
rect 2629 -626 2675 -615
rect 2833 -81 2879 -70
rect 2833 -626 2879 -615
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2.8 l 0.5 m 2 nf 28 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
