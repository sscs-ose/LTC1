magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6123 -2128 6123 2128
<< nwell >>
rect -4123 -128 4123 128
<< nsubdiff >>
rect -4040 23 4040 45
rect -4040 -23 -4018 23
rect 4018 -23 4040 23
rect -4040 -45 4040 -23
<< nsubdiffcont >>
rect -4018 -23 4018 23
<< metal1 >>
rect -4029 23 4029 34
rect -4029 -23 -4018 23
rect 4018 -23 4029 23
rect -4029 -34 4029 -23
<< end >>
