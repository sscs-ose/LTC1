magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2231 -2045 2231 2045
<< psubdiff >>
rect -231 23 231 45
rect -231 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 231 23
rect -231 -45 231 -23
<< psubdiffcont >>
rect -209 -23 -163 23
rect -85 -23 -39 23
rect 39 -23 85 23
rect 163 -23 209 23
<< metal1 >>
rect -220 23 220 34
rect -220 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 220 23
rect -220 -34 220 -23
<< end >>
