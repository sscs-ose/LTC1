magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2530 -2298 2530 2298
<< nwell >>
rect -530 -298 530 298
<< pmos >>
rect -356 68 -256 168
rect -152 68 -52 168
rect 52 68 152 168
rect 256 68 356 168
rect -356 -168 -256 -68
rect -152 -168 -52 -68
rect 52 -168 152 -68
rect 256 -168 356 -68
<< pdiff >>
rect -444 141 -356 168
rect -444 95 -431 141
rect -385 95 -356 141
rect -444 68 -356 95
rect -256 141 -152 168
rect -256 95 -227 141
rect -181 95 -152 141
rect -256 68 -152 95
rect -52 141 52 168
rect -52 95 -23 141
rect 23 95 52 141
rect -52 68 52 95
rect 152 141 256 168
rect 152 95 181 141
rect 227 95 256 141
rect 152 68 256 95
rect 356 141 444 168
rect 356 95 385 141
rect 431 95 444 141
rect 356 68 444 95
rect -444 -95 -356 -68
rect -444 -141 -431 -95
rect -385 -141 -356 -95
rect -444 -168 -356 -141
rect -256 -95 -152 -68
rect -256 -141 -227 -95
rect -181 -141 -152 -95
rect -256 -168 -152 -141
rect -52 -95 52 -68
rect -52 -141 -23 -95
rect 23 -141 52 -95
rect -52 -168 52 -141
rect 152 -95 256 -68
rect 152 -141 181 -95
rect 227 -141 256 -95
rect 152 -168 256 -141
rect 356 -95 444 -68
rect 356 -141 385 -95
rect 431 -141 444 -95
rect 356 -168 444 -141
<< pdiffc >>
rect -431 95 -385 141
rect -227 95 -181 141
rect -23 95 23 141
rect 181 95 227 141
rect 385 95 431 141
rect -431 -141 -385 -95
rect -227 -141 -181 -95
rect -23 -141 23 -95
rect 181 -141 227 -95
rect 385 -141 431 -95
<< polysilicon >>
rect -356 168 -256 212
rect -152 168 -52 212
rect 52 168 152 212
rect 256 168 356 212
rect -356 24 -256 68
rect -152 24 -52 68
rect 52 24 152 68
rect 256 24 356 68
rect -356 -68 -256 -24
rect -152 -68 -52 -24
rect 52 -68 152 -24
rect 256 -68 356 -24
rect -356 -212 -256 -168
rect -152 -212 -52 -168
rect 52 -212 152 -168
rect 256 -212 356 -168
<< metal1 >>
rect -431 141 -385 166
rect -431 70 -385 95
rect -227 141 -181 166
rect -227 70 -181 95
rect -23 141 23 166
rect -23 70 23 95
rect 181 141 227 166
rect 181 70 227 95
rect 385 141 431 166
rect 385 70 431 95
rect -431 -95 -385 -70
rect -431 -166 -385 -141
rect -227 -95 -181 -70
rect -227 -166 -181 -141
rect -23 -95 23 -70
rect -23 -166 23 -141
rect 181 -95 227 -70
rect 181 -166 227 -141
rect 385 -95 431 -70
rect 385 -166 431 -141
<< end >>
