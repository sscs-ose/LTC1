* NGSPICE file created from CM_LSB_mod_flat.ext - technology: gf180mcuC

.subckt pex_CM_LSB_mod ITAIL VSS OUT_1 OUT_2 VDD OUT_3 OUT_4 OUT_5 OUT_6
X0 OUT_6 ITAIL_1.t24 SD3_1.t42 VSS.t107 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 G2_1 ITAIL.t0 ITAIL.t1 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X2 VDD G1_1.t10 G1_1.t11 VDD.t37 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 OUT_6 ITAIL_1.t25 SD3_1.t41 VSS.t106 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X4 VSS G2_1.t3 SD2_4.t7 VSS.t141 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X5 OUT_4 ITAIL.t2 SD2_5.t3 VSS.t195 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 ITAIL_1 ITAIL_1.t19 SD0_2.t7 VSS.t37 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 SD0_2 SD0_2.t22 VSS.t164 VSS.t103 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X8 SD3_1 SD0_2.t25 VSS.t165 VSS.t86 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 SD3_1 ITAIL_1.t27 OUT_6.t29 VSS.t105 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 SD2_5 G2_1.t4 VSS.t175 VSS.t174 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 VSS G2_1.t5 SD2_5.t14 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X12 OUT_5 ITAIL_1.t28 SD0_1.t7 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X13 SD2_1 G2_1.t6 VSS.t148 VSS.t147 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X14 OUT_4 ITAIL.t3 SD2_5.t2 VSS.t195 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 SD0_1 SD0_2.t26 VSS.t149 VSS.t70 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X16 G1_1 G1_1.t14 VDD.t36 VDD.t35 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 VSS G2_1.t7 SD2_2.t1 VSS.t25 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X18 VSS SD0_2.t27 SD0_1.t30 VSS.t100 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X19 SD0_2 ITAIL_1.t15 ITAIL_1.t16 VSS.t104 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X20 VDD G1_1.t8 G1_1.t9 VDD.t32 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X21 SD0_2 ITAIL_1.t13 ITAIL_1.t14 VSS.t103 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X22 SD0_1 ITAIL_1.t29 OUT_5.t14 VSS.t102 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X23 OUT_6 ITAIL_1.t30 SD3_1.t40 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X24 VSS SD0_2.t28 SD3_1.t52 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X25 VSS SD0_2.t29 SD0_1.t29 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 SD2_5 G2_1.t8 VSS.t192 VSS.t174 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X27 ITAIL_1 ITAIL_1.t17 SD0_2.t4 VSS.t101 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X28 OUT_6 ITAIL_1.t32 SD3_1.t39 VSS.t60 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 SD3_1 ITAIL_1.t33 OUT_6.t26 VSS.t56 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X30 OUT_5 ITAIL_1.t34 SD0_1.t6 VSS.t100 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 SD0_2 SD0_2.t20 VSS.t168 VSS.t104 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X32 SD2_1 G2_1.t9 VSS.t157 VSS.t147 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X33 VSS SD0_2.t31 SD3_1.t7 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X34 VSS SD0_2.t32 SD3_1.t46 VSS.t79 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X35 SD3_1 SD0_2.t33 VSS.t126 VSS.t80 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X36 SD3_1 ITAIL_1.t35 OUT_6.t25 VSS.t58 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X37 SD2_2 ITAIL.t4 OUT_1.t0 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X38 SD0_1 SD0_2.t34 VSS.t127 VSS.t102 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X39 OUT_3 ITAIL.t5 SD2_4.t3 VSS.t52 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X40 SD3_1 SD0_2.t35 VSS.t1 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X41 G1_1 G1_1.t12 VDD.t31 VDD.t30 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X42 OUT_5 ITAIL_1.t36 SD0_1.t5 VSS.t99 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X43 VSS SD0_2.t36 SD3_1.t1 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X44 SD3_1 SD0_2.t37 VSS.t110 VSS.t78 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X45 VSS SD0_2.t18 SD0_2.t19 VSS.t101 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X46 VSS G2_1.t10 SD2_5.t12 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X47 SD3_1 ITAIL_1.t37 OUT_6.t24 VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X48 OUT_6 ITAIL_1.t38 SD3_1.t38 VSS.t98 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X49 G1_2 ITAIL.t6 SD2_1.t7 VSS.t115 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X50 SD2_1 ITAIL.t7 G1_2.t6 VSS.t144 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X51 VSS SD0_2.t38 SD0_1.t27 VSS.t97 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X52 VSS G2_1.t11 SD2_5.t11 VSS.t17 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X53 G1_2 G1_2.t22 G1_1.t21 VDD.t50 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X54 SD0_1 SD0_2.t39 VSS.t138 VSS.t95 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X55 OUT_2 ITAIL.t8 SD2_3.t0 VSS.t48 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X56 VSS SD0_2.t40 SD0_1.t25 VSS.t99 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X57 VSS G2_1.t12 SD2_1.t13 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X58 SD1_1 G1_1.t26 VDD.t29 VDD.t28 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X59 SD2_4 ITAIL.t9 OUT_3.t2 VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X60 SD2_5 G2_1.t13 VSS.t119 VSS.t15 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X61 ITAIL_1 G1_2.t25 SD1_1.t15 VDD.t51 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X62 VSS SD0_2.t41 SD3_1.t2 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X63 OUT_5 ITAIL_1.t39 SD0_1.t4 VSS.t97 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X64 VSS SD0_2.t16 SD0_2.t17 VSS.t87 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X65 SD3_1 SD0_2.t42 VSS.t14 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X66 SD3_1 ITAIL_1.t40 OUT_6.t22 VSS.t96 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X67 SD0_1 ITAIL_1.t41 OUT_5.t10 VSS.t95 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X68 OUT_5 ITAIL_1.t42 SD0_1.t3 VSS.t94 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X69 VSS G2_1.t14 SD2_4.t6 VSS.t141 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X70 SD3_1 ITAIL_1.t43 OUT_6.t21 VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X71 SD3_1 SD0_2.t43 VSS.t31 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X72 G1_1 G1_2.t20 G1_2.t21 VDD.t49 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X73 VDD G1_1.t6 G1_1.t7 VDD.t25 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X74 VSS SD0_2.t44 SD3_1.t6 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X75 VSS SD0_2.t45 SD3_1.t61 VSS.t75 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X76 SD0_2 SD0_2.t14 VSS.t191 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X77 OUT_6 ITAIL_1.t44 SD3_1.t37 VSS.t92 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X78 VDD G1_1.t27 SD1_1.t6 VDD.t22 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X79 OUT_6 ITAIL_1.t45 SD3_1.t36 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X80 SD3_1 ITAIL_1.t46 OUT_6.t18 VSS.t90 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X81 SD2_1 ITAIL.t10 G1_2.t5 VSS.t144 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X82 ITAIL_1 G1_2.t26 SD1_1.t14 VDD.t52 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X83 OUT_6 ITAIL_1.t47 SD3_1.t35 VSS.t89 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X84 SD2_1 ITAIL.t11 G1_2.t4 VSS.t145 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X85 SD3_1 ITAIL_1.t48 OUT_6.t16 VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X86 SD3_1 ITAIL_1.t49 OUT_6.t15 VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X87 SD3_1 SD0_2.t47 VSS.t158 VSS.t73 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X88 SD0_1 SD0_2.t48 VSS.t159 VSS.t82 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X89 VSS SD0_2.t49 SD3_1.t54 VSS.t72 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X90 SD2_4 G2_1.t15 VSS.t114 VSS.t113 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X91 ITAIL_1 ITAIL_1.t7 SD0_2.t3 VSS.t87 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X92 VSS G2_1.t16 SD2_1.t12 VSS.t20 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X93 SD2_4 G2_1.t17 VSS.t178 VSS.t113 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X94 SD1_1 G1_1.t28 VDD.t21 VDD.t20 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X95 VSS SD0_2.t50 SD0_1.t23 VSS.t94 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X96 SD1_1 G1_1.t29 VDD.t19 VDD.t18 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X97 SD3_1 ITAIL_1.t51 OUT_6.t14 VSS.t86 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X98 SD3_1 SD0_2.t51 VSS.t186 VSS.t105 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X99 SD0_2 ITAIL_1.t11 ITAIL_1.t12 VSS.t85 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X100 VSS SD0_2.t52 SD3_1.t48 VSS.t107 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X101 VSS SD0_2.t53 SD3_1.t49 VSS.t106 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X102 G1_1 G1_2.t18 G1_2.t19 VDD.t55 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X103 G1_2 G1_2.t16 G1_1.t22 VDD.t54 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X104 ITAIL_1 ITAIL_1.t5 SD0_2.t1 VSS.t84 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X105 VSS G2_1.t18 SD2_3.t3 VSS.t48 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X106 SD1_1 G1_2.t28 ITAIL_1.t23 VDD.t53 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X107 SD0_1 ITAIL_1.t53 OUT_5.t8 VSS.t83 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X108 SD0_1 ITAIL_1.t54 OUT_5.t7 VSS.t82 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X109 SD1_1 G1_2.t29 ITAIL_1.t0 VDD.t42 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X110 VDD G1_1.t30 SD1_1.t3 VDD.t9 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X111 SD2_5 G2_1.t19 VSS.t16 VSS.t15 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X112 ITAIL_1 G1_2.t30 SD1_1.t11 VDD.t43 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X113 SD2_5 ITAIL.t12 OUT_4.t5 VSS.t108 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X114 SD2_3 G2_1.t20 VSS.t9 VSS.t8 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X115 SD1_1 G1_1.t31 VDD.t16 VDD.t15 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X116 VDD G1_1.t4 G1_1.t5 VDD.t12 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X117 OUT_6 ITAIL_1.t55 SD3_1.t34 VSS.t81 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X118 VSS SD0_2.t12 SD0_2.t13 VSS.t84 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X119 OUT_5 ITAIL_1.t56 SD0_1.t2 VSS.t63 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X120 SD0_1 SD0_2.t54 VSS.t154 VSS.t83 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X121 VDD G1_1.t32 SD1_1.t1 VDD.t7 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X122 VSS SD0_2.t55 SD0_1.t21 VSS.t77 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X123 G1_1 G1_1.t2 VDD.t3 VDD.t2 pfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X124 VSS SD0_2.t56 SD3_1.t8 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X125 SD0_2 ITAIL_1.t9 ITAIL_1.t10 VSS.t40 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X126 SD2_1 G2_1.t21 VSS.t137 VSS.t136 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X127 SD1_1 G1_2.t31 ITAIL_1.t2 VDD.t44 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X128 SD3_1 SD0_2.t57 VSS.t57 VSS.t56 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X129 G1_1 G1_2.t14 G1_2.t15 VDD.t41 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X130 SD3_1 ITAIL_1.t57 OUT_6.t12 VSS.t80 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X131 SD1_1 G1_2.t32 ITAIL_1.t3 VDD.t47 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X132 SD3_1 SD0_2.t58 VSS.t59 VSS.t58 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X133 G1_1 G1_1.t0 VDD.t6 VDD.t5 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X134 VSS SD0_2.t59 SD3_1.t11 VSS.t60 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X135 VSS G2_1.t22 SD2_5.t8 VSS.t5 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X136 G1_2 ITAIL.t13 SD2_1.t6 VSS.t109 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X137 G1_2 ITAIL.t14 SD2_1.t5 VSS.t109 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X138 OUT_6 ITAIL_1.t58 SD3_1.t33 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X139 OUT_6 ITAIL_1.t59 SD3_1.t32 VSS.t79 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X140 VSS SD0_2.t60 SD0_1.t20 VSS.t63 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X141 SD3_1 ITAIL_1.t60 OUT_6.t9 VSS.t78 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X142 OUT_5 ITAIL_1.t61 SD0_1.t1 VSS.t77 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X143 SD2_1 ITAIL.t15 G1_2.t1 VSS.t145 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X144 SD3_1 ITAIL_1.t62 OUT_6.t8 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X145 SD0_1 SD0_2.t61 VSS.t67 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X146 SD3_1 SD0_2.t62 VSS.t69 VSS.t68 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X147 VSS G2_1.t1 G2_1.t2 VSS.t25 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X148 OUT_4 ITAIL.t16 SD2_5.t1 VSS.t128 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X149 OUT_6 ITAIL_1.t63 SD3_1.t31 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X150 SD0_2 SD0_2.t10 VSS.t41 VSS.t40 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X151 VSS SD0_2.t64 SD3_1.t62 VSS.t98 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X152 SD2_3 ITAIL.t17 OUT_2.t0 VSS.t8 nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
X153 ITAIL_1 G1_2.t33 SD1_1.t8 VDD.t48 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X154 G1_2 ITAIL.t18 SD2_1.t4 VSS.t115 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X155 SD2_5 ITAIL.t19 OUT_4.t3 VSS.t36 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X156 SD2_5 ITAIL.t20 OUT_4.t2 VSS.t108 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X157 VDD G1_1.t35 SD1_1.t0 VDD.t0 pfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X158 G1_2 G1_2.t12 G1_1.t16 VDD.t40 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X159 VSS SD0_2.t65 SD0_1.t18 VSS.t74 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X160 SD0_1 ITAIL_1.t64 OUT_5.t4 VSS.t66 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X161 SD0_1 ITAIL_1.t65 OUT_5.t3 VSS.t76 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X162 SD3_1 SD0_2.t66 VSS.t200 VSS.t96 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X163 OUT_4 ITAIL.t21 SD2_5.t0 VSS.t128 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X164 G1_1 G1_2.t10 G1_2.t11 VDD.t46 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X165 SD3_1 ITAIL_1.t66 OUT_6.t6 VSS.t30 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X166 SD0_1 SD0_2.t67 VSS.t171 VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X167 SD2_4 ITAIL.t22 OUT_3.t1 VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X168 OUT_6 ITAIL_1.t67 SD3_1.t30 VSS.t10 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X169 OUT_6 ITAIL_1.t68 SD3_1.t29 VSS.t75 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X170 OUT_5 ITAIL_1.t69 SD0_1.t0 VSS.t74 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X171 VSS SD0_2.t68 SD3_1.t56 VSS.t92 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X172 SD3_1 ITAIL_1.t70 OUT_6.t3 VSS.t13 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X173 SD2_5 ITAIL.t23 OUT_4.t0 VSS.t36 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X174 SD3_1 SD0_2.t69 VSS.t179 VSS.t88 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X175 VSS SD0_2.t70 SD3_1.t58 VSS.t89 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X176 SD3_1 SD0_2.t71 VSS.t187 VSS.t93 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X177 VSS SD0_2.t8 SD0_2.t9 VSS.t37 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X178 SD3_1 ITAIL_1.t71 OUT_6.t2 VSS.t73 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X179 OUT_6 ITAIL_1.t72 SD3_1.t28 VSS.t32 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X180 VSS G2_1.t23 SD2_1.t10 VSS.t116 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X181 OUT_6 ITAIL_1.t73 SD3_1.t27 VSS.t72 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X182 SD0_1 SD0_2.t72 VSS.t188 VSS.t76 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X183 OUT_3 ITAIL.t24 SD2_4.t2 VSS.t52 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X184 VSS G2_1.t24 SD2_1.t9 VSS.t116 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X185 VSS SD0_2.t73 SD3_1.t50 VSS.t91 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X186 SD3_1 SD0_2.t74 VSS.t135 VSS.t90 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X187 G1_2 G1_2.t8 G1_1.t18 VDD.t45 pfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X188 SD3_1 SD0_2.t75 VSS.t29 VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X189 SD2_1 G2_1.t25 VSS.t146 VSS.t136 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X190 SD0_1 ITAIL_1.t74 OUT_5.t1 VSS.t71 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X191 SD0_1 ITAIL_1.t75 OUT_5.t0 VSS.t70 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
R0 ITAIL_1.n86 ITAIL_1.n85 132.385
R1 ITAIL_1.n80 ITAIL_1.n79 131.189
R2 ITAIL_1.n2 ITAIL_1.t25 117.838
R3 ITAIL_1.n59 ITAIL_1.n58 108.54
R4 ITAIL_1.n64 ITAIL_1.n63 106.138
R5 ITAIL_1.n53 ITAIL_1.n52 105.632
R6 ITAIL_1.n16 ITAIL_1.n15 105.126
R7 ITAIL_1.n4 ITAIL_1.n3 103.823
R8 ITAIL_1.n6 ITAIL_1.n5 103.823
R9 ITAIL_1.n8 ITAIL_1.n7 103.823
R10 ITAIL_1.n10 ITAIL_1.n9 103.823
R11 ITAIL_1.n12 ITAIL_1.n11 103.823
R12 ITAIL_1.n14 ITAIL_1.n13 103.823
R13 ITAIL_1.n39 ITAIL_1.n38 103.823
R14 ITAIL_1.n78 ITAIL_1.n77 103.823
R15 ITAIL_1.n33 ITAIL_1.n32 103.823
R16 ITAIL_1.n31 ITAIL_1.n30 103.823
R17 ITAIL_1.n29 ITAIL_1.n28 103.823
R18 ITAIL_1.n27 ITAIL_1.n26 103.823
R19 ITAIL_1.n25 ITAIL_1.n24 103.823
R20 ITAIL_1.n46 ITAIL_1.n45 103.823
R21 ITAIL_1.n55 ITAIL_1.n54 103.823
R22 ITAIL_1.n71 ITAIL_1.n70 103.823
R23 ITAIL_1.n69 ITAIL_1.n68 103.823
R24 ITAIL_1.n72 ITAIL_1.n71 36.3254
R25 ITAIL_1.n77 ITAIL_1.t53 34.7404
R26 ITAIL_1.n57 ITAIL_1.n55 33.2561
R27 ITAIL_1.n47 ITAIL_1.n46 22.0563
R28 ITAIL_1.n40 ITAIL_1.n39 21.6519
R29 ITAIL_1.n3 ITAIL_1.n2 21.0894
R30 ITAIL_1.n5 ITAIL_1.n4 21.0894
R31 ITAIL_1.n7 ITAIL_1.n6 21.0894
R32 ITAIL_1.n9 ITAIL_1.n8 21.0894
R33 ITAIL_1.n11 ITAIL_1.n10 21.0894
R34 ITAIL_1.n13 ITAIL_1.n12 21.0894
R35 ITAIL_1.n15 ITAIL_1.n14 21.0894
R36 ITAIL_1.n79 ITAIL_1.n78 21.0894
R37 ITAIL_1.n34 ITAIL_1.n33 21.0894
R38 ITAIL_1.n32 ITAIL_1.n31 21.0894
R39 ITAIL_1.n30 ITAIL_1.n29 21.0894
R40 ITAIL_1.n28 ITAIL_1.n27 21.0894
R41 ITAIL_1.n26 ITAIL_1.n25 21.0894
R42 ITAIL_1.n24 ITAIL_1.n23 21.0894
R43 ITAIL_1.n45 ITAIL_1.n44 21.0894
R44 ITAIL_1.n54 ITAIL_1.n53 21.0894
R45 ITAIL_1.n70 ITAIL_1.n69 21.0894
R46 ITAIL_1.n2 ITAIL_1.t71 14.0165
R47 ITAIL_1.n3 ITAIL_1.t32 14.0165
R48 ITAIL_1.n4 ITAIL_1.t48 14.0165
R49 ITAIL_1.n5 ITAIL_1.t55 14.0165
R50 ITAIL_1.n6 ITAIL_1.t66 14.0165
R51 ITAIL_1.n7 ITAIL_1.t30 14.0165
R52 ITAIL_1.n8 ITAIL_1.t46 14.0165
R53 ITAIL_1.n9 ITAIL_1.t73 14.0165
R54 ITAIL_1.n10 ITAIL_1.t43 14.0165
R55 ITAIL_1.n11 ITAIL_1.t68 14.0165
R56 ITAIL_1.n12 ITAIL_1.t57 14.0165
R57 ITAIL_1.n13 ITAIL_1.t45 14.0165
R58 ITAIL_1.n14 ITAIL_1.t51 14.0165
R59 ITAIL_1.n15 ITAIL_1.t24 14.0165
R60 ITAIL_1.n33 ITAIL_1.t37 14.0165
R61 ITAIL_1.n32 ITAIL_1.t72 14.0165
R62 ITAIL_1.n31 ITAIL_1.t49 14.0165
R63 ITAIL_1.n30 ITAIL_1.t58 14.0165
R64 ITAIL_1.n29 ITAIL_1.t70 14.0165
R65 ITAIL_1.n28 ITAIL_1.t44 14.0165
R66 ITAIL_1.n27 ITAIL_1.t62 14.0165
R67 ITAIL_1.n26 ITAIL_1.t47 14.0165
R68 ITAIL_1.n25 ITAIL_1.t33 14.0165
R69 ITAIL_1.n24 ITAIL_1.t67 14.0165
R70 ITAIL_1.n23 ITAIL_1.t40 14.0165
R71 ITAIL_1.n44 ITAIL_1.t59 14.0165
R72 ITAIL_1.n45 ITAIL_1.t35 14.0165
R73 ITAIL_1.n46 ITAIL_1.t38 14.0165
R74 ITAIL_1.n53 ITAIL_1.t41 13.7245
R75 ITAIL_1.n54 ITAIL_1.t69 13.7245
R76 ITAIL_1.n55 ITAIL_1.t64 13.7245
R77 ITAIL_1.n71 ITAIL_1.t34 13.7245
R78 ITAIL_1.n70 ITAIL_1.t74 13.7245
R79 ITAIL_1.n69 ITAIL_1.t61 13.7245
R80 ITAIL_1.n39 ITAIL_1.t29 13.6515
R81 ITAIL_1.n38 ITAIL_1.t42 13.6515
R82 ITAIL_1.n85 ITAIL_1.t65 13.6515
R83 ITAIL_1.n77 ITAIL_1.t28 13.6515
R84 ITAIL_1.n78 ITAIL_1.t75 13.6515
R85 ITAIL_1.n79 ITAIL_1.t36 13.6515
R86 ITAIL_1.n40 ITAIL_1.t56 13.0378
R87 ITAIL_1.n87 ITAIL_1.t15 12.6295
R88 ITAIL_1.n86 ITAIL_1.t5 12.6295
R89 ITAIL_1.n0 ITAIL_1.t54 12.6295
R90 ITAIL_1.n59 ITAIL_1.t11 12.5565
R91 ITAIL_1.n63 ITAIL_1.t19 12.5565
R92 ITAIL_1.n81 ITAIL_1.t17 12.3375
R93 ITAIL_1.n80 ITAIL_1.t9 12.3375
R94 ITAIL_1.n64 ITAIL_1.t13 12.1915
R95 ITAIL_1.n52 ITAIL_1.t39 10.8639
R96 ITAIL_1.n48 ITAIL_1.t27 10.4542
R97 ITAIL_1.n22 ITAIL_1.t63 10.4093
R98 ITAIL_1.n57 ITAIL_1.n56 10.1427
R99 ITAIL_1.n18 ITAIL_1.t60 9.3445
R100 ITAIL_1.n58 ITAIL_1.t7 7.7385
R101 ITAIL_1.n62 ITAIL_1.n61 7.45611
R102 ITAIL_1.n106 ITAIL_1.n105 7.24501
R103 ITAIL_1.n58 ITAIL_1.n57 6.3515
R104 ITAIL_1.n41 ITAIL_1.t14 6.33405
R105 ITAIL_1.n52 ITAIL_1.n51 6.07308
R106 ITAIL_1.n88 ITAIL_1.n86 4.63315
R107 ITAIL_1.n73 ITAIL_1.n72 4.5005
R108 ITAIL_1.n62 ITAIL_1.n59 4.33237
R109 ITAIL_1.n82 ITAIL_1.n80 4.19412
R110 ITAIL_1.n88 ITAIL_1.n87 4.03194
R111 ITAIL_1.n63 ITAIL_1.n62 4.01149
R112 ITAIL_1.n82 ITAIL_1.n81 3.88348
R113 ITAIL_1.n105 ITAIL_1.n102 3.67213
R114 ITAIL_1.n96 ITAIL_1.n40 3.64368
R115 ITAIL_1.n49 ITAIL_1.n47 3.54502
R116 ITAIL_1.n49 ITAIL_1.n48 3.51942
R117 ITAIL_1.n92 ITAIL_1.n91 3.43549
R118 ITAIL_1.n83 ITAIL_1.n76 3.41085
R119 ITAIL_1.n37 ITAIL_1.n20 3.14528
R120 ITAIL_1.n102 ITAIL_1.t3 3.03383
R121 ITAIL_1.n102 ITAIL_1.n101 3.03383
R122 ITAIL_1.n104 ITAIL_1.t0 3.03383
R123 ITAIL_1.n104 ITAIL_1.n103 3.03383
R124 ITAIL_1.n100 ITAIL_1.t23 3.03383
R125 ITAIL_1.n100 ITAIL_1.n99 3.03383
R126 ITAIL_1.n98 ITAIL_1.t2 3.03383
R127 ITAIL_1.n98 ITAIL_1.n97 3.03383
R128 ITAIL_1.n20 ITAIL_1.n19 2.88564
R129 ITAIL_1.n51 ITAIL_1.n50 2.88451
R130 ITAIL_1.n111 ITAIL_1.n1 2.8805
R131 ITAIL_1.n106 ITAIL_1.n100 2.82159
R132 ITAIL_1.n107 ITAIL_1.n98 2.82159
R133 ITAIL_1.n105 ITAIL_1.n104 2.81922
R134 ITAIL_1.n61 ITAIL_1.t12 2.7305
R135 ITAIL_1.n61 ITAIL_1.n60 2.7305
R136 ITAIL_1.n91 ITAIL_1.t16 2.7305
R137 ITAIL_1.n91 ITAIL_1.n90 2.7305
R138 ITAIL_1.n76 ITAIL_1.t10 2.7305
R139 ITAIL_1.n76 ITAIL_1.n75 2.7305
R140 ITAIL_1.n19 ITAIL_1.n18 2.3365
R141 ITAIL_1.n37 ITAIL_1.n36 2.25242
R142 ITAIL_1.n93 ITAIL_1.n92 2.24675
R143 ITAIL_1.n17 ITAIL_1.n16 2.23635
R144 ITAIL_1.n36 ITAIL_1.n35 2.12238
R145 ITAIL_1.n83 ITAIL_1.n82 2.11998
R146 ITAIL_1.n35 ITAIL_1.n34 2.1175
R147 ITAIL_1.n66 ITAIL_1.n65 1.90845
R148 ITAIL_1.n108 ITAIL_1.n107 1.44061
R149 ITAIL_1.n84 ITAIL_1.n83 1.3863
R150 ITAIL_1.n89 ITAIL_1.n88 1.32705
R151 ITAIL_1.n35 ITAIL_1.n22 1.21129
R152 ITAIL_1.n74 ITAIL_1.n73 1.13048
R153 ITAIL_1.n96 ITAIL_1.n95 1.01644
R154 ITAIL_1.n111 ITAIL_1.n110 0.89823
R155 ITAIL_1.n65 ITAIL_1.n64 0.747091
R156 ITAIL_1.n109 ITAIL_1.n37 0.710424
R157 ITAIL_1.n1 ITAIL_1.n0 0.6575
R158 ITAIL_1.n72 ITAIL_1.n66 0.581182
R159 ITAIL_1.n107 ITAIL_1.n106 0.525071
R160 ITAIL_1.n109 ITAIL_1.n108 0.400171
R161 ITAIL_1.n68 ITAIL_1.n67 0.3655
R162 ITAIL_1.n95 ITAIL_1.n74 0.286359
R163 ITAIL_1.n95 ITAIL_1.n94 0.166826
R164 ITAIL_1.n108 ITAIL_1.n96 0.0964132
R165 ITAIL_1.n67 ITAIL_1.n1 0.0735
R166 ITAIL_1.n110 ITAIL_1.n109 0.0336328
R167 ITAIL_1.n42 ITAIL_1.n41 0.0250455
R168 ITAIL_1.n92 ITAIL_1.n89 0.0151731
R169 ITAIL_1.n94 ITAIL_1.n93 0.00905634
R170 ITAIL_1.n36 ITAIL_1.n21 0.00457413
R171 ITAIL_1 ITAIL_1.n111 0.00375301
R172 ITAIL_1.n73 ITAIL_1.n43 0.00356818
R173 ITAIL_1.n43 ITAIL_1.n42 0.00356818
R174 ITAIL_1.n51 ITAIL_1.n49 0.0025
R175 ITAIL_1.n20 ITAIL_1.n17 0.0015
R176 ITAIL_1.n93 ITAIL_1.n84 0.000816901
R177 SD3_1.n97 SD3_1.n7 3.48971
R178 SD3_1.n109 SD3_1.n3 3.48281
R179 SD3_1.n56 SD3_1.n55 3.07792
R180 SD3_1.n85 SD3_1.n27 3.07726
R181 SD3_1.n88 SD3_1.n22 3.07632
R182 SD3_1.n121 SD3_1.n118 3.07564
R183 SD3_1.n76 SD3_1.n42 3.0732
R184 SD3_1.n82 SD3_1.n32 3.07118
R185 SD3_1.n79 SD3_1.n37 3.06982
R186 SD3_1.n70 SD3_1.n44 3.06866
R187 SD3_1.n91 SD3_1.n17 3.06533
R188 SD3_1.n64 SD3_1.n49 3.06484
R189 SD3_1 SD3_1.n1 3.06384
R190 SD3_1.n58 SD3_1.n51 3.05987
R191 SD3_1.n100 SD3_1.n5 3.05915
R192 SD3_1.n94 SD3_1.n12 3.05307
R193 SD3_1.n12 SD3_1.n11 2.90211
R194 SD3_1.n102 SD3_1.n101 2.90208
R195 SD3_1.n120 SD3_1.t1 2.7305
R196 SD3_1.n120 SD3_1.n119 2.7305
R197 SD3_1.n118 SD3_1.t31 2.7305
R198 SD3_1.n118 SD3_1.n117 2.7305
R199 SD3_1.n106 SD3_1.t6 2.7305
R200 SD3_1.n106 SD3_1.n105 2.7305
R201 SD3_1.n9 SD3_1.t7 2.7305
R202 SD3_1.n9 SD3_1.n8 2.7305
R203 SD3_1.n14 SD3_1.t29 2.7305
R204 SD3_1.n14 SD3_1.n13 2.7305
R205 SD3_1.n19 SD3_1.t56 2.7305
R206 SD3_1.n19 SD3_1.n18 2.7305
R207 SD3_1.n24 SD3_1.t27 2.7305
R208 SD3_1.n24 SD3_1.n23 2.7305
R209 SD3_1.n29 SD3_1.t58 2.7305
R210 SD3_1.n29 SD3_1.n28 2.7305
R211 SD3_1.n34 SD3_1.t40 2.7305
R212 SD3_1.n34 SD3_1.n33 2.7305
R213 SD3_1.n39 SD3_1.t2 2.7305
R214 SD3_1.n39 SD3_1.n38 2.7305
R215 SD3_1.n73 SD3_1.t34 2.7305
R216 SD3_1.n73 SD3_1.n72 2.7305
R217 SD3_1.n46 SD3_1.t46 2.7305
R218 SD3_1.n46 SD3_1.n45 2.7305
R219 SD3_1.n66 SD3_1.t39 2.7305
R220 SD3_1.n66 SD3_1.n65 2.7305
R221 SD3_1.n60 SD3_1.t62 2.7305
R222 SD3_1.n60 SD3_1.n59 2.7305
R223 SD3_1.n53 SD3_1.t41 2.7305
R224 SD3_1.n53 SD3_1.n52 2.7305
R225 SD3_1.n55 SD3_1.t49 2.7305
R226 SD3_1.n55 SD3_1.n54 2.7305
R227 SD3_1.n51 SD3_1.t38 2.7305
R228 SD3_1.n51 SD3_1.n50 2.7305
R229 SD3_1.n49 SD3_1.t11 2.7305
R230 SD3_1.n49 SD3_1.n48 2.7305
R231 SD3_1.n44 SD3_1.t32 2.7305
R232 SD3_1.n44 SD3_1.n43 2.7305
R233 SD3_1.n42 SD3_1.t52 2.7305
R234 SD3_1.n42 SD3_1.n41 2.7305
R235 SD3_1.n37 SD3_1.t30 2.7305
R236 SD3_1.n37 SD3_1.n36 2.7305
R237 SD3_1.n32 SD3_1.t8 2.7305
R238 SD3_1.n32 SD3_1.n31 2.7305
R239 SD3_1.n27 SD3_1.t35 2.7305
R240 SD3_1.n27 SD3_1.n26 2.7305
R241 SD3_1.n22 SD3_1.t54 2.7305
R242 SD3_1.n22 SD3_1.n21 2.7305
R243 SD3_1.n17 SD3_1.t37 2.7305
R244 SD3_1.n17 SD3_1.n16 2.7305
R245 SD3_1.n7 SD3_1.t33 2.7305
R246 SD3_1.n7 SD3_1.n6 2.7305
R247 SD3_1.n5 SD3_1.t50 2.7305
R248 SD3_1.n5 SD3_1.n4 2.7305
R249 SD3_1.n3 SD3_1.t28 2.7305
R250 SD3_1.n3 SD3_1.n2 2.7305
R251 SD3_1.n1 SD3_1.t48 2.7305
R252 SD3_1.n1 SD3_1.n0 2.7305
R253 SD3_1.n113 SD3_1.t42 2.7305
R254 SD3_1.n113 SD3_1.n112 2.7305
R255 SD3_1.n56 SD3_1.n53 2.5571
R256 SD3_1.n121 SD3_1.n120 2.55706
R257 SD3_1.n102 SD3_1.t36 2.40707
R258 SD3_1.n12 SD3_1.t61 2.40704
R259 SD3_1.n108 SD3_1.n107 2.24937
R260 SD3_1.n104 SD3_1.n103 2.24505
R261 SD3_1.n62 SD3_1.n61 2.24478
R262 SD3_1.n68 SD3_1.n67 2.24478
R263 SD3_1.n75 SD3_1.n74 1.49476
R264 SD3_1.n87 SD3_1.n25 1.49463
R265 SD3_1.n116 SD3_1.n115 1.49463
R266 SD3_1.n81 SD3_1.n35 1.49463
R267 SD3_1.n90 SD3_1.n20 1.49463
R268 SD3_1.n69 SD3_1.n47 1.49439
R269 SD3_1.n84 SD3_1.n30 1.49439
R270 SD3_1.n78 SD3_1.n40 1.49439
R271 SD3_1.n93 SD3_1.n15 1.49439
R272 SD3_1.n96 SD3_1.n10 1.49439
R273 SD3_1.n40 SD3_1.n39 1.43788
R274 SD3_1.n74 SD3_1.n73 1.43788
R275 SD3_1.n10 SD3_1.n9 1.43741
R276 SD3_1.n25 SD3_1.n24 1.43741
R277 SD3_1.n30 SD3_1.n29 1.43741
R278 SD3_1.n47 SD3_1.n46 1.43741
R279 SD3_1.n20 SD3_1.n19 1.43705
R280 SD3_1.n107 SD3_1.n106 1.43694
R281 SD3_1.n35 SD3_1.n34 1.43694
R282 SD3_1.n67 SD3_1.n66 1.43694
R283 SD3_1.n15 SD3_1.n14 1.43673
R284 SD3_1.n61 SD3_1.n60 1.43673
R285 SD3_1.n114 SD3_1.n113 1.43607
R286 SD3_1.n103 SD3_1.n102 1.01023
R287 SD3_1.n108 SD3_1.n104 0.593824
R288 SD3_1.n57 SD3_1.n56 0.593282
R289 SD3_1.n69 SD3_1.n68 0.586829
R290 SD3_1.n99 SD3_1.n98 0.583544
R291 SD3_1.n63 SD3_1.n62 0.581823
R292 SD3_1.n78 SD3_1.n77 0.579925
R293 SD3_1.n122 SD3_1.n121 0.577695
R294 SD3_1.n93 SD3_1.n92 0.577272
R295 SD3_1.n84 SD3_1.n83 0.576023
R296 SD3_1.n90 SD3_1.n89 0.575664
R297 SD3_1.n96 SD3_1.n95 0.575142
R298 SD3_1.n81 SD3_1.n80 0.573011
R299 SD3_1.n87 SD3_1.n86 0.572285
R300 SD3_1.n116 SD3_1.n110 0.571741
R301 SD3_1.n75 SD3_1.n71 0.569825
R302 SD3_1.n71 SD3_1.n70 0.0254398
R303 SD3_1.n92 SD3_1.n91 0.0254398
R304 SD3_1 SD3_1.n122 0.0243554
R305 SD3_1.n80 SD3_1.n79 0.0232711
R306 SD3_1.n98 SD3_1.n97 0.0232711
R307 SD3_1.n110 SD3_1.n109 0.0232711
R308 SD3_1.n88 SD3_1.n87 0.0218667
R309 SD3_1.n86 SD3_1.n85 0.0211024
R310 SD3_1.n95 SD3_1.n94 0.0211024
R311 SD3_1.n82 SD3_1.n81 0.0200598
R312 SD3_1.n77 SD3_1.n76 0.0200181
R313 SD3_1.n76 SD3_1.n75 0.0190332
R314 SD3_1.n83 SD3_1.n82 0.0189337
R315 SD3_1.n85 SD3_1.n84 0.0186111
R316 SD3_1.n94 SD3_1.n93 0.0178882
R317 SD3_1.n89 SD3_1.n88 0.0178494
R318 SD3_1.n58 SD3_1.n57 0.0166884
R319 SD3_1.n68 SD3_1.n64 0.0166884
R320 SD3_1.n79 SD3_1.n78 0.0157195
R321 SD3_1.n97 SD3_1.n96 0.0157195
R322 SD3_1.n62 SD3_1.n58 0.0156041
R323 SD3_1.n64 SD3_1.n63 0.0156041
R324 SD3_1.n104 SD3_1.n100 0.0150649
R325 SD3_1 SD3_1.n116 0.0143027
R326 SD3_1.n70 SD3_1.n69 0.0142737
R327 SD3_1.n91 SD3_1.n90 0.0135538
R328 SD3_1.n109 SD3_1.n108 0.00641934
R329 SD3_1.n100 SD3_1.n99 0.00592169
R330 SD3_1.n114 SD3_1.n111 0.00585128
R331 SD3_1.n115 SD3_1.n114 0.00242298
R332 OUT_6.n31 OUT_6.t9 6.52669
R333 OUT_6.n46 OUT_6.n0 6.10941
R334 OUT_6.n31 OUT_6.n30 3.52028
R335 OUT_6.n33 OUT_6.n26 3.52028
R336 OUT_6.n35 OUT_6.n22 3.52028
R337 OUT_6.n37 OUT_6.n18 3.52028
R338 OUT_6.n39 OUT_6.n14 3.52028
R339 OUT_6.n41 OUT_6.n10 3.52028
R340 OUT_6.n43 OUT_6.n6 3.52028
R341 OUT_6.n45 OUT_6.n2 3.52028
R342 OUT_6.n44 OUT_6.n4 3.37941
R343 OUT_6.n42 OUT_6.n8 3.37941
R344 OUT_6.n40 OUT_6.n12 3.37941
R345 OUT_6.n38 OUT_6.n16 3.37941
R346 OUT_6.n36 OUT_6.n20 3.37941
R347 OUT_6.n34 OUT_6.n24 3.37941
R348 OUT_6.n32 OUT_6.n28 3.37941
R349 OUT_6.n4 OUT_6.t2 2.7305
R350 OUT_6.n4 OUT_6.n3 2.7305
R351 OUT_6.n8 OUT_6.t16 2.7305
R352 OUT_6.n8 OUT_6.n7 2.7305
R353 OUT_6.n12 OUT_6.t6 2.7305
R354 OUT_6.n12 OUT_6.n11 2.7305
R355 OUT_6.n16 OUT_6.t18 2.7305
R356 OUT_6.n16 OUT_6.n15 2.7305
R357 OUT_6.n20 OUT_6.t21 2.7305
R358 OUT_6.n20 OUT_6.n19 2.7305
R359 OUT_6.n24 OUT_6.t12 2.7305
R360 OUT_6.n24 OUT_6.n23 2.7305
R361 OUT_6.n28 OUT_6.t14 2.7305
R362 OUT_6.n28 OUT_6.n27 2.7305
R363 OUT_6.n30 OUT_6.t24 2.7305
R364 OUT_6.n30 OUT_6.n29 2.7305
R365 OUT_6.n26 OUT_6.t15 2.7305
R366 OUT_6.n26 OUT_6.n25 2.7305
R367 OUT_6.n22 OUT_6.t3 2.7305
R368 OUT_6.n22 OUT_6.n21 2.7305
R369 OUT_6.n18 OUT_6.t8 2.7305
R370 OUT_6.n18 OUT_6.n17 2.7305
R371 OUT_6.n14 OUT_6.t26 2.7305
R372 OUT_6.n14 OUT_6.n13 2.7305
R373 OUT_6.n10 OUT_6.t22 2.7305
R374 OUT_6.n10 OUT_6.n9 2.7305
R375 OUT_6.n6 OUT_6.t25 2.7305
R376 OUT_6.n6 OUT_6.n5 2.7305
R377 OUT_6.n2 OUT_6.t29 2.7305
R378 OUT_6.n2 OUT_6.n1 2.7305
R379 OUT_6.n46 OUT_6.n45 0.417773
R380 OUT_6.n45 OUT_6.n44 0.417773
R381 OUT_6.n44 OUT_6.n43 0.417773
R382 OUT_6.n43 OUT_6.n42 0.417773
R383 OUT_6.n42 OUT_6.n41 0.417773
R384 OUT_6.n41 OUT_6.n40 0.417773
R385 OUT_6.n40 OUT_6.n39 0.417773
R386 OUT_6.n39 OUT_6.n38 0.417773
R387 OUT_6.n38 OUT_6.n37 0.417773
R388 OUT_6.n37 OUT_6.n36 0.417773
R389 OUT_6.n36 OUT_6.n35 0.417773
R390 OUT_6.n35 OUT_6.n34 0.417773
R391 OUT_6.n34 OUT_6.n33 0.417773
R392 OUT_6.n33 OUT_6.n32 0.417773
R393 OUT_6.n32 OUT_6.n31 0.417773
R394 OUT_6 OUT_6.n46 0.133455
R395 VSS.t108 VSS.t109 733.941
R396 VSS.t128 VSS.t145 714.571
R397 VSS.t52 VSS.t36 714.571
R398 VSS.t8 VSS.t113 714.571
R399 VSS.t51 VSS.t48 714.571
R400 VSS.t48 VSS.t141 714.571
R401 VSS.t35 VSS.t195 714.571
R402 VSS.n217 VSS.t8 523.014
R403 VSS.t136 VSS.t115 439.074
R404 VSS.t20 VSS.t136 439.074
R405 VSS.t145 VSS.t20 439.074
R406 VSS.t174 VSS.t128 439.074
R407 VSS.t17 VSS.t174 439.074
R408 VSS.t36 VSS.t17 439.074
R409 VSS.t113 VSS.t52 439.074
R410 VSS.t141 VSS.t35 439.074
R411 VSS.t195 VSS.t15 439.074
R412 VSS.t15 VSS.t5 439.074
R413 VSS.t5 VSS.t108 439.074
R414 VSS.t109 VSS.t147 439.074
R415 VSS.t147 VSS.t116 439.074
R416 VSS.t116 VSS.t144 439.074
R417 VSS.n203 VSS.t51 391.723
R418 VSS.n73 VSS.t78 106.175
R419 VSS.n174 VSS.t82 100.996
R420 VSS.n63 VSS.t88 95.8172
R421 VSS.t71 VSS.t80 93.2276
R422 VSS.t77 VSS.t91 93.2276
R423 VSS.n160 VSS.t45 90.638
R424 VSS.t93 VSS.t103 82.869
R425 VSS.n170 VSS.t63 80.2794
R426 VSS.n248 VSS.t56 75.1001
R427 VSS.n43 VSS.t81 72.5105
R428 VSS.n72 VSS.t2 72.5105
R429 VSS.n126 VSS.t70 71.2156
R430 VSS.n156 VSS.t13 67.3312
R431 VSS.n49 VSS.t53 62.1519
R432 VSS.n66 VSS.t32 62.1519
R433 VSS.n167 VSS.t102 59.5623
R434 VSS.n250 VSS.t89 54.383
R435 VSS.n123 VSS.t74 50.4985
R436 VSS.n58 VSS.t84 49.2037
R437 VSS.n203 VSS.t25 47.3515
R438 VSS.n44 VSS.t96 38.8451
R439 VSS.n165 VSS.t77 38.8451
R440 VSS.n69 VSS.t68 38.8451
R441 VSS.n252 VSS.t90 33.6658
R442 VSS.n59 VSS.t75 33.6658
R443 VSS.n121 VSS.t95 29.7814
R444 VSS.n28 VSS.t106 28.4866
R445 VSS.n48 VSS.t30 28.4866
R446 VSS.n141 VSS.t85 28.4866
R447 VSS.n67 VSS.t86 28.4866
R448 VSS.n36 VSS.t98 23.3073
R449 VSS.n264 VSS.t100 23.3073
R450 VSS.n54 VSS.t37 18.128
R451 VSS.n162 VSS.t71 18.128
R452 VSS.n55 VSS.t104 15.5383
R453 VSS.t42 VSS.t58 14.2435
R454 VSS.t95 VSS.t79 14.2435
R455 VSS.t74 VSS.t28 14.2435
R456 VSS.t96 VSS.t99 14.2435
R457 VSS.t10 VSS.t66 14.2435
R458 VSS.n246 VSS.t87 12.9487
R459 VSS.n255 VSS.t72 12.9487
R460 VSS.n227 VSS.t97 11.6539
R461 VSS.n33 VSS.t105 10.3591
R462 VSS.n229 VSS.t83 9.06425
R463 VSS.n119 VSS.t42 9.06425
R464 VSS.n226 VSS.n225 8.54246
R465 VSS.n248 VSS.t40 7.76942
R466 VSS.n139 VSS.t101 7.76942
R467 VSS.n257 VSS.t0 7.76942
R468 VSS.n149 VSS.t92 7.76942
R469 VSS.n283 VSS.t110 7.64137
R470 VSS.n200 VSS.n199 7.09117
R471 VSS.n112 VSS.n26 6.51634
R472 VSS.n196 VSS.t114 6.41395
R473 VSS.n262 VSS.t164 6.41267
R474 VSS.n226 VSS.n185 6.41267
R475 VSS.n242 VSS.t67 6.41267
R476 VSS.n245 VSS.n182 6.41267
R477 VSS.n263 VSS.n179 6.41267
R478 VSS.n282 VSS.t159 6.41267
R479 VSS.n200 VSS.t9 6.26682
R480 VSS.n218 VSS.n217 6.21469
R481 VSS.n218 VSS.n216 5.8805
R482 VSS.n219 VSS.n215 5.8805
R483 VSS.n201 VSS.n198 5.8805
R484 VSS.n202 VSS.n197 5.8805
R485 VSS.n196 VSS.t178 5.8805
R486 VSS.n74 VSS.n73 5.32155
R487 VSS.n221 VSS.n203 5.2005
R488 VSS.n228 VSS.n227 5.2005
R489 VSS.n230 VSS.n229 5.2005
R490 VSS.n232 VSS.n231 5.2005
R491 VSS.n234 VSS.n233 5.2005
R492 VSS.n237 VSS.n236 5.2005
R493 VSS.n239 VSS.n238 5.2005
R494 VSS.n241 VSS.n240 5.2005
R495 VSS.n244 VSS.n243 5.2005
R496 VSS.n247 VSS.n246 5.2005
R497 VSS.n249 VSS.n248 5.2005
R498 VSS.n251 VSS.n250 5.2005
R499 VSS.n253 VSS.n252 5.2005
R500 VSS.n256 VSS.n255 5.2005
R501 VSS.n258 VSS.n257 5.2005
R502 VSS.n260 VSS.n259 5.2005
R503 VSS.n262 VSS.n261 5.2005
R504 VSS.n265 VSS.n264 5.2005
R505 VSS.n267 VSS.n266 5.2005
R506 VSS.n269 VSS.n268 5.2005
R507 VSS.n272 VSS.n271 5.2005
R508 VSS.n275 VSS.n274 5.2005
R509 VSS.n277 VSS.n276 5.2005
R510 VSS.n279 VSS.n278 5.2005
R511 VSS.n281 VSS.n280 5.2005
R512 VSS.n30 VSS.n28 5.2005
R513 VSS.n108 VSS.n33 5.2005
R514 VSS.n106 VSS.n36 5.2005
R515 VSS.n105 VSS.n37 5.2005
R516 VSS.n104 VSS.n38 5.2005
R517 VSS.n103 VSS.n39 5.2005
R518 VSS.n101 VSS.n42 5.2005
R519 VSS.n100 VSS.n43 5.2005
R520 VSS.n99 VSS.n44 5.2005
R521 VSS.n97 VSS.n47 5.2005
R522 VSS.n96 VSS.n48 5.2005
R523 VSS.n95 VSS.n49 5.2005
R524 VSS.n94 VSS.n50 5.2005
R525 VSS.n92 VSS.n53 5.2005
R526 VSS.n91 VSS.n54 5.2005
R527 VSS.n90 VSS.n55 5.2005
R528 VSS.n88 VSS.n58 5.2005
R529 VSS.n87 VSS.t93 5.2005
R530 VSS.n86 VSS.n59 5.2005
R531 VSS.n83 VSS.n62 5.2005
R532 VSS.n81 VSS.n63 5.2005
R533 VSS.n79 VSS.n66 5.2005
R534 VSS.n78 VSS.n67 5.2005
R535 VSS.n77 VSS.n68 5.2005
R536 VSS.n76 VSS.n69 5.2005
R537 VSS.n74 VSS.n72 5.2005
R538 VSS.n114 VSS.n113 5.2005
R539 VSS.n117 VSS.n116 5.2005
R540 VSS.n120 VSS.n119 5.2005
R541 VSS.n122 VSS.n121 5.2005
R542 VSS.n124 VSS.n123 5.2005
R543 VSS.n127 VSS.n126 5.2005
R544 VSS.n130 VSS.n129 5.2005
R545 VSS.n132 VSS.n131 5.2005
R546 VSS.n135 VSS.n134 5.2005
R547 VSS.n137 VSS.n136 5.2005
R548 VSS.n140 VSS.n139 5.2005
R549 VSS.n142 VSS.n141 5.2005
R550 VSS.n145 VSS.n144 5.2005
R551 VSS.n147 VSS.n146 5.2005
R552 VSS.n150 VSS.n149 5.2005
R553 VSS.n152 VSS.n151 5.2005
R554 VSS.n155 VSS.n154 5.2005
R555 VSS.n158 VSS.n157 5.2005
R556 VSS.n161 VSS.n160 5.2005
R557 VSS.n163 VSS.n162 5.2005
R558 VSS.n166 VSS.n165 5.2005
R559 VSS.n168 VSS.n167 5.2005
R560 VSS.n171 VSS.n170 5.2005
R561 VSS.n47 VSS.t10 5.17978
R562 VSS.n68 VSS.t107 5.17978
R563 VSS.n112 VSS.n111 4.99464
R564 VSS.n30 VSS.n29 4.5005
R565 VSS.n213 VSS.n212 3.78833
R566 VSS.n190 VSS.n189 3.78833
R567 VSS.n169 VSS.n3 3.7355
R568 VSS.n159 VSS.n7 3.7355
R569 VSS.n148 VSS.n11 3.7355
R570 VSS.n138 VSS.n15 3.7355
R571 VSS.n128 VSS.n19 3.7355
R572 VSS.n118 VSS.n23 3.7355
R573 VSS.n195 VSS.n194 3.71473
R574 VSS.n115 VSS.n25 3.7042
R575 VSS.n125 VSS.n21 3.7042
R576 VSS.n133 VSS.n17 3.7042
R577 VSS.n143 VSS.n13 3.7042
R578 VSS.n153 VSS.n9 3.7042
R579 VSS.n164 VSS.n5 3.7042
R580 VSS.n172 VSS.n1 3.7042
R581 VSS.n235 VSS.n184 3.68267
R582 VSS.n254 VSS.n181 3.68267
R583 VSS.n273 VSS.n178 3.68267
R584 VSS.n208 VSS.n207 3.67443
R585 VSS.n75 VSS.n71 3.64941
R586 VSS.n80 VSS.n65 3.64941
R587 VSS.n84 VSS.n61 3.64941
R588 VSS.n89 VSS.n57 3.64941
R589 VSS.n93 VSS.n52 3.64941
R590 VSS.n98 VSS.n46 3.64941
R591 VSS.n102 VSS.n41 3.64941
R592 VSS.n107 VSS.n35 3.64941
R593 VSS.n213 VSS.n210 3.1505
R594 VSS.n208 VSS.n205 3.1505
R595 VSS.n190 VSS.n187 3.1505
R596 VSS.n195 VSS.n192 3.1505
R597 VSS.n210 VSS.t148 2.7305
R598 VSS.n210 VSS.n209 2.7305
R599 VSS.n212 VSS.t157 2.7305
R600 VSS.n212 VSS.n211 2.7305
R601 VSS.n207 VSS.t16 2.7305
R602 VSS.n207 VSS.n206 2.7305
R603 VSS.n205 VSS.t119 2.7305
R604 VSS.n205 VSS.n204 2.7305
R605 VSS.n184 VSS.t138 2.7305
R606 VSS.n184 VSS.n183 2.7305
R607 VSS.n181 VSS.t191 2.7305
R608 VSS.n181 VSS.n180 2.7305
R609 VSS.n178 VSS.t171 2.7305
R610 VSS.n178 VSS.n177 2.7305
R611 VSS.n187 VSS.t137 2.7305
R612 VSS.n187 VSS.n186 2.7305
R613 VSS.n189 VSS.t146 2.7305
R614 VSS.n189 VSS.n188 2.7305
R615 VSS.n194 VSS.t175 2.7305
R616 VSS.n194 VSS.n193 2.7305
R617 VSS.n192 VSS.t192 2.7305
R618 VSS.n192 VSS.n191 2.7305
R619 VSS.n71 VSS.t69 2.7305
R620 VSS.n71 VSS.n70 2.7305
R621 VSS.n65 VSS.t179 2.7305
R622 VSS.n65 VSS.n64 2.7305
R623 VSS.n61 VSS.t14 2.7305
R624 VSS.n61 VSS.n60 2.7305
R625 VSS.n57 VSS.t1 2.7305
R626 VSS.n57 VSS.n56 2.7305
R627 VSS.n52 VSS.t57 2.7305
R628 VSS.n52 VSS.n51 2.7305
R629 VSS.n46 VSS.t200 2.7305
R630 VSS.n46 VSS.n45 2.7305
R631 VSS.n41 VSS.t59 2.7305
R632 VSS.n41 VSS.n40 2.7305
R633 VSS.n35 VSS.t186 2.7305
R634 VSS.n35 VSS.n34 2.7305
R635 VSS.n25 VSS.t158 2.7305
R636 VSS.n25 VSS.n24 2.7305
R637 VSS.n21 VSS.t29 2.7305
R638 VSS.n21 VSS.n20 2.7305
R639 VSS.n17 VSS.t31 2.7305
R640 VSS.n17 VSS.n16 2.7305
R641 VSS.n13 VSS.t135 2.7305
R642 VSS.n13 VSS.n12 2.7305
R643 VSS.n9 VSS.t187 2.7305
R644 VSS.n9 VSS.n8 2.7305
R645 VSS.n5 VSS.t126 2.7305
R646 VSS.n5 VSS.n4 2.7305
R647 VSS.n1 VSS.t165 2.7305
R648 VSS.n1 VSS.n0 2.7305
R649 VSS.n3 VSS.t127 2.7305
R650 VSS.n3 VSS.n2 2.7305
R651 VSS.n7 VSS.t188 2.7305
R652 VSS.n7 VSS.n6 2.7305
R653 VSS.n11 VSS.t168 2.7305
R654 VSS.n11 VSS.n10 2.7305
R655 VSS.n15 VSS.t41 2.7305
R656 VSS.n15 VSS.n14 2.7305
R657 VSS.n19 VSS.t149 2.7305
R658 VSS.n19 VSS.n18 2.7305
R659 VSS.n23 VSS.t154 2.7305
R660 VSS.n23 VSS.n22 2.7305
R661 VSS.n32 VSS.n31 2.60175
R662 VSS.n110 VSS.n32 2.601
R663 VSS.n176 VSS.n175 2.6005
R664 VSS.n175 VSS.n174 2.6005
R665 VSS.n227 VSS.t73 2.59014
R666 VSS.n116 VSS.t60 2.59014
R667 VSS.n157 VSS.n156 2.59014
R668 VSS.n266 VSS.t76 2.59014
R669 VSS.n160 VSS.t94 2.59014
R670 VSS.n271 VSS.n270 2.59014
R671 VSS.n30 VSS.n27 2.15773
R672 VSS.n283 VSS.n282 1.43392
R673 VSS.n214 VSS.n213 0.96262
R674 VSS.n114 VSS.n112 0.661796
R675 VSS.n175 VSS.n173 0.655471
R676 VSS.n219 VSS.n218 0.5873
R677 VSS.n202 VSS.n201 0.506362
R678 VSS.n225 VSS.n190 0.491587
R679 VSS.n224 VSS.n223 0.4638
R680 VSS.n220 VSS.n214 0.46349
R681 VSS.n225 VSS.n224 0.462607
R682 VSS.n220 VSS.n219 0.4559
R683 VSS.n224 VSS.n195 0.438385
R684 VSS.n32 VSS.n30 0.426384
R685 VSS.n223 VSS.n196 0.4145
R686 VSS.n214 VSS.n208 0.407107
R687 VSS.n222 VSS.n202 0.393086
R688 VSS.n221 VSS.n220 0.36591
R689 VSS.n201 VSS.n200 0.230155
R690 VSS.n223 VSS.n222 0.225254
R691 VSS VSS.n283 0.183461
R692 VSS.n106 VSS.n105 0.121553
R693 VSS.n105 VSS.n104 0.121553
R694 VSS.n104 VSS.n103 0.121553
R695 VSS.n101 VSS.n100 0.121553
R696 VSS.n100 VSS.n99 0.121553
R697 VSS.n97 VSS.n96 0.121553
R698 VSS.n96 VSS.n95 0.121553
R699 VSS.n95 VSS.n94 0.121553
R700 VSS.n92 VSS.n91 0.121553
R701 VSS.n91 VSS.n90 0.121553
R702 VSS.n88 VSS.n87 0.121553
R703 VSS.n87 VSS.n86 0.121553
R704 VSS.n86 VSS.n85 0.121553
R705 VSS.n83 VSS.n82 0.121553
R706 VSS.n82 VSS.n81 0.121553
R707 VSS.n79 VSS.n78 0.121553
R708 VSS.n78 VSS.n77 0.121553
R709 VSS.n77 VSS.n76 0.121553
R710 VSS.n102 VSS.n101 0.118395
R711 VSS.n230 VSS.n228 0.116289
R712 VSS.n232 VSS.n230 0.116289
R713 VSS.n234 VSS.n232 0.116289
R714 VSS.n239 VSS.n237 0.116289
R715 VSS.n241 VSS.n239 0.116289
R716 VSS.n249 VSS.n247 0.116289
R717 VSS.n251 VSS.n249 0.116289
R718 VSS.n253 VSS.n251 0.116289
R719 VSS.n258 VSS.n256 0.116289
R720 VSS.n260 VSS.n258 0.116289
R721 VSS.n262 VSS.n260 0.116289
R722 VSS.n267 VSS.n265 0.116289
R723 VSS.n269 VSS.n267 0.116289
R724 VSS.n272 VSS.n269 0.116289
R725 VSS.n277 VSS.n275 0.116289
R726 VSS.n279 VSS.n277 0.116289
R727 VSS.n281 VSS.n279 0.116289
R728 VSS.n122 VSS.n120 0.116289
R729 VSS.n124 VSS.n122 0.116289
R730 VSS.n132 VSS.n130 0.116289
R731 VSS.n137 VSS.n135 0.116289
R732 VSS.n142 VSS.n140 0.116289
R733 VSS.n147 VSS.n145 0.116289
R734 VSS.n152 VSS.n150 0.116289
R735 VSS.n158 VSS.n155 0.116289
R736 VSS.n163 VSS.n161 0.116289
R737 VSS.n168 VSS.n166 0.116289
R738 VSS.n242 VSS.n241 0.115763
R739 VSS.n109 VSS.n108 0.115237
R740 VSS.n133 VSS.n132 0.109974
R741 VSS.n166 VSS.n164 0.107868
R742 VSS.n93 VSS.n92 0.106816
R743 VSS.n84 VSS.n83 0.0952368
R744 VSS.n81 VSS.n80 0.0931316
R745 VSS.n130 VSS.n128 0.0915526
R746 VSS.n150 VSS.n148 0.0910263
R747 VSS.n172 VSS.n171 0.0910263
R748 VSS.n127 VSS.n125 0.0889211
R749 VSS.n171 VSS.n169 0.0868158
R750 VSS.n75 VSS.n74 0.0836579
R751 VSS.n237 VSS.n235 0.0831316
R752 VSS.n256 VSS.n254 0.0826053
R753 VSS.n90 VSS.n89 0.0815526
R754 VSS.n275 VSS.n273 0.0783947
R755 VSS.n143 VSS.n142 0.0762895
R756 VSS.n155 VSS.n153 0.0741842
R757 VSS.n263 VSS.n262 0.0720789
R758 VSS.n99 VSS.n98 0.0699737
R759 VSS.n245 VSS.n244 0.0678684
R760 VSS.n107 VSS.n106 0.0636579
R761 VSS.n159 VSS.n158 0.0636579
R762 VSS.n222 VSS.n221 0.062959
R763 VSS.n115 VSS.n114 0.0615526
R764 VSS.n138 VSS.n137 0.0594474
R765 VSS.n118 VSS.n117 0.058921
R766 VSS.n108 VSS.n107 0.0583947
R767 VSS.n120 VSS.n118 0.0578684
R768 VSS.n140 VSS.n138 0.0573421
R769 VSS.n117 VSS.n115 0.0552368
R770 VSS.n161 VSS.n159 0.0531316
R771 VSS.n98 VSS.n97 0.052079
R772 VSS.n228 VSS.n226 0.0494474
R773 VSS.n247 VSS.n245 0.0489211
R774 VSS.n265 VSS.n263 0.0447105
R775 VSS.n153 VSS.n152 0.0426053
R776 VSS.n89 VSS.n88 0.0405
R777 VSS.n145 VSS.n143 0.0405
R778 VSS.n273 VSS.n272 0.0383947
R779 VSS.n76 VSS.n75 0.0383947
R780 VSS.n254 VSS.n253 0.0341842
R781 VSS.n235 VSS.n234 0.0336579
R782 VSS.n169 VSS.n168 0.0299737
R783 VSS.n80 VSS.n79 0.0289211
R784 VSS.n125 VSS.n124 0.0278684
R785 VSS.n85 VSS.n84 0.0268158
R786 VSS.n148 VSS.n147 0.0257632
R787 VSS.n176 VSS.n172 0.0257632
R788 VSS.n128 VSS.n127 0.0252368
R789 VSS.n111 VSS.n110 0.0231316
R790 VSS.n94 VSS.n93 0.0152368
R791 VSS.n164 VSS.n163 0.00892105
R792 VSS VSS.n176 0.00892105
R793 VSS.n110 VSS.n109 0.00681579
R794 VSS.n135 VSS.n133 0.00681579
R795 VSS.n282 VSS.n281 0.00471053
R796 VSS.n103 VSS.n102 0.00365789
R797 VSS.n244 VSS.n242 0.00102632
R798 ITAIL.n11 ITAIL.n6 333.663
R799 ITAIL.n7 ITAIL.t7 116.817
R800 ITAIL.n9 ITAIL.n8 103.823
R801 ITAIL.n2 ITAIL.t6 97.648
R802 ITAIL.n6 ITAIL.n5 90.8936
R803 ITAIL.n11 ITAIL.n10 88.6306
R804 ITAIL.n4 ITAIL.n3 84.9459
R805 ITAIL.n8 ITAIL.n7 48.8699
R806 ITAIL.n10 ITAIL.n9 47.0449
R807 ITAIL.n3 ITAIL.n2 38.4914
R808 ITAIL.n5 ITAIL.n4 38.4914
R809 ITAIL ITAIL.t8 27.414
R810 ITAIL.t7 ITAIL.t10 23.7985
R811 ITAIL.t14 ITAIL.t13 23.7985
R812 ITAIL.t12 ITAIL.t20 23.7985
R813 ITAIL.t2 ITAIL.t3 23.7985
R814 ITAIL.t9 ITAIL.t22 23.7985
R815 ITAIL.t6 ITAIL.t18 23.7985
R816 ITAIL.t11 ITAIL.t15 23.7985
R817 ITAIL.t16 ITAIL.t21 23.7985
R818 ITAIL.t23 ITAIL.t19 23.7985
R819 ITAIL.t5 ITAIL.t24 23.7985
R820 ITAIL.n7 ITAIL.t14 12.9945
R821 ITAIL.n8 ITAIL.t12 12.9945
R822 ITAIL.n9 ITAIL.t2 12.9945
R823 ITAIL.n10 ITAIL.t9 12.9945
R824 ITAIL.t8 ITAIL.n11 12.7755
R825 ITAIL.n2 ITAIL.t11 12.7025
R826 ITAIL.n3 ITAIL.t16 12.7025
R827 ITAIL.n4 ITAIL.t23 12.7025
R828 ITAIL.n5 ITAIL.t5 12.7025
R829 ITAIL.n6 ITAIL.t17 10.8045
R830 ITAIL.n1 ITAIL.t1 10.1411
R831 ITAIL.n0 ITAIL.t0 8.6875
R832 ITAIL.n0 ITAIL.t4 7.3735
R833 ITAIL ITAIL.n1 4.95899
R834 ITAIL.n1 ITAIL.n0 2.47975
R835 G2_1.n3 G2_1.n2 102.993
R836 G2_1.n5 G2_1.n4 101.566
R837 G2_1.n8 G2_1.n7 99.4048
R838 G2_1.n10 G2_1.n9 99.4048
R839 G2_1.n12 G2_1.n6 70.7294
R840 G2_1.n11 G2_1.n10 39.5325
R841 G2_1.n12 G2_1.n11 39.4595
R842 G2_1.n6 G2_1.n5 37.7091
R843 G2_1.n2 G2_1.t24 29.4988
R844 G2_1.n7 G2_1.t25 29.1477
R845 G2_1.t24 G2_1.t23 23.7985
R846 G2_1.t9 G2_1.t6 23.7985
R847 G2_1.t5 G2_1.t22 23.7985
R848 G2_1.t19 G2_1.t13 23.7985
R849 G2_1.t14 G2_1.t3 23.7985
R850 G2_1.t25 G2_1.t21 23.7985
R851 G2_1.t16 G2_1.t12 23.7985
R852 G2_1.t4 G2_1.t8 23.7985
R853 G2_1.t11 G2_1.t10 23.7985
R854 G2_1.t15 G2_1.t17 23.7985
R855 G2_1.n4 G2_1.n3 16.5048
R856 G2_1.n9 G2_1.n8 16.1537
R857 G2_1.n11 G2_1.t20 13.1405
R858 G2_1.n6 G2_1.t18 13.0675
R859 G2_1.t1 G2_1.n12 13.0675
R860 G2_1.n2 G2_1.t9 12.9945
R861 G2_1.n3 G2_1.t5 12.9945
R862 G2_1.n4 G2_1.t19 12.9945
R863 G2_1.n5 G2_1.t14 12.9945
R864 G2_1.n7 G2_1.t16 12.9945
R865 G2_1.n8 G2_1.t4 12.9945
R866 G2_1.n9 G2_1.t11 12.9945
R867 G2_1.n10 G2_1.t15 12.9945
R868 G2_1.n14 G2_1.t7 12.6295
R869 G2_1.n13 G2_1.t1 10.8045
R870 G2_1.n15 G2_1.n14 4.0005
R871 G2_1.n15 G2_1.n1 3.43609
R872 G2_1.n1 G2_1.t2 2.7305
R873 G2_1.n1 G2_1.n0 2.7305
R874 G2_1.n14 G2_1.n13 0.3655
R875 G2_1 G2_1.n15 0.0065
R876 G1_1.n25 G1_1.t35 113.573
R877 G1_1.n0 G1_1.t31 113.573
R878 G1_1.n27 G1_1.n26 101.016
R879 G1_1.n31 G1_1.n30 101.016
R880 G1_1.n29 G1_1.n28 101.016
R881 G1_1.n4 G1_1.n3 101.016
R882 G1_1.n2 G1_1.n1 101.016
R883 G1_1.n6 G1_1.n5 101.016
R884 G1_1.n6 G1_1.n2 67.0816
R885 G1_1.n31 G1_1.n27 62.3464
R886 G1_1.n26 G1_1.n25 20.5194
R887 G1_1.n30 G1_1.n29 20.5194
R888 G1_1.n5 G1_1.n4 20.5194
R889 G1_1.n1 G1_1.n0 20.5194
R890 G1_1.n25 G1_1.t29 12.5565
R891 G1_1.n26 G1_1.t32 12.5565
R892 G1_1.n27 G1_1.t26 12.5565
R893 G1_1.n30 G1_1.t0 12.5565
R894 G1_1.n29 G1_1.t4 12.5565
R895 G1_1.n28 G1_1.t12 12.5565
R896 G1_1.n3 G1_1.t8 12.5565
R897 G1_1.n4 G1_1.t14 12.5565
R898 G1_1.n5 G1_1.t6 12.5565
R899 G1_1.n0 G1_1.t30 12.5565
R900 G1_1.n1 G1_1.t28 12.5565
R901 G1_1.n2 G1_1.t27 12.5565
R902 G1_1.n32 G1_1.t10 10.2935
R903 G1_1.n7 G1_1.t2 10.2205
R904 G1_1.n33 G1_1.n32 4.12693
R905 G1_1 G1_1.n8 4.0015
R906 G1_1.n10 G1_1.t22 3.03383
R907 G1_1.n10 G1_1.n9 3.03383
R908 G1_1.n12 G1_1.t7 3.03383
R909 G1_1.n12 G1_1.n11 3.03383
R910 G1_1.n14 G1_1.t18 3.03383
R911 G1_1.n14 G1_1.n13 3.03383
R912 G1_1.n16 G1_1.t9 3.03383
R913 G1_1.n16 G1_1.n15 3.03383
R914 G1_1.n18 G1_1.t21 3.03383
R915 G1_1.n18 G1_1.n17 3.03383
R916 G1_1.n20 G1_1.t5 3.03383
R917 G1_1.n20 G1_1.n19 3.03383
R918 G1_1.n22 G1_1.t16 3.03383
R919 G1_1.n22 G1_1.n21 3.03383
R920 G1_1.n24 G1_1.t11 3.03383
R921 G1_1.n24 G1_1.n23 3.03383
R922 G1_1.n39 G1_1.n12 2.82159
R923 G1_1.n38 G1_1.n14 2.82159
R924 G1_1.n37 G1_1.n16 2.82159
R925 G1_1.n36 G1_1.n18 2.82159
R926 G1_1.n35 G1_1.n20 2.82159
R927 G1_1.n34 G1_1.n22 2.82159
R928 G1_1.n40 G1_1.n10 2.78833
R929 G1_1.n33 G1_1.n24 2.78833
R930 G1_1.n32 G1_1.n31 2.2635
R931 G1_1.n8 G1_1.n6 2.2635
R932 G1_1.n35 G1_1.n34 0.798761
R933 G1_1.n36 G1_1.n35 0.798761
R934 G1_1.n37 G1_1.n36 0.798761
R935 G1_1.n38 G1_1.n37 0.798761
R936 G1_1.n39 G1_1.n38 0.798761
R937 G1_1.n40 G1_1.n39 0.786618
R938 G1_1.n34 G1_1.n33 0.786618
R939 G1_1 G1_1.n40 0.0949286
R940 G1_1.n8 G1_1.n7 0.0735
R941 VDD.n78 VDD.t55 166.102
R942 VDD.n96 VDD.t22 161.018
R943 VDD.n64 VDD.t45 159.322
R944 VDD.n80 VDD.t54 155.933
R945 VDD.n97 VDD.t53 150.847
R946 VDD.n62 VDD.t41 149.154
R947 VDD.n82 VDD.t2 145.763
R948 VDD.n98 VDD.t51 140.679
R949 VDD.n60 VDD.t32 138.983
R950 VDD.n3 VDD.t0 135.114
R951 VDD.n99 VDD.t20 130.508
R952 VDD.n102 VDD.t9 120.34
R953 VDD.n75 VDD.t25 118.865
R954 VDD.n4 VDD.t47 118.644
R955 VDD.n46 VDD.t50 118.644
R956 VDD.n73 VDD.t35 111.865
R957 VDD.n103 VDD.t44 110.169
R958 VDD.n6 VDD.t43 108.475
R959 VDD.n44 VDD.t49 108.475
R960 VDD.n104 VDD.t48 100.001
R961 VDD.n8 VDD.t18 98.3056
R962 VDD.n42 VDD.t12 98.3056
R963 VDD.n51 VDD.t30 98.3056
R964 VDD.n105 VDD.t15 89.831
R965 VDD.n11 VDD.t7 88.1361
R966 VDD.n13 VDD.t42 77.9666
R967 VDD.n28 VDD.t40 77.9666
R968 VDD.n15 VDD.t52 67.7971
R969 VDD.n26 VDD.t46 67.7971
R970 VDD.n33 VDD.t5 67.7971
R971 VDD.n17 VDD.t28 57.6276
R972 VDD.n24 VDD.t37 57.6276
R973 VDD.n23 VDD.n22 8.30127
R974 VDD.n84 VDD.t3 7.67003
R975 VDD.n76 VDD.n73 6.3005
R976 VDD.n52 VDD.n51 6.3005
R977 VDD.n34 VDD.n33 6.3005
R978 VDD.n5 VDD.n4 6.3005
R979 VDD.n7 VDD.n6 6.3005
R980 VDD.n9 VDD.n8 6.3005
R981 VDD.n12 VDD.n11 6.3005
R982 VDD.n14 VDD.n13 6.3005
R983 VDD.n16 VDD.n15 6.3005
R984 VDD.n18 VDD.n17 6.3005
R985 VDD.n21 VDD.n20 6.3005
R986 VDD.n25 VDD.n24 6.3005
R987 VDD.n27 VDD.n26 6.3005
R988 VDD.n29 VDD.n28 6.3005
R989 VDD.n43 VDD.n42 6.3005
R990 VDD.n45 VDD.n44 6.3005
R991 VDD.n47 VDD.n46 6.3005
R992 VDD.n61 VDD.n60 6.3005
R993 VDD.n63 VDD.n62 6.3005
R994 VDD.n65 VDD.n64 6.3005
R995 VDD.n79 VDD.n78 6.3005
R996 VDD.n81 VDD.n80 6.3005
R997 VDD.n83 VDD.n82 6.3005
R998 VDD.n114 VDD.n96 6.3005
R999 VDD.n113 VDD.n97 6.3005
R1000 VDD.n112 VDD.n98 6.3005
R1001 VDD.n111 VDD.n99 6.3005
R1002 VDD.n109 VDD.n102 6.3005
R1003 VDD.n108 VDD.n103 6.3005
R1004 VDD.n107 VDD.n104 6.3005
R1005 VDD.n106 VDD.n105 6.3005
R1006 VDD.n90 VDD.n87 6.3005
R1007 VDD.n93 VDD.n86 6.3005
R1008 VDD.n106 VDD.t16 6.18063
R1009 VDD.n3 VDD.n2 6.10984
R1010 VDD.n115 VDD.n95 6.09557
R1011 VDD.n19 VDD.t29 6.09557
R1012 VDD.n72 VDD.n71 4.98502
R1013 VDD.n52 VDD.n50 4.5005
R1014 VDD.n34 VDD.n32 4.5005
R1015 VDD.n90 VDD.n89 4.5005
R1016 VDD.n59 VDD.n58 4.26092
R1017 VDD.n41 VDD.n40 4.24066
R1018 VDD.n58 VDD.n57 3.2271
R1019 VDD.n40 VDD.n39 3.20234
R1020 VDD.n71 VDD.n70 3.17695
R1021 VDD.n54 VDD.n53 3.15175
R1022 VDD.n93 VDD.n92 3.15175
R1023 VDD.n69 VDD.n68 3.15175
R1024 VDD.n36 VDD.n35 3.15175
R1025 VDD.n37 VDD.n36 3.151
R1026 VDD.n92 VDD.n91 3.151
R1027 VDD.n55 VDD.n54 3.151
R1028 VDD.n68 VDD.n67 3.151
R1029 VDD.n110 VDD.n101 3.06224
R1030 VDD.n10 VDD.n1 3.06224
R1031 VDD.n101 VDD.t21 3.03383
R1032 VDD.n101 VDD.n100 3.03383
R1033 VDD.n1 VDD.t19 3.03383
R1034 VDD.n1 VDD.n0 3.03383
R1035 VDD.n71 VDD.t36 2.69573
R1036 VDD.n40 VDD.t6 2.66058
R1037 VDD.n58 VDD.t31 2.62483
R1038 VDD.n77 VDD.n76 2.62147
R1039 VDD.n34 VDD.n31 1.88512
R1040 VDD.n76 VDD.n74 1.83127
R1041 VDD.n88 VDD.n86 1.72358
R1042 VDD.n52 VDD.n49 1.56204
R1043 VDD.n54 VDD.n52 1.12174
R1044 VDD.n92 VDD.n90 0.724621
R1045 VDD.n36 VDD.n34 0.525399
R1046 VDD.n76 VDD.n75 0.415309
R1047 VDD.n5 VDD.n3 0.115744
R1048 VDD.n7 VDD.n5 0.115744
R1049 VDD.n9 VDD.n7 0.115744
R1050 VDD.n14 VDD.n12 0.115744
R1051 VDD.n16 VDD.n14 0.115744
R1052 VDD.n18 VDD.n16 0.115744
R1053 VDD.n27 VDD.n25 0.115744
R1054 VDD.n29 VDD.n27 0.115744
R1055 VDD.n45 VDD.n43 0.115744
R1056 VDD.n47 VDD.n45 0.115744
R1057 VDD.n63 VDD.n61 0.115744
R1058 VDD.n65 VDD.n63 0.115744
R1059 VDD.n81 VDD.n79 0.115744
R1060 VDD.n83 VDD.n81 0.115744
R1061 VDD.n114 VDD.n113 0.115744
R1062 VDD.n113 VDD.n112 0.115744
R1063 VDD.n112 VDD.n111 0.115744
R1064 VDD.n109 VDD.n108 0.115744
R1065 VDD.n108 VDD.n107 0.115744
R1066 VDD.n107 VDD.n106 0.115744
R1067 VDD.n30 VDD.n29 0.109159
R1068 VDD.n79 VDD.n77 0.106804
R1069 VDD.n48 VDD.n47 0.105866
R1070 VDD.n111 VDD.n110 0.0987317
R1071 VDD.n66 VDD.n65 0.0970854
R1072 VDD VDD.n115 0.0959878
R1073 VDD.n61 VDD.n59 0.0957073
R1074 VDD.n84 VDD.n83 0.0953491
R1075 VDD.n43 VDD.n41 0.0913202
R1076 VDD.n10 VDD.n9 0.0883049
R1077 VDD.n25 VDD.n23 0.0789756
R1078 VDD.n19 VDD.n18 0.0751341
R1079 VDD.n23 VDD.n21 0.0723902
R1080 VDD.n90 VDD.n88 0.0543462
R1081 VDD.n21 VDD.n19 0.0411098
R1082 VDD.n12 VDD.n10 0.027939
R1083 VDD.n69 VDD.n66 0.0191585
R1084 VDD.n38 VDD.n37 0.018061
R1085 VDD.n110 VDD.n109 0.0175122
R1086 VDD.n93 VDD.n85 0.0153171
R1087 VDD.n56 VDD.n55 0.0147683
R1088 VDD VDD.n94 0.013122
R1089 VDD.n55 VDD.n48 0.010378
R1090 VDD.n94 VDD.n93 0.00982927
R1091 VDD.n41 VDD.n38 0.00933668
R1092 VDD.n77 VDD.n72 0.00876098
R1093 VDD.n59 VDD.n56 0.00824116
R1094 VDD.n85 VDD.n84 0.00805275
R1095 VDD.n37 VDD.n30 0.00708537
R1096 VDD.n115 VDD.n114 0.00434146
R1097 VDD.n72 VDD.n69 0.00214634
R1098 SD2_4.n11 SD2_4.n4 5.11704
R1099 SD2_4.n4 SD2_4.n1 3.44424
R1100 SD2_4.n7 SD2_4.n6 3.41802
R1101 SD2_4.n10 SD2_4.n9 3.37323
R1102 SD2_4.n4 SD2_4.n3 3.33687
R1103 SD2_4.n1 SD2_4.t3 2.7305
R1104 SD2_4.n1 SD2_4.n0 2.7305
R1105 SD2_4.n3 SD2_4.t2 2.7305
R1106 SD2_4.n3 SD2_4.n2 2.7305
R1107 SD2_4.n6 SD2_4.t7 2.7305
R1108 SD2_4.n6 SD2_4.n5 2.7305
R1109 SD2_4.n9 SD2_4.t6 2.7305
R1110 SD2_4.n9 SD2_4.n8 2.7305
R1111 SD2_4.n11 SD2_4.n10 2.2505
R1112 SD2_4.n10 SD2_4.n7 0.015125
R1113 SD2_4 SD2_4.n11 0.00261765
R1114 SD2_5 SD2_5.n10 4.78409
R1115 SD2_5.n4 SD2_5.n3 3.44212
R1116 SD2_5.n9 SD2_5.n8 3.43911
R1117 SD2_5.n15 SD2_5.n12 3.41246
R1118 SD2_5.n18 SD2_5.n17 3.41088
R1119 SD2_5.n21 SD2_5.n20 3.38757
R1120 SD2_5.n15 SD2_5.n14 3.38387
R1121 SD2_5.n4 SD2_5.n1 3.38278
R1122 SD2_5.n9 SD2_5.n6 3.38274
R1123 SD2_5.n10 SD2_5.n4 2.87871
R1124 SD2_5.n22 SD2_5.n15 2.87758
R1125 SD2_5.n12 SD2_5.t8 2.7305
R1126 SD2_5.n12 SD2_5.n11 2.7305
R1127 SD2_5.n14 SD2_5.t14 2.7305
R1128 SD2_5.n14 SD2_5.n13 2.7305
R1129 SD2_5.n6 SD2_5.t12 2.7305
R1130 SD2_5.n6 SD2_5.n5 2.7305
R1131 SD2_5.n8 SD2_5.t11 2.7305
R1132 SD2_5.n8 SD2_5.n7 2.7305
R1133 SD2_5.n1 SD2_5.t1 2.7305
R1134 SD2_5.n1 SD2_5.n0 2.7305
R1135 SD2_5.n3 SD2_5.t0 2.7305
R1136 SD2_5.n3 SD2_5.n2 2.7305
R1137 SD2_5.n17 SD2_5.t3 2.7305
R1138 SD2_5.n17 SD2_5.n16 2.7305
R1139 SD2_5.n20 SD2_5.t2 2.7305
R1140 SD2_5.n20 SD2_5.n19 2.7305
R1141 SD2_5.n10 SD2_5.n9 2.2505
R1142 SD2_5.n22 SD2_5.n21 2.2505
R1143 SD2_5.n21 SD2_5.n18 0.00543151
R1144 SD2_5 SD2_5.n22 0.00283766
R1145 OUT_4.n8 OUT_4.n7 11.6572
R1146 OUT_4.n5 OUT_4.t0 6.44473
R1147 OUT_4.n2 OUT_4.n0 6.42383
R1148 OUT_4.n2 OUT_4.n1 5.8805
R1149 OUT_4.n8 OUT_4.t5 5.8805
R1150 OUT_4.n9 OUT_4.t2 5.8805
R1151 OUT_4.n6 OUT_4.n4 5.8805
R1152 OUT_4.n7 OUT_4.n3 5.8805
R1153 OUT_4.n5 OUT_4.t3 5.8805
R1154 OUT_4 OUT_4.n9 1.88642
R1155 OUT_4.n6 OUT_4.n5 1.79955
R1156 OUT_4.n9 OUT_4.n8 0.599276
R1157 OUT_4.n7 OUT_4.n6 0.575794
R1158 OUT_4 OUT_4.n2 0.0205
R1159 SD0_2.n34 SD0_2.n33 133.643
R1160 SD0_2.n42 SD0_2.n41 48.6672
R1161 SD0_2.n69 SD0_2.n68 47.4505
R1162 SD0_2.n3 SD0_2.t53 35.1054
R1163 SD0_2.n62 SD0_2.t38 34.0104
R1164 SD0_2.n72 SD0_2.n71 21.2922
R1165 SD0_2.n63 SD0_2.n62 21.0894
R1166 SD0_2.n64 SD0_2.n63 21.0894
R1167 SD0_2.n65 SD0_2.n64 21.0894
R1168 SD0_2.n66 SD0_2.n65 21.0894
R1169 SD0_2.n67 SD0_2.n66 21.0894
R1170 SD0_2.n68 SD0_2.n67 21.0894
R1171 SD0_2.n70 SD0_2.n69 21.0894
R1172 SD0_2.n72 SD0_2.n70 21.0894
R1173 SD0_2.n44 SD0_2.n43 21.0894
R1174 SD0_2.n4 SD0_2.n3 21.0894
R1175 SD0_2.n5 SD0_2.n4 21.0894
R1176 SD0_2.n6 SD0_2.n5 21.0894
R1177 SD0_2.n7 SD0_2.n6 21.0894
R1178 SD0_2.n8 SD0_2.n7 21.0894
R1179 SD0_2.n9 SD0_2.n8 21.0894
R1180 SD0_2.n10 SD0_2.n9 21.0894
R1181 SD0_2.n11 SD0_2.n10 21.0894
R1182 SD0_2.n12 SD0_2.n11 21.0894
R1183 SD0_2.n13 SD0_2.n12 21.0894
R1184 SD0_2.n14 SD0_2.n13 21.0894
R1185 SD0_2.n15 SD0_2.n14 21.0894
R1186 SD0_2.n16 SD0_2.n15 21.0894
R1187 SD0_2.n17 SD0_2.n16 21.0894
R1188 SD0_2.n18 SD0_2.n17 21.0894
R1189 SD0_2.n19 SD0_2.n18 21.0894
R1190 SD0_2.n20 SD0_2.n19 21.0894
R1191 SD0_2.n21 SD0_2.n20 21.0894
R1192 SD0_2.n22 SD0_2.n21 21.0894
R1193 SD0_2.n23 SD0_2.n22 21.0894
R1194 SD0_2.n24 SD0_2.n23 21.0894
R1195 SD0_2.n25 SD0_2.n24 21.0894
R1196 SD0_2.n26 SD0_2.n25 21.0894
R1197 SD0_2.n27 SD0_2.n26 21.0894
R1198 SD0_2.n28 SD0_2.n27 21.0894
R1199 SD0_2.n29 SD0_2.n28 21.0894
R1200 SD0_2.n30 SD0_2.n29 21.0894
R1201 SD0_2.n31 SD0_2.n30 21.0894
R1202 SD0_2.n32 SD0_2.n31 21.0894
R1203 SD0_2.n33 SD0_2.n32 21.0894
R1204 SD0_2.n35 SD0_2.n34 21.0894
R1205 SD0_2.n36 SD0_2.n35 21.0894
R1206 SD0_2.n37 SD0_2.n36 21.0894
R1207 SD0_2.n38 SD0_2.n37 21.0894
R1208 SD0_2.n39 SD0_2.n38 21.0894
R1209 SD0_2.n40 SD0_2.n39 21.0894
R1210 SD0_2.n41 SD0_2.n40 21.0894
R1211 SD0_2.n45 SD0_2.n42 21.0894
R1212 SD0_2.n45 SD0_2.n44 21.0894
R1213 SD0_2.n3 SD0_2.t51 14.7465
R1214 SD0_2.n4 SD0_2.t64 14.7465
R1215 SD0_2.n7 SD0_2.t58 14.7465
R1216 SD0_2.n8 SD0_2.t32 14.7465
R1217 SD0_2.n11 SD0_2.t66 14.7465
R1218 SD0_2.n12 SD0_2.t41 14.7465
R1219 SD0_2.n15 SD0_2.t57 14.7465
R1220 SD0_2.n16 SD0_2.t70 14.7465
R1221 SD0_2.n19 SD0_2.t35 14.7465
R1222 SD0_2.n20 SD0_2.t68 14.7465
R1223 SD0_2.n23 SD0_2.t42 14.7465
R1224 SD0_2.n24 SD0_2.t31 14.7465
R1225 SD0_2.n27 SD0_2.t69 14.7465
R1226 SD0_2.n28 SD0_2.t44 14.7465
R1227 SD0_2.n31 SD0_2.t62 14.7465
R1228 SD0_2.n32 SD0_2.t36 14.7465
R1229 SD0_2.n62 SD0_2.t54 14.3815
R1230 SD0_2.n63 SD0_2.t29 14.3815
R1231 SD0_2.n66 SD0_2.t26 14.3815
R1232 SD0_2.n67 SD0_2.t40 14.3815
R1233 SD0_2.n70 SD0_2.t10 14.3815
R1234 SD0_2.n44 SD0_2.t20 14.3815
R1235 SD0_2.n35 SD0_2.t60 14.3815
R1236 SD0_2.n36 SD0_2.t34 14.3815
R1237 SD0_2.n39 SD0_2.t50 14.3815
R1238 SD0_2.n40 SD0_2.t72 14.3815
R1239 SD0_2.n5 SD0_2.t47 14.0165
R1240 SD0_2.n6 SD0_2.t59 14.0165
R1241 SD0_2.n9 SD0_2.t75 14.0165
R1242 SD0_2.n10 SD0_2.t28 14.0165
R1243 SD0_2.n13 SD0_2.t43 14.0165
R1244 SD0_2.n14 SD0_2.t56 14.0165
R1245 SD0_2.n17 SD0_2.t74 14.0165
R1246 SD0_2.n18 SD0_2.t49 14.0165
R1247 SD0_2.n21 SD0_2.t71 14.0165
R1248 SD0_2.n22 SD0_2.t45 14.0165
R1249 SD0_2.n25 SD0_2.t33 14.0165
R1250 SD0_2.n26 SD0_2.t73 14.0165
R1251 SD0_2.n29 SD0_2.t25 14.0165
R1252 SD0_2.n30 SD0_2.t52 14.0165
R1253 SD0_2.n33 SD0_2.t37 14.0165
R1254 SD0_2.n69 SD0_2.t16 12.9916
R1255 SD0_2.n71 SD0_2.t14 12.9916
R1256 SD0_2.n43 SD0_2.t8 12.9916
R1257 SD0_2.n64 SD0_2.t39 12.9215
R1258 SD0_2.n65 SD0_2.t65 12.9215
R1259 SD0_2.n68 SD0_2.t61 12.9215
R1260 SD0_2.n34 SD0_2.t48 12.9215
R1261 SD0_2.n37 SD0_2.t55 12.9215
R1262 SD0_2.n38 SD0_2.t67 12.9215
R1263 SD0_2.n41 SD0_2.t27 12.9215
R1264 SD0_2.n42 SD0_2.t22 12.9215
R1265 SD0_2.n74 SD0_2.t18 10.7743
R1266 SD0_2.n47 SD0_2.t12 10.7743
R1267 SD0_2.n75 SD0_2.n73 3.54502
R1268 SD0_2.n48 SD0_2.n46 3.54477
R1269 SD0_2.n75 SD0_2.n74 3.50535
R1270 SD0_2.n48 SD0_2.n47 3.50535
R1271 SD0_2.n59 SD0_2.n56 3.07598
R1272 SD0_2.n85 SD0_2.n52 3.01065
R1273 SD0_2.n54 SD0_2.n53 2.90221
R1274 SD0_2.n82 SD0_2.n81 2.90214
R1275 SD0_2.n77 SD0_2.n76 2.88451
R1276 SD0_2.n49 SD0_2.n2 2.88438
R1277 SD0_2.n61 SD0_2.n60 2.87834
R1278 SD0_2.n56 SD0_2.n55 2.87828
R1279 SD0_2.n58 SD0_2.n57 2.87828
R1280 SD0_2.n52 SD0_2.n51 2.82902
R1281 SD0_2.n50 SD0_2.n1 2.76772
R1282 SD0_2.n78 SD0_2.n61 2.75462
R1283 SD0_2.n1 SD0_2.t1 2.7305
R1284 SD0_2.n1 SD0_2.n0 2.7305
R1285 SD0_2.n90 SD0_2.t13 2.7305
R1286 SD0_2.n90 SD0_2.n89 2.7305
R1287 SD0_2.n59 SD0_2.n58 2.50797
R1288 SD0_2.n80 SD0_2.n54 2.50522
R1289 SD0_2.n52 SD0_2.t9 2.49942
R1290 SD0_2.n58 SD0_2.t3 2.43824
R1291 SD0_2.n56 SD0_2.t17 2.43824
R1292 SD0_2.n61 SD0_2.t4 2.4382
R1293 SD0_2.n82 SD0_2.t7 2.40701
R1294 SD0_2.n54 SD0_2.t19 2.40696
R1295 SD0_2.n78 SD0_2.n77 2.35277
R1296 SD0_2.n50 SD0_2.n49 2.3515
R1297 SD0_2.n84 SD0_2.n83 2.24989
R1298 SD0_2.n94 SD0_2.n93 1.50283
R1299 SD0_2.n92 SD0_2.n90 1.43792
R1300 SD0_2.n83 SD0_2.n82 1.0106
R1301 SD0_2.n46 SD0_2.n45 0.967483
R1302 SD0_2.n73 SD0_2.n72 0.96743
R1303 SD0_2.n84 SD0_2.n80 0.610728
R1304 SD0_2.n79 SD0_2.n59 0.564953
R1305 SD0_2.n87 SD0_2.n86 0.560976
R1306 SD0_2.n79 SD0_2.n78 0.141929
R1307 SD0_2.n88 SD0_2.n50 0.119429
R1308 SD0_2.n88 SD0_2.n87 0.0205
R1309 SD0_2.n86 SD0_2.n85 0.0171667
R1310 SD0_2.n80 SD0_2.n79 0.013514
R1311 SD0_2.n85 SD0_2.n84 0.0109989
R1312 SD0_2.n94 SD0_2.n88 0.00943873
R1313 SD0_2.n49 SD0_2.n48 0.0045
R1314 SD0_2.n92 SD0_2.n91 0.00371009
R1315 SD0_2 SD0_2.n94 0.00355856
R1316 SD0_2.n77 SD0_2.n75 0.0025
R1317 SD0_2.n93 SD0_2.n92 0.0017949
R1318 SD0_1.n39 SD0_1.n36 4.73161
R1319 SD0_1.n35 SD0_1.n34 3.08659
R1320 SD0_1.n42 SD0_1.n41 3.04854
R1321 SD0_1.n26 SD0_1.n11 3.04726
R1322 SD0_1.n18 SD0_1.n17 3.04688
R1323 SD0_1.n53 SD0_1.n7 3.04375
R1324 SD0_1.n44 SD0_1.n9 3.04171
R1325 SD0_1.n20 SD0_1.n13 3.03541
R1326 SD0_1.n41 SD0_1.n40 2.9021
R1327 SD0_1.n5 SD0_1.t4 2.7305
R1328 SD0_1.n5 SD0_1.n4 2.7305
R1329 SD0_1.n50 SD0_1.t29 2.7305
R1330 SD0_1.n50 SD0_1.n49 2.7305
R1331 SD0_1.n46 SD0_1.t0 2.7305
R1332 SD0_1.n46 SD0_1.n45 2.7305
R1333 SD0_1.n38 SD0_1.t25 2.7305
R1334 SD0_1.n38 SD0_1.n37 2.7305
R1335 SD0_1.n32 SD0_1.t6 2.7305
R1336 SD0_1.n32 SD0_1.n31 2.7305
R1337 SD0_1.n28 SD0_1.t23 2.7305
R1338 SD0_1.n28 SD0_1.n27 2.7305
R1339 SD0_1.n22 SD0_1.t1 2.7305
R1340 SD0_1.n22 SD0_1.n21 2.7305
R1341 SD0_1.n15 SD0_1.t20 2.7305
R1342 SD0_1.n15 SD0_1.n14 2.7305
R1343 SD0_1.n17 SD0_1.t2 2.7305
R1344 SD0_1.n17 SD0_1.n16 2.7305
R1345 SD0_1.n13 SD0_1.t21 2.7305
R1346 SD0_1.n13 SD0_1.n12 2.7305
R1347 SD0_1.n11 SD0_1.t3 2.7305
R1348 SD0_1.n11 SD0_1.n10 2.7305
R1349 SD0_1.n34 SD0_1.t30 2.7305
R1350 SD0_1.n34 SD0_1.n33 2.7305
R1351 SD0_1.n9 SD0_1.t18 2.7305
R1352 SD0_1.n9 SD0_1.n8 2.7305
R1353 SD0_1.n7 SD0_1.t7 2.7305
R1354 SD0_1.n7 SD0_1.n6 2.7305
R1355 SD0_1.n1 SD0_1.t27 2.7305
R1356 SD0_1.n1 SD0_1.n0 2.7305
R1357 SD0_1.n18 SD0_1.n15 2.56247
R1358 SD0_1.n39 SD0_1.n38 2.56221
R1359 SD0_1.n35 SD0_1.n32 2.562
R1360 SD0_1.n55 SD0_1.n5 2.55991
R1361 SD0_1.n41 SD0_1.t5 2.40706
R1362 SD0_1.n52 SD0_1.n51 1.49447
R1363 SD0_1.n24 SD0_1.n23 1.49447
R1364 SD0_1.n30 SD0_1.n29 1.49423
R1365 SD0_1.n48 SD0_1.n47 1.49423
R1366 SD0_1.n3 SD0_1.n1 1.43789
R1367 SD0_1.n51 SD0_1.n50 1.43787
R1368 SD0_1.n29 SD0_1.n28 1.43765
R1369 SD0_1.n47 SD0_1.n46 1.43732
R1370 SD0_1.n23 SD0_1.n22 1.437
R1371 SD0_1.n56 SD0_1.n3 1.12934
R1372 SD0_1.n52 SD0_1.n48 0.58072
R1373 SD0_1.n19 SD0_1.n18 0.575838
R1374 SD0_1.n25 SD0_1.n24 0.574178
R1375 SD0_1.n55 SD0_1.n54 0.566624
R1376 SD0_1.n36 SD0_1.n30 0.554675
R1377 SD0_1.n43 SD0_1.n42 0.513212
R1378 SD0_1.n56 SD0_1.n55 0.482617
R1379 SD0_1.n20 SD0_1.n19 0.0271667
R1380 SD0_1.n54 SD0_1.n53 0.0249444
R1381 SD0_1.n48 SD0_1.n44 0.0212506
R1382 SD0_1.n26 SD0_1.n25 0.0205
R1383 SD0_1.n30 SD0_1.n26 0.0201395
R1384 SD0_1.n44 SD0_1.n43 0.0193889
R1385 SD0_1.n53 SD0_1.n52 0.0153623
R1386 SD0_1.n24 SD0_1.n20 0.0134755
R1387 SD0_1.n36 SD0_1.n35 0.0132059
R1388 SD0_1 SD0_1.n56 0.00682738
R1389 SD0_1.n42 SD0_1.n39 0.00579412
R1390 SD0_1.n3 SD0_1.n2 0.00157825
R1391 OUT_5.n18 OUT_5.n17 11.1462
R1392 OUT_5.n10 OUT_5.n9 6.90515
R1393 OUT_5.n15 OUT_5.t7 6.48993
R1394 OUT_5.n18 OUT_5.t4 6.12071
R1395 OUT_5.n22 OUT_5.n0 6.11137
R1396 OUT_5.n10 OUT_5.n8 3.54767
R1397 OUT_5.n15 OUT_5.n14 3.46159
R1398 OUT_5.n19 OUT_5.n6 3.46159
R1399 OUT_5.n21 OUT_5.n2 3.46159
R1400 OUT_5.n16 OUT_5.n12 3.38137
R1401 OUT_5.n20 OUT_5.n4 3.38137
R1402 OUT_5.n12 OUT_5.t1 2.7305
R1403 OUT_5.n12 OUT_5.n11 2.7305
R1404 OUT_5.n14 OUT_5.t14 2.7305
R1405 OUT_5.n14 OUT_5.n13 2.7305
R1406 OUT_5.n8 OUT_5.t3 2.7305
R1407 OUT_5.n8 OUT_5.n7 2.7305
R1408 OUT_5.n4 OUT_5.t10 2.7305
R1409 OUT_5.n4 OUT_5.n3 2.7305
R1410 OUT_5.n6 OUT_5.t0 2.7305
R1411 OUT_5.n6 OUT_5.n5 2.7305
R1412 OUT_5.n2 OUT_5.t8 2.7305
R1413 OUT_5.n2 OUT_5.n1 2.7305
R1414 OUT_5.n17 OUT_5.n16 0.379057
R1415 OUT_5.n16 OUT_5.n15 0.379057
R1416 OUT_5.n22 OUT_5.n21 0.379057
R1417 OUT_5.n21 OUT_5.n20 0.379057
R1418 OUT_5.n20 OUT_5.n19 0.379057
R1419 OUT_5.n19 OUT_5.n18 0.370706
R1420 OUT_5 OUT_5.n22 0.136892
R1421 OUT_5.n17 OUT_5.n10 0.00235567
R1422 SD2_1 SD2_1.n20 9.24575
R1423 SD2_1 SD2_1.n9 4.5005
R1424 SD2_1 SD2_1.n9 4.5005
R1425 SD2_1.n19 SD2_1.n18 3.45039
R1426 SD2_1.n14 SD2_1.n13 3.44985
R1427 SD2_1.n9 SD2_1.n8 3.44969
R1428 SD2_1.n4 SD2_1.n3 3.44925
R1429 SD2_1.n14 SD2_1.n11 3.4367
R1430 SD2_1.n19 SD2_1.n16 3.43615
R1431 SD2_1.n4 SD2_1.n1 3.43133
R1432 SD2_1.n9 SD2_1.n6 3.43013
R1433 SD2_1.n20 SD2_1.n19 2.87896
R1434 SD2_1 SD2_1.n4 2.8298
R1435 SD2_1.n11 SD2_1.t13 2.7305
R1436 SD2_1.n11 SD2_1.n10 2.7305
R1437 SD2_1.n13 SD2_1.t12 2.7305
R1438 SD2_1.n13 SD2_1.n12 2.7305
R1439 SD2_1.n16 SD2_1.t7 2.7305
R1440 SD2_1.n16 SD2_1.n15 2.7305
R1441 SD2_1.n18 SD2_1.t4 2.7305
R1442 SD2_1.n18 SD2_1.n17 2.7305
R1443 SD2_1.n1 SD2_1.t10 2.7305
R1444 SD2_1.n1 SD2_1.n0 2.7305
R1445 SD2_1.n3 SD2_1.t9 2.7305
R1446 SD2_1.n3 SD2_1.n2 2.7305
R1447 SD2_1.n6 SD2_1.t5 2.7305
R1448 SD2_1.n6 SD2_1.n5 2.7305
R1449 SD2_1.n8 SD2_1.t6 2.7305
R1450 SD2_1.n8 SD2_1.n7 2.7305
R1451 SD2_1.n20 SD2_1.n14 2.25147
R1452 SD2_2 SD2_2.n1 3.20697
R1453 SD2_2.n1 SD2_2.t1 2.7305
R1454 SD2_2.n1 SD2_2.n0 2.7305
R1455 OUT_1 OUT_1.t0 5.96093
R1456 OUT_3.n3 OUT_3.n2 8.66766
R1457 OUT_3.n2 OUT_3.n0 6.45579
R1458 OUT_3.n4 OUT_3.t2 5.8805
R1459 OUT_3.n3 OUT_3.t1 5.8805
R1460 OUT_3.n2 OUT_3.n1 5.8805
R1461 OUT_3.n4 OUT_3.n3 0.564731
R1462 OUT_3 OUT_3.n4 0.0558846
R1463 G1_2.n20 G1_2.n16 147.578
R1464 G1_2.n39 G1_2.n35 142.844
R1465 G1_2.n34 G1_2.n33 101.016
R1466 G1_2.n38 G1_2.n37 101.016
R1467 G1_2.n19 G1_2.n18 101.016
R1468 G1_2.n15 G1_2.n14 101.016
R1469 G1_2.n33 G1_2.t32 33.5864
R1470 G1_2.n14 G1_2.t33 33.5864
R1471 G1_2.n35 G1_2.n34 20.5194
R1472 G1_2.n39 G1_2.n38 20.5194
R1473 G1_2.n37 G1_2.n36 20.5194
R1474 G1_2.n18 G1_2.n17 20.5194
R1475 G1_2.n16 G1_2.n15 20.5194
R1476 G1_2.n20 G1_2.n19 20.5194
R1477 G1_2.n33 G1_2.t30 13.0675
R1478 G1_2.n34 G1_2.t29 13.0675
R1479 G1_2.n35 G1_2.t26 13.0675
R1480 G1_2.n38 G1_2.t12 13.0675
R1481 G1_2.n37 G1_2.t20 13.0675
R1482 G1_2.n36 G1_2.t22 13.0675
R1483 G1_2.n17 G1_2.t14 13.0675
R1484 G1_2.n18 G1_2.t8 13.0675
R1485 G1_2.n19 G1_2.t18 13.0675
R1486 G1_2.n14 G1_2.t31 13.0675
R1487 G1_2.n15 G1_2.t25 13.0675
R1488 G1_2.n16 G1_2.t28 13.0675
R1489 G1_2.n30 G1_2.t10 8.3225
R1490 G1_2.n13 G1_2.t16 8.1765
R1491 G1_2.n13 G1_2.n0 8.0005
R1492 G1_2.n48 G1_2.n47 8.0005
R1493 G1_2.n9 G1_2.n7 6.51833
R1494 G1_2.n3 G1_2.t4 6.51833
R1495 G1_2.n11 G1_2.t6 5.8805
R1496 G1_2.n10 G1_2.t5 5.8805
R1497 G1_2.n9 G1_2.n8 5.8805
R1498 G1_2.n5 G1_2.n1 5.8805
R1499 G1_2.n4 G1_2.n2 5.8805
R1500 G1_2.n3 G1_2.t1 5.8805
R1501 G1_2.n12 G1_2.n11 5.81863
R1502 G1_2.n6 G1_2.n5 5.52662
R1503 G1_2.n49 G1_2.n48 4.5005
R1504 G1_2.n12 G1_2.n6 4.28996
R1505 G1_2.n21 G1_2.n0 3.53359
R1506 G1_2.n41 G1_2.n40 3.50535
R1507 G1_2.n23 G1_2.t19 3.03383
R1508 G1_2.n23 G1_2.n22 3.03383
R1509 G1_2.n27 G1_2.t21 3.03383
R1510 G1_2.n27 G1_2.n26 3.03383
R1511 G1_2.n25 G1_2.t15 3.03383
R1512 G1_2.n25 G1_2.n24 3.03383
R1513 G1_2.n29 G1_2.t11 3.03383
R1514 G1_2.n29 G1_2.n28 3.03383
R1515 G1_2.n32 G1_2.n31 2.88425
R1516 G1_2.n44 G1_2.n27 2.8392
R1517 G1_2.n45 G1_2.n25 2.8392
R1518 G1_2.n46 G1_2.n23 2.80007
R1519 G1_2.n43 G1_2.n29 2.80007
R1520 G1_2.n31 G1_2.n30 2.1905
R1521 G1_2.n10 G1_2.n9 2.07441
R1522 G1_2.n48 G1_2.n13 2.0445
R1523 G1_2.n4 G1_2.n3 2.0118
R1524 G1_2.n49 G1_2.n12 1.80063
R1525 G1_2.n45 G1_2.n44 1.59702
R1526 G1_2.n46 G1_2.n45 1.58339
R1527 G1_2.n44 G1_2.n43 1.58339
R1528 G1_2.n48 G1_2.n21 1.44681
R1529 G1_2.n21 G1_2.n20 1.15481
R1530 G1_2.n40 G1_2.n39 1.06529
R1531 G1_2.n11 G1_2.n10 0.638326
R1532 G1_2.n5 G1_2.n4 0.638326
R1533 G1_2.n47 G1_2.n46 0.0972273
R1534 G1_2.n43 G1_2.n42 0.0932273
R1535 G1_2.n42 G1_2.n41 0.0305
R1536 G1_2.n47 G1_2.n0 0.0265
R1537 G1_2 G1_2.n0 0.0085
R1538 G1_2.n41 G1_2.n32 0.0055
R1539 G1_2 G1_2.n49 0.0025
R1540 SD2_3.n3 SD2_3.n2 6.50095
R1541 SD2_3.n2 SD2_3.n0 6.4673
R1542 SD2_3 SD2_3.t0 6.15396
R1543 SD2_3.n3 SD2_3.t3 5.8805
R1544 SD2_3.n2 SD2_3.n1 5.8805
R1545 SD2_3 SD2_3.n3 0.291269
R1546 OUT_2.n1 OUT_2.t0 11.8383
R1547 OUT_2.n1 OUT_2.n0 5.8805
R1548 OUT_2 OUT_2.n1 0.068
R1549 SD1_1.n16 SD1_1.n15 7.78572
R1550 SD1_1.n10 SD1_1.n9 3.20235
R1551 SD1_1.n18 SD1_1.n17 3.17681
R1552 SD1_1.n23 SD1_1.t15 3.03383
R1553 SD1_1.n23 SD1_1.n22 3.03383
R1554 SD1_1.n20 SD1_1.t3 3.03383
R1555 SD1_1.n20 SD1_1.n19 3.03383
R1556 SD1_1.n14 SD1_1.t14 3.03383
R1557 SD1_1.n14 SD1_1.n13 3.03383
R1558 SD1_1.n6 SD1_1.t1 3.03383
R1559 SD1_1.n6 SD1_1.n5 3.03383
R1560 SD1_1.n8 SD1_1.t11 3.03383
R1561 SD1_1.n8 SD1_1.n7 3.03383
R1562 SD1_1.n1 SD1_1.t6 3.03383
R1563 SD1_1.n1 SD1_1.n0 3.03383
R1564 SD1_1.n21 SD1_1.n18 2.97146
R1565 SD1_1.n11 SD1_1.n10 2.94829
R1566 SD1_1.n11 SD1_1.n8 2.75112
R1567 SD1_1.n18 SD1_1.t8 2.69498
R1568 SD1_1.n10 SD1_1.t0 2.66057
R1569 SD1_1.n15 SD1_1.n14 2.38615
R1570 SD1_1.n24 SD1_1.n23 2.37424
R1571 SD1_1.n21 SD1_1.n20 2.37412
R1572 SD1_1.n12 SD1_1.n6 2.37207
R1573 SD1_1.n3 SD1_1.n1 1.65597
R1574 SD1_1.n16 SD1_1.n4 1.12886
R1575 SD1_1.n24 SD1_1.n21 0.626727
R1576 SD1_1.n12 SD1_1.n11 0.613463
R1577 SD1_1.n15 SD1_1.n12 0.609042
R1578 SD1_1.n25 SD1_1.n24 0.584266
R1579 SD1_1 SD1_1.n25 0.0265
R1580 SD1_1 SD1_1.n16 0.00686644
R1581 SD1_1.n4 SD1_1.n3 0.00289542
R1582 SD1_1.n3 SD1_1.n2 0.00210331
C0 OUT_4 G1_2 2.04f
C1 OUT_1 SD2_2 0.037f
C2 OUT_4 SD2_3 0.00229f
C3 SD2_5 SD2_4 0.31f
C4 OUT_3 ITAIL_1 9.92e-21
C5 OUT_3 G1_2 0.00637f
C6 OUT_4 ITAIL 0.345f
C7 G1_2 ITAIL_1 2.95f
C8 G1_1 SD0_2 0.0117f
C9 G1_1 SD1_1 0.278f
C10 SD2_5 OUT_2 0.357f
C11 OUT_3 SD2_3 0.401f
C12 OUT_4 OUT_5 3.28e-20
C13 ITAIL_1 OUT_6 0.783f
C14 OUT_3 ITAIL 0.115f
C15 OUT_4 SD2_1 0.0577f
C16 SD2_3 G1_2 8.28e-20
C17 SD2_5 G2_1 0.248f
C18 OUT_2 G1_1 0.00111f
C19 ITAIL ITAIL_1 0.0238f
C20 SD1_1 SD0_2 0.0268f
C21 G1_2 ITAIL 0.404f
C22 VDD G1_1 8.09f
C23 SD2_4 OUT_2 0.278f
C24 OUT_2 SD0_2 1.91e-19
C25 ITAIL_1 OUT_5 0.966f
C26 SD0_2 SD3_1 0.714f
C27 SD2_4 G2_1 0.162f
C28 OUT_3 SD2_1 1.03f
C29 OUT_2 SD1_1 1.34e-19
C30 SD2_3 ITAIL 0.0655f
C31 OUT_1 SD2_5 0.548f
C32 G1_1 SD0_1 0.00111f
C33 G1_2 OUT_5 0.0145f
C34 SD2_1 ITAIL_1 0.00647f
C35 VDD SD0_2 0.0482f
C36 G1_2 SD2_1 0.908f
C37 OUT_1 G1_1 2.47e-19
C38 VDD SD1_1 1.81f
C39 OUT_6 OUT_5 0.0108f
C40 SD0_2 SD0_1 0.578f
C41 OUT_2 G2_1 0.0405f
C42 OUT_1 SD2_4 0.00368f
C43 OUT_2 VDD 0.00143f
C44 SD1_1 SD0_1 0.0888f
C45 OUT_1 SD0_2 3.23e-19
C46 ITAIL SD2_1 0.159f
C47 OUT_1 SD1_1 1.66e-19
C48 SD3_1 SD0_1 0.297f
C49 OUT_1 OUT_2 0.119f
C50 VDD SD0_1 0.00435f
C51 OUT_1 G2_1 0.0181f
C52 SD2_2 ITAIL 0.00992f
C53 OUT_1 VDD 0.00414f
C54 OUT_4 SD2_5 1.05f
C55 OUT_1 SD0_1 4.34e-20
C56 OUT_4 G1_1 0.00299f
C57 SD2_5 OUT_3 0.182f
C58 OUT_4 SD2_4 0.00348f
C59 OUT_4 SD0_2 7.89e-19
C60 OUT_4 SD1_1 0.00292f
C61 SD2_5 G1_2 0.00259f
C62 OUT_3 G1_1 5.15e-21
C63 G1_1 ITAIL_1 0.378f
C64 G1_1 G1_2 2.47f
C65 OUT_3 SD2_4 0.373f
C66 OUT_4 OUT_2 0.0432f
C67 SD2_5 SD2_3 0.0442f
C68 ITAIL_1 SD0_2 4.05f
C69 OUT_3 SD1_1 3.89e-21
C70 SD2_5 ITAIL 0.265f
C71 SD2_4 G1_2 2.28e-19
C72 OUT_4 G2_1 0.246f
C73 SD1_1 ITAIL_1 2.15f
C74 OUT_4 VDD 0.00942f
C75 G1_2 SD1_1 0.643f
C76 OUT_3 OUT_2 0.00229f
C77 SD2_4 SD2_3 0.461f
C78 OUT_4 SD0_1 3e-19
C79 OUT_2 ITAIL_1 0.00111f
C80 ITAIL_1 SD3_1 1.01f
C81 SD0_2 OUT_6 1.22f
C82 SD2_4 ITAIL 0.124f
C83 OUT_3 G2_1 0.115f
C84 SD2_5 SD2_1 0.0861f
C85 OUT_2 G1_2 0.0172f
C86 OUT_1 OUT_4 0.93f
C87 OUT_3 VDD 1.31e-20
C88 G1_1 OUT_5 0.0179f
C89 G2_1 ITAIL_1 0.00126f
C90 VDD ITAIL_1 1.31f
C91 G1_2 G2_1 0.192f
C92 VDD G1_2 3.52f
C93 SD2_3 OUT_2 0.159f
C94 ITAIL_1 SD0_1 1.01f
C95 SD0_2 OUT_5 0.921f
C96 OUT_6 SD3_1 3.97f
C97 OUT_2 ITAIL 0.144f
C98 SD2_4 SD2_1 0.00249f
C99 SD2_3 G2_1 0.0979f
C100 OUT_1 OUT_3 0.0247f
C101 SD2_2 SD2_5 0.0175f
C102 SD1_1 OUT_5 0.0217f
C103 G1_2 SD0_1 5.13e-19
C104 OUT_1 ITAIL_1 0.00116f
C105 ITAIL G2_1 1.17f
C106 OUT_1 G1_2 0.0105f
C107 OUT_2 OUT_5 0.00243f
C108 OUT_6 SD0_1 0.0272f
C109 SD3_1 OUT_5 0.00851f
C110 OUT_2 SD2_1 3.54e-19
C111 OUT_1 SD2_3 0.00462f
C112 VDD OUT_5 0.0363f
C113 G2_1 SD2_1 0.212f
C114 OUT_1 ITAIL 0.149f
C115 OUT_5 SD0_1 2.11f
C116 SD2_2 OUT_2 0.00234f
C117 SD2_2 G2_1 0.0436f
C118 OUT_1 SD2_1 7.09e-19
C119 OUT_4 OUT_3 0.783f
C120 OUT_4 ITAIL_1 0.00434f
.ends

