magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1703 -1133 1703 1133
<< metal1 >>
rect -703 127 703 133
rect -703 101 -697 127
rect -671 101 -621 127
rect -595 101 -545 127
rect -519 101 -469 127
rect -443 101 -393 127
rect -367 101 -317 127
rect -291 101 -241 127
rect -215 101 -165 127
rect -139 101 -89 127
rect -63 101 -13 127
rect 13 101 63 127
rect 89 101 139 127
rect 165 101 215 127
rect 241 101 291 127
rect 317 101 367 127
rect 393 101 443 127
rect 469 101 519 127
rect 545 101 595 127
rect 621 101 671 127
rect 697 101 703 127
rect -703 51 703 101
rect -703 25 -697 51
rect -671 25 -621 51
rect -595 25 -545 51
rect -519 25 -469 51
rect -443 25 -393 51
rect -367 25 -317 51
rect -291 25 -241 51
rect -215 25 -165 51
rect -139 25 -89 51
rect -63 25 -13 51
rect 13 25 63 51
rect 89 25 139 51
rect 165 25 215 51
rect 241 25 291 51
rect 317 25 367 51
rect 393 25 443 51
rect 469 25 519 51
rect 545 25 595 51
rect 621 25 671 51
rect 697 25 703 51
rect -703 -25 703 25
rect -703 -51 -697 -25
rect -671 -51 -621 -25
rect -595 -51 -545 -25
rect -519 -51 -469 -25
rect -443 -51 -393 -25
rect -367 -51 -317 -25
rect -291 -51 -241 -25
rect -215 -51 -165 -25
rect -139 -51 -89 -25
rect -63 -51 -13 -25
rect 13 -51 63 -25
rect 89 -51 139 -25
rect 165 -51 215 -25
rect 241 -51 291 -25
rect 317 -51 367 -25
rect 393 -51 443 -25
rect 469 -51 519 -25
rect 545 -51 595 -25
rect 621 -51 671 -25
rect 697 -51 703 -25
rect -703 -101 703 -51
rect -703 -127 -697 -101
rect -671 -127 -621 -101
rect -595 -127 -545 -101
rect -519 -127 -469 -101
rect -443 -127 -393 -101
rect -367 -127 -317 -101
rect -291 -127 -241 -101
rect -215 -127 -165 -101
rect -139 -127 -89 -101
rect -63 -127 -13 -101
rect 13 -127 63 -101
rect 89 -127 139 -101
rect 165 -127 215 -101
rect 241 -127 291 -101
rect 317 -127 367 -101
rect 393 -127 443 -101
rect 469 -127 519 -101
rect 545 -127 595 -101
rect 621 -127 671 -101
rect 697 -127 703 -101
rect -703 -133 703 -127
<< via1 >>
rect -697 101 -671 127
rect -621 101 -595 127
rect -545 101 -519 127
rect -469 101 -443 127
rect -393 101 -367 127
rect -317 101 -291 127
rect -241 101 -215 127
rect -165 101 -139 127
rect -89 101 -63 127
rect -13 101 13 127
rect 63 101 89 127
rect 139 101 165 127
rect 215 101 241 127
rect 291 101 317 127
rect 367 101 393 127
rect 443 101 469 127
rect 519 101 545 127
rect 595 101 621 127
rect 671 101 697 127
rect -697 25 -671 51
rect -621 25 -595 51
rect -545 25 -519 51
rect -469 25 -443 51
rect -393 25 -367 51
rect -317 25 -291 51
rect -241 25 -215 51
rect -165 25 -139 51
rect -89 25 -63 51
rect -13 25 13 51
rect 63 25 89 51
rect 139 25 165 51
rect 215 25 241 51
rect 291 25 317 51
rect 367 25 393 51
rect 443 25 469 51
rect 519 25 545 51
rect 595 25 621 51
rect 671 25 697 51
rect -697 -51 -671 -25
rect -621 -51 -595 -25
rect -545 -51 -519 -25
rect -469 -51 -443 -25
rect -393 -51 -367 -25
rect -317 -51 -291 -25
rect -241 -51 -215 -25
rect -165 -51 -139 -25
rect -89 -51 -63 -25
rect -13 -51 13 -25
rect 63 -51 89 -25
rect 139 -51 165 -25
rect 215 -51 241 -25
rect 291 -51 317 -25
rect 367 -51 393 -25
rect 443 -51 469 -25
rect 519 -51 545 -25
rect 595 -51 621 -25
rect 671 -51 697 -25
rect -697 -127 -671 -101
rect -621 -127 -595 -101
rect -545 -127 -519 -101
rect -469 -127 -443 -101
rect -393 -127 -367 -101
rect -317 -127 -291 -101
rect -241 -127 -215 -101
rect -165 -127 -139 -101
rect -89 -127 -63 -101
rect -13 -127 13 -101
rect 63 -127 89 -101
rect 139 -127 165 -101
rect 215 -127 241 -101
rect 291 -127 317 -101
rect 367 -127 393 -101
rect 443 -127 469 -101
rect 519 -127 545 -101
rect 595 -127 621 -101
rect 671 -127 697 -101
<< metal2 >>
rect -703 127 703 133
rect -703 101 -697 127
rect -671 101 -621 127
rect -595 101 -545 127
rect -519 101 -469 127
rect -443 101 -393 127
rect -367 101 -317 127
rect -291 101 -241 127
rect -215 101 -165 127
rect -139 101 -89 127
rect -63 101 -13 127
rect 13 101 63 127
rect 89 101 139 127
rect 165 101 215 127
rect 241 101 291 127
rect 317 101 367 127
rect 393 101 443 127
rect 469 101 519 127
rect 545 101 595 127
rect 621 101 671 127
rect 697 101 703 127
rect -703 51 703 101
rect -703 25 -697 51
rect -671 25 -621 51
rect -595 25 -545 51
rect -519 25 -469 51
rect -443 25 -393 51
rect -367 25 -317 51
rect -291 25 -241 51
rect -215 25 -165 51
rect -139 25 -89 51
rect -63 25 -13 51
rect 13 25 63 51
rect 89 25 139 51
rect 165 25 215 51
rect 241 25 291 51
rect 317 25 367 51
rect 393 25 443 51
rect 469 25 519 51
rect 545 25 595 51
rect 621 25 671 51
rect 697 25 703 51
rect -703 -25 703 25
rect -703 -51 -697 -25
rect -671 -51 -621 -25
rect -595 -51 -545 -25
rect -519 -51 -469 -25
rect -443 -51 -393 -25
rect -367 -51 -317 -25
rect -291 -51 -241 -25
rect -215 -51 -165 -25
rect -139 -51 -89 -25
rect -63 -51 -13 -25
rect 13 -51 63 -25
rect 89 -51 139 -25
rect 165 -51 215 -25
rect 241 -51 291 -25
rect 317 -51 367 -25
rect 393 -51 443 -25
rect 469 -51 519 -25
rect 545 -51 595 -25
rect 621 -51 671 -25
rect 697 -51 703 -25
rect -703 -101 703 -51
rect -703 -127 -697 -101
rect -671 -127 -621 -101
rect -595 -127 -545 -101
rect -519 -127 -469 -101
rect -443 -127 -393 -101
rect -367 -127 -317 -101
rect -291 -127 -241 -101
rect -215 -127 -165 -101
rect -139 -127 -89 -101
rect -63 -127 -13 -101
rect 13 -127 63 -101
rect 89 -127 139 -101
rect 165 -127 215 -101
rect 241 -127 291 -101
rect 317 -127 367 -101
rect 393 -127 443 -101
rect 469 -127 519 -101
rect 545 -127 595 -101
rect 621 -127 671 -101
rect 697 -127 703 -101
rect -703 -133 703 -127
<< end >>
