magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2278 -14728 2278 14728
<< nwell >>
rect -278 -12728 278 12728
<< nsubdiff >>
rect -195 12623 195 12645
rect -195 -12623 -173 12623
rect 173 -12623 195 12623
rect -195 -12645 195 -12623
<< nsubdiffcont >>
rect -173 -12623 173 12623
<< metal1 >>
rect -184 12623 184 12634
rect -184 -12623 -173 12623
rect 173 -12623 184 12623
rect -184 -12634 184 -12623
<< end >>
