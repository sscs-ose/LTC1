magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -2309 -1022 989 1022
<< metal4 >>
rect -1306 14 -14 19
rect -1306 -14 -1301 14
rect -1273 -14 -1235 14
rect -1207 -14 -1169 14
rect -1141 -14 -1103 14
rect -1075 -14 -1037 14
rect -1009 -14 -971 14
rect -943 -14 -905 14
rect -877 -14 -839 14
rect -811 -14 -773 14
rect -745 -14 -707 14
rect -679 -14 -641 14
rect -613 -14 -575 14
rect -547 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 -14 14
rect -1306 -19 -14 -14
<< via4 >>
rect -1301 -14 -1273 14
rect -1235 -14 -1207 14
rect -1169 -14 -1141 14
rect -1103 -14 -1075 14
rect -1037 -14 -1009 14
rect -971 -14 -943 14
rect -905 -14 -877 14
rect -839 -14 -811 14
rect -773 -14 -745 14
rect -707 -14 -679 14
rect -641 -14 -613 14
rect -575 -14 -547 14
rect -509 -14 -481 14
rect -443 -14 -415 14
rect -377 -14 -349 14
rect -311 -14 -283 14
rect -245 -14 -217 14
rect -179 -14 -151 14
rect -113 -14 -85 14
rect -47 -14 -19 14
<< metal5 >>
rect -1309 14 -11 22
rect -1309 -14 -1301 14
rect -1273 -14 -1235 14
rect -1207 -14 -1169 14
rect -1141 -14 -1103 14
rect -1075 -14 -1037 14
rect -1009 -14 -971 14
rect -943 -14 -905 14
rect -877 -14 -839 14
rect -811 -14 -773 14
rect -745 -14 -707 14
rect -679 -14 -641 14
rect -613 -14 -575 14
rect -547 -14 -509 14
rect -481 -14 -443 14
rect -415 -14 -377 14
rect -349 -14 -311 14
rect -283 -14 -245 14
rect -217 -14 -179 14
rect -151 -14 -113 14
rect -85 -14 -47 14
rect -19 -14 -11 14
rect -1309 -22 -11 -14
<< end >>
