magic
tech gf180mcuC
magscale 1 10
timestamp 1714554054
<< nwell >>
rect -60 831 344 1012
rect 114 556 171 558
<< psubdiff >>
rect -20 141 293 156
rect -20 94 17 141
rect 250 94 293 141
rect -20 80 293 94
<< nsubdiff >>
rect 18 938 277 951
rect 18 937 217 938
rect 18 891 40 937
rect 86 892 217 937
rect 263 892 277 938
rect 86 891 277 892
rect 18 878 277 891
<< psubdiffcont >>
rect 17 94 250 141
<< nsubdiffcont >>
rect 40 891 86 937
rect 217 892 263 938
<< polysilicon >>
rect 114 556 171 558
rect 114 511 170 556
rect 75 498 170 511
rect 75 442 89 498
rect 144 442 170 498
rect 75 428 170 442
rect 114 383 170 428
<< polycontact >>
rect 89 442 144 498
<< metal1 >>
rect -61 938 344 1028
rect -61 937 217 938
rect -61 891 40 937
rect 86 892 217 937
rect 263 892 344 938
rect 86 891 344 892
rect -61 857 344 891
rect 33 612 85 857
rect 75 498 152 511
rect 75 496 89 498
rect -61 446 89 496
rect 75 442 89 446
rect 144 446 152 498
rect 199 499 248 760
rect 199 446 338 499
rect 144 442 151 446
rect 75 428 151 442
rect 20 172 84 349
rect 199 294 248 446
rect -61 141 344 172
rect -61 94 17 141
rect 250 94 344 141
rect -61 58 344 94
use nmos_3p3_DDNVWA  nmos_3p3_DDNVWA_0
timestamp 1714126980
transform 1 0 142 0 1 317
box -144 -97 144 97
use pmos_3p3_MQGBLR  pmos_3p3_MQGBLR_0
timestamp 1714474474
transform 1 0 143 0 1 682
box -202 -210 202 210
<< labels >>
flabel psubdiffcont 134 118 134 118 0 FreeSans 480 0 0 0 VSS
port 6 nsew
flabel metal1 -37 469 -37 469 0 FreeSans 320 0 0 0 IN
port 8 nsew
flabel metal1 307 471 307 471 0 FreeSans 320 0 0 0 OUT
port 9 nsew
<< end >>
