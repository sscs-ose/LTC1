* NGSPICE file created from CM_MSB.ext - technology: gf180mcuC

.subckt nmos_3p3_AGPLV7 a_n138_n60# a_50_n60# a_n50_n104# VSUBS
X0 a_50_n60# a_n50_n104# a_n138_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt nmos_3p3_AQEADK a_n138_n60# a_50_n60# a_n50_n104# VSUBS
X0 a_50_n60# a_n50_n104# a_n138_n60# VSUBS nfet_03v3 ad=0.264p pd=2.08u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt MSB_Unit_Cell_p1 m1_0_435# m1_37_n24# a_316_n447# m1_0_n631# a_316_26# a_84_242#
+ a_3095_69# VSUBS
Xnmos_3p3_AGPLV7_5 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_6 a_3095_69# m1_37_n24# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_7 m1_37_n24# a_3095_69# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_8 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_9 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_0 a_3095_69# m1_0_435# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_1 m1_37_n24# a_3095_69# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_2 a_3095_69# m1_0_435# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_30 a_3095_69# m1_37_n24# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_4 a_3095_69# m1_37_n24# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_3 m1_0_435# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_31 m1_0_435# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_20 a_3095_69# m1_37_n24# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_5 m1_37_n24# a_3095_69# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_21 m1_37_n24# a_3095_69# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_10 a_3095_69# m1_37_n24# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_6 a_3095_69# m1_0_435# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_22 a_3095_69# m1_0_435# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_11 m1_0_435# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_7 m1_0_435# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_23 m1_0_435# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_12 a_3095_69# m1_37_n24# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_8 a_3095_69# m1_37_n24# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_30 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_24 a_3095_69# m1_37_n24# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_13 m1_37_n24# a_3095_69# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_9 m1_37_n24# a_3095_69# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_31 m1_37_n24# a_3095_69# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_20 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_26 a_3095_69# m1_0_435# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_25 m1_37_n24# a_3095_69# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_15 m1_0_435# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_14 a_3095_69# m1_0_435# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_21 a_3095_69# m1_37_n24# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_10 a_3095_69# m1_37_n24# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_27 a_3095_69# m1_0_435# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_16 m1_0_435# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_22 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_23 m1_37_n24# a_3095_69# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_12 a_3095_69# m1_37_n24# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_11 m1_37_n24# a_3095_69# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_28 a_3095_69# m1_37_n24# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_17 m1_37_n24# a_3095_69# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_24 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_13 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_29 m1_37_n24# a_3095_69# a_84_242# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AQEADK_18 a_3095_69# m1_0_435# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_25 m1_37_n24# a_3095_69# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_14 m1_37_n24# a_3095_69# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AQEADK_19 m1_0_435# a_3095_69# a_316_26# VSUBS nmos_3p3_AQEADK
Xnmos_3p3_AGPLV7_26 a_3095_69# m1_37_n24# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_15 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_27 a_3095_69# m1_37_n24# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_16 a_3095_69# m1_37_n24# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_28 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_17 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_29 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_18 m1_37_n24# a_3095_69# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_19 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_0 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_1 m1_0_n631# a_3095_69# a_316_26# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_2 a_3095_69# m1_37_n24# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_3 m1_37_n24# a_3095_69# a_316_n447# VSUBS nmos_3p3_AGPLV7
Xnmos_3p3_AGPLV7_4 a_3095_69# m1_0_n631# a_316_26# VSUBS nmos_3p3_AGPLV7
.ends

.subckt CM_MSB OUT VSS IM IM_T
XMSB_Unit_Cell_p1_0 VSS OUT IM_T VSS IM IM_T m2_630_2002# VSS MSB_Unit_Cell_p1
XMSB_Unit_Cell_p1_1 VSS OUT IM_T VSS IM IM_T m2_630_2002# VSS MSB_Unit_Cell_p1
.ends

