** sch_path: /home/shahid/GF180Projects/Divider/Xschem/dec_3x8_test.sch
**.subckt dec_3x8_test
x1 IN1 VSS VDD D0 D1 D2 D3 D4 D5 D6 D7 IN3 IN2 dec_3x8
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 IN1 VSS pulse(3.3 0 0 100p 100p 200n 400n)
.save i(v3)
V4 IN2 VSS pulse(3.3 0 0 100p 100p 100n 200n)
.save i(v4)
V5 IN3 VSS pulse(3.3 0 0 100p 100p 50n 100n)
.save i(v5)
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.control
save all
tran 50p 500n
plot v(IN1) v(IN2)+3.5 v(IN3)+7 v(D0)+10.5 v(D1)+14 v(D2)+17.5 v(D3)+21 v(D4)+24.5 v(D5)+28
+ v(D6)+31.5 v(D7)+35



*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  dec_3x8.sym # of pins=13
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/dec_3x8.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/dec_3x8.sch
.subckt dec_3x8 IN1 VSS VDD D0 D1 D2 D3 D4 D5 D6 D7 IN3 IN2
x1 VSS IN1 IN1B VDD inv_my
x2 VSS IN2 IN2B VDD inv_my
x3 VSS IN3 IN3B VDD inv_my
x4 IN1B VSS VDD D0 IN2B IN3B and_3
x5 IN1B VSS VDD D0 IN2B IN3 and_3
x6 IN1B VSS VDD D0 IN2 IN3B and_3
x7 IN1B VSS VDD D0 IN2 IN3 and_3
x8 IN1 VSS VDD D0 IN2B IN3B and_3
x9 IN1 VSS VDD D0 IN2B IN3 and_3
x10 IN1 VSS VDD D0 IN2 IN3B and_3
x11 IN1 VSS VDD D0 IN2 IN3 and_3
.ends


* expanding   symbol:  inv_my.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/inv_my.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/inv_my.sch
.subckt inv_my VSS IN OUT VDD
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  and_3.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/and_3.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/and_3.sch
.subckt and_3 IN1 VSS VDD OUT IN3 IN2
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin OUT
*.ipin IN3
XM3 net2 IN3 VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=3
XM4 net1 IN1 net3 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=3
XM5 OUT net1 VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 OUT net1 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM1 net1 IN3 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM2 net1 IN1 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM7 net3 IN2 net2 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=3
XM8 net1 IN2 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
.ends

.GLOBAL GND
.end
