magic
tech gf180mcuD
magscale 1 10
timestamp 1701146377
<< error_s >>
rect -1010 61760 -821 61846
rect 3787 61760 3976 61846
rect 4206 61760 4395 61846
rect 9003 61760 9192 61846
rect -927 61743 -926 61760
rect -927 61730 -913 61743
rect -907 61730 -821 61760
rect -940 61717 -821 61730
rect -928 61697 -821 61717
rect -940 61684 -821 61697
rect -927 61671 -913 61684
rect -927 61652 -926 61671
rect -907 61652 -821 61684
rect -927 61651 -821 61652
rect 3873 61652 3874 61760
rect 3893 61743 3976 61760
rect 3879 61671 3976 61743
rect 4289 61743 4290 61760
rect 4289 61730 4303 61743
rect 4309 61730 4395 61760
rect 4276 61717 4395 61730
rect 4288 61697 4395 61717
rect 4276 61684 4395 61697
rect 3893 61652 3976 61671
rect 3873 61651 3976 61652
rect 4289 61671 4303 61684
rect 4289 61652 4290 61671
rect 4309 61652 4395 61684
rect 4289 61651 4395 61652
rect 9089 61652 9090 61760
rect 9109 61743 9192 61760
rect 9095 61671 9192 61743
rect 10266 61697 10447 61730
rect 9109 61652 9192 61671
rect 9089 61651 9192 61652
rect 10252 61644 10447 61697
rect 13690 61715 13871 61748
rect 13690 61662 13885 61715
rect 14764 61697 14945 61730
rect -1010 61548 -821 61634
rect 4206 61548 4395 61634
rect 10252 61611 10353 61644
rect -986 61440 -985 61548
rect -907 61440 -821 61548
rect -986 61439 -821 61440
rect 4230 61440 4231 61548
rect 4309 61440 4395 61548
rect 10338 61550 10339 61611
rect 10338 61537 10352 61550
rect 10361 61537 10447 61644
rect 10325 61524 10447 61537
rect 10337 61504 10447 61524
rect 10325 61491 10447 61504
rect 4230 61439 4395 61440
rect 10338 61478 10352 61491
rect 10338 61372 10339 61478
rect 10361 61372 10447 61491
rect 13776 61390 13777 61662
rect 13785 61629 13885 61662
rect 13799 61568 13885 61629
rect 14750 61644 14945 61697
rect 18188 61715 18369 61748
rect 18188 61662 18383 61715
rect 14750 61611 14851 61644
rect 13785 61496 13885 61568
rect 14836 61550 14837 61611
rect 14836 61537 14850 61550
rect 14859 61537 14945 61644
rect 14823 61524 14945 61537
rect 14835 61504 14945 61524
rect 13799 61390 13885 61496
rect 14823 61491 14945 61504
rect 13776 61389 13885 61390
rect 14836 61478 14850 61491
rect 10338 61371 10447 61372
rect 14836 61372 14837 61478
rect 14859 61372 14945 61491
rect 18274 61390 18275 61662
rect 18283 61629 18383 61662
rect 18297 61568 18383 61629
rect 18283 61496 18383 61568
rect 18297 61390 18383 61496
rect 18274 61389 18383 61390
rect 14836 61371 14945 61372
rect 10242 60442 10432 60528
rect 13705 60460 13895 60546
rect 10314 60397 10315 60442
rect 10346 60414 10432 60442
rect 13791 60432 13792 60460
rect 10314 60384 10328 60397
rect 10333 60384 10432 60414
rect 10301 60371 10432 60384
rect 10313 60351 10432 60371
rect 10301 60338 10432 60351
rect 13705 60402 13804 60432
rect 13823 60415 13895 60460
rect 14740 60442 14930 60528
rect 18203 60460 18393 60546
rect 13809 60402 13895 60415
rect 13705 60392 13895 60402
rect 13705 60356 13804 60392
rect 13705 60346 13805 60356
rect 10314 60325 10328 60338
rect 10333 60328 10432 60338
rect 10314 60288 10315 60325
rect 10346 60288 10432 60328
rect 13791 60306 13792 60346
rect 13809 60343 13895 60392
rect 14812 60397 14813 60442
rect 14844 60414 14930 60442
rect 18289 60432 18290 60460
rect 14812 60384 14826 60397
rect 14831 60384 14930 60414
rect 14799 60371 14930 60384
rect 14811 60351 14930 60371
rect 13823 60306 13895 60343
rect 14799 60338 14930 60351
rect 18203 60402 18302 60432
rect 18321 60415 18393 60460
rect 18307 60402 18393 60415
rect 18203 60392 18393 60402
rect 18203 60356 18302 60392
rect 18203 60346 18303 60356
rect 13791 60305 13895 60306
rect 14812 60325 14826 60338
rect 14831 60328 14930 60338
rect 10314 60287 10432 60288
rect 14812 60288 14813 60325
rect 14844 60288 14930 60328
rect 18289 60306 18290 60346
rect 18307 60343 18393 60392
rect 18321 60306 18393 60343
rect 18289 60305 18393 60306
rect 14812 60287 14930 60288
rect 10266 59434 10447 59467
rect 10252 59381 10447 59434
rect 13690 59452 13871 59485
rect 13690 59399 13885 59452
rect 14764 59434 14945 59467
rect 10252 59348 10353 59381
rect 10338 59287 10339 59348
rect 10338 59274 10352 59287
rect 10361 59274 10447 59381
rect 10325 59261 10447 59274
rect 10337 59241 10447 59261
rect 10325 59228 10447 59241
rect 10338 59215 10352 59228
rect 10338 59109 10339 59215
rect 10361 59109 10447 59228
rect 13776 59127 13777 59399
rect 13785 59366 13885 59399
rect 13799 59305 13885 59366
rect 14750 59381 14945 59434
rect 18188 59452 18369 59485
rect 18188 59399 18383 59452
rect 14750 59348 14851 59381
rect 13785 59233 13885 59305
rect 14836 59287 14837 59348
rect 14836 59274 14850 59287
rect 14859 59274 14945 59381
rect 14823 59261 14945 59274
rect 14835 59241 14945 59261
rect 13799 59127 13885 59233
rect 14823 59228 14945 59241
rect 13776 59126 13885 59127
rect 14836 59215 14850 59228
rect 10338 59108 10447 59109
rect 14836 59109 14837 59215
rect 14859 59109 14945 59228
rect 18274 59127 18275 59399
rect 18283 59366 18383 59399
rect 18297 59305 18383 59366
rect 18283 59233 18383 59305
rect 18297 59127 18383 59233
rect 18274 59126 18383 59127
rect 14836 59108 14945 59109
rect 10266 58202 10447 58235
rect 10252 58149 10447 58202
rect 13690 58220 13871 58253
rect 13690 58167 13885 58220
rect 14764 58202 14945 58235
rect 10252 58116 10353 58149
rect 10338 58055 10339 58116
rect 10338 58042 10352 58055
rect 10361 58042 10447 58149
rect 10325 58029 10447 58042
rect 10337 58009 10447 58029
rect 10325 57996 10447 58009
rect 10338 57983 10352 57996
rect 10338 57877 10339 57983
rect 10361 57877 10447 57996
rect 13776 57895 13777 58167
rect 13785 58134 13885 58167
rect 13799 58073 13885 58134
rect 14750 58149 14945 58202
rect 18188 58220 18369 58253
rect 18188 58167 18383 58220
rect 14750 58116 14851 58149
rect 13785 58001 13885 58073
rect 14836 58055 14837 58116
rect 14836 58042 14850 58055
rect 14859 58042 14945 58149
rect 14823 58029 14945 58042
rect 14835 58009 14945 58029
rect 13799 57895 13885 58001
rect 14823 57996 14945 58009
rect 13776 57894 13885 57895
rect 14836 57983 14850 57996
rect 10338 57876 10447 57877
rect 14836 57877 14837 57983
rect 14859 57877 14945 57996
rect 18274 57895 18275 58167
rect 18283 58134 18383 58167
rect 18297 58073 18383 58134
rect 18283 58001 18383 58073
rect 18297 57895 18383 58001
rect 18274 57894 18383 57895
rect 14836 57876 14945 57877
rect 3787 57784 3976 57870
rect 9003 57784 9192 57870
rect 3873 57676 3874 57784
rect 3893 57767 3976 57784
rect 3879 57695 3976 57767
rect 3893 57676 3976 57695
rect 3873 57675 3976 57676
rect 9089 57676 9090 57784
rect 9109 57767 9192 57784
rect 9095 57695 9192 57767
rect 9109 57676 9192 57695
rect 9089 57675 9192 57676
rect 10242 56947 10432 57033
rect 13705 56965 13895 57051
rect 10314 56902 10315 56947
rect 10346 56919 10432 56947
rect 13791 56937 13792 56965
rect 10314 56889 10328 56902
rect 10333 56889 10432 56919
rect 10301 56876 10432 56889
rect 10313 56856 10432 56876
rect 10301 56843 10432 56856
rect 13705 56907 13804 56937
rect 13823 56920 13895 56965
rect 14740 56947 14930 57033
rect 18203 56965 18393 57051
rect 13809 56907 13895 56920
rect 13705 56897 13895 56907
rect 13705 56861 13804 56897
rect 13705 56851 13805 56861
rect 10314 56830 10328 56843
rect 10333 56833 10432 56843
rect 10314 56793 10315 56830
rect 10346 56793 10432 56833
rect 13791 56811 13792 56851
rect 13809 56848 13895 56897
rect 14812 56902 14813 56947
rect 14844 56919 14930 56947
rect 18289 56937 18290 56965
rect 14812 56889 14826 56902
rect 14831 56889 14930 56919
rect 14799 56876 14930 56889
rect 14811 56856 14930 56876
rect 13823 56811 13895 56848
rect 14799 56843 14930 56856
rect 18203 56907 18302 56937
rect 18321 56920 18393 56965
rect 18307 56907 18393 56920
rect 18203 56897 18393 56907
rect 18203 56861 18302 56897
rect 18203 56851 18303 56861
rect 13791 56810 13895 56811
rect 14812 56830 14826 56843
rect 14831 56833 14930 56843
rect 10314 56792 10432 56793
rect 14812 56793 14813 56830
rect 14844 56793 14930 56833
rect 18289 56811 18290 56851
rect 18307 56848 18393 56897
rect 18321 56811 18393 56848
rect 18289 56810 18393 56811
rect 14812 56792 14930 56793
rect 10266 55939 10447 55972
rect 10252 55886 10447 55939
rect 13690 55957 13871 55990
rect 13690 55904 13885 55957
rect 14764 55939 14945 55972
rect 10252 55853 10353 55886
rect 10338 55792 10339 55853
rect 10338 55779 10352 55792
rect 10361 55779 10447 55886
rect 10325 55766 10447 55779
rect 10337 55746 10447 55766
rect 10325 55733 10447 55746
rect 10338 55720 10352 55733
rect 10338 55614 10339 55720
rect 10361 55614 10447 55733
rect 13776 55632 13777 55904
rect 13785 55871 13885 55904
rect 13799 55810 13885 55871
rect 14750 55886 14945 55939
rect 18188 55957 18369 55990
rect 18188 55904 18383 55957
rect 14750 55853 14851 55886
rect 13785 55738 13885 55810
rect 14836 55792 14837 55853
rect 14836 55779 14850 55792
rect 14859 55779 14945 55886
rect 14823 55766 14945 55779
rect 14835 55746 14945 55766
rect 13799 55632 13885 55738
rect 14823 55733 14945 55746
rect 13776 55631 13885 55632
rect 14836 55720 14850 55733
rect 10338 55613 10447 55614
rect 14836 55614 14837 55720
rect 14859 55614 14945 55733
rect 18274 55632 18275 55904
rect 18283 55871 18383 55904
rect 18297 55810 18383 55871
rect 18283 55738 18383 55810
rect 18297 55632 18383 55738
rect 18274 55631 18383 55632
rect 14836 55613 14945 55614
rect 13690 54733 13871 54766
rect 18188 54733 18369 54766
rect 13690 54680 13885 54733
rect 18188 54680 18383 54733
rect 10266 54613 10447 54646
rect 10252 54560 10447 54613
rect 10252 54527 10353 54560
rect 10338 54466 10339 54527
rect 10338 54453 10352 54466
rect 10361 54453 10447 54560
rect 10325 54440 10447 54453
rect 10337 54420 10447 54440
rect 10325 54407 10447 54420
rect 13776 54408 13777 54680
rect 13785 54647 13885 54680
rect 13799 54586 13885 54647
rect 14764 54613 14945 54646
rect 13785 54514 13885 54586
rect 14750 54560 14945 54613
rect 14750 54527 14851 54560
rect 13799 54408 13885 54514
rect 14836 54466 14837 54527
rect 14836 54453 14850 54466
rect 14859 54453 14945 54560
rect 14823 54440 14945 54453
rect 14835 54420 14945 54440
rect 13776 54407 13885 54408
rect 14823 54407 14945 54420
rect 18274 54408 18275 54680
rect 18283 54647 18383 54680
rect 18297 54586 18383 54647
rect 18283 54514 18383 54586
rect 18297 54408 18383 54514
rect 18274 54407 18383 54408
rect 10338 54394 10352 54407
rect 10338 54288 10339 54394
rect 10361 54288 10447 54407
rect 10338 54287 10447 54288
rect 14836 54394 14850 54407
rect 14836 54288 14837 54394
rect 14859 54288 14945 54407
rect 14836 54287 14945 54288
rect 13705 53478 13895 53564
rect 18203 53478 18393 53564
rect 13791 53450 13792 53478
rect 10242 53358 10432 53444
rect 13705 53420 13804 53450
rect 13823 53433 13895 53478
rect 18289 53450 18290 53478
rect 13809 53420 13895 53433
rect 13705 53410 13895 53420
rect 13705 53374 13804 53410
rect 13705 53364 13805 53374
rect 10314 53313 10315 53358
rect 10346 53330 10432 53358
rect 10314 53300 10328 53313
rect 10333 53300 10432 53330
rect 13791 53324 13792 53364
rect 13809 53361 13895 53410
rect 13823 53324 13895 53361
rect 14740 53358 14930 53444
rect 18203 53420 18302 53450
rect 18321 53433 18393 53478
rect 18307 53420 18393 53433
rect 18203 53410 18393 53420
rect 18203 53374 18302 53410
rect 18203 53364 18303 53374
rect 13791 53323 13895 53324
rect 14812 53313 14813 53358
rect 14844 53330 14930 53358
rect 14812 53300 14826 53313
rect 14831 53300 14930 53330
rect 18289 53324 18290 53364
rect 18307 53361 18393 53410
rect 18321 53324 18393 53361
rect 18289 53323 18393 53324
rect 10301 53287 10432 53300
rect 14799 53287 14930 53300
rect 10313 53267 10432 53287
rect 14811 53267 14930 53287
rect 10301 53254 10432 53267
rect 14799 53254 14930 53267
rect 10314 53241 10328 53254
rect 10333 53244 10432 53254
rect 10314 53204 10315 53241
rect 10346 53204 10432 53244
rect 10314 53203 10432 53204
rect 14812 53241 14826 53254
rect 14831 53244 14930 53254
rect 14812 53204 14813 53241
rect 14844 53204 14930 53244
rect 14812 53203 14930 53204
rect 13690 52470 13871 52503
rect 18188 52470 18369 52503
rect 13690 52417 13885 52470
rect 18188 52417 18383 52470
rect 10266 52350 10447 52383
rect 10252 52297 10447 52350
rect -1011 52205 -822 52291
rect 4206 52205 4395 52291
rect 10252 52264 10353 52297
rect -928 52185 -927 52205
rect -928 52172 -914 52185
rect -908 52172 -822 52205
rect 4289 52185 4290 52205
rect 4289 52172 4303 52185
rect 4309 52172 4395 52205
rect 10338 52203 10339 52264
rect 10338 52190 10352 52203
rect 10361 52190 10447 52297
rect 10325 52177 10447 52190
rect -941 52159 -822 52172
rect 4276 52159 4395 52172
rect -929 52139 -822 52159
rect 4288 52139 4395 52159
rect 10337 52157 10447 52177
rect 10325 52144 10447 52157
rect 13776 52145 13777 52417
rect 13785 52384 13885 52417
rect 13799 52323 13885 52384
rect 14764 52350 14945 52383
rect 13785 52251 13885 52323
rect 14750 52297 14945 52350
rect 14750 52264 14851 52297
rect 13799 52145 13885 52251
rect 14836 52203 14837 52264
rect 14836 52190 14850 52203
rect 14859 52190 14945 52297
rect 14823 52177 14945 52190
rect 14835 52157 14945 52177
rect 13776 52144 13885 52145
rect 14823 52144 14945 52157
rect 18274 52145 18275 52417
rect 18283 52384 18383 52417
rect 18297 52323 18383 52384
rect 18283 52251 18383 52323
rect 18297 52145 18383 52251
rect 18274 52144 18383 52145
rect -941 52126 -822 52139
rect 4276 52126 4395 52139
rect -928 52113 -914 52126
rect -928 52097 -927 52113
rect -908 52097 -822 52126
rect -928 52096 -822 52097
rect 4289 52113 4303 52126
rect 4289 52097 4290 52113
rect 4309 52097 4395 52126
rect 4289 52096 4395 52097
rect 10338 52131 10352 52144
rect 10338 52025 10339 52131
rect 10361 52025 10447 52144
rect 10338 52024 10447 52025
rect 14836 52131 14850 52144
rect 14836 52025 14837 52131
rect 14859 52025 14945 52144
rect 14836 52024 14945 52025
rect 13690 51082 13871 51115
rect 18188 51082 18369 51115
rect 13690 51029 13885 51082
rect 18188 51029 18383 51082
rect 10042 50733 10233 50819
rect 13776 50757 13777 51029
rect 13785 50996 13885 51029
rect 13799 50935 13885 50996
rect 13785 50863 13885 50935
rect 13799 50757 13885 50863
rect 13776 50756 13885 50757
rect 14540 50733 14731 50819
rect 18274 50757 18275 51029
rect 18283 50996 18383 51029
rect 18297 50935 18383 50996
rect 18283 50863 18383 50935
rect 18297 50757 18383 50863
rect 18274 50756 18383 50757
rect 10093 50692 10094 50733
rect 10093 50679 10107 50692
rect 10087 50666 10140 50679
rect 10092 50646 10140 50666
rect 10087 50633 10140 50646
rect 10093 50620 10107 50633
rect 10093 50589 10094 50620
rect 10147 50589 10233 50733
rect 14591 50692 14592 50733
rect 14591 50679 14605 50692
rect 14585 50666 14638 50679
rect 14590 50646 14638 50666
rect 14585 50633 14638 50646
rect 10093 50588 10233 50589
rect 14591 50620 14605 50633
rect 14591 50589 14592 50620
rect 14645 50589 14731 50733
rect 14591 50588 14731 50589
rect 13705 49827 13895 49913
rect 18203 49827 18393 49913
rect 13791 49799 13792 49827
rect 13705 49769 13804 49799
rect 13823 49782 13895 49827
rect 18289 49799 18290 49827
rect 13809 49769 13895 49782
rect 13705 49759 13895 49769
rect 13705 49723 13804 49759
rect 13705 49713 13805 49723
rect 13791 49673 13792 49713
rect 13809 49710 13895 49759
rect 18203 49769 18302 49799
rect 18321 49782 18393 49827
rect 18307 49769 18393 49782
rect 18203 49759 18393 49769
rect 18203 49723 18302 49759
rect 18203 49713 18303 49723
rect 13823 49673 13895 49710
rect 13791 49672 13895 49673
rect 18289 49673 18290 49713
rect 18307 49710 18393 49759
rect 18321 49673 18393 49710
rect 18289 49672 18393 49673
rect 13690 48819 13871 48852
rect 18188 48819 18369 48852
rect 13690 48766 13885 48819
rect 18188 48766 18383 48819
rect 10042 48672 10233 48758
rect 10093 48631 10094 48672
rect 10093 48618 10107 48631
rect 10087 48605 10140 48618
rect 10092 48585 10140 48605
rect 10087 48572 10140 48585
rect 10093 48559 10107 48572
rect 10093 48528 10094 48559
rect 10147 48528 10233 48672
rect 10093 48527 10233 48528
rect 3786 48441 3975 48527
rect 9003 48441 9192 48527
rect 13776 48494 13777 48766
rect 13785 48733 13885 48766
rect 13799 48672 13885 48733
rect 14540 48672 14731 48758
rect 13785 48600 13885 48672
rect 14591 48631 14592 48672
rect 14591 48618 14605 48631
rect 14585 48605 14638 48618
rect 13799 48494 13885 48600
rect 14590 48585 14638 48605
rect 14585 48572 14638 48585
rect 14591 48559 14605 48572
rect 14591 48528 14592 48559
rect 14645 48528 14731 48672
rect 14591 48527 14731 48528
rect 13776 48493 13885 48494
rect 18274 48494 18275 48766
rect 18283 48733 18383 48766
rect 18297 48672 18383 48733
rect 18283 48600 18383 48672
rect 18297 48494 18383 48600
rect 18274 48493 18383 48494
rect 3872 48333 3873 48441
rect 3951 48333 3975 48441
rect 3872 48332 3975 48333
rect 9089 48333 9090 48441
rect 9168 48333 9192 48441
rect 9089 48332 9192 48333
rect -1011 48229 -822 48315
rect 3786 48229 3975 48315
rect 4206 48229 4395 48315
rect 9003 48229 9192 48315
rect -928 48209 -927 48229
rect -928 48196 -914 48209
rect -908 48196 -822 48229
rect -941 48183 -822 48196
rect -929 48163 -822 48183
rect -941 48150 -822 48163
rect -928 48137 -914 48150
rect -928 48121 -927 48137
rect -908 48121 -822 48150
rect -928 48120 -822 48121
rect 3872 48121 3873 48229
rect 3892 48209 3975 48229
rect 3878 48137 3975 48209
rect 4289 48209 4290 48229
rect 4289 48196 4303 48209
rect 4309 48196 4395 48229
rect 4276 48183 4395 48196
rect 4288 48163 4395 48183
rect 4276 48150 4395 48163
rect 3892 48121 3975 48137
rect 3872 48120 3975 48121
rect 4289 48137 4303 48150
rect 4289 48121 4290 48137
rect 4309 48121 4395 48150
rect 4289 48120 4395 48121
rect 9089 48121 9090 48229
rect 9109 48209 9192 48229
rect 9095 48137 9192 48209
rect 9109 48121 9192 48137
rect 9089 48120 9192 48121
rect -1011 47104 -822 47190
rect 3786 47104 3975 47190
rect 4206 47104 4395 47190
rect 9003 47104 9192 47190
rect -928 47087 -927 47104
rect -928 47074 -914 47087
rect -908 47074 -822 47104
rect -941 47061 -822 47074
rect -929 47041 -822 47061
rect -941 47028 -822 47041
rect -928 47015 -914 47028
rect -928 46996 -927 47015
rect -908 46996 -822 47028
rect -928 46995 -822 46996
rect 3872 46996 3873 47104
rect 3892 47087 3975 47104
rect 3878 47015 3975 47087
rect 4289 47087 4290 47104
rect 4289 47074 4303 47087
rect 4309 47074 4395 47104
rect 4276 47061 4395 47074
rect 4288 47041 4395 47061
rect 4276 47028 4395 47041
rect 3892 46996 3975 47015
rect 3872 46995 3975 46996
rect 4289 47015 4303 47028
rect 4289 46996 4290 47015
rect 4309 46996 4395 47028
rect 4289 46995 4395 46996
rect 9089 46996 9090 47104
rect 9109 47087 9192 47104
rect 9095 47015 9192 47087
rect 9109 46996 9192 47015
rect 9089 46995 9192 46996
rect 3786 46892 3975 46978
rect 9003 46892 9192 46978
rect 3872 46860 3975 46892
rect 3872 46814 3888 46860
rect 3951 46814 3975 46860
rect 3872 46800 3975 46814
rect 3872 46791 3950 46800
rect 3951 46791 3975 46800
rect 3872 46783 3975 46791
rect 9089 46784 9090 46892
rect 9168 46784 9192 46892
rect 10065 46815 10246 46848
rect 14559 46815 14740 46848
rect 9089 46783 9192 46784
rect 10051 46762 10246 46815
rect 10051 46729 10152 46762
rect 10137 46668 10138 46729
rect 10137 46655 10151 46668
rect 10160 46655 10246 46762
rect 14545 46762 14740 46815
rect 14545 46729 14646 46762
rect 14631 46668 14632 46729
rect 14631 46655 14645 46668
rect 14654 46655 14740 46762
rect 10124 46642 10246 46655
rect 14618 46642 14740 46655
rect 10136 46622 10246 46642
rect 14630 46622 14740 46642
rect 10124 46609 10246 46622
rect 14618 46609 14740 46622
rect 10137 46596 10151 46609
rect 10137 46490 10138 46596
rect 10160 46490 10246 46609
rect 10137 46489 10246 46490
rect 14631 46596 14645 46609
rect 14631 46490 14632 46596
rect 14654 46490 14740 46609
rect 14631 46489 14740 46490
rect 10065 45731 10246 45764
rect 14559 45731 14740 45764
rect 10051 45678 10246 45731
rect 10051 45645 10152 45678
rect 10137 45584 10138 45645
rect 10137 45571 10151 45584
rect 10160 45571 10246 45678
rect 14545 45678 14740 45731
rect 14545 45645 14646 45678
rect 14631 45584 14632 45645
rect 14631 45571 14645 45584
rect 14654 45571 14740 45678
rect 10124 45558 10246 45571
rect 14618 45558 14740 45571
rect 10136 45538 10246 45558
rect 14630 45538 14740 45558
rect 10124 45525 10246 45538
rect 14618 45525 14740 45538
rect 10137 45512 10151 45525
rect 10137 45406 10138 45512
rect 10160 45406 10246 45525
rect 10137 45405 10246 45406
rect 14631 45512 14645 45525
rect 14631 45406 14632 45512
rect 14654 45406 14740 45525
rect 14631 45405 14740 45406
rect 12191 44714 12386 44800
rect 16685 44714 16880 44800
rect 12277 44442 12278 44714
rect 12300 44607 12386 44714
rect 12286 44535 12386 44607
rect 12300 44475 12386 44535
rect 12286 44474 12386 44475
rect 12286 44442 12372 44474
rect 12277 44441 12372 44442
rect 16771 44442 16772 44714
rect 16794 44607 16880 44714
rect 16780 44535 16880 44607
rect 16794 44475 16880 44535
rect 16780 44474 16880 44475
rect 16780 44442 16866 44474
rect 16771 44441 16866 44442
rect 18188 44251 18369 44284
rect 18188 44198 18383 44251
rect 18274 43926 18275 44198
rect 18283 44165 18383 44198
rect 18297 44104 18383 44165
rect 18283 44032 18383 44104
rect 18297 43926 18383 44032
rect 18274 43925 18383 43926
rect 10065 43780 10246 43813
rect 14559 43780 14740 43813
rect 10051 43727 10246 43780
rect 10051 43694 10152 43727
rect 10137 43633 10138 43694
rect 10137 43620 10151 43633
rect 10160 43620 10246 43727
rect 12199 43649 12394 43735
rect 14545 43727 14740 43780
rect 14545 43694 14646 43727
rect 10124 43607 10246 43620
rect 10136 43587 10246 43607
rect 10124 43574 10246 43587
rect 10137 43561 10151 43574
rect 10137 43455 10138 43561
rect 10160 43455 10246 43574
rect 10137 43454 10246 43455
rect 12285 43377 12286 43649
rect 12308 43542 12394 43649
rect 14631 43633 14632 43694
rect 14631 43620 14645 43633
rect 14654 43620 14740 43727
rect 16693 43649 16888 43735
rect 14618 43607 14740 43620
rect 14630 43587 14740 43607
rect 14618 43574 14740 43587
rect 12294 43470 12394 43542
rect 12308 43410 12394 43470
rect 14631 43561 14645 43574
rect 14631 43455 14632 43561
rect 14654 43455 14740 43574
rect 14631 43454 14740 43455
rect 12294 43409 12394 43410
rect 12294 43377 12380 43409
rect 12285 43376 12380 43377
rect 16779 43377 16780 43649
rect 16802 43542 16888 43649
rect 16788 43470 16888 43542
rect 16802 43410 16888 43470
rect 16788 43409 16888 43410
rect 16788 43377 16874 43409
rect 16779 43376 16874 43377
rect -1011 43128 -822 43214
rect 4206 43128 4395 43214
rect -928 43111 -927 43128
rect -928 43098 -914 43111
rect -908 43098 -822 43128
rect 4289 43111 4290 43128
rect 4289 43098 4303 43111
rect 4309 43098 4395 43128
rect -941 43085 -822 43098
rect 4276 43085 4395 43098
rect -929 43065 -822 43085
rect 4288 43065 4395 43085
rect -941 43052 -822 43065
rect 4276 43052 4395 43065
rect -928 43039 -914 43052
rect -928 43020 -927 43039
rect -908 43020 -822 43052
rect -928 43019 -822 43020
rect 4289 43039 4303 43052
rect 4289 43020 4290 43039
rect 4309 43020 4395 43052
rect 4289 43019 4395 43020
rect 10066 42517 10247 42550
rect 14560 42517 14741 42550
rect 10052 42464 10247 42517
rect 10052 42431 10153 42464
rect 10138 42370 10139 42431
rect 10138 42357 10152 42370
rect 10161 42357 10247 42464
rect 14546 42464 14741 42517
rect 14546 42431 14647 42464
rect 14632 42370 14633 42431
rect 14632 42357 14646 42370
rect 14655 42357 14741 42464
rect 10125 42344 10247 42357
rect 14619 42344 14741 42357
rect 10137 42324 10247 42344
rect 14631 42324 14741 42344
rect 10125 42311 10247 42324
rect 14619 42311 14741 42324
rect 10138 42298 10152 42311
rect 10138 42192 10139 42298
rect 10161 42192 10247 42311
rect 10138 42191 10247 42192
rect 14632 42298 14646 42311
rect 14632 42192 14633 42298
rect 14655 42192 14741 42311
rect 14632 42191 14741 42192
rect 12191 41500 12386 41586
rect 16685 41500 16880 41586
rect 12277 41228 12278 41500
rect 12300 41393 12386 41500
rect 12286 41321 12386 41393
rect 12300 41261 12386 41321
rect 12286 41260 12386 41261
rect 12286 41228 12372 41260
rect 12277 41227 12372 41228
rect 16771 41228 16772 41500
rect 16794 41393 16880 41500
rect 16780 41321 16880 41393
rect 16794 41261 16880 41321
rect 16780 41260 16880 41261
rect 16780 41228 16866 41260
rect 16771 41227 16866 41228
rect 10058 40517 10239 40550
rect 14552 40517 14733 40550
rect 10044 40464 10239 40517
rect 10044 40431 10145 40464
rect 10130 40370 10131 40431
rect 10130 40357 10144 40370
rect 10153 40357 10239 40464
rect 12199 40392 12394 40478
rect 14538 40464 14733 40517
rect 14538 40431 14639 40464
rect 10117 40344 10239 40357
rect 10129 40324 10239 40344
rect 10117 40311 10239 40324
rect 10130 40298 10144 40311
rect 10130 40192 10131 40298
rect 10153 40192 10239 40311
rect 10130 40191 10239 40192
rect 12285 40120 12286 40392
rect 12308 40285 12394 40392
rect 14624 40370 14625 40431
rect 14624 40357 14638 40370
rect 14647 40357 14733 40464
rect 16693 40392 16888 40478
rect 14611 40344 14733 40357
rect 14623 40324 14733 40344
rect 14611 40311 14733 40324
rect 12294 40213 12394 40285
rect 12308 40153 12394 40213
rect 14624 40298 14638 40311
rect 14624 40192 14625 40298
rect 14647 40192 14733 40311
rect 14624 40191 14733 40192
rect 12294 40152 12394 40153
rect 12294 40120 12380 40152
rect 12285 40119 12380 40120
rect 16779 40120 16780 40392
rect 16802 40285 16888 40392
rect 16788 40213 16888 40285
rect 16802 40153 16888 40213
rect 16788 40152 16888 40153
rect 16788 40120 16874 40152
rect 16779 40119 16874 40120
rect 3786 39355 3975 39441
rect 3872 39216 3873 39355
rect 3921 39269 3933 39315
rect 3934 39216 3975 39355
rect 3872 39215 3975 39216
rect 10058 38465 10239 38498
rect 10044 38412 10239 38465
rect 10044 38379 10145 38412
rect 10130 38318 10131 38379
rect 10130 38305 10144 38318
rect 10153 38305 10239 38412
rect 10117 38292 10239 38305
rect 10129 38272 10239 38292
rect 10117 38259 10239 38272
rect 10130 38246 10144 38259
rect 10130 38140 10131 38246
rect 10153 38140 10239 38259
rect 10130 38139 10239 38140
rect 50 38040 241 38126
rect 101 37999 102 38040
rect 101 37986 115 37999
rect 95 37973 148 37986
rect 100 37953 148 37973
rect 95 37940 148 37953
rect 101 37927 115 37940
rect 101 37896 102 37927
rect 155 37896 241 38040
rect 101 37895 241 37896
rect -1393 37797 -1202 37883
rect -1341 37778 -1340 37797
rect -1341 37765 -1327 37778
rect -1353 37752 -1294 37765
rect -1342 37732 -1294 37752
rect -1353 37719 -1294 37732
rect -1341 37706 -1327 37719
rect -1341 37682 -1340 37706
rect -1288 37682 -1202 37797
rect -1341 37681 -1202 37682
rect 9003 37358 9192 37444
rect 10058 37381 10239 37414
rect 9089 37250 9090 37358
rect 9109 37338 9192 37358
rect 9095 37266 9192 37338
rect 10044 37328 10239 37381
rect 10044 37295 10145 37328
rect 9109 37250 9192 37266
rect 9089 37249 9192 37250
rect 10130 37234 10131 37295
rect 10130 37221 10144 37234
rect 10153 37221 10239 37328
rect 14560 37277 14741 37310
rect 10117 37208 10239 37221
rect 10129 37188 10239 37208
rect 14546 37224 14741 37277
rect 14546 37191 14647 37224
rect 10117 37175 10239 37188
rect 10130 37162 10144 37175
rect 10130 37056 10131 37162
rect 10153 37056 10239 37175
rect 14632 37130 14633 37191
rect 14632 37117 14646 37130
rect 14655 37117 14741 37224
rect 14619 37104 14741 37117
rect 14631 37084 14741 37104
rect 14619 37071 14741 37084
rect 10130 37055 10239 37056
rect 14632 37058 14646 37071
rect 14632 36952 14633 37058
rect 14655 36952 14741 37071
rect 14632 36951 14741 36952
rect 12184 36364 12379 36450
rect 1636 36329 1817 36362
rect 73 36292 254 36325
rect 59 36239 254 36292
rect 1622 36276 1817 36329
rect 1622 36243 1723 36276
rect 59 36206 160 36239
rect 145 36145 146 36206
rect 145 36132 159 36145
rect 168 36132 254 36239
rect 1708 36182 1709 36243
rect 1708 36169 1722 36182
rect 1731 36169 1817 36276
rect 1695 36156 1817 36169
rect 1707 36136 1817 36156
rect 132 36119 254 36132
rect 1695 36123 1817 36136
rect 144 36099 254 36119
rect 132 36086 254 36099
rect 145 36073 159 36086
rect 145 35967 146 36073
rect 168 35967 254 36086
rect 1708 36110 1722 36123
rect 1708 36004 1709 36110
rect 1731 36004 1817 36123
rect 12270 36092 12271 36364
rect 12293 36257 12379 36364
rect 12279 36185 12379 36257
rect 14560 36193 14741 36226
rect 12293 36125 12379 36185
rect 12279 36124 12379 36125
rect 14546 36140 14741 36193
rect 12279 36092 12365 36124
rect 14546 36107 14647 36140
rect 12270 36091 12365 36092
rect 14632 36046 14633 36107
rect 14632 36033 14646 36046
rect 14655 36033 14741 36140
rect 14619 36020 14741 36033
rect 1708 36003 1817 36004
rect 14631 36000 14741 36020
rect 14619 35987 14741 36000
rect 145 35966 254 35967
rect 14632 35974 14646 35987
rect 14632 35868 14633 35974
rect 14655 35868 14741 35987
rect 14632 35867 14741 35868
rect 10058 35430 10239 35463
rect 10044 35377 10239 35430
rect 10044 35344 10145 35377
rect 10130 35283 10131 35344
rect 1636 35245 1817 35278
rect 10130 35270 10144 35283
rect 10153 35270 10239 35377
rect 12192 35299 12387 35385
rect 10117 35257 10239 35270
rect 1622 35192 1817 35245
rect 10129 35237 10239 35257
rect 10117 35224 10239 35237
rect 1622 35159 1723 35192
rect 1708 35098 1709 35159
rect 1708 35085 1722 35098
rect 1731 35085 1817 35192
rect 10130 35211 10144 35224
rect 10130 35105 10131 35211
rect 10153 35105 10239 35224
rect 10130 35104 10239 35105
rect 1695 35072 1817 35085
rect 1707 35052 1817 35072
rect 1695 35039 1817 35052
rect 1708 35026 1722 35039
rect 1708 34920 1709 35026
rect 1731 34920 1817 35039
rect 12278 35027 12279 35299
rect 12301 35192 12387 35299
rect 12287 35120 12387 35192
rect 16686 35176 16881 35262
rect 12301 35060 12387 35120
rect 12287 35059 12387 35060
rect 12287 35027 12373 35059
rect 12278 35026 12373 35027
rect 1708 34919 1817 34920
rect 16772 34904 16773 35176
rect 16795 35069 16881 35176
rect 16781 34997 16881 35069
rect 16795 34937 16881 34997
rect 16781 34936 16881 34937
rect 16781 34904 16867 34936
rect 16772 34903 16867 34904
rect 3762 34228 3957 34314
rect 14560 34242 14741 34275
rect 3848 33956 3849 34228
rect 3871 34121 3957 34228
rect 10059 34167 10240 34200
rect 3857 34049 3957 34121
rect 10045 34114 10240 34167
rect 14546 34189 14741 34242
rect 14546 34156 14647 34189
rect 10045 34081 10146 34114
rect 3871 33989 3957 34049
rect 10131 34020 10132 34081
rect 10131 34007 10145 34020
rect 10154 34007 10240 34114
rect 14632 34095 14633 34156
rect 14632 34082 14646 34095
rect 14655 34082 14741 34189
rect 16694 34111 16889 34197
rect 14619 34069 14741 34082
rect 14631 34049 14741 34069
rect 14619 34036 14741 34049
rect 10118 33994 10240 34007
rect 3857 33988 3957 33989
rect 3857 33956 3943 33988
rect 10130 33974 10240 33994
rect 10118 33961 10240 33974
rect 3848 33955 3943 33956
rect 10131 33948 10145 33961
rect 10131 33842 10132 33948
rect 10154 33842 10240 33961
rect 14632 34023 14646 34036
rect 14632 33917 14633 34023
rect 14655 33917 14741 34036
rect 14632 33916 14741 33917
rect 10131 33841 10240 33842
rect 16780 33839 16781 34111
rect 16803 34004 16889 34111
rect 16789 33932 16889 34004
rect 16803 33872 16889 33932
rect 16789 33871 16889 33872
rect 16789 33839 16875 33871
rect 16780 33838 16875 33839
rect 4206 33594 4395 33680
rect 4230 33486 4231 33594
rect 4309 33486 4395 33594
rect 4230 33485 4395 33486
rect 4206 33382 4395 33468
rect 9003 33382 9192 33468
rect 4289 33362 4290 33382
rect 4289 33349 4303 33362
rect 4309 33349 4395 33382
rect 4276 33336 4395 33349
rect 1636 33294 1817 33327
rect 4288 33316 4395 33336
rect 4276 33303 4395 33316
rect 1622 33241 1817 33294
rect 4289 33290 4303 33303
rect 4289 33274 4290 33290
rect 4309 33274 4395 33303
rect 4289 33273 4395 33274
rect 9089 33274 9090 33382
rect 9109 33362 9192 33382
rect 9095 33290 9192 33362
rect 9109 33274 9192 33290
rect 9089 33273 9192 33274
rect -249 33152 -56 33238
rect 1622 33208 1723 33241
rect -222 33026 -221 33152
rect -142 33026 -56 33152
rect 1708 33147 1709 33208
rect 1708 33134 1722 33147
rect 1731 33134 1817 33241
rect 3770 33163 3965 33249
rect 1695 33121 1817 33134
rect 1707 33101 1817 33121
rect 1695 33088 1817 33101
rect -222 33025 -56 33026
rect 1708 33075 1722 33088
rect 1708 32969 1709 33075
rect 1731 32969 1817 33088
rect 1708 32968 1817 32969
rect 3856 32891 3857 33163
rect 3879 33056 3965 33163
rect 12184 33150 12379 33236
rect 3865 32984 3965 33056
rect 3879 32924 3965 32984
rect 3865 32923 3965 32924
rect 3865 32891 3951 32923
rect 3856 32890 3951 32891
rect 12270 32878 12271 33150
rect 12293 33043 12379 33150
rect 12279 32971 12379 33043
rect 14561 32979 14742 33012
rect 12293 32911 12379 32971
rect 12279 32910 12379 32911
rect 14547 32926 14742 32979
rect 12279 32878 12365 32910
rect 14547 32893 14648 32926
rect 12270 32877 12365 32878
rect 14633 32832 14634 32893
rect 14633 32819 14647 32832
rect 14656 32819 14742 32926
rect 14620 32806 14742 32819
rect 14632 32786 14742 32806
rect 14620 32773 14742 32786
rect 14633 32760 14647 32773
rect 14633 32654 14634 32760
rect 14656 32654 14742 32773
rect 14633 32653 14742 32654
rect 10051 32167 10232 32200
rect 10037 32114 10232 32167
rect 10037 32081 10138 32114
rect 1637 32031 1818 32064
rect 1623 31978 1818 32031
rect 10123 32020 10124 32081
rect 10123 32007 10137 32020
rect 10146 32007 10232 32114
rect 12192 32042 12387 32128
rect 10110 31994 10232 32007
rect 1623 31945 1724 31978
rect 1709 31884 1710 31945
rect 1709 31871 1723 31884
rect 1732 31871 1818 31978
rect 10122 31974 10232 31994
rect 10110 31961 10232 31974
rect 1696 31858 1818 31871
rect 1708 31838 1818 31858
rect 10123 31948 10137 31961
rect 10123 31842 10124 31948
rect 10146 31842 10232 31961
rect 10123 31841 10232 31842
rect 1696 31825 1818 31838
rect 1709 31812 1723 31825
rect 1709 31706 1710 31812
rect 1732 31706 1818 31825
rect 12278 31770 12279 32042
rect 12301 31935 12387 32042
rect 16686 31962 16881 32048
rect 12287 31863 12387 31935
rect 12301 31803 12387 31863
rect 12287 31802 12387 31803
rect 12287 31770 12373 31802
rect 12278 31769 12373 31770
rect 1709 31705 1818 31706
rect 16772 31690 16773 31962
rect 16795 31855 16881 31962
rect 16781 31783 16881 31855
rect 16795 31723 16881 31783
rect 16781 31722 16881 31723
rect 16781 31690 16867 31722
rect 16772 31689 16867 31690
rect 6567 31362 6748 31395
rect 6553 31309 6748 31362
rect 6553 31276 6654 31309
rect 6639 31215 6640 31276
rect 6639 31202 6653 31215
rect 6662 31202 6748 31309
rect 6626 31189 6748 31202
rect 6638 31169 6748 31189
rect 6626 31156 6748 31169
rect 6639 31143 6653 31156
rect 3762 31014 3957 31100
rect 6639 31037 6640 31143
rect 6662 31037 6748 31156
rect 6639 31036 6748 31037
rect 3848 30742 3849 31014
rect 3871 30907 3957 31014
rect 14553 30979 14734 31012
rect 3857 30835 3957 30907
rect 14539 30926 14734 30979
rect 14539 30893 14640 30926
rect 3871 30775 3957 30835
rect 14625 30832 14626 30893
rect 14625 30819 14639 30832
rect 14648 30819 14734 30926
rect 16694 30854 16889 30940
rect 14612 30806 14734 30819
rect 14624 30786 14734 30806
rect 3857 30774 3957 30775
rect 3857 30742 3943 30774
rect 14612 30773 14734 30786
rect 3848 30741 3943 30742
rect 14625 30760 14639 30773
rect 14625 30654 14626 30760
rect 14648 30654 14734 30773
rect 14625 30653 14734 30654
rect 16780 30582 16781 30854
rect 16803 30747 16889 30854
rect 16789 30675 16889 30747
rect 16803 30615 16889 30675
rect 16789 30614 16889 30615
rect 16789 30582 16875 30614
rect 16780 30581 16875 30582
rect 10027 30353 10216 30439
rect 10110 30336 10111 30353
rect 10110 30323 10124 30336
rect 10130 30323 10216 30353
rect 6567 30278 6748 30311
rect 10097 30310 10216 30323
rect 10109 30290 10216 30310
rect 6553 30225 6748 30278
rect 10097 30277 10216 30290
rect 10110 30264 10124 30277
rect 10110 30245 10111 30264
rect 10130 30245 10216 30277
rect 10110 30244 10216 30245
rect 6553 30192 6654 30225
rect 6639 30131 6640 30192
rect 6639 30118 6653 30131
rect 6662 30118 6748 30225
rect 6626 30105 6748 30118
rect 6638 30085 6748 30105
rect 6626 30072 6748 30085
rect 1629 30031 1810 30064
rect 1615 29978 1810 30031
rect 6639 30059 6653 30072
rect 1615 29945 1716 29978
rect 1701 29884 1702 29945
rect 1701 29871 1715 29884
rect 1724 29871 1810 29978
rect 3770 29906 3965 29992
rect 6639 29953 6640 30059
rect 6662 29953 6748 30072
rect 6639 29952 6748 29953
rect 1688 29858 1810 29871
rect 1700 29838 1810 29858
rect 1688 29825 1810 29838
rect 1701 29812 1715 29825
rect 1701 29706 1702 29812
rect 1724 29706 1810 29825
rect 1701 29705 1810 29706
rect 3856 29634 3857 29906
rect 3879 29799 3965 29906
rect 3865 29727 3965 29799
rect 3879 29667 3965 29727
rect 3865 29666 3965 29667
rect 3865 29634 3951 29666
rect 3856 29633 3951 29634
rect 8693 29261 8888 29347
rect 8779 28989 8780 29261
rect 8802 29154 8888 29261
rect 8788 29082 8888 29154
rect 8802 29022 8888 29082
rect 8788 29021 8888 29022
rect 8788 28989 8874 29021
rect 8779 28988 8874 28989
rect 6567 28327 6748 28360
rect 6553 28274 6748 28327
rect 6553 28241 6654 28274
rect 6639 28180 6640 28241
rect 6639 28167 6653 28180
rect 6662 28167 6748 28274
rect 8701 28196 8896 28282
rect 6626 28154 6748 28167
rect 6638 28134 6748 28154
rect 6626 28121 6748 28134
rect 6639 28108 6653 28121
rect 6639 28002 6640 28108
rect 6662 28002 6748 28121
rect 6639 28001 6748 28002
rect 8787 27924 8788 28196
rect 8810 28089 8896 28196
rect 8796 28017 8896 28089
rect 8810 27957 8896 28017
rect 8796 27956 8896 27957
rect 8796 27924 8882 27956
rect 8787 27923 8882 27924
rect 1792 27775 2141 27829
rect 1558 27773 2196 27775
rect 1878 27740 1879 27773
rect 1930 27760 2002 27773
rect 1943 27742 1989 27752
rect 2055 27740 2141 27773
rect 1878 27739 2141 27740
rect 1878 27731 1965 27739
rect 6568 27064 6749 27097
rect 6554 27011 6749 27064
rect 6554 26978 6655 27011
rect 6640 26917 6641 26978
rect 6640 26904 6654 26917
rect 6663 26904 6749 27011
rect 6627 26891 6749 26904
rect 6639 26871 6749 26891
rect 6627 26858 6749 26871
rect 6640 26845 6654 26858
rect 6640 26739 6641 26845
rect 6663 26739 6749 26858
rect 6640 26738 6749 26739
rect 8693 26047 8888 26133
rect 8779 25775 8780 26047
rect 8802 25940 8888 26047
rect 8788 25868 8888 25940
rect 8802 25808 8888 25868
rect 8788 25807 8888 25808
rect 8788 25775 8874 25807
rect 8779 25774 8874 25775
rect 6560 25064 6741 25097
rect 6546 25011 6741 25064
rect 6546 24978 6647 25011
rect 6632 24917 6633 24978
rect 6632 24904 6646 24917
rect 6655 24904 6741 25011
rect 8701 24939 8896 25025
rect 6619 24891 6741 24904
rect 6631 24871 6741 24891
rect 6619 24858 6741 24871
rect 6632 24845 6646 24858
rect 6632 24739 6633 24845
rect 6655 24739 6741 24858
rect 6632 24738 6741 24739
rect 8787 24667 8788 24939
rect 8810 24832 8896 24939
rect 8796 24760 8896 24832
rect 8810 24700 8896 24760
rect 8796 24699 8896 24700
rect 8796 24667 8882 24699
rect 8787 24666 8882 24667
rect 67978 12810 73842 12820
rect 7959 11559 8308 11613
rect 7725 11557 8363 11559
rect 8045 11524 8046 11557
rect 8097 11544 8169 11557
rect 8110 11526 8156 11536
rect 8222 11524 8308 11557
rect 8045 11523 8308 11524
rect 8045 11515 8132 11523
rect 18773 11428 18774 11457
rect 21502 11426 21503 11455
rect 36908 11056 36909 11085
rect 39637 11054 39638 11083
rect 27703 10341 27704 10370
rect 30432 10343 30433 10372
rect 53190 9051 53539 9105
rect 61151 9058 61500 9112
rect 61096 9056 61734 9058
rect 53135 9049 53773 9051
rect 53276 9016 53277 9049
rect 53329 9036 53401 9049
rect 53342 9018 53388 9028
rect 53276 9015 53452 9016
rect 53453 9015 53539 9049
rect 61237 9023 61238 9056
rect 61290 9043 61362 9056
rect 61303 9025 61349 9035
rect 61237 9022 61413 9023
rect 61414 9022 61500 9056
rect 53452 9007 53539 9015
rect 61413 9014 61500 9022
rect 18731 8871 18732 8900
rect 21460 8873 21461 8902
rect 27646 7335 27647 7364
rect 30375 7337 30376 7366
rect 9138 6922 9487 6976
rect 67978 6966 67988 12810
rect 73832 6966 73842 12810
rect 67978 6956 73842 6966
rect 74592 12810 80456 12820
rect 74592 6966 74602 12810
rect 80446 6966 80456 12810
rect 74592 6956 80456 6966
rect 81206 12810 87070 12820
rect 81206 6966 81216 12810
rect 87060 6966 87070 12810
rect 81206 6956 87070 6966
rect 9036 6920 9542 6922
rect 9224 6887 9225 6920
rect 9276 6907 9348 6920
rect 9289 6889 9335 6899
rect 9401 6887 9487 6920
rect 9224 6886 9487 6887
rect 9224 6878 9311 6886
rect 67978 6450 73842 6460
rect 42986 5835 42987 5864
rect 45715 5837 45716 5866
rect 53370 4374 53719 4428
rect 53315 4372 53953 4374
rect 53456 4339 53457 4372
rect 53509 4359 53581 4372
rect 53522 4341 53568 4351
rect 53456 4338 53632 4339
rect 53633 4338 53719 4372
rect 53632 4330 53719 4338
rect 34091 2146 34189 2147
rect 45273 1478 45274 1507
rect 42102 1439 42103 1468
rect 29971 1366 30069 1367
rect 67978 606 67988 6450
rect 73832 606 73842 6450
rect 67978 596 73842 606
rect 74592 6450 80456 6460
rect 74592 606 74602 6450
rect 80446 606 80456 6450
rect 74592 596 80456 606
rect 81206 6450 87070 6460
rect 81206 606 81216 6450
rect 87060 606 87070 6450
rect 91847 4018 92196 4072
rect 91613 4016 92251 4018
rect 91933 3983 91934 4016
rect 91985 4003 92057 4016
rect 91998 3985 92044 3995
rect 92110 3983 92196 4016
rect 91933 3982 92196 3983
rect 91933 3974 92020 3982
rect 81206 596 87070 606
rect 42102 -40 42103 -11
rect 45273 -19 45274 10
rect 17203 -2071 17204 -2042
rect 19932 -2069 19933 -2040
rect 30726 -5935 31014 -5884
rect 81876 -5915 82164 -5864
rect 81552 -5917 82164 -5915
rect 30402 -5937 31014 -5935
rect 30812 -5988 30813 -5937
rect 30831 -5950 30903 -5937
rect 30928 -5988 31014 -5937
rect 81962 -5968 81963 -5917
rect 81981 -5930 82053 -5917
rect 82078 -5968 82164 -5917
rect 81962 -5969 82164 -5968
rect 30812 -5989 31014 -5988
rect 6763 -6291 7256 -6267
rect 6763 -6349 7044 -6291
rect 7061 -6349 7062 -6291
rect 6698 -6351 7093 -6349
rect 6849 -6369 6850 -6351
rect 6866 -6364 6938 -6351
rect 6958 -6369 7044 -6351
rect 6849 -6370 7044 -6369
rect 7061 -6369 7062 -6351
rect 7170 -6369 7256 -6291
rect 16318 -6348 16599 -6266
rect 20294 -6348 20575 -6266
rect 21419 -6348 21700 -6266
rect 25395 -6348 25676 -6266
rect 57913 -6271 58406 -6247
rect 57913 -6329 58194 -6271
rect 58211 -6329 58212 -6271
rect 57848 -6331 58243 -6329
rect 15886 -6350 17952 -6348
rect 19862 -6350 20780 -6348
rect 21214 -6350 22132 -6348
rect 24042 -6350 26108 -6348
rect 57999 -6349 58000 -6331
rect 58016 -6344 58088 -6331
rect 58108 -6349 58194 -6331
rect 57999 -6350 58194 -6349
rect 58211 -6349 58212 -6331
rect 58320 -6349 58406 -6271
rect 67468 -6328 67749 -6246
rect 71444 -6328 71725 -6246
rect 72569 -6328 72850 -6246
rect 76545 -6328 76826 -6246
rect 67036 -6330 69102 -6328
rect 71012 -6330 71930 -6328
rect 72364 -6330 73282 -6328
rect 75192 -6330 77258 -6328
rect 67554 -6348 67555 -6330
rect 67574 -6343 67646 -6330
rect 67663 -6348 67749 -6330
rect 67554 -6349 67749 -6348
rect 71530 -6348 71531 -6330
rect 71550 -6343 71622 -6330
rect 71639 -6348 71725 -6330
rect 71530 -6349 71725 -6348
rect 72655 -6348 72656 -6330
rect 72672 -6343 72744 -6330
rect 72764 -6348 72850 -6330
rect 72655 -6349 72850 -6348
rect 76631 -6348 76632 -6330
rect 76648 -6343 76720 -6330
rect 76740 -6348 76826 -6330
rect 76631 -6349 76826 -6348
rect 58211 -6350 58406 -6349
rect 16404 -6368 16405 -6350
rect 16424 -6363 16496 -6350
rect 16513 -6368 16599 -6350
rect 16404 -6369 16599 -6368
rect 20380 -6368 20381 -6350
rect 20400 -6363 20472 -6350
rect 20489 -6368 20575 -6350
rect 20380 -6369 20575 -6368
rect 21505 -6368 21506 -6350
rect 21522 -6363 21594 -6350
rect 21614 -6368 21700 -6350
rect 21505 -6369 21700 -6368
rect 25481 -6368 25482 -6350
rect 25498 -6363 25570 -6350
rect 25590 -6368 25676 -6350
rect 25481 -6369 25676 -6368
rect 7061 -6370 7256 -6369
rect 35371 -7055 35670 -7028
rect 86521 -7035 86820 -7008
rect 35457 -7134 35458 -7055
rect 35584 -7134 35670 -7055
rect 86607 -7114 86608 -7035
rect 86734 -7114 86820 -7035
rect 86607 -7115 86820 -7114
rect 35457 -7135 35670 -7134
rect 30483 -7377 30800 -7327
rect 32317 -7350 32729 -7336
rect 30218 -7379 31328 -7377
rect 30569 -7431 30570 -7379
rect 30610 -7392 30682 -7379
rect 30714 -7431 30800 -7379
rect 32284 -7421 32729 -7350
rect 81633 -7357 81950 -7307
rect 83467 -7330 83879 -7316
rect 81368 -7359 82478 -7357
rect 81719 -7411 81720 -7359
rect 81760 -7372 81832 -7359
rect 81864 -7411 81950 -7359
rect 83434 -7401 83879 -7330
rect 83348 -7403 84156 -7401
rect 81719 -7412 81950 -7411
rect 83434 -7416 83554 -7403
rect 83614 -7416 83686 -7403
rect 32198 -7423 33006 -7421
rect 30569 -7432 30800 -7431
rect 32284 -7436 32404 -7423
rect 32464 -7436 32536 -7423
rect 32370 -7444 32371 -7436
rect 32643 -7444 32729 -7423
rect 83520 -7424 83521 -7416
rect 83793 -7424 83879 -7403
rect 83520 -7425 83879 -7424
rect 32370 -7445 32729 -7444
rect 32280 -8913 32692 -8899
rect 33364 -8913 33776 -8899
rect 35315 -8913 35727 -8899
rect 32247 -8984 32692 -8913
rect 33331 -8984 33776 -8913
rect 35282 -8984 35727 -8913
rect 36578 -8914 36990 -8900
rect 38578 -8906 38990 -8892
rect 83430 -8893 83842 -8879
rect 84514 -8893 84926 -8879
rect 86465 -8893 86877 -8879
rect 36545 -8977 36990 -8914
rect 38545 -8977 38990 -8906
rect 83397 -8964 83842 -8893
rect 84481 -8964 84926 -8893
rect 86432 -8964 86877 -8893
rect 87728 -8894 88140 -8880
rect 89728 -8886 90140 -8872
rect 87695 -8957 88140 -8894
rect 89695 -8957 90140 -8886
rect 87695 -8959 90364 -8957
rect 83227 -8966 85203 -8964
rect 86189 -8966 87154 -8964
rect 87695 -8965 88140 -8959
rect 36545 -8979 39214 -8977
rect 83397 -8979 83517 -8966
rect 83577 -8979 83649 -8966
rect 32077 -8986 34053 -8984
rect 35039 -8986 36004 -8984
rect 36545 -8985 36990 -8979
rect 32247 -8999 32367 -8986
rect 32427 -8999 32499 -8986
rect 32333 -9007 32334 -8999
rect 32606 -9007 32692 -8986
rect 33331 -8999 33451 -8986
rect 33511 -8999 33583 -8986
rect 32333 -9008 32692 -9007
rect 33417 -9007 33418 -8999
rect 33690 -9007 33776 -8986
rect 35282 -8999 35402 -8986
rect 35462 -8999 35534 -8986
rect 33417 -9008 33776 -9007
rect 35368 -9007 35369 -8999
rect 35641 -9007 35727 -8986
rect 36302 -8987 37267 -8985
rect 36545 -9000 36665 -8987
rect 36725 -9000 36797 -8987
rect 35368 -9008 35727 -9007
rect 36631 -9008 36632 -9000
rect 36904 -9008 36990 -8987
rect 38545 -8992 38665 -8979
rect 38725 -8992 38797 -8979
rect 38631 -9000 38632 -8992
rect 38904 -9000 38990 -8979
rect 83483 -8987 83484 -8979
rect 83756 -8987 83842 -8966
rect 84481 -8979 84601 -8966
rect 84661 -8979 84733 -8966
rect 83483 -8988 83842 -8987
rect 84567 -8987 84568 -8979
rect 84840 -8987 84926 -8966
rect 86432 -8979 86552 -8966
rect 86612 -8979 86684 -8966
rect 84567 -8988 84926 -8987
rect 86518 -8987 86519 -8979
rect 86791 -8987 86877 -8966
rect 87452 -8967 88417 -8965
rect 87695 -8980 87815 -8967
rect 87875 -8980 87947 -8967
rect 86518 -8988 86877 -8987
rect 87781 -8988 87782 -8980
rect 88054 -8988 88140 -8967
rect 89695 -8972 89815 -8959
rect 89875 -8972 89947 -8959
rect 89781 -8980 89782 -8972
rect 90054 -8980 90140 -8959
rect 89781 -8981 90140 -8980
rect 87781 -8989 88140 -8988
rect 38631 -9001 38990 -9000
rect 36631 -9009 36990 -9008
rect 51854 -11027 52027 -11019
rect 6763 -11150 7044 -11064
rect 10739 -11150 11020 -11064
rect 20082 -11149 20575 -11063
rect 21419 -11149 21809 -11063
rect 21818 -11149 21912 -11063
rect 29168 -11149 29480 -11063
rect 34295 -11125 34740 -11039
rect 34381 -11147 34382 -11125
rect 34501 -11134 34547 -11125
rect 34654 -11133 34740 -11125
rect 35360 -11133 35805 -11047
rect 37509 -11125 37954 -11039
rect 34621 -11134 34740 -11133
rect 34488 -11147 34560 -11134
rect 34621 -11147 34707 -11134
rect 34018 -11149 34983 -11147
rect 6849 -11169 6850 -11150
rect 6879 -11156 6925 -11150
rect 6866 -11169 6938 -11156
rect 6958 -11169 7044 -11150
rect 10825 -11169 10826 -11150
rect 10855 -11156 10901 -11150
rect 10842 -11169 10914 -11156
rect 10934 -11169 11020 -11150
rect 6558 -11170 7044 -11169
rect 6558 -11171 6984 -11170
rect 9386 -11171 11452 -11169
rect 6879 -11183 6892 -11171
rect 6912 -11183 6925 -11171
rect 10855 -11183 10868 -11171
rect 10888 -11183 10901 -11171
rect 20168 -11227 20169 -11149
rect 20277 -11168 20363 -11149
rect 20380 -11168 20381 -11149
rect 20413 -11155 20459 -11149
rect 20400 -11168 20472 -11155
rect 20489 -11168 20575 -11149
rect 21505 -11168 21506 -11149
rect 21535 -11155 21581 -11149
rect 21522 -11168 21594 -11155
rect 21614 -11168 21700 -11149
rect 21717 -11165 21818 -11149
rect 21717 -11168 21749 -11165
rect 20245 -11170 20640 -11168
rect 21354 -11170 21749 -11168
rect 20277 -11227 20363 -11170
rect 20413 -11182 20426 -11170
rect 20446 -11182 20459 -11170
rect 21535 -11182 21548 -11170
rect 21568 -11182 21581 -11170
rect 20168 -11228 20363 -11227
rect 21717 -11211 21749 -11170
rect 21809 -11211 21818 -11165
rect 21717 -11227 21818 -11211
rect 21826 -11227 21912 -11149
rect 29254 -11210 29255 -11149
rect 29294 -11210 29340 -11198
rect 29394 -11210 29480 -11149
rect 34501 -11161 34514 -11149
rect 34534 -11155 34547 -11149
rect 35446 -11155 35447 -11133
rect 35566 -11142 35612 -11133
rect 35719 -11141 35805 -11133
rect 35686 -11142 35805 -11141
rect 35553 -11155 35625 -11142
rect 35686 -11155 35772 -11142
rect 37595 -11147 37596 -11125
rect 37715 -11134 37761 -11125
rect 37868 -11133 37954 -11125
rect 38617 -11133 39062 -11047
rect 51678 -11113 52027 -11027
rect 37835 -11134 37954 -11133
rect 37702 -11147 37774 -11134
rect 37835 -11147 37921 -11134
rect 38703 -11147 38704 -11133
rect 38823 -11142 38869 -11133
rect 38976 -11141 39062 -11133
rect 38943 -11142 39062 -11141
rect 38810 -11147 38882 -11142
rect 37232 -11149 38882 -11147
rect 37715 -11155 37728 -11149
rect 34534 -11157 37728 -11155
rect 34534 -11161 34547 -11157
rect 35566 -11169 35579 -11157
rect 35599 -11169 35612 -11157
rect 37715 -11161 37728 -11157
rect 37748 -11155 37761 -11149
rect 38703 -11155 38704 -11149
rect 38810 -11155 38882 -11149
rect 38943 -11155 39029 -11142
rect 51764 -11147 51765 -11113
rect 51830 -11134 51876 -11113
rect 51817 -11147 51889 -11134
rect 51941 -11147 52027 -11113
rect 57913 -11130 58194 -11044
rect 61889 -11130 62170 -11044
rect 71232 -11129 71725 -11043
rect 72569 -11129 72959 -11043
rect 72968 -11129 73062 -11043
rect 80318 -11129 80630 -11043
rect 85445 -11105 85890 -11019
rect 85531 -11127 85532 -11105
rect 85651 -11114 85697 -11105
rect 85804 -11113 85890 -11105
rect 86510 -11113 86955 -11027
rect 88659 -11105 89104 -11019
rect 85771 -11114 85890 -11113
rect 85638 -11127 85710 -11114
rect 85771 -11127 85857 -11114
rect 85168 -11129 86133 -11127
rect 51623 -11149 52261 -11147
rect 57999 -11149 58000 -11130
rect 58029 -11136 58075 -11130
rect 58016 -11149 58088 -11136
rect 58108 -11149 58194 -11130
rect 61975 -11149 61976 -11130
rect 62005 -11136 62051 -11130
rect 61992 -11149 62064 -11136
rect 62084 -11149 62170 -11130
rect 37748 -11157 39220 -11155
rect 37748 -11161 37761 -11157
rect 38823 -11169 38836 -11157
rect 38856 -11169 38869 -11157
rect 51830 -11161 51843 -11149
rect 51863 -11161 51876 -11149
rect 57708 -11150 58194 -11149
rect 57708 -11151 58134 -11150
rect 60536 -11151 62602 -11149
rect 58029 -11163 58042 -11151
rect 58062 -11163 58075 -11151
rect 62005 -11163 62018 -11151
rect 62038 -11163 62051 -11151
rect 71318 -11207 71319 -11129
rect 71427 -11148 71513 -11129
rect 71530 -11148 71531 -11129
rect 71563 -11135 71609 -11129
rect 71550 -11148 71622 -11135
rect 71639 -11148 71725 -11129
rect 72655 -11148 72656 -11129
rect 72685 -11135 72731 -11129
rect 72672 -11148 72744 -11135
rect 72764 -11148 72850 -11129
rect 72867 -11145 72968 -11129
rect 72867 -11148 72899 -11145
rect 71395 -11150 71790 -11148
rect 72504 -11150 72899 -11148
rect 71427 -11207 71513 -11150
rect 71563 -11162 71576 -11150
rect 71596 -11162 71609 -11150
rect 72685 -11162 72698 -11150
rect 72718 -11162 72731 -11150
rect 71318 -11208 71513 -11207
rect 72867 -11191 72899 -11150
rect 72959 -11191 72968 -11145
rect 72867 -11207 72968 -11191
rect 72976 -11207 73062 -11129
rect 80404 -11190 80405 -11129
rect 80444 -11190 80490 -11178
rect 80544 -11190 80630 -11129
rect 85651 -11141 85664 -11129
rect 85684 -11135 85697 -11129
rect 86596 -11135 86597 -11113
rect 86716 -11122 86762 -11113
rect 86869 -11121 86955 -11113
rect 86836 -11122 86955 -11121
rect 86703 -11135 86775 -11122
rect 86836 -11135 86922 -11122
rect 88745 -11127 88746 -11105
rect 88865 -11114 88911 -11105
rect 89018 -11113 89104 -11105
rect 89767 -11113 90212 -11027
rect 88985 -11114 89104 -11113
rect 88852 -11127 88924 -11114
rect 88985 -11127 89071 -11114
rect 89853 -11127 89854 -11113
rect 89973 -11122 90019 -11113
rect 90126 -11121 90212 -11113
rect 90093 -11122 90212 -11121
rect 89960 -11127 90032 -11122
rect 88382 -11129 90032 -11127
rect 88865 -11135 88878 -11129
rect 85684 -11137 88878 -11135
rect 85684 -11141 85697 -11137
rect 86716 -11149 86729 -11137
rect 86749 -11149 86762 -11137
rect 88865 -11141 88878 -11137
rect 88898 -11135 88911 -11129
rect 89853 -11135 89854 -11129
rect 89960 -11135 90032 -11129
rect 90093 -11135 90179 -11122
rect 88898 -11137 90370 -11135
rect 88898 -11141 88911 -11137
rect 89973 -11149 89986 -11137
rect 90006 -11149 90019 -11137
rect 80404 -11191 80630 -11190
rect 72867 -11208 73062 -11207
rect 29254 -11211 29480 -11210
rect 21717 -11228 21912 -11227
rect 6763 -11507 7256 -11483
rect 6763 -11565 7044 -11507
rect 6698 -11566 7044 -11565
rect 7061 -11566 7062 -11507
rect 6698 -11567 7093 -11566
rect 6849 -11585 6850 -11567
rect 6866 -11580 6938 -11567
rect 6958 -11585 7044 -11567
rect 6849 -11586 7044 -11585
rect 7061 -11585 7062 -11567
rect 7170 -11585 7256 -11507
rect 16318 -11565 16599 -11483
rect 20294 -11565 20575 -11483
rect 21419 -11565 21700 -11483
rect 25395 -11565 25676 -11483
rect 34929 -11507 35422 -11483
rect 15886 -11567 17952 -11565
rect 19862 -11567 20780 -11565
rect 21214 -11567 22132 -11565
rect 24042 -11567 26108 -11565
rect 7061 -11586 7256 -11585
rect 16404 -11585 16405 -11567
rect 16424 -11580 16496 -11567
rect 16513 -11585 16599 -11567
rect 16404 -11586 16599 -11585
rect 20380 -11585 20381 -11567
rect 20400 -11580 20472 -11567
rect 20489 -11585 20575 -11567
rect 20380 -11586 20575 -11585
rect 21505 -11585 21506 -11567
rect 21522 -11580 21594 -11567
rect 21614 -11585 21700 -11567
rect 21505 -11586 21700 -11585
rect 25481 -11585 25482 -11567
rect 25498 -11580 25570 -11567
rect 25590 -11585 25676 -11567
rect 25481 -11586 25676 -11585
rect 35015 -11585 35016 -11507
rect 35124 -11565 35422 -11507
rect 57913 -11487 58406 -11463
rect 57913 -11545 58194 -11487
rect 57848 -11546 58194 -11545
rect 58211 -11546 58212 -11487
rect 57848 -11547 58243 -11546
rect 57999 -11565 58000 -11547
rect 58016 -11560 58088 -11547
rect 58108 -11565 58194 -11547
rect 35092 -11567 35487 -11565
rect 57999 -11566 58194 -11565
rect 58211 -11565 58212 -11547
rect 58320 -11565 58406 -11487
rect 67468 -11545 67749 -11463
rect 71444 -11545 71725 -11463
rect 72569 -11545 72850 -11463
rect 76545 -11545 76826 -11463
rect 86079 -11487 86572 -11463
rect 67036 -11547 69102 -11545
rect 71012 -11547 71930 -11545
rect 72364 -11547 73282 -11545
rect 75192 -11547 77258 -11545
rect 58211 -11566 58406 -11565
rect 67554 -11565 67555 -11547
rect 67574 -11560 67646 -11547
rect 67663 -11565 67749 -11547
rect 67554 -11566 67749 -11565
rect 71530 -11565 71531 -11547
rect 71550 -11560 71622 -11547
rect 71639 -11565 71725 -11547
rect 71530 -11566 71725 -11565
rect 72655 -11565 72656 -11547
rect 72672 -11560 72744 -11547
rect 72764 -11565 72850 -11547
rect 72655 -11566 72850 -11565
rect 76631 -11565 76632 -11547
rect 76648 -11560 76720 -11547
rect 76740 -11565 76826 -11547
rect 76631 -11566 76826 -11565
rect 86165 -11565 86166 -11487
rect 86274 -11545 86572 -11487
rect 86242 -11547 86637 -11545
rect 86274 -11565 86360 -11547
rect 86165 -11566 86360 -11565
rect 86377 -11565 86378 -11547
rect 86397 -11560 86469 -11547
rect 86486 -11565 86572 -11547
rect 86377 -11566 86572 -11565
rect 35124 -11585 35210 -11567
rect 35015 -11586 35210 -11585
rect 35227 -11585 35228 -11567
rect 35247 -11580 35319 -11567
rect 35336 -11585 35422 -11567
rect 35227 -11586 35422 -11585
rect 37247 -13844 37659 -13830
rect 38331 -13844 38743 -13830
rect 40282 -13844 40694 -13830
rect 37214 -13915 37659 -13844
rect 38298 -13915 38743 -13844
rect 40249 -13915 40694 -13844
rect 41545 -13845 41957 -13831
rect 43545 -13837 43957 -13823
rect 88397 -13824 88809 -13810
rect 89481 -13824 89893 -13810
rect 91432 -13824 91844 -13810
rect 41512 -13908 41957 -13845
rect 43512 -13908 43957 -13837
rect 88364 -13895 88809 -13824
rect 89448 -13895 89893 -13824
rect 91399 -13895 91844 -13824
rect 92695 -13825 93107 -13811
rect 94695 -13817 95107 -13803
rect 92662 -13888 93107 -13825
rect 94662 -13888 95107 -13817
rect 92662 -13890 95331 -13888
rect 88194 -13897 90170 -13895
rect 91156 -13897 92121 -13895
rect 92662 -13896 93107 -13890
rect 41512 -13910 44181 -13908
rect 88364 -13910 88484 -13897
rect 88544 -13910 88616 -13897
rect 37044 -13917 39020 -13915
rect 40006 -13917 40971 -13915
rect 41512 -13916 41957 -13910
rect 37214 -13930 37334 -13917
rect 37394 -13930 37466 -13917
rect 37300 -13938 37301 -13930
rect 37573 -13938 37659 -13917
rect 38298 -13930 38418 -13917
rect 38478 -13930 38550 -13917
rect 37300 -13939 37659 -13938
rect 38384 -13938 38385 -13930
rect 38657 -13938 38743 -13917
rect 40249 -13930 40369 -13917
rect 40429 -13930 40501 -13917
rect 38384 -13939 38743 -13938
rect 40335 -13938 40336 -13930
rect 40608 -13938 40694 -13917
rect 41269 -13918 42234 -13916
rect 41512 -13931 41632 -13918
rect 41692 -13931 41764 -13918
rect 40335 -13939 40694 -13938
rect 41598 -13939 41599 -13931
rect 41871 -13939 41957 -13918
rect 43512 -13923 43632 -13910
rect 43692 -13923 43764 -13910
rect 43598 -13931 43599 -13923
rect 43871 -13931 43957 -13910
rect 88450 -13918 88451 -13910
rect 88723 -13918 88809 -13897
rect 89448 -13910 89568 -13897
rect 89628 -13910 89700 -13897
rect 88450 -13919 88809 -13918
rect 89534 -13918 89535 -13910
rect 89807 -13918 89893 -13897
rect 91399 -13910 91519 -13897
rect 91579 -13910 91651 -13897
rect 89534 -13919 89893 -13918
rect 91485 -13918 91486 -13910
rect 91758 -13918 91844 -13897
rect 92419 -13898 93384 -13896
rect 92662 -13911 92782 -13898
rect 92842 -13911 92914 -13898
rect 91485 -13919 91844 -13918
rect 92748 -13919 92749 -13911
rect 93021 -13919 93107 -13898
rect 94662 -13903 94782 -13890
rect 94842 -13903 94914 -13890
rect 94748 -13911 94749 -13903
rect 95021 -13911 95107 -13890
rect 94748 -13912 95107 -13911
rect 92748 -13920 93107 -13919
rect 43598 -13932 43957 -13931
rect 41598 -13940 41957 -13939
rect 39262 -16056 39707 -15970
rect 39348 -16078 39349 -16056
rect 39468 -16065 39514 -16056
rect 39621 -16064 39707 -16056
rect 40327 -16064 40772 -15978
rect 42476 -16056 42921 -15970
rect 39588 -16065 39707 -16064
rect 39455 -16078 39527 -16065
rect 39588 -16078 39674 -16065
rect 38985 -16080 39950 -16078
rect 39468 -16092 39481 -16080
rect 39501 -16086 39514 -16080
rect 40413 -16086 40414 -16064
rect 40533 -16073 40579 -16064
rect 40686 -16072 40772 -16064
rect 40653 -16073 40772 -16072
rect 40520 -16086 40592 -16073
rect 40653 -16086 40739 -16073
rect 42562 -16078 42563 -16056
rect 42682 -16065 42728 -16056
rect 42835 -16064 42921 -16056
rect 43584 -16064 44029 -15978
rect 90412 -16036 90857 -15950
rect 90498 -16058 90499 -16036
rect 90618 -16045 90664 -16036
rect 90771 -16044 90857 -16036
rect 91477 -16044 91922 -15958
rect 93626 -16036 94071 -15950
rect 90738 -16045 90857 -16044
rect 90605 -16058 90677 -16045
rect 90738 -16058 90824 -16045
rect 90135 -16060 91100 -16058
rect 42802 -16065 42921 -16064
rect 42669 -16078 42741 -16065
rect 42802 -16078 42888 -16065
rect 43670 -16078 43671 -16064
rect 43790 -16073 43836 -16064
rect 43943 -16072 44029 -16064
rect 90618 -16072 90631 -16060
rect 90651 -16066 90664 -16060
rect 91563 -16066 91564 -16044
rect 91683 -16053 91729 -16044
rect 91836 -16052 91922 -16044
rect 91803 -16053 91922 -16052
rect 91670 -16066 91742 -16053
rect 91803 -16066 91889 -16053
rect 93712 -16058 93713 -16036
rect 93832 -16045 93878 -16036
rect 93985 -16044 94071 -16036
rect 94734 -16044 95179 -15958
rect 93952 -16045 94071 -16044
rect 93819 -16058 93891 -16045
rect 93952 -16058 94038 -16045
rect 94820 -16058 94821 -16044
rect 94940 -16053 94986 -16044
rect 95093 -16052 95179 -16044
rect 95060 -16053 95179 -16052
rect 94927 -16058 94999 -16053
rect 93349 -16060 94999 -16058
rect 93832 -16066 93845 -16060
rect 90651 -16068 93845 -16066
rect 90651 -16072 90664 -16068
rect 43910 -16073 44029 -16072
rect 43777 -16078 43849 -16073
rect 42199 -16080 43849 -16078
rect 42682 -16086 42695 -16080
rect 39501 -16088 42695 -16086
rect 39501 -16092 39514 -16088
rect 40533 -16100 40546 -16088
rect 40566 -16100 40579 -16088
rect 42682 -16092 42695 -16088
rect 42715 -16086 42728 -16080
rect 43670 -16086 43671 -16080
rect 43777 -16086 43849 -16080
rect 43910 -16086 43996 -16073
rect 91683 -16080 91696 -16068
rect 91716 -16080 91729 -16068
rect 93832 -16072 93845 -16068
rect 93865 -16066 93878 -16060
rect 94820 -16066 94821 -16060
rect 94927 -16066 94999 -16060
rect 95060 -16066 95146 -16053
rect 93865 -16068 95337 -16066
rect 93865 -16072 93878 -16068
rect 94940 -16080 94953 -16068
rect 94973 -16080 94986 -16068
rect 42715 -16088 44187 -16086
rect 42715 -16092 42728 -16088
rect 43790 -16100 43803 -16088
rect 43823 -16100 43836 -16088
rect 6763 -16366 7044 -16280
rect 10739 -16366 11020 -16280
rect 20082 -16366 20575 -16280
rect 21419 -16366 21912 -16280
rect 31165 -16366 31446 -16280
rect 35141 -16366 35422 -16280
rect 57913 -16346 58194 -16260
rect 61889 -16346 62170 -16260
rect 71232 -16346 71725 -16260
rect 72569 -16346 73062 -16260
rect 82315 -16346 82596 -16260
rect 86291 -16346 86572 -16260
rect 57999 -16365 58000 -16346
rect 58029 -16352 58075 -16346
rect 58016 -16365 58088 -16352
rect 58108 -16365 58194 -16346
rect 61975 -16365 61976 -16346
rect 62005 -16352 62051 -16346
rect 61992 -16365 62064 -16352
rect 62084 -16365 62170 -16346
rect 6849 -16385 6850 -16366
rect 6879 -16372 6925 -16366
rect 6866 -16385 6938 -16372
rect 6958 -16385 7044 -16366
rect 10825 -16385 10826 -16366
rect 10855 -16372 10901 -16366
rect 10842 -16385 10914 -16372
rect 10934 -16385 11020 -16366
rect 6558 -16387 7476 -16385
rect 9386 -16387 11452 -16385
rect 6879 -16399 6892 -16387
rect 6912 -16399 6925 -16387
rect 10855 -16399 10868 -16387
rect 10888 -16399 10901 -16387
rect 20168 -16444 20169 -16366
rect 20277 -16385 20363 -16366
rect 20380 -16385 20381 -16366
rect 20413 -16372 20459 -16366
rect 20400 -16385 20472 -16372
rect 20489 -16385 20575 -16366
rect 21505 -16385 21506 -16366
rect 21535 -16372 21581 -16366
rect 21522 -16385 21594 -16372
rect 21614 -16385 21700 -16366
rect 21717 -16385 21718 -16366
rect 20245 -16387 20640 -16385
rect 21500 -16387 21749 -16385
rect 20277 -16444 20363 -16387
rect 20413 -16399 20426 -16387
rect 20446 -16399 20459 -16387
rect 21535 -16399 21548 -16387
rect 21568 -16399 21581 -16387
rect 20168 -16445 20363 -16444
rect 21717 -16444 21718 -16387
rect 21826 -16444 21912 -16366
rect 31251 -16385 31252 -16366
rect 31284 -16372 31330 -16366
rect 31271 -16385 31343 -16372
rect 31360 -16385 31446 -16366
rect 35227 -16385 35228 -16366
rect 35260 -16372 35306 -16366
rect 35247 -16385 35319 -16372
rect 35336 -16385 35422 -16366
rect 57708 -16367 58626 -16365
rect 60536 -16367 62602 -16365
rect 58029 -16379 58042 -16367
rect 58062 -16379 58075 -16367
rect 62005 -16379 62018 -16367
rect 62038 -16379 62051 -16367
rect 30733 -16387 32000 -16385
rect 34709 -16387 35627 -16385
rect 31284 -16399 31297 -16387
rect 31317 -16399 31330 -16387
rect 35260 -16399 35273 -16387
rect 35293 -16399 35306 -16387
rect 71318 -16424 71319 -16346
rect 71427 -16365 71513 -16346
rect 71530 -16365 71531 -16346
rect 71563 -16352 71609 -16346
rect 71550 -16365 71622 -16352
rect 71639 -16365 71725 -16346
rect 72655 -16365 72656 -16346
rect 72685 -16352 72731 -16346
rect 72672 -16365 72744 -16352
rect 72764 -16365 72850 -16346
rect 72867 -16365 72868 -16346
rect 71395 -16367 71790 -16365
rect 72650 -16367 72899 -16365
rect 71427 -16424 71513 -16367
rect 71563 -16379 71576 -16367
rect 71596 -16379 71609 -16367
rect 72685 -16379 72698 -16367
rect 72718 -16379 72731 -16367
rect 71318 -16425 71513 -16424
rect 72867 -16424 72868 -16367
rect 72976 -16424 73062 -16346
rect 82401 -16365 82402 -16346
rect 82434 -16352 82480 -16346
rect 82421 -16365 82493 -16352
rect 82510 -16365 82596 -16346
rect 86377 -16365 86378 -16346
rect 86410 -16352 86456 -16346
rect 86397 -16365 86469 -16352
rect 86486 -16365 86572 -16346
rect 81883 -16367 83949 -16365
rect 85859 -16367 86777 -16365
rect 82434 -16379 82447 -16367
rect 82467 -16379 82480 -16367
rect 86410 -16379 86423 -16367
rect 86443 -16379 86456 -16367
rect 72867 -16425 73062 -16424
rect 21717 -16445 21912 -16444
rect 17790 -17369 18107 -17319
rect 19851 -17369 20168 -17319
rect 21794 -17342 22206 -17328
rect 22878 -17342 23290 -17328
rect 24829 -17342 25241 -17328
rect 16832 -17371 18569 -17369
rect 19786 -17371 20700 -17369
rect 17876 -17423 17877 -17371
rect 17917 -17384 17989 -17371
rect 18021 -17423 18107 -17371
rect 17876 -17424 18107 -17423
rect 19937 -17423 19938 -17371
rect 19978 -17384 20050 -17371
rect 20082 -17423 20168 -17371
rect 21761 -17413 22206 -17342
rect 22845 -17413 23290 -17342
rect 24796 -17413 25241 -17342
rect 26092 -17343 26504 -17329
rect 28092 -17335 28504 -17321
rect 30144 -17335 30556 -17321
rect 31228 -17335 31640 -17321
rect 33179 -17335 33591 -17321
rect 26059 -17406 26504 -17343
rect 28059 -17406 28504 -17335
rect 30111 -17406 30556 -17335
rect 31195 -17406 31640 -17335
rect 33146 -17406 33591 -17335
rect 34442 -17336 34854 -17322
rect 36442 -17328 36854 -17314
rect 34409 -17399 34854 -17336
rect 36409 -17399 36854 -17328
rect 38170 -17386 38451 -17304
rect 68940 -17349 69257 -17299
rect 71001 -17349 71318 -17299
rect 72944 -17322 73356 -17308
rect 74028 -17322 74440 -17308
rect 75979 -17322 76391 -17308
rect 67982 -17351 69719 -17349
rect 70936 -17351 71850 -17349
rect 37965 -17388 38883 -17386
rect 34409 -17401 37078 -17399
rect 26059 -17408 28728 -17406
rect 29941 -17408 31917 -17406
rect 32903 -17408 33868 -17406
rect 34409 -17407 34854 -17401
rect 21591 -17415 23567 -17413
rect 24553 -17415 25518 -17413
rect 26059 -17414 26504 -17408
rect 19937 -17424 20168 -17423
rect 21761 -17428 21881 -17415
rect 21941 -17428 22013 -17415
rect 21847 -17436 21848 -17428
rect 22120 -17436 22206 -17415
rect 22845 -17428 22965 -17415
rect 23025 -17428 23097 -17415
rect 21847 -17437 22206 -17436
rect 22931 -17436 22932 -17428
rect 23204 -17436 23290 -17415
rect 24796 -17428 24916 -17415
rect 24976 -17428 25048 -17415
rect 22931 -17437 23290 -17436
rect 24882 -17436 24883 -17428
rect 25155 -17436 25241 -17415
rect 25816 -17416 26781 -17414
rect 26059 -17429 26179 -17416
rect 26239 -17429 26311 -17416
rect 24882 -17437 25241 -17436
rect 26145 -17437 26146 -17429
rect 26418 -17437 26504 -17416
rect 28059 -17421 28179 -17408
rect 28239 -17421 28311 -17408
rect 28145 -17429 28146 -17421
rect 28418 -17429 28504 -17408
rect 30111 -17421 30231 -17408
rect 30291 -17421 30363 -17408
rect 28145 -17430 28504 -17429
rect 30197 -17429 30198 -17421
rect 30470 -17429 30556 -17408
rect 31195 -17421 31315 -17408
rect 31375 -17421 31447 -17408
rect 30197 -17430 30556 -17429
rect 31281 -17429 31282 -17421
rect 31554 -17429 31640 -17408
rect 33146 -17421 33266 -17408
rect 33326 -17421 33398 -17408
rect 31281 -17430 31640 -17429
rect 33232 -17429 33233 -17421
rect 33505 -17429 33591 -17408
rect 34166 -17409 35131 -17407
rect 34409 -17422 34529 -17409
rect 34589 -17422 34661 -17409
rect 33232 -17430 33591 -17429
rect 34495 -17430 34496 -17422
rect 34768 -17430 34854 -17409
rect 36409 -17414 36529 -17401
rect 36589 -17414 36661 -17401
rect 36495 -17422 36496 -17414
rect 36768 -17422 36854 -17401
rect 38256 -17406 38257 -17388
rect 38273 -17401 38345 -17388
rect 38365 -17406 38451 -17388
rect 69026 -17403 69027 -17351
rect 69067 -17364 69139 -17351
rect 69171 -17403 69257 -17351
rect 69026 -17404 69257 -17403
rect 71087 -17403 71088 -17351
rect 71128 -17364 71200 -17351
rect 71232 -17403 71318 -17351
rect 72911 -17393 73356 -17322
rect 73995 -17393 74440 -17322
rect 75946 -17393 76391 -17322
rect 77242 -17323 77654 -17309
rect 79242 -17315 79654 -17301
rect 81294 -17315 81706 -17301
rect 82378 -17315 82790 -17301
rect 84329 -17315 84741 -17301
rect 77209 -17386 77654 -17323
rect 79209 -17386 79654 -17315
rect 81261 -17386 81706 -17315
rect 82345 -17386 82790 -17315
rect 84296 -17386 84741 -17315
rect 85592 -17316 86004 -17302
rect 87592 -17308 88004 -17294
rect 85559 -17379 86004 -17316
rect 87559 -17379 88004 -17308
rect 89320 -17366 89601 -17284
rect 89115 -17368 90033 -17366
rect 85559 -17381 88228 -17379
rect 77209 -17388 79878 -17386
rect 81091 -17388 83067 -17386
rect 84053 -17388 85018 -17386
rect 85559 -17387 86004 -17381
rect 72741 -17395 74717 -17393
rect 75703 -17395 76668 -17393
rect 77209 -17394 77654 -17388
rect 71087 -17404 71318 -17403
rect 38256 -17407 38451 -17406
rect 72911 -17408 73031 -17395
rect 73091 -17408 73163 -17395
rect 72997 -17416 72998 -17408
rect 73270 -17416 73356 -17395
rect 73995 -17408 74115 -17395
rect 74175 -17408 74247 -17395
rect 72997 -17417 73356 -17416
rect 74081 -17416 74082 -17408
rect 74354 -17416 74440 -17395
rect 75946 -17408 76066 -17395
rect 76126 -17408 76198 -17395
rect 74081 -17417 74440 -17416
rect 76032 -17416 76033 -17408
rect 76305 -17416 76391 -17395
rect 76966 -17396 77931 -17394
rect 77209 -17409 77329 -17396
rect 77389 -17409 77461 -17396
rect 76032 -17417 76391 -17416
rect 77295 -17417 77296 -17409
rect 77568 -17417 77654 -17396
rect 79209 -17401 79329 -17388
rect 79389 -17401 79461 -17388
rect 79295 -17409 79296 -17401
rect 79568 -17409 79654 -17388
rect 81261 -17401 81381 -17388
rect 81441 -17401 81513 -17388
rect 79295 -17410 79654 -17409
rect 81347 -17409 81348 -17401
rect 81620 -17409 81706 -17388
rect 82345 -17401 82465 -17388
rect 82525 -17401 82597 -17388
rect 81347 -17410 81706 -17409
rect 82431 -17409 82432 -17401
rect 82704 -17409 82790 -17388
rect 84296 -17401 84416 -17388
rect 84476 -17401 84548 -17388
rect 82431 -17410 82790 -17409
rect 84382 -17409 84383 -17401
rect 84655 -17409 84741 -17388
rect 85316 -17389 86281 -17387
rect 85559 -17402 85679 -17389
rect 85739 -17402 85811 -17389
rect 84382 -17410 84741 -17409
rect 85645 -17410 85646 -17402
rect 85918 -17410 86004 -17389
rect 87559 -17394 87679 -17381
rect 87739 -17394 87811 -17381
rect 87645 -17402 87646 -17394
rect 87918 -17402 88004 -17381
rect 89406 -17386 89407 -17368
rect 89423 -17381 89495 -17368
rect 89515 -17386 89601 -17368
rect 89406 -17387 89601 -17386
rect 87645 -17403 88004 -17402
rect 85645 -17411 86004 -17410
rect 77295 -17418 77654 -17417
rect 36495 -17423 36854 -17422
rect 34495 -17431 34854 -17430
rect 26145 -17438 26504 -17437
rect 6912 -17543 7324 -17529
rect 6879 -17590 7324 -17543
rect 8081 -17590 8408 -17519
rect 9175 -17543 9587 -17529
rect 10407 -17543 10819 -17529
rect 9142 -17590 9587 -17543
rect 6879 -17592 9587 -17590
rect 6879 -17614 7324 -17592
rect 8167 -17614 8168 -17592
rect 8212 -17605 8284 -17592
rect 8225 -17610 8235 -17605
rect 8271 -17610 8281 -17609
rect 8235 -17614 8321 -17610
rect 8322 -17614 8408 -17592
rect 9142 -17614 9587 -17592
rect 10374 -17590 10819 -17543
rect 11576 -17590 11903 -17519
rect 12670 -17543 13082 -17529
rect 13996 -17543 14408 -17529
rect 12637 -17590 13082 -17543
rect 10374 -17592 13082 -17590
rect 10374 -17614 10819 -17592
rect 11662 -17614 11663 -17592
rect 11707 -17605 11779 -17592
rect 11720 -17610 11730 -17605
rect 11766 -17610 11776 -17609
rect 11730 -17614 11816 -17610
rect 11817 -17614 11903 -17592
rect 12637 -17614 13082 -17592
rect 13963 -17590 14408 -17543
rect 15165 -17590 15492 -17519
rect 58062 -17523 58474 -17509
rect 16259 -17543 16671 -17529
rect 16226 -17590 16671 -17543
rect 13963 -17592 16671 -17590
rect 13963 -17614 14408 -17592
rect 15251 -17614 15252 -17592
rect 15296 -17605 15368 -17592
rect 15309 -17610 15319 -17605
rect 15355 -17610 15365 -17609
rect 15319 -17614 15405 -17610
rect 15406 -17614 15492 -17592
rect 16226 -17614 16671 -17592
rect 58029 -17570 58474 -17523
rect 59231 -17570 59558 -17499
rect 60325 -17523 60737 -17509
rect 61557 -17523 61969 -17509
rect 60292 -17570 60737 -17523
rect 58029 -17572 60737 -17570
rect 58029 -17594 58474 -17572
rect 59317 -17594 59318 -17572
rect 59362 -17585 59434 -17572
rect 59375 -17590 59385 -17585
rect 59421 -17590 59431 -17589
rect 59385 -17594 59471 -17590
rect 59472 -17594 59558 -17572
rect 60292 -17594 60737 -17572
rect 61524 -17570 61969 -17523
rect 62726 -17570 63053 -17499
rect 63820 -17523 64232 -17509
rect 65146 -17523 65558 -17509
rect 63787 -17570 64232 -17523
rect 61524 -17572 64232 -17570
rect 61524 -17594 61969 -17572
rect 62812 -17594 62813 -17572
rect 62857 -17585 62929 -17572
rect 62870 -17590 62880 -17585
rect 62916 -17590 62926 -17589
rect 62880 -17594 62966 -17590
rect 62967 -17594 63053 -17572
rect 63787 -17594 64232 -17572
rect 65113 -17570 65558 -17523
rect 66315 -17570 66642 -17499
rect 67409 -17523 67821 -17509
rect 67376 -17570 67821 -17523
rect 65113 -17572 67821 -17570
rect 65113 -17594 65558 -17572
rect 66401 -17594 66402 -17572
rect 66446 -17585 66518 -17572
rect 66459 -17590 66469 -17585
rect 66505 -17590 66515 -17589
rect 66469 -17594 66555 -17590
rect 66556 -17594 66642 -17572
rect 67376 -17594 67821 -17572
rect 57431 -17596 68098 -17594
rect 58029 -17609 58149 -17596
rect 58209 -17609 58281 -17596
rect 6281 -17616 16948 -17614
rect 6879 -17629 6999 -17616
rect 7059 -17629 7131 -17616
rect 6965 -17637 6966 -17629
rect 7238 -17637 7324 -17616
rect 8167 -17622 8168 -17616
rect 8235 -17622 8321 -17616
rect 8322 -17622 8408 -17616
rect 8167 -17623 8408 -17622
rect 9142 -17629 9262 -17616
rect 9322 -17629 9394 -17616
rect 6965 -17638 7324 -17637
rect 9228 -17637 9229 -17629
rect 9501 -17637 9587 -17616
rect 10374 -17629 10494 -17616
rect 10554 -17629 10626 -17616
rect 9228 -17638 9587 -17637
rect 10460 -17637 10461 -17629
rect 10733 -17637 10819 -17616
rect 11662 -17622 11663 -17616
rect 11730 -17622 11816 -17616
rect 11817 -17622 11903 -17616
rect 11662 -17623 11903 -17622
rect 12637 -17629 12757 -17616
rect 12817 -17629 12889 -17616
rect 10460 -17638 10819 -17637
rect 12723 -17637 12724 -17629
rect 12996 -17637 13082 -17616
rect 13963 -17629 14083 -17616
rect 14143 -17629 14215 -17616
rect 12723 -17638 13082 -17637
rect 14049 -17637 14050 -17629
rect 14322 -17637 14408 -17616
rect 15251 -17622 15252 -17616
rect 15319 -17622 15405 -17616
rect 15406 -17622 15492 -17616
rect 15251 -17623 15492 -17622
rect 16226 -17629 16346 -17616
rect 16406 -17629 16478 -17616
rect 14049 -17638 14408 -17637
rect 16312 -17637 16313 -17629
rect 16585 -17637 16671 -17616
rect 58115 -17617 58116 -17609
rect 58388 -17617 58474 -17596
rect 59317 -17602 59318 -17596
rect 59385 -17602 59471 -17596
rect 59472 -17602 59558 -17596
rect 59317 -17603 59558 -17602
rect 60292 -17609 60412 -17596
rect 60472 -17609 60544 -17596
rect 58115 -17618 58474 -17617
rect 60378 -17617 60379 -17609
rect 60651 -17617 60737 -17596
rect 61524 -17609 61644 -17596
rect 61704 -17609 61776 -17596
rect 60378 -17618 60737 -17617
rect 61610 -17617 61611 -17609
rect 61883 -17617 61969 -17596
rect 62812 -17602 62813 -17596
rect 62880 -17602 62966 -17596
rect 62967 -17602 63053 -17596
rect 62812 -17603 63053 -17602
rect 63787 -17609 63907 -17596
rect 63967 -17609 64039 -17596
rect 61610 -17618 61969 -17617
rect 63873 -17617 63874 -17609
rect 64146 -17617 64232 -17596
rect 65113 -17609 65233 -17596
rect 65293 -17609 65365 -17596
rect 63873 -17618 64232 -17617
rect 65199 -17617 65200 -17609
rect 65472 -17617 65558 -17596
rect 66401 -17602 66402 -17596
rect 66469 -17602 66555 -17596
rect 66556 -17602 66642 -17596
rect 66401 -17603 66642 -17602
rect 67376 -17609 67496 -17596
rect 67556 -17609 67628 -17596
rect 65199 -17618 65558 -17617
rect 67462 -17617 67463 -17609
rect 67735 -17617 67821 -17596
rect 67462 -17618 67821 -17617
rect 16312 -17638 16671 -17637
rect 23809 -19554 24254 -19468
rect 23895 -19576 23896 -19554
rect 24015 -19563 24061 -19554
rect 24168 -19562 24254 -19554
rect 24874 -19562 25319 -19476
rect 27023 -19554 27468 -19468
rect 24135 -19563 24254 -19562
rect 24002 -19576 24074 -19563
rect 24135 -19576 24221 -19563
rect 23532 -19578 24497 -19576
rect 24015 -19590 24028 -19578
rect 24048 -19584 24061 -19578
rect 24960 -19584 24961 -19562
rect 25080 -19571 25126 -19562
rect 25233 -19570 25319 -19562
rect 25200 -19571 25319 -19570
rect 25067 -19584 25139 -19571
rect 25200 -19584 25286 -19571
rect 27109 -19576 27110 -19554
rect 27229 -19563 27275 -19554
rect 27382 -19562 27468 -19554
rect 28131 -19562 28576 -19476
rect 32159 -19547 32604 -19461
rect 27349 -19563 27468 -19562
rect 27216 -19576 27288 -19563
rect 27349 -19576 27435 -19563
rect 26746 -19578 28016 -19576
rect 27229 -19584 27242 -19578
rect 24048 -19586 27242 -19584
rect 24048 -19590 24061 -19586
rect 25080 -19598 25093 -19586
rect 25113 -19598 25126 -19586
rect 27229 -19590 27242 -19586
rect 27262 -19590 27275 -19578
rect 28217 -19584 28218 -19562
rect 28337 -19571 28383 -19562
rect 28490 -19570 28576 -19562
rect 32245 -19569 32246 -19547
rect 32365 -19556 32411 -19547
rect 32518 -19555 32604 -19547
rect 33224 -19555 33669 -19469
rect 35373 -19547 35818 -19461
rect 32485 -19556 32604 -19555
rect 32352 -19569 32424 -19556
rect 32485 -19569 32571 -19556
rect 28457 -19571 28576 -19570
rect 32000 -19571 32847 -19569
rect 28324 -19584 28396 -19571
rect 28457 -19584 28543 -19571
rect 32365 -19583 32378 -19571
rect 32398 -19577 32411 -19571
rect 33310 -19577 33311 -19555
rect 33430 -19564 33476 -19555
rect 33583 -19563 33669 -19555
rect 33550 -19564 33669 -19563
rect 33417 -19577 33489 -19564
rect 33550 -19577 33636 -19564
rect 35459 -19569 35460 -19547
rect 35579 -19556 35625 -19547
rect 35732 -19555 35818 -19547
rect 36481 -19555 36926 -19469
rect 74959 -19534 75404 -19448
rect 35699 -19556 35818 -19555
rect 35566 -19569 35638 -19556
rect 35699 -19569 35785 -19556
rect 36567 -19569 36568 -19555
rect 36687 -19564 36733 -19555
rect 36840 -19563 36926 -19555
rect 75045 -19556 75046 -19534
rect 75165 -19543 75211 -19534
rect 75318 -19542 75404 -19534
rect 76024 -19542 76469 -19456
rect 78173 -19534 78618 -19448
rect 75285 -19543 75404 -19542
rect 75152 -19556 75224 -19543
rect 75285 -19556 75371 -19543
rect 74682 -19558 75647 -19556
rect 36807 -19564 36926 -19563
rect 36674 -19569 36746 -19564
rect 35096 -19571 36746 -19569
rect 35579 -19577 35592 -19571
rect 32398 -19579 35592 -19577
rect 32398 -19583 32411 -19579
rect 28217 -19585 28734 -19584
rect 28223 -19586 28734 -19585
rect 28337 -19598 28350 -19586
rect 28370 -19598 28383 -19586
rect 33430 -19591 33443 -19579
rect 33463 -19591 33476 -19579
rect 35579 -19583 35592 -19579
rect 35612 -19577 35625 -19571
rect 36567 -19577 36568 -19571
rect 36674 -19577 36746 -19571
rect 36807 -19577 36893 -19564
rect 75165 -19570 75178 -19558
rect 75198 -19564 75211 -19558
rect 76110 -19564 76111 -19542
rect 76230 -19551 76276 -19542
rect 76383 -19550 76469 -19542
rect 76350 -19551 76469 -19550
rect 76217 -19564 76289 -19551
rect 76350 -19564 76436 -19551
rect 78259 -19556 78260 -19534
rect 78379 -19543 78425 -19534
rect 78532 -19542 78618 -19534
rect 79281 -19542 79726 -19456
rect 83309 -19527 83754 -19441
rect 78499 -19543 78618 -19542
rect 78366 -19556 78438 -19543
rect 78499 -19556 78585 -19543
rect 77896 -19558 79166 -19556
rect 78379 -19564 78392 -19558
rect 75198 -19566 78392 -19564
rect 75198 -19570 75211 -19566
rect 35612 -19579 37084 -19577
rect 76230 -19578 76243 -19566
rect 76263 -19578 76276 -19566
rect 78379 -19570 78392 -19566
rect 78412 -19570 78425 -19558
rect 79367 -19564 79368 -19542
rect 79487 -19551 79533 -19542
rect 79640 -19550 79726 -19542
rect 83395 -19549 83396 -19527
rect 83515 -19536 83561 -19527
rect 83668 -19535 83754 -19527
rect 84374 -19535 84819 -19449
rect 86523 -19527 86968 -19441
rect 83635 -19536 83754 -19535
rect 83502 -19549 83574 -19536
rect 83635 -19549 83721 -19536
rect 79607 -19551 79726 -19550
rect 83032 -19551 83997 -19549
rect 79474 -19564 79546 -19551
rect 79607 -19564 79693 -19551
rect 83515 -19563 83528 -19551
rect 83548 -19557 83561 -19551
rect 84460 -19557 84461 -19535
rect 84580 -19544 84626 -19535
rect 84733 -19543 84819 -19535
rect 84700 -19544 84819 -19543
rect 84567 -19557 84639 -19544
rect 84700 -19557 84786 -19544
rect 86609 -19549 86610 -19527
rect 86729 -19536 86775 -19527
rect 86882 -19535 86968 -19527
rect 87631 -19535 88076 -19449
rect 86849 -19536 86968 -19535
rect 86716 -19549 86788 -19536
rect 86849 -19549 86935 -19536
rect 87717 -19549 87718 -19535
rect 87837 -19544 87883 -19535
rect 87990 -19543 88076 -19535
rect 87957 -19544 88076 -19543
rect 87824 -19549 87896 -19544
rect 86246 -19551 87896 -19549
rect 86729 -19557 86742 -19551
rect 83548 -19559 86742 -19557
rect 83548 -19563 83561 -19559
rect 79367 -19565 79884 -19564
rect 79373 -19566 79884 -19565
rect 79487 -19578 79500 -19566
rect 79520 -19578 79533 -19566
rect 84580 -19571 84593 -19559
rect 84613 -19571 84626 -19559
rect 86729 -19563 86742 -19559
rect 86762 -19557 86775 -19551
rect 87717 -19557 87718 -19551
rect 87824 -19557 87896 -19551
rect 87957 -19557 88043 -19544
rect 86762 -19559 88234 -19557
rect 86762 -19563 86775 -19559
rect 87837 -19571 87850 -19559
rect 87870 -19571 87883 -19559
rect 35612 -19583 35625 -19579
rect 36687 -19591 36700 -19579
rect 36720 -19591 36733 -19579
rect 6861 -21053 7306 -20967
rect 6947 -21061 6948 -21053
rect 6947 -21062 6980 -21061
rect 7054 -21062 7100 -21053
rect 6980 -21075 6981 -21062
rect 7041 -21075 7113 -21062
rect 7220 -21075 7306 -21053
rect 8063 -21068 8390 -20982
rect 9124 -21053 9569 -20967
rect 10356 -21053 10801 -20967
rect 9210 -21061 9211 -21053
rect 9210 -21062 9243 -21061
rect 9317 -21062 9363 -21053
rect 8149 -21075 8150 -21068
rect 8207 -21075 8303 -21068
rect 8304 -21075 8390 -21068
rect 9243 -21075 9244 -21062
rect 9304 -21075 9376 -21062
rect 9483 -21075 9569 -21053
rect 10442 -21061 10443 -21053
rect 10442 -21062 10475 -21061
rect 10549 -21062 10595 -21053
rect 10475 -21075 10476 -21062
rect 10536 -21075 10608 -21062
rect 10715 -21075 10801 -21053
rect 11558 -21068 11885 -20982
rect 12619 -21053 13064 -20967
rect 13843 -21053 14288 -20967
rect 12705 -21061 12706 -21053
rect 12705 -21062 12738 -21061
rect 12812 -21062 12858 -21053
rect 11644 -21075 11645 -21068
rect 11702 -21075 11798 -21068
rect 11799 -21075 11885 -21068
rect 12738 -21075 12739 -21062
rect 12799 -21075 12871 -21062
rect 12978 -21075 13064 -21053
rect 13929 -21061 13930 -21053
rect 13929 -21062 13962 -21061
rect 14036 -21062 14082 -21053
rect 13962 -21075 13963 -21062
rect 14023 -21075 14095 -21062
rect 14202 -21075 14288 -21053
rect 15045 -21068 15372 -20982
rect 16106 -21053 16551 -20967
rect 17494 -21053 17939 -20967
rect 16192 -21061 16193 -21053
rect 16192 -21062 16225 -21061
rect 16299 -21062 16345 -21053
rect 15131 -21075 15132 -21068
rect 15189 -21075 15285 -21068
rect 15286 -21075 15372 -21068
rect 16225 -21075 16226 -21062
rect 16286 -21075 16358 -21062
rect 16465 -21075 16551 -21053
rect 17580 -21061 17581 -21053
rect 17580 -21062 17613 -21061
rect 17687 -21062 17733 -21053
rect 17613 -21075 17614 -21062
rect 17674 -21075 17746 -21062
rect 17853 -21075 17939 -21053
rect 18696 -21068 19023 -20982
rect 19757 -21053 20202 -20967
rect 58011 -21033 58456 -20947
rect 58097 -21041 58098 -21033
rect 58097 -21042 58130 -21041
rect 58204 -21042 58250 -21033
rect 19843 -21061 19844 -21053
rect 19843 -21062 19876 -21061
rect 19950 -21062 19996 -21053
rect 18782 -21075 18783 -21068
rect 18840 -21075 18936 -21068
rect 18937 -21075 19023 -21068
rect 19876 -21075 19877 -21062
rect 19937 -21075 20009 -21062
rect 20116 -21075 20202 -21053
rect 58130 -21055 58131 -21042
rect 58191 -21055 58263 -21042
rect 58370 -21055 58456 -21033
rect 59213 -21048 59540 -20962
rect 60274 -21033 60719 -20947
rect 61506 -21033 61951 -20947
rect 60360 -21041 60361 -21033
rect 60360 -21042 60393 -21041
rect 60467 -21042 60513 -21033
rect 59299 -21055 59300 -21048
rect 59357 -21055 59453 -21048
rect 59454 -21055 59540 -21048
rect 60393 -21055 60394 -21042
rect 60454 -21055 60526 -21042
rect 60633 -21055 60719 -21033
rect 61592 -21041 61593 -21033
rect 61592 -21042 61625 -21041
rect 61699 -21042 61745 -21033
rect 61625 -21055 61626 -21042
rect 61686 -21055 61758 -21042
rect 61865 -21055 61951 -21033
rect 62708 -21048 63035 -20962
rect 63769 -21033 64214 -20947
rect 64993 -21033 65438 -20947
rect 63855 -21041 63856 -21033
rect 63855 -21042 63888 -21041
rect 63962 -21042 64008 -21033
rect 62794 -21055 62795 -21048
rect 62852 -21055 62948 -21048
rect 62949 -21055 63035 -21048
rect 63888 -21055 63889 -21042
rect 63949 -21055 64021 -21042
rect 64128 -21055 64214 -21033
rect 65079 -21041 65080 -21033
rect 65079 -21042 65112 -21041
rect 65186 -21042 65232 -21033
rect 65112 -21055 65113 -21042
rect 65173 -21055 65245 -21042
rect 65352 -21055 65438 -21033
rect 66195 -21048 66522 -20962
rect 67256 -21033 67701 -20947
rect 68644 -21033 69089 -20947
rect 67342 -21041 67343 -21033
rect 67342 -21042 67375 -21041
rect 67449 -21042 67495 -21033
rect 66281 -21055 66282 -21048
rect 66339 -21055 66435 -21048
rect 66436 -21055 66522 -21048
rect 67375 -21055 67376 -21042
rect 67436 -21055 67508 -21042
rect 67615 -21055 67701 -21033
rect 68730 -21041 68731 -21033
rect 68730 -21042 68763 -21041
rect 68837 -21042 68883 -21033
rect 68763 -21055 68764 -21042
rect 68824 -21055 68896 -21042
rect 69003 -21055 69089 -21033
rect 69846 -21048 70173 -20962
rect 70907 -21033 71352 -20947
rect 70993 -21041 70994 -21033
rect 70993 -21042 71026 -21041
rect 71100 -21042 71146 -21033
rect 69932 -21055 69933 -21048
rect 69990 -21055 70086 -21048
rect 70087 -21055 70173 -21048
rect 71026 -21055 71027 -21042
rect 71087 -21055 71159 -21042
rect 71266 -21055 71352 -21033
rect 57431 -21057 74935 -21055
rect 58204 -21069 58217 -21057
rect 58237 -21069 58250 -21057
rect 6281 -21077 23785 -21075
rect 7054 -21089 7067 -21077
rect 7087 -21089 7100 -21077
rect 8149 -21099 8150 -21077
rect 8207 -21081 8303 -21077
rect 8207 -21086 8253 -21081
rect 8194 -21099 8266 -21086
rect 8304 -21099 8390 -21077
rect 9317 -21089 9330 -21077
rect 9350 -21089 9363 -21077
rect 10549 -21089 10562 -21077
rect 10582 -21089 10595 -21077
rect 11644 -21099 11645 -21077
rect 11702 -21081 11798 -21077
rect 11702 -21086 11748 -21081
rect 11689 -21099 11761 -21086
rect 11799 -21099 11885 -21077
rect 12812 -21089 12825 -21077
rect 12845 -21089 12858 -21077
rect 14036 -21089 14049 -21077
rect 14069 -21089 14082 -21077
rect 15131 -21099 15132 -21077
rect 15189 -21081 15285 -21077
rect 15189 -21086 15235 -21081
rect 15176 -21099 15248 -21086
rect 15286 -21099 15372 -21077
rect 16299 -21089 16312 -21077
rect 16332 -21089 16345 -21077
rect 17687 -21089 17700 -21077
rect 17720 -21089 17733 -21077
rect 18782 -21099 18783 -21077
rect 18840 -21081 18936 -21077
rect 18840 -21086 18886 -21081
rect 18827 -21099 18899 -21086
rect 18937 -21099 19023 -21077
rect 19950 -21089 19963 -21077
rect 19983 -21089 19996 -21077
rect 59299 -21079 59300 -21057
rect 59357 -21061 59453 -21057
rect 59357 -21066 59403 -21061
rect 59344 -21079 59416 -21066
rect 59454 -21079 59540 -21057
rect 60467 -21069 60480 -21057
rect 60500 -21069 60513 -21057
rect 61699 -21069 61712 -21057
rect 61732 -21069 61745 -21057
rect 62794 -21079 62795 -21057
rect 62852 -21061 62948 -21057
rect 62852 -21066 62898 -21061
rect 62839 -21079 62911 -21066
rect 62949 -21079 63035 -21057
rect 63962 -21069 63975 -21057
rect 63995 -21069 64008 -21057
rect 65186 -21069 65199 -21057
rect 65219 -21069 65232 -21057
rect 66281 -21079 66282 -21057
rect 66339 -21061 66435 -21057
rect 66339 -21066 66385 -21061
rect 66326 -21079 66398 -21066
rect 66436 -21079 66522 -21057
rect 67449 -21069 67462 -21057
rect 67482 -21069 67495 -21057
rect 68837 -21069 68850 -21057
rect 68870 -21069 68883 -21057
rect 69932 -21079 69933 -21057
rect 69990 -21061 70086 -21057
rect 69990 -21066 70036 -21061
rect 69977 -21079 70049 -21066
rect 70087 -21079 70173 -21057
rect 71100 -21069 71113 -21057
rect 71133 -21069 71146 -21057
rect 58250 -21081 60467 -21079
rect 61745 -21080 63035 -21079
rect 61745 -21081 62959 -21080
rect 65232 -21081 67449 -21079
rect 68883 -21081 71100 -21079
rect 59357 -21093 59370 -21081
rect 59390 -21093 59403 -21081
rect 62852 -21093 62865 -21081
rect 62885 -21093 62898 -21081
rect 66339 -21093 66352 -21081
rect 66372 -21093 66385 -21081
rect 69990 -21093 70003 -21081
rect 70023 -21093 70036 -21081
rect 7100 -21101 9317 -21099
rect 10595 -21100 11885 -21099
rect 10595 -21101 11809 -21100
rect 14082 -21101 16299 -21099
rect 17733 -21101 19950 -21099
rect 8207 -21113 8220 -21101
rect 8240 -21113 8253 -21101
rect 11702 -21113 11715 -21101
rect 11735 -21113 11748 -21101
rect 15189 -21113 15202 -21101
rect 15222 -21113 15235 -21101
rect 18840 -21113 18853 -21101
rect 18873 -21113 18886 -21101
rect 17790 -21867 18107 -21817
rect 19851 -21867 20168 -21817
rect 21794 -21836 22206 -21822
rect 22878 -21836 23290 -21822
rect 24829 -21836 25241 -21822
rect 16832 -21869 18569 -21867
rect 19786 -21869 20700 -21867
rect 17876 -21921 17877 -21869
rect 17917 -21882 17989 -21869
rect 18021 -21921 18107 -21869
rect 17876 -21922 18107 -21921
rect 19937 -21921 19938 -21869
rect 19978 -21882 20050 -21869
rect 20082 -21921 20168 -21869
rect 21761 -21907 22206 -21836
rect 22845 -21907 23290 -21836
rect 24796 -21907 25241 -21836
rect 26092 -21837 26504 -21823
rect 28092 -21829 28504 -21815
rect 21591 -21909 23567 -21907
rect 24553 -21909 25518 -21907
rect 26059 -21908 26504 -21837
rect 28059 -21900 28504 -21829
rect 31332 -21837 31744 -21823
rect 32416 -21837 32828 -21823
rect 34367 -21837 34779 -21823
rect 28059 -21901 28528 -21900
rect 19937 -21922 20168 -21921
rect 21761 -21922 21881 -21909
rect 21941 -21922 22013 -21909
rect 21847 -21930 21848 -21922
rect 22120 -21930 22206 -21909
rect 22845 -21922 22965 -21909
rect 23025 -21922 23097 -21909
rect 21847 -21931 22206 -21930
rect 22931 -21930 22932 -21922
rect 23204 -21930 23290 -21909
rect 24796 -21922 24916 -21909
rect 24976 -21922 25048 -21909
rect 22931 -21931 23290 -21930
rect 24882 -21930 24883 -21922
rect 25155 -21930 25241 -21909
rect 25816 -21910 26781 -21908
rect 26059 -21923 26179 -21910
rect 26239 -21923 26311 -21910
rect 24882 -21931 25241 -21930
rect 26145 -21931 26146 -21923
rect 26418 -21931 26504 -21910
rect 28059 -21915 28179 -21901
rect 28189 -21902 28528 -21901
rect 28239 -21915 28311 -21902
rect 28145 -21923 28146 -21915
rect 28418 -21923 28504 -21902
rect 31299 -21908 31744 -21837
rect 32383 -21908 32828 -21837
rect 34334 -21908 34779 -21837
rect 35630 -21838 36042 -21824
rect 37630 -21830 38042 -21816
rect 35597 -21901 36042 -21838
rect 37597 -21901 38042 -21830
rect 68940 -21847 69257 -21797
rect 71001 -21847 71318 -21797
rect 72944 -21816 73356 -21802
rect 74028 -21816 74440 -21802
rect 75979 -21816 76391 -21802
rect 67982 -21849 69719 -21847
rect 70936 -21849 71850 -21847
rect 69026 -21901 69027 -21849
rect 69067 -21862 69139 -21849
rect 69171 -21901 69257 -21849
rect 35597 -21903 38266 -21901
rect 69026 -21902 69257 -21901
rect 71087 -21901 71088 -21849
rect 71128 -21862 71200 -21849
rect 71232 -21901 71318 -21849
rect 72911 -21887 73356 -21816
rect 73995 -21887 74440 -21816
rect 75946 -21887 76391 -21816
rect 77242 -21817 77654 -21803
rect 79242 -21809 79654 -21795
rect 72741 -21889 74717 -21887
rect 75703 -21889 76668 -21887
rect 77209 -21888 77654 -21817
rect 79209 -21880 79654 -21809
rect 82482 -21817 82894 -21803
rect 83566 -21817 83978 -21803
rect 85517 -21817 85929 -21803
rect 79209 -21881 79678 -21880
rect 71087 -21902 71318 -21901
rect 72911 -21902 73031 -21889
rect 73091 -21902 73163 -21889
rect 31129 -21910 33105 -21908
rect 34091 -21910 35056 -21908
rect 35597 -21909 36042 -21903
rect 31299 -21923 31419 -21910
rect 31479 -21923 31551 -21910
rect 28145 -21924 28504 -21923
rect 26145 -21932 26504 -21931
rect 31385 -21931 31386 -21923
rect 31658 -21931 31744 -21910
rect 32383 -21923 32503 -21910
rect 32563 -21923 32635 -21910
rect 31385 -21932 31744 -21931
rect 32469 -21931 32470 -21923
rect 32742 -21931 32828 -21910
rect 34334 -21923 34454 -21910
rect 34514 -21923 34586 -21910
rect 32469 -21932 32828 -21931
rect 34420 -21931 34421 -21923
rect 34693 -21931 34779 -21910
rect 35354 -21911 36319 -21909
rect 35597 -21924 35717 -21911
rect 35777 -21924 35849 -21911
rect 34420 -21932 34779 -21931
rect 35683 -21932 35684 -21924
rect 35956 -21932 36042 -21911
rect 37597 -21916 37717 -21903
rect 37777 -21916 37849 -21903
rect 37683 -21924 37684 -21916
rect 37956 -21924 38042 -21903
rect 72997 -21910 72998 -21902
rect 73270 -21910 73356 -21889
rect 73995 -21902 74115 -21889
rect 74175 -21902 74247 -21889
rect 72997 -21911 73356 -21910
rect 74081 -21910 74082 -21902
rect 74354 -21910 74440 -21889
rect 75946 -21902 76066 -21889
rect 76126 -21902 76198 -21889
rect 74081 -21911 74440 -21910
rect 76032 -21910 76033 -21902
rect 76305 -21910 76391 -21889
rect 76966 -21890 77931 -21888
rect 77209 -21903 77329 -21890
rect 77389 -21903 77461 -21890
rect 76032 -21911 76391 -21910
rect 77295 -21911 77296 -21903
rect 77568 -21911 77654 -21890
rect 79209 -21895 79329 -21881
rect 79339 -21882 79678 -21881
rect 79389 -21895 79461 -21882
rect 79295 -21903 79296 -21895
rect 79568 -21903 79654 -21882
rect 82449 -21888 82894 -21817
rect 83533 -21888 83978 -21817
rect 85484 -21888 85929 -21817
rect 86780 -21818 87192 -21804
rect 88780 -21810 89192 -21796
rect 86747 -21881 87192 -21818
rect 88747 -21881 89192 -21810
rect 86747 -21883 89416 -21881
rect 82279 -21890 84255 -21888
rect 85241 -21890 86206 -21888
rect 86747 -21889 87192 -21883
rect 82449 -21903 82569 -21890
rect 82629 -21903 82701 -21890
rect 79295 -21904 79654 -21903
rect 77295 -21912 77654 -21911
rect 82535 -21911 82536 -21903
rect 82808 -21911 82894 -21890
rect 83533 -21903 83653 -21890
rect 83713 -21903 83785 -21890
rect 82535 -21912 82894 -21911
rect 83619 -21911 83620 -21903
rect 83892 -21911 83978 -21890
rect 85484 -21903 85604 -21890
rect 85664 -21903 85736 -21890
rect 83619 -21912 83978 -21911
rect 85570 -21911 85571 -21903
rect 85843 -21911 85929 -21890
rect 86504 -21891 87469 -21889
rect 86747 -21904 86867 -21891
rect 86927 -21904 86999 -21891
rect 85570 -21912 85929 -21911
rect 86833 -21912 86834 -21904
rect 87106 -21912 87192 -21891
rect 88747 -21896 88867 -21883
rect 88927 -21896 88999 -21883
rect 88833 -21904 88834 -21896
rect 89106 -21904 89192 -21883
rect 88833 -21905 89192 -21904
rect 86833 -21913 87192 -21912
rect 37683 -21925 38042 -21924
rect 35683 -21933 36042 -21932
rect 6912 -22041 7324 -22027
rect 6879 -22088 7324 -22041
rect 8081 -22088 8408 -22017
rect 9175 -22041 9587 -22027
rect 10407 -22041 10819 -22027
rect 9142 -22088 9587 -22041
rect 6879 -22090 9587 -22088
rect 6879 -22112 7324 -22090
rect 8167 -22112 8168 -22090
rect 8212 -22103 8284 -22090
rect 8225 -22108 8235 -22103
rect 8271 -22108 8281 -22107
rect 8235 -22112 8321 -22108
rect 8322 -22112 8408 -22090
rect 9142 -22112 9587 -22090
rect 10374 -22088 10819 -22041
rect 11576 -22088 11903 -22017
rect 12670 -22041 13082 -22027
rect 13996 -22041 14408 -22027
rect 12637 -22088 13082 -22041
rect 10374 -22090 13082 -22088
rect 10374 -22112 10819 -22090
rect 11662 -22112 11663 -22090
rect 11707 -22103 11779 -22090
rect 11720 -22108 11730 -22103
rect 11766 -22108 11776 -22107
rect 11730 -22112 11816 -22108
rect 11817 -22112 11903 -22090
rect 12637 -22112 13082 -22090
rect 13963 -22088 14408 -22041
rect 15165 -22088 15492 -22017
rect 58062 -22021 58474 -22007
rect 16259 -22041 16671 -22027
rect 16226 -22088 16671 -22041
rect 13963 -22090 16671 -22088
rect 13963 -22112 14408 -22090
rect 15251 -22112 15252 -22090
rect 15296 -22103 15368 -22090
rect 15309 -22108 15319 -22103
rect 15355 -22108 15365 -22107
rect 15319 -22112 15405 -22108
rect 15406 -22112 15492 -22090
rect 16226 -22112 16671 -22090
rect 58029 -22068 58474 -22021
rect 59231 -22068 59558 -21997
rect 60325 -22021 60737 -22007
rect 61557 -22021 61969 -22007
rect 60292 -22068 60737 -22021
rect 58029 -22070 60737 -22068
rect 58029 -22092 58474 -22070
rect 59317 -22092 59318 -22070
rect 59362 -22083 59434 -22070
rect 59375 -22088 59385 -22083
rect 59421 -22088 59431 -22087
rect 59385 -22092 59471 -22088
rect 59472 -22092 59558 -22070
rect 60292 -22092 60737 -22070
rect 61524 -22068 61969 -22021
rect 62726 -22068 63053 -21997
rect 63820 -22021 64232 -22007
rect 65146 -22021 65558 -22007
rect 63787 -22068 64232 -22021
rect 61524 -22070 64232 -22068
rect 61524 -22092 61969 -22070
rect 62812 -22092 62813 -22070
rect 62857 -22083 62929 -22070
rect 62870 -22088 62880 -22083
rect 62916 -22088 62926 -22087
rect 62880 -22092 62966 -22088
rect 62967 -22092 63053 -22070
rect 63787 -22092 64232 -22070
rect 65113 -22068 65558 -22021
rect 66315 -22068 66642 -21997
rect 67409 -22021 67821 -22007
rect 67376 -22068 67821 -22021
rect 65113 -22070 67821 -22068
rect 65113 -22092 65558 -22070
rect 66401 -22092 66402 -22070
rect 66446 -22083 66518 -22070
rect 66459 -22088 66469 -22083
rect 66505 -22088 66515 -22087
rect 66469 -22092 66555 -22088
rect 66556 -22092 66642 -22070
rect 67376 -22092 67821 -22070
rect 57431 -22094 68098 -22092
rect 58029 -22107 58149 -22094
rect 58209 -22107 58281 -22094
rect 6281 -22114 16948 -22112
rect 6879 -22127 6999 -22114
rect 7059 -22127 7131 -22114
rect 6965 -22135 6966 -22127
rect 7238 -22135 7324 -22114
rect 8167 -22120 8168 -22114
rect 8235 -22120 8321 -22114
rect 8322 -22120 8408 -22114
rect 8167 -22121 8408 -22120
rect 9142 -22127 9262 -22114
rect 9322 -22127 9394 -22114
rect 6965 -22136 7324 -22135
rect 9228 -22135 9229 -22127
rect 9501 -22135 9587 -22114
rect 10374 -22127 10494 -22114
rect 10554 -22127 10626 -22114
rect 9228 -22136 9587 -22135
rect 10460 -22135 10461 -22127
rect 10733 -22135 10819 -22114
rect 11662 -22120 11663 -22114
rect 11730 -22120 11816 -22114
rect 11817 -22120 11903 -22114
rect 11662 -22121 11903 -22120
rect 12637 -22127 12757 -22114
rect 12817 -22127 12889 -22114
rect 10460 -22136 10819 -22135
rect 12723 -22135 12724 -22127
rect 12996 -22135 13082 -22114
rect 13963 -22127 14083 -22114
rect 14143 -22127 14215 -22114
rect 12723 -22136 13082 -22135
rect 14049 -22135 14050 -22127
rect 14322 -22135 14408 -22114
rect 15251 -22120 15252 -22114
rect 15319 -22120 15405 -22114
rect 15406 -22120 15492 -22114
rect 15251 -22121 15492 -22120
rect 16226 -22127 16346 -22114
rect 16406 -22127 16478 -22114
rect 14049 -22136 14408 -22135
rect 16312 -22135 16313 -22127
rect 16585 -22135 16671 -22114
rect 58115 -22115 58116 -22107
rect 58388 -22115 58474 -22094
rect 59317 -22100 59318 -22094
rect 59385 -22100 59471 -22094
rect 59472 -22100 59558 -22094
rect 59317 -22101 59558 -22100
rect 60292 -22107 60412 -22094
rect 60472 -22107 60544 -22094
rect 58115 -22116 58474 -22115
rect 60378 -22115 60379 -22107
rect 60651 -22115 60737 -22094
rect 61524 -22107 61644 -22094
rect 61704 -22107 61776 -22094
rect 60378 -22116 60737 -22115
rect 61610 -22115 61611 -22107
rect 61883 -22115 61969 -22094
rect 62812 -22100 62813 -22094
rect 62880 -22100 62966 -22094
rect 62967 -22100 63053 -22094
rect 62812 -22101 63053 -22100
rect 63787 -22107 63907 -22094
rect 63967 -22107 64039 -22094
rect 61610 -22116 61969 -22115
rect 63873 -22115 63874 -22107
rect 64146 -22115 64232 -22094
rect 65113 -22107 65233 -22094
rect 65293 -22107 65365 -22094
rect 63873 -22116 64232 -22115
rect 65199 -22115 65200 -22107
rect 65472 -22115 65558 -22094
rect 66401 -22100 66402 -22094
rect 66469 -22100 66555 -22094
rect 66556 -22100 66642 -22094
rect 66401 -22101 66642 -22100
rect 67376 -22107 67496 -22094
rect 67556 -22107 67628 -22094
rect 65199 -22116 65558 -22115
rect 67462 -22115 67463 -22107
rect 67735 -22115 67821 -22094
rect 67462 -22116 67821 -22115
rect 16312 -22136 16671 -22135
rect 23809 -24048 24254 -23962
rect 23895 -24070 23896 -24048
rect 24015 -24057 24061 -24048
rect 24168 -24056 24254 -24048
rect 24874 -24056 25319 -23970
rect 27023 -24048 27468 -23962
rect 24135 -24057 24254 -24056
rect 24002 -24070 24074 -24057
rect 24135 -24070 24221 -24057
rect 23532 -24072 24497 -24070
rect 24015 -24084 24028 -24072
rect 24048 -24078 24061 -24072
rect 24960 -24078 24961 -24056
rect 25080 -24065 25126 -24056
rect 25233 -24064 25319 -24056
rect 25200 -24065 25319 -24064
rect 25067 -24078 25139 -24065
rect 25200 -24078 25286 -24065
rect 27109 -24070 27110 -24048
rect 27229 -24057 27275 -24048
rect 27382 -24056 27468 -24048
rect 28131 -24056 28576 -23970
rect 33347 -24049 33792 -23963
rect 27349 -24057 27468 -24056
rect 27216 -24070 27288 -24057
rect 27349 -24070 27435 -24057
rect 28217 -24070 28218 -24056
rect 28337 -24065 28383 -24056
rect 28490 -24064 28576 -24056
rect 28457 -24065 28576 -24064
rect 28324 -24070 28396 -24065
rect 26746 -24072 28396 -24070
rect 27229 -24078 27242 -24072
rect 24048 -24080 27242 -24078
rect 24048 -24084 24061 -24080
rect 25080 -24092 25093 -24080
rect 25113 -24092 25126 -24080
rect 27229 -24084 27242 -24080
rect 27262 -24078 27275 -24072
rect 28217 -24078 28218 -24072
rect 28324 -24078 28396 -24072
rect 28457 -24078 28543 -24065
rect 33433 -24071 33434 -24049
rect 33553 -24058 33599 -24049
rect 33706 -24057 33792 -24049
rect 34412 -24057 34857 -23971
rect 36561 -24049 37006 -23963
rect 33673 -24058 33792 -24057
rect 33540 -24071 33612 -24058
rect 33673 -24071 33759 -24058
rect 33070 -24073 34035 -24071
rect 27262 -24080 28616 -24078
rect 27262 -24084 27275 -24080
rect 28337 -24092 28350 -24080
rect 28370 -24092 28383 -24080
rect 33553 -24085 33566 -24073
rect 33586 -24079 33599 -24073
rect 34498 -24079 34499 -24057
rect 34618 -24066 34664 -24057
rect 34771 -24065 34857 -24057
rect 34738 -24066 34857 -24065
rect 34605 -24079 34677 -24066
rect 34738 -24079 34824 -24066
rect 36647 -24071 36648 -24049
rect 36767 -24058 36813 -24049
rect 36920 -24057 37006 -24049
rect 37669 -24057 38114 -23971
rect 74959 -24028 75404 -23942
rect 75045 -24050 75046 -24028
rect 75165 -24037 75211 -24028
rect 75318 -24036 75404 -24028
rect 76024 -24036 76469 -23950
rect 78173 -24028 78618 -23942
rect 75285 -24037 75404 -24036
rect 75152 -24050 75224 -24037
rect 75285 -24050 75371 -24037
rect 74682 -24052 75647 -24050
rect 36887 -24058 37006 -24057
rect 36754 -24071 36826 -24058
rect 36887 -24071 36973 -24058
rect 37755 -24071 37756 -24057
rect 37875 -24066 37921 -24057
rect 38028 -24065 38114 -24057
rect 75165 -24064 75178 -24052
rect 75198 -24058 75211 -24052
rect 76110 -24058 76111 -24036
rect 76230 -24045 76276 -24036
rect 76383 -24044 76469 -24036
rect 76350 -24045 76469 -24044
rect 76217 -24058 76289 -24045
rect 76350 -24058 76436 -24045
rect 78259 -24050 78260 -24028
rect 78379 -24037 78425 -24028
rect 78532 -24036 78618 -24028
rect 79281 -24036 79726 -23950
rect 84497 -24029 84942 -23943
rect 78499 -24037 78618 -24036
rect 78366 -24050 78438 -24037
rect 78499 -24050 78585 -24037
rect 79367 -24050 79368 -24036
rect 79487 -24045 79533 -24036
rect 79640 -24044 79726 -24036
rect 79607 -24045 79726 -24044
rect 79474 -24050 79546 -24045
rect 77896 -24052 79546 -24050
rect 78379 -24058 78392 -24052
rect 75198 -24060 78392 -24058
rect 75198 -24064 75211 -24060
rect 37995 -24066 38114 -24065
rect 37862 -24071 37934 -24066
rect 36284 -24073 37934 -24071
rect 36767 -24079 36780 -24073
rect 33586 -24081 36780 -24079
rect 33586 -24085 33599 -24081
rect 34618 -24093 34631 -24081
rect 34651 -24093 34664 -24081
rect 36767 -24085 36780 -24081
rect 36800 -24079 36813 -24073
rect 37755 -24079 37756 -24073
rect 37862 -24079 37934 -24073
rect 37995 -24079 38081 -24066
rect 76230 -24072 76243 -24060
rect 76263 -24072 76276 -24060
rect 78379 -24064 78392 -24060
rect 78412 -24058 78425 -24052
rect 79367 -24058 79368 -24052
rect 79474 -24058 79546 -24052
rect 79607 -24058 79693 -24045
rect 84583 -24051 84584 -24029
rect 84703 -24038 84749 -24029
rect 84856 -24037 84942 -24029
rect 85562 -24037 86007 -23951
rect 87711 -24029 88156 -23943
rect 84823 -24038 84942 -24037
rect 84690 -24051 84762 -24038
rect 84823 -24051 84909 -24038
rect 84220 -24053 85185 -24051
rect 78412 -24060 79766 -24058
rect 78412 -24064 78425 -24060
rect 79487 -24072 79500 -24060
rect 79520 -24072 79533 -24060
rect 84703 -24065 84716 -24053
rect 84736 -24059 84749 -24053
rect 85648 -24059 85649 -24037
rect 85768 -24046 85814 -24037
rect 85921 -24045 86007 -24037
rect 85888 -24046 86007 -24045
rect 85755 -24059 85827 -24046
rect 85888 -24059 85974 -24046
rect 87797 -24051 87798 -24029
rect 87917 -24038 87963 -24029
rect 88070 -24037 88156 -24029
rect 88819 -24037 89264 -23951
rect 88037 -24038 88156 -24037
rect 87904 -24051 87976 -24038
rect 88037 -24051 88123 -24038
rect 88905 -24051 88906 -24037
rect 89025 -24046 89071 -24037
rect 89178 -24045 89264 -24037
rect 89145 -24046 89264 -24045
rect 89012 -24051 89084 -24046
rect 87434 -24053 89084 -24051
rect 87917 -24059 87930 -24053
rect 84736 -24061 87930 -24059
rect 84736 -24065 84749 -24061
rect 85768 -24073 85781 -24061
rect 85801 -24073 85814 -24061
rect 87917 -24065 87930 -24061
rect 87950 -24059 87963 -24053
rect 88905 -24059 88906 -24053
rect 89012 -24059 89084 -24053
rect 89145 -24059 89231 -24046
rect 87950 -24061 89422 -24059
rect 87950 -24065 87963 -24061
rect 89025 -24073 89038 -24061
rect 89058 -24073 89071 -24061
rect 36800 -24081 38272 -24079
rect 36800 -24085 36813 -24081
rect 37875 -24093 37888 -24081
rect 37908 -24093 37921 -24081
rect 6861 -25551 7306 -25465
rect 6947 -25559 6948 -25551
rect 6947 -25560 6980 -25559
rect 7054 -25560 7100 -25551
rect 6980 -25573 6981 -25560
rect 7041 -25573 7113 -25560
rect 7220 -25573 7306 -25551
rect 8063 -25566 8390 -25480
rect 9124 -25551 9569 -25465
rect 10356 -25551 10801 -25465
rect 9210 -25559 9211 -25551
rect 9210 -25560 9243 -25559
rect 9317 -25560 9363 -25551
rect 8149 -25573 8150 -25566
rect 8207 -25573 8303 -25566
rect 8304 -25573 8390 -25566
rect 9243 -25573 9244 -25560
rect 9304 -25573 9376 -25560
rect 9483 -25573 9569 -25551
rect 10442 -25559 10443 -25551
rect 10442 -25560 10475 -25559
rect 10549 -25560 10595 -25551
rect 10475 -25573 10476 -25560
rect 10536 -25573 10608 -25560
rect 10715 -25573 10801 -25551
rect 11558 -25566 11885 -25480
rect 12619 -25551 13064 -25465
rect 13843 -25551 14288 -25465
rect 12705 -25559 12706 -25551
rect 12705 -25560 12738 -25559
rect 12812 -25560 12858 -25551
rect 11644 -25573 11645 -25566
rect 11702 -25573 11798 -25566
rect 11799 -25573 11885 -25566
rect 12738 -25573 12739 -25560
rect 12799 -25573 12871 -25560
rect 12978 -25573 13064 -25551
rect 13929 -25559 13930 -25551
rect 13929 -25560 13962 -25559
rect 14036 -25560 14082 -25551
rect 13962 -25573 13963 -25560
rect 14023 -25573 14095 -25560
rect 14202 -25573 14288 -25551
rect 15045 -25566 15372 -25480
rect 16106 -25551 16551 -25465
rect 17494 -25551 17939 -25465
rect 16192 -25559 16193 -25551
rect 16192 -25560 16225 -25559
rect 16299 -25560 16345 -25551
rect 15131 -25573 15132 -25566
rect 15189 -25573 15285 -25566
rect 15286 -25573 15372 -25566
rect 16225 -25573 16226 -25560
rect 16286 -25573 16358 -25560
rect 16465 -25573 16551 -25551
rect 17580 -25559 17581 -25551
rect 17580 -25560 17613 -25559
rect 17687 -25560 17733 -25551
rect 17613 -25573 17614 -25560
rect 17674 -25573 17746 -25560
rect 17853 -25573 17939 -25551
rect 18696 -25566 19023 -25480
rect 19757 -25551 20202 -25465
rect 24325 -25551 24770 -25465
rect 58011 -25531 58456 -25445
rect 58097 -25539 58098 -25531
rect 58097 -25540 58130 -25539
rect 58204 -25540 58250 -25531
rect 19843 -25559 19844 -25551
rect 19843 -25560 19876 -25559
rect 19950 -25560 19996 -25551
rect 18782 -25573 18783 -25566
rect 18840 -25573 18936 -25566
rect 18937 -25573 19023 -25566
rect 19876 -25573 19877 -25560
rect 19937 -25573 20009 -25560
rect 20116 -25573 20202 -25551
rect 24411 -25559 24412 -25551
rect 24411 -25560 24444 -25559
rect 24518 -25560 24564 -25551
rect 24444 -25573 24445 -25560
rect 24505 -25573 24577 -25560
rect 24684 -25573 24770 -25551
rect 58130 -25553 58131 -25540
rect 58191 -25553 58263 -25540
rect 58370 -25553 58456 -25531
rect 59213 -25546 59540 -25460
rect 60274 -25531 60719 -25445
rect 61506 -25531 61951 -25445
rect 60360 -25539 60361 -25531
rect 60360 -25540 60393 -25539
rect 60467 -25540 60513 -25531
rect 59299 -25553 59300 -25546
rect 59357 -25553 59453 -25546
rect 59454 -25553 59540 -25546
rect 60393 -25553 60394 -25540
rect 60454 -25553 60526 -25540
rect 60633 -25553 60719 -25531
rect 61592 -25539 61593 -25531
rect 61592 -25540 61625 -25539
rect 61699 -25540 61745 -25531
rect 61625 -25553 61626 -25540
rect 61686 -25553 61758 -25540
rect 61865 -25553 61951 -25531
rect 62708 -25546 63035 -25460
rect 63769 -25531 64214 -25445
rect 64993 -25531 65438 -25445
rect 63855 -25539 63856 -25531
rect 63855 -25540 63888 -25539
rect 63962 -25540 64008 -25531
rect 62794 -25553 62795 -25546
rect 62852 -25553 62948 -25546
rect 62949 -25553 63035 -25546
rect 63888 -25553 63889 -25540
rect 63949 -25553 64021 -25540
rect 64128 -25553 64214 -25531
rect 65079 -25539 65080 -25531
rect 65079 -25540 65112 -25539
rect 65186 -25540 65232 -25531
rect 65112 -25553 65113 -25540
rect 65173 -25553 65245 -25540
rect 65352 -25553 65438 -25531
rect 66195 -25546 66522 -25460
rect 67256 -25531 67701 -25445
rect 68644 -25531 69089 -25445
rect 67342 -25539 67343 -25531
rect 67342 -25540 67375 -25539
rect 67449 -25540 67495 -25531
rect 66281 -25553 66282 -25546
rect 66339 -25553 66435 -25546
rect 66436 -25553 66522 -25546
rect 67375 -25553 67376 -25540
rect 67436 -25553 67508 -25540
rect 67615 -25553 67701 -25531
rect 68730 -25539 68731 -25531
rect 68730 -25540 68763 -25539
rect 68837 -25540 68883 -25531
rect 68763 -25553 68764 -25540
rect 68824 -25553 68896 -25540
rect 69003 -25553 69089 -25531
rect 69846 -25546 70173 -25460
rect 70907 -25531 71352 -25445
rect 75475 -25531 75920 -25445
rect 70993 -25539 70994 -25531
rect 70993 -25540 71026 -25539
rect 71100 -25540 71146 -25531
rect 69932 -25553 69933 -25546
rect 69990 -25553 70086 -25546
rect 70087 -25553 70173 -25546
rect 71026 -25553 71027 -25540
rect 71087 -25553 71159 -25540
rect 71266 -25553 71352 -25531
rect 75561 -25539 75562 -25531
rect 75561 -25540 75594 -25539
rect 75668 -25540 75714 -25531
rect 75594 -25553 75595 -25540
rect 75655 -25553 75727 -25540
rect 75834 -25553 75920 -25531
rect 57431 -25555 76197 -25553
rect 58204 -25567 58217 -25555
rect 58237 -25567 58250 -25555
rect 6281 -25575 25047 -25573
rect 7054 -25587 7067 -25575
rect 7087 -25587 7100 -25575
rect 8149 -25597 8150 -25575
rect 8207 -25579 8303 -25575
rect 8207 -25584 8253 -25579
rect 8194 -25597 8266 -25584
rect 8304 -25597 8390 -25575
rect 9317 -25587 9330 -25575
rect 9350 -25587 9363 -25575
rect 10549 -25587 10562 -25575
rect 10582 -25587 10595 -25575
rect 11644 -25597 11645 -25575
rect 11702 -25579 11798 -25575
rect 11702 -25584 11748 -25579
rect 11689 -25597 11761 -25584
rect 11799 -25597 11885 -25575
rect 12812 -25587 12825 -25575
rect 12845 -25587 12858 -25575
rect 14036 -25587 14049 -25575
rect 14069 -25587 14082 -25575
rect 15131 -25597 15132 -25575
rect 15189 -25579 15285 -25575
rect 15189 -25584 15235 -25579
rect 15176 -25597 15248 -25584
rect 15286 -25597 15372 -25575
rect 16299 -25587 16312 -25575
rect 16332 -25587 16345 -25575
rect 17687 -25587 17700 -25575
rect 17720 -25587 17733 -25575
rect 18782 -25597 18783 -25575
rect 18840 -25579 18936 -25575
rect 18840 -25584 18886 -25579
rect 18827 -25597 18899 -25584
rect 18937 -25597 19023 -25575
rect 19950 -25587 19963 -25575
rect 19983 -25587 19996 -25575
rect 24518 -25587 24531 -25575
rect 24551 -25587 24564 -25575
rect 59299 -25577 59300 -25555
rect 59357 -25559 59453 -25555
rect 59357 -25564 59403 -25559
rect 59344 -25577 59416 -25564
rect 59454 -25577 59540 -25555
rect 60467 -25567 60480 -25555
rect 60500 -25567 60513 -25555
rect 61699 -25567 61712 -25555
rect 61732 -25567 61745 -25555
rect 62794 -25577 62795 -25555
rect 62852 -25559 62948 -25555
rect 62852 -25564 62898 -25559
rect 62839 -25577 62911 -25564
rect 62949 -25577 63035 -25555
rect 63962 -25567 63975 -25555
rect 63995 -25567 64008 -25555
rect 65186 -25567 65199 -25555
rect 65219 -25567 65232 -25555
rect 66281 -25577 66282 -25555
rect 66339 -25559 66435 -25555
rect 66339 -25564 66385 -25559
rect 66326 -25577 66398 -25564
rect 66436 -25577 66522 -25555
rect 67449 -25567 67462 -25555
rect 67482 -25567 67495 -25555
rect 68837 -25567 68850 -25555
rect 68870 -25567 68883 -25555
rect 69932 -25577 69933 -25555
rect 69990 -25559 70086 -25555
rect 69990 -25564 70036 -25559
rect 69977 -25577 70049 -25564
rect 70087 -25577 70173 -25555
rect 71100 -25567 71113 -25555
rect 71133 -25567 71146 -25555
rect 75668 -25567 75681 -25555
rect 75701 -25567 75714 -25555
rect 58250 -25579 60467 -25577
rect 61745 -25579 63962 -25577
rect 65232 -25579 67449 -25577
rect 68883 -25579 71100 -25577
rect 59357 -25591 59370 -25579
rect 59390 -25591 59403 -25579
rect 62852 -25591 62865 -25579
rect 62885 -25591 62898 -25579
rect 66339 -25591 66352 -25579
rect 66372 -25591 66385 -25579
rect 69990 -25591 70003 -25579
rect 70023 -25591 70036 -25579
rect 7100 -25599 9317 -25597
rect 10595 -25599 12812 -25597
rect 14082 -25599 16299 -25597
rect 17733 -25599 19950 -25597
rect 8207 -25611 8220 -25599
rect 8240 -25611 8253 -25599
rect 11702 -25611 11715 -25599
rect 11735 -25611 11748 -25599
rect 15189 -25611 15202 -25599
rect 15222 -25611 15235 -25599
rect 18840 -25611 18853 -25599
rect 18873 -25611 18886 -25599
<< nwell >>
rect 8578 11491 8995 11493
rect 8561 11488 8995 11491
<< metal1 >>
rect 18808 63061 19203 63067
rect -3079 62798 -2804 62816
rect -3079 62746 -3050 62798
rect -2998 62796 -2804 62798
rect -2998 62746 -2886 62796
rect -3079 62744 -2886 62746
rect -2834 62744 -2804 62796
rect -3079 62684 -2804 62744
rect -3079 62677 -2884 62684
rect -3390 62671 -2884 62677
rect -3390 62619 -3050 62671
rect -2998 62632 -2884 62671
rect -2832 62632 -2804 62684
rect -2998 62619 -2804 62632
rect -3390 62549 -2804 62619
rect -3079 62544 -2804 62549
rect -3079 62533 -2879 62544
rect -3079 62481 -3050 62533
rect -2998 62492 -2879 62533
rect -2827 62492 -2804 62544
rect -2998 62481 -2804 62492
rect -3079 62466 -2804 62481
rect -1982 62677 19203 63061
rect -4059 61402 -3689 61414
rect -4411 61370 -3689 61402
rect -4411 61357 -3843 61370
rect -4411 61305 -4009 61357
rect -3957 61318 -3843 61357
rect -3791 61318 -3689 61370
rect -3957 61305 -3689 61318
rect -4411 61237 -3689 61305
rect -4059 61230 -3689 61237
rect -4059 61219 -3838 61230
rect -4059 61167 -4009 61219
rect -3957 61178 -3838 61219
rect -3786 61178 -3689 61230
rect -3957 61167 -3689 61178
rect -4059 61136 -3689 61167
rect -2698 52726 -2423 52744
rect -2698 52674 -2669 52726
rect -2617 52724 -2423 52726
rect -2617 52674 -2505 52724
rect -2698 52672 -2505 52674
rect -2453 52672 -2423 52724
rect -2698 52639 -2423 52672
rect -3477 52612 -2423 52639
rect -3477 52599 -2503 52612
rect -3477 52547 -2669 52599
rect -2617 52560 -2503 52599
rect -2451 52560 -2423 52612
rect -2617 52547 -2423 52560
rect -3477 52491 -2423 52547
rect -2698 52472 -2423 52491
rect -2698 52461 -2498 52472
rect -2698 52409 -2669 52461
rect -2617 52420 -2498 52461
rect -2446 52420 -2423 52472
rect -2617 52409 -2423 52420
rect -2698 52394 -2423 52409
rect -3907 52246 -3537 52258
rect -4131 52214 -3537 52246
rect -4131 52201 -3691 52214
rect -4131 52149 -3857 52201
rect -3805 52162 -3691 52201
rect -3639 52162 -3537 52214
rect -3805 52149 -3537 52162
rect -4131 52081 -3537 52149
rect -3907 52074 -3537 52081
rect -3907 52063 -3686 52074
rect -3907 52011 -3857 52063
rect -3805 52022 -3686 52063
rect -3634 52022 -3537 52074
rect -3805 52011 -3537 52022
rect -3907 51980 -3537 52011
rect -2388 44200 -2113 44218
rect -2388 44148 -2359 44200
rect -2307 44198 -2113 44200
rect -2307 44148 -2195 44198
rect -2388 44146 -2195 44148
rect -2143 44146 -2113 44198
rect -2388 44086 -2113 44146
rect -2388 44073 -2193 44086
rect -3246 44021 -2359 44073
rect -2307 44034 -2193 44073
rect -2141 44034 -2113 44086
rect -2307 44021 -2113 44034
rect -3246 43946 -2113 44021
rect -3246 43935 -2188 43946
rect -3246 43925 -2359 43935
rect -2388 43883 -2359 43925
rect -2307 43894 -2188 43935
rect -2136 43894 -2113 43946
rect -2307 43883 -2113 43894
rect -2388 43868 -2113 43883
rect -2381 43659 -2106 43677
rect -2381 43607 -2352 43659
rect -2300 43657 -2106 43659
rect -2300 43607 -2188 43657
rect -2381 43605 -2188 43607
rect -2136 43605 -2106 43657
rect -2381 43547 -2106 43605
rect -3246 43545 -2106 43547
rect -3246 43532 -2186 43545
rect -3246 43480 -2352 43532
rect -2300 43493 -2186 43532
rect -2134 43493 -2106 43545
rect -2300 43480 -2106 43493
rect -3246 43405 -2106 43480
rect -3246 43399 -2181 43405
rect -2381 43394 -2181 43399
rect -2381 43342 -2352 43394
rect -2300 43353 -2181 43394
rect -2129 43353 -2106 43405
rect -2300 43342 -2106 43353
rect -2381 43327 -2106 43342
rect -2489 36766 -2214 36784
rect -2489 36714 -2460 36766
rect -2408 36764 -2214 36766
rect -2408 36714 -2296 36764
rect -2489 36712 -2296 36714
rect -2244 36712 -2214 36764
rect -2489 36680 -2214 36712
rect -3157 36652 -2214 36680
rect -3157 36639 -2294 36652
rect -3157 36587 -2460 36639
rect -2408 36600 -2294 36639
rect -2242 36600 -2214 36652
rect -2408 36587 -2214 36600
rect -3157 36532 -2214 36587
rect -2489 36512 -2214 36532
rect -2489 36501 -2289 36512
rect -2489 36449 -2460 36501
rect -2408 36460 -2289 36501
rect -2237 36460 -2214 36512
rect -2408 36449 -2214 36460
rect -2489 36434 -2214 36449
rect -3588 25040 -3261 25051
rect -3588 24988 -3571 25040
rect -3519 24988 -3451 25040
rect -3399 24988 -3331 25040
rect -3279 24988 -3261 25040
rect -3588 24965 -3261 24988
rect -3896 24920 -3261 24965
rect -3896 24868 -3571 24920
rect -3519 24868 -3451 24920
rect -3399 24868 -3331 24920
rect -3279 24868 -3261 24920
rect -3896 24824 -3261 24868
rect -3588 24800 -3261 24824
rect -3588 24748 -3571 24800
rect -3519 24748 -3451 24800
rect -3399 24748 -3331 24800
rect -3279 24748 -3261 24800
rect -3588 24732 -3261 24748
rect -1982 24212 -1598 62677
rect -734 55462 -180 55520
rect 4523 55463 5059 55511
rect 2762 54729 2988 54776
rect 8386 54369 8903 54424
rect -1113 48238 -1066 48601
rect 7285 41464 7336 42465
rect 7526 40566 7997 40618
rect 61 39776 236 39866
rect 4351 39720 4955 39766
rect 2010 28025 2740 28118
rect 2010 28017 2609 28025
rect 2010 27965 2043 28017
rect 2095 28014 2419 28017
rect 2095 27965 2222 28014
rect 2010 27962 2222 27965
rect 2274 27965 2419 28014
rect 2471 27973 2609 28017
rect 2661 27973 2740 28025
rect 2471 27965 2740 27973
rect 2274 27962 2740 27965
rect 2010 27890 2740 27962
rect 2010 27838 2046 27890
rect 2098 27882 2609 27890
rect 2098 27879 2411 27882
rect 2098 27838 2222 27879
rect 2010 27827 2222 27838
rect 2274 27830 2411 27879
rect 2463 27838 2609 27882
rect 2661 27838 2740 27890
rect 2463 27830 2740 27838
rect 2274 27827 2740 27830
rect 2010 27720 2740 27827
rect 5020 26011 5999 26363
rect -1982 24059 -1230 24212
rect -1982 23938 -1598 24059
rect -1383 23938 -1230 24059
rect -1982 23785 -806 23938
rect -1982 22452 -1598 23785
rect 5647 23168 5999 26011
rect 2715 22816 11131 23168
rect 18808 22570 19203 62677
rect 18790 22452 19220 22570
rect -1982 22068 19220 22452
rect 18790 21990 19220 22068
rect 9800 17596 10310 17660
rect 9800 17544 9836 17596
rect 9888 17544 9964 17596
rect 10016 17593 10310 17596
rect 10016 17544 10115 17593
rect 9800 17541 10115 17544
rect 10167 17541 10310 17593
rect 9800 17482 10310 17541
rect 7638 17437 10310 17482
rect 7638 17385 9834 17437
rect 9886 17435 10181 17437
rect 9886 17385 10005 17435
rect 7638 17383 10005 17385
rect 10057 17385 10181 17435
rect 10233 17385 10310 17437
rect 10057 17383 10310 17385
rect 7638 17338 10310 17383
rect 7638 16685 7782 17338
rect 9800 17274 10310 17338
rect 9800 17258 10197 17274
rect 9800 17253 10048 17258
rect 9800 17201 9846 17253
rect 9898 17206 10048 17253
rect 10100 17222 10197 17258
rect 10249 17222 10310 17274
rect 10100 17206 10310 17222
rect 9898 17201 10310 17206
rect 9800 17160 10310 17201
rect 13355 17337 25065 18084
rect 4098 16541 7782 16685
rect 9750 16933 10260 16990
rect 9750 16926 10054 16933
rect 9750 16923 9923 16926
rect 9750 16871 9795 16923
rect 9847 16874 9923 16923
rect 9975 16881 10054 16926
rect 10106 16881 10260 16933
rect 9975 16874 10260 16881
rect 9847 16871 10260 16874
rect 9750 16749 10260 16871
rect 9750 16744 10107 16749
rect 9750 16726 9959 16744
rect 9750 16674 9790 16726
rect 9842 16692 9959 16726
rect 10011 16697 10107 16744
rect 10159 16697 10260 16749
rect 10011 16692 10260 16697
rect 9842 16674 10260 16692
rect 9750 16616 10260 16674
rect 9750 16606 10141 16616
rect 9750 16575 9964 16606
rect 9750 16523 9767 16575
rect 9819 16554 9964 16575
rect 10016 16564 10141 16606
rect 10193 16564 10260 16616
rect 10016 16554 10260 16564
rect 9819 16523 10260 16554
rect 9750 16490 10260 16523
rect 1520 15970 1593 16058
rect 1320 15880 1398 15964
rect 1740 15510 1998 15563
rect 1863 15507 1996 15510
rect 9778 15355 9980 16490
rect 1530 15295 2126 15296
rect 1530 15240 2128 15295
rect 1532 15239 2128 15240
rect 3928 15153 9980 15355
rect 11733 14403 11992 14405
rect 2167 13969 7519 14172
rect 5930 11533 6133 13969
rect 6482 11515 6685 13969
rect 7316 11533 7519 13969
rect 9781 13966 11992 14403
rect 9781 11862 10218 13966
rect 11532 13843 11992 13966
rect 13355 13958 14102 17337
rect 22731 16826 23374 16880
rect 22731 16802 22815 16826
rect 22672 16774 22815 16802
rect 22867 16774 22935 16826
rect 22987 16774 23055 16826
rect 23107 16774 23175 16826
rect 23227 16774 23295 16826
rect 23347 16774 23374 16826
rect 22672 16706 23374 16774
rect 22672 16654 22815 16706
rect 22867 16654 22935 16706
rect 22987 16654 23055 16706
rect 23107 16654 23175 16706
rect 23227 16654 23295 16706
rect 23347 16654 23374 16706
rect 22672 16626 23374 16654
rect 22731 16591 23374 16626
rect 22735 16431 23393 16495
rect 22735 16430 22822 16431
rect 22669 16379 22822 16430
rect 22874 16379 22942 16431
rect 22994 16379 23062 16431
rect 23114 16379 23182 16431
rect 23234 16379 23302 16431
rect 23354 16379 23393 16431
rect 22669 16311 23393 16379
rect 22669 16259 22822 16311
rect 22874 16259 22942 16311
rect 22994 16259 23062 16311
rect 23114 16259 23182 16311
rect 23234 16259 23302 16311
rect 23354 16259 23393 16311
rect 22669 16232 23393 16259
rect 22735 16213 23393 16232
rect 22738 16210 23393 16213
rect 24318 16043 25065 17337
rect 55673 16043 56135 16047
rect 24318 15847 67173 16043
rect 67680 15847 88740 15857
rect 24318 15482 88740 15847
rect 24318 15472 68127 15482
rect 24318 15296 67173 15472
rect 22079 15270 22652 15272
rect 21918 15250 22652 15270
rect 21918 15198 22094 15250
rect 22146 15198 22214 15250
rect 22266 15198 22334 15250
rect 22386 15198 22454 15250
rect 22506 15198 22574 15250
rect 22626 15198 22652 15250
rect 21918 15130 22652 15198
rect 21918 15078 22094 15130
rect 22146 15078 22214 15130
rect 22266 15078 22334 15130
rect 22386 15078 22454 15130
rect 22506 15078 22574 15130
rect 22626 15078 22652 15130
rect 21918 15051 22652 15078
rect 21918 15049 22491 15051
rect 55490 14890 56420 15296
rect 22045 14662 22661 14694
rect 21999 14632 22694 14662
rect 21999 14580 22063 14632
rect 22115 14580 22183 14632
rect 22235 14580 22303 14632
rect 22355 14580 22423 14632
rect 22475 14580 22543 14632
rect 22595 14580 22694 14632
rect 21999 14512 22694 14580
rect 21999 14470 22063 14512
rect 17927 14293 18154 14470
rect 22045 14460 22063 14470
rect 22115 14460 22183 14512
rect 22235 14460 22303 14512
rect 22355 14460 22423 14512
rect 22475 14460 22543 14512
rect 22595 14470 22694 14512
rect 22595 14460 22661 14470
rect 22045 14427 22661 14460
rect 17890 14268 18200 14293
rect 17890 14008 17931 14268
rect 18191 14008 18200 14268
rect 19228 14168 19380 14254
rect 10844 13450 11116 13516
rect 10844 13398 10858 13450
rect 10910 13398 10996 13450
rect 11048 13398 11116 13450
rect 10844 13323 11116 13398
rect 10844 13271 10861 13323
rect 10913 13321 11116 13323
rect 10913 13271 11000 13321
rect 10844 13269 11000 13271
rect 11052 13269 11116 13321
rect 10844 13252 11116 13269
rect 10844 13212 11222 13252
rect 12351 13241 12512 13253
rect 10844 13179 11335 13212
rect 12222 13195 12512 13241
rect 12351 13184 12512 13195
rect 10844 13170 11000 13179
rect 10844 13118 10860 13170
rect 10912 13127 11000 13170
rect 11052 13140 11335 13179
rect 11052 13127 11222 13140
rect 10912 13118 11222 13127
rect 10844 13100 11222 13118
rect 11365 12706 11683 12801
rect 11365 12654 11401 12706
rect 11453 12703 11683 12706
rect 11453 12654 11585 12703
rect 11365 12651 11585 12654
rect 11637 12651 11683 12703
rect 11365 12578 11683 12651
rect 11365 12526 11398 12578
rect 11450 12570 11683 12578
rect 11450 12526 11583 12570
rect 11365 12518 11583 12526
rect 11635 12518 11683 12570
rect 11365 12433 11683 12518
rect 12387 12469 12512 13184
rect 11365 12381 11399 12433
rect 11451 12381 11576 12433
rect 11628 12381 11683 12433
rect 11365 12334 11683 12381
rect 12257 12415 12529 12469
rect 12257 12363 12271 12415
rect 12323 12363 12409 12415
rect 12461 12363 12529 12415
rect 12257 12288 12529 12363
rect 12257 12236 12274 12288
rect 12326 12286 12529 12288
rect 12326 12236 12413 12286
rect 12257 12234 12413 12236
rect 12465 12234 12529 12286
rect 12257 12217 12529 12234
rect 12257 12144 12533 12217
rect 12257 12135 12413 12144
rect 12257 12083 12273 12135
rect 12325 12092 12413 12135
rect 12465 12092 12533 12144
rect 12325 12083 12533 12092
rect 12257 12065 12533 12083
rect 8578 11665 8995 11731
rect 8578 11662 8876 11665
rect 8578 11661 8731 11662
rect 8578 11609 8609 11661
rect 8661 11610 8731 11661
rect 8783 11613 8876 11662
rect 8928 11613 8995 11665
rect 8783 11610 8995 11613
rect 8661 11609 8995 11610
rect 8578 11550 8995 11609
rect 9781 11564 12433 11862
rect 8578 11549 8746 11550
rect 8578 11497 8615 11549
rect 8667 11498 8746 11549
rect 8798 11498 8885 11550
rect 8937 11498 8995 11550
rect 8667 11497 8995 11498
rect 8578 11491 8995 11497
rect 9959 11492 12433 11564
rect 8561 11488 8995 11491
rect 1646 10690 2266 10779
rect 2407 10345 2529 10437
rect -63 7610 319 10120
rect 11236 9990 11632 10070
rect 11236 9979 11521 9990
rect 11236 9927 11344 9979
rect 11396 9938 11521 9979
rect 11573 9938 11632 9990
rect 11396 9927 11632 9938
rect 11236 9858 11632 9927
rect 11236 9848 11414 9858
rect 11236 9796 11278 9848
rect 11330 9806 11414 9848
rect 11466 9853 11632 9858
rect 11466 9806 11561 9853
rect 11330 9801 11561 9806
rect 11613 9801 11632 9853
rect 11330 9796 11632 9801
rect 11236 9772 11632 9796
rect 4086 9217 5247 9311
rect 12063 8509 12433 11492
rect 11423 7982 11671 8029
rect 11423 7930 11440 7982
rect 11492 7930 11574 7982
rect 11626 7930 11671 7982
rect 11423 7894 11671 7930
rect 12747 7909 13129 7920
rect 11423 7874 11740 7894
rect 11423 7868 11837 7874
rect 11423 7816 11435 7868
rect 11487 7856 11837 7868
rect 11487 7816 11564 7856
rect 11423 7804 11564 7816
rect 11616 7804 11837 7856
rect 12692 7851 13129 7909
rect 11423 7802 11837 7804
rect 11423 7782 11740 7802
rect 12747 7798 13129 7851
rect 11423 7781 11671 7782
rect 5268 7610 6063 7709
rect -63 7564 6063 7610
rect -63 7560 5731 7564
rect -63 7544 5592 7560
rect -63 7492 5395 7544
rect 5447 7508 5592 7544
rect 5644 7512 5731 7560
rect 5783 7560 6063 7564
rect 5783 7512 5875 7560
rect 5644 7508 5875 7512
rect 5927 7508 6063 7560
rect 5447 7492 6063 7508
rect -63 7440 6063 7492
rect -63 7426 5854 7440
rect -63 7419 5680 7426
rect -63 7414 5507 7419
rect -63 7362 5358 7414
rect 5410 7367 5507 7414
rect 5559 7374 5680 7419
rect 5732 7388 5854 7426
rect 5906 7388 6063 7440
rect 5732 7374 6063 7388
rect 5559 7367 6063 7374
rect 5410 7362 6063 7367
rect -63 7311 6063 7362
rect 10683 7569 11112 7726
rect 10683 7355 11727 7569
rect 10753 7354 11727 7355
rect 13007 7311 13129 7798
rect -63 7306 5943 7311
rect -63 7302 5641 7306
rect -63 7294 5478 7302
rect -63 7242 5327 7294
rect 5379 7250 5478 7294
rect 5530 7254 5641 7302
rect 5693 7254 5802 7306
rect 5854 7259 5943 7306
rect 5995 7259 6063 7311
rect 5854 7254 6063 7259
rect 5530 7250 6063 7254
rect 5379 7242 6063 7250
rect -63 7228 6063 7242
rect 5268 7226 6063 7228
rect 12940 7305 13192 7311
rect 12940 7253 12966 7305
rect 13018 7253 13102 7305
rect 13154 7253 13192 7305
rect 12940 7192 13192 7253
rect 12940 7140 12961 7192
rect 13013 7185 13192 7192
rect 13013 7140 13097 7185
rect 8560 7073 9108 7137
rect 12940 7133 13097 7140
rect 13149 7133 13192 7185
rect 12940 7111 13192 7133
rect 8560 7068 8953 7073
rect 8560 7016 8598 7068
rect 8650 7016 8741 7068
rect 8793 7021 8953 7068
rect 9005 7021 9108 7073
rect 8793 7016 9108 7021
rect 8560 6956 9108 7016
rect 8560 6904 8598 6956
rect 8650 6904 8746 6956
rect 8798 6904 8984 6956
rect 9036 6904 9108 6956
rect 8560 6879 9108 6904
rect 12397 5486 12483 5488
rect 12397 5403 12791 5486
rect 12397 5392 12679 5403
rect 12397 5340 12502 5392
rect 12554 5351 12679 5392
rect 12731 5351 12791 5403
rect 12554 5340 12791 5351
rect 12397 5271 12791 5340
rect 12397 5261 12572 5271
rect 12397 5209 12436 5261
rect 12488 5219 12572 5261
rect 12624 5266 12791 5271
rect 12624 5219 12719 5266
rect 12488 5214 12719 5219
rect 12771 5214 12791 5266
rect 12488 5209 12791 5214
rect 12397 5185 12791 5209
rect 5586 4579 6428 4675
rect 4778 -990 5148 -932
rect 4778 -1042 4828 -990
rect 4880 -992 5148 -990
rect 4880 -1042 4992 -992
rect 4778 -1044 4992 -1042
rect 5044 -1044 5148 -992
rect 4778 -1072 5148 -1044
rect 4422 -1104 5148 -1072
rect 4422 -1117 4994 -1104
rect 4422 -1169 4828 -1117
rect 4880 -1156 4994 -1117
rect 5046 -1156 5148 -1104
rect 4880 -1169 5148 -1156
rect 4422 -1237 5148 -1169
rect 4778 -1244 5148 -1237
rect 4778 -1255 4999 -1244
rect 4778 -1307 4828 -1255
rect 4880 -1296 4999 -1255
rect 5051 -1296 5148 -1244
rect 4880 -1307 5148 -1296
rect 4778 -1338 5148 -1307
rect 4844 -1524 5214 -1512
rect 4488 -1556 5214 -1524
rect 4488 -1569 5060 -1556
rect 4488 -1621 4894 -1569
rect 4946 -1608 5060 -1569
rect 5112 -1608 5214 -1556
rect 4946 -1621 5214 -1608
rect 4488 -1689 5214 -1621
rect 4844 -1696 5214 -1689
rect 4844 -1707 5065 -1696
rect 4844 -1759 4894 -1707
rect 4946 -1748 5065 -1707
rect 5117 -1748 5214 -1696
rect 4946 -1759 5214 -1748
rect 4844 -1790 5214 -1759
rect 4506 -2253 4874 -2240
rect 4506 -2305 4796 -2253
rect 4848 -2305 4874 -2253
rect 4506 -2330 4874 -2305
rect 4377 -2356 4874 -2330
rect 4377 -2408 4547 -2356
rect 4599 -2408 4687 -2356
rect 4739 -2408 4874 -2356
rect 4377 -2441 4874 -2408
rect 4506 -2477 4874 -2441
rect 4506 -2529 4549 -2477
rect 4601 -2480 4874 -2477
rect 4601 -2529 4695 -2480
rect 4506 -2532 4695 -2529
rect 4747 -2485 4874 -2480
rect 4747 -2532 4815 -2485
rect 4506 -2537 4815 -2532
rect 4867 -2537 4874 -2485
rect 4506 -2563 4874 -2537
rect 5001 -2620 5371 -2608
rect 4645 -2652 5371 -2620
rect 4645 -2665 5217 -2652
rect 4645 -2717 5051 -2665
rect 5103 -2704 5217 -2665
rect 5269 -2704 5371 -2652
rect 5103 -2717 5371 -2704
rect 4645 -2785 5371 -2717
rect 5001 -2792 5371 -2785
rect 5001 -2803 5222 -2792
rect 5001 -2855 5051 -2803
rect 5103 -2844 5222 -2803
rect 5274 -2844 5371 -2792
rect 5103 -2855 5371 -2844
rect 5001 -2886 5371 -2855
rect 4905 -3038 5275 -3026
rect 4549 -3070 5275 -3038
rect 4549 -3083 5121 -3070
rect 4549 -3135 4955 -3083
rect 5007 -3122 5121 -3083
rect 5173 -3122 5275 -3070
rect 5007 -3135 5275 -3122
rect 4549 -3203 5275 -3135
rect 4905 -3210 5275 -3203
rect 4905 -3221 5126 -3210
rect 4905 -3273 4955 -3221
rect 5007 -3262 5126 -3221
rect 5178 -3262 5275 -3210
rect 5007 -3273 5275 -3262
rect 4905 -3304 5275 -3273
rect 4882 -3452 5252 -3440
rect 4526 -3484 5252 -3452
rect 4526 -3497 5098 -3484
rect 4526 -3549 4932 -3497
rect 4984 -3536 5098 -3497
rect 5150 -3536 5252 -3484
rect 4984 -3549 5252 -3536
rect 4526 -3617 5252 -3549
rect 4882 -3624 5252 -3617
rect 4882 -3635 5103 -3624
rect 4882 -3687 4932 -3635
rect 4984 -3676 5103 -3635
rect 5155 -3676 5252 -3624
rect 4984 -3687 5252 -3676
rect 4882 -3718 5252 -3687
rect 4928 -3931 5298 -3919
rect 4572 -3963 5298 -3931
rect 4572 -3976 5144 -3963
rect 4572 -4028 4978 -3976
rect 5030 -4015 5144 -3976
rect 5196 -4015 5298 -3963
rect 5030 -4028 5298 -4015
rect 4572 -4096 5298 -4028
rect 4928 -4103 5298 -4096
rect 4928 -4114 5149 -4103
rect 4928 -4166 4978 -4114
rect 5030 -4155 5149 -4114
rect 5201 -4155 5298 -4103
rect 5030 -4166 5298 -4155
rect 4928 -4197 5298 -4166
rect 5033 -4474 5403 -4462
rect 4677 -4506 5403 -4474
rect 4677 -4519 5249 -4506
rect 4677 -4571 5083 -4519
rect 5135 -4558 5249 -4519
rect 5301 -4558 5403 -4506
rect 5135 -4571 5403 -4558
rect 4677 -4639 5403 -4571
rect 5033 -4646 5403 -4639
rect 5033 -4657 5254 -4646
rect 5033 -4709 5083 -4657
rect 5135 -4698 5254 -4657
rect 5306 -4698 5403 -4646
rect 5135 -4709 5403 -4698
rect 5033 -4740 5403 -4709
rect 5638 -5420 5862 -5418
rect 8579 -5420 9022 3070
rect 9531 -5420 9974 3070
rect 10350 -5420 10793 3070
rect 13382 -3641 14075 13958
rect 17890 13943 18200 14008
rect 17890 13787 17919 13943
rect 18179 13787 18200 13943
rect 17890 13738 18200 13787
rect 19198 14114 19410 14168
rect 20406 14143 20600 14210
rect 28009 14158 45862 14382
rect 20393 14129 20705 14143
rect 19198 13750 19222 14114
rect 19378 13750 19410 14114
rect 20370 14091 20705 14129
rect 20370 13831 20393 14091
rect 20653 13831 20705 14091
rect 22087 14087 23144 14135
rect 21918 14084 23144 14087
rect 21918 13928 22116 14084
rect 22272 13928 22498 14084
rect 22654 13928 22917 14084
rect 23073 13928 23144 14084
rect 21918 13926 23144 13928
rect 22087 13904 23144 13926
rect 28009 14106 37935 14158
rect 37987 14106 38055 14158
rect 38107 14106 38175 14158
rect 38227 14106 38295 14158
rect 38347 14106 38415 14158
rect 38467 14106 45862 14158
rect 28009 14038 45862 14106
rect 28009 13986 37935 14038
rect 37987 13986 38055 14038
rect 38107 13986 38175 14038
rect 38227 13986 38295 14038
rect 38347 13986 38415 14038
rect 38467 13986 45862 14038
rect 28009 13917 45862 13986
rect 20370 13811 20705 13831
rect 19198 13738 19410 13750
rect 21938 13658 22849 13700
rect 21833 13616 22849 13658
rect 21833 13564 22006 13616
rect 22058 13564 22429 13616
rect 22481 13564 22720 13616
rect 22772 13564 22849 13616
rect 21833 13522 22849 13564
rect 21938 13497 22849 13522
rect 21781 13239 22530 13292
rect 21781 13187 21838 13239
rect 21890 13187 22077 13239
rect 22129 13187 22410 13239
rect 22462 13187 22530 13239
rect 21781 13142 22530 13187
rect 28009 13000 28474 13917
rect 29826 13325 30426 13389
rect 29826 13323 29830 13325
rect 29802 13273 29830 13323
rect 29882 13273 29950 13325
rect 30002 13273 30070 13325
rect 30122 13273 30190 13325
rect 30242 13273 30310 13325
rect 30362 13323 30426 13325
rect 30362 13273 31638 13323
rect 29802 13205 31638 13273
rect 29802 13153 29830 13205
rect 29882 13153 29950 13205
rect 30002 13153 30070 13205
rect 30122 13153 30190 13205
rect 30242 13153 30310 13205
rect 30362 13153 31638 13205
rect 29802 13134 31638 13153
rect 28009 12882 28470 13000
rect 22767 12489 24077 12615
rect 25831 12525 28470 12882
rect 22767 12487 23800 12489
rect 22767 12486 23246 12487
rect 22823 12412 22947 12486
rect 23122 12412 23246 12486
rect 23406 12412 23530 12487
rect 23676 12412 23800 12487
rect 23953 12412 24077 12489
rect 25830 12503 28470 12525
rect 25830 12433 26744 12503
rect 24624 12412 24967 12413
rect 25540 12412 25770 12413
rect 25830 12412 26545 12433
rect 16702 12108 17532 12110
rect 16702 11903 18051 12108
rect 22793 11960 26545 12412
rect 16702 11653 17532 11903
rect 16702 11448 18065 11653
rect 26224 11549 26277 11586
rect 16702 11170 17532 11448
rect 22449 11211 22560 11220
rect 19654 11188 19738 11204
rect 16702 10965 18065 11170
rect 19654 11136 19670 11188
rect 19722 11136 19738 11188
rect 19654 11121 19738 11136
rect 19895 11193 19979 11209
rect 19895 11141 19911 11193
rect 19963 11141 19979 11193
rect 19895 11126 19979 11141
rect 20134 11195 20218 11211
rect 20134 11143 20150 11195
rect 20202 11143 20218 11195
rect 20134 11139 20218 11143
rect 20206 11128 20218 11139
rect 20361 11195 20445 11211
rect 20361 11143 20377 11195
rect 20429 11143 20445 11195
rect 20361 11128 20445 11143
rect 22449 11167 22956 11211
rect 22449 11115 22481 11167
rect 22533 11115 22956 11167
rect 22449 11110 22956 11115
rect 22449 11023 22560 11110
rect 22449 10971 22476 11023
rect 22528 10971 22560 11023
rect 16702 10715 17532 10965
rect 22449 10942 22560 10971
rect 16702 10510 18070 10715
rect 16702 9691 17532 10510
rect 20845 10390 21011 10561
rect 21224 10390 21390 10578
rect 21511 10390 21677 10561
rect 20845 10386 21677 10390
rect 21966 10388 22132 10574
rect 21966 10386 23117 10388
rect 20845 10224 23117 10386
rect 21511 10222 23117 10224
rect 31449 10181 31638 13134
rect 31886 11708 32351 13917
rect 44097 13154 44562 13917
rect 44130 13150 44562 13154
rect 45397 13145 45862 13917
rect 64769 13772 65603 13916
rect 64769 13720 64929 13772
rect 64981 13768 65603 13772
rect 64981 13720 65188 13768
rect 64769 13718 65188 13720
rect 47691 13716 65188 13718
rect 65240 13716 65603 13768
rect 47691 13703 65603 13716
rect 47691 13651 65429 13703
rect 65481 13651 65603 13703
rect 47691 13621 65603 13651
rect 47691 13569 64933 13621
rect 64985 13591 65603 13621
rect 64985 13569 65200 13591
rect 47691 13539 65200 13569
rect 65252 13550 65603 13591
rect 65252 13539 65424 13550
rect 47691 13498 65424 13539
rect 65476 13498 65603 13550
rect 47691 13454 65603 13498
rect 47691 13452 65190 13454
rect 47691 13400 64932 13452
rect 64984 13402 65190 13452
rect 65242 13407 65603 13454
rect 65242 13402 65422 13407
rect 64984 13400 65422 13402
rect 47691 13355 65422 13400
rect 65474 13355 65603 13407
rect 47691 13277 65603 13355
rect 47691 13225 64982 13277
rect 65034 13272 65603 13277
rect 65034 13225 65184 13272
rect 47691 13220 65184 13225
rect 65236 13260 65603 13272
rect 65236 13220 65347 13260
rect 47691 13208 65347 13220
rect 65399 13208 65603 13260
rect 47691 13149 65603 13208
rect 41677 12634 41885 12734
rect 41677 12582 41755 12634
rect 41807 12582 41885 12634
rect 41677 12384 41885 12582
rect 41677 12332 41755 12384
rect 41807 12332 41885 12384
rect 41677 12214 41885 12332
rect 41677 12160 42058 12214
rect 41677 12108 41755 12160
rect 41807 12108 42058 12160
rect 41677 12061 42058 12108
rect 37793 10784 38571 10840
rect 37793 10732 37877 10784
rect 37929 10732 37997 10784
rect 38049 10732 38117 10784
rect 38169 10732 38237 10784
rect 38289 10732 38357 10784
rect 38409 10732 38571 10784
rect 37793 10664 38571 10732
rect 37793 10612 37877 10664
rect 37929 10612 37997 10664
rect 38049 10612 38117 10664
rect 38169 10612 38237 10664
rect 38289 10612 38357 10664
rect 38409 10612 38571 10664
rect 37793 10547 38571 10612
rect 19888 9897 22600 10122
rect 31449 10073 32313 10181
rect 31449 9975 31638 10073
rect 28770 9909 28848 9964
rect 29009 9914 29087 9964
rect 29248 9916 29326 9964
rect 29474 9916 29552 9964
rect 16702 9264 17980 9691
rect 22373 9505 22600 9897
rect 28768 9893 28852 9909
rect 28768 9841 28784 9893
rect 28836 9841 28852 9893
rect 28768 9826 28852 9841
rect 29009 9898 29093 9914
rect 29009 9846 29025 9898
rect 29077 9846 29093 9898
rect 29009 9831 29093 9846
rect 29248 9900 29332 9916
rect 29248 9848 29264 9900
rect 29316 9848 29332 9900
rect 29248 9833 29332 9848
rect 29474 9900 29559 9916
rect 29474 9848 29491 9900
rect 29543 9848 29559 9900
rect 29474 9833 29559 9848
rect 28770 9794 28848 9826
rect 29009 9794 29087 9831
rect 29248 9794 29326 9833
rect 29474 9794 29552 9833
rect 22373 9472 22743 9505
rect 22373 9390 22985 9472
rect 22373 9358 22743 9390
rect 16702 8606 17532 9264
rect 19614 9158 19692 9209
rect 19853 9163 19931 9209
rect 20318 9165 20396 9209
rect 19612 9142 19696 9158
rect 19612 9090 19628 9142
rect 19680 9090 19696 9142
rect 19612 9075 19696 9090
rect 19853 9147 19937 9163
rect 19853 9095 19869 9147
rect 19921 9095 19937 9147
rect 19853 9080 19937 9095
rect 20092 9149 20176 9153
rect 20092 9097 20108 9149
rect 20160 9097 20176 9149
rect 20092 9082 20176 9097
rect 20318 9149 20403 9165
rect 20318 9097 20335 9149
rect 20387 9097 20403 9149
rect 20318 9082 20403 9097
rect 19614 9039 19692 9075
rect 19853 9039 19931 9080
rect 20092 9039 20170 9082
rect 20318 9039 20396 9082
rect 26167 8889 26249 8932
rect 16702 8179 18037 8606
rect 27648 8585 27807 9468
rect 27901 8593 28060 9476
rect 28305 8593 28464 9476
rect 28660 8589 28819 9472
rect 30473 8717 30883 9048
rect 26351 8450 26523 8578
rect 16702 4973 17532 8179
rect 22865 7922 22989 8384
rect 23323 7922 23447 8384
rect 24418 7922 24542 8396
rect 25281 7922 25405 8393
rect 25975 7922 26099 8413
rect 26224 8326 26523 8450
rect 26343 8324 26523 8326
rect 26351 7922 26523 8324
rect 22840 7881 26523 7922
rect 22840 7879 23419 7881
rect 22840 7874 23180 7879
rect 22840 7822 22939 7874
rect 22991 7827 23180 7874
rect 23232 7829 23419 7879
rect 23471 7829 23646 7881
rect 23698 7829 26523 7881
rect 23232 7827 26523 7829
rect 22991 7822 26523 7827
rect 22840 7798 26523 7822
rect 26351 7706 26523 7798
rect 18490 7270 18630 7520
rect 28714 6915 28792 6970
rect 28953 6920 29031 6970
rect 29192 6922 29270 6970
rect 29418 6922 29496 6970
rect 28712 6899 28796 6915
rect 17937 6751 18038 6809
rect 22095 6791 22546 6850
rect 28712 6847 28728 6899
rect 28780 6847 28796 6899
rect 28712 6832 28796 6847
rect 28953 6904 29037 6920
rect 28953 6852 28969 6904
rect 29021 6852 29037 6904
rect 28953 6837 29037 6852
rect 29192 6906 29276 6922
rect 29192 6854 29208 6906
rect 29260 6854 29276 6906
rect 29192 6839 29276 6854
rect 29418 6906 29503 6922
rect 29418 6854 29435 6906
rect 29487 6854 29503 6906
rect 29418 6839 29503 6854
rect 28714 6800 28792 6832
rect 28953 6800 29031 6837
rect 29192 6800 29270 6839
rect 29418 6800 29496 6839
rect 21988 6789 22546 6791
rect 17937 6711 19507 6751
rect 21988 6737 22134 6789
rect 22186 6737 22430 6789
rect 22482 6737 22546 6789
rect 17937 6670 19508 6711
rect 21988 6705 22546 6737
rect 22085 6683 22546 6705
rect 17937 6646 18072 6670
rect 17938 6618 18072 6646
rect 18124 6618 18192 6670
rect 18244 6618 18312 6670
rect 18364 6618 18432 6670
rect 18484 6618 18552 6670
rect 18604 6618 18672 6670
rect 18724 6618 18792 6670
rect 18844 6618 18912 6670
rect 18964 6618 19032 6670
rect 19084 6618 19152 6670
rect 19204 6618 19272 6670
rect 19324 6618 19392 6670
rect 19444 6618 19508 6670
rect 17938 6585 19508 6618
rect 26889 5053 27137 6444
rect 27452 5078 27700 6469
rect 27937 5086 28185 6477
rect 28962 6257 29078 6331
rect 31485 6257 31602 9975
rect 32011 9879 32303 9911
rect 32011 9827 32075 9879
rect 32127 9827 32303 9879
rect 32011 9792 32303 9827
rect 28962 6141 31602 6257
rect 33295 9275 33729 9309
rect 36032 9299 36466 10247
rect 36737 9299 37171 10223
rect 36032 9275 37171 9299
rect 33295 8865 37171 9275
rect 33295 8841 36466 8865
rect 32225 5373 32329 5795
rect 33295 5113 33729 8841
rect 47691 8256 48260 13149
rect 64769 13020 65603 13149
rect 55240 9830 56170 9840
rect 47615 8228 48260 8256
rect 47615 8176 47793 8228
rect 47845 8176 47949 8228
rect 48001 8176 48260 8228
rect 47615 8150 48260 8176
rect 47690 7940 48260 8150
rect 50084 9609 57840 9830
rect 50084 7719 50305 9609
rect 53921 9316 54794 9377
rect 53921 9315 54374 9316
rect 53921 9314 54252 9315
rect 53921 9262 54014 9314
rect 54066 9262 54133 9314
rect 54185 9263 54252 9314
rect 54304 9264 54374 9315
rect 54426 9315 54794 9316
rect 54426 9264 54492 9315
rect 54304 9263 54492 9264
rect 54544 9263 54794 9315
rect 54185 9262 54794 9263
rect 53921 9199 54794 9262
rect 53921 9197 54374 9199
rect 53921 9196 54254 9197
rect 53921 9144 54014 9196
rect 54066 9144 54133 9196
rect 54185 9145 54254 9196
rect 54306 9147 54374 9197
rect 54426 9195 54794 9199
rect 54426 9147 54493 9195
rect 54306 9145 54493 9147
rect 54185 9144 54493 9145
rect 53921 9143 54493 9144
rect 54545 9143 54794 9195
rect 53921 9088 54794 9143
rect 50084 7338 50292 7719
rect 43227 7112 43321 7123
rect 46153 7119 46241 7191
rect 46418 7119 46522 7199
rect 46706 7119 46809 7195
rect 46908 7119 47009 7188
rect 48084 7130 50292 7338
rect 57619 7531 57840 9609
rect 61491 9323 62361 9385
rect 61491 9322 61944 9323
rect 61491 9321 61822 9322
rect 61491 9269 61584 9321
rect 61636 9269 61703 9321
rect 61755 9270 61822 9321
rect 61874 9271 61944 9322
rect 61996 9322 62361 9323
rect 61996 9271 62062 9322
rect 61874 9270 62062 9271
rect 62114 9270 62361 9322
rect 61755 9269 62361 9270
rect 61491 9206 62361 9269
rect 61491 9204 61944 9206
rect 61491 9203 61824 9204
rect 61491 9151 61584 9203
rect 61636 9151 61703 9203
rect 61755 9152 61824 9203
rect 61876 9154 61944 9204
rect 61996 9202 62361 9206
rect 61996 9154 62063 9202
rect 61876 9152 62063 9154
rect 61755 9151 62063 9152
rect 61491 9150 62063 9151
rect 62115 9150 62361 9202
rect 61491 9099 62361 9150
rect 58049 7531 58270 8320
rect 66783 7933 67158 15296
rect 57619 7310 58270 7531
rect 43227 7111 43449 7112
rect 43820 7111 43992 7112
rect 43227 7104 44714 7111
rect 43227 6948 43285 7104
rect 43441 6948 43828 7104
rect 43984 6948 44538 7104
rect 44694 6948 44714 7104
rect 46136 7078 47059 7119
rect 46136 7073 46937 7078
rect 46136 7021 46195 7073
rect 46247 7070 46937 7073
rect 46247 7068 46721 7070
rect 46247 7021 46441 7068
rect 46136 7016 46441 7021
rect 46493 7018 46721 7068
rect 46773 7026 46937 7070
rect 46989 7026 47059 7078
rect 46773 7018 47059 7026
rect 46493 7016 47059 7018
rect 46136 6961 47059 7016
rect 43227 6941 44714 6948
rect 43227 6940 43449 6941
rect 43820 6940 43992 6941
rect 43227 6919 43321 6940
rect 38263 6633 39669 6671
rect 38263 6608 39913 6633
rect 38263 6452 39342 6608
rect 39498 6452 39913 6608
rect 38263 6430 39913 6452
rect 38287 6427 39913 6430
rect 38287 6418 39669 6427
rect 38287 6414 38493 6418
rect 43759 6074 44718 6127
rect 43759 6022 43825 6074
rect 43877 6061 44718 6074
rect 43877 6022 44074 6061
rect 43759 6009 44074 6022
rect 44126 6060 44718 6061
rect 44126 6056 44530 6060
rect 44126 6009 44308 6056
rect 43759 6004 44308 6009
rect 44360 6008 44530 6056
rect 44582 6008 44718 6060
rect 44360 6004 44718 6008
rect 43759 5971 44718 6004
rect 16702 4546 24378 4973
rect 40140 4953 42232 5122
rect 16702 3267 17532 4546
rect 21250 3267 21677 4546
rect 30400 4487 30604 4659
rect 27094 4405 27485 4463
rect 27094 4353 27149 4405
rect 27201 4353 27381 4405
rect 27433 4353 27485 4405
rect 27094 4209 27485 4353
rect 30400 4435 30470 4487
rect 30522 4435 30604 4487
rect 30400 4263 30604 4435
rect 27094 4157 27146 4209
rect 27198 4157 27381 4209
rect 27433 4157 27485 4209
rect 27094 4108 27485 4157
rect 30300 4226 30604 4263
rect 42800 4230 42910 4490
rect 30300 4174 30470 4226
rect 30522 4174 30604 4226
rect 43290 4210 43400 4470
rect 30300 4138 30604 4174
rect 30400 4129 30604 4138
rect 27110 3940 27240 4108
rect 16702 2840 24359 3267
rect 16702 1379 17532 2840
rect 21227 1379 21654 2840
rect 44729 2789 45104 4670
rect 48084 2343 48292 7130
rect 50084 6664 50292 7130
rect 56251 6721 56621 6792
rect 58049 6680 58270 7310
rect 66784 6887 67156 7933
rect 64336 6799 67156 6887
rect 64234 6728 67156 6799
rect 64336 6639 67156 6728
rect 66784 6577 67156 6639
rect 49311 5107 64328 5157
rect 48076 2220 48292 2343
rect 48596 4954 64328 5107
rect 48596 4904 49514 4954
rect 48596 1659 48799 4904
rect 49311 4006 49514 4904
rect 49799 4761 50002 4954
rect 51438 4912 51796 4954
rect 51593 4761 51796 4912
rect 49799 4558 51796 4761
rect 53695 4662 54568 4724
rect 53695 4661 54148 4662
rect 53695 4660 54026 4661
rect 53695 4608 53788 4660
rect 53840 4608 53907 4660
rect 53959 4609 54026 4660
rect 54078 4610 54148 4661
rect 54200 4661 54568 4662
rect 54200 4610 54266 4661
rect 54078 4609 54266 4610
rect 54318 4609 54568 4661
rect 53959 4608 54568 4609
rect 49799 4006 50002 4558
rect 53695 4545 54568 4608
rect 53695 4543 54148 4545
rect 53695 4542 54028 4543
rect 53695 4490 53788 4542
rect 53840 4490 53907 4542
rect 53959 4491 54028 4542
rect 54080 4493 54148 4543
rect 54200 4541 54568 4545
rect 54200 4493 54267 4541
rect 54080 4491 54267 4493
rect 53959 4490 54267 4491
rect 53695 4489 54267 4490
rect 54319 4489 54568 4541
rect 53695 4412 54568 4489
rect 53695 4319 54344 4412
rect 53701 4315 54344 4319
rect 53701 4314 54194 4315
rect 49311 3803 50002 4006
rect 49311 1659 49514 3803
rect 50335 2374 50478 3627
rect 47450 1456 49514 1659
rect 50081 2231 50478 2374
rect 16702 952 24382 1379
rect 47945 1007 48083 1256
rect 50081 1007 50224 2231
rect 50335 1992 50478 2231
rect 56403 2041 56855 2118
rect 16702 -1185 17532 952
rect 19771 -1203 20198 952
rect 47943 864 50224 1007
rect 50715 -448 51181 505
rect 52024 -448 52490 458
rect 53443 -448 53909 458
rect 54484 -448 54950 458
rect 74047 -448 74513 -207
rect 47429 -914 74513 -448
rect 88322 -822 88697 15482
rect 98848 4719 99160 4739
rect 98848 4667 98889 4719
rect 98941 4713 99160 4719
rect 98941 4667 99064 4713
rect 98848 4661 99064 4667
rect 99116 4661 99160 4713
rect 98848 4660 99160 4661
rect 98848 4564 99482 4660
rect 98848 4560 99065 4564
rect 98848 4508 98887 4560
rect 98939 4512 99065 4560
rect 99117 4512 99482 4564
rect 98939 4508 99482 4512
rect 98848 4440 99482 4508
rect 98848 4395 99160 4440
rect 98848 4343 98890 4395
rect 98942 4390 99160 4395
rect 98942 4343 99078 4390
rect 98848 4338 99078 4343
rect 99130 4338 99160 4390
rect 91327 4255 92059 4316
rect 98848 4305 99160 4338
rect 91327 4254 91780 4255
rect 91327 4253 91658 4254
rect 91327 4201 91420 4253
rect 91472 4201 91539 4253
rect 91591 4202 91658 4253
rect 91710 4203 91780 4254
rect 91832 4254 92059 4255
rect 91832 4203 91898 4254
rect 91710 4202 91898 4203
rect 91950 4202 92059 4254
rect 91591 4201 92059 4202
rect 91327 4138 92059 4201
rect 91327 4136 91780 4138
rect 91327 4135 91660 4136
rect 91327 4083 91420 4135
rect 91472 4083 91539 4135
rect 91591 4084 91660 4135
rect 91712 4086 91780 4136
rect 91832 4134 92059 4138
rect 91832 4086 91899 4134
rect 91712 4084 91899 4086
rect 91591 4083 91899 4084
rect 91327 4082 91899 4083
rect 91951 4082 92059 4134
rect 91327 4051 92059 4082
rect 95080 2666 95620 2970
rect 95080 2614 95236 2666
rect 95288 2614 95356 2666
rect 95408 2614 95476 2666
rect 95528 2614 95620 2666
rect 95080 2546 95620 2614
rect 95080 2494 95236 2546
rect 95288 2494 95356 2546
rect 95408 2494 95476 2546
rect 95528 2494 95620 2546
rect 95080 2426 95620 2494
rect 95080 2374 95236 2426
rect 95288 2374 95356 2426
rect 95408 2374 95476 2426
rect 95528 2374 95620 2426
rect 95080 2270 95620 2374
rect 90062 -69 90216 161
rect 90062 -223 91541 -69
rect 90062 -240 90357 -223
rect 89933 -302 90357 -240
rect 89933 -314 90131 -302
rect 89933 -366 90007 -314
rect 90059 -354 90131 -314
rect 90183 -354 90357 -302
rect 90059 -366 90357 -354
rect 89933 -410 90357 -366
rect 91387 -410 91541 -223
rect 93502 -410 93656 120
rect 89933 -431 93656 -410
rect 89933 -483 90025 -431
rect 90077 -443 93656 -431
rect 90077 -483 90149 -443
rect 89933 -495 90149 -483
rect 90201 -495 93656 -443
rect 89933 -564 93656 -495
rect 89933 -570 90316 -564
rect 50307 -915 50773 -914
rect 52557 -915 53023 -914
rect 55367 -915 55833 -914
rect 18080 -1534 18860 -1470
rect 18080 -1541 18702 -1534
rect 18080 -1546 18452 -1541
rect 18080 -1598 18145 -1546
rect 18197 -1593 18452 -1546
rect 18504 -1586 18702 -1541
rect 18754 -1586 18860 -1534
rect 18504 -1593 18860 -1586
rect 18197 -1598 18860 -1593
rect 18080 -1660 18860 -1598
rect 58411 -2964 58526 -2610
rect 58344 -3015 58612 -2964
rect 58344 -3040 58527 -3015
rect 58344 -3092 58357 -3040
rect 58409 -3067 58527 -3040
rect 58579 -3067 58612 -3015
rect 58409 -3092 58612 -3067
rect 58344 -3213 58612 -3092
rect 58344 -3214 58522 -3213
rect 58344 -3266 58356 -3214
rect 58408 -3265 58522 -3214
rect 58574 -3265 58612 -3213
rect 58408 -3266 58612 -3265
rect 58344 -3325 58612 -3266
rect 20040 -3641 20542 -3449
rect 13382 -3920 20542 -3641
rect 13382 -4128 14075 -3920
rect 60197 -5340 60663 -914
rect 64717 -5340 65183 -914
rect 66293 -5340 66759 -914
rect 68159 -3641 68520 -3628
rect 68159 -3693 68218 -3641
rect 68270 -3642 68520 -3641
rect 68270 -3693 68392 -3642
rect 68159 -3694 68392 -3693
rect 68444 -3694 68520 -3642
rect 68159 -3695 68520 -3694
rect 68159 -3807 69109 -3695
rect 68159 -3859 68219 -3807
rect 68271 -3810 69109 -3807
rect 68271 -3812 68520 -3810
rect 68271 -3859 68417 -3812
rect 68159 -3864 68417 -3859
rect 68469 -3864 68520 -3812
rect 68159 -3896 68520 -3864
rect 70747 -5340 71213 -914
rect 73441 -5340 73907 -914
rect 87273 -1197 88697 -822
rect 98561 -762 98873 -742
rect 98561 -814 98602 -762
rect 98654 -768 98873 -762
rect 98654 -814 98777 -768
rect 98561 -820 98777 -814
rect 98829 -820 98873 -768
rect 98561 -900 98873 -820
rect 98561 -917 99246 -900
rect 98561 -921 98778 -917
rect 98561 -973 98600 -921
rect 98652 -969 98778 -921
rect 98830 -969 99246 -917
rect 98652 -973 99246 -969
rect 98561 -1057 99246 -973
rect 98561 -1086 98873 -1057
rect 98561 -1138 98603 -1086
rect 98655 -1091 98873 -1086
rect 98655 -1138 98791 -1091
rect 98561 -1143 98791 -1138
rect 98843 -1143 98873 -1091
rect 98561 -1181 98873 -1143
rect 87273 -4550 87648 -1197
rect 98576 -1966 98937 -1953
rect 98576 -2018 98635 -1966
rect 98687 -1967 98937 -1966
rect 98687 -2018 98809 -1967
rect 98576 -2019 98809 -2018
rect 98861 -2019 98937 -1967
rect 98576 -2020 98937 -2019
rect 98576 -2132 99239 -2020
rect 98576 -2184 98636 -2132
rect 98688 -2135 99239 -2132
rect 98688 -2137 98937 -2135
rect 98688 -2184 98834 -2137
rect 98576 -2189 98834 -2184
rect 98886 -2189 98937 -2137
rect 98576 -2221 98937 -2189
rect 98546 -2863 98907 -2850
rect 98546 -2915 98605 -2863
rect 98657 -2864 98907 -2863
rect 98657 -2915 98779 -2864
rect 98546 -2916 98779 -2915
rect 98831 -2916 98907 -2864
rect 98546 -2917 98907 -2916
rect 98546 -3029 99209 -2917
rect 98546 -3081 98606 -3029
rect 98658 -3032 99209 -3029
rect 98658 -3034 98907 -3032
rect 98658 -3081 98804 -3034
rect 98546 -3086 98804 -3081
rect 98856 -3086 98907 -3034
rect 98546 -3118 98907 -3086
rect 98538 -3346 98899 -3333
rect 98538 -3398 98597 -3346
rect 98649 -3347 98899 -3346
rect 98649 -3398 98771 -3347
rect 98538 -3399 98771 -3398
rect 98823 -3399 98899 -3347
rect 98538 -3400 98899 -3399
rect 98538 -3512 99201 -3400
rect 98538 -3564 98598 -3512
rect 98650 -3515 99201 -3512
rect 98650 -3517 98899 -3515
rect 98650 -3564 98796 -3517
rect 98538 -3569 98796 -3564
rect 98848 -3569 98899 -3517
rect 98538 -3601 98899 -3569
rect 98576 -3898 98937 -3885
rect 98576 -3950 98635 -3898
rect 98687 -3899 98937 -3898
rect 98687 -3950 98809 -3899
rect 98576 -3951 98809 -3950
rect 98861 -3951 98937 -3899
rect 98576 -3952 98937 -3951
rect 98576 -4064 99239 -3952
rect 98576 -4116 98636 -4064
rect 98688 -4067 99239 -4064
rect 98688 -4069 98937 -4067
rect 98688 -4116 98834 -4069
rect 98576 -4121 98834 -4116
rect 98886 -4121 98937 -4069
rect 98576 -4153 98937 -4121
rect 87090 -4724 87760 -4550
rect 87090 -4776 87136 -4724
rect 87188 -4776 87256 -4724
rect 87308 -4776 87376 -4724
rect 87428 -4776 87760 -4724
rect 87090 -4844 87760 -4776
rect 87090 -4896 87136 -4844
rect 87188 -4896 87256 -4844
rect 87308 -4896 87376 -4844
rect 87428 -4896 87760 -4844
rect 87090 -4964 87760 -4896
rect 87090 -5016 87136 -4964
rect 87188 -5016 87256 -4964
rect 87308 -5016 87376 -4964
rect 87428 -5016 87760 -4964
rect 87090 -5090 87760 -5016
rect 5638 -5640 46550 -5420
rect 5638 -26120 5862 -5640
rect 46330 -7116 46550 -5640
rect 56830 -5580 97660 -5340
rect 56830 -7113 57070 -5580
rect 46330 -7305 49145 -7116
rect 6386 -8123 6433 -7467
rect 13089 -7874 13136 -7507
rect 28743 -7995 28833 -7665
rect 13833 -10333 13879 -9997
rect 13098 -12624 13146 -12186
rect 28843 -12493 28889 -11707
rect 25725 -14613 27275 -14562
rect 14185 -16057 14240 -15620
rect 27991 -15636 28043 -14884
rect 28905 -18073 28951 -17807
rect 42594 -18574 45406 -18222
rect 46330 -26120 46550 -7305
rect 54749 -7361 57070 -7113
rect 54726 -8904 56321 -8804
rect 48724 -9293 48793 -9131
rect 48405 -9341 48793 -9293
rect 48405 -9393 48446 -9341
rect 48498 -9353 48793 -9341
rect 48498 -9393 48585 -9353
rect 48405 -9405 48585 -9393
rect 48637 -9405 48793 -9353
rect 48405 -9457 48793 -9405
rect 48405 -9509 48440 -9457
rect 48492 -9478 48793 -9457
rect 48492 -9509 48588 -9478
rect 48405 -9530 48588 -9509
rect 48640 -9530 48793 -9478
rect 48405 -9571 48793 -9530
rect 48405 -9623 48443 -9571
rect 48495 -9594 48793 -9571
rect 48495 -9623 48588 -9594
rect 48405 -9646 48588 -9623
rect 48640 -9646 48793 -9594
rect 48405 -9663 48793 -9646
rect 48724 -10104 48793 -9663
rect 52279 -11322 53565 -11166
rect 52279 -11368 53571 -11322
rect 52279 -11371 53319 -11368
rect 52279 -11379 53077 -11371
rect 52279 -11381 52808 -11379
rect 52279 -11394 52553 -11381
rect 52279 -11446 52348 -11394
rect 52400 -11433 52553 -11394
rect 52605 -11431 52808 -11381
rect 52860 -11423 53077 -11379
rect 53129 -11420 53319 -11371
rect 53371 -11420 53571 -11368
rect 53129 -11423 53571 -11420
rect 52860 -11431 53571 -11423
rect 52605 -11433 53571 -11431
rect 52400 -11446 53571 -11433
rect 52279 -11550 53571 -11446
rect 52279 -11551 53406 -11550
rect 52279 -11563 53247 -11551
rect 52279 -11566 53034 -11563
rect 52279 -11576 52789 -11566
rect 52279 -11584 52556 -11576
rect 52279 -11636 52350 -11584
rect 52402 -11628 52556 -11584
rect 52608 -11618 52789 -11576
rect 52841 -11615 53034 -11566
rect 53086 -11603 53247 -11563
rect 53299 -11602 53406 -11551
rect 53458 -11602 53571 -11550
rect 53299 -11603 53571 -11602
rect 53086 -11615 53571 -11603
rect 52841 -11618 53571 -11615
rect 52608 -11628 53571 -11618
rect 52402 -11636 53571 -11628
rect 52279 -11736 53571 -11636
rect 52279 -11744 53355 -11736
rect 52279 -11754 53157 -11744
rect 52279 -11757 52918 -11754
rect 52279 -11759 52707 -11757
rect 52279 -11760 52509 -11759
rect 52279 -11812 52341 -11760
rect 52393 -11811 52509 -11760
rect 52561 -11809 52707 -11759
rect 52759 -11806 52918 -11757
rect 52970 -11796 53157 -11754
rect 53209 -11788 53355 -11744
rect 53407 -11788 53571 -11736
rect 53209 -11796 53571 -11788
rect 52970 -11806 53571 -11796
rect 52759 -11809 53571 -11806
rect 52561 -11811 53571 -11809
rect 52393 -11812 53571 -11811
rect 52279 -11848 53571 -11812
rect 48991 -14110 49554 -14074
rect 56118 -14110 56321 -8904
rect 48991 -14140 56322 -14110
rect 48789 -14156 56322 -14140
rect 48789 -14208 49199 -14156
rect 49251 -14208 49319 -14156
rect 49371 -14208 49439 -14156
rect 49491 -14208 56322 -14156
rect 48789 -14276 56322 -14208
rect 48789 -14328 49199 -14276
rect 49251 -14328 49319 -14276
rect 49371 -14328 49439 -14276
rect 49491 -14315 56322 -14276
rect 49491 -14328 49554 -14315
rect 48789 -14335 49554 -14328
rect 48991 -14450 49554 -14335
rect 5638 -26332 46550 -26120
rect 5780 -26340 46550 -26332
rect 56830 -26120 57070 -7361
rect 57536 -8443 57583 -7347
rect 64239 -8183 64286 -7477
rect 79893 -8205 79983 -7375
rect 64983 -10117 65030 -10037
rect 64983 -10164 65333 -10117
rect 64983 -10343 65030 -10164
rect 64248 -12534 64296 -11606
rect 79993 -12443 80039 -11737
rect 77165 -14593 77995 -14542
rect 65335 -15997 65390 -15493
rect 65336 -16516 65388 -15997
rect 79141 -16316 79193 -14894
rect 79617 -17833 80103 -17787
rect 80055 -18003 80101 -17833
rect 93784 -18554 96726 -18202
rect 97420 -26120 97660 -5580
rect 98574 -7474 98910 -7460
rect 98574 -7526 98606 -7474
rect 98658 -7526 98726 -7474
rect 98778 -7526 98846 -7474
rect 98898 -7526 98910 -7474
rect 98574 -7530 98910 -7526
rect 98574 -7594 99250 -7530
rect 98574 -7646 98606 -7594
rect 98658 -7646 98726 -7594
rect 98778 -7646 98846 -7594
rect 98898 -7646 99250 -7594
rect 98574 -7690 99250 -7646
rect 98574 -7714 98910 -7690
rect 98574 -7766 98606 -7714
rect 98658 -7766 98726 -7714
rect 98778 -7766 98846 -7714
rect 98898 -7766 98910 -7714
rect 98574 -7800 98910 -7766
rect 56830 -26360 97660 -26120
<< via1 >>
rect -3050 62746 -2998 62798
rect -2886 62744 -2834 62796
rect -3050 62619 -2998 62671
rect -2884 62632 -2832 62684
rect -3050 62481 -2998 62533
rect -2879 62492 -2827 62544
rect -4009 61305 -3957 61357
rect -3843 61318 -3791 61370
rect -4009 61167 -3957 61219
rect -3838 61178 -3786 61230
rect -2669 52674 -2617 52726
rect -2505 52672 -2453 52724
rect -2669 52547 -2617 52599
rect -2503 52560 -2451 52612
rect -2669 52409 -2617 52461
rect -2498 52420 -2446 52472
rect -3857 52149 -3805 52201
rect -3691 52162 -3639 52214
rect -3857 52011 -3805 52063
rect -3686 52022 -3634 52074
rect -2359 44148 -2307 44200
rect -2195 44146 -2143 44198
rect -2359 44021 -2307 44073
rect -2193 44034 -2141 44086
rect -2359 43883 -2307 43935
rect -2188 43894 -2136 43946
rect -2352 43607 -2300 43659
rect -2188 43605 -2136 43657
rect -2352 43480 -2300 43532
rect -2186 43493 -2134 43545
rect -2352 43342 -2300 43394
rect -2181 43353 -2129 43405
rect -2460 36714 -2408 36766
rect -2296 36712 -2244 36764
rect -2460 36587 -2408 36639
rect -2294 36600 -2242 36652
rect -2460 36449 -2408 36501
rect -2289 36460 -2237 36512
rect -3571 24988 -3519 25040
rect -3451 24988 -3399 25040
rect -3331 24988 -3279 25040
rect -3571 24868 -3519 24920
rect -3451 24868 -3399 24920
rect -3331 24868 -3279 24920
rect -3571 24748 -3519 24800
rect -3451 24748 -3399 24800
rect -3331 24748 -3279 24800
rect 2043 27965 2095 28017
rect 2222 27962 2274 28014
rect 2419 27965 2471 28017
rect 2609 27973 2661 28025
rect 2046 27838 2098 27890
rect 2222 27827 2274 27879
rect 2411 27830 2463 27882
rect 2609 27838 2661 27890
rect 9836 17544 9888 17596
rect 9964 17544 10016 17596
rect 10115 17541 10167 17593
rect 9834 17385 9886 17437
rect 10005 17383 10057 17435
rect 10181 17385 10233 17437
rect 9846 17201 9898 17253
rect 10048 17206 10100 17258
rect 10197 17222 10249 17274
rect 9795 16871 9847 16923
rect 9923 16874 9975 16926
rect 10054 16881 10106 16933
rect 9790 16674 9842 16726
rect 9959 16692 10011 16744
rect 10107 16697 10159 16749
rect 9767 16523 9819 16575
rect 9964 16554 10016 16606
rect 10141 16564 10193 16616
rect 22815 16774 22867 16826
rect 22935 16774 22987 16826
rect 23055 16774 23107 16826
rect 23175 16774 23227 16826
rect 23295 16774 23347 16826
rect 22815 16654 22867 16706
rect 22935 16654 22987 16706
rect 23055 16654 23107 16706
rect 23175 16654 23227 16706
rect 23295 16654 23347 16706
rect 22822 16379 22874 16431
rect 22942 16379 22994 16431
rect 23062 16379 23114 16431
rect 23182 16379 23234 16431
rect 23302 16379 23354 16431
rect 22822 16259 22874 16311
rect 22942 16259 22994 16311
rect 23062 16259 23114 16311
rect 23182 16259 23234 16311
rect 23302 16259 23354 16311
rect 22094 15198 22146 15250
rect 22214 15198 22266 15250
rect 22334 15198 22386 15250
rect 22454 15198 22506 15250
rect 22574 15198 22626 15250
rect 22094 15078 22146 15130
rect 22214 15078 22266 15130
rect 22334 15078 22386 15130
rect 22454 15078 22506 15130
rect 22574 15078 22626 15130
rect 22063 14580 22115 14632
rect 22183 14580 22235 14632
rect 22303 14580 22355 14632
rect 22423 14580 22475 14632
rect 22543 14580 22595 14632
rect 22063 14460 22115 14512
rect 22183 14460 22235 14512
rect 22303 14460 22355 14512
rect 22423 14460 22475 14512
rect 22543 14460 22595 14512
rect 17931 14008 18191 14268
rect 10858 13398 10910 13450
rect 10996 13398 11048 13450
rect 10861 13271 10913 13323
rect 11000 13269 11052 13321
rect 10860 13118 10912 13170
rect 11000 13127 11052 13179
rect 11401 12654 11453 12706
rect 11585 12651 11637 12703
rect 11398 12526 11450 12578
rect 11583 12518 11635 12570
rect 11399 12381 11451 12433
rect 11576 12381 11628 12433
rect 12271 12363 12323 12415
rect 12409 12363 12461 12415
rect 12274 12236 12326 12288
rect 12413 12234 12465 12286
rect 12273 12083 12325 12135
rect 12413 12092 12465 12144
rect 8609 11609 8661 11661
rect 8731 11610 8783 11662
rect 8876 11613 8928 11665
rect 8615 11497 8667 11549
rect 8746 11498 8798 11550
rect 8885 11498 8937 11550
rect 11344 9927 11396 9979
rect 11521 9938 11573 9990
rect 11278 9796 11330 9848
rect 11414 9806 11466 9858
rect 11561 9801 11613 9853
rect 11440 7930 11492 7982
rect 11574 7930 11626 7982
rect 11435 7816 11487 7868
rect 11564 7804 11616 7856
rect 5395 7492 5447 7544
rect 5592 7508 5644 7560
rect 5731 7512 5783 7564
rect 5875 7508 5927 7560
rect 5358 7362 5410 7414
rect 5507 7367 5559 7419
rect 5680 7374 5732 7426
rect 5854 7388 5906 7440
rect 5327 7242 5379 7294
rect 5478 7250 5530 7302
rect 5641 7254 5693 7306
rect 5802 7254 5854 7306
rect 5943 7259 5995 7311
rect 12966 7253 13018 7305
rect 13102 7253 13154 7305
rect 12961 7140 13013 7192
rect 13097 7133 13149 7185
rect 8598 7016 8650 7068
rect 8741 7016 8793 7068
rect 8953 7021 9005 7073
rect 8598 6904 8650 6956
rect 8746 6904 8798 6956
rect 8984 6904 9036 6956
rect 12502 5340 12554 5392
rect 12679 5351 12731 5403
rect 12436 5209 12488 5261
rect 12572 5219 12624 5271
rect 12719 5214 12771 5266
rect 4828 -1042 4880 -990
rect 4992 -1044 5044 -992
rect 4828 -1169 4880 -1117
rect 4994 -1156 5046 -1104
rect 4828 -1307 4880 -1255
rect 4999 -1296 5051 -1244
rect 4894 -1621 4946 -1569
rect 5060 -1608 5112 -1556
rect 4894 -1759 4946 -1707
rect 5065 -1748 5117 -1696
rect 4796 -2305 4848 -2253
rect 4547 -2408 4599 -2356
rect 4687 -2408 4739 -2356
rect 4549 -2529 4601 -2477
rect 4695 -2532 4747 -2480
rect 4815 -2537 4867 -2485
rect 5051 -2717 5103 -2665
rect 5217 -2704 5269 -2652
rect 5051 -2855 5103 -2803
rect 5222 -2844 5274 -2792
rect 4955 -3135 5007 -3083
rect 5121 -3122 5173 -3070
rect 4955 -3273 5007 -3221
rect 5126 -3262 5178 -3210
rect 4932 -3549 4984 -3497
rect 5098 -3536 5150 -3484
rect 4932 -3687 4984 -3635
rect 5103 -3676 5155 -3624
rect 4978 -4028 5030 -3976
rect 5144 -4015 5196 -3963
rect 4978 -4166 5030 -4114
rect 5149 -4155 5201 -4103
rect 5083 -4571 5135 -4519
rect 5249 -4558 5301 -4506
rect 5083 -4709 5135 -4657
rect 5254 -4698 5306 -4646
rect 17919 13787 18179 13943
rect 19222 13750 19378 14114
rect 20393 13831 20653 14091
rect 22116 13928 22272 14084
rect 22498 13928 22654 14084
rect 22917 13928 23073 14084
rect 37935 14106 37987 14158
rect 38055 14106 38107 14158
rect 38175 14106 38227 14158
rect 38295 14106 38347 14158
rect 38415 14106 38467 14158
rect 37935 13986 37987 14038
rect 38055 13986 38107 14038
rect 38175 13986 38227 14038
rect 38295 13986 38347 14038
rect 38415 13986 38467 14038
rect 22006 13564 22058 13616
rect 22429 13564 22481 13616
rect 22720 13564 22772 13616
rect 21838 13187 21890 13239
rect 22077 13187 22129 13239
rect 22410 13187 22462 13239
rect 29830 13273 29882 13325
rect 29950 13273 30002 13325
rect 30070 13273 30122 13325
rect 30190 13273 30242 13325
rect 30310 13273 30362 13325
rect 29830 13153 29882 13205
rect 29950 13153 30002 13205
rect 30070 13153 30122 13205
rect 30190 13153 30242 13205
rect 30310 13153 30362 13205
rect 19670 11136 19722 11188
rect 19911 11141 19963 11193
rect 20150 11143 20202 11195
rect 20377 11143 20429 11195
rect 22481 11115 22533 11167
rect 22476 10971 22528 11023
rect 64929 13720 64981 13772
rect 65188 13716 65240 13768
rect 65429 13651 65481 13703
rect 64933 13569 64985 13621
rect 65200 13539 65252 13591
rect 65424 13498 65476 13550
rect 64932 13400 64984 13452
rect 65190 13402 65242 13454
rect 65422 13355 65474 13407
rect 64982 13225 65034 13277
rect 65184 13220 65236 13272
rect 65347 13208 65399 13260
rect 41755 12582 41807 12634
rect 41755 12332 41807 12384
rect 41755 12108 41807 12160
rect 37877 10732 37929 10784
rect 37997 10732 38049 10784
rect 38117 10732 38169 10784
rect 38237 10732 38289 10784
rect 38357 10732 38409 10784
rect 37877 10612 37929 10664
rect 37997 10612 38049 10664
rect 38117 10612 38169 10664
rect 38237 10612 38289 10664
rect 38357 10612 38409 10664
rect 28784 9841 28836 9893
rect 29025 9846 29077 9898
rect 29264 9848 29316 9900
rect 29491 9848 29543 9900
rect 19628 9090 19680 9142
rect 19869 9095 19921 9147
rect 20108 9097 20160 9149
rect 20335 9097 20387 9149
rect 22939 7822 22991 7874
rect 23180 7827 23232 7879
rect 23419 7829 23471 7881
rect 23646 7829 23698 7881
rect 28728 6847 28780 6899
rect 28969 6852 29021 6904
rect 29208 6854 29260 6906
rect 29435 6854 29487 6906
rect 22134 6737 22186 6789
rect 22430 6737 22482 6789
rect 18072 6618 18124 6670
rect 18192 6618 18244 6670
rect 18312 6618 18364 6670
rect 18432 6618 18484 6670
rect 18552 6618 18604 6670
rect 18672 6618 18724 6670
rect 18792 6618 18844 6670
rect 18912 6618 18964 6670
rect 19032 6618 19084 6670
rect 19152 6618 19204 6670
rect 19272 6618 19324 6670
rect 19392 6618 19444 6670
rect 32075 9827 32127 9879
rect 47793 8176 47845 8228
rect 47949 8176 48001 8228
rect 54014 9262 54066 9314
rect 54133 9262 54185 9314
rect 54252 9263 54304 9315
rect 54374 9264 54426 9316
rect 54492 9263 54544 9315
rect 54014 9144 54066 9196
rect 54133 9144 54185 9196
rect 54254 9145 54306 9197
rect 54374 9147 54426 9199
rect 54493 9143 54545 9195
rect 61584 9269 61636 9321
rect 61703 9269 61755 9321
rect 61822 9270 61874 9322
rect 61944 9271 61996 9323
rect 62062 9270 62114 9322
rect 61584 9151 61636 9203
rect 61703 9151 61755 9203
rect 61824 9152 61876 9204
rect 61944 9154 61996 9206
rect 62063 9150 62115 9202
rect 43285 6948 43441 7104
rect 43828 6948 43984 7104
rect 44538 6948 44694 7104
rect 46195 7021 46247 7073
rect 46441 7016 46493 7068
rect 46721 7018 46773 7070
rect 46937 7026 46989 7078
rect 39342 6452 39498 6608
rect 43825 6022 43877 6074
rect 44074 6009 44126 6061
rect 44308 6004 44360 6056
rect 44530 6008 44582 6060
rect 27149 4353 27201 4405
rect 27381 4353 27433 4405
rect 30470 4435 30522 4487
rect 27146 4157 27198 4209
rect 27381 4157 27433 4209
rect 30470 4174 30522 4226
rect 53788 4608 53840 4660
rect 53907 4608 53959 4660
rect 54026 4609 54078 4661
rect 54148 4610 54200 4662
rect 54266 4609 54318 4661
rect 53788 4490 53840 4542
rect 53907 4490 53959 4542
rect 54028 4491 54080 4543
rect 54148 4493 54200 4545
rect 54267 4489 54319 4541
rect 98889 4667 98941 4719
rect 99064 4661 99116 4713
rect 98887 4508 98939 4560
rect 99065 4512 99117 4564
rect 98890 4343 98942 4395
rect 99078 4338 99130 4390
rect 91420 4201 91472 4253
rect 91539 4201 91591 4253
rect 91658 4202 91710 4254
rect 91780 4203 91832 4255
rect 91898 4202 91950 4254
rect 91420 4083 91472 4135
rect 91539 4083 91591 4135
rect 91660 4084 91712 4136
rect 91780 4086 91832 4138
rect 91899 4082 91951 4134
rect 95236 2614 95288 2666
rect 95356 2614 95408 2666
rect 95476 2614 95528 2666
rect 95236 2494 95288 2546
rect 95356 2494 95408 2546
rect 95476 2494 95528 2546
rect 95236 2374 95288 2426
rect 95356 2374 95408 2426
rect 95476 2374 95528 2426
rect 90007 -366 90059 -314
rect 90131 -354 90183 -302
rect 90025 -483 90077 -431
rect 90149 -495 90201 -443
rect 18145 -1598 18197 -1546
rect 18452 -1593 18504 -1541
rect 18702 -1586 18754 -1534
rect 58357 -3092 58409 -3040
rect 58527 -3067 58579 -3015
rect 58356 -3266 58408 -3214
rect 58522 -3265 58574 -3213
rect 68218 -3693 68270 -3641
rect 68392 -3694 68444 -3642
rect 68219 -3859 68271 -3807
rect 68417 -3864 68469 -3812
rect 98602 -814 98654 -762
rect 98777 -820 98829 -768
rect 98600 -973 98652 -921
rect 98778 -969 98830 -917
rect 98603 -1138 98655 -1086
rect 98791 -1143 98843 -1091
rect 98635 -2018 98687 -1966
rect 98809 -2019 98861 -1967
rect 98636 -2184 98688 -2132
rect 98834 -2189 98886 -2137
rect 98605 -2915 98657 -2863
rect 98779 -2916 98831 -2864
rect 98606 -3081 98658 -3029
rect 98804 -3086 98856 -3034
rect 98597 -3398 98649 -3346
rect 98771 -3399 98823 -3347
rect 98598 -3564 98650 -3512
rect 98796 -3569 98848 -3517
rect 98635 -3950 98687 -3898
rect 98809 -3951 98861 -3899
rect 98636 -4116 98688 -4064
rect 98834 -4121 98886 -4069
rect 87136 -4776 87188 -4724
rect 87256 -4776 87308 -4724
rect 87376 -4776 87428 -4724
rect 87136 -4896 87188 -4844
rect 87256 -4896 87308 -4844
rect 87376 -4896 87428 -4844
rect 87136 -5016 87188 -4964
rect 87256 -5016 87308 -4964
rect 87376 -5016 87428 -4964
rect 48446 -9393 48498 -9341
rect 48585 -9405 48637 -9353
rect 48440 -9509 48492 -9457
rect 48588 -9530 48640 -9478
rect 48443 -9623 48495 -9571
rect 48588 -9646 48640 -9594
rect 52348 -11446 52400 -11394
rect 52553 -11433 52605 -11381
rect 52808 -11431 52860 -11379
rect 53077 -11423 53129 -11371
rect 53319 -11420 53371 -11368
rect 52350 -11636 52402 -11584
rect 52556 -11628 52608 -11576
rect 52789 -11618 52841 -11566
rect 53034 -11615 53086 -11563
rect 53247 -11603 53299 -11551
rect 53406 -11602 53458 -11550
rect 52341 -11812 52393 -11760
rect 52509 -11811 52561 -11759
rect 52707 -11809 52759 -11757
rect 52918 -11806 52970 -11754
rect 53157 -11796 53209 -11744
rect 53355 -11788 53407 -11736
rect 49199 -14208 49251 -14156
rect 49319 -14208 49371 -14156
rect 49439 -14208 49491 -14156
rect 49199 -14328 49251 -14276
rect 49319 -14328 49371 -14276
rect 49439 -14328 49491 -14276
rect 98606 -7526 98658 -7474
rect 98726 -7526 98778 -7474
rect 98846 -7526 98898 -7474
rect 98606 -7646 98658 -7594
rect 98726 -7646 98778 -7594
rect 98846 -7646 98898 -7594
rect 98606 -7766 98658 -7714
rect 98726 -7766 98778 -7714
rect 98846 -7766 98898 -7714
<< metal2 >>
rect -3079 62800 -2804 62816
rect -3079 62744 -3052 62800
rect -2996 62798 -2804 62800
rect -2996 62744 -2888 62798
rect -3079 62742 -2888 62744
rect -2832 62742 -2804 62798
rect -3079 62686 -2804 62742
rect -3079 62673 -2886 62686
rect -3079 62617 -3052 62673
rect -2996 62630 -2886 62673
rect -2830 62630 -2804 62686
rect -2996 62617 -2804 62630
rect -3079 62546 -2804 62617
rect -3079 62535 -2881 62546
rect -3079 62479 -3052 62535
rect -2996 62490 -2881 62535
rect -2825 62490 -2804 62546
rect -2996 62479 -2804 62490
rect -3079 62466 -2804 62479
rect -4059 61372 -3689 61414
rect -4059 61359 -3845 61372
rect -4059 61303 -4011 61359
rect -3955 61316 -3845 61359
rect -3789 61316 -3689 61372
rect -3955 61303 -3689 61316
rect -4059 61232 -3689 61303
rect -4059 61221 -3840 61232
rect -4059 61165 -4011 61221
rect -3955 61176 -3840 61221
rect -3784 61176 -3689 61232
rect -3955 61165 -3689 61176
rect -4059 61136 -3689 61165
rect -2698 52728 -2423 52744
rect -2698 52672 -2671 52728
rect -2615 52726 -2423 52728
rect -2615 52672 -2507 52726
rect -2698 52670 -2507 52672
rect -2451 52670 -2423 52726
rect -2698 52614 -2423 52670
rect -2698 52601 -2505 52614
rect -2698 52545 -2671 52601
rect -2615 52558 -2505 52601
rect -2449 52558 -2423 52614
rect -2615 52545 -2423 52558
rect -2698 52474 -2423 52545
rect -2698 52463 -2500 52474
rect -2698 52407 -2671 52463
rect -2615 52418 -2500 52463
rect -2444 52418 -2423 52474
rect -2615 52407 -2423 52418
rect -2698 52394 -2423 52407
rect -3907 52216 -3537 52258
rect -3907 52203 -3693 52216
rect -3907 52147 -3859 52203
rect -3803 52160 -3693 52203
rect -3637 52160 -3537 52216
rect -3803 52147 -3537 52160
rect -3907 52076 -3537 52147
rect -3907 52065 -3688 52076
rect -3907 52009 -3859 52065
rect -3803 52020 -3688 52065
rect -3632 52020 -3537 52076
rect -3803 52009 -3537 52020
rect -3907 51980 -3537 52009
rect -2388 44202 -2113 44218
rect -2388 44146 -2361 44202
rect -2305 44200 -2113 44202
rect -2305 44146 -2197 44200
rect -2388 44144 -2197 44146
rect -2141 44144 -2113 44200
rect -2388 44088 -2113 44144
rect -2388 44075 -2195 44088
rect -2388 44019 -2361 44075
rect -2305 44032 -2195 44075
rect -2139 44032 -2113 44088
rect -2305 44019 -2113 44032
rect -2388 43948 -2113 44019
rect -2388 43937 -2190 43948
rect -2388 43881 -2361 43937
rect -2305 43892 -2190 43937
rect -2134 43892 -2113 43948
rect -2305 43881 -2113 43892
rect -2388 43868 -2113 43881
rect -2381 43661 -2106 43677
rect -2381 43605 -2354 43661
rect -2298 43659 -2106 43661
rect -2298 43605 -2190 43659
rect -2381 43603 -2190 43605
rect -2134 43603 -2106 43659
rect -2381 43547 -2106 43603
rect -2381 43534 -2188 43547
rect -2381 43478 -2354 43534
rect -2298 43491 -2188 43534
rect -2132 43491 -2106 43547
rect -2298 43478 -2106 43491
rect -2381 43407 -2106 43478
rect -2381 43396 -2183 43407
rect -2381 43340 -2354 43396
rect -2298 43351 -2183 43396
rect -2127 43351 -2106 43407
rect -2298 43340 -2106 43351
rect -2381 43327 -2106 43340
rect -2489 36768 -2214 36784
rect -2489 36712 -2462 36768
rect -2406 36766 -2214 36768
rect -2406 36712 -2298 36766
rect -2489 36710 -2298 36712
rect -2242 36710 -2214 36766
rect -2489 36654 -2214 36710
rect -2489 36641 -2296 36654
rect -2489 36585 -2462 36641
rect -2406 36598 -2296 36641
rect -2240 36598 -2214 36654
rect -2406 36585 -2214 36598
rect -2489 36514 -2214 36585
rect -2489 36503 -2291 36514
rect -2489 36447 -2462 36503
rect -2406 36458 -2291 36503
rect -2235 36458 -2214 36514
rect -2406 36447 -2214 36458
rect -2489 36434 -2214 36447
rect 2010 28027 2740 28118
rect 2010 28019 2607 28027
rect 2010 27963 2041 28019
rect 2097 28016 2417 28019
rect 2097 27963 2220 28016
rect 2010 27960 2220 27963
rect 2276 27963 2417 28016
rect 2473 27971 2607 28019
rect 2663 27971 2740 28027
rect 2473 27963 2740 27971
rect 2276 27960 2740 27963
rect 2010 27892 2740 27960
rect 2010 27836 2044 27892
rect 2100 27884 2607 27892
rect 2100 27881 2409 27884
rect 2100 27836 2220 27881
rect 2010 27825 2220 27836
rect 2276 27828 2409 27881
rect 2465 27836 2607 27884
rect 2663 27836 2740 27892
rect 2465 27828 2740 27836
rect 2276 27825 2740 27828
rect 2010 27720 2740 27825
rect -3588 25044 -3261 25051
rect -3592 25043 -3165 25044
rect -3592 25040 -1026 25043
rect -3592 24988 -3571 25040
rect -3519 24988 -3451 25040
rect -3399 24988 -3331 25040
rect -3279 24988 -1026 25040
rect -3592 24951 -1026 24988
rect -3592 24920 -464 24951
rect -3592 24868 -3571 24920
rect -3519 24868 -3451 24920
rect -3399 24868 -3331 24920
rect -3279 24868 -464 24920
rect -3592 24840 -464 24868
rect -3592 24800 -1026 24840
rect -3592 24748 -3571 24800
rect -3519 24748 -3451 24800
rect -3399 24748 -3331 24800
rect -3279 24748 -1026 24800
rect -3592 24732 -3165 24748
rect -1775 20749 -1405 23311
rect 8582 21777 9071 21859
rect 8582 21757 8980 21777
rect 8582 21701 8765 21757
rect 8821 21721 8980 21757
rect 9036 21721 9071 21777
rect 8821 21701 9071 21721
rect 8582 21604 9071 21701
rect 8582 21594 8916 21604
rect 8582 21538 8654 21594
rect 8710 21548 8916 21594
rect 8972 21548 9071 21604
rect 8710 21538 9071 21548
rect 8582 21353 9071 21538
rect 8582 21343 8892 21353
rect 8582 21287 8672 21343
rect 8728 21297 8892 21343
rect 8948 21297 9071 21353
rect 8728 21287 9071 21297
rect 8582 21236 9071 21287
rect -265 20749 1066 20974
rect -1794 20711 1066 20749
rect -1794 20691 377 20711
rect -1794 20635 162 20691
rect 218 20655 377 20691
rect 433 20655 1066 20711
rect 218 20635 1066 20655
rect -1794 20538 1066 20635
rect -1794 20528 313 20538
rect -1794 20472 51 20528
rect 107 20482 313 20528
rect 369 20482 1066 20538
rect 107 20472 1066 20482
rect -1794 20340 1066 20472
rect -265 20287 1066 20340
rect -265 20277 289 20287
rect -265 20221 69 20277
rect 125 20231 289 20277
rect 345 20231 1066 20287
rect 125 20221 1066 20231
rect -265 19888 1066 20221
rect 2458 16522 2515 16888
rect -198 15447 -142 15448
rect -298 15391 -132 15447
rect -198 15252 -142 15391
rect 2503 15111 2561 15299
rect 1122 14386 1678 14442
rect 2080 14352 2136 14528
rect 919 13812 975 14048
rect 1943 11782 1999 12188
rect 8582 11731 8987 21236
rect 41677 20265 44259 20474
rect 9800 17596 10310 17660
rect 9800 17544 9836 17596
rect 9888 17544 9964 17596
rect 10016 17593 10310 17596
rect 10016 17544 10115 17593
rect 9800 17541 10115 17544
rect 10167 17541 10310 17593
rect 9800 17470 10310 17541
rect 9800 17437 21600 17470
rect 9800 17385 9834 17437
rect 9886 17435 10181 17437
rect 9886 17385 10005 17435
rect 9800 17383 10005 17385
rect 10057 17385 10181 17435
rect 10233 17385 21600 17437
rect 10057 17383 21600 17385
rect 9800 17274 21600 17383
rect 9800 17258 10197 17274
rect 9800 17253 10048 17258
rect 9800 17201 9846 17253
rect 9898 17206 10048 17253
rect 10100 17222 10197 17258
rect 10249 17250 21600 17274
rect 10249 17222 10310 17250
rect 10100 17206 10310 17222
rect 9898 17201 10310 17206
rect 9800 17160 10310 17201
rect 9750 16933 10260 16990
rect 9750 16926 10054 16933
rect 9750 16923 9923 16926
rect 9750 16871 9795 16923
rect 9847 16874 9923 16923
rect 9975 16881 10054 16926
rect 10106 16914 10260 16933
rect 10106 16881 20684 16914
rect 9975 16874 20684 16881
rect 9847 16871 20684 16874
rect 9750 16749 20684 16871
rect 9750 16744 10107 16749
rect 9750 16726 9959 16744
rect 9750 16674 9790 16726
rect 9842 16692 9959 16726
rect 10011 16697 10107 16744
rect 10159 16697 20684 16749
rect 10011 16692 20684 16697
rect 9842 16674 20684 16692
rect 9750 16646 20684 16674
rect 9750 16616 10260 16646
rect 9750 16606 10141 16616
rect 9750 16575 9964 16606
rect 9750 16523 9767 16575
rect 9819 16554 9964 16575
rect 10016 16564 10141 16606
rect 10193 16564 10260 16616
rect 10016 16554 10260 16564
rect 9819 16523 10260 16554
rect 9750 16490 10260 16523
rect 12240 16138 19962 16431
rect 12240 14461 12533 16138
rect 19669 15309 19962 16138
rect 20416 15743 20684 16646
rect 21380 16095 21600 17250
rect 22731 16826 23374 16880
rect 22731 16774 22815 16826
rect 22867 16774 22935 16826
rect 22987 16774 23055 16826
rect 23107 16774 23175 16826
rect 23227 16774 23295 16826
rect 23347 16799 23374 16826
rect 23347 16774 37528 16799
rect 22731 16706 37528 16774
rect 22731 16654 22815 16706
rect 22867 16654 22935 16706
rect 22987 16654 23055 16706
rect 23107 16654 23175 16706
rect 23227 16654 23295 16706
rect 23347 16654 37528 16706
rect 22731 16594 37528 16654
rect 22731 16591 23374 16594
rect 22735 16494 23393 16495
rect 22735 16431 36567 16494
rect 22735 16379 22822 16431
rect 22874 16379 22942 16431
rect 22994 16379 23062 16431
rect 23114 16379 23182 16431
rect 23234 16379 23302 16431
rect 23354 16379 36567 16431
rect 22735 16311 36567 16379
rect 22735 16259 22822 16311
rect 22874 16259 22942 16311
rect 22994 16259 23062 16311
rect 23114 16259 23182 16311
rect 23234 16259 23302 16311
rect 23354 16289 36567 16311
rect 23354 16259 23393 16289
rect 22735 16213 23393 16259
rect 22738 16210 23393 16213
rect 21380 16087 24210 16095
rect 21380 15884 35629 16087
rect 21380 15875 24210 15884
rect 20416 15712 24234 15743
rect 20416 15506 33629 15712
rect 20416 15475 24234 15506
rect 19669 15286 23314 15309
rect 19669 15250 31910 15286
rect 19669 15198 22094 15250
rect 22146 15198 22214 15250
rect 22266 15198 22334 15250
rect 22386 15198 22454 15250
rect 22506 15198 22574 15250
rect 22626 15198 31910 15250
rect 19669 15130 31910 15198
rect 10823 14168 12533 14461
rect 12941 14846 19271 15094
rect 19669 15078 22094 15130
rect 22146 15078 22214 15130
rect 22266 15078 22334 15130
rect 22386 15078 22454 15130
rect 22506 15078 22574 15130
rect 22626 15078 31910 15130
rect 19669 15039 31910 15078
rect 19669 15016 23314 15039
rect 10823 13450 11116 14168
rect 10823 13398 10858 13450
rect 10910 13398 10996 13450
rect 11048 13398 11116 13450
rect 10823 13323 11116 13398
rect 10823 13271 10861 13323
rect 10913 13321 11116 13323
rect 10913 13271 11000 13321
rect 10823 13269 11000 13271
rect 11052 13269 11116 13321
rect 10823 13179 11116 13269
rect 10823 13170 11000 13179
rect 10823 13118 10860 13170
rect 10912 13127 11000 13170
rect 11052 13127 11116 13179
rect 10912 13118 11116 13127
rect 10823 13099 11116 13118
rect 11365 12708 11683 12801
rect 11365 12652 11399 12708
rect 11455 12705 11683 12708
rect 11455 12652 11583 12705
rect 11365 12649 11583 12652
rect 11639 12649 11683 12705
rect 11365 12580 11683 12649
rect 11365 12524 11396 12580
rect 11452 12572 11683 12580
rect 11452 12524 11581 12572
rect 11365 12516 11581 12524
rect 11637 12516 11683 12572
rect 11365 12435 11683 12516
rect 11365 12379 11397 12435
rect 11453 12379 11574 12435
rect 11630 12379 11683 12435
rect 11365 12334 11683 12379
rect 12236 12459 12529 12469
rect 12236 12415 12533 12459
rect 12236 12363 12271 12415
rect 12323 12363 12409 12415
rect 12461 12363 12533 12415
rect 12236 12288 12533 12363
rect 12236 12236 12274 12288
rect 12326 12286 12533 12288
rect 12326 12236 12413 12286
rect 12236 12234 12413 12236
rect 12465 12234 12533 12286
rect 12236 12144 12533 12234
rect 12236 12135 12413 12144
rect 12236 12083 12273 12135
rect 12325 12092 12413 12135
rect 12465 12092 12533 12144
rect 12325 12083 12533 12092
rect 12236 12064 12533 12083
rect 8578 11667 8995 11731
rect 8578 11664 8873 11667
rect 8578 11663 8727 11664
rect 8578 11607 8607 11663
rect 8663 11608 8727 11663
rect 8783 11611 8873 11664
rect 8929 11611 8995 11667
rect 8783 11608 8995 11611
rect 8663 11607 8995 11608
rect 8578 11552 8995 11607
rect 8578 11496 8612 11552
rect 8668 11496 8743 11552
rect 8799 11496 8883 11552
rect 8939 11496 8995 11552
rect 8578 11488 8995 11496
rect 11239 10062 11632 10070
rect 12240 10062 12533 12064
rect 11238 10056 12533 10062
rect 11236 9990 12533 10056
rect 11236 9979 11521 9990
rect 11236 9927 11344 9979
rect 11396 9938 11521 9979
rect 11573 9938 12533 9990
rect 11396 9927 12533 9938
rect 11236 9858 12533 9927
rect 11236 9848 11414 9858
rect 11236 9796 11278 9848
rect 11330 9806 11414 9848
rect 11466 9853 12533 9858
rect 11466 9806 11561 9853
rect 11330 9801 11561 9806
rect 11613 9801 12533 9853
rect 11330 9796 12533 9801
rect 11236 9772 12533 9796
rect 11238 9769 12533 9772
rect 12941 8826 13189 14846
rect 19023 14678 19271 14846
rect 22059 14694 22659 14696
rect 22045 14678 22661 14694
rect 19023 14632 30057 14678
rect 19023 14580 22063 14632
rect 22115 14580 22183 14632
rect 22235 14580 22303 14632
rect 22355 14580 22423 14632
rect 22475 14580 22543 14632
rect 22595 14580 30057 14632
rect 19023 14512 30057 14580
rect 19023 14460 22063 14512
rect 22115 14460 22183 14512
rect 22235 14460 22303 14512
rect 22355 14460 22423 14512
rect 22475 14460 22543 14512
rect 22595 14460 30057 14512
rect 19023 14430 30057 14460
rect 22045 14427 22661 14430
rect 17357 14268 18262 14318
rect 17357 14180 17931 14268
rect 17357 14160 17795 14180
rect 17357 14104 17580 14160
rect 17636 14124 17795 14160
rect 17851 14124 17931 14180
rect 17636 14104 17931 14124
rect 17357 14008 17931 14104
rect 18191 14008 18262 14268
rect 17357 14007 18262 14008
rect 17357 13997 17731 14007
rect 17357 13941 17469 13997
rect 17525 13951 17731 13997
rect 17787 13951 18262 14007
rect 17525 13945 18262 13951
rect 17525 13943 17920 13945
rect 17976 13943 18262 13945
rect 17525 13941 17919 13943
rect 17357 13787 17919 13941
rect 18179 13787 18262 13943
rect 17357 13756 18262 13787
rect 17357 13746 17707 13756
rect 17357 13690 17487 13746
rect 17543 13700 17707 13746
rect 17763 13700 18262 13756
rect 19198 14114 19410 14168
rect 19198 13750 19222 14114
rect 19378 13750 19410 14114
rect 20130 14145 20656 14238
rect 20130 14104 20725 14145
rect 20130 14094 20480 14104
rect 20130 14038 20260 14094
rect 20316 14091 20480 14094
rect 20536 14091 20725 14104
rect 20316 14038 20393 14091
rect 20130 13905 20393 14038
rect 20130 13849 20251 13905
rect 20307 13849 20393 13905
rect 20130 13831 20393 13849
rect 20653 13831 20725 14091
rect 22087 14087 23144 14135
rect 22087 14084 28904 14087
rect 22087 13928 22116 14084
rect 22272 13928 22498 14084
rect 22654 13928 22917 14084
rect 23073 13928 28904 14084
rect 22087 13926 28904 13928
rect 22087 13904 23144 13926
rect 20130 13787 20725 13831
rect 19198 13738 19410 13750
rect 17543 13695 18262 13700
rect 17543 13690 17924 13695
rect 17357 13639 17924 13690
rect 17980 13639 18262 13695
rect 17357 13551 18262 13639
rect 11423 8578 13189 8826
rect 13467 13461 13922 13516
rect 17357 13495 17705 13551
rect 17761 13495 18262 13551
rect 17357 13461 18262 13495
rect 13467 13285 18262 13461
rect 13467 13116 18226 13285
rect 11423 7982 11671 8578
rect 11423 7930 11440 7982
rect 11492 7930 11574 7982
rect 11626 7930 11671 7982
rect 11423 7868 11671 7930
rect 11423 7816 11435 7868
rect 11487 7856 11671 7868
rect 11487 7816 11564 7856
rect 11423 7804 11564 7816
rect 11616 7804 11671 7856
rect 11423 7781 11671 7804
rect 5268 7566 6063 7709
rect 5268 7562 5729 7566
rect 5268 7546 5590 7562
rect 5268 7490 5393 7546
rect 5449 7506 5590 7546
rect 5646 7510 5729 7562
rect 5785 7562 6063 7566
rect 5785 7510 5873 7562
rect 5646 7506 5873 7510
rect 5929 7506 6063 7562
rect 5449 7490 6063 7506
rect 5268 7442 6063 7490
rect 5268 7428 5852 7442
rect 5268 7421 5678 7428
rect 5268 7416 5505 7421
rect 5268 7360 5356 7416
rect 5412 7365 5505 7416
rect 5561 7372 5678 7421
rect 5734 7386 5852 7428
rect 5908 7386 6063 7442
rect 5734 7372 6063 7386
rect 5561 7365 6063 7372
rect 5412 7360 6063 7365
rect 5268 7313 6063 7360
rect 5268 7308 5941 7313
rect 5268 7304 5639 7308
rect 5268 7296 5476 7304
rect 5268 7240 5325 7296
rect 5381 7248 5476 7296
rect 5532 7252 5639 7304
rect 5695 7252 5800 7308
rect 5856 7257 5941 7308
rect 5997 7257 6063 7313
rect 5856 7252 6063 7257
rect 5532 7248 6063 7252
rect 5381 7240 6063 7248
rect 5268 7226 6063 7240
rect 12940 7305 13192 7311
rect 12940 7253 12966 7305
rect 13018 7253 13102 7305
rect 13154 7253 13192 7305
rect 12940 7192 13192 7253
rect 12940 7140 12961 7192
rect 13013 7185 13192 7192
rect 13013 7140 13097 7185
rect 8560 7075 9108 7137
rect 12940 7133 13097 7140
rect 13149 7133 13192 7185
rect 12940 7111 13192 7133
rect 8560 7068 8951 7075
rect 8560 7012 8590 7068
rect 8650 7016 8731 7068
rect 8793 7019 8951 7068
rect 9007 7019 9108 7075
rect 8793 7016 9108 7019
rect 8646 7012 8731 7016
rect 8787 7012 9108 7016
rect 8560 6958 9108 7012
rect 8560 6902 8596 6958
rect 8652 6956 9108 6958
rect 8652 6953 8746 6956
rect 8798 6953 8984 6956
rect 8652 6902 8737 6953
rect 8798 6904 8977 6953
rect 9036 6904 9108 6956
rect 8560 6897 8737 6902
rect 8793 6897 8977 6904
rect 9033 6897 9108 6904
rect 8560 6879 9108 6897
rect 12397 5486 12483 5488
rect 12397 5469 12848 5486
rect 12382 5466 12848 5469
rect 12941 5466 13189 7111
rect 12382 5403 13189 5466
rect 12382 5392 12679 5403
rect 12382 5340 12502 5392
rect 12554 5351 12679 5392
rect 12731 5351 13189 5403
rect 12554 5340 13189 5351
rect 12382 5271 13189 5340
rect 12382 5261 12572 5271
rect 12382 5209 12436 5261
rect 12488 5219 12572 5261
rect 12624 5266 13189 5271
rect 12624 5219 12719 5266
rect 12488 5214 12719 5219
rect 12771 5218 13189 5266
rect 12771 5214 12848 5218
rect 12488 5209 12848 5214
rect 12382 5176 12848 5209
rect 4778 -988 5148 -932
rect 4778 -1044 4826 -988
rect 4882 -990 5148 -988
rect 4882 -1044 4990 -990
rect 4778 -1046 4990 -1044
rect 5046 -1046 5148 -990
rect 4778 -1102 5148 -1046
rect 4778 -1115 4992 -1102
rect 4778 -1171 4826 -1115
rect 4882 -1158 4992 -1115
rect 5048 -1158 5148 -1102
rect 4882 -1171 5148 -1158
rect 4778 -1242 5148 -1171
rect 4778 -1253 4997 -1242
rect 4778 -1309 4826 -1253
rect 4882 -1298 4997 -1253
rect 5053 -1298 5148 -1242
rect 4882 -1309 5148 -1298
rect 4778 -1338 5148 -1309
rect 4844 -1554 5214 -1512
rect 4844 -1567 5058 -1554
rect 4844 -1623 4892 -1567
rect 4948 -1610 5058 -1567
rect 5114 -1610 5214 -1554
rect 4948 -1623 5214 -1610
rect 4844 -1694 5214 -1623
rect 4844 -1705 5063 -1694
rect 4844 -1761 4892 -1705
rect 4948 -1750 5063 -1705
rect 5119 -1750 5214 -1694
rect 4948 -1761 5214 -1750
rect 4844 -1790 5214 -1761
rect 4506 -2253 4874 -2240
rect 4506 -2305 4796 -2253
rect 4848 -2255 4874 -2253
rect 4848 -2305 11467 -2255
rect 4506 -2356 11467 -2305
rect 4506 -2408 4547 -2356
rect 4599 -2408 4687 -2356
rect 4739 -2408 11467 -2356
rect 4506 -2455 11467 -2408
rect 4506 -2477 4874 -2455
rect 4506 -2529 4549 -2477
rect 4601 -2480 4874 -2477
rect 4601 -2529 4695 -2480
rect 4506 -2532 4695 -2529
rect 4747 -2485 4874 -2480
rect 4747 -2532 4815 -2485
rect 4506 -2537 4815 -2532
rect 4867 -2537 4874 -2485
rect 4506 -2563 4874 -2537
rect 5001 -2650 5371 -2608
rect 5001 -2663 5215 -2650
rect 5001 -2719 5049 -2663
rect 5105 -2706 5215 -2663
rect 5271 -2706 5371 -2650
rect 5105 -2719 5371 -2706
rect 5001 -2790 5371 -2719
rect 5001 -2801 5220 -2790
rect 5001 -2857 5049 -2801
rect 5105 -2846 5220 -2801
rect 5276 -2846 5371 -2790
rect 5105 -2857 5371 -2846
rect 5001 -2886 5371 -2857
rect 4905 -3068 5275 -3026
rect 4905 -3081 5119 -3068
rect 4905 -3137 4953 -3081
rect 5009 -3124 5119 -3081
rect 5175 -3124 5275 -3068
rect 5009 -3137 5275 -3124
rect 4905 -3208 5275 -3137
rect 4905 -3219 5124 -3208
rect 4905 -3275 4953 -3219
rect 5009 -3264 5124 -3219
rect 5180 -3264 5275 -3208
rect 5009 -3275 5275 -3264
rect 4905 -3304 5275 -3275
rect 4882 -3482 5252 -3440
rect 4882 -3495 5096 -3482
rect 4882 -3551 4930 -3495
rect 4986 -3538 5096 -3495
rect 5152 -3538 5252 -3482
rect 4986 -3551 5252 -3538
rect 4882 -3622 5252 -3551
rect 4882 -3633 5101 -3622
rect 4882 -3689 4930 -3633
rect 4986 -3678 5101 -3633
rect 5157 -3678 5252 -3622
rect 4986 -3689 5252 -3678
rect 4882 -3718 5252 -3689
rect 11285 -3874 11467 -2455
rect 13467 -3380 13922 13116
rect 17908 12969 18198 13116
rect 19228 12977 19380 13738
rect 20406 12980 20725 13787
rect 21938 13658 22849 13700
rect 25430 13658 26138 13671
rect 21938 13618 26138 13658
rect 21938 13616 25520 13618
rect 21938 13564 22006 13616
rect 22058 13564 22429 13616
rect 22481 13564 22720 13616
rect 22772 13564 25520 13616
rect 21938 13562 25520 13564
rect 25576 13562 25708 13618
rect 25764 13562 25903 13618
rect 25959 13562 26138 13618
rect 21938 13522 26138 13562
rect 21938 13497 22849 13522
rect 25430 13504 26138 13522
rect 25430 13503 26015 13504
rect 21799 13290 22548 13292
rect 21799 13239 25263 13290
rect 21799 13187 21838 13239
rect 21890 13187 22077 13239
rect 22129 13187 22410 13239
rect 22462 13187 25263 13239
rect 21799 13142 25263 13187
rect 22003 13130 25263 13142
rect 17908 12820 18711 12969
rect 19228 12825 19543 12977
rect 19391 12008 19543 12825
rect 20406 12807 22149 12980
rect 21976 12098 22149 12807
rect 25103 12633 25263 13130
rect 25103 12473 28368 12633
rect 21863 11925 22149 12098
rect 27026 11727 27558 11886
rect 28208 11854 28368 12473
rect 28743 12234 28904 13926
rect 29809 13377 30057 14430
rect 29808 13325 30422 13377
rect 29808 13273 29830 13325
rect 29882 13273 29950 13325
rect 30002 13273 30070 13325
rect 30122 13273 30190 13325
rect 30242 13273 30310 13325
rect 30362 13273 30422 13325
rect 29808 13205 30422 13273
rect 29808 13153 29830 13205
rect 29882 13153 29950 13205
rect 30002 13153 30070 13205
rect 30122 13153 30190 13205
rect 30242 13153 30310 13205
rect 30362 13153 30422 13205
rect 29808 13140 30422 13153
rect 28743 12073 30776 12234
rect 30615 11894 30776 12073
rect 27026 11650 27185 11727
rect 28208 11694 30139 11854
rect 30615 11733 30983 11894
rect 26304 11491 27236 11650
rect 19654 11190 19738 11204
rect 19654 11134 19668 11190
rect 19724 11134 19738 11190
rect 19654 11121 19738 11134
rect 19895 11195 19979 11209
rect 19895 11139 19909 11195
rect 19965 11139 19979 11195
rect 19895 11126 19979 11139
rect 20120 11197 20230 11220
rect 20120 11141 20148 11197
rect 20204 11141 20230 11197
rect 20120 11110 20230 11141
rect 20361 11197 20445 11211
rect 20361 11141 20375 11197
rect 20431 11141 20445 11197
rect 20361 11128 20445 11141
rect 22449 11208 22560 11220
rect 22449 11167 22574 11208
rect 21983 11113 22080 11125
rect 22449 11115 22481 11167
rect 22533 11115 22574 11167
rect 22449 11113 22574 11115
rect 21983 11072 22574 11113
rect 21983 11023 22575 11072
rect 21983 10971 22476 11023
rect 22528 10971 22575 11023
rect 21983 10919 22575 10971
rect 21984 10918 22575 10919
rect 27077 11032 27236 11491
rect 27077 10873 27324 11032
rect 29660 10913 29767 11694
rect 30822 10849 30983 11733
rect 31663 9951 31910 15039
rect 33423 12307 33629 15506
rect 33149 12101 33629 12307
rect 33423 11895 33629 12101
rect 28768 9895 28852 9909
rect 28768 9839 28782 9895
rect 28838 9839 28852 9895
rect 28768 9826 28852 9839
rect 29009 9900 29093 9914
rect 29009 9844 29023 9900
rect 29079 9844 29093 9900
rect 29009 9831 29093 9844
rect 29248 9902 29332 9916
rect 29248 9846 29262 9902
rect 29318 9846 29332 9902
rect 29248 9833 29332 9846
rect 29475 9902 29559 9916
rect 29475 9846 29489 9902
rect 29545 9846 29559 9902
rect 29475 9833 29559 9846
rect 30909 9879 32327 9951
rect 35426 9902 35629 15884
rect 36362 11499 36567 16289
rect 37323 12528 37528 16594
rect 41677 15783 41886 20265
rect 37851 14158 38494 14212
rect 37851 14106 37935 14158
rect 37987 14106 38055 14158
rect 38107 14106 38175 14158
rect 38227 14106 38295 14158
rect 38347 14106 38415 14158
rect 38467 14106 38494 14158
rect 37851 14038 38494 14106
rect 37851 13986 37935 14038
rect 37987 13986 38055 14038
rect 38107 13986 38175 14038
rect 38227 13986 38295 14038
rect 38347 13986 38415 14038
rect 38467 13986 38494 14038
rect 37851 13923 38494 13986
rect 37852 10840 37971 13923
rect 38108 10840 38227 13923
rect 38374 10840 38493 13923
rect 41677 12634 41885 15783
rect 64769 13772 65603 13916
rect 64769 13720 64929 13772
rect 64981 13768 65603 13772
rect 64981 13720 65188 13768
rect 64769 13716 65188 13720
rect 65240 13759 65603 13768
rect 65240 13716 71106 13759
rect 64769 13703 71106 13716
rect 64769 13651 65429 13703
rect 65481 13651 71106 13703
rect 64769 13621 71106 13651
rect 64769 13569 64933 13621
rect 64985 13591 71106 13621
rect 64985 13569 65200 13591
rect 64769 13539 65200 13569
rect 65252 13550 71106 13591
rect 65252 13539 65424 13550
rect 64769 13498 65424 13539
rect 65476 13498 71106 13550
rect 64769 13454 71106 13498
rect 64769 13452 65190 13454
rect 64769 13400 64932 13452
rect 64984 13402 65190 13452
rect 65242 13407 71106 13454
rect 65242 13402 65422 13407
rect 64984 13400 65422 13402
rect 64769 13355 65422 13400
rect 65474 13355 71106 13407
rect 64769 13318 71106 13355
rect 64769 13277 65603 13318
rect 64769 13225 64982 13277
rect 65034 13272 65603 13277
rect 65034 13225 65184 13272
rect 64769 13220 65184 13225
rect 65236 13260 65603 13272
rect 65236 13220 65347 13260
rect 64769 13208 65347 13220
rect 65399 13208 65603 13260
rect 64769 13020 65603 13208
rect 39735 12603 41562 12604
rect 39735 12349 41564 12603
rect 37793 10784 38571 10840
rect 37793 10732 37877 10784
rect 37929 10732 37997 10784
rect 38049 10732 38117 10784
rect 38169 10732 38237 10784
rect 38289 10732 38357 10784
rect 38409 10732 38571 10784
rect 37793 10664 38571 10732
rect 37793 10612 37877 10664
rect 37929 10612 37997 10664
rect 38049 10612 38117 10664
rect 38169 10612 38237 10664
rect 38289 10612 38357 10664
rect 38409 10612 38571 10664
rect 37793 10547 38571 10612
rect 38124 10314 38319 10344
rect 30909 9827 32075 9879
rect 32127 9827 32327 9879
rect 30909 9794 32327 9827
rect 34743 9821 35629 9902
rect 31663 9749 31910 9794
rect 32011 9792 32327 9794
rect 32170 9693 32327 9792
rect 35426 9791 35629 9821
rect 38116 9812 38319 10314
rect 35450 9784 35605 9791
rect 35021 9697 35271 9715
rect 34756 9668 35271 9697
rect 34756 9620 35439 9668
rect 34858 9581 35439 9620
rect 38116 9581 38311 9812
rect 34858 9492 38311 9581
rect 29769 9190 31596 9392
rect 35150 9389 38311 9492
rect 35367 9386 38311 9389
rect 41307 9609 41564 12349
rect 41677 12582 41755 12634
rect 41807 12582 41885 12634
rect 41677 12384 41885 12582
rect 41677 12332 41755 12384
rect 41807 12332 41885 12384
rect 41677 12214 41885 12332
rect 41677 12160 42058 12214
rect 41677 12108 41755 12160
rect 41807 12108 42058 12160
rect 41677 12061 42058 12108
rect 19612 9144 19696 9158
rect 19612 9088 19626 9144
rect 19682 9088 19696 9144
rect 19612 9075 19696 9088
rect 19853 9149 19937 9163
rect 19853 9093 19867 9149
rect 19923 9093 19937 9149
rect 19853 9080 19937 9093
rect 20060 9151 20200 9180
rect 20060 9095 20106 9151
rect 20162 9095 20200 9151
rect 20060 9070 20200 9095
rect 20319 9151 20403 9165
rect 20319 9095 20333 9151
rect 20389 9095 20403 9151
rect 20319 9082 20403 9095
rect 26250 8881 27154 9033
rect 29769 8898 29971 9190
rect 30473 9032 30883 9048
rect 30473 9019 30667 9032
rect 30473 8963 30535 9019
rect 30591 8976 30667 9019
rect 30723 9031 30883 9032
rect 30723 8976 30792 9031
rect 30591 8975 30792 8976
rect 30848 8975 30883 9031
rect 30591 8963 30883 8975
rect 30473 8922 30883 8963
rect 30473 8906 30665 8922
rect 21824 8205 22125 8362
rect 19342 7505 19505 8018
rect 21968 7600 22125 8205
rect 27002 8017 27154 8881
rect 29614 8696 30098 8898
rect 30473 8850 30532 8906
rect 30588 8866 30665 8906
rect 30721 8866 30792 8922
rect 30848 8866 30883 8922
rect 30588 8850 30883 8866
rect 30473 8795 30883 8850
rect 30473 8793 30654 8795
rect 30473 8737 30529 8793
rect 30585 8739 30654 8793
rect 30710 8739 30792 8795
rect 30848 8739 30883 8795
rect 30585 8737 30883 8739
rect 30473 8717 30883 8737
rect 22923 7876 23007 7890
rect 22923 7820 22937 7876
rect 22993 7820 23007 7876
rect 22923 7807 23007 7820
rect 23164 7881 23248 7895
rect 23164 7825 23178 7881
rect 23234 7825 23248 7881
rect 23164 7812 23248 7825
rect 23403 7883 23487 7897
rect 23403 7827 23417 7883
rect 23473 7827 23487 7883
rect 23403 7814 23487 7827
rect 23630 7883 23714 7897
rect 23630 7827 23644 7883
rect 23700 7827 23714 7883
rect 27002 7865 27262 8017
rect 23630 7814 23714 7827
rect 19076 7342 19505 7505
rect 21969 7489 22125 7600
rect 21177 7488 22125 7489
rect 19076 6748 19239 7342
rect 20972 7320 22125 7488
rect 17938 6711 19507 6748
rect 17938 6670 19508 6711
rect 17938 6618 18072 6670
rect 18124 6618 18192 6670
rect 18244 6618 18312 6670
rect 18364 6618 18432 6670
rect 18484 6618 18552 6670
rect 18604 6618 18672 6670
rect 18724 6618 18792 6670
rect 18844 6618 18912 6670
rect 18964 6618 19032 6670
rect 19084 6618 19152 6670
rect 19204 6618 19272 6670
rect 19324 6618 19392 6670
rect 19444 6618 19508 6670
rect 17938 6585 19508 6618
rect 20972 6253 21508 7320
rect 22095 6791 26596 6907
rect 28712 6901 28796 6915
rect 28712 6845 28726 6901
rect 28782 6845 28796 6901
rect 28712 6832 28796 6845
rect 28953 6906 29037 6920
rect 28953 6850 28967 6906
rect 29023 6850 29037 6906
rect 28953 6837 29037 6850
rect 29192 6908 29276 6922
rect 29192 6852 29206 6908
rect 29262 6852 29276 6908
rect 29192 6839 29276 6852
rect 29419 6908 29503 6922
rect 29419 6852 29433 6908
rect 29489 6852 29503 6908
rect 29419 6839 29503 6852
rect 22083 6789 26596 6791
rect 22083 6737 22134 6789
rect 22186 6737 22430 6789
rect 22482 6737 26596 6789
rect 22083 6707 26596 6737
rect 22085 6705 26596 6707
rect 22085 6683 22546 6705
rect 20972 5718 22844 6253
rect 18271 -774 18995 -726
rect 18271 -830 18331 -774
rect 18387 -830 18995 -774
rect 18271 -916 18995 -830
rect 18271 -935 18795 -916
rect 18271 -991 18536 -935
rect 18592 -972 18795 -935
rect 18851 -972 18995 -916
rect 18592 -991 18995 -972
rect 18271 -1063 18995 -991
rect 18080 -1531 18860 -1470
rect 18080 -1534 18706 -1531
rect 18080 -1541 18702 -1534
rect 18080 -1544 18452 -1541
rect 18504 -1544 18702 -1541
rect 18080 -1600 18143 -1544
rect 18199 -1600 18452 -1544
rect 18508 -1586 18702 -1544
rect 18508 -1587 18706 -1586
rect 18762 -1587 18860 -1531
rect 18508 -1600 18860 -1587
rect 18080 -1660 18860 -1600
rect 22309 -2588 22844 5718
rect 26394 5828 26596 6705
rect 31394 5828 31596 9190
rect 38043 7647 38298 9386
rect 41307 9354 48122 9609
rect 47867 8256 48122 9354
rect 53921 9318 54794 9377
rect 53921 9317 54372 9318
rect 53921 9314 54248 9317
rect 53921 9258 54012 9314
rect 54068 9258 54131 9314
rect 54187 9261 54248 9314
rect 54304 9262 54372 9317
rect 54428 9317 54794 9318
rect 54428 9262 54489 9317
rect 54304 9261 54489 9262
rect 54545 9261 54794 9317
rect 54187 9258 54794 9261
rect 53921 9204 54794 9258
rect 53921 9200 54373 9204
rect 53921 9198 54253 9200
rect 53921 9142 54012 9198
rect 54068 9142 54130 9198
rect 54186 9144 54253 9198
rect 54309 9148 54373 9200
rect 54429 9197 54794 9204
rect 54429 9148 54491 9197
rect 54309 9147 54374 9148
rect 54426 9147 54491 9148
rect 54309 9144 54491 9147
rect 54186 9142 54491 9144
rect 53921 9141 54491 9142
rect 54547 9141 54794 9197
rect 53921 9088 54794 9141
rect 61491 9325 62361 9385
rect 61491 9324 61942 9325
rect 61491 9321 61818 9324
rect 61491 9265 61582 9321
rect 61638 9265 61701 9321
rect 61757 9268 61818 9321
rect 61874 9269 61942 9324
rect 61998 9324 62361 9325
rect 61998 9269 62059 9324
rect 61874 9268 62059 9269
rect 62115 9268 62361 9324
rect 61757 9265 62361 9268
rect 61491 9211 62361 9265
rect 61491 9207 61943 9211
rect 61491 9205 61823 9207
rect 61491 9149 61582 9205
rect 61638 9149 61700 9205
rect 61756 9151 61823 9205
rect 61879 9155 61943 9207
rect 61999 9204 62361 9211
rect 61999 9155 62061 9204
rect 61879 9154 61944 9155
rect 61996 9154 62061 9155
rect 61879 9151 62061 9154
rect 61756 9149 62061 9151
rect 61491 9148 62061 9149
rect 62117 9148 62361 9204
rect 61491 9099 62361 9148
rect 47615 8252 48122 8256
rect 47615 8228 48258 8252
rect 47615 8176 47793 8228
rect 47845 8176 47949 8228
rect 48001 8176 48258 8228
rect 47615 8150 48258 8176
rect 47690 8137 48258 8150
rect 47690 7940 48260 8137
rect 47852 7647 48122 7648
rect 38043 7392 48122 7647
rect 44110 7124 44460 7130
rect 43227 7106 44715 7124
rect 43227 6946 43283 7106
rect 43443 6946 43826 7106
rect 43986 6946 44536 7106
rect 44696 6946 44715 7106
rect 46136 7080 47059 7119
rect 46136 7075 46935 7080
rect 46136 7019 46193 7075
rect 46249 7072 46935 7075
rect 46249 7070 46719 7072
rect 46249 7019 46439 7070
rect 46136 7014 46439 7019
rect 46495 7016 46719 7070
rect 46775 7024 46935 7072
rect 46991 7024 47059 7080
rect 47852 7063 48122 7392
rect 46775 7016 47059 7024
rect 46495 7014 47059 7016
rect 46136 6961 47059 7014
rect 43227 6919 44715 6946
rect 44110 6850 44480 6919
rect 44110 6810 44460 6850
rect 38263 6610 39669 6671
rect 38263 6450 38310 6610
rect 38470 6608 39669 6610
rect 38470 6452 39342 6608
rect 39498 6452 39669 6608
rect 38470 6450 39669 6452
rect 38263 6430 39669 6450
rect 38287 6418 39669 6430
rect 38287 6414 38493 6418
rect 43759 6076 44718 6127
rect 43759 6020 43823 6076
rect 43879 6063 44718 6076
rect 43879 6020 44072 6063
rect 44128 6062 44718 6063
rect 43759 6007 44072 6020
rect 44128 6058 44528 6062
rect 44128 6007 44306 6058
rect 43759 6002 44306 6007
rect 44362 6006 44528 6058
rect 44584 6006 44718 6062
rect 44362 6002 44718 6006
rect 43759 5971 44718 6002
rect 26394 5626 31596 5828
rect 30400 4489 30604 4659
rect 47853 4548 48122 7063
rect 27094 4407 27485 4463
rect 27094 4351 27147 4407
rect 27203 4351 27379 4407
rect 27435 4351 27485 4407
rect 27094 4211 27485 4351
rect 27094 4155 27144 4211
rect 27200 4155 27379 4211
rect 27435 4155 27485 4211
rect 27094 4108 27485 4155
rect 30400 4433 30468 4489
rect 30524 4433 30604 4489
rect 30400 4228 30604 4433
rect 45792 4279 48122 4548
rect 53695 4664 54568 4724
rect 53695 4663 54146 4664
rect 53695 4660 54022 4663
rect 53695 4604 53786 4660
rect 53842 4604 53905 4660
rect 53961 4607 54022 4660
rect 54078 4608 54146 4663
rect 54202 4663 54568 4664
rect 54202 4608 54263 4663
rect 54078 4607 54263 4608
rect 54319 4607 54568 4663
rect 53961 4604 54568 4607
rect 53695 4550 54568 4604
rect 53695 4546 54147 4550
rect 53695 4544 54027 4546
rect 53695 4488 53786 4544
rect 53842 4488 53904 4544
rect 53960 4490 54027 4544
rect 54083 4494 54147 4546
rect 54203 4543 54568 4550
rect 54203 4494 54265 4543
rect 54083 4493 54148 4494
rect 54200 4493 54265 4494
rect 54083 4490 54265 4493
rect 53960 4488 54265 4490
rect 53695 4487 54265 4488
rect 54321 4487 54568 4543
rect 53695 4412 54568 4487
rect 98848 4723 99160 4739
rect 98848 4667 98889 4723
rect 98945 4717 99160 4723
rect 98945 4667 99064 4717
rect 98848 4661 99064 4667
rect 99120 4661 99160 4717
rect 98848 4568 99160 4661
rect 98848 4564 99065 4568
rect 98848 4508 98887 4564
rect 98943 4512 99065 4564
rect 99121 4512 99160 4568
rect 98943 4508 99160 4512
rect 53695 4319 54344 4412
rect 53701 4315 54344 4319
rect 98848 4399 99160 4508
rect 98848 4343 98890 4399
rect 98946 4394 99160 4399
rect 98946 4343 99078 4394
rect 98848 4338 99078 4343
rect 99134 4338 99160 4394
rect 53701 4314 54194 4315
rect 30400 4172 30468 4228
rect 30524 4172 30604 4228
rect 30400 4129 30604 4172
rect 91327 4257 92059 4316
rect 98848 4305 99160 4338
rect 91327 4256 91778 4257
rect 91327 4253 91654 4256
rect 91327 4197 91418 4253
rect 91474 4197 91537 4253
rect 91593 4200 91654 4253
rect 91710 4201 91778 4256
rect 91834 4256 92059 4257
rect 91834 4201 91895 4256
rect 91710 4200 91895 4201
rect 91951 4200 92059 4256
rect 91593 4197 92059 4200
rect 91327 4143 92059 4197
rect 91327 4139 91779 4143
rect 91327 4137 91659 4139
rect 91327 4081 91418 4137
rect 91474 4081 91536 4137
rect 91592 4083 91659 4137
rect 91715 4087 91779 4139
rect 91835 4136 92059 4143
rect 91835 4087 91897 4136
rect 91715 4086 91780 4087
rect 91832 4086 91897 4087
rect 91715 4083 91897 4086
rect 91592 4081 91897 4083
rect 91327 4080 91897 4081
rect 91953 4080 92059 4136
rect 91327 4051 92059 4080
rect 95080 2785 95620 2970
rect 95080 2666 96818 2785
rect 95080 2614 95236 2666
rect 95288 2614 95356 2666
rect 95408 2614 95476 2666
rect 95528 2614 96818 2666
rect 95080 2546 96818 2614
rect 95080 2494 95236 2546
rect 95288 2494 95356 2546
rect 95408 2494 95476 2546
rect 95528 2494 96818 2546
rect 95080 2426 96818 2494
rect 95080 2374 95236 2426
rect 95288 2374 95356 2426
rect 95408 2374 95476 2426
rect 95528 2390 96818 2426
rect 95528 2374 95620 2390
rect 95080 2270 95620 2374
rect 94369 368 94922 651
rect 89933 -302 90316 -240
rect 89933 -314 90131 -302
rect 89933 -317 90007 -314
rect 86599 -366 90007 -317
rect 90059 -354 90131 -314
rect 90183 -354 90316 -302
rect 90059 -366 90316 -354
rect 86599 -431 90316 -366
rect 86599 -483 90025 -431
rect 90077 -443 90316 -431
rect 90077 -483 90149 -443
rect 86599 -495 90149 -483
rect 90201 -495 90316 -443
rect 86599 -523 90316 -495
rect 89933 -570 90316 -523
rect 22309 -3123 47333 -2588
rect 58344 -3011 58612 -2964
rect 58344 -3036 58524 -3011
rect 58344 -3092 58354 -3036
rect 58410 -3067 58524 -3036
rect 58580 -3067 58612 -3011
rect 58410 -3092 58612 -3067
rect 13467 -3705 17126 -3380
rect 17805 -3874 17987 -3316
rect 4928 -3961 5298 -3919
rect 4928 -3974 5142 -3961
rect 4928 -4030 4976 -3974
rect 5032 -4017 5142 -3974
rect 5198 -4017 5298 -3961
rect 5032 -4030 5298 -4017
rect 4928 -4101 5298 -4030
rect 11285 -4056 17987 -3874
rect 11296 -4081 17960 -4056
rect 4928 -4112 5147 -4101
rect 4928 -4168 4976 -4112
rect 5032 -4157 5147 -4112
rect 5203 -4157 5298 -4101
rect 5032 -4168 5298 -4157
rect 4928 -4197 5298 -4168
rect 5033 -4504 5403 -4462
rect 5033 -4517 5247 -4504
rect 5033 -4573 5081 -4517
rect 5137 -4560 5247 -4517
rect 5303 -4560 5403 -4504
rect 5137 -4573 5403 -4560
rect 5033 -4644 5403 -4573
rect 5033 -4655 5252 -4644
rect 5033 -4711 5081 -4655
rect 5137 -4700 5252 -4655
rect 5308 -4700 5403 -4644
rect 5137 -4711 5403 -4700
rect 5033 -4740 5403 -4711
rect 46962 -5017 47332 -3123
rect 58344 -3209 58612 -3092
rect 58344 -3210 58519 -3209
rect 58344 -3266 58353 -3210
rect 58409 -3265 58519 -3210
rect 58575 -3265 58612 -3209
rect 58409 -3266 58612 -3265
rect 58344 -3325 58612 -3266
rect 68159 -3637 68520 -3628
rect 68159 -3693 68218 -3637
rect 68274 -3638 68520 -3637
rect 68274 -3693 68392 -3638
rect 68159 -3694 68392 -3693
rect 68448 -3694 68520 -3638
rect 68159 -3803 68520 -3694
rect 68159 -3859 68219 -3803
rect 68275 -3808 68520 -3803
rect 68275 -3859 68417 -3808
rect 68159 -3864 68417 -3859
rect 68473 -3864 68520 -3808
rect 68159 -3896 68520 -3864
rect 87090 -4722 87760 -4550
rect 87090 -4778 87132 -4722
rect 87188 -4778 87252 -4722
rect 87308 -4778 87372 -4722
rect 87428 -4778 87760 -4722
rect 87090 -4842 87760 -4778
rect 87090 -4898 87132 -4842
rect 87188 -4898 87252 -4842
rect 87308 -4898 87372 -4842
rect 87428 -4898 87760 -4842
rect 87090 -4962 87760 -4898
rect 45298 -5387 48300 -5017
rect 87090 -5018 87134 -4962
rect 87190 -5018 87252 -4962
rect 87308 -5018 87372 -4962
rect 87428 -5018 87760 -4962
rect 87090 -5090 87760 -5018
rect 47930 -9293 48300 -5387
rect 94639 -7468 94922 368
rect 96448 -5325 96818 2390
rect 98561 -758 98873 -742
rect 98561 -814 98602 -758
rect 98658 -764 98873 -758
rect 98658 -814 98777 -764
rect 98561 -820 98777 -814
rect 98833 -820 98873 -764
rect 98561 -913 98873 -820
rect 98561 -917 98778 -913
rect 98561 -973 98600 -917
rect 98656 -969 98778 -917
rect 98834 -969 98873 -913
rect 98656 -973 98873 -969
rect 98561 -1082 98873 -973
rect 98561 -1138 98603 -1082
rect 98659 -1087 98873 -1082
rect 98659 -1138 98791 -1087
rect 98561 -1143 98791 -1138
rect 98847 -1143 98873 -1087
rect 98561 -1181 98873 -1143
rect 98576 -1962 98937 -1953
rect 98576 -2018 98635 -1962
rect 98691 -1963 98937 -1962
rect 98691 -2018 98809 -1963
rect 98576 -2019 98809 -2018
rect 98865 -2019 98937 -1963
rect 98576 -2128 98937 -2019
rect 98576 -2184 98636 -2128
rect 98692 -2133 98937 -2128
rect 98692 -2184 98834 -2133
rect 98576 -2189 98834 -2184
rect 98890 -2189 98937 -2133
rect 98576 -2221 98937 -2189
rect 98546 -2859 98907 -2850
rect 98546 -2915 98605 -2859
rect 98661 -2860 98907 -2859
rect 98661 -2915 98779 -2860
rect 98546 -2916 98779 -2915
rect 98835 -2916 98907 -2860
rect 98546 -3025 98907 -2916
rect 98546 -3081 98606 -3025
rect 98662 -3030 98907 -3025
rect 98662 -3081 98804 -3030
rect 98546 -3086 98804 -3081
rect 98860 -3086 98907 -3030
rect 98546 -3118 98907 -3086
rect 98538 -3342 98899 -3333
rect 98538 -3398 98597 -3342
rect 98653 -3343 98899 -3342
rect 98653 -3398 98771 -3343
rect 98538 -3399 98771 -3398
rect 98827 -3399 98899 -3343
rect 98538 -3508 98899 -3399
rect 98538 -3564 98598 -3508
rect 98654 -3513 98899 -3508
rect 98654 -3564 98796 -3513
rect 98538 -3569 98796 -3564
rect 98852 -3569 98899 -3513
rect 98538 -3601 98899 -3569
rect 98576 -3894 98937 -3885
rect 98576 -3950 98635 -3894
rect 98691 -3895 98937 -3894
rect 98691 -3950 98809 -3895
rect 98576 -3951 98809 -3950
rect 98865 -3951 98937 -3895
rect 98576 -4060 98937 -3951
rect 98576 -4116 98636 -4060
rect 98692 -4065 98937 -4060
rect 98692 -4116 98834 -4065
rect 98576 -4121 98834 -4116
rect 98890 -4121 98937 -4065
rect 98576 -4153 98937 -4121
rect 98574 -7468 98910 -7460
rect 94639 -7474 98910 -7468
rect 94639 -7526 98606 -7474
rect 98658 -7526 98726 -7474
rect 98778 -7526 98846 -7474
rect 98898 -7526 98910 -7474
rect 94639 -7594 98910 -7526
rect 94639 -7646 98606 -7594
rect 98658 -7646 98726 -7594
rect 98778 -7646 98846 -7594
rect 98898 -7646 98910 -7594
rect 94639 -7714 98910 -7646
rect 94639 -7751 98606 -7714
rect 98574 -7766 98606 -7751
rect 98658 -7766 98726 -7714
rect 98778 -7766 98846 -7714
rect 98898 -7766 98910 -7714
rect 98574 -7800 98910 -7766
rect 47930 -9341 48775 -9293
rect 47930 -9393 48446 -9341
rect 48498 -9353 48775 -9341
rect 48498 -9393 48585 -9353
rect 47930 -9405 48585 -9393
rect 48637 -9405 48775 -9353
rect 47930 -9457 48775 -9405
rect 47930 -9509 48440 -9457
rect 48492 -9478 48775 -9457
rect 48492 -9509 48588 -9478
rect 47930 -9530 48588 -9509
rect 48640 -9530 48775 -9478
rect 47930 -9571 48775 -9530
rect 47930 -9623 48443 -9571
rect 48495 -9594 48775 -9571
rect 48495 -9623 48588 -9594
rect 47930 -9646 48588 -9623
rect 48640 -9646 48775 -9594
rect 47930 -9663 48775 -9646
rect 52279 -11322 53565 -11166
rect 52279 -11366 53571 -11322
rect 52279 -11369 53317 -11366
rect 52279 -11377 53075 -11369
rect 52279 -11379 52806 -11377
rect 52279 -11392 52551 -11379
rect 52279 -11448 52346 -11392
rect 52402 -11435 52551 -11392
rect 52607 -11433 52806 -11379
rect 52862 -11425 53075 -11377
rect 53131 -11422 53317 -11369
rect 53373 -11422 53571 -11366
rect 53131 -11425 53571 -11422
rect 52862 -11433 53571 -11425
rect 52607 -11435 53571 -11433
rect 52402 -11448 53571 -11435
rect 52279 -11548 53571 -11448
rect 52279 -11549 53404 -11548
rect 52279 -11561 53245 -11549
rect 52279 -11564 53032 -11561
rect 52279 -11574 52787 -11564
rect 52279 -11582 52554 -11574
rect 52279 -11638 52348 -11582
rect 52404 -11630 52554 -11582
rect 52610 -11620 52787 -11574
rect 52843 -11617 53032 -11564
rect 53088 -11605 53245 -11561
rect 53301 -11604 53404 -11549
rect 53460 -11604 53571 -11548
rect 53301 -11605 53571 -11604
rect 53088 -11617 53571 -11605
rect 52843 -11620 53571 -11617
rect 52610 -11630 53571 -11620
rect 52404 -11638 53571 -11630
rect 52279 -11734 53571 -11638
rect 52279 -11742 53353 -11734
rect 52279 -11752 53155 -11742
rect 52279 -11755 52916 -11752
rect 52279 -11757 52705 -11755
rect 52279 -11758 52507 -11757
rect 52279 -11814 52339 -11758
rect 52395 -11813 52507 -11758
rect 52563 -11811 52705 -11757
rect 52761 -11808 52916 -11755
rect 52972 -11798 53155 -11752
rect 53211 -11790 53353 -11742
rect 53409 -11790 53571 -11734
rect 53211 -11798 53571 -11790
rect 52972 -11808 53571 -11798
rect 52761 -11811 53571 -11808
rect 52563 -11813 53571 -11811
rect 52395 -11814 53571 -11813
rect 52279 -11848 53571 -11814
rect 48991 -14156 49554 -14074
rect 48991 -14208 49199 -14156
rect 49251 -14208 49319 -14156
rect 49371 -14208 49439 -14156
rect 49491 -14208 49554 -14156
rect 48991 -14276 49554 -14208
rect 48991 -14328 49199 -14276
rect 49251 -14328 49319 -14276
rect 49371 -14328 49439 -14276
rect 49491 -14328 49554 -14276
rect 48991 -14450 49554 -14328
<< via2 >>
rect -3052 62798 -2996 62800
rect -3052 62746 -3050 62798
rect -3050 62746 -2998 62798
rect -2998 62746 -2996 62798
rect -3052 62744 -2996 62746
rect -2888 62796 -2832 62798
rect -2888 62744 -2886 62796
rect -2886 62744 -2834 62796
rect -2834 62744 -2832 62796
rect -2888 62742 -2832 62744
rect -2886 62684 -2830 62686
rect -3052 62671 -2996 62673
rect -3052 62619 -3050 62671
rect -3050 62619 -2998 62671
rect -2998 62619 -2996 62671
rect -2886 62632 -2884 62684
rect -2884 62632 -2832 62684
rect -2832 62632 -2830 62684
rect -2886 62630 -2830 62632
rect -3052 62617 -2996 62619
rect -2881 62544 -2825 62546
rect -3052 62533 -2996 62535
rect -3052 62481 -3050 62533
rect -3050 62481 -2998 62533
rect -2998 62481 -2996 62533
rect -2881 62492 -2879 62544
rect -2879 62492 -2827 62544
rect -2827 62492 -2825 62544
rect -2881 62490 -2825 62492
rect -3052 62479 -2996 62481
rect -3845 61370 -3789 61372
rect -4011 61357 -3955 61359
rect -4011 61305 -4009 61357
rect -4009 61305 -3957 61357
rect -3957 61305 -3955 61357
rect -3845 61318 -3843 61370
rect -3843 61318 -3791 61370
rect -3791 61318 -3789 61370
rect -3845 61316 -3789 61318
rect -4011 61303 -3955 61305
rect -3840 61230 -3784 61232
rect -4011 61219 -3955 61221
rect -4011 61167 -4009 61219
rect -4009 61167 -3957 61219
rect -3957 61167 -3955 61219
rect -3840 61178 -3838 61230
rect -3838 61178 -3786 61230
rect -3786 61178 -3784 61230
rect -3840 61176 -3784 61178
rect -4011 61165 -3955 61167
rect -2671 52726 -2615 52728
rect -2671 52674 -2669 52726
rect -2669 52674 -2617 52726
rect -2617 52674 -2615 52726
rect -2671 52672 -2615 52674
rect -2507 52724 -2451 52726
rect -2507 52672 -2505 52724
rect -2505 52672 -2453 52724
rect -2453 52672 -2451 52724
rect -2507 52670 -2451 52672
rect -2505 52612 -2449 52614
rect -2671 52599 -2615 52601
rect -2671 52547 -2669 52599
rect -2669 52547 -2617 52599
rect -2617 52547 -2615 52599
rect -2505 52560 -2503 52612
rect -2503 52560 -2451 52612
rect -2451 52560 -2449 52612
rect -2505 52558 -2449 52560
rect -2671 52545 -2615 52547
rect -2500 52472 -2444 52474
rect -2671 52461 -2615 52463
rect -2671 52409 -2669 52461
rect -2669 52409 -2617 52461
rect -2617 52409 -2615 52461
rect -2500 52420 -2498 52472
rect -2498 52420 -2446 52472
rect -2446 52420 -2444 52472
rect -2500 52418 -2444 52420
rect -2671 52407 -2615 52409
rect -3693 52214 -3637 52216
rect -3859 52201 -3803 52203
rect -3859 52149 -3857 52201
rect -3857 52149 -3805 52201
rect -3805 52149 -3803 52201
rect -3693 52162 -3691 52214
rect -3691 52162 -3639 52214
rect -3639 52162 -3637 52214
rect -3693 52160 -3637 52162
rect -3859 52147 -3803 52149
rect -3688 52074 -3632 52076
rect -3859 52063 -3803 52065
rect -3859 52011 -3857 52063
rect -3857 52011 -3805 52063
rect -3805 52011 -3803 52063
rect -3688 52022 -3686 52074
rect -3686 52022 -3634 52074
rect -3634 52022 -3632 52074
rect -3688 52020 -3632 52022
rect -3859 52009 -3803 52011
rect -2361 44200 -2305 44202
rect -2361 44148 -2359 44200
rect -2359 44148 -2307 44200
rect -2307 44148 -2305 44200
rect -2361 44146 -2305 44148
rect -2197 44198 -2141 44200
rect -2197 44146 -2195 44198
rect -2195 44146 -2143 44198
rect -2143 44146 -2141 44198
rect -2197 44144 -2141 44146
rect -2195 44086 -2139 44088
rect -2361 44073 -2305 44075
rect -2361 44021 -2359 44073
rect -2359 44021 -2307 44073
rect -2307 44021 -2305 44073
rect -2195 44034 -2193 44086
rect -2193 44034 -2141 44086
rect -2141 44034 -2139 44086
rect -2195 44032 -2139 44034
rect -2361 44019 -2305 44021
rect -2190 43946 -2134 43948
rect -2361 43935 -2305 43937
rect -2361 43883 -2359 43935
rect -2359 43883 -2307 43935
rect -2307 43883 -2305 43935
rect -2190 43894 -2188 43946
rect -2188 43894 -2136 43946
rect -2136 43894 -2134 43946
rect -2190 43892 -2134 43894
rect -2361 43881 -2305 43883
rect -2354 43659 -2298 43661
rect -2354 43607 -2352 43659
rect -2352 43607 -2300 43659
rect -2300 43607 -2298 43659
rect -2354 43605 -2298 43607
rect -2190 43657 -2134 43659
rect -2190 43605 -2188 43657
rect -2188 43605 -2136 43657
rect -2136 43605 -2134 43657
rect -2190 43603 -2134 43605
rect -2188 43545 -2132 43547
rect -2354 43532 -2298 43534
rect -2354 43480 -2352 43532
rect -2352 43480 -2300 43532
rect -2300 43480 -2298 43532
rect -2188 43493 -2186 43545
rect -2186 43493 -2134 43545
rect -2134 43493 -2132 43545
rect -2188 43491 -2132 43493
rect -2354 43478 -2298 43480
rect -2183 43405 -2127 43407
rect -2354 43394 -2298 43396
rect -2354 43342 -2352 43394
rect -2352 43342 -2300 43394
rect -2300 43342 -2298 43394
rect -2183 43353 -2181 43405
rect -2181 43353 -2129 43405
rect -2129 43353 -2127 43405
rect -2183 43351 -2127 43353
rect -2354 43340 -2298 43342
rect -2462 36766 -2406 36768
rect -2462 36714 -2460 36766
rect -2460 36714 -2408 36766
rect -2408 36714 -2406 36766
rect -2462 36712 -2406 36714
rect -2298 36764 -2242 36766
rect -2298 36712 -2296 36764
rect -2296 36712 -2244 36764
rect -2244 36712 -2242 36764
rect -2298 36710 -2242 36712
rect -2296 36652 -2240 36654
rect -2462 36639 -2406 36641
rect -2462 36587 -2460 36639
rect -2460 36587 -2408 36639
rect -2408 36587 -2406 36639
rect -2296 36600 -2294 36652
rect -2294 36600 -2242 36652
rect -2242 36600 -2240 36652
rect -2296 36598 -2240 36600
rect -2462 36585 -2406 36587
rect -2291 36512 -2235 36514
rect -2462 36501 -2406 36503
rect -2462 36449 -2460 36501
rect -2460 36449 -2408 36501
rect -2408 36449 -2406 36501
rect -2291 36460 -2289 36512
rect -2289 36460 -2237 36512
rect -2237 36460 -2235 36512
rect -2291 36458 -2235 36460
rect -2462 36447 -2406 36449
rect 2607 28025 2663 28027
rect 2041 28017 2097 28019
rect 2041 27965 2043 28017
rect 2043 27965 2095 28017
rect 2095 27965 2097 28017
rect 2417 28017 2473 28019
rect 2041 27963 2097 27965
rect 2220 28014 2276 28016
rect 2220 27962 2222 28014
rect 2222 27962 2274 28014
rect 2274 27962 2276 28014
rect 2417 27965 2419 28017
rect 2419 27965 2471 28017
rect 2471 27965 2473 28017
rect 2607 27973 2609 28025
rect 2609 27973 2661 28025
rect 2661 27973 2663 28025
rect 2607 27971 2663 27973
rect 2417 27963 2473 27965
rect 2220 27960 2276 27962
rect 2044 27890 2100 27892
rect 2044 27838 2046 27890
rect 2046 27838 2098 27890
rect 2098 27838 2100 27890
rect 2607 27890 2663 27892
rect 2409 27882 2465 27884
rect 2044 27836 2100 27838
rect 2220 27879 2276 27881
rect 2220 27827 2222 27879
rect 2222 27827 2274 27879
rect 2274 27827 2276 27879
rect 2409 27830 2411 27882
rect 2411 27830 2463 27882
rect 2463 27830 2465 27882
rect 2607 27838 2609 27890
rect 2609 27838 2661 27890
rect 2661 27838 2663 27890
rect 2607 27836 2663 27838
rect 2409 27828 2465 27830
rect 2220 27825 2276 27827
rect 8765 21701 8821 21757
rect 8980 21721 9036 21777
rect 8654 21538 8710 21594
rect 8916 21548 8972 21604
rect 8672 21287 8728 21343
rect 8892 21297 8948 21353
rect 162 20635 218 20691
rect 377 20655 433 20711
rect 51 20472 107 20528
rect 313 20482 369 20538
rect 69 20221 125 20277
rect 289 20231 345 20287
rect 11399 12706 11455 12708
rect 11399 12654 11401 12706
rect 11401 12654 11453 12706
rect 11453 12654 11455 12706
rect 11399 12652 11455 12654
rect 11583 12703 11639 12705
rect 11583 12651 11585 12703
rect 11585 12651 11637 12703
rect 11637 12651 11639 12703
rect 11583 12649 11639 12651
rect 11396 12578 11452 12580
rect 11396 12526 11398 12578
rect 11398 12526 11450 12578
rect 11450 12526 11452 12578
rect 11396 12524 11452 12526
rect 11581 12570 11637 12572
rect 11581 12518 11583 12570
rect 11583 12518 11635 12570
rect 11635 12518 11637 12570
rect 11581 12516 11637 12518
rect 11397 12433 11453 12435
rect 11397 12381 11399 12433
rect 11399 12381 11451 12433
rect 11451 12381 11453 12433
rect 11397 12379 11453 12381
rect 11574 12433 11630 12435
rect 11574 12381 11576 12433
rect 11576 12381 11628 12433
rect 11628 12381 11630 12433
rect 11574 12379 11630 12381
rect 8873 11665 8929 11667
rect 8607 11661 8663 11663
rect 8607 11609 8609 11661
rect 8609 11609 8661 11661
rect 8661 11609 8663 11661
rect 8607 11607 8663 11609
rect 8727 11662 8783 11664
rect 8727 11610 8731 11662
rect 8731 11610 8783 11662
rect 8873 11613 8876 11665
rect 8876 11613 8928 11665
rect 8928 11613 8929 11665
rect 8873 11611 8929 11613
rect 8727 11608 8783 11610
rect 8612 11549 8668 11552
rect 8612 11497 8615 11549
rect 8615 11497 8667 11549
rect 8667 11497 8668 11549
rect 8612 11496 8668 11497
rect 8743 11550 8799 11552
rect 8743 11498 8746 11550
rect 8746 11498 8798 11550
rect 8798 11498 8799 11550
rect 8743 11496 8799 11498
rect 8883 11550 8939 11552
rect 8883 11498 8885 11550
rect 8885 11498 8937 11550
rect 8937 11498 8939 11550
rect 8883 11496 8939 11498
rect 17580 14104 17636 14160
rect 17795 14124 17851 14180
rect 18056 14056 18112 14112
rect 17469 13941 17525 13997
rect 17731 13951 17787 14007
rect 17920 13943 17976 13945
rect 17920 13889 17976 13943
rect 17487 13690 17543 13746
rect 17707 13700 17763 13756
rect 20260 14038 20316 14094
rect 20480 14091 20536 14104
rect 20480 14048 20536 14091
rect 20251 13849 20307 13905
rect 20478 13843 20534 13899
rect 17924 13639 17980 13695
rect 17705 13495 17761 13551
rect 5729 7564 5785 7566
rect 5590 7560 5646 7562
rect 5393 7544 5449 7546
rect 5393 7492 5395 7544
rect 5395 7492 5447 7544
rect 5447 7492 5449 7544
rect 5590 7508 5592 7560
rect 5592 7508 5644 7560
rect 5644 7508 5646 7560
rect 5729 7512 5731 7564
rect 5731 7512 5783 7564
rect 5783 7512 5785 7564
rect 5729 7510 5785 7512
rect 5873 7560 5929 7562
rect 5590 7506 5646 7508
rect 5873 7508 5875 7560
rect 5875 7508 5927 7560
rect 5927 7508 5929 7560
rect 5873 7506 5929 7508
rect 5393 7490 5449 7492
rect 5852 7440 5908 7442
rect 5678 7426 5734 7428
rect 5505 7419 5561 7421
rect 5356 7414 5412 7416
rect 5356 7362 5358 7414
rect 5358 7362 5410 7414
rect 5410 7362 5412 7414
rect 5505 7367 5507 7419
rect 5507 7367 5559 7419
rect 5559 7367 5561 7419
rect 5678 7374 5680 7426
rect 5680 7374 5732 7426
rect 5732 7374 5734 7426
rect 5852 7388 5854 7440
rect 5854 7388 5906 7440
rect 5906 7388 5908 7440
rect 5852 7386 5908 7388
rect 5678 7372 5734 7374
rect 5505 7365 5561 7367
rect 5356 7360 5412 7362
rect 5941 7311 5997 7313
rect 5639 7306 5695 7308
rect 5476 7302 5532 7304
rect 5325 7294 5381 7296
rect 5325 7242 5327 7294
rect 5327 7242 5379 7294
rect 5379 7242 5381 7294
rect 5476 7250 5478 7302
rect 5478 7250 5530 7302
rect 5530 7250 5532 7302
rect 5639 7254 5641 7306
rect 5641 7254 5693 7306
rect 5693 7254 5695 7306
rect 5639 7252 5695 7254
rect 5800 7306 5856 7308
rect 5800 7254 5802 7306
rect 5802 7254 5854 7306
rect 5854 7254 5856 7306
rect 5941 7259 5943 7311
rect 5943 7259 5995 7311
rect 5995 7259 5997 7311
rect 5941 7257 5997 7259
rect 5800 7252 5856 7254
rect 5476 7248 5532 7250
rect 5325 7240 5381 7242
rect 8951 7073 9007 7075
rect 8590 7016 8598 7068
rect 8598 7016 8646 7068
rect 8731 7016 8741 7068
rect 8741 7016 8787 7068
rect 8951 7021 8953 7073
rect 8953 7021 9005 7073
rect 9005 7021 9007 7073
rect 8951 7019 9007 7021
rect 8590 7012 8646 7016
rect 8731 7012 8787 7016
rect 8596 6956 8652 6958
rect 8596 6904 8598 6956
rect 8598 6904 8650 6956
rect 8650 6904 8652 6956
rect 8596 6902 8652 6904
rect 8737 6904 8746 6953
rect 8746 6904 8793 6953
rect 8977 6904 8984 6953
rect 8984 6904 9033 6953
rect 8737 6897 8793 6904
rect 8977 6897 9033 6904
rect 4826 -990 4882 -988
rect 4826 -1042 4828 -990
rect 4828 -1042 4880 -990
rect 4880 -1042 4882 -990
rect 4826 -1044 4882 -1042
rect 4990 -992 5046 -990
rect 4990 -1044 4992 -992
rect 4992 -1044 5044 -992
rect 5044 -1044 5046 -992
rect 4990 -1046 5046 -1044
rect 4992 -1104 5048 -1102
rect 4826 -1117 4882 -1115
rect 4826 -1169 4828 -1117
rect 4828 -1169 4880 -1117
rect 4880 -1169 4882 -1117
rect 4992 -1156 4994 -1104
rect 4994 -1156 5046 -1104
rect 5046 -1156 5048 -1104
rect 4992 -1158 5048 -1156
rect 4826 -1171 4882 -1169
rect 4997 -1244 5053 -1242
rect 4826 -1255 4882 -1253
rect 4826 -1307 4828 -1255
rect 4828 -1307 4880 -1255
rect 4880 -1307 4882 -1255
rect 4997 -1296 4999 -1244
rect 4999 -1296 5051 -1244
rect 5051 -1296 5053 -1244
rect 4997 -1298 5053 -1296
rect 4826 -1309 4882 -1307
rect 5058 -1556 5114 -1554
rect 4892 -1569 4948 -1567
rect 4892 -1621 4894 -1569
rect 4894 -1621 4946 -1569
rect 4946 -1621 4948 -1569
rect 5058 -1608 5060 -1556
rect 5060 -1608 5112 -1556
rect 5112 -1608 5114 -1556
rect 5058 -1610 5114 -1608
rect 4892 -1623 4948 -1621
rect 5063 -1696 5119 -1694
rect 4892 -1707 4948 -1705
rect 4892 -1759 4894 -1707
rect 4894 -1759 4946 -1707
rect 4946 -1759 4948 -1707
rect 5063 -1748 5065 -1696
rect 5065 -1748 5117 -1696
rect 5117 -1748 5119 -1696
rect 5063 -1750 5119 -1748
rect 4892 -1761 4948 -1759
rect 5215 -2652 5271 -2650
rect 5049 -2665 5105 -2663
rect 5049 -2717 5051 -2665
rect 5051 -2717 5103 -2665
rect 5103 -2717 5105 -2665
rect 5215 -2704 5217 -2652
rect 5217 -2704 5269 -2652
rect 5269 -2704 5271 -2652
rect 5215 -2706 5271 -2704
rect 5049 -2719 5105 -2717
rect 5220 -2792 5276 -2790
rect 5049 -2803 5105 -2801
rect 5049 -2855 5051 -2803
rect 5051 -2855 5103 -2803
rect 5103 -2855 5105 -2803
rect 5220 -2844 5222 -2792
rect 5222 -2844 5274 -2792
rect 5274 -2844 5276 -2792
rect 5220 -2846 5276 -2844
rect 5049 -2857 5105 -2855
rect 5119 -3070 5175 -3068
rect 4953 -3083 5009 -3081
rect 4953 -3135 4955 -3083
rect 4955 -3135 5007 -3083
rect 5007 -3135 5009 -3083
rect 5119 -3122 5121 -3070
rect 5121 -3122 5173 -3070
rect 5173 -3122 5175 -3070
rect 5119 -3124 5175 -3122
rect 4953 -3137 5009 -3135
rect 5124 -3210 5180 -3208
rect 4953 -3221 5009 -3219
rect 4953 -3273 4955 -3221
rect 4955 -3273 5007 -3221
rect 5007 -3273 5009 -3221
rect 5124 -3262 5126 -3210
rect 5126 -3262 5178 -3210
rect 5178 -3262 5180 -3210
rect 5124 -3264 5180 -3262
rect 4953 -3275 5009 -3273
rect 5096 -3484 5152 -3482
rect 4930 -3497 4986 -3495
rect 4930 -3549 4932 -3497
rect 4932 -3549 4984 -3497
rect 4984 -3549 4986 -3497
rect 5096 -3536 5098 -3484
rect 5098 -3536 5150 -3484
rect 5150 -3536 5152 -3484
rect 5096 -3538 5152 -3536
rect 4930 -3551 4986 -3549
rect 5101 -3624 5157 -3622
rect 4930 -3635 4986 -3633
rect 4930 -3687 4932 -3635
rect 4932 -3687 4984 -3635
rect 4984 -3687 4986 -3635
rect 5101 -3676 5103 -3624
rect 5103 -3676 5155 -3624
rect 5155 -3676 5157 -3624
rect 5101 -3678 5157 -3676
rect 4930 -3689 4986 -3687
rect 25520 13562 25576 13618
rect 25708 13562 25764 13618
rect 25903 13562 25959 13618
rect 19668 11188 19724 11190
rect 19668 11136 19670 11188
rect 19670 11136 19722 11188
rect 19722 11136 19724 11188
rect 19668 11134 19724 11136
rect 19909 11193 19965 11195
rect 19909 11141 19911 11193
rect 19911 11141 19963 11193
rect 19963 11141 19965 11193
rect 19909 11139 19965 11141
rect 20148 11195 20204 11197
rect 20148 11143 20150 11195
rect 20150 11143 20202 11195
rect 20202 11143 20204 11195
rect 20148 11141 20204 11143
rect 20375 11195 20431 11197
rect 20375 11143 20377 11195
rect 20377 11143 20429 11195
rect 20429 11143 20431 11195
rect 20375 11141 20431 11143
rect 28782 9893 28838 9895
rect 28782 9841 28784 9893
rect 28784 9841 28836 9893
rect 28836 9841 28838 9893
rect 28782 9839 28838 9841
rect 29023 9898 29079 9900
rect 29023 9846 29025 9898
rect 29025 9846 29077 9898
rect 29077 9846 29079 9898
rect 29023 9844 29079 9846
rect 29262 9900 29318 9902
rect 29262 9848 29264 9900
rect 29264 9848 29316 9900
rect 29316 9848 29318 9900
rect 29262 9846 29318 9848
rect 29489 9900 29545 9902
rect 29489 9848 29491 9900
rect 29491 9848 29543 9900
rect 29543 9848 29545 9900
rect 29489 9846 29545 9848
rect 19626 9142 19682 9144
rect 19626 9090 19628 9142
rect 19628 9090 19680 9142
rect 19680 9090 19682 9142
rect 19626 9088 19682 9090
rect 19867 9147 19923 9149
rect 19867 9095 19869 9147
rect 19869 9095 19921 9147
rect 19921 9095 19923 9147
rect 19867 9093 19923 9095
rect 20106 9149 20162 9151
rect 20106 9097 20108 9149
rect 20108 9097 20160 9149
rect 20160 9097 20162 9149
rect 20106 9095 20162 9097
rect 20333 9149 20389 9151
rect 20333 9097 20335 9149
rect 20335 9097 20387 9149
rect 20387 9097 20389 9149
rect 20333 9095 20389 9097
rect 30535 8963 30591 9019
rect 30667 8976 30723 9032
rect 30792 8975 30848 9031
rect 30532 8850 30588 8906
rect 30665 8866 30721 8922
rect 30792 8866 30848 8922
rect 30529 8737 30585 8793
rect 30654 8739 30710 8795
rect 30792 8739 30848 8795
rect 22937 7874 22993 7876
rect 22937 7822 22939 7874
rect 22939 7822 22991 7874
rect 22991 7822 22993 7874
rect 22937 7820 22993 7822
rect 23178 7879 23234 7881
rect 23178 7827 23180 7879
rect 23180 7827 23232 7879
rect 23232 7827 23234 7879
rect 23178 7825 23234 7827
rect 23417 7881 23473 7883
rect 23417 7829 23419 7881
rect 23419 7829 23471 7881
rect 23471 7829 23473 7881
rect 23417 7827 23473 7829
rect 23644 7881 23700 7883
rect 23644 7829 23646 7881
rect 23646 7829 23698 7881
rect 23698 7829 23700 7881
rect 23644 7827 23700 7829
rect 28726 6899 28782 6901
rect 28726 6847 28728 6899
rect 28728 6847 28780 6899
rect 28780 6847 28782 6899
rect 28726 6845 28782 6847
rect 28967 6904 29023 6906
rect 28967 6852 28969 6904
rect 28969 6852 29021 6904
rect 29021 6852 29023 6904
rect 28967 6850 29023 6852
rect 29206 6906 29262 6908
rect 29206 6854 29208 6906
rect 29208 6854 29260 6906
rect 29260 6854 29262 6906
rect 29206 6852 29262 6854
rect 29433 6906 29489 6908
rect 29433 6854 29435 6906
rect 29435 6854 29487 6906
rect 29487 6854 29489 6906
rect 29433 6852 29489 6854
rect 18331 -830 18387 -774
rect 18536 -991 18592 -935
rect 18795 -972 18851 -916
rect 18706 -1534 18762 -1531
rect 18143 -1546 18199 -1544
rect 18143 -1598 18145 -1546
rect 18145 -1598 18197 -1546
rect 18197 -1598 18199 -1546
rect 18143 -1600 18199 -1598
rect 18452 -1593 18504 -1544
rect 18504 -1593 18508 -1544
rect 18706 -1586 18754 -1534
rect 18754 -1586 18762 -1534
rect 18706 -1587 18762 -1586
rect 18452 -1600 18508 -1593
rect 54248 9315 54304 9317
rect 54012 9262 54014 9314
rect 54014 9262 54066 9314
rect 54066 9262 54068 9314
rect 54012 9258 54068 9262
rect 54131 9262 54133 9314
rect 54133 9262 54185 9314
rect 54185 9262 54187 9314
rect 54131 9258 54187 9262
rect 54248 9263 54252 9315
rect 54252 9263 54304 9315
rect 54248 9261 54304 9263
rect 54372 9316 54428 9318
rect 54372 9264 54374 9316
rect 54374 9264 54426 9316
rect 54426 9264 54428 9316
rect 54372 9262 54428 9264
rect 54489 9315 54545 9317
rect 54489 9263 54492 9315
rect 54492 9263 54544 9315
rect 54544 9263 54545 9315
rect 54489 9261 54545 9263
rect 54012 9196 54068 9198
rect 54012 9144 54014 9196
rect 54014 9144 54066 9196
rect 54066 9144 54068 9196
rect 54012 9142 54068 9144
rect 54130 9196 54186 9198
rect 54130 9144 54133 9196
rect 54133 9144 54185 9196
rect 54185 9144 54186 9196
rect 54253 9197 54309 9200
rect 54253 9145 54254 9197
rect 54254 9145 54306 9197
rect 54306 9145 54309 9197
rect 54373 9199 54429 9204
rect 54373 9148 54374 9199
rect 54374 9148 54426 9199
rect 54426 9148 54429 9199
rect 54491 9195 54547 9197
rect 54253 9144 54309 9145
rect 54130 9142 54186 9144
rect 54491 9143 54493 9195
rect 54493 9143 54545 9195
rect 54545 9143 54547 9195
rect 54491 9141 54547 9143
rect 61818 9322 61874 9324
rect 61582 9269 61584 9321
rect 61584 9269 61636 9321
rect 61636 9269 61638 9321
rect 61582 9265 61638 9269
rect 61701 9269 61703 9321
rect 61703 9269 61755 9321
rect 61755 9269 61757 9321
rect 61701 9265 61757 9269
rect 61818 9270 61822 9322
rect 61822 9270 61874 9322
rect 61818 9268 61874 9270
rect 61942 9323 61998 9325
rect 61942 9271 61944 9323
rect 61944 9271 61996 9323
rect 61996 9271 61998 9323
rect 61942 9269 61998 9271
rect 62059 9322 62115 9324
rect 62059 9270 62062 9322
rect 62062 9270 62114 9322
rect 62114 9270 62115 9322
rect 62059 9268 62115 9270
rect 61582 9203 61638 9205
rect 61582 9151 61584 9203
rect 61584 9151 61636 9203
rect 61636 9151 61638 9203
rect 61582 9149 61638 9151
rect 61700 9203 61756 9205
rect 61700 9151 61703 9203
rect 61703 9151 61755 9203
rect 61755 9151 61756 9203
rect 61823 9204 61879 9207
rect 61823 9152 61824 9204
rect 61824 9152 61876 9204
rect 61876 9152 61879 9204
rect 61943 9206 61999 9211
rect 61943 9155 61944 9206
rect 61944 9155 61996 9206
rect 61996 9155 61999 9206
rect 62061 9202 62117 9204
rect 61823 9151 61879 9152
rect 61700 9149 61756 9151
rect 62061 9150 62063 9202
rect 62063 9150 62115 9202
rect 62115 9150 62117 9202
rect 62061 9148 62117 9150
rect 43283 7104 43443 7106
rect 43283 6948 43285 7104
rect 43285 6948 43441 7104
rect 43441 6948 43443 7104
rect 43283 6946 43443 6948
rect 43826 7104 43986 7106
rect 43826 6948 43828 7104
rect 43828 6948 43984 7104
rect 43984 6948 43986 7104
rect 43826 6946 43986 6948
rect 44536 7104 44696 7106
rect 44536 6948 44538 7104
rect 44538 6948 44694 7104
rect 44694 6948 44696 7104
rect 44536 6946 44696 6948
rect 46935 7078 46991 7080
rect 46193 7073 46249 7075
rect 46193 7021 46195 7073
rect 46195 7021 46247 7073
rect 46247 7021 46249 7073
rect 46719 7070 46775 7072
rect 46193 7019 46249 7021
rect 46439 7068 46495 7070
rect 46439 7016 46441 7068
rect 46441 7016 46493 7068
rect 46493 7016 46495 7068
rect 46719 7018 46721 7070
rect 46721 7018 46773 7070
rect 46773 7018 46775 7070
rect 46935 7026 46937 7078
rect 46937 7026 46989 7078
rect 46989 7026 46991 7078
rect 46935 7024 46991 7026
rect 46719 7016 46775 7018
rect 46439 7014 46495 7016
rect 38310 6450 38470 6610
rect 43823 6074 43879 6076
rect 43823 6022 43825 6074
rect 43825 6022 43877 6074
rect 43877 6022 43879 6074
rect 43823 6020 43879 6022
rect 44072 6061 44128 6063
rect 44072 6009 44074 6061
rect 44074 6009 44126 6061
rect 44126 6009 44128 6061
rect 44528 6060 44584 6062
rect 44072 6007 44128 6009
rect 44306 6056 44362 6058
rect 44306 6004 44308 6056
rect 44308 6004 44360 6056
rect 44360 6004 44362 6056
rect 44528 6008 44530 6060
rect 44530 6008 44582 6060
rect 44582 6008 44584 6060
rect 44528 6006 44584 6008
rect 44306 6002 44362 6004
rect 27147 4405 27203 4407
rect 27147 4353 27149 4405
rect 27149 4353 27201 4405
rect 27201 4353 27203 4405
rect 27147 4351 27203 4353
rect 27379 4405 27435 4407
rect 27379 4353 27381 4405
rect 27381 4353 27433 4405
rect 27433 4353 27435 4405
rect 27379 4351 27435 4353
rect 27144 4209 27200 4211
rect 27144 4157 27146 4209
rect 27146 4157 27198 4209
rect 27198 4157 27200 4209
rect 27144 4155 27200 4157
rect 27379 4209 27435 4211
rect 27379 4157 27381 4209
rect 27381 4157 27433 4209
rect 27433 4157 27435 4209
rect 27379 4155 27435 4157
rect 30468 4487 30524 4489
rect 30468 4435 30470 4487
rect 30470 4435 30522 4487
rect 30522 4435 30524 4487
rect 30468 4433 30524 4435
rect 54022 4661 54078 4663
rect 53786 4608 53788 4660
rect 53788 4608 53840 4660
rect 53840 4608 53842 4660
rect 53786 4604 53842 4608
rect 53905 4608 53907 4660
rect 53907 4608 53959 4660
rect 53959 4608 53961 4660
rect 53905 4604 53961 4608
rect 54022 4609 54026 4661
rect 54026 4609 54078 4661
rect 54022 4607 54078 4609
rect 54146 4662 54202 4664
rect 54146 4610 54148 4662
rect 54148 4610 54200 4662
rect 54200 4610 54202 4662
rect 54146 4608 54202 4610
rect 54263 4661 54319 4663
rect 54263 4609 54266 4661
rect 54266 4609 54318 4661
rect 54318 4609 54319 4661
rect 54263 4607 54319 4609
rect 53786 4542 53842 4544
rect 53786 4490 53788 4542
rect 53788 4490 53840 4542
rect 53840 4490 53842 4542
rect 53786 4488 53842 4490
rect 53904 4542 53960 4544
rect 53904 4490 53907 4542
rect 53907 4490 53959 4542
rect 53959 4490 53960 4542
rect 54027 4543 54083 4546
rect 54027 4491 54028 4543
rect 54028 4491 54080 4543
rect 54080 4491 54083 4543
rect 54147 4545 54203 4550
rect 54147 4494 54148 4545
rect 54148 4494 54200 4545
rect 54200 4494 54203 4545
rect 54265 4541 54321 4543
rect 54027 4490 54083 4491
rect 53904 4488 53960 4490
rect 54265 4489 54267 4541
rect 54267 4489 54319 4541
rect 54319 4489 54321 4541
rect 54265 4487 54321 4489
rect 98889 4719 98945 4723
rect 98889 4667 98941 4719
rect 98941 4667 98945 4719
rect 99064 4713 99120 4717
rect 99064 4661 99116 4713
rect 99116 4661 99120 4713
rect 99065 4564 99121 4568
rect 98887 4560 98943 4564
rect 98887 4508 98939 4560
rect 98939 4508 98943 4560
rect 99065 4512 99117 4564
rect 99117 4512 99121 4564
rect 98890 4395 98946 4399
rect 98890 4343 98942 4395
rect 98942 4343 98946 4395
rect 99078 4390 99134 4394
rect 99078 4338 99130 4390
rect 99130 4338 99134 4390
rect 30468 4226 30524 4228
rect 30468 4174 30470 4226
rect 30470 4174 30522 4226
rect 30522 4174 30524 4226
rect 30468 4172 30524 4174
rect 91654 4254 91710 4256
rect 91418 4201 91420 4253
rect 91420 4201 91472 4253
rect 91472 4201 91474 4253
rect 91418 4197 91474 4201
rect 91537 4201 91539 4253
rect 91539 4201 91591 4253
rect 91591 4201 91593 4253
rect 91537 4197 91593 4201
rect 91654 4202 91658 4254
rect 91658 4202 91710 4254
rect 91654 4200 91710 4202
rect 91778 4255 91834 4257
rect 91778 4203 91780 4255
rect 91780 4203 91832 4255
rect 91832 4203 91834 4255
rect 91778 4201 91834 4203
rect 91895 4254 91951 4256
rect 91895 4202 91898 4254
rect 91898 4202 91950 4254
rect 91950 4202 91951 4254
rect 91895 4200 91951 4202
rect 91418 4135 91474 4137
rect 91418 4083 91420 4135
rect 91420 4083 91472 4135
rect 91472 4083 91474 4135
rect 91418 4081 91474 4083
rect 91536 4135 91592 4137
rect 91536 4083 91539 4135
rect 91539 4083 91591 4135
rect 91591 4083 91592 4135
rect 91659 4136 91715 4139
rect 91659 4084 91660 4136
rect 91660 4084 91712 4136
rect 91712 4084 91715 4136
rect 91779 4138 91835 4143
rect 91779 4087 91780 4138
rect 91780 4087 91832 4138
rect 91832 4087 91835 4138
rect 91897 4134 91953 4136
rect 91659 4083 91715 4084
rect 91536 4081 91592 4083
rect 91897 4082 91899 4134
rect 91899 4082 91951 4134
rect 91951 4082 91953 4134
rect 91897 4080 91953 4082
rect 58524 -3015 58580 -3011
rect 58354 -3040 58410 -3036
rect 58354 -3092 58357 -3040
rect 58357 -3092 58409 -3040
rect 58409 -3092 58410 -3040
rect 58524 -3067 58527 -3015
rect 58527 -3067 58579 -3015
rect 58579 -3067 58580 -3015
rect 5142 -3963 5198 -3961
rect 4976 -3976 5032 -3974
rect 4976 -4028 4978 -3976
rect 4978 -4028 5030 -3976
rect 5030 -4028 5032 -3976
rect 5142 -4015 5144 -3963
rect 5144 -4015 5196 -3963
rect 5196 -4015 5198 -3963
rect 5142 -4017 5198 -4015
rect 4976 -4030 5032 -4028
rect 5147 -4103 5203 -4101
rect 4976 -4114 5032 -4112
rect 4976 -4166 4978 -4114
rect 4978 -4166 5030 -4114
rect 5030 -4166 5032 -4114
rect 5147 -4155 5149 -4103
rect 5149 -4155 5201 -4103
rect 5201 -4155 5203 -4103
rect 5147 -4157 5203 -4155
rect 4976 -4168 5032 -4166
rect 5247 -4506 5303 -4504
rect 5081 -4519 5137 -4517
rect 5081 -4571 5083 -4519
rect 5083 -4571 5135 -4519
rect 5135 -4571 5137 -4519
rect 5247 -4558 5249 -4506
rect 5249 -4558 5301 -4506
rect 5301 -4558 5303 -4506
rect 5247 -4560 5303 -4558
rect 5081 -4573 5137 -4571
rect 5252 -4646 5308 -4644
rect 5081 -4657 5137 -4655
rect 5081 -4709 5083 -4657
rect 5083 -4709 5135 -4657
rect 5135 -4709 5137 -4657
rect 5252 -4698 5254 -4646
rect 5254 -4698 5306 -4646
rect 5306 -4698 5308 -4646
rect 5252 -4700 5308 -4698
rect 5081 -4711 5137 -4709
rect 58353 -3214 58409 -3210
rect 58353 -3266 58356 -3214
rect 58356 -3266 58408 -3214
rect 58408 -3266 58409 -3214
rect 58519 -3213 58575 -3209
rect 58519 -3265 58522 -3213
rect 58522 -3265 58574 -3213
rect 58574 -3265 58575 -3213
rect 68218 -3641 68274 -3637
rect 68218 -3693 68270 -3641
rect 68270 -3693 68274 -3641
rect 68392 -3642 68448 -3638
rect 68392 -3694 68444 -3642
rect 68444 -3694 68448 -3642
rect 68219 -3807 68275 -3803
rect 68219 -3859 68271 -3807
rect 68271 -3859 68275 -3807
rect 68417 -3812 68473 -3808
rect 68417 -3864 68469 -3812
rect 68469 -3864 68473 -3812
rect 87132 -4724 87188 -4722
rect 87132 -4776 87136 -4724
rect 87136 -4776 87188 -4724
rect 87132 -4778 87188 -4776
rect 87252 -4724 87308 -4722
rect 87252 -4776 87256 -4724
rect 87256 -4776 87308 -4724
rect 87252 -4778 87308 -4776
rect 87372 -4724 87428 -4722
rect 87372 -4776 87376 -4724
rect 87376 -4776 87428 -4724
rect 87372 -4778 87428 -4776
rect 87132 -4844 87188 -4842
rect 87132 -4896 87136 -4844
rect 87136 -4896 87188 -4844
rect 87132 -4898 87188 -4896
rect 87252 -4844 87308 -4842
rect 87252 -4896 87256 -4844
rect 87256 -4896 87308 -4844
rect 87252 -4898 87308 -4896
rect 87372 -4844 87428 -4842
rect 87372 -4896 87376 -4844
rect 87376 -4896 87428 -4844
rect 87372 -4898 87428 -4896
rect 87134 -4964 87190 -4962
rect 87134 -5016 87136 -4964
rect 87136 -5016 87188 -4964
rect 87188 -5016 87190 -4964
rect 87134 -5018 87190 -5016
rect 87252 -4964 87308 -4962
rect 87252 -5016 87256 -4964
rect 87256 -5016 87308 -4964
rect 87252 -5018 87308 -5016
rect 87372 -4964 87428 -4962
rect 87372 -5016 87376 -4964
rect 87376 -5016 87428 -4964
rect 87372 -5018 87428 -5016
rect 98602 -762 98658 -758
rect 98602 -814 98654 -762
rect 98654 -814 98658 -762
rect 98777 -768 98833 -764
rect 98777 -820 98829 -768
rect 98829 -820 98833 -768
rect 98778 -917 98834 -913
rect 98600 -921 98656 -917
rect 98600 -973 98652 -921
rect 98652 -973 98656 -921
rect 98778 -969 98830 -917
rect 98830 -969 98834 -917
rect 98603 -1086 98659 -1082
rect 98603 -1138 98655 -1086
rect 98655 -1138 98659 -1086
rect 98791 -1091 98847 -1087
rect 98791 -1143 98843 -1091
rect 98843 -1143 98847 -1091
rect 98635 -1966 98691 -1962
rect 98635 -2018 98687 -1966
rect 98687 -2018 98691 -1966
rect 98809 -1967 98865 -1963
rect 98809 -2019 98861 -1967
rect 98861 -2019 98865 -1967
rect 98636 -2132 98692 -2128
rect 98636 -2184 98688 -2132
rect 98688 -2184 98692 -2132
rect 98834 -2137 98890 -2133
rect 98834 -2189 98886 -2137
rect 98886 -2189 98890 -2137
rect 98605 -2863 98661 -2859
rect 98605 -2915 98657 -2863
rect 98657 -2915 98661 -2863
rect 98779 -2864 98835 -2860
rect 98779 -2916 98831 -2864
rect 98831 -2916 98835 -2864
rect 98606 -3029 98662 -3025
rect 98606 -3081 98658 -3029
rect 98658 -3081 98662 -3029
rect 98804 -3034 98860 -3030
rect 98804 -3086 98856 -3034
rect 98856 -3086 98860 -3034
rect 98597 -3346 98653 -3342
rect 98597 -3398 98649 -3346
rect 98649 -3398 98653 -3346
rect 98771 -3347 98827 -3343
rect 98771 -3399 98823 -3347
rect 98823 -3399 98827 -3347
rect 98598 -3512 98654 -3508
rect 98598 -3564 98650 -3512
rect 98650 -3564 98654 -3512
rect 98796 -3517 98852 -3513
rect 98796 -3569 98848 -3517
rect 98848 -3569 98852 -3517
rect 98635 -3898 98691 -3894
rect 98635 -3950 98687 -3898
rect 98687 -3950 98691 -3898
rect 98809 -3899 98865 -3895
rect 98809 -3951 98861 -3899
rect 98861 -3951 98865 -3899
rect 98636 -4064 98692 -4060
rect 98636 -4116 98688 -4064
rect 98688 -4116 98692 -4064
rect 98834 -4069 98890 -4065
rect 98834 -4121 98886 -4069
rect 98886 -4121 98890 -4069
rect 53317 -11368 53373 -11366
rect 53075 -11371 53131 -11369
rect 52806 -11379 52862 -11377
rect 52551 -11381 52607 -11379
rect 52346 -11394 52402 -11392
rect 52346 -11446 52348 -11394
rect 52348 -11446 52400 -11394
rect 52400 -11446 52402 -11394
rect 52551 -11433 52553 -11381
rect 52553 -11433 52605 -11381
rect 52605 -11433 52607 -11381
rect 52806 -11431 52808 -11379
rect 52808 -11431 52860 -11379
rect 52860 -11431 52862 -11379
rect 53075 -11423 53077 -11371
rect 53077 -11423 53129 -11371
rect 53129 -11423 53131 -11371
rect 53317 -11420 53319 -11368
rect 53319 -11420 53371 -11368
rect 53371 -11420 53373 -11368
rect 53317 -11422 53373 -11420
rect 53075 -11425 53131 -11423
rect 52806 -11433 52862 -11431
rect 52551 -11435 52607 -11433
rect 52346 -11448 52402 -11446
rect 53245 -11551 53301 -11549
rect 53032 -11563 53088 -11561
rect 52787 -11566 52843 -11564
rect 52554 -11576 52610 -11574
rect 52348 -11584 52404 -11582
rect 52348 -11636 52350 -11584
rect 52350 -11636 52402 -11584
rect 52402 -11636 52404 -11584
rect 52554 -11628 52556 -11576
rect 52556 -11628 52608 -11576
rect 52608 -11628 52610 -11576
rect 52787 -11618 52789 -11566
rect 52789 -11618 52841 -11566
rect 52841 -11618 52843 -11566
rect 53032 -11615 53034 -11563
rect 53034 -11615 53086 -11563
rect 53086 -11615 53088 -11563
rect 53245 -11603 53247 -11551
rect 53247 -11603 53299 -11551
rect 53299 -11603 53301 -11551
rect 53245 -11605 53301 -11603
rect 53404 -11550 53460 -11548
rect 53404 -11602 53406 -11550
rect 53406 -11602 53458 -11550
rect 53458 -11602 53460 -11550
rect 53404 -11604 53460 -11602
rect 53032 -11617 53088 -11615
rect 52787 -11620 52843 -11618
rect 52554 -11630 52610 -11628
rect 52348 -11638 52404 -11636
rect 53353 -11736 53409 -11734
rect 53155 -11744 53211 -11742
rect 52916 -11754 52972 -11752
rect 52705 -11757 52761 -11755
rect 52339 -11760 52395 -11758
rect 52339 -11812 52341 -11760
rect 52341 -11812 52393 -11760
rect 52393 -11812 52395 -11760
rect 52339 -11814 52395 -11812
rect 52507 -11759 52563 -11757
rect 52507 -11811 52509 -11759
rect 52509 -11811 52561 -11759
rect 52561 -11811 52563 -11759
rect 52705 -11809 52707 -11757
rect 52707 -11809 52759 -11757
rect 52759 -11809 52761 -11757
rect 52916 -11806 52918 -11754
rect 52918 -11806 52970 -11754
rect 52970 -11806 52972 -11754
rect 53155 -11796 53157 -11744
rect 53157 -11796 53209 -11744
rect 53209 -11796 53211 -11744
rect 53353 -11788 53355 -11736
rect 53355 -11788 53407 -11736
rect 53407 -11788 53409 -11736
rect 53353 -11790 53409 -11788
rect 53155 -11798 53211 -11796
rect 52916 -11808 52972 -11806
rect 52705 -11811 52761 -11809
rect 52507 -11813 52563 -11811
<< metal3 >>
rect -3079 62800 -2804 62816
rect -3079 62744 -3052 62800
rect -2996 62798 -2804 62800
rect -2996 62744 -2888 62798
rect -3079 62742 -2888 62744
rect -2832 62742 -2804 62798
rect -3079 62739 -2804 62742
rect -3089 62686 7594 62739
rect -3089 62673 -2886 62686
rect -3089 62617 -3052 62673
rect -2996 62630 -2886 62673
rect -2830 62630 7594 62686
rect -2996 62617 7594 62630
rect -3089 62546 7594 62617
rect -3089 62535 -2881 62546
rect -3089 62487 -3052 62535
rect -3079 62479 -3052 62487
rect -2996 62490 -2881 62535
rect -2825 62490 7594 62546
rect -2996 62487 7594 62490
rect -2996 62479 -2804 62487
rect -3079 62466 -2804 62479
rect -4059 61382 -3685 61414
rect -4059 61372 -2311 61382
rect -4059 61359 -3845 61372
rect -4059 61303 -4011 61359
rect -3955 61316 -3845 61359
rect -3789 61316 -2311 61372
rect -3955 61303 -2311 61316
rect -4059 61232 -2311 61303
rect -4059 61221 -3840 61232
rect -4059 61165 -4011 61221
rect -3955 61176 -3840 61221
rect -3784 61176 -2311 61232
rect -3955 61165 -2311 61176
rect -4059 61157 -2311 61165
rect -4059 61153 -3685 61157
rect -4059 61136 -3689 61153
rect -2118 60500 -1893 60774
rect -2698 52728 -2423 52744
rect -2698 52672 -2671 52728
rect -2615 52726 -2423 52728
rect -2615 52672 -2507 52726
rect -2698 52670 -2507 52672
rect -2451 52670 -2423 52726
rect -2698 52614 -2423 52670
rect -2698 52601 -2505 52614
rect -2698 52545 -2671 52601
rect -2615 52558 -2505 52601
rect -2449 52575 -2423 52614
rect -2449 52558 861 52575
rect -2615 52545 861 52558
rect -2698 52474 861 52545
rect -2698 52463 -2500 52474
rect -2698 52407 -2671 52463
rect -2615 52418 -2500 52463
rect -2444 52418 861 52474
rect -2615 52407 861 52418
rect -2698 52399 861 52407
rect -2698 52394 -2423 52399
rect -3907 52216 -3536 52258
rect -3907 52203 -3693 52216
rect -3907 52147 -3859 52203
rect -3803 52160 -3693 52203
rect -3637 52195 -3536 52216
rect -3637 52160 1088 52195
rect -3803 52147 1088 52160
rect -3907 52076 1088 52147
rect -3907 52065 -3688 52076
rect -3907 52009 -3859 52065
rect -3803 52020 -3688 52065
rect -3632 52020 1088 52076
rect -3803 52009 1088 52020
rect -3907 51994 1088 52009
rect -3907 51980 -3537 51994
rect -2076 51992 -1875 51994
rect -2076 50862 -1875 51119
rect -2388 44202 -2113 44218
rect -2388 44146 -2361 44202
rect -2305 44200 -2113 44202
rect -2305 44146 -2197 44200
rect -2388 44144 -2197 44146
rect -2141 44144 -2113 44200
rect -2388 44088 -2113 44144
rect -2388 44075 -2195 44088
rect -2388 44019 -2361 44075
rect -2305 44032 -2195 44075
rect -2139 44032 -2113 44088
rect -2305 44019 -2113 44032
rect -2388 43948 -2113 44019
rect -2388 43937 -2190 43948
rect -2388 43881 -2361 43937
rect -2305 43892 -2190 43937
rect -2134 43933 -2113 43948
rect 1490 43933 1578 44198
rect -2134 43892 1578 43933
rect -2305 43881 1578 43892
rect -2388 43868 1578 43881
rect -2336 43845 1578 43868
rect -2336 43798 -2269 43845
rect 1490 43798 1578 43845
rect -2381 43661 -2106 43677
rect -2381 43605 -2354 43661
rect -2298 43659 -2106 43661
rect -2298 43605 -2190 43659
rect -2381 43603 -2190 43605
rect -2134 43603 -2106 43659
rect -2381 43547 -2106 43603
rect -2381 43534 -2188 43547
rect -2381 43478 -2354 43534
rect -2298 43491 -2188 43534
rect -2132 43491 -2106 43547
rect -2298 43478 -2106 43491
rect -2381 43407 -2106 43478
rect -2381 43396 -2183 43407
rect -2381 43340 -2354 43396
rect -2298 43351 -2183 43396
rect -2127 43351 -2106 43407
rect -2298 43340 -2106 43351
rect -2381 43327 -2106 43340
rect -2489 36768 -2214 36784
rect -2489 36712 -2462 36768
rect -2406 36766 -2214 36768
rect -2406 36712 -2298 36766
rect -2489 36710 -2298 36712
rect -2242 36710 -2214 36766
rect -2489 36654 -2214 36710
rect -2489 36641 -2296 36654
rect -2489 36585 -2462 36641
rect -2406 36598 -2296 36641
rect -2240 36598 -2214 36654
rect -2406 36585 -2214 36598
rect -2489 36514 -2214 36585
rect -2489 36503 -2291 36514
rect -2489 36447 -2462 36503
rect -2406 36458 -2291 36503
rect -2235 36458 -2214 36514
rect -2406 36447 -2214 36458
rect -2489 36434 -2214 36447
rect 6888 32662 7411 33451
rect -4689 32139 7411 32662
rect -4689 18858 -4166 32139
rect 2010 28027 2740 28118
rect 2010 28019 2607 28027
rect 2010 27963 2041 28019
rect 2097 28016 2417 28019
rect 2097 27963 2220 28016
rect 2010 27960 2220 27963
rect 2276 27963 2417 28016
rect 2473 27971 2607 28019
rect 2663 27971 2740 28027
rect 2473 27963 2740 27971
rect 2276 27960 2740 27963
rect 2010 27892 2740 27960
rect 2010 27836 2044 27892
rect 2100 27884 2607 27892
rect 2100 27881 2409 27884
rect 2100 27836 2220 27881
rect 2010 27825 2220 27836
rect 2276 27828 2409 27881
rect 2465 27836 2607 27884
rect 2663 27836 2740 27892
rect 2465 27828 2740 27836
rect 2276 27825 2740 27828
rect 2010 27720 2740 27825
rect 2011 21918 2709 27720
rect 2011 21777 22718 21918
rect 2011 21757 8980 21777
rect 2011 21701 8765 21757
rect 8821 21721 8980 21757
rect 9036 21721 22718 21777
rect 8821 21701 22718 21721
rect 2011 21604 22718 21701
rect 2011 21594 8916 21604
rect 2011 21538 8654 21594
rect 8710 21548 8916 21594
rect 8972 21548 22718 21604
rect 8710 21538 22718 21548
rect 2011 21353 22718 21538
rect 2011 21343 8892 21353
rect 2011 21287 8672 21343
rect 8728 21297 8892 21343
rect 8948 21297 22718 21353
rect 8728 21287 22718 21297
rect 2011 21220 22718 21287
rect -265 20781 1066 20974
rect -265 20711 20745 20781
rect -265 20691 377 20711
rect -265 20635 162 20691
rect 218 20655 377 20691
rect 433 20655 20745 20711
rect 218 20635 20745 20655
rect -265 20538 20745 20635
rect -265 20528 313 20538
rect -265 20472 51 20528
rect 107 20482 313 20528
rect 369 20482 20745 20538
rect 107 20472 20745 20482
rect -265 20287 20745 20472
rect -265 20277 289 20287
rect -265 20221 69 20277
rect 125 20231 289 20277
rect 345 20231 20745 20287
rect 125 20221 20745 20231
rect -265 20107 20745 20221
rect -265 19888 1066 20107
rect -4689 18335 17883 18858
rect 17360 14316 17883 18335
rect 17360 14180 18261 14316
rect 17360 14160 17795 14180
rect 17360 14104 17580 14160
rect 17636 14124 17795 14160
rect 17851 14124 18261 14180
rect 17636 14112 18261 14124
rect 17636 14104 18056 14112
rect 17360 14056 18056 14104
rect 18112 14056 18261 14112
rect 17360 14007 18261 14056
rect 17360 13997 17731 14007
rect 17360 13941 17469 13997
rect 17525 13951 17731 13997
rect 17787 13951 18261 14007
rect 17525 13945 18261 13951
rect 17525 13941 17920 13945
rect 17360 13889 17920 13941
rect 17976 13889 18261 13945
rect 17360 13756 18261 13889
rect 17360 13746 17707 13756
rect 17360 13690 17487 13746
rect 17543 13700 17707 13746
rect 17763 13700 18261 13756
rect 20071 14104 20745 20107
rect 22020 17766 22718 21220
rect 22020 17741 49711 17766
rect 22020 17109 91956 17741
rect 22020 17094 55075 17109
rect 22020 17068 49711 17094
rect 20071 14094 20480 14104
rect 20071 14038 20260 14094
rect 20316 14048 20480 14094
rect 20536 14048 20745 14104
rect 20316 14038 20745 14048
rect 20071 13905 20745 14038
rect 20071 13849 20251 13905
rect 20307 13899 20745 13905
rect 20307 13849 20478 13899
rect 20071 13843 20478 13849
rect 20534 13843 20745 13899
rect 20071 13708 20745 13843
rect 17543 13695 18261 13700
rect 17543 13690 17924 13695
rect 17360 13639 17924 13690
rect 17980 13639 18261 13695
rect 26035 13671 26139 13672
rect 25430 13657 26202 13671
rect 17360 13551 18261 13639
rect 17360 13495 17705 13551
rect 17761 13495 18261 13551
rect 17360 13289 18261 13495
rect 25426 13618 26202 13657
rect 25426 13562 25520 13618
rect 25576 13562 25708 13618
rect 25764 13562 25903 13618
rect 25959 13562 26202 13618
rect 25426 13428 26202 13562
rect 11365 12714 11683 12801
rect 5394 12708 11683 12714
rect 5394 12652 11399 12708
rect 11455 12705 11683 12708
rect 11455 12652 11583 12705
rect 5394 12649 11583 12652
rect 11639 12649 11683 12705
rect 5394 12580 11683 12649
rect 5394 12524 11396 12580
rect 11452 12572 11683 12580
rect 11452 12524 11581 12572
rect 5394 12516 11581 12524
rect 11637 12516 11683 12572
rect 5394 12461 11683 12516
rect 5394 12458 5607 12461
rect 5394 12402 5434 12458
rect 5490 12405 5607 12458
rect 5663 12435 11683 12461
rect 5663 12405 11397 12435
rect 5490 12402 11397 12405
rect 5394 12379 11397 12402
rect 11453 12379 11574 12435
rect 11630 12379 11683 12435
rect 5394 12363 11683 12379
rect 5394 12267 5745 12363
rect 11365 12334 11683 12363
rect 5394 12211 5433 12267
rect 5489 12265 5745 12267
rect 5489 12211 5594 12265
rect 5394 12209 5594 12211
rect 5650 12209 5745 12265
rect 5394 12132 5745 12209
rect 8578 11667 8996 11732
rect 8578 11664 8873 11667
rect 8578 11663 8727 11664
rect 8578 11607 8607 11663
rect 8663 11608 8727 11663
rect 8783 11611 8873 11664
rect 8929 11611 8996 11667
rect 8783 11608 8996 11611
rect 8663 11607 8996 11608
rect 8578 11552 8996 11607
rect 8578 11496 8612 11552
rect 8668 11496 8743 11552
rect 8799 11496 8883 11552
rect 8939 11496 8996 11552
rect 8578 11488 8996 11496
rect 5268 7566 6063 7709
rect 5268 7562 5729 7566
rect 5268 7546 5590 7562
rect 5268 7490 5393 7546
rect 5449 7506 5590 7546
rect 5646 7510 5729 7562
rect 5785 7562 6063 7566
rect 5785 7510 5873 7562
rect 5646 7506 5873 7510
rect 5929 7506 6063 7562
rect 5449 7490 6063 7506
rect 5268 7442 6063 7490
rect 5268 7428 5852 7442
rect 5268 7421 5678 7428
rect 5268 7416 5505 7421
rect 5268 7360 5356 7416
rect 5412 7365 5505 7416
rect 5561 7372 5678 7421
rect 5734 7386 5852 7428
rect 5908 7386 6063 7442
rect 5734 7372 6063 7386
rect 5561 7365 6063 7372
rect 5412 7360 6063 7365
rect 5268 7313 6063 7360
rect 5268 7308 5941 7313
rect 5268 7304 5639 7308
rect 5268 7296 5476 7304
rect 5268 7240 5325 7296
rect 5381 7248 5476 7296
rect 5532 7252 5639 7304
rect 5695 7252 5800 7308
rect 5856 7257 5941 7308
rect 5997 7257 6063 7313
rect 5856 7252 6063 7257
rect 5532 7248 6063 7252
rect 5381 7240 6063 7248
rect 5268 7226 6063 7240
rect 8648 7137 8897 11488
rect 19634 11244 19861 11247
rect 19622 11197 20513 11244
rect 19622 11195 20148 11197
rect 19622 11190 19909 11195
rect 19622 11134 19668 11190
rect 19724 11139 19909 11190
rect 19965 11141 20148 11195
rect 20204 11141 20375 11197
rect 20431 11141 20513 11197
rect 19965 11139 20513 11141
rect 19724 11134 20513 11139
rect 19622 11090 20513 11134
rect 19634 9198 19861 11090
rect 20286 9198 20513 11090
rect 19580 9187 19979 9198
rect 20206 9187 20513 9198
rect 19580 9151 20513 9187
rect 19580 9149 20106 9151
rect 19580 9144 19867 9149
rect 19580 9088 19626 9144
rect 19682 9093 19867 9144
rect 19923 9095 20106 9149
rect 20162 9095 20333 9151
rect 20389 9095 20513 9151
rect 19923 9093 20513 9095
rect 19682 9088 20513 9093
rect 19580 9044 20513 9088
rect 20286 8003 20513 9044
rect 25973 9080 26202 13428
rect 28727 10002 32041 10065
rect 28718 9902 32041 10002
rect 28718 9900 29262 9902
rect 28718 9895 29023 9900
rect 28718 9839 28782 9895
rect 28838 9844 29023 9895
rect 29079 9846 29262 9900
rect 29318 9846 29489 9902
rect 29545 9846 32041 9902
rect 29079 9844 32041 9846
rect 28838 9839 32041 9844
rect 28718 9814 32041 9839
rect 28718 9777 29681 9814
rect 30509 9080 30918 9085
rect 25973 9032 30918 9080
rect 25973 9019 30667 9032
rect 25973 8963 30535 9019
rect 30591 8976 30667 9019
rect 30723 9031 30918 9032
rect 30723 8976 30792 9031
rect 30591 8975 30792 8976
rect 30848 8975 30918 9031
rect 30591 8963 30918 8975
rect 25973 8922 30918 8963
rect 25973 8906 30665 8922
rect 25973 8851 30532 8906
rect 30355 8850 30532 8851
rect 30588 8866 30665 8906
rect 30721 8866 30792 8922
rect 30848 8866 30918 8922
rect 30588 8850 30918 8866
rect 30355 8795 30918 8850
rect 30355 8793 30654 8795
rect 30355 8737 30529 8793
rect 30585 8739 30654 8793
rect 30710 8739 30792 8795
rect 30848 8739 30918 8795
rect 30585 8737 30918 8739
rect 30355 8672 30918 8737
rect 20286 7955 20641 8003
rect 20286 7883 26699 7955
rect 20286 7881 23417 7883
rect 20286 7876 23178 7881
rect 20286 7820 22937 7876
rect 22993 7825 23178 7876
rect 23234 7827 23417 7881
rect 23473 7827 23644 7883
rect 23700 7827 26699 7883
rect 23234 7825 26699 7827
rect 22993 7820 26699 7825
rect 20286 7728 26699 7820
rect 8560 7075 9108 7137
rect 8560 7068 8951 7075
rect 8560 7012 8590 7068
rect 8646 7012 8731 7068
rect 8787 7019 8951 7068
rect 9007 7019 9108 7075
rect 8787 7012 9108 7019
rect 8560 6958 9108 7012
rect 8560 6902 8596 6958
rect 8652 6953 9108 6958
rect 8652 6902 8737 6953
rect 8560 6897 8737 6902
rect 8793 6897 8977 6953
rect 9033 6897 9108 6953
rect 8560 6879 9108 6897
rect 20318 352 20641 7728
rect 26472 6980 26699 7728
rect 31790 6980 32041 9814
rect 49039 9313 49671 17068
rect 53921 9318 54794 9377
rect 53921 9317 54372 9318
rect 53921 9314 54248 9317
rect 53921 9313 54012 9314
rect 49039 9258 54012 9313
rect 54068 9258 54131 9314
rect 54187 9261 54248 9314
rect 54304 9262 54372 9317
rect 54428 9317 54794 9318
rect 54428 9262 54489 9317
rect 54304 9261 54489 9262
rect 54545 9313 54794 9317
rect 61491 9325 62361 9385
rect 61491 9324 61942 9325
rect 61491 9321 61818 9324
rect 61491 9313 61582 9321
rect 54545 9265 61582 9313
rect 61638 9265 61701 9321
rect 61757 9268 61818 9321
rect 61874 9269 61942 9324
rect 61998 9324 62361 9325
rect 61998 9269 62059 9324
rect 61874 9268 62059 9269
rect 62115 9313 62361 9324
rect 62115 9268 62375 9313
rect 61757 9265 62375 9268
rect 54545 9261 62375 9265
rect 54187 9258 62375 9261
rect 49039 9211 62375 9258
rect 49039 9207 61943 9211
rect 49039 9205 61823 9207
rect 49039 9204 61582 9205
rect 49039 9200 54373 9204
rect 49039 9198 54253 9200
rect 49039 9142 54012 9198
rect 54068 9142 54130 9198
rect 54186 9144 54253 9198
rect 54309 9148 54373 9200
rect 54429 9197 61582 9204
rect 54429 9148 54491 9197
rect 54309 9144 54491 9148
rect 54186 9142 54491 9144
rect 49039 9141 54491 9142
rect 54547 9149 61582 9197
rect 61638 9149 61700 9205
rect 61756 9151 61823 9205
rect 61879 9155 61943 9207
rect 61999 9204 62375 9211
rect 61999 9155 62061 9204
rect 61879 9151 62061 9155
rect 61756 9149 62061 9151
rect 54547 9148 62061 9149
rect 62117 9148 62375 9204
rect 54547 9141 62375 9148
rect 49039 9087 62375 9141
rect 26472 6908 32041 6980
rect 26472 6906 29206 6908
rect 26472 6901 28967 6906
rect 26472 6845 28726 6901
rect 28782 6850 28967 6901
rect 29023 6852 29206 6906
rect 29262 6852 29433 6908
rect 29489 6852 32041 6908
rect 29023 6850 32041 6852
rect 28782 6845 32041 6850
rect 26472 6753 32041 6845
rect 27167 4463 27415 6753
rect 31790 6741 32041 6753
rect 32327 7125 32533 7128
rect 32327 7124 43272 7125
rect 44110 7124 44460 7130
rect 32327 7106 44715 7124
rect 32327 6946 43283 7106
rect 43443 6946 43826 7106
rect 43986 6946 44536 7106
rect 44696 6946 44715 7106
rect 46136 7080 47059 7119
rect 46136 7075 46935 7080
rect 46136 7019 46193 7075
rect 46249 7072 46935 7075
rect 46249 7070 46719 7072
rect 46249 7019 46439 7070
rect 46136 7014 46439 7019
rect 46495 7016 46719 7070
rect 46775 7024 46935 7072
rect 46991 7024 47059 7080
rect 46775 7016 47059 7024
rect 46495 7014 47059 7016
rect 46136 6961 47059 7014
rect 32327 6919 44715 6946
rect 30400 5978 30606 5983
rect 32327 5978 32533 6919
rect 38287 6610 38493 6919
rect 44110 6850 44480 6919
rect 44110 6810 44460 6850
rect 38287 6450 38310 6610
rect 38470 6450 38493 6610
rect 38287 6414 38493 6450
rect 46593 6163 46752 6961
rect 47454 6163 47743 6195
rect 46512 6130 47745 6163
rect 30400 5772 32533 5978
rect 43759 6076 47745 6130
rect 43759 6020 43823 6076
rect 43879 6063 47745 6076
rect 43879 6020 44072 6063
rect 43759 6007 44072 6020
rect 44128 6062 47745 6063
rect 44128 6058 44528 6062
rect 44128 6007 44306 6058
rect 43759 6002 44306 6007
rect 44362 6006 44528 6058
rect 44584 6006 47745 6062
rect 44362 6002 47745 6006
rect 43759 5971 47745 6002
rect 46512 5937 47745 5971
rect 30400 4489 30606 5772
rect 27094 4407 27485 4463
rect 27094 4351 27147 4407
rect 27203 4351 27379 4407
rect 27435 4351 27485 4407
rect 27094 4211 27485 4351
rect 27094 4155 27144 4211
rect 27200 4155 27379 4211
rect 27435 4155 27485 4211
rect 27094 4108 27485 4155
rect 30400 4433 30468 4489
rect 30524 4433 30606 4489
rect 30400 4228 30606 4433
rect 30400 4172 30468 4228
rect 30524 4172 30606 4228
rect 30400 4129 30606 4172
rect 47454 3849 47743 5937
rect 49039 4545 49671 9087
rect 91324 4952 91956 17109
rect 53695 4664 54568 4724
rect 53695 4663 54146 4664
rect 53695 4660 54022 4663
rect 53695 4604 53786 4660
rect 53842 4604 53905 4660
rect 53961 4607 54022 4660
rect 54078 4608 54146 4663
rect 54202 4663 54568 4664
rect 54202 4608 54263 4663
rect 54078 4607 54263 4608
rect 54319 4607 54568 4663
rect 53961 4604 54568 4607
rect 53695 4550 54568 4604
rect 53695 4546 54147 4550
rect 53695 4545 54027 4546
rect 49039 4544 54027 4545
rect 49039 4488 53786 4544
rect 53842 4488 53904 4544
rect 53960 4490 54027 4544
rect 54083 4494 54147 4546
rect 54203 4545 54568 4550
rect 91324 4723 99215 4952
rect 91324 4667 98889 4723
rect 98945 4717 99215 4723
rect 98945 4667 99064 4717
rect 91324 4661 99064 4667
rect 99120 4661 99215 4717
rect 91324 4568 99215 4661
rect 91324 4564 99065 4568
rect 54203 4543 57420 4545
rect 54203 4494 54265 4543
rect 54083 4490 54265 4494
rect 53960 4488 54265 4490
rect 49039 4487 54265 4488
rect 54321 4487 57420 4543
rect 49039 4319 57420 4487
rect 49039 4304 49671 4319
rect 49161 4303 49588 4304
rect 49161 3849 49588 3854
rect 47454 3560 49588 3849
rect 17589 29 20641 352
rect 4778 -988 5148 -932
rect 4778 -1044 4826 -988
rect 4882 -990 5148 -988
rect 4882 -1044 4990 -990
rect 4778 -1046 4990 -1044
rect 5046 -1004 5148 -990
rect 5046 -1046 15958 -1004
rect 4778 -1102 15958 -1046
rect 4778 -1115 4992 -1102
rect 4778 -1171 4826 -1115
rect 4882 -1158 4992 -1115
rect 5048 -1158 15958 -1102
rect 4882 -1171 15958 -1158
rect 4778 -1242 15958 -1171
rect 4778 -1253 4997 -1242
rect 4778 -1309 4826 -1253
rect 4882 -1298 4997 -1253
rect 5053 -1298 15958 -1242
rect 4882 -1309 15958 -1298
rect 4778 -1321 15958 -1309
rect 4778 -1338 5148 -1321
rect 4844 -1554 14921 -1512
rect 4844 -1567 5058 -1554
rect 4844 -1623 4892 -1567
rect 4948 -1610 5058 -1567
rect 5114 -1610 14921 -1554
rect 4948 -1623 14921 -1610
rect 4844 -1694 14921 -1623
rect 4844 -1705 5063 -1694
rect 4844 -1761 4892 -1705
rect 4948 -1750 5063 -1705
rect 5119 -1750 14921 -1694
rect 4948 -1756 14921 -1750
rect 4948 -1761 5222 -1756
rect 4844 -1773 5222 -1761
rect 4844 -1790 5214 -1773
rect 14677 -2260 14921 -1756
rect 15641 -1813 15958 -1321
rect 17649 -1459 17851 29
rect 18284 -774 21310 -725
rect 18284 -830 18331 -774
rect 18387 -830 21310 -774
rect 18284 -916 21310 -830
rect 18284 -935 18795 -916
rect 18284 -991 18536 -935
rect 18592 -972 18795 -935
rect 18851 -972 21310 -916
rect 18592 -991 21310 -972
rect 18284 -1061 21310 -991
rect 20974 -1269 21310 -1061
rect 17649 -1531 18861 -1459
rect 17649 -1544 18706 -1531
rect 17649 -1600 18143 -1544
rect 18199 -1600 18452 -1544
rect 18508 -1587 18706 -1544
rect 18762 -1587 18861 -1531
rect 18508 -1600 18861 -1587
rect 17649 -1661 18861 -1600
rect 20974 -1605 26713 -1269
rect 15641 -2130 25855 -1813
rect 24985 -2260 25196 -2248
rect 14677 -2504 25212 -2260
rect 5001 -2623 5379 -2608
rect 4971 -2650 24848 -2623
rect 4971 -2663 5215 -2650
rect 4971 -2719 5049 -2663
rect 5105 -2706 5215 -2663
rect 5271 -2706 24848 -2650
rect 5105 -2719 24848 -2706
rect 4971 -2774 24848 -2719
rect 5001 -2790 5379 -2774
rect 5001 -2801 5220 -2790
rect 5001 -2857 5049 -2801
rect 5105 -2846 5220 -2801
rect 5276 -2846 5379 -2790
rect 5105 -2857 5379 -2846
rect 5001 -2869 5379 -2857
rect 5001 -2886 5371 -2869
rect 4975 -3026 16639 -2983
rect 4905 -3068 16639 -3026
rect 4905 -3081 5119 -3068
rect 4905 -3137 4953 -3081
rect 5009 -3124 5119 -3081
rect 5175 -3124 16639 -3068
rect 5009 -3137 16639 -3124
rect 4905 -3208 16639 -3137
rect 4905 -3219 5124 -3208
rect 4905 -3275 4953 -3219
rect 5009 -3264 5124 -3219
rect 5180 -3232 16639 -3208
rect 5180 -3264 5283 -3232
rect 5009 -3275 5283 -3264
rect 4905 -3287 5283 -3275
rect 4905 -3304 5275 -3287
rect 4882 -3462 5260 -3440
rect 4882 -3482 16212 -3462
rect 4882 -3495 5096 -3482
rect 4882 -3551 4930 -3495
rect 4986 -3538 5096 -3495
rect 5152 -3538 16212 -3482
rect 4986 -3551 16212 -3538
rect 4882 -3622 16212 -3551
rect 4882 -3633 5101 -3622
rect 4882 -3689 4930 -3633
rect 4986 -3678 5101 -3633
rect 5157 -3643 16212 -3622
rect 5157 -3678 5260 -3643
rect 4986 -3689 5260 -3678
rect 4882 -3701 5260 -3689
rect 4882 -3718 5252 -3701
rect 5001 -3919 7452 -3878
rect 4928 -3961 7452 -3919
rect 4928 -3974 5142 -3961
rect 4928 -4030 4976 -3974
rect 5032 -4017 5142 -3974
rect 5198 -4017 7452 -3961
rect 5032 -4030 7452 -4017
rect 4928 -4101 7452 -4030
rect 4928 -4112 5147 -4101
rect 4928 -4168 4976 -4112
rect 5032 -4157 5147 -4112
rect 5203 -4103 7452 -4101
rect 5203 -4157 5306 -4103
rect 5032 -4168 5306 -4157
rect 4928 -4180 5306 -4168
rect 4928 -4197 5298 -4180
rect 7227 -4372 7452 -4103
rect 5070 -4462 6102 -4418
rect 5033 -4504 6102 -4462
rect 5033 -4517 5247 -4504
rect 5033 -4573 5081 -4517
rect 5137 -4560 5247 -4517
rect 5303 -4560 6102 -4504
rect 5137 -4573 6102 -4560
rect 5033 -4630 6102 -4573
rect 5033 -4644 5411 -4630
rect 5033 -4655 5252 -4644
rect 5033 -4711 5081 -4655
rect 5137 -4700 5252 -4655
rect 5308 -4700 5411 -4644
rect 5137 -4711 5411 -4700
rect 5033 -4723 5411 -4711
rect 5033 -4740 5403 -4723
rect 16031 -5048 16212 -3643
rect 16390 -5174 16639 -3232
rect 24697 -5269 24848 -2774
rect 24985 -5303 25196 -2504
rect 25538 -3786 25855 -2130
rect 26377 -2241 26713 -1605
rect 49161 -1981 49588 3560
rect 57127 213 57420 4319
rect 91324 4508 98887 4564
rect 98943 4512 99065 4564
rect 99121 4512 99215 4568
rect 98943 4508 99215 4512
rect 91324 4399 99215 4508
rect 91324 4343 98890 4399
rect 98946 4394 99215 4399
rect 98946 4343 99078 4394
rect 91324 4338 99078 4343
rect 99134 4338 99215 4394
rect 91324 4320 99215 4338
rect 91324 4257 92059 4320
rect 98838 4305 99160 4320
rect 91324 4256 91778 4257
rect 91324 4253 91654 4256
rect 91324 4197 91418 4253
rect 91474 4197 91537 4253
rect 91593 4200 91654 4253
rect 91710 4201 91778 4256
rect 91834 4256 92059 4257
rect 91834 4201 91895 4256
rect 91710 4200 91895 4201
rect 91951 4200 92059 4256
rect 91593 4197 92059 4200
rect 91324 4143 92059 4197
rect 91324 4139 91779 4143
rect 91324 4137 91659 4139
rect 91324 4081 91418 4137
rect 91474 4081 91536 4137
rect 91592 4083 91659 4137
rect 91715 4087 91779 4139
rect 91835 4136 92059 4143
rect 91835 4087 91897 4136
rect 91715 4083 91897 4087
rect 91592 4081 91897 4083
rect 91324 4080 91897 4081
rect 91953 4080 92059 4136
rect 91324 4051 92059 4080
rect 91324 4026 91956 4051
rect 55465 -151 57420 213
rect 26377 -2577 36376 -2241
rect 49161 -2408 51945 -1981
rect 25538 -4103 32240 -3786
rect 31923 -5255 32240 -4103
rect 36040 -6541 36376 -2577
rect 51518 -4201 51945 -2408
rect 51284 -4246 52067 -4201
rect 51284 -4273 51585 -4246
rect 51284 -4329 51344 -4273
rect 51400 -4302 51585 -4273
rect 51641 -4277 52067 -4246
rect 51641 -4302 51860 -4277
rect 51400 -4329 51860 -4302
rect 51284 -4333 51860 -4329
rect 51916 -4333 52067 -4277
rect 51284 -4396 52067 -4333
rect 51284 -4415 51571 -4396
rect 51284 -4471 51328 -4415
rect 51384 -4452 51571 -4415
rect 51627 -4427 52067 -4396
rect 51627 -4452 51833 -4427
rect 51384 -4471 51833 -4452
rect 51284 -4483 51833 -4471
rect 51889 -4483 52067 -4427
rect 51284 -4573 52067 -4483
rect 51284 -4577 51559 -4573
rect 51284 -4633 51313 -4577
rect 51369 -4629 51559 -4577
rect 51615 -4577 52067 -4573
rect 51615 -4629 51867 -4577
rect 51369 -4633 51867 -4629
rect 51923 -4633 52067 -4577
rect 51284 -4719 52067 -4633
rect 36093 -14454 36324 -6662
rect 52279 -11322 53565 -11166
rect 52279 -11366 53571 -11322
rect 52279 -11369 53317 -11366
rect 52279 -11377 53075 -11369
rect 52279 -11379 52806 -11377
rect 52279 -11392 52551 -11379
rect 52279 -11448 52346 -11392
rect 52402 -11435 52551 -11392
rect 52607 -11433 52806 -11379
rect 52862 -11425 53075 -11377
rect 53131 -11422 53317 -11369
rect 53373 -11422 53571 -11366
rect 53131 -11425 53571 -11422
rect 52862 -11433 53571 -11425
rect 52607 -11435 53571 -11433
rect 52402 -11448 53571 -11435
rect 52279 -11479 53571 -11448
rect 55465 -11479 55829 -151
rect 98561 -757 98873 -742
rect 56983 -758 98873 -757
rect 56983 -814 98602 -758
rect 98658 -764 98873 -758
rect 98658 -814 98777 -764
rect 56983 -820 98777 -814
rect 98833 -820 98873 -764
rect 56983 -913 98873 -820
rect 56983 -917 98778 -913
rect 56983 -973 98600 -917
rect 98656 -969 98778 -917
rect 98834 -969 98873 -913
rect 98656 -973 98873 -969
rect 56983 -1082 98873 -973
rect 56983 -1138 98603 -1082
rect 98659 -1087 98873 -1082
rect 98659 -1138 98791 -1087
rect 56983 -1143 98791 -1138
rect 98847 -1143 98873 -1087
rect 56983 -1181 98873 -1143
rect 56983 -1186 98866 -1181
rect 56983 -5243 57309 -1186
rect 67147 -1962 98964 -1936
rect 67147 -2018 98635 -1962
rect 98691 -1963 98964 -1962
rect 98691 -2018 98809 -1963
rect 67147 -2019 98809 -2018
rect 98865 -2019 98964 -1963
rect 67147 -2128 98964 -2019
rect 67147 -2184 98636 -2128
rect 98692 -2133 98964 -2128
rect 98692 -2184 98834 -2133
rect 67147 -2189 98834 -2184
rect 98890 -2189 98964 -2133
rect 67147 -2230 98964 -2189
rect 58351 -2964 58627 -2793
rect 58344 -3011 58627 -2964
rect 58344 -3036 58524 -3011
rect 58344 -3092 58354 -3036
rect 58410 -3067 58524 -3036
rect 58580 -3067 58627 -3011
rect 58410 -3092 58627 -3067
rect 58344 -3209 58627 -3092
rect 58344 -3210 58519 -3209
rect 58344 -3266 58353 -3210
rect 58409 -3265 58519 -3210
rect 58575 -3265 58627 -3209
rect 58409 -3266 58627 -3265
rect 58344 -3325 58627 -3266
rect 58351 -3328 58627 -3325
rect 58377 -5154 58602 -3328
rect 67147 -4968 67396 -2230
rect 98546 -2859 98907 -2850
rect 98546 -2905 98605 -2859
rect 75818 -2915 98605 -2905
rect 98661 -2860 98907 -2859
rect 98661 -2915 98779 -2860
rect 75818 -2916 98779 -2915
rect 98835 -2916 98907 -2860
rect 75818 -3025 98907 -2916
rect 75818 -3081 98606 -3025
rect 98662 -3030 98907 -3025
rect 98662 -3081 98804 -3030
rect 75818 -3086 98804 -3081
rect 98860 -3086 98907 -3030
rect 75818 -3114 98907 -3086
rect 68159 -3635 68520 -3628
rect 68156 -3637 68691 -3635
rect 68156 -3661 68218 -3637
rect 68107 -3683 68218 -3661
rect 67579 -3693 68218 -3683
rect 68274 -3638 68691 -3637
rect 68274 -3693 68392 -3638
rect 67579 -3694 68392 -3693
rect 68448 -3694 68691 -3638
rect 67579 -3803 68691 -3694
rect 67579 -3854 68219 -3803
rect 67579 -5030 67750 -3854
rect 68107 -3859 68219 -3854
rect 68275 -3808 68691 -3803
rect 68275 -3859 68417 -3808
rect 68107 -3864 68417 -3859
rect 68473 -3864 68691 -3808
rect 68107 -3886 68691 -3864
rect 68156 -3911 68691 -3886
rect 57040 -5346 57252 -5243
rect 68640 -5267 69133 -5096
rect 75848 -5104 75996 -3114
rect 98546 -3118 98907 -3114
rect 76086 -3342 98994 -3305
rect 76086 -3398 98597 -3342
rect 98653 -3343 98994 -3342
rect 98653 -3398 98771 -3343
rect 76086 -3399 98771 -3398
rect 98827 -3399 98994 -3343
rect 76086 -3508 98994 -3399
rect 76086 -3564 98598 -3508
rect 98654 -3513 98994 -3508
rect 98654 -3564 98796 -3513
rect 76086 -3569 98796 -3564
rect 98852 -3569 98994 -3513
rect 76086 -3614 98994 -3569
rect 75883 -5179 75961 -5104
rect 76158 -5181 76323 -3614
rect 98576 -3892 98937 -3885
rect 83093 -3894 99108 -3892
rect 83093 -3950 98635 -3894
rect 98691 -3895 99108 -3894
rect 98691 -3950 98809 -3895
rect 83093 -3951 98809 -3950
rect 98865 -3951 99108 -3895
rect 83093 -4060 99108 -3951
rect 83093 -4116 98636 -4060
rect 98692 -4065 99108 -4060
rect 98692 -4116 98834 -4065
rect 83093 -4121 98834 -4116
rect 98890 -4121 99108 -4065
rect 83093 -4168 99108 -4121
rect 83093 -5156 83369 -4168
rect 87090 -4722 87760 -4550
rect 87090 -4778 87132 -4722
rect 87188 -4778 87252 -4722
rect 87308 -4778 87372 -4722
rect 87428 -4778 87760 -4722
rect 87090 -4842 87760 -4778
rect 87090 -4898 87132 -4842
rect 87188 -4898 87252 -4842
rect 87308 -4898 87372 -4842
rect 87428 -4898 87760 -4842
rect 87090 -4962 87760 -4898
rect 87090 -5018 87134 -4962
rect 87190 -5018 87252 -4962
rect 87308 -5018 87372 -4962
rect 87428 -5018 87760 -4962
rect 87090 -5090 87760 -5018
rect 52279 -11548 55829 -11479
rect 52279 -11549 53404 -11548
rect 52279 -11561 53245 -11549
rect 52279 -11564 53032 -11561
rect 52279 -11574 52787 -11564
rect 52279 -11582 52554 -11574
rect 52279 -11638 52348 -11582
rect 52404 -11630 52554 -11582
rect 52610 -11620 52787 -11574
rect 52843 -11617 53032 -11564
rect 53088 -11605 53245 -11561
rect 53301 -11604 53404 -11549
rect 53460 -11604 55829 -11548
rect 53301 -11605 55829 -11604
rect 53088 -11617 55829 -11605
rect 52843 -11620 55829 -11617
rect 52610 -11630 55829 -11620
rect 52404 -11638 55829 -11630
rect 52279 -11734 55829 -11638
rect 52279 -11742 53353 -11734
rect 52279 -11752 53155 -11742
rect 52279 -11755 52916 -11752
rect 52279 -11757 52705 -11755
rect 52279 -11758 52507 -11757
rect 52279 -11814 52339 -11758
rect 52395 -11813 52507 -11758
rect 52563 -11811 52705 -11757
rect 52761 -11808 52916 -11755
rect 52972 -11798 53155 -11752
rect 53211 -11790 53353 -11742
rect 53409 -11790 55829 -11734
rect 53211 -11798 55829 -11790
rect 52972 -11808 55829 -11798
rect 52761 -11811 55829 -11808
rect 52563 -11813 55829 -11811
rect 52395 -11814 55829 -11813
rect 52279 -11843 55829 -11814
rect 52279 -11848 53571 -11843
rect 87243 -14434 87474 -5992
rect 34855 -14685 36324 -14454
rect 78405 -14665 87474 -14434
<< via3 >>
rect 5434 12402 5490 12458
rect 5607 12405 5663 12461
rect 5433 12211 5489 12267
rect 5594 12209 5650 12265
rect 5393 7490 5449 7546
rect 5590 7506 5646 7562
rect 5729 7510 5785 7566
rect 5873 7506 5929 7562
rect 5356 7360 5412 7416
rect 5505 7365 5561 7421
rect 5678 7372 5734 7428
rect 5852 7386 5908 7442
rect 5325 7240 5381 7296
rect 5476 7248 5532 7304
rect 5639 7252 5695 7308
rect 5800 7252 5856 7308
rect 5941 7257 5997 7313
rect 51344 -4329 51400 -4273
rect 51585 -4302 51641 -4246
rect 51860 -4333 51916 -4277
rect 51328 -4471 51384 -4415
rect 51571 -4452 51627 -4396
rect 51833 -4483 51889 -4427
rect 51313 -4633 51369 -4577
rect 51559 -4629 51615 -4573
rect 51867 -4633 51923 -4577
<< metal4 >>
rect -7940 41508 -7091 41515
rect -7940 41159 -2689 41508
rect -7940 40575 -2522 41159
rect -7940 -27439 -7091 40575
rect 5385 12461 5993 29177
rect 27663 28397 28023 28607
rect 27811 28389 28023 28397
rect 5385 12458 5607 12461
rect 5385 12402 5434 12458
rect 5490 12405 5607 12458
rect 5663 12405 5993 12461
rect 5490 12402 5993 12405
rect 5385 12267 5993 12402
rect 5385 12211 5433 12267
rect 5489 12265 5993 12267
rect 5489 12211 5594 12265
rect 5385 12209 5594 12211
rect 5650 12209 5993 12265
rect 5385 7709 5993 12209
rect 5268 7566 6063 7709
rect 5268 7562 5729 7566
rect 5268 7546 5590 7562
rect 5268 7490 5393 7546
rect 5449 7506 5590 7546
rect 5646 7510 5729 7562
rect 5785 7562 6063 7566
rect 5785 7510 5873 7562
rect 5646 7506 5873 7510
rect 5929 7506 6063 7562
rect 5449 7490 6063 7506
rect 5268 7442 6063 7490
rect 5268 7428 5852 7442
rect 5268 7421 5678 7428
rect 5268 7416 5505 7421
rect 5268 7360 5356 7416
rect 5412 7365 5505 7416
rect 5561 7372 5678 7421
rect 5734 7386 5852 7428
rect 5908 7386 6063 7442
rect 5734 7372 6063 7386
rect 5561 7365 6063 7372
rect 5412 7360 6063 7365
rect 5268 7313 6063 7360
rect 5268 7308 5941 7313
rect 5268 7304 5639 7308
rect 5268 7296 5476 7304
rect 5268 7240 5325 7296
rect 5381 7248 5476 7296
rect 5532 7252 5639 7304
rect 5695 7252 5800 7308
rect 5856 7257 5941 7308
rect 5997 7257 6063 7313
rect 5856 7252 6063 7257
rect 5532 7248 6063 7252
rect 5381 7240 6063 7248
rect 5268 7226 6063 7240
rect 5385 -5287 5993 7226
rect 51271 -4204 52095 -4173
rect 27683 -4246 64047 -4204
rect 27683 -4273 51585 -4246
rect 27683 -4329 51344 -4273
rect 51400 -4302 51585 -4273
rect 51641 -4277 64047 -4246
rect 51641 -4302 51860 -4277
rect 51400 -4329 51860 -4302
rect 27683 -4333 51860 -4329
rect 51916 -4333 64047 -4277
rect 27683 -4396 64047 -4333
rect 27683 -4415 51571 -4396
rect 27683 -4471 51328 -4415
rect 51384 -4452 51571 -4415
rect 51627 -4427 64047 -4396
rect 51627 -4452 51833 -4427
rect 51384 -4471 51833 -4452
rect 27683 -4483 51833 -4471
rect 51889 -4483 64047 -4427
rect 27683 -4573 64047 -4483
rect 27683 -4577 51559 -4573
rect 27683 -4633 51313 -4577
rect 51369 -4629 51559 -4577
rect 51615 -4577 64047 -4573
rect 51615 -4629 51867 -4577
rect 51369 -4633 51867 -4629
rect 51923 -4633 64047 -4577
rect 27683 -4719 64047 -4633
rect 5385 -5895 8343 -5287
rect 39445 -6852 59430 -6272
rect 11279 -27389 12128 -26499
rect 21483 -27389 22332 -26499
rect 11279 -27439 22332 -27389
rect -7940 -27686 22332 -27439
rect 28864 -27686 29713 -26251
rect 62449 -27498 66334 -26649
rect 62449 -27686 63298 -27498
rect -7940 -28288 63298 -27686
rect 21483 -28535 63298 -28288
rect 65485 -27544 66334 -27498
rect 72203 -27544 73052 -26649
rect 65485 -27594 73052 -27544
rect 80015 -27594 80864 -26550
rect 65485 -28393 80864 -27594
rect 72203 -28443 80864 -28393
<< metal5 >>
rect 27811 28210 28023 28746
rect 95916 21264 96692 22542
rect 95916 20488 98134 21264
rect 97352 20450 98134 20488
rect 97352 118 98128 20450
rect 87362 -658 98128 118
use 7b_divider_magic  7b_divider_magic_0
timestamp 1697518002
transform 1 0 57381 0 1 -16876
box -441 -10214 40218 12749
use 7b_divider_magic  7b_divider_magic_1
timestamp 1697518002
transform 0 -1 9619 -1 0 62378
box -441 -10214 40218 12749
use 7b_divider_magic  7b_divider_magic_2
timestamp 1697518002
transform 1 0 6231 0 1 -16896
box -441 -10214 40218 12749
use A_MUX  A_MUX_0
timestamp 1697518002
transform 1 0 42495 0 1 4782
box -285 -452 3979 2227
use A_MUX  A_MUX_1
timestamp 1697518002
transform 1 0 18282 0 -1 12510
box -285 -452 3979 2227
use A_MUX  A_MUX_2
timestamp 1697518002
transform 1 0 18240 0 1 7818
box -285 -452 3979 2227
use A_MUX  A_MUX_3
timestamp 1697518002
transform -1 0 30924 0 -1 11425
box -285 -452 3979 2227
use A_MUX  A_MUX_4
timestamp 1697518002
transform -1 0 30867 0 -1 8419
box -285 -452 3979 2227
use A_MUX  A_MUX_5
timestamp 1697518002
transform 1 0 16712 0 1 -3124
box -285 -452 3979 2227
use A_MUX  A_MUX_6
timestamp 1697518002
transform 1 0 36417 0 -1 12138
box -285 -452 3979 2227
use cap_11p  cap_11p_0
timestamp 1697518002
transform 1 0 94240 0 1 13088
box -26450 -13708 -6739 632
use cap_240p  cap_240p_0
timestamp 1697518021
transform 1 0 89483 0 -1 28277
box -68140 -68970 6839 8429
use CP_1  CP_1_0
timestamp 1697518002
transform 1 0 33105 0 1 10459
box -1133 -1188 2101 1774
use Current_Mirror_Top  Current_Mirror_Top_0
timestamp 1697518002
transform -1 0 2228 0 1 10249
box -1992 -209 4486 7070
use INV_2  INV_2_0
timestamp 1697518002
transform 1 0 11673 0 1 7901
box 21 -485 1081 648
use INV_2  INV_2_1
timestamp 1697518002
transform 1 0 11228 0 1 13239
box 21 -485 1081 648
use PFD_T2  PFD_T2_0
timestamp 1697518002
transform 1 0 22661 0 1 8437
box -28 -113 4062 3793
use RES_74k  RES_74k_1
timestamp 1697518002
transform -1 0 51462 0 -1 12102
box 3672 -1094 9598 4966
use Tappered_Buffer  Tappered_Buffer_0
timestamp 1697518002
transform 1 0 50570 0 1 3553
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_1
timestamp 1697518002
transform 1 0 50390 0 1 8230
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_2
timestamp 1697518002
transform 1 0 58351 0 1 8237
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_4
timestamp 1697518002
transform -1 0 94996 0 1 3197
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_5
timestamp 1697518002
transform 1 0 48878 0 -1 -10328
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_6
timestamp 1697518002
transform -1 0 4941 0 1 26954
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_7
timestamp 1697518002
transform -1 0 11108 0 1 10738
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_8
timestamp 1697518002
transform -1 0 12287 0 1 6101
box -161 -3147 5956 876
use VCO_DFF_C  VCO_DFF_C_0
timestamp 1697518002
transform 1 0 24282 0 1 -1600
box 0 -27 23932 7170
<< labels >>
flabel metal1 s 1578 15993 1578 15993 0 FreeSans 600 180 0 0 G_source_up
port 1 nsew
flabel metal1 s 1382 15902 1382 15902 0 FreeSans 600 180 0 0 G_source_dn
port 2 nsew
flabel metal1 s 1916 15531 1916 15531 0 FreeSans 600 180 0 0 G_sink_up
port 3 nsew
flabel metal1 s 1919 15268 1919 15268 0 FreeSans 600 180 0 0 G_sink_dn
port 4 nsew
flabel metal1 s 22036 6756 22036 6756 0 FreeSans 2000 0 0 0 S3
port 5 nsew
flabel metal1 s 21788 13207 21788 13207 0 FreeSans 2000 0 0 0 S2
port 6 nsew
flabel metal1 s 19290 14218 19290 14218 0 FreeSans 2000 0 0 0 S1
port 7 nsew
flabel metal1 s 17988 6714 17988 6714 0 FreeSans 2000 0 0 0 S6
port 8 nsew
flabel metal1 s 21995 13993 21995 13993 0 FreeSans 2000 0 0 0 UP_INPUT
port 9 nsew
flabel metal1 s 21858 13590 21858 13590 0 FreeSans 2000 0 0 0 DN_INPUT
port 10 nsew
flabel metal1 s 18022 14399 18022 14399 0 FreeSans 2000 0 0 0 F_IN
port 11 nsew
flabel metal1 s 32279 5743 32279 5743 0 FreeSans 2000 0 0 0 VCTRL2
port 12 nsew
flabel metal1 s 33470 8331 33470 8331 0 FreeSans 2000 0 0 0 VSS
port 13 nsew
flabel metal1 s 30024 14122 30024 14122 0 FreeSans 2000 0 0 0 VDD
port 14 nsew
flabel metal1 s 42870 4240 42870 4240 0 FreeSans 2000 0 0 0 VCTRL_IN
port 15 nsew
flabel metal1 s 43370 4280 43370 4280 0 FreeSans 2000 0 0 0 S4
port 16 nsew
flabel metal1 s 26249 11574 26249 11574 0 FreeSans 2000 0 0 0 UP1
port 17 nsew
flabel metal1 s 26214 8908 26214 8908 0 FreeSans 2000 0 0 0 DN1
port 18 nsew
flabel metal1 s 22703 16344 22703 16344 0 FreeSans 2000 0 0 0 LF_OFFCHIP
port 19 nsew
flabel metal1 s 22694 16690 22694 16690 0 FreeSans 2000 0 0 0 S5
port 20 nsew
flabel metal1 s 56568 6749 56568 6749 0 FreeSans 2000 0 0 0 OUTB
port 21 nsew
flabel metal1 s 56817 2078 56817 2078 0 FreeSans 2000 0 0 0 OUT
port 22 nsew
flabel metal1 s 99070 -7610 99070 -7610 0 FreeSans 2000 0 0 0 OUT1
port 23 nsew
flabel metal1 s 99167 -991 99167 -991 0 FreeSans 2000 0 0 0 D16
port 24 nsew
flabel metal1 s 99137 -2090 99137 -2090 0 FreeSans 2000 0 0 0 D13
port 25 nsew
flabel metal1 s 99090 -2966 99090 -2966 0 FreeSans 2000 0 0 0 D12
port 26 nsew
flabel metal1 s 99146 -3471 99146 -3471 0 FreeSans 2000 0 0 0 D14
port 27 nsew
flabel metal1 s 99171 -4022 99171 -4022 0 FreeSans 2000 0 0 0 D15
port 28 nsew
flabel metal1 s 4423 -2365 4423 -2365 0 FreeSans 2000 0 0 0 S7
port 29 nsew
flabel metal1 s 4793 -4573 4793 -4573 0 FreeSans 2000 0 0 0 D4
port 30 nsew
flabel metal1 s 4742 -4063 4742 -4063 0 FreeSans 2000 0 0 0 D6
port 31 nsew
flabel metal1 s 4675 -3537 4675 -3537 0 FreeSans 2000 0 0 0 D1
port 32 nsew
flabel metal1 s 4723 -3078 4723 -3078 0 FreeSans 2000 0 0 0 D5
port 33 nsew
flabel metal1 s 4752 -2715 4752 -2715 0 FreeSans 2000 0 0 0 D0
port 34 nsew
flabel metal1 s 4646 -1595 4646 -1595 0 FreeSans 2000 0 0 0 D2
port 35 nsew
flabel metal1 s 4579 -1155 4579 -1155 0 FreeSans 2000 0 0 0 D3
port 36 nsew
flabel metal1 s -3298 62608 -3298 62608 0 FreeSans 2000 0 0 0 D11
port 37 nsew
flabel metal1 s -3395 52547 -3395 52547 0 FreeSans 2000 0 0 0 D8
port 38 nsew
flabel metal1 s -3154 44010 -3154 44010 0 FreeSans 2000 0 0 0 D7
port 39 nsew
flabel metal1 s -3184 43467 -3184 43467 0 FreeSans 2000 0 0 0 D9
port 40 nsew
flabel metal1 s -3049 36634 -3049 36634 0 FreeSans 2000 0 0 0 D10
port 41 nsew
flabel metal1 s -3814 24857 -3814 24857 0 FreeSans 2000 0 0 0 PRE_SCALAR
port 42 nsew
flabel metal1 s 4188 9245 4188 9245 0 FreeSans 2000 0 0 0 UP_OUT
port 43 nsew
flabel metal1 s 5730 4634 5730 4634 0 FreeSans 2000 0 0 0 DN_OUT
port 44 nsew
flabel metal2 s 21999 15127 21999 15127 0 FreeSans 2000 0 0 0 UP
port 45 nsew
flabel metal2 s 22016 14545 22016 14545 0 FreeSans 2000 0 0 0 DN
port 46 nsew
flabel metal1 s 99365 4556 99365 4556 0 FreeSans 2000 0 0 0 VDD_TEST
port 47 nsew
flabel metal1 s 39830 6510 39830 6510 0 FreeSans 2000 0 0 0 VCTRL_OBV
port 48 nsew
flabel metal1 s 18550 7330 18550 7330 0 FreeSans 2000 0 0 0 DIV_OUT2
port 49 nsew
flabel metal1 s 13110 -7700 13110 -7700 0 FreeSans 2000 0 0 0 Q02
port 50 nsew
flabel metal1 s 13860 -10180 13860 -10180 0 FreeSans 2000 0 0 0 Q07
port 51 nsew
flabel metal1 s 28770 -7800 28770 -7800 0 FreeSans 2000 0 0 0 Q01
port 52 nsew
flabel metal1 s 14210 -15910 14210 -15910 0 FreeSans 2000 0 0 0 Q05
port 53 nsew
flabel metal1 s 13110 -12310 13110 -12310 0 FreeSans 2000 0 0 0 Q06
port 54 nsew
flabel metal1 s 28860 -12250 28860 -12250 0 FreeSans 2000 0 0 0 Q03
port 55 nsew
flabel metal1 s 28010 -15010 28010 -15010 0 FreeSans 2000 0 0 0 Q04
port 56 nsew
flabel metal1 s 28920 -18000 28920 -18000 0 FreeSans 2000 0 0 0 P02
port 57 nsew
flabel metal1 s 6410 -8020 6410 -8020 0 FreeSans 2000 0 0 0 LD0
port 58 nsew
flabel metal1 s 43780 -18390 43780 -18390 0 FreeSans 2000 0 0 0 OUT01
port 59 nsew
flabel metal1 s 95190 -18410 95190 -18410 0 FreeSans 4000 0 0 0 OUT11
port 60 nsew
flabel metal1 s 57550 -8180 57550 -8180 0 FreeSans 4000 0 0 0 LD1
port 61 nsew
flabel metal1 s 64250 -7650 64250 -7650 0 FreeSans 4000 0 0 0 Q12
port 62 nsew
flabel metal1 s 79910 -7950 79910 -7950 0 FreeSans 4000 0 0 0 Q11
port 63 nsew
flabel metal1 s 64260 -11900 64260 -11900 0 FreeSans 4000 0 0 0 Q16
port 64 nsew
flabel metal1 s 80010 -12090 80010 -12090 0 FreeSans 4000 0 0 0 Q13
port 65 nsew
flabel metal1 s 65360 -15960 65360 -15960 0 FreeSans 4000 0 0 0 Q15
port 66 nsew
flabel metal1 s 79160 -15880 79160 -15880 0 FreeSans 4000 0 0 0 Q14
port 67 nsew
flabel metal1 s 65000 -10230 65000 -10230 0 FreeSans 4000 0 0 0 Q17
port 68 nsew
flabel metal1 s 80070 -17980 80070 -17980 0 FreeSans 4000 0 0 0 P12
port 69 nsew
flabel metal1 s 58470 -2667 58470 -2667 0 FreeSans 4000 0 0 0 D17G
port 70 nsew
flabel metal1 s 69038 -3769 69038 -3769 0 FreeSans 4000 0 0 0 D16G
port 71 nsew
flabel metal1 s -4324 61270 -4324 61270 0 FreeSans 4000 0 0 0 D27G
port 72 nsew
flabel metal1 s -4077 52130 -4077 52130 0 FreeSans 4000 0 0 0 D26G
port 73 nsew
flabel metal1 s 8667 22935 8667 22935 0 FreeSans 4000 0 0 0 OUT21
port 74 nsew
flabel metal1 s 4687 55482 4687 55482 0 FreeSans 4000 0 0 0 Q26
port 75 nsew
flabel metal1 s 2862 54749 2862 54749 0 FreeSans 4000 0 0 0 Q27
port 76 nsew
flabel metal1 s 8628 54398 8628 54398 0 FreeSans 4000 0 0 0 Q25
port 77 nsew
flabel metal1 s -561 55487 -561 55487 0 FreeSans 4000 0 0 0 Q22
port 78 nsew
flabel metal1 s -1095 48432 -1095 48432 0 FreeSans 4000 0 0 0 LD2
port 79 nsew
flabel metal1 s 137 39812 137 39812 0 FreeSans 4000 0 0 0 Q21
port 80 nsew
flabel metal1 s 4469 39744 4469 39744 0 FreeSans 4000 0 0 0 Q23
port 81 nsew
flabel metal1 s 7673 40583 7673 40583 0 FreeSans 4000 0 0 0 Q24
port 82 nsew
flabel metal1 s 48873 -14249 48873 -14249 0 FreeSans 2000 0 0 0 DIV_OUT
port 83 nsew
flabel metal1 s 2488 10382 2488 10382 0 FreeSans 2000 0 0 0 ITAIL
port 84 nsew
flabel metal1 s 5149 16633 5149 16633 0 FreeSans 2000 0 0 0 ITAIL_SRC
port 85 nsew
flabel metal1 s 5143 15231 5143 15231 0 FreeSans 2000 0 0 0 ITAIL_SINK
port 86 nsew
flabel metal1 s 53770 15520 53770 15520 0 FreeSans 2000 0 0 0 A1
port 87 nsew
flabel metal2 s 2480 16670 2480 16670 0 FreeSans 2000 0 0 0 A0
port 88 nsew
flabel metal2 s 2530 15190 2530 15190 0 FreeSans 2000 0 0 0 A3
port 89 nsew
flabel metal2 s 2100 14450 2100 14450 0 FreeSans 2000 0 0 0 G1_2
port 90 nsew
flabel metal2 s 1230 14410 1230 14410 0 FreeSans 2000 0 0 0 SD0_1
port 91 nsew
flabel metal2 s 1970 11950 1970 11950 0 FreeSans 2000 0 0 0 SD2_1
port 92 nsew
flabel metal1 s 1720 10740 1720 10740 0 FreeSans 2000 0 0 0 G2_1
port 93 nsew
flabel metal2 s 940 13900 940 13900 0 FreeSans 2000 0 0 0 G1_1
port 94 nsew
flabel metal2 s -170 15280 -170 15280 0 FreeSans 2000 0 0 0 SD01
port 95 nsew
<< properties >>
string GDS_END 15057316
string GDS_FILE PLL_TOP_MUX_7-t.gds
string GDS_START 14927958
<< end >>
