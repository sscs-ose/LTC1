magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1050 -1081 1050 1081
<< metal1 >>
rect -50 75 50 81
rect -50 49 -44 75
rect -18 49 18 75
rect 44 49 50 75
rect -50 13 50 49
rect -50 -13 -44 13
rect -18 -13 18 13
rect 44 -13 50 13
rect -50 -49 50 -13
rect -50 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 50 -49
rect -50 -81 50 -75
<< via1 >>
rect -44 49 -18 75
rect 18 49 44 75
rect -44 -13 -18 13
rect 18 -13 44 13
rect -44 -75 -18 -49
rect 18 -75 44 -49
<< metal2 >>
rect -50 75 50 81
rect -50 49 -44 75
rect -18 49 18 75
rect 44 49 50 75
rect -50 13 50 49
rect -50 -13 -44 13
rect -18 -13 18 13
rect 44 -13 50 13
rect -50 -49 50 -13
rect -50 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 50 -49
rect -50 -81 50 -75
<< end >>
