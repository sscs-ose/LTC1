magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1046 -1073 1046 1073
<< metal1 >>
rect -46 67 46 73
rect -46 41 -40 67
rect -14 41 14 67
rect 40 41 46 67
rect -46 13 46 41
rect -46 -13 -40 13
rect -14 -13 14 13
rect 40 -13 46 13
rect -46 -41 46 -13
rect -46 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 46 -41
rect -46 -73 46 -67
<< via1 >>
rect -40 41 -14 67
rect 14 41 40 67
rect -40 -13 -14 13
rect 14 -13 40 13
rect -40 -67 -14 -41
rect 14 -67 40 -41
<< metal2 >>
rect -46 67 46 73
rect -46 41 -40 67
rect -14 41 14 67
rect 40 41 46 67
rect -46 13 46 41
rect -46 -13 -40 13
rect -14 -13 14 13
rect 40 -13 46 13
rect -46 -41 46 -13
rect -46 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 46 -41
rect -46 -73 46 -67
<< end >>
