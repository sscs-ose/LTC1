magic
tech gf180mcuC
magscale 1 10
timestamp 1695306401
<< metal1 >>
rect 399 1612 436 1649
rect 2650 1607 2726 1656
rect 139 1506 199 1561
rect 1267 1504 1327 1559
rect 3300 1504 3534 1553
rect 4425 1513 4462 1550
rect 49 -978 116 991
rect 3689 675 3726 712
rect 957 451 1004 498
rect 2096 448 2156 503
rect 4322 498 4399 503
rect 4322 446 4334 498
rect 4386 446 4399 498
rect 4322 442 4399 446
rect 3377 161 3564 162
rect 3377 11 3732 161
rect 1129 -5 1304 11
rect 3545 10 3732 11
rect 2259 -4 2423 6
rect 4309 -49 4391 -46
rect 4309 -58 4323 -49
rect 1931 -138 2007 -89
rect 3439 -102 4323 -58
rect 4375 -102 4391 -49
rect 3439 -108 4391 -102
rect 3439 -340 3492 -108
rect 4309 -113 4391 -108
rect 2091 -444 2151 -442
rect 966 -502 1026 -447
rect 2091 -497 2159 -444
rect 3439 -495 3491 -340
rect 2099 -499 2159 -497
rect 1402 -1037 1571 -956
rect 3438 -1368 3491 -495
rect 146 -1558 206 -1503
rect 3438 -1504 3490 -1368
rect 1267 -1563 1327 -1508
rect 3301 -1545 3490 -1504
rect 3301 -1554 3489 -1545
<< via1 >>
rect 4334 446 4386 498
rect 4323 -102 4375 -49
<< metal2 >>
rect 313 -737 377 739
rect 2567 347 2627 743
rect 4322 498 4399 503
rect 4322 446 4334 498
rect 4386 446 4399 498
rect 4322 442 4399 446
rect 2567 337 2643 347
rect 2567 281 2577 337
rect 2633 281 2643 337
rect 2567 271 2643 281
rect 4328 -46 4391 442
rect 4309 -49 4391 -46
rect 4309 -102 4323 -49
rect 4375 -102 4391 -49
rect 4309 -113 4391 -102
rect 2567 -283 2643 -274
rect 2567 -339 2577 -283
rect 2633 -339 2643 -283
rect 2567 -350 2643 -339
rect 2567 -746 2627 -350
<< via2 >>
rect 2577 281 2633 337
rect 2577 -339 2633 -283
<< metal3 >>
rect 2567 337 2643 347
rect 2567 281 2577 337
rect 2633 281 2643 337
rect 2567 271 2643 281
rect 2567 -274 2627 271
rect 2567 -283 2643 -274
rect 2567 -339 2577 -283
rect 2633 -339 2643 -283
rect 2567 -350 2643 -339
use mux_2x1_ibr  mux_2x1_ibr_0
timestamp 1695127730
transform 1 0 3377 0 1 1051
box 0 -1051 1135 1051
use mux_4x1_ibr  mux_4x1_ibr_0
timestamp 1695306401
transform 1 0 1194 0 1 -5
box -1194 5 2193 2107
use mux_4x1_ibr  mux_4x1_ibr_1
timestamp 1695306401
transform 1 0 1194 0 -1 5
box -1194 5 2193 2107
<< labels >>
flabel metal1 984 -474 984 -474 0 FreeSans 640 0 0 0 I0
port 0 nsew
flabel metal1 169 -1539 169 -1539 0 FreeSans 640 0 0 0 I1
port 1 nsew
flabel metal1 2110 -474 2110 -474 0 FreeSans 640 0 0 0 I2
port 2 nsew
flabel metal1 1299 -1535 1299 -1535 0 FreeSans 640 0 0 0 I3
port 3 nsew
flabel metal1 979 476 979 476 0 FreeSans 640 0 0 0 I4
port 4 nsew
flabel metal1 169 1537 169 1537 0 FreeSans 640 0 0 0 I5
port 5 nsew
flabel metal1 2106 476 2106 476 0 FreeSans 640 0 0 0 I6
port 6 nsew
flabel metal1 1299 1532 1299 1532 0 FreeSans 640 0 0 0 I7
port 7 nsew
flabel metal1 1489 -993 1489 -993 0 FreeSans 640 0 0 0 VSS
port 8 nsew
flabel metal1 1966 -117 1966 -117 0 FreeSans 640 0 0 0 VDD
port 9 nsew
flabel metal1 4445 1528 4445 1528 0 FreeSans 640 0 0 0 OUT
port 10 nsew
flabel metal1 414 1634 414 1634 0 FreeSans 640 0 0 0 S0
port 11 nsew
flabel metal1 2675 1634 2675 1634 0 FreeSans 640 0 0 0 S1
port 12 nsew
flabel metal1 3713 689 3713 689 0 FreeSans 640 0 0 0 S2
port 13 nsew
<< end >>
