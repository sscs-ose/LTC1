magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3068 -2128 3068 2128
<< nwell >>
rect -1068 -128 1068 128
<< nsubdiff >>
rect -985 23 985 45
rect -985 -23 -963 23
rect 963 -23 985 23
rect -985 -45 985 -23
<< nsubdiffcont >>
rect -963 -23 963 23
<< metal1 >>
rect -974 23 974 34
rect -974 -23 -963 23
rect 963 -23 974 23
rect -974 -34 974 -23
<< end >>
