* NGSPICE file created from AND_flat.ext - technology: gf180mcuC

.subckt AND_flat VDD VSS B A OUT
X0 OUT Inverter_0.IN VSS.t1 VSS.t0 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X1 Inverter_0.IN B.t0 a_250_78# VSS.t2 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 OUT Inverter_0.IN VDD.t1 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X3 a_250_78# A.t0 VSS.t4 VSS.t3 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X4 VDD B.t1 Inverter_0.IN VDD.t2 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X5 Inverter_0.IN A.t1 VDD.t6 VDD.t5 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 VSS.n3 VSS.t2 1563.68
R1 VSS.n3 VSS.t3 1533.02
R2 VSS.n1 VSS.n0 996.279
R3 VSS.n0 VSS.t0 455.748
R4 VSS.n6 VSS.t1 8.96939
R5 VSS VSS.t4 6.91394
R6 VSS VSS.n1 2.6005
R7 VSS.n5 VSS.n4 2.6005
R8 VSS.n4 VSS.n3 2.6005
R9 VSS.n4 VSS.n2 1.72653
R10 VSS.n6 VSS.n5 0.400161
R11 VSS VSS.n6 0.0689956
R12 VSS.n5 VSS 0.0142288
R13 OUT.n2 OUT.n1 9.02722
R14 OUT.n2 OUT.n0 6.48941
R15 OUT OUT.n2 0.130713
R16 B B.n0 33.3896
R17 B.n0 B.t1 31.5469
R18 B.n0 B.t0 12.6451
R19 VDD.n5 VDD.t2 443.255
R20 VDD.t2 VDD.n4 432.548
R21 VDD.n5 VDD.t5 421.842
R22 VDD.n4 VDD 315.707
R23 VDD.n4 VDD.t0 116.338
R24 VDD VDD.t6 6.73971
R25 VDD.n1 VDD.n0 6.57115
R26 VDD.n3 VDD.t1 6.40636
R27 VDD.n6 VDD.n2 4.2005
R28 VDD.n7 VDD.n6 3.1505
R29 VDD.n6 VDD.n5 3.1505
R30 VDD.n7 VDD.n1 0.219398
R31 VDD.n3 VDD.n1 0.145855
R32 VDD VDD.n7 0.0432119
R33 VDD VDD.n3 0.0353691
R34 A.n0 A.t0 31.938
R35 A.n2 A.n0 28.718
R36 A.n0 A.t1 12.2541
R37 A A.n2 4.00671
R38 A.n2 A.n1 0.503948
C0 a_250_78# A 8.64e-19
C1 VDD B 0.226f
C2 VDD Inverter_0.IN 0.574f
C3 VDD OUT 0.124f
C4 Inverter_0.IN B 0.124f
C5 B OUT 2.17e-19
C6 Inverter_0.IN OUT 0.113f
C7 VDD A 0.249f
C8 B A 0.104f
C9 Inverter_0.IN A 0.00979f
C10 OUT A 1.57e-20
C11 VDD a_250_78# 0.00253f
C12 B a_250_78# 0.155f
C13 Inverter_0.IN a_250_78# 0.0608f
C14 B VSS 0.414f
C15 A VSS 0.296f
C16 a_250_78# VSS 0.188f
C17 OUT VSS 0.177f
C18 Inverter_0.IN VSS 0.418f
C19 VDD VSS 2.01f
.ends

