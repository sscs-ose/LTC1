* NGSPICE file created from A_MUX_flat.ext - technology: gf180mcuC

.subckt A_MUX_pex VDD VSS IN1 IN2 SEL OUT 
X0 OUT SEL.t0 IN2.t5 VSS.t10 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1 VSS SEL.t1 Tr_Gate_1.CLK.t6 VSS.t16 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X2 VSS SEL.t2 Tr_Gate_1.CLK.t5 VSS.t13 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X3 Tr_Gate_1.CLK SEL.t3 VDD.t35 VDD.t22 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X4 Tr_Gate_1.CLK SEL.t4 VSS.t12 VSS.t11 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X5 VDD SEL.t5 Tr_Gate_1.CLK.t10 VDD.t19 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X6 OUT a_2663_557.t6 IN1.t3 VDD.t9 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X7 VDD SEL.t6 Tr_Gate_1.CLK.t9 VDD.t16 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X8 IN2 SEL.t7 OUT.t10 VSS.t7 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X9 OUT a_2663_557.t7 IN1.t2 VDD.t7 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X10 VDD SEL.t8 a_268_897.t5 VDD.t28 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X11 IN1 a_2663_557.t8 OUT.t7 VDD.t4 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X12 Tr_Gate_1.CLK SEL.t9 VDD.t27 VDD.t13 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X13 OUT SEL.t10 IN2.t4 VSS.t5 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X14 VDD Tr_Gate_1.CLK.t12 a_2663_557.t5 VDD.t1 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X15 IN1 a_2663_557.t9 OUT.t1 VDD.t1 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X16 IN1 Tr_Gate_1.CLK.t13 OUT.t13 VSS.t19 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X17 OUT SEL.t11 IN2.t3 VSS.t10 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X18 IN1 Tr_Gate_1.CLK.t15 OUT.t14 VSS.t0 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X19 VDD SEL.t12 a_268_897.t4 VDD.t3 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X20 OUT Tr_Gate_1.CLK.t16 IN1.t5 VSS.t1 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X21 OUT a_268_897.t6 IN2.t0 VDD.t0 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X22 IN2 a_268_897.t7 OUT.t15 VDD.t28 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X23 Tr_Gate_1.CLK SEL.t14 VDD.t23 VDD.t22 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X24 VDD SEL.t15 Tr_Gate_1.CLK.t8 VDD.t19 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X25 VSS SEL.t16 a_268_897.t1 VSS.t7 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X26 VDD SEL.t17 Tr_Gate_1.CLK.t7 VDD.t16 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X27 OUT a_268_897.t8 IN2.t1 VDD.t2 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X28 IN2 a_268_897.t9 OUT.t3 VDD.t3 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X29 Tr_Gate_1.CLK SEL.t20 VDD.t14 VDD.t13 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X30 VSS Tr_Gate_1.CLK.t17 a_2663_557.t1 VSS.t19 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X31 IN1 Tr_Gate_1.CLK.t19 OUT.t4 VSS.t0 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X32 VDD Tr_Gate_1.CLK.t20 a_2663_557.t2 VDD.t4 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X33 Tr_Gate_1.CLK SEL.t21 VSS.t4 VSS.t3 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
R0 SEL.n14 SEL.t0 45.6363
R1 SEL.n0 SEL.t13 29.6446
R2 SEL.t12 SEL.n1 29.6446
R3 SEL.n2 SEL.t16 24.6117
R4 SEL.n8 SEL.t15 23.6945
R5 SEL.n9 SEL.t14 23.6945
R6 SEL.n1 SEL.n0 22.2047
R7 SEL.t0 SEL.t11 22.1925
R8 SEL.n15 SEL.n14 20.9314
R9 SEL.n9 SEL.n8 18.8035
R10 SEL SEL.t12 18.5175
R11 SEL.n6 SEL.n3 15.8172
R12 SEL.n12 SEL.n11 15.8172
R13 SEL.n11 SEL.n3 15.8172
R14 SEL.t5 SEL.n6 14.8925
R15 SEL.t9 SEL.n3 14.8925
R16 SEL.n11 SEL.t6 14.8925
R17 SEL.n10 SEL.n4 12.2457
R18 SEL.n10 SEL.n5 12.2457
R19 SEL.n7 SEL.n5 12.2457
R20 SEL.n13 SEL.t3 11.6285
R21 SEL.t15 SEL.n7 8.9065
R22 SEL.t20 SEL.n5 8.9065
R23 SEL.n10 SEL.t17 8.9065
R24 SEL.t14 SEL.n4 8.9065
R25 SEL.n6 SEL.t1 8.6145
R26 SEL.n3 SEL.t4 8.6145
R27 SEL.n11 SEL.t2 8.6145
R28 SEL.n12 SEL.t21 8.59715
R29 SEL.n7 SEL.t5 8.3225
R30 SEL.n5 SEL.t9 8.3225
R31 SEL.t6 SEL.n10 8.3225
R32 SEL.n4 SEL.t3 8.3225
R33 SEL.n2 SEL.t18 6.1325
R34 SEL.n0 SEL.t8 6.1325
R35 SEL.n1 SEL.t19 6.1325
R36 SEL.n14 SEL.t7 6.1325
R37 SEL.n15 SEL.t10 6.1325
R38 SEL.n16 SEL.n15 4.86779
R39 SEL.n18 SEL.n2 4.79907
R40 SEL SEL.n13 4.223
R41 SEL.n8 SEL.t20 3.6505
R42 SEL.t17 SEL.n9 3.6505
R43 SEL.n13 SEL.n12 3.1807
R44 SEL.n16 SEL 2.68257
R45 SEL SEL.n18 0.640368
R46 SEL.n17 SEL 0.1655
R47 SEL.n17 SEL.n16 0.109537
R48 SEL.n18 SEL.n17 0.0592755
R49 IN2.n3 IN2.n2 5.81586
R50 IN2.n5 IN2.t3 5.10208
R51 IN2.n8 IN2.t5 5.10194
R52 IN2.n4 IN2.t0 5.08021
R53 IN2.n8 IN2.n7 4.66114
R54 IN2.n3 IN2.n1 2.85093
R55 IN2.n1 IN2.t1 2.16717
R56 IN2.n1 IN2.n0 2.16717
R57 IN2.n7 IN2.t4 1.9505
R58 IN2.n7 IN2.n6 1.9505
R59 IN2.n4 IN2.n3 0.644196
R60 IN2.n5 IN2.n4 0.449473
R61 IN2.n9 IN2.n8 0.21214
R62 IN2.n9 IN2.n5 0.198571
R63 IN2 IN2.n9 0.0718949
R64 OUT.n24 OUT.t13 6.74332
R65 OUT.n7 OUT.n6 6.74326
R66 OUT.n9 OUT.n8 5.1005
R67 OUT.n25 OUT.t14 5.1005
R68 OUT.n4 OUT.n1 3.57508
R69 OUT.n18 OUT.n17 3.56654
R70 OUT.n7 OUT.t10 3.40075
R71 OUT.n24 OUT.n23 3.40011
R72 OUT.n26 OUT.t4 3.00158
R73 OUT.n10 OUT.n5 3.00032
R74 OUT.n13 OUT 2.60907
R75 OUT.n22 OUT.n15 2.41287
R76 OUT.n13 OUT.n12 2.36206
R77 OUT.n30 OUT.n13 2.30849
R78 OUT.n29 OUT.n22 2.26352
R79 OUT.n3 OUT.t15 2.16717
R80 OUT.n3 OUT.n2 2.16717
R81 OUT.n1 OUT.t3 2.16717
R82 OUT.n1 OUT.n0 2.16717
R83 OUT.n17 OUT.t1 2.16717
R84 OUT.n17 OUT.n16 2.16717
R85 OUT.n15 OUT.t7 2.16717
R86 OUT.n15 OUT.n14 2.16717
R87 OUT.n11 OUT.n10 1.84797
R88 OUT.n27 OUT.n26 1.82978
R89 OUT.n4 OUT.n3 1.25233
R90 OUT.n11 OUT.n4 1.12574
R91 OUT.n12 OUT 0.751569
R92 OUT OUT.n30 0.736653
R93 OUT.n10 OUT.n9 0.446259
R94 OUT.n26 OUT.n25 0.445613
R95 OUT.n30 OUT.n29 0.366541
R96 OUT.n12 OUT.n11 0.33941
R97 OUT.n25 OUT.n24 0.11326
R98 OUT.n9 OUT.n7 0.112615
R99 OUT.n19 OUT.n18 0.0556613
R100 OUT.n20 OUT.n19 0.0382419
R101 OUT.n21 OUT.n20 0.0324355
R102 OUT.n22 OUT.n21 0.0208226
R103 OUT.n29 OUT.n28 0.0160394
R104 OUT.n28 OUT.n27 0.0132434
R105 VSS.n244 VSS.n243 209.026
R106 VSS.n197 VSS.t7 162.114
R107 VSS.n109 VSS.t19 146.444
R108 VSS.n27 VSS.n26 142.726
R109 VSS.n117 VSS.t1 100.198
R110 VSS.n158 VSS.t16 91.2286
R111 VSS.n117 VSS.n116 87.3523
R112 VSS.n186 VSS.t5 84.9174
R113 VSS.n4 VSS.n3 79.6448
R114 VSS.n126 VSS.t0 69.3681
R115 VSS.n298 VSS.t10 66.9047
R116 VSS.n151 VSS.t11 57.018
R117 VSS.n216 VSS.n215 47.576
R118 VSS.n173 VSS.t3 45.6145
R119 VSS.n284 VSS.n283 25.7329
R120 VSS.n97 VSS.n96 10.2772
R121 VSS.t0 VSS.n125 10.2772
R122 VSS.n141 VSS.n2 6.65541
R123 VSS.n314 VSS.t4 6.65541
R124 VSS.n11 VSS.n10 5.2005
R125 VSS.n134 VSS.n133 5.2005
R126 VSS.n136 VSS.n135 5.2005
R127 VSS.n13 VSS.n12 5.2005
R128 VSS.n310 VSS.n168 5.2005
R129 VSS.n309 VSS.n169 5.2005
R130 VSS.n307 VSS.n193 5.2005
R131 VSS.n306 VSS.n305 5.2005
R132 VSS.n305 VSS.n304 5.2005
R133 VSS.n303 VSS.n302 5.2005
R134 VSS.n302 VSS.n301 5.2005
R135 VSS.n128 VSS.n9 4.88533
R136 VSS.n128 VSS.n127 4.5005
R137 VSS.n127 VSS.n126 4.5005
R138 VSS.n300 VSS.n299 4.5005
R139 VSS.n299 VSS.n298 4.5005
R140 VSS.n196 VSS.n195 3.95358
R141 VSS.n325 VSS.t13 3.80167
R142 VSS.n154 VSS.n1 3.37941
R143 VSS.n1 VSS.t12 3.2765
R144 VSS.n1 VSS.n0 3.2765
R145 VSS.n127 VSS.n13 2.9883
R146 VSS.n56 VSS.n55 2.6005
R147 VSS.n55 VSS.n54 2.6005
R148 VSS.n53 VSS.n52 2.6005
R149 VSS.n52 VSS.n51 2.6005
R150 VSS.n50 VSS.n49 2.6005
R151 VSS.n49 VSS.n48 2.6005
R152 VSS.n47 VSS.n46 2.6005
R153 VSS.n46 VSS.n45 2.6005
R154 VSS.n44 VSS.n43 2.6005
R155 VSS.n43 VSS.n42 2.6005
R156 VSS.n41 VSS.n40 2.6005
R157 VSS.n40 VSS.n39 2.6005
R158 VSS.n38 VSS.n37 2.6005
R159 VSS.n37 VSS.n36 2.6005
R160 VSS.n35 VSS.n34 2.6005
R161 VSS.n34 VSS.n33 2.6005
R162 VSS.n32 VSS.n31 2.6005
R163 VSS.n31 VSS.n30 2.6005
R164 VSS.n77 VSS.n76 2.6005
R165 VSS.n76 VSS.n75 2.6005
R166 VSS.n74 VSS.n73 2.6005
R167 VSS.n73 VSS.n72 2.6005
R168 VSS.n71 VSS.n70 2.6005
R169 VSS.n70 VSS.n69 2.6005
R170 VSS.n68 VSS.n67 2.6005
R171 VSS.n67 VSS.n66 2.6005
R172 VSS.n65 VSS.n64 2.6005
R173 VSS.n64 VSS.n63 2.6005
R174 VSS.n62 VSS.n61 2.6005
R175 VSS.n61 VSS.n60 2.6005
R176 VSS.n59 VSS.n58 2.6005
R177 VSS.n58 VSS.n57 2.6005
R178 VSS.n95 VSS.n94 2.6005
R179 VSS.n91 VSS.n90 2.6005
R180 VSS.n88 VSS.n87 2.6005
R181 VSS.n85 VSS.n84 2.6005
R182 VSS.n82 VSS.n81 2.6005
R183 VSS.n80 VSS.n79 2.6005
R184 VSS.n29 VSS.n28 2.6005
R185 VSS.n28 VSS.n27 2.6005
R186 VSS.n25 VSS.n24 2.6005
R187 VSS.n24 VSS.n23 2.6005
R188 VSS.n22 VSS.n21 2.6005
R189 VSS.n21 VSS.n20 2.6005
R190 VSS.n19 VSS.n18 2.6005
R191 VSS.n18 VSS.n17 2.6005
R192 VSS.n16 VSS.n15 2.6005
R193 VSS.n15 VSS.n14 2.6005
R194 VSS.n208 VSS.n207 2.6005
R195 VSS.n207 VSS.n206 2.6005
R196 VSS.n211 VSS.n210 2.6005
R197 VSS.n210 VSS.n209 2.6005
R198 VSS.n214 VSS.n213 2.6005
R199 VSS.n213 VSS.n212 2.6005
R200 VSS.n218 VSS.n217 2.6005
R201 VSS.n217 VSS.n216 2.6005
R202 VSS.n248 VSS.n247 2.6005
R203 VSS.n221 VSS.n220 2.6005
R204 VSS.n220 VSS.n219 2.6005
R205 VSS.n224 VSS.n223 2.6005
R206 VSS.n223 VSS.n222 2.6005
R207 VSS.n227 VSS.n226 2.6005
R208 VSS.n226 VSS.n225 2.6005
R209 VSS.n230 VSS.n229 2.6005
R210 VSS.n229 VSS.n228 2.6005
R211 VSS.n233 VSS.n232 2.6005
R212 VSS.n232 VSS.n231 2.6005
R213 VSS.n236 VSS.n235 2.6005
R214 VSS.n235 VSS.n234 2.6005
R215 VSS.n239 VSS.n238 2.6005
R216 VSS.n238 VSS.n237 2.6005
R217 VSS.n242 VSS.n241 2.6005
R218 VSS.n241 VSS.n240 2.6005
R219 VSS.n246 VSS.n245 2.6005
R220 VSS.n251 VSS.n250 2.6005
R221 VSS.n250 VSS.n249 2.6005
R222 VSS.n254 VSS.n253 2.6005
R223 VSS.n253 VSS.n252 2.6005
R224 VSS.n257 VSS.n256 2.6005
R225 VSS.n256 VSS.n255 2.6005
R226 VSS.n260 VSS.n259 2.6005
R227 VSS.n259 VSS.n258 2.6005
R228 VSS.n263 VSS.n262 2.6005
R229 VSS.n262 VSS.n261 2.6005
R230 VSS.n266 VSS.n265 2.6005
R231 VSS.n265 VSS.n264 2.6005
R232 VSS.n268 VSS.n267 2.6005
R233 VSS.n271 VSS.n270 2.6005
R234 VSS.n273 VSS.n272 2.6005
R235 VSS.n276 VSS.n275 2.6005
R236 VSS.n278 VSS.n277 2.6005
R237 VSS.n282 VSS.n281 2.6005
R238 VSS.n289 VSS.n288 2.6005
R239 VSS.n288 VSS.n287 2.6005
R240 VSS.n286 VSS.n285 2.6005
R241 VSS.n285 VSS.n284 2.6005
R242 VSS.n102 VSS.n101 2.6005
R243 VSS.n101 VSS.n100 2.6005
R244 VSS.n105 VSS.n104 2.6005
R245 VSS.n104 VSS.n103 2.6005
R246 VSS.n124 VSS.n123 2.6005
R247 VSS.n125 VSS.n124 2.6005
R248 VSS.n122 VSS.n121 2.6005
R249 VSS.n121 VSS.n120 2.6005
R250 VSS.n119 VSS.n118 2.6005
R251 VSS.n118 VSS.n117 2.6005
R252 VSS.n114 VSS.n113 2.6005
R253 VSS.n113 VSS.n112 2.6005
R254 VSS.n111 VSS.n110 2.6005
R255 VSS.n110 VSS.n109 2.6005
R256 VSS.n108 VSS.n107 2.6005
R257 VSS.n107 VSS.n106 2.6005
R258 VSS.n6 VSS.n5 2.6005
R259 VSS.n5 VSS.n4 2.6005
R260 VSS.n157 VSS.n156 2.6005
R261 VSS.n156 VSS.n155 2.6005
R262 VSS.n160 VSS.n159 2.6005
R263 VSS.n159 VSS.n158 2.6005
R264 VSS.n163 VSS.n162 2.6005
R265 VSS.n162 VSS.n161 2.6005
R266 VSS.n166 VSS.n165 2.6005
R267 VSS.n165 VSS.n164 2.6005
R268 VSS.n172 VSS.n171 2.6005
R269 VSS.n171 VSS.n170 2.6005
R270 VSS.n175 VSS.n174 2.6005
R271 VSS.n174 VSS.n173 2.6005
R272 VSS.n178 VSS.n177 2.6005
R273 VSS.n177 VSS.n176 2.6005
R274 VSS.n182 VSS.n181 2.6005
R275 VSS.n181 VSS.n180 2.6005
R276 VSS.n185 VSS.n184 2.6005
R277 VSS.n184 VSS.n183 2.6005
R278 VSS.n188 VSS.n187 2.6005
R279 VSS.n187 VSS.n186 2.6005
R280 VSS.n191 VSS.n190 2.6005
R281 VSS.n190 VSS.n189 2.6005
R282 VSS.n199 VSS.n198 2.6005
R283 VSS.n198 VSS.n197 2.6005
R284 VSS.n202 VSS.n201 2.6005
R285 VSS.n201 VSS.n200 2.6005
R286 VSS.n205 VSS.n204 2.6005
R287 VSS.n204 VSS.n203 2.6005
R288 VSS.n292 VSS.n291 2.6005
R289 VSS.n291 VSS.n290 2.6005
R290 VSS.n99 VSS.n98 2.6005
R291 VSS.n98 VSS.n97 2.6005
R292 VSS.n144 VSS.n143 2.6005
R293 VSS.n143 VSS.n142 2.6005
R294 VSS.n147 VSS.n146 2.6005
R295 VSS.n146 VSS.n145 2.6005
R296 VSS.n150 VSS.n149 2.6005
R297 VSS.n149 VSS.n148 2.6005
R298 VSS.n153 VSS.n152 2.6005
R299 VSS.n152 VSS.n151 2.6005
R300 VSS VSS.n329 2.6005
R301 VSS.n329 VSS.n328 2.6005
R302 VSS.n327 VSS.n326 2.6005
R303 VSS.n326 VSS.n325 2.6005
R304 VSS.n323 VSS.n322 2.6005
R305 VSS.n322 VSS.n321 2.6005
R306 VSS.n320 VSS.n319 2.6005
R307 VSS.n319 VSS.n318 2.6005
R308 VSS.n317 VSS.n316 2.6005
R309 VSS.n316 VSS.n315 2.6005
R310 VSS.n313 VSS.n312 2.6005
R311 VSS.n312 VSS.n311 2.6005
R312 VSS.n140 VSS.n139 2.6005
R313 VSS.n139 VSS.n138 2.6005
R314 VSS.n180 VSS.n179 2.57374
R315 VSS.n84 VSS.n83 2.48961
R316 VSS.n87 VSS.n86 2.48961
R317 VSS.n90 VSS.n89 2.48961
R318 VSS.n297 VSS.n296 2.24725
R319 VSS.n295 VSS.n196 2.24654
R320 VSS.n9 VSS.t2 2.02837
R321 VSS.n195 VSS.n194 2.00969
R322 VSS.n195 VSS.t6 1.82525
R323 VSS.n9 VSS.n8 1.80405
R324 VSS.n270 VSS.n269 1.68421
R325 VSS.n275 VSS.n274 1.68411
R326 VSS.n281 VSS.n280 1.68411
R327 VSS.n79 VSS.n78 1.43195
R328 VSS.n94 VSS.n93 1.43182
R329 VSS.n13 VSS.n11 1.02489
R330 VSS.n93 VSS.n92 0.780455
R331 VSS.n280 VSS.n279 0.459446
R332 VSS VSS.n310 0.243106
R333 VSS.n59 VSS.n56 0.188
R334 VSS.n137 VSS.n136 0.169688
R335 VSS.n136 VSS.n134 0.161214
R336 VSS.n310 VSS.n309 0.161214
R337 VSS.n286 VSS.n282 0.15275
R338 VSS.n131 VSS.n130 0.151571
R339 VSS.n307 VSS.n306 0.150768
R340 VSS.n140 VSS.n137 0.148402
R341 VSS.n294 VSS.n293 0.139082
R342 VSS.n99 VSS.n95 0.12841
R343 VSS.n248 VSS.n246 0.128
R344 VSS.n102 VSS.n99 0.113945
R345 VSS.n105 VSS.n102 0.113945
R346 VSS.n123 VSS.n105 0.113945
R347 VSS.n123 VSS.n122 0.113945
R348 VSS.n122 VSS.n119 0.113945
R349 VSS.n114 VSS.n111 0.113945
R350 VSS.n111 VSS.n108 0.113945
R351 VSS.n160 VSS.n157 0.113945
R352 VSS.n163 VSS.n160 0.113945
R353 VSS.n166 VSS.n163 0.113945
R354 VSS.n175 VSS.n172 0.113945
R355 VSS.n178 VSS.n175 0.113945
R356 VSS.n182 VSS.n178 0.113945
R357 VSS.n185 VSS.n182 0.113945
R358 VSS.n188 VSS.n185 0.113945
R359 VSS.n191 VSS.n188 0.113945
R360 VSS.n202 VSS.n199 0.113945
R361 VSS.n205 VSS.n202 0.113945
R362 VSS.n292 VSS.n289 0.113933
R363 VSS.n289 VSS.n286 0.113
R364 VSS.n251 VSS.n248 0.113
R365 VSS.n254 VSS.n251 0.113
R366 VSS.n257 VSS.n254 0.113
R367 VSS.n260 VSS.n257 0.113
R368 VSS.n263 VSS.n260 0.113
R369 VSS.n266 VSS.n263 0.113
R370 VSS.n268 VSS.n266 0.113
R371 VSS.n271 VSS.n268 0.113
R372 VSS.n273 VSS.n271 0.113
R373 VSS.n276 VSS.n273 0.113
R374 VSS.n278 VSS.n276 0.113
R375 VSS.n282 VSS.n278 0.113
R376 VSS.n62 VSS.n59 0.113
R377 VSS.n65 VSS.n62 0.113
R378 VSS.n68 VSS.n65 0.113
R379 VSS.n71 VSS.n68 0.113
R380 VSS.n74 VSS.n71 0.113
R381 VSS.n77 VSS.n74 0.113
R382 VSS.n80 VSS.n77 0.113
R383 VSS.n82 VSS.n80 0.113
R384 VSS.n85 VSS.n82 0.113
R385 VSS.n88 VSS.n85 0.113
R386 VSS.n91 VSS.n88 0.113
R387 VSS.n95 VSS.n91 0.113
R388 VSS.n56 VSS.n53 0.113
R389 VSS.n53 VSS.n50 0.113
R390 VSS.n50 VSS.n47 0.113
R391 VSS.n47 VSS.n44 0.113
R392 VSS.n44 VSS.n41 0.113
R393 VSS.n41 VSS.n38 0.113
R394 VSS.n38 VSS.n35 0.113
R395 VSS.n35 VSS.n32 0.113
R396 VSS.n32 VSS.n29 0.113
R397 VSS.n29 VSS.n25 0.113
R398 VSS.n25 VSS.n22 0.113
R399 VSS.n22 VSS.n19 0.113
R400 VSS.n19 VSS.n16 0.113
R401 VSS.n211 VSS.n208 0.113
R402 VSS.n214 VSS.n211 0.113
R403 VSS.n218 VSS.n214 0.113
R404 VSS.n221 VSS.n218 0.113
R405 VSS.n224 VSS.n221 0.113
R406 VSS.n227 VSS.n224 0.113
R407 VSS.n230 VSS.n227 0.113
R408 VSS.n233 VSS.n230 0.113
R409 VSS.n236 VSS.n233 0.113
R410 VSS.n239 VSS.n236 0.113
R411 VSS.n242 VSS.n239 0.113
R412 VSS.n246 VSS.n242 0.113
R413 VSS.n167 VSS.n166 0.107895
R414 VSS.n134 VSS.n132 0.0808571
R415 VSS.n309 VSS.n308 0.0808571
R416 VSS.n137 VSS.n7 0.07925
R417 VSS.n313 VSS 0.07925
R418 VSS.n132 VSS 0.0760357
R419 VSS.n324 VSS.n167 0.0755
R420 VSS.n108 VSS.n7 0.0753739
R421 VSS.n308 VSS 0.0752321
R422 VSS.n293 VSS.n205 0.0715924
R423 VSS.n199 VSS.n192 0.0678109
R424 VSS.n115 VSS.n114 0.0640294
R425 VSS.n308 VSS.n192 0.0639286
R426 VSS.n147 VSS.n144 0.0596608
R427 VSS.n150 VSS.n147 0.0596608
R428 VSS.n153 VSS.n150 0.0596608
R429 VSS VSS.n327 0.0596608
R430 VSS.n323 VSS.n320 0.0596608
R431 VSS.n320 VSS.n317 0.0596608
R432 VSS.n154 VSS.n153 0.0552552
R433 VSS.n119 VSS.n115 0.050416
R434 VSS.n192 VSS.n191 0.0466345
R435 VSS.n314 VSS.n313 0.0439266
R436 VSS.n293 VSS.n292 0.0428529
R437 VSS.n7 VSS.n6 0.0390714
R438 VSS.n327 VSS.n324 0.0376329
R439 VSS.n245 VSS.n244 0.0373597
R440 VSS.n141 VSS.n140 0.0351154
R441 VSS.n129 VSS.n128 0.028625
R442 VSS.n303 VSS.n300 0.028625
R443 VSS.n144 VSS.n141 0.0250455
R444 VSS.n324 VSS.n323 0.022528
R445 VSS.n297 VSS.n295 0.0174458
R446 VSS.n300 VSS.n297 0.0173807
R447 VSS.n317 VSS.n314 0.0162343
R448 VSS.n306 VSS.n303 0.0109464
R449 VSS.n130 VSS.n129 0.0101429
R450 VSS.n295 VSS.n294 0.0101429
R451 VSS.n172 VSS.n167 0.00655042
R452 VSS VSS.n307 0.006125
R453 VSS VSS.n131 0.00532143
R454 VSS VSS.n154 0.00490559
R455 Tr_Gate_1.CLK.n3 Tr_Gate_1.CLK.t15 45.6363
R456 Tr_Gate_1.CLK.n5 Tr_Gate_1.CLK.t20 29.6446
R457 Tr_Gate_1.CLK.t18 Tr_Gate_1.CLK.n6 29.6446
R458 Tr_Gate_1.CLK.n7 Tr_Gate_1.CLK.t21 24.6117
R459 Tr_Gate_1.CLK.n6 Tr_Gate_1.CLK.n5 22.2047
R460 Tr_Gate_1.CLK.t15 Tr_Gate_1.CLK.t19 22.1925
R461 Tr_Gate_1.CLK.n4 Tr_Gate_1.CLK.n3 20.9314
R462 Tr_Gate_1.CLK Tr_Gate_1.CLK.t18 18.5231
R463 Tr_Gate_1.CLK.n7 Tr_Gate_1.CLK.t17 6.1325
R464 Tr_Gate_1.CLK.n5 Tr_Gate_1.CLK.t14 6.1325
R465 Tr_Gate_1.CLK.n6 Tr_Gate_1.CLK.t12 6.1325
R466 Tr_Gate_1.CLK.n3 Tr_Gate_1.CLK.t16 6.1325
R467 Tr_Gate_1.CLK.n4 Tr_Gate_1.CLK.t13 6.1325
R468 Tr_Gate_1.CLK.n2 Tr_Gate_1.CLK.n4 5.28481
R469 Tr_Gate_1.CLK.n2 Tr_Gate_1.CLK.n7 4.89628
R470 Tr_Gate_1.CLK.n17 Tr_Gate_1.CLK.t8 3.6405
R471 Tr_Gate_1.CLK.n17 Tr_Gate_1.CLK.n16 3.6405
R472 Tr_Gate_1.CLK.n13 Tr_Gate_1.CLK.t9 3.6405
R473 Tr_Gate_1.CLK.n13 Tr_Gate_1.CLK.n12 3.6405
R474 Tr_Gate_1.CLK.n11 Tr_Gate_1.CLK.t7 3.6405
R475 Tr_Gate_1.CLK.n11 Tr_Gate_1.CLK.n10 3.6405
R476 Tr_Gate_1.CLK.n19 Tr_Gate_1.CLK.t10 3.6405
R477 Tr_Gate_1.CLK.n19 Tr_Gate_1.CLK.n18 3.6405
R478 Tr_Gate_1.CLK.n1 Tr_Gate_1.CLK.n9 3.50463
R479 Tr_Gate_1.CLK.n0 Tr_Gate_1.CLK.n15 3.50463
R480 Tr_Gate_1.CLK.n9 Tr_Gate_1.CLK.t6 3.2765
R481 Tr_Gate_1.CLK.n9 Tr_Gate_1.CLK.n8 3.2765
R482 Tr_Gate_1.CLK.n15 Tr_Gate_1.CLK.t5 3.2765
R483 Tr_Gate_1.CLK.n15 Tr_Gate_1.CLK.n14 3.2765
R484 Tr_Gate_1.CLK.n0 Tr_Gate_1.CLK.n11 3.06224
R485 Tr_Gate_1.CLK.n1 Tr_Gate_1.CLK.n17 3.06224
R486 Tr_Gate_1.CLK.n0 Tr_Gate_1.CLK.n13 2.6005
R487 Tr_Gate_1.CLK.n1 Tr_Gate_1.CLK.n19 2.6005
R488 Tr_Gate_1.CLK.n1 Tr_Gate_1.CLK.n0 0.98463
R489 Tr_Gate_1.CLK Tr_Gate_1.CLK.n1 0.747891
R490 Tr_Gate_1.CLK.n2 Tr_Gate_1.CLK 0.629606
R491 Tr_Gate_1.CLK Tr_Gate_1.CLK.n2 0.253378
R492 VDD.n40 VDD.t28 122.1
R493 VDD.t9 VDD.n15 121.091
R494 VDD.t2 VDD.n38 116.044
R495 VDD.n39 VDD.t2 105.954
R496 VDD.n16 VDD.t1 104.945
R497 VDD.n16 VDD.t9 100.909
R498 VDD.t28 VDD.n39 99.8996
R499 VDD.n38 VDD.t3 89.8088
R500 VDD.n18 VDD.t7 88.7997
R501 VDD.n15 VDD.t4 84.7634
R502 VDD.n40 VDD.t0 83.7543
R503 VDD.n55 VDD.t22 39.6722
R504 VDD.n58 VDD.n36 23.2342
R505 VDD.n63 VDD.t16 21.8883
R506 VDD.n58 VDD.n37 20.3898
R507 VDD.n5 VDD.t19 13.6804
R508 VDD.n2 VDD.n1 6.70224
R509 VDD.n37 VDD.t35 6.65503
R510 VDD.n48 VDD.n38 6.3005
R511 VDD VDD.n39 6.3005
R512 VDD.n47 VDD.n40 6.3005
R513 VDD.n15 VDD.n14 6.3005
R514 VDD.n17 VDD.n16 6.3005
R515 VDD.n19 VDD.n18 6.3005
R516 VDD.n37 VDD.t23 6.2405
R517 VDD.n2 VDD.n0 6.2405
R518 VDD.n44 VDD.n43 5.77744
R519 VDD.n10 VDD.t8 5.77744
R520 VDD.n45 VDD.t24 5.07264
R521 VDD.n12 VDD.n11 5.07264
R522 VDD.n26 VDD.t13 4.10447
R523 VDD.n33 VDD.t14 3.6405
R524 VDD.n33 VDD.n32 3.6405
R525 VDD.n35 VDD.t27 3.6405
R526 VDD.n35 VDD.n34 3.6405
R527 VDD.n7 VDD.n6 3.1505
R528 VDD.n6 VDD.n5 3.1505
R529 VDD.n25 VDD.n24 3.1505
R530 VDD.n24 VDD.n23 3.1505
R531 VDD.n28 VDD.n27 3.1505
R532 VDD.n27 VDD.n26 3.1505
R533 VDD VDD.n67 3.1505
R534 VDD.n67 VDD.n66 3.1505
R535 VDD.n65 VDD.n64 3.1505
R536 VDD.n64 VDD.n63 3.1505
R537 VDD.n62 VDD.n61 3.1505
R538 VDD.n61 VDD.n60 3.1505
R539 VDD.n57 VDD.n56 3.1505
R540 VDD.n56 VDD.n55 3.1505
R541 VDD.n54 VDD.n53 3.1505
R542 VDD.n4 VDD.n3 3.1505
R543 VDD.n36 VDD.n35 3.06224
R544 VDD.n44 VDD.n42 2.87637
R545 VDD.n10 VDD.n9 2.87637
R546 VDD.n36 VDD.n33 2.6005
R547 VDD.n42 VDD.t15 2.16717
R548 VDD.n42 VDD.n41 2.16717
R549 VDD.n9 VDD.t10 2.16717
R550 VDD.n9 VDD.n8 2.16717
R551 VDD.n30 VDD.n29 0.662808
R552 VDD.n59 VDD.n31 0.662808
R553 VDD.n51 VDD.n50 0.662808
R554 VDD.n22 VDD.n21 0.662808
R555 VDD.n45 VDD.n44 0.6395
R556 VDD.n12 VDD.n10 0.6395
R557 VDD.n21 VDD.n20 0.597767
R558 VDD.n4 VDD.n2 0.389323
R559 VDD.n50 VDD.n49 0.388557
R560 VDD VDD.n30 0.215115
R561 VDD.n53 VDD.n52 0.182274
R562 VDD.n48 VDD 0.174184
R563 VDD VDD.n47 0.174184
R564 VDD.n19 VDD.n17 0.174184
R565 VDD.n14 VDD 0.173395
R566 VDD.n49 VDD.n48 0.158395
R567 VDD.n20 VDD.n19 0.158395
R568 VDD.n14 VDD.n13 0.1355
R569 VDD.n47 VDD.n46 0.134711
R570 VDD.n46 VDD.n45 0.0893158
R571 VDD.n13 VDD.n12 0.0893158
R572 VDD.n65 VDD.n62 0.0714756
R573 VDD.n57 VDD.n54 0.0714756
R574 VDD.n7 VDD.n4 0.0692805
R575 VDD.n28 VDD.n25 0.0692805
R576 VDD VDD.n65 0.0692805
R577 VDD.n31 VDD 0.0616538
R578 VDD.n29 VDD.n28 0.0561098
R579 VDD.n54 VDD.n51 0.055378
R580 VDD.n25 VDD.n22 0.0414756
R581 VDD.n59 VDD.n58 0.0326951
R582 VDD.n22 VDD.n7 0.0305
R583 VDD.n62 VDD.n59 0.0202561
R584 VDD.n58 VDD.n57 0.0173293
R585 VDD VDD.n29 0.0158659
R586 VDD.n17 VDD 0.00128947
R587 a_2663_557.n2 a_2663_557.t7 29.2961
R588 a_2663_557.n3 a_2663_557.n2 21.9292
R589 a_2663_557.n4 a_2663_557.n3 18.1271
R590 a_2663_557.n4 a_2663_557.t8 11.1695
R591 a_2663_557.n2 a_2663_557.t9 6.1325
R592 a_2663_557.n3 a_2663_557.t6 6.1325
R593 a_2663_557.n7 a_2663_557.n6 4.93252
R594 a_2663_557.n7 a_2663_557.t1 4.70348
R595 a_2663_557.n5 a_2663_557.n4 4.6311
R596 a_2663_557.n5 a_2663_557.n1 2.85093
R597 a_2663_557.n1 a_2663_557.t2 2.16717
R598 a_2663_557.n1 a_2663_557.n0 2.16717
R599 a_2663_557.t5 a_2663_557.n10 2.16717
R600 a_2663_557.n10 a_2663_557.n9 2.16717
R601 a_2663_557.n8 a_2663_557.n7 1.58583
R602 a_2663_557.n10 a_2663_557.n8 1.24398
R603 a_2663_557.n8 a_2663_557.n5 0.971047
R604 IN1.n6 IN1.t2 5.81586
R605 IN1.n3 IN1.n0 5.10148
R606 IN1.n10 IN1.n9 5.10115
R607 IN1.n8 IN1.n7 5.08021
R608 IN1.n3 IN1.n2 4.66166
R609 IN1.n6 IN1.n5 2.85093
R610 IN1.n5 IN1.t3 2.16717
R611 IN1.n5 IN1.n4 2.16717
R612 IN1.n2 IN1.t5 1.9505
R613 IN1.n2 IN1.n1 1.9505
R614 IN1.n8 IN1.n6 0.644196
R615 IN1.n10 IN1.n8 0.45084
R616 IN1.n11 IN1.n3 0.309585
R617 IN1.n11 IN1.n10 0.274999
R618 IN1 IN1.n11 0.0936034
R619 a_268_897.n5 a_268_897.t9 29.2961
R620 a_268_897.n6 a_268_897.n5 21.9292
R621 a_268_897.n7 a_268_897.n6 18.1271
R622 a_268_897.n7 a_268_897.t6 11.1695
R623 a_268_897.n3 a_268_897.t1 10.2143
R624 a_268_897.n5 a_268_897.t8 6.1325
R625 a_268_897.n6 a_268_897.t7 6.1325
R626 a_268_897.n3 a_268_897.n2 4.68517
R627 a_268_897.n8 a_268_897.n7 4.6311
R628 a_268_897.n10 a_268_897.n8 2.85093
R629 a_268_897.n1 a_268_897.t4 2.16717
R630 a_268_897.n1 a_268_897.n0 2.16717
R631 a_268_897.t5 a_268_897.n10 2.16717
R632 a_268_897.n10 a_268_897.n9 2.16717
R633 a_268_897.n4 a_268_897.n3 1.58582
R634 a_268_897.n4 a_268_897.n1 1.24371
R635 a_268_897.n8 a_268_897.n4 0.971051
C0 IN1 VDD 0.112f
C1 OUT IN2 1.25f
C2 SEL IN2 0.53f
C3 OUT Tr_Gate_1.CLK 0.425f
C4 Tr_Gate_1.CLK SEL 0.403f
C5 OUT VDD 1.01f
C6 VDD SEL 2.75f
C7 OUT IN1 1.25f
C8 IN1 SEL 8.5e-19
C9 VDD IN2 0.112f
C10 Tr_Gate_1.CLK VDD 1.84f
C11 IN1 Tr_Gate_1.CLK 0.49f
C12 OUT SEL 0.52f
.ends

