magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2195 -3545 2195 3545
<< ndiff >>
rect -195 1523 195 1545
rect -195 -1523 -173 1523
rect 173 -1523 195 1523
rect -195 -1545 195 -1523
<< ndiffc >>
rect -173 -1523 173 1523
<< metal1 >>
rect -184 1523 184 1534
rect -184 -1523 -173 1523
rect 173 -1523 184 1523
rect -184 -1534 184 -1523
<< end >>
