* NGSPICE file created from Output_Div_Mag.ext - technology: gf180mcuC

.subckt pmos_3p3_M8SWPS a_n28_n124# a_n116_n80# a_28_n80# w_n202_n210#
X0 a_28_n80# a_n28_n124# a_n116_n80# w_n202_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
.ends

.subckt nmos_3p3_5QNVWA a_n116_n44# a_28_n44# a_n28_n88# VSUBS
X0 a_28_n44# a_n28_n88# a_n116_n44# VSUBS nfet_03v3 ad=0.194p pd=1.76u as=0.194p ps=1.76u w=0.44u l=0.28u
.ends

.subckt nand2 VDD IN2 IN1 OUT VSS m1_186_70#
Xpmos_3p3_M8SWPS_0 IN1 OUT VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD OUT VDD pmos_3p3_M8SWPS
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# OUT IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt pmos_3p3_MQGBLR a_n28_n124# a_n116_n80# a_28_n80# w_n202_n210#
X0 a_28_n80# a_n28_n124# a_n116_n80# w_n202_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
.ends

.subckt nmos_3p3_DDNVWA a_n120_n36# a_28_n22# a_n28_n66# VSUBS
X0 a_28_n22# a_n28_n66# a_n120_n36# VSUBS nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
.ends

.subckt nverterlayout VDD VSS OUT IN
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt mux_2x1 Sel I0 I1 VDD OUT VSS
Xnand2_0 VDD I1 Sel nand2_1/IN2 VSS nand2_0/m1_186_70# nand2
Xnand2_1 VDD nand2_1/IN2 nand2_2/OUT OUT VSS nand2_1/m1_186_70# nand2
Xnand2_2 VDD nand2_2/IN2 I0 nand2_2/OUT VSS nand2_2/m1_186_70# nand2
Xnverterlayout_0 VDD VSS nand2_2/IN2 Sel nverterlayout
.ends

.subckt mux_4x1 I0 I1 I2 I3 S1 S0 OUT VDD VSS mux_2x1_1/I0
Xmux_2x1_0 S0 I2 I3 VDD mux_2x1_1/I1 VSS mux_2x1
Xmux_2x1_1 S1 mux_2x1_1/I0 mux_2x1_1/I1 VDD OUT VSS mux_2x1
Xmux_2x1_2 S0 I0 I1 VDD mux_2x1_1/I0 VSS mux_2x1
.ends

.subckt nand2_ibr VDD IN2 IN1 OUT VSS m1_186_70#
Xpmos_3p3_M8SWPS_0 IN1 OUT VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD OUT VDD pmos_3p3_M8SWPS
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# OUT IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt nverterlayout_ibr VDD VSS OUT IN
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt and_2_ibr VDD IN2 OUT IN1 nand2_ibr_0/OUT nand2_ibr_0/m1_186_70# VSS
Xnand2_ibr_0 VDD IN2 IN1 nand2_ibr_0/OUT VSS nand2_ibr_0/m1_186_70# nand2_ibr
Xnverterlayout_ibr_0 VDD VSS OUT nand2_ibr_0/OUT nverterlayout_ibr
.ends

.subckt dec_2x4_ibr_mag IN1 IN2 D0 D1 D2 D3 VSS VDD
Xand_2_ibr_0 VDD nand2_2/IN2 D0 nand2_1/IN1 nand2_0/OUT nand2_0/m1_186_70# VSS and_2_ibr
Xand_2_ibr_1 VDD IN1 D1 nand2_1/IN1 nand2_1/OUT nand2_1/m1_186_70# VSS and_2_ibr
Xand_2_ibr_3 VDD IN1 D3 IN2 nand2_3/OUT nand2_3/m1_186_70# VSS and_2_ibr
Xand_2_ibr_2 VDD nand2_2/IN2 D2 IN2 nand2_2/OUT nand2_2/m1_186_70# VSS and_2_ibr
Xnverterlayout_ibr_0 VDD VSS nand2_2/IN2 IN1 nverterlayout_ibr
Xnverterlayout_ibr_1 VDD VSS nand2_1/IN1 IN2 nverterlayout_ibr
Xnand2_0 VDD nand2_2/IN2 nand2_1/IN1 nand2_0/OUT VSS nand2_0/m1_186_70# nand2
Xnand2_2 VDD nand2_2/IN2 IN2 nand2_2/OUT VSS nand2_2/m1_186_70# nand2
Xnand2_1 VDD IN1 nand2_1/IN1 nand2_1/OUT VSS nand2_1/m1_186_70# nand2
Xnand2_3 VDD IN1 IN2 nand2_3/OUT VSS nand2_3/m1_186_70# nand2
.ends

.subckt nand2_mag IN2 OUT IN1 VDD VSS
Xpmos_3p3_M8SWPS_0 IN1 OUT VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD OUT VDD pmos_3p3_M8SWPS
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# OUT IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt nmos_3p3_VGTVWA a_n116_n66# a_28_n66# a_n28_n110# VSUBS
X0 a_28_n66# a_n28_n110# a_n116_n66# VSUBS nfet_03v3 ad=0.29p pd=2.2u as=0.29p ps=2.2u w=0.66u l=0.28u
.ends

.subckt nand3_mag IN3 IN2 IN1 VDD VSS OUT
Xnmos_3p3_VGTVWA_0 nmos_3p3_VGTVWA_1/a_28_n66# nmos_3p3_VGTVWA_0/a_28_n66# IN2 VSS
+ nmos_3p3_VGTVWA
Xnmos_3p3_VGTVWA_1 VSS nmos_3p3_VGTVWA_1/a_28_n66# IN3 VSS nmos_3p3_VGTVWA
Xnmos_3p3_VGTVWA_2 nmos_3p3_VGTVWA_0/a_28_n66# OUT IN1 VSS nmos_3p3_VGTVWA
Xpmos_3p3_M8SWPS_0 IN1 VDD OUT VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN3 VDD OUT VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_2 IN2 OUT VDD VDD pmos_3p3_M8SWPS
.ends

.subckt GF_INV_MAG VDD VSS IN OUT
Xpmos_3p3_MQGBLR_0 IN VDD OUT VDD pmos_3p3_MQGBLR
Xnmos_3p3_DDNVWA_0 VSS OUT IN VSS nmos_3p3_DDNVWA
.ends

.subckt JK_FF_mag CLK RST Q QB J K nand2_mag_4/IN2 nand3_mag_2/OUT nand3_mag_0/OUT
+ nand3_mag_1/OUT VDD VSS
Xnand2_mag_1 nand2_mag_1/IN2 Q QB VDD VSS nand2_mag
Xnand3_mag_2 J CLK Q VDD VSS nand3_mag_2/OUT nand3_mag
Xnand2_mag_2 nand3_mag_0/OUT nand3_mag_1/IN1 nand3_mag_1/OUT VDD VSS nand2_mag
Xnand2_mag_3 nand3_mag_1/OUT nand2_mag_4/IN2 nand2_mag_3/IN1 VDD VSS nand2_mag
Xnand2_mag_4 nand2_mag_4/IN2 QB Q VDD VSS nand2_mag
XGF_INV_MAG_0 VDD VSS CLK nand2_mag_3/IN1 GF_INV_MAG
Xnand3_mag_0 K CLK QB VDD VSS nand3_mag_0/OUT nand3_mag
Xnand2_mag_0 nand3_mag_1/IN1 nand2_mag_1/IN2 nand2_mag_3/IN1 VDD VSS nand2_mag
Xnand3_mag_1 nand3_mag_2/OUT RST nand3_mag_1/IN1 VDD VSS nand3_mag_1/OUT nand3_mag
.ends

.subckt CLK_div_2_mag Vdiv2 CLK JK_FF_mag_0/nand3_mag_0/OUT JK_FF_mag_0/nand3_mag_1/OUT
+ RST VSS JK_FF_mag_0/nand3_mag_2/OUT VDD
XJK_FF_mag_0 CLK RST Vdiv2 JK_FF_mag_0/QB VDD VDD JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_2/OUT
+ JK_FF_mag_0/nand3_mag_0/OUT JK_FF_mag_0/nand3_mag_1/OUT VDD VSS JK_FF_mag
.ends

.subckt CLK_div_4_mag Vdiv4 RST CLK CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_1/OUT
+ CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_2/OUT CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT
+ VDD CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_0/OUT
+ VSS
XCLK_div_2_mag_0 CLK_div_2_mag_1/CLK CLK CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT
+ CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT RST VSS CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT
+ VDD CLK_div_2_mag
XCLK_div_2_mag_1 Vdiv4 CLK_div_2_mag_1/CLK CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_0/OUT
+ CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_1/OUT RST VSS CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_2/OUT
+ VDD CLK_div_2_mag
.ends

.subckt pmos_3p3_M8QNDR w_n202_n290# a_28_n160# a_n116_n160# a_n28_n204#
X0 a_28_n160# a_n28_n204# a_n116_n160# w_n202_n290# pfet_03v3 ad=0.704p pd=4.08u as=0.704p ps=4.08u w=1.6u l=0.28u
.ends

.subckt pmos_3p3_M4YALR w_n202_n290# a_28_n160# a_n116_n160# a_n28_n204#
X0 a_28_n160# a_n28_n204# a_n116_n160# w_n202_n290# pfet_03v3 ad=0.704p pd=4.08u as=0.704p ps=4.08u w=1.6u l=0.28u
.ends

.subckt or_2_mag VSS VDD IN2 IN1 OUT
Xpmos_3p3_M8QNDR_0 VDD pmos_3p3_M8QNDR_0/a_28_n160# VDD IN2 pmos_3p3_M8QNDR
XGF_INV_MAG_1 VDD VSS GF_INV_MAG_1/IN OUT GF_INV_MAG
Xpmos_3p3_M4YALR_0 VDD GF_INV_MAG_1/IN pmos_3p3_M8QNDR_0/a_28_n160# IN1 pmos_3p3_M4YALR
Xnmos_3p3_DDNVWA_0 GF_INV_MAG_1/IN VSS IN1 VSS nmos_3p3_DDNVWA
Xnmos_3p3_DDNVWA_1 VSS GF_INV_MAG_1/IN IN2 VSS nmos_3p3_DDNVWA
.ends

.subckt and2_mag IN2 IN1 OUT VSS VDD
Xpmos_3p3_M8SWPS_0 IN1 GF_INV_MAG_0/IN VDD VDD pmos_3p3_M8SWPS
Xpmos_3p3_M8SWPS_1 IN2 VDD GF_INV_MAG_0/IN VDD pmos_3p3_M8SWPS
XGF_INV_MAG_0 VDD VSS GF_INV_MAG_0/IN OUT GF_INV_MAG
Xnmos_3p3_5QNVWA_0 VSS m1_186_70# IN2 VSS nmos_3p3_5QNVWA
Xnmos_3p3_5QNVWA_1 m1_186_70# GF_INV_MAG_0/IN IN1 VSS nmos_3p3_5QNVWA
.ends

.subckt CLK_div_3_mag Q1 Q0 Vdiv3 CLK RST JK_FF_mag_1/nand3_mag_0/OUT JK_FF_mag_0/nand3_mag_0/OUT
+ JK_FF_mag_1/nand3_mag_1/OUT JK_FF_mag_0/nand3_mag_1/OUT JK_FF_mag_1/nand3_mag_2/OUT
+ VDD VSS JK_FF_mag_0/nand3_mag_2/OUT
XJK_FF_mag_0 CLK RST Q0 JK_FF_mag_1/K VDD Q1 JK_FF_mag_0/nand2_mag_4/IN2 JK_FF_mag_0/nand3_mag_2/OUT
+ JK_FF_mag_0/nand3_mag_0/OUT JK_FF_mag_0/nand3_mag_1/OUT VDD VSS JK_FF_mag
XJK_FF_mag_1 CLK RST Q1 JK_FF_mag_1/QB VDD JK_FF_mag_1/K JK_FF_mag_1/nand2_mag_4/IN2
+ JK_FF_mag_1/nand3_mag_2/OUT JK_FF_mag_1/nand3_mag_0/OUT JK_FF_mag_1/nand3_mag_1/OUT
+ VDD VSS JK_FF_mag
Xor_2_mag_0 VSS VDD or_2_mag_0/IN2 Q0 Vdiv3 or_2_mag
Xand2_mag_0 CLK Q1 or_2_mag_0/IN2 VSS VDD and2_mag
.ends

.subckt pmos_3p3_MW53B7 a_n188_n80# a_n100_n124# a_100_n80# w_n274_n210#
X0 a_100_n80# a_n100_n124# a_n188_n80# w_n274_n210# pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
.ends

.subckt nmos_3p3_MGBSF7 a_100_n22# a_n100_n66# a_n192_n36# VSUBS
X0 a_100_n22# a_n100_n66# a_n192_n36# VSUBS nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
.ends

.subckt Inverter_delayed_mag VDD VSS IN OUT
Xpmos_3p3_MW53B7_0 VDD IN OUT VDD pmos_3p3_MW53B7
Xnmos_3p3_MGBSF7_0 OUT IN VSS VSS nmos_3p3_MGBSF7
.ends

.subckt Buffer_delayed_mag IN OUT VDD VSS
Xpmos_3p3_MW53B7_0 VDD IN Inverter_delayed_mag_0/IN VDD pmos_3p3_MW53B7
XInverter_delayed_mag_0 VDD VSS Inverter_delayed_mag_0/IN OUT Inverter_delayed_mag
Xnmos_3p3_MGBSF7_0 Inverter_delayed_mag_0/IN IN VSS VSS nmos_3p3_MGBSF7
.ends

.subckt Output_Div_Mag OPA0 OPA1 Vdiv VDD VSS CLK RST
Xmux_4x1_0 mux_4x1_0/I0 mux_4x1_0/I1 mux_4x1_0/I2 mux_4x1_0/I3 OPA1 OPA0 Vdiv VDD
+ VSS mux_4x1_0/mux_2x1_1/I0 mux_4x1
Xdec_2x4_ibr_mag_0 OPA0 OPA1 dec_2x4_ibr_mag_0/D0 CLK_div_2_mag_0/VDD CLK_div_3_mag_0/VDD
+ CLK_div_4_mag_0/VDD VSS VDD dec_2x4_ibr_mag
XCLK_div_4_mag_0 mux_4x1_0/I3 RST CLK CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT
+ CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_2/OUT
+ CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_4_mag_0/VDD
+ CLK_div_4_mag_0/CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_4_mag_0/CLK_div_2_mag_1/JK_FF_mag_0/nand3_mag_0/OUT
+ VSS CLK_div_4_mag
XCLK_div_3_mag_0 CLK_div_3_mag_0/Q1 CLK_div_3_mag_0/Q0 mux_4x1_0/I2 CLK RST CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_0/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_1/OUT
+ CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_1/OUT CLK_div_3_mag_0/JK_FF_mag_1/nand3_mag_2/OUT
+ CLK_div_3_mag_0/VDD VSS CLK_div_3_mag_0/JK_FF_mag_0/nand3_mag_2/OUT CLK_div_3_mag
XCLK_div_2_mag_0 mux_4x1_0/I1 CLK CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_0/OUT CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_1/OUT
+ RST VSS CLK_div_2_mag_0/JK_FF_mag_0/nand3_mag_2/OUT CLK_div_2_mag_0/VDD CLK_div_2_mag
XBuffer_delayed_mag_0 CLK mux_4x1_0/I0 dec_2x4_ibr_mag_0/D0 VSS Buffer_delayed_mag
.ends

