magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1235 -1046 1235 1046
<< metal1 >>
rect -235 40 235 46
rect -235 14 -229 40
rect -203 14 -175 40
rect -149 14 -121 40
rect -95 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 95 40
rect 121 14 149 40
rect 175 14 203 40
rect 229 14 235 40
rect -235 -14 235 14
rect -235 -40 -229 -14
rect -203 -40 -175 -14
rect -149 -40 -121 -14
rect -95 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 95 -14
rect 121 -40 149 -14
rect 175 -40 203 -14
rect 229 -40 235 -14
rect -235 -46 235 -40
<< via1 >>
rect -229 14 -203 40
rect -175 14 -149 40
rect -121 14 -95 40
rect -67 14 -41 40
rect -13 14 13 40
rect 41 14 67 40
rect 95 14 121 40
rect 149 14 175 40
rect 203 14 229 40
rect -229 -40 -203 -14
rect -175 -40 -149 -14
rect -121 -40 -95 -14
rect -67 -40 -41 -14
rect -13 -40 13 -14
rect 41 -40 67 -14
rect 95 -40 121 -14
rect 149 -40 175 -14
rect 203 -40 229 -14
<< metal2 >>
rect -235 40 235 46
rect -235 14 -229 40
rect -203 14 -175 40
rect -149 14 -121 40
rect -95 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 95 40
rect 121 14 149 40
rect 175 14 203 40
rect 229 14 235 40
rect -235 -14 235 14
rect -235 -40 -229 -14
rect -203 -40 -175 -14
rect -149 -40 -121 -14
rect -95 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 95 -14
rect 121 -40 149 -14
rect 175 -40 203 -14
rect 229 -40 235 -14
rect -235 -46 235 -40
<< end >>
