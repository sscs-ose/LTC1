magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -4959 2045 4959
<< psubdiff >>
rect -45 2937 45 2959
rect -45 2891 -23 2937
rect 23 2891 45 2937
rect -45 2813 45 2891
rect -45 2767 -23 2813
rect 23 2767 45 2813
rect -45 2689 45 2767
rect -45 2643 -23 2689
rect 23 2643 45 2689
rect -45 2565 45 2643
rect -45 2519 -23 2565
rect 23 2519 45 2565
rect -45 2441 45 2519
rect -45 2395 -23 2441
rect 23 2395 45 2441
rect -45 2317 45 2395
rect -45 2271 -23 2317
rect 23 2271 45 2317
rect -45 2193 45 2271
rect -45 2147 -23 2193
rect 23 2147 45 2193
rect -45 2069 45 2147
rect -45 2023 -23 2069
rect 23 2023 45 2069
rect -45 1945 45 2023
rect -45 1899 -23 1945
rect 23 1899 45 1945
rect -45 1821 45 1899
rect -45 1775 -23 1821
rect 23 1775 45 1821
rect -45 1697 45 1775
rect -45 1651 -23 1697
rect 23 1651 45 1697
rect -45 1573 45 1651
rect -45 1527 -23 1573
rect 23 1527 45 1573
rect -45 1449 45 1527
rect -45 1403 -23 1449
rect 23 1403 45 1449
rect -45 1325 45 1403
rect -45 1279 -23 1325
rect 23 1279 45 1325
rect -45 1201 45 1279
rect -45 1155 -23 1201
rect 23 1155 45 1201
rect -45 1077 45 1155
rect -45 1031 -23 1077
rect 23 1031 45 1077
rect -45 953 45 1031
rect -45 907 -23 953
rect 23 907 45 953
rect -45 829 45 907
rect -45 783 -23 829
rect 23 783 45 829
rect -45 705 45 783
rect -45 659 -23 705
rect 23 659 45 705
rect -45 581 45 659
rect -45 535 -23 581
rect 23 535 45 581
rect -45 457 45 535
rect -45 411 -23 457
rect 23 411 45 457
rect -45 333 45 411
rect -45 287 -23 333
rect 23 287 45 333
rect -45 209 45 287
rect -45 163 -23 209
rect 23 163 45 209
rect -45 85 45 163
rect -45 39 -23 85
rect 23 39 45 85
rect -45 -39 45 39
rect -45 -85 -23 -39
rect 23 -85 45 -39
rect -45 -163 45 -85
rect -45 -209 -23 -163
rect 23 -209 45 -163
rect -45 -287 45 -209
rect -45 -333 -23 -287
rect 23 -333 45 -287
rect -45 -411 45 -333
rect -45 -457 -23 -411
rect 23 -457 45 -411
rect -45 -535 45 -457
rect -45 -581 -23 -535
rect 23 -581 45 -535
rect -45 -659 45 -581
rect -45 -705 -23 -659
rect 23 -705 45 -659
rect -45 -783 45 -705
rect -45 -829 -23 -783
rect 23 -829 45 -783
rect -45 -907 45 -829
rect -45 -953 -23 -907
rect 23 -953 45 -907
rect -45 -1031 45 -953
rect -45 -1077 -23 -1031
rect 23 -1077 45 -1031
rect -45 -1155 45 -1077
rect -45 -1201 -23 -1155
rect 23 -1201 45 -1155
rect -45 -1279 45 -1201
rect -45 -1325 -23 -1279
rect 23 -1325 45 -1279
rect -45 -1403 45 -1325
rect -45 -1449 -23 -1403
rect 23 -1449 45 -1403
rect -45 -1527 45 -1449
rect -45 -1573 -23 -1527
rect 23 -1573 45 -1527
rect -45 -1651 45 -1573
rect -45 -1697 -23 -1651
rect 23 -1697 45 -1651
rect -45 -1775 45 -1697
rect -45 -1821 -23 -1775
rect 23 -1821 45 -1775
rect -45 -1899 45 -1821
rect -45 -1945 -23 -1899
rect 23 -1945 45 -1899
rect -45 -2023 45 -1945
rect -45 -2069 -23 -2023
rect 23 -2069 45 -2023
rect -45 -2147 45 -2069
rect -45 -2193 -23 -2147
rect 23 -2193 45 -2147
rect -45 -2271 45 -2193
rect -45 -2317 -23 -2271
rect 23 -2317 45 -2271
rect -45 -2395 45 -2317
rect -45 -2441 -23 -2395
rect 23 -2441 45 -2395
rect -45 -2519 45 -2441
rect -45 -2565 -23 -2519
rect 23 -2565 45 -2519
rect -45 -2643 45 -2565
rect -45 -2689 -23 -2643
rect 23 -2689 45 -2643
rect -45 -2767 45 -2689
rect -45 -2813 -23 -2767
rect 23 -2813 45 -2767
rect -45 -2891 45 -2813
rect -45 -2937 -23 -2891
rect 23 -2937 45 -2891
rect -45 -2959 45 -2937
<< psubdiffcont >>
rect -23 2891 23 2937
rect -23 2767 23 2813
rect -23 2643 23 2689
rect -23 2519 23 2565
rect -23 2395 23 2441
rect -23 2271 23 2317
rect -23 2147 23 2193
rect -23 2023 23 2069
rect -23 1899 23 1945
rect -23 1775 23 1821
rect -23 1651 23 1697
rect -23 1527 23 1573
rect -23 1403 23 1449
rect -23 1279 23 1325
rect -23 1155 23 1201
rect -23 1031 23 1077
rect -23 907 23 953
rect -23 783 23 829
rect -23 659 23 705
rect -23 535 23 581
rect -23 411 23 457
rect -23 287 23 333
rect -23 163 23 209
rect -23 39 23 85
rect -23 -85 23 -39
rect -23 -209 23 -163
rect -23 -333 23 -287
rect -23 -457 23 -411
rect -23 -581 23 -535
rect -23 -705 23 -659
rect -23 -829 23 -783
rect -23 -953 23 -907
rect -23 -1077 23 -1031
rect -23 -1201 23 -1155
rect -23 -1325 23 -1279
rect -23 -1449 23 -1403
rect -23 -1573 23 -1527
rect -23 -1697 23 -1651
rect -23 -1821 23 -1775
rect -23 -1945 23 -1899
rect -23 -2069 23 -2023
rect -23 -2193 23 -2147
rect -23 -2317 23 -2271
rect -23 -2441 23 -2395
rect -23 -2565 23 -2519
rect -23 -2689 23 -2643
rect -23 -2813 23 -2767
rect -23 -2937 23 -2891
<< metal1 >>
rect -34 2937 34 2948
rect -34 2891 -23 2937
rect 23 2891 34 2937
rect -34 2813 34 2891
rect -34 2767 -23 2813
rect 23 2767 34 2813
rect -34 2689 34 2767
rect -34 2643 -23 2689
rect 23 2643 34 2689
rect -34 2565 34 2643
rect -34 2519 -23 2565
rect 23 2519 34 2565
rect -34 2441 34 2519
rect -34 2395 -23 2441
rect 23 2395 34 2441
rect -34 2317 34 2395
rect -34 2271 -23 2317
rect 23 2271 34 2317
rect -34 2193 34 2271
rect -34 2147 -23 2193
rect 23 2147 34 2193
rect -34 2069 34 2147
rect -34 2023 -23 2069
rect 23 2023 34 2069
rect -34 1945 34 2023
rect -34 1899 -23 1945
rect 23 1899 34 1945
rect -34 1821 34 1899
rect -34 1775 -23 1821
rect 23 1775 34 1821
rect -34 1697 34 1775
rect -34 1651 -23 1697
rect 23 1651 34 1697
rect -34 1573 34 1651
rect -34 1527 -23 1573
rect 23 1527 34 1573
rect -34 1449 34 1527
rect -34 1403 -23 1449
rect 23 1403 34 1449
rect -34 1325 34 1403
rect -34 1279 -23 1325
rect 23 1279 34 1325
rect -34 1201 34 1279
rect -34 1155 -23 1201
rect 23 1155 34 1201
rect -34 1077 34 1155
rect -34 1031 -23 1077
rect 23 1031 34 1077
rect -34 953 34 1031
rect -34 907 -23 953
rect 23 907 34 953
rect -34 829 34 907
rect -34 783 -23 829
rect 23 783 34 829
rect -34 705 34 783
rect -34 659 -23 705
rect 23 659 34 705
rect -34 581 34 659
rect -34 535 -23 581
rect 23 535 34 581
rect -34 457 34 535
rect -34 411 -23 457
rect 23 411 34 457
rect -34 333 34 411
rect -34 287 -23 333
rect 23 287 34 333
rect -34 209 34 287
rect -34 163 -23 209
rect 23 163 34 209
rect -34 85 34 163
rect -34 39 -23 85
rect 23 39 34 85
rect -34 -39 34 39
rect -34 -85 -23 -39
rect 23 -85 34 -39
rect -34 -163 34 -85
rect -34 -209 -23 -163
rect 23 -209 34 -163
rect -34 -287 34 -209
rect -34 -333 -23 -287
rect 23 -333 34 -287
rect -34 -411 34 -333
rect -34 -457 -23 -411
rect 23 -457 34 -411
rect -34 -535 34 -457
rect -34 -581 -23 -535
rect 23 -581 34 -535
rect -34 -659 34 -581
rect -34 -705 -23 -659
rect 23 -705 34 -659
rect -34 -783 34 -705
rect -34 -829 -23 -783
rect 23 -829 34 -783
rect -34 -907 34 -829
rect -34 -953 -23 -907
rect 23 -953 34 -907
rect -34 -1031 34 -953
rect -34 -1077 -23 -1031
rect 23 -1077 34 -1031
rect -34 -1155 34 -1077
rect -34 -1201 -23 -1155
rect 23 -1201 34 -1155
rect -34 -1279 34 -1201
rect -34 -1325 -23 -1279
rect 23 -1325 34 -1279
rect -34 -1403 34 -1325
rect -34 -1449 -23 -1403
rect 23 -1449 34 -1403
rect -34 -1527 34 -1449
rect -34 -1573 -23 -1527
rect 23 -1573 34 -1527
rect -34 -1651 34 -1573
rect -34 -1697 -23 -1651
rect 23 -1697 34 -1651
rect -34 -1775 34 -1697
rect -34 -1821 -23 -1775
rect 23 -1821 34 -1775
rect -34 -1899 34 -1821
rect -34 -1945 -23 -1899
rect 23 -1945 34 -1899
rect -34 -2023 34 -1945
rect -34 -2069 -23 -2023
rect 23 -2069 34 -2023
rect -34 -2147 34 -2069
rect -34 -2193 -23 -2147
rect 23 -2193 34 -2147
rect -34 -2271 34 -2193
rect -34 -2317 -23 -2271
rect 23 -2317 34 -2271
rect -34 -2395 34 -2317
rect -34 -2441 -23 -2395
rect 23 -2441 34 -2395
rect -34 -2519 34 -2441
rect -34 -2565 -23 -2519
rect 23 -2565 34 -2519
rect -34 -2643 34 -2565
rect -34 -2689 -23 -2643
rect 23 -2689 34 -2643
rect -34 -2767 34 -2689
rect -34 -2813 -23 -2767
rect 23 -2813 34 -2767
rect -34 -2891 34 -2813
rect -34 -2937 -23 -2891
rect 23 -2937 34 -2891
rect -34 -2948 34 -2937
<< end >>
