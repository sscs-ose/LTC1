magic
tech gf180mcuC
magscale 1 10
timestamp 1694088395
<< nwell >>
rect -864 -1121 864 1121
<< nsubdiff >>
rect -840 1025 840 1097
rect -840 981 -768 1025
rect -840 -981 -827 981
rect -781 -981 -768 981
rect 768 981 840 1025
rect -840 -1025 -768 -981
rect 768 -981 781 981
rect 827 -981 840 981
rect 768 -1025 840 -981
rect -840 -1097 840 -1025
<< nsubdiffcont >>
rect -827 -981 -781 981
rect 781 -981 827 981
<< polysilicon >>
rect -680 924 -520 937
rect -680 878 -667 924
rect -533 878 -520 924
rect -680 834 -520 878
rect -680 -878 -520 -834
rect -680 -924 -667 -878
rect -533 -924 -520 -878
rect -680 -937 -520 -924
rect -440 924 -280 937
rect -440 878 -427 924
rect -293 878 -280 924
rect -440 834 -280 878
rect -440 -878 -280 -834
rect -440 -924 -427 -878
rect -293 -924 -280 -878
rect -440 -937 -280 -924
rect -200 924 -40 937
rect -200 878 -187 924
rect -53 878 -40 924
rect -200 834 -40 878
rect -200 -878 -40 -834
rect -200 -924 -187 -878
rect -53 -924 -40 -878
rect -200 -937 -40 -924
rect 40 924 200 937
rect 40 878 53 924
rect 187 878 200 924
rect 40 834 200 878
rect 40 -878 200 -834
rect 40 -924 53 -878
rect 187 -924 200 -878
rect 40 -937 200 -924
rect 280 924 440 937
rect 280 878 293 924
rect 427 878 440 924
rect 280 834 440 878
rect 280 -878 440 -834
rect 280 -924 293 -878
rect 427 -924 440 -878
rect 280 -937 440 -924
rect 520 924 680 937
rect 520 878 533 924
rect 667 878 680 924
rect 520 834 680 878
rect 520 -878 680 -834
rect 520 -924 533 -878
rect 667 -924 680 -878
rect 520 -937 680 -924
<< polycontact >>
rect -667 878 -533 924
rect -667 -924 -533 -878
rect -427 878 -293 924
rect -427 -924 -293 -878
rect -187 878 -53 924
rect -187 -924 -53 -878
rect 53 878 187 924
rect 53 -924 187 -878
rect 293 878 427 924
rect 293 -924 427 -878
rect 533 878 667 924
rect 533 -924 667 -878
<< ppolyres >>
rect -680 -834 -520 834
rect -440 -834 -280 834
rect -200 -834 -40 834
rect 40 -834 200 834
rect 280 -834 440 834
rect 520 -834 680 834
<< metal1 >>
rect -827 1038 827 1084
rect -827 981 -781 1038
rect 781 981 827 1038
rect -678 878 -667 924
rect -533 878 -522 924
rect -438 878 -427 924
rect -293 878 -282 924
rect -198 878 -187 924
rect -53 878 -42 924
rect 42 878 53 924
rect 187 878 198 924
rect 282 878 293 924
rect 427 878 438 924
rect 522 878 533 924
rect 667 878 678 924
rect -678 -924 -667 -878
rect -533 -924 -522 -878
rect -438 -924 -427 -878
rect -293 -924 -282 -878
rect -198 -924 -187 -878
rect -53 -924 -42 -878
rect 42 -924 53 -878
rect 187 -924 198 -878
rect 282 -924 293 -878
rect 427 -924 438 -878
rect 522 -924 533 -878
rect 667 -924 678 -878
rect -827 -1038 -781 -981
rect 781 -1038 827 -981
rect -827 -1084 827 -1038
<< properties >>
string FIXED_BBOX -804 -1061 804 1061
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 8.343 m 1 nx 6 wmin 0.80 lmin 1.00 rho 315 val 3.6k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1
<< end >>
