magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1085 -1646 1085 1646
<< metal2 >>
rect -85 641 85 646
rect -85 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 85 641
rect -85 575 85 613
rect -85 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 85 575
rect -85 509 85 547
rect -85 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 85 509
rect -85 443 85 481
rect -85 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 85 443
rect -85 377 85 415
rect -85 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 85 377
rect -85 311 85 349
rect -85 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 85 311
rect -85 245 85 283
rect -85 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 85 245
rect -85 179 85 217
rect -85 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 85 179
rect -85 113 85 151
rect -85 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 85 113
rect -85 47 85 85
rect -85 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 85 47
rect -85 -19 85 19
rect -85 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 85 -19
rect -85 -85 85 -47
rect -85 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 85 -85
rect -85 -151 85 -113
rect -85 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 85 -151
rect -85 -217 85 -179
rect -85 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 85 -217
rect -85 -283 85 -245
rect -85 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 85 -283
rect -85 -349 85 -311
rect -85 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 85 -349
rect -85 -415 85 -377
rect -85 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 85 -415
rect -85 -481 85 -443
rect -85 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 85 -481
rect -85 -547 85 -509
rect -85 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 85 -547
rect -85 -613 85 -575
rect -85 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 85 -613
rect -85 -646 85 -641
<< via2 >>
rect -80 613 -52 641
rect -14 613 14 641
rect 52 613 80 641
rect -80 547 -52 575
rect -14 547 14 575
rect 52 547 80 575
rect -80 481 -52 509
rect -14 481 14 509
rect 52 481 80 509
rect -80 415 -52 443
rect -14 415 14 443
rect 52 415 80 443
rect -80 349 -52 377
rect -14 349 14 377
rect 52 349 80 377
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect -80 -377 -52 -349
rect -14 -377 14 -349
rect 52 -377 80 -349
rect -80 -443 -52 -415
rect -14 -443 14 -415
rect 52 -443 80 -415
rect -80 -509 -52 -481
rect -14 -509 14 -481
rect 52 -509 80 -481
rect -80 -575 -52 -547
rect -14 -575 14 -547
rect 52 -575 80 -547
rect -80 -641 -52 -613
rect -14 -641 14 -613
rect 52 -641 80 -613
<< metal3 >>
rect -85 641 85 646
rect -85 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 85 641
rect -85 575 85 613
rect -85 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 85 575
rect -85 509 85 547
rect -85 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 85 509
rect -85 443 85 481
rect -85 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 85 443
rect -85 377 85 415
rect -85 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 85 377
rect -85 311 85 349
rect -85 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 85 311
rect -85 245 85 283
rect -85 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 85 245
rect -85 179 85 217
rect -85 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 85 179
rect -85 113 85 151
rect -85 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 85 113
rect -85 47 85 85
rect -85 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 85 47
rect -85 -19 85 19
rect -85 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 85 -19
rect -85 -85 85 -47
rect -85 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 85 -85
rect -85 -151 85 -113
rect -85 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 85 -151
rect -85 -217 85 -179
rect -85 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 85 -217
rect -85 -283 85 -245
rect -85 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 85 -283
rect -85 -349 85 -311
rect -85 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 85 -349
rect -85 -415 85 -377
rect -85 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 85 -415
rect -85 -481 85 -443
rect -85 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 85 -481
rect -85 -547 85 -509
rect -85 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 85 -547
rect -85 -613 85 -575
rect -85 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 85 -613
rect -85 -646 85 -641
<< end >>
