* NGSPICE file created from nverterlayout_flat.ext - technology: gf180mcuC

.subckt nverterlayout_flat VDD VSS OUT IN
X0 OUT IN.t0 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1 OUT IN.t1 VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 IN.n1 IN.t1 25.7638
R1 IN.n0 IN.t0 13.214
R2 IN IN.n1 4.00252
R3 IN.n1 IN.n0 0.0834545
R4 VSS.n1 VSS.t0 1426.49
R5 VSS VSS.t1 9.40995
R6 VSS VSS.n1 2.60126
R7 VSS.n1 VSS.n0 0.039174
R8 OUT OUT.n1 9.44217
R9 OUT OUT.n0 5.13104
R10 VDD.n1 VDD.t0 678.894
R11 VDD.n2 VDD.t1 5.16824
R12 VDD.n2 VDD.n1 3.1505
R13 VDD.n1 VDD.n0 0.0358933
R14 VDD VDD.n2 0.00094665
C0 OUT VDD 0.12f
C1 IN OUT 0.116f
C2 IN VDD 0.144f
.ends

