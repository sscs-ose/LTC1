magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1453 -1174 1453 1174
<< metal1 >>
rect -453 168 453 174
rect -453 142 -447 168
rect -421 142 -385 168
rect -359 142 -323 168
rect -297 142 -261 168
rect -235 142 -199 168
rect -173 142 -137 168
rect -111 142 -75 168
rect -49 142 -13 168
rect 13 142 49 168
rect 75 142 111 168
rect 137 142 173 168
rect 199 142 235 168
rect 261 142 297 168
rect 323 142 359 168
rect 385 142 421 168
rect 447 142 453 168
rect -453 106 453 142
rect -453 80 -447 106
rect -421 80 -385 106
rect -359 80 -323 106
rect -297 80 -261 106
rect -235 80 -199 106
rect -173 80 -137 106
rect -111 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 111 106
rect 137 80 173 106
rect 199 80 235 106
rect 261 80 297 106
rect 323 80 359 106
rect 385 80 421 106
rect 447 80 453 106
rect -453 44 453 80
rect -453 18 -447 44
rect -421 18 -385 44
rect -359 18 -323 44
rect -297 18 -261 44
rect -235 18 -199 44
rect -173 18 -137 44
rect -111 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 111 44
rect 137 18 173 44
rect 199 18 235 44
rect 261 18 297 44
rect 323 18 359 44
rect 385 18 421 44
rect 447 18 453 44
rect -453 -18 453 18
rect -453 -44 -447 -18
rect -421 -44 -385 -18
rect -359 -44 -323 -18
rect -297 -44 -261 -18
rect -235 -44 -199 -18
rect -173 -44 -137 -18
rect -111 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 111 -18
rect 137 -44 173 -18
rect 199 -44 235 -18
rect 261 -44 297 -18
rect 323 -44 359 -18
rect 385 -44 421 -18
rect 447 -44 453 -18
rect -453 -80 453 -44
rect -453 -106 -447 -80
rect -421 -106 -385 -80
rect -359 -106 -323 -80
rect -297 -106 -261 -80
rect -235 -106 -199 -80
rect -173 -106 -137 -80
rect -111 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 111 -80
rect 137 -106 173 -80
rect 199 -106 235 -80
rect 261 -106 297 -80
rect 323 -106 359 -80
rect 385 -106 421 -80
rect 447 -106 453 -80
rect -453 -142 453 -106
rect -453 -168 -447 -142
rect -421 -168 -385 -142
rect -359 -168 -323 -142
rect -297 -168 -261 -142
rect -235 -168 -199 -142
rect -173 -168 -137 -142
rect -111 -168 -75 -142
rect -49 -168 -13 -142
rect 13 -168 49 -142
rect 75 -168 111 -142
rect 137 -168 173 -142
rect 199 -168 235 -142
rect 261 -168 297 -142
rect 323 -168 359 -142
rect 385 -168 421 -142
rect 447 -168 453 -142
rect -453 -174 453 -168
<< via1 >>
rect -447 142 -421 168
rect -385 142 -359 168
rect -323 142 -297 168
rect -261 142 -235 168
rect -199 142 -173 168
rect -137 142 -111 168
rect -75 142 -49 168
rect -13 142 13 168
rect 49 142 75 168
rect 111 142 137 168
rect 173 142 199 168
rect 235 142 261 168
rect 297 142 323 168
rect 359 142 385 168
rect 421 142 447 168
rect -447 80 -421 106
rect -385 80 -359 106
rect -323 80 -297 106
rect -261 80 -235 106
rect -199 80 -173 106
rect -137 80 -111 106
rect -75 80 -49 106
rect -13 80 13 106
rect 49 80 75 106
rect 111 80 137 106
rect 173 80 199 106
rect 235 80 261 106
rect 297 80 323 106
rect 359 80 385 106
rect 421 80 447 106
rect -447 18 -421 44
rect -385 18 -359 44
rect -323 18 -297 44
rect -261 18 -235 44
rect -199 18 -173 44
rect -137 18 -111 44
rect -75 18 -49 44
rect -13 18 13 44
rect 49 18 75 44
rect 111 18 137 44
rect 173 18 199 44
rect 235 18 261 44
rect 297 18 323 44
rect 359 18 385 44
rect 421 18 447 44
rect -447 -44 -421 -18
rect -385 -44 -359 -18
rect -323 -44 -297 -18
rect -261 -44 -235 -18
rect -199 -44 -173 -18
rect -137 -44 -111 -18
rect -75 -44 -49 -18
rect -13 -44 13 -18
rect 49 -44 75 -18
rect 111 -44 137 -18
rect 173 -44 199 -18
rect 235 -44 261 -18
rect 297 -44 323 -18
rect 359 -44 385 -18
rect 421 -44 447 -18
rect -447 -106 -421 -80
rect -385 -106 -359 -80
rect -323 -106 -297 -80
rect -261 -106 -235 -80
rect -199 -106 -173 -80
rect -137 -106 -111 -80
rect -75 -106 -49 -80
rect -13 -106 13 -80
rect 49 -106 75 -80
rect 111 -106 137 -80
rect 173 -106 199 -80
rect 235 -106 261 -80
rect 297 -106 323 -80
rect 359 -106 385 -80
rect 421 -106 447 -80
rect -447 -168 -421 -142
rect -385 -168 -359 -142
rect -323 -168 -297 -142
rect -261 -168 -235 -142
rect -199 -168 -173 -142
rect -137 -168 -111 -142
rect -75 -168 -49 -142
rect -13 -168 13 -142
rect 49 -168 75 -142
rect 111 -168 137 -142
rect 173 -168 199 -142
rect 235 -168 261 -142
rect 297 -168 323 -142
rect 359 -168 385 -142
rect 421 -168 447 -142
<< metal2 >>
rect -453 168 453 174
rect -453 142 -447 168
rect -421 142 -385 168
rect -359 142 -323 168
rect -297 142 -261 168
rect -235 142 -199 168
rect -173 142 -137 168
rect -111 142 -75 168
rect -49 142 -13 168
rect 13 142 49 168
rect 75 142 111 168
rect 137 142 173 168
rect 199 142 235 168
rect 261 142 297 168
rect 323 142 359 168
rect 385 142 421 168
rect 447 142 453 168
rect -453 106 453 142
rect -453 80 -447 106
rect -421 80 -385 106
rect -359 80 -323 106
rect -297 80 -261 106
rect -235 80 -199 106
rect -173 80 -137 106
rect -111 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 111 106
rect 137 80 173 106
rect 199 80 235 106
rect 261 80 297 106
rect 323 80 359 106
rect 385 80 421 106
rect 447 80 453 106
rect -453 44 453 80
rect -453 18 -447 44
rect -421 18 -385 44
rect -359 18 -323 44
rect -297 18 -261 44
rect -235 18 -199 44
rect -173 18 -137 44
rect -111 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 111 44
rect 137 18 173 44
rect 199 18 235 44
rect 261 18 297 44
rect 323 18 359 44
rect 385 18 421 44
rect 447 18 453 44
rect -453 -18 453 18
rect -453 -44 -447 -18
rect -421 -44 -385 -18
rect -359 -44 -323 -18
rect -297 -44 -261 -18
rect -235 -44 -199 -18
rect -173 -44 -137 -18
rect -111 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 111 -18
rect 137 -44 173 -18
rect 199 -44 235 -18
rect 261 -44 297 -18
rect 323 -44 359 -18
rect 385 -44 421 -18
rect 447 -44 453 -18
rect -453 -80 453 -44
rect -453 -106 -447 -80
rect -421 -106 -385 -80
rect -359 -106 -323 -80
rect -297 -106 -261 -80
rect -235 -106 -199 -80
rect -173 -106 -137 -80
rect -111 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 111 -80
rect 137 -106 173 -80
rect 199 -106 235 -80
rect 261 -106 297 -80
rect 323 -106 359 -80
rect 385 -106 421 -80
rect 447 -106 453 -80
rect -453 -142 453 -106
rect -453 -168 -447 -142
rect -421 -168 -385 -142
rect -359 -168 -323 -142
rect -297 -168 -261 -142
rect -235 -168 -199 -142
rect -173 -168 -137 -142
rect -111 -168 -75 -142
rect -49 -168 -13 -142
rect 13 -168 49 -142
rect 75 -168 111 -142
rect 137 -168 173 -142
rect 199 -168 235 -142
rect 261 -168 297 -142
rect 323 -168 359 -142
rect 385 -168 421 -142
rect 447 -168 453 -142
rect -453 -174 453 -168
<< end >>
