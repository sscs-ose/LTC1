* NGSPICE file created from nand2_mag_flat.ext - technology: gf180mcuC

.subckt pex_nand2_mag IN1 VSS VDD OUT IN2
X0 OUT IN1.t0 a_168_68# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1 OUT IN2.t0 VDD.t4 VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 a_168_68# IN2.t1 VSS.t2 VSS.t1 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3 VDD IN1.t1 OUT.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 IN1.n0 IN1.t0 31.528
R1 IN1.n0 IN1.t1 15.3826
R2 IN1 IN1.n0 8.88964
R3 OUT.n3 OUT.n0 7.11377
R4 OUT.n3 OUT.n2 3.25706
R5 OUT.n2 OUT.t1 2.2755
R6 OUT.n2 OUT.n1 2.2755
R7 OUT OUT.n3 0.191955
R8 VSS.n1 VSS.t0 596.558
R9 VSS.n1 VSS.t1 397.707
R10 VSS.n3 VSS.t2 7.30963
R11 VSS.n3 VSS.n2 2.6005
R12 VSS.n2 VSS.n1 2.6005
R13 VSS.n2 VSS.n0 0.553132
R14 VSS VSS.n3 0.00545413
R15 IN2.n0 IN2.t0 30.9379
R16 IN2.n0 IN2.t1 21.6422
R17 IN2 IN2.n0 4.12052
R18 VDD.n2 VDD.t0 193.183
R19 VDD.n2 VDD.t3 109.849
R20 VDD.n4 VDD.n0 5.23971
R21 VDD VDD.t4 5.21184
R22 VDD.n4 VDD.n3 3.1505
R23 VDD.n3 VDD.n2 3.1505
R24 VDD.n3 VDD.n1 0.089483
R25 VDD VDD.n4 0.00166129
C0 a_168_68# IN2 0.00347f
C1 OUT IN2 0.0929f
C2 IN1 IN2 0.0466f
C3 VDD a_168_68# 3.14e-19
C4 VDD OUT 0.209f
C5 VDD IN1 0.225f
C6 OUT a_168_68# 0.069f
C7 IN1 a_168_68# 0.00348f
C8 VDD IN2 0.158f
C9 OUT IN1 0.256f
.ends

