magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -4336 -1112 4336 1112
<< metal2 >>
rect -3336 107 3336 112
rect -3336 79 -3331 107
rect -3303 79 -3269 107
rect -3241 79 -3207 107
rect -3179 79 -3145 107
rect -3117 79 -3083 107
rect -3055 79 -3021 107
rect -2993 79 -2959 107
rect -2931 79 -2897 107
rect -2869 79 -2835 107
rect -2807 79 -2773 107
rect -2745 79 -2711 107
rect -2683 79 -2649 107
rect -2621 79 -2587 107
rect -2559 79 -2525 107
rect -2497 79 -2463 107
rect -2435 79 -2401 107
rect -2373 79 -2339 107
rect -2311 79 -2277 107
rect -2249 79 -2215 107
rect -2187 79 -2153 107
rect -2125 79 -2091 107
rect -2063 79 -2029 107
rect -2001 79 -1967 107
rect -1939 79 -1905 107
rect -1877 79 -1843 107
rect -1815 79 -1781 107
rect -1753 79 -1719 107
rect -1691 79 -1657 107
rect -1629 79 -1595 107
rect -1567 79 -1533 107
rect -1505 79 -1471 107
rect -1443 79 -1409 107
rect -1381 79 -1347 107
rect -1319 79 -1285 107
rect -1257 79 -1223 107
rect -1195 79 -1161 107
rect -1133 79 -1099 107
rect -1071 79 -1037 107
rect -1009 79 -975 107
rect -947 79 -913 107
rect -885 79 -851 107
rect -823 79 -789 107
rect -761 79 -727 107
rect -699 79 -665 107
rect -637 79 -603 107
rect -575 79 -541 107
rect -513 79 -479 107
rect -451 79 -417 107
rect -389 79 -355 107
rect -327 79 -293 107
rect -265 79 -231 107
rect -203 79 -169 107
rect -141 79 -107 107
rect -79 79 -45 107
rect -17 79 17 107
rect 45 79 79 107
rect 107 79 141 107
rect 169 79 203 107
rect 231 79 265 107
rect 293 79 327 107
rect 355 79 389 107
rect 417 79 451 107
rect 479 79 513 107
rect 541 79 575 107
rect 603 79 637 107
rect 665 79 699 107
rect 727 79 761 107
rect 789 79 823 107
rect 851 79 885 107
rect 913 79 947 107
rect 975 79 1009 107
rect 1037 79 1071 107
rect 1099 79 1133 107
rect 1161 79 1195 107
rect 1223 79 1257 107
rect 1285 79 1319 107
rect 1347 79 1381 107
rect 1409 79 1443 107
rect 1471 79 1505 107
rect 1533 79 1567 107
rect 1595 79 1629 107
rect 1657 79 1691 107
rect 1719 79 1753 107
rect 1781 79 1815 107
rect 1843 79 1877 107
rect 1905 79 1939 107
rect 1967 79 2001 107
rect 2029 79 2063 107
rect 2091 79 2125 107
rect 2153 79 2187 107
rect 2215 79 2249 107
rect 2277 79 2311 107
rect 2339 79 2373 107
rect 2401 79 2435 107
rect 2463 79 2497 107
rect 2525 79 2559 107
rect 2587 79 2621 107
rect 2649 79 2683 107
rect 2711 79 2745 107
rect 2773 79 2807 107
rect 2835 79 2869 107
rect 2897 79 2931 107
rect 2959 79 2993 107
rect 3021 79 3055 107
rect 3083 79 3117 107
rect 3145 79 3179 107
rect 3207 79 3241 107
rect 3269 79 3303 107
rect 3331 79 3336 107
rect -3336 45 3336 79
rect -3336 17 -3331 45
rect -3303 17 -3269 45
rect -3241 17 -3207 45
rect -3179 17 -3145 45
rect -3117 17 -3083 45
rect -3055 17 -3021 45
rect -2993 17 -2959 45
rect -2931 17 -2897 45
rect -2869 17 -2835 45
rect -2807 17 -2773 45
rect -2745 17 -2711 45
rect -2683 17 -2649 45
rect -2621 17 -2587 45
rect -2559 17 -2525 45
rect -2497 17 -2463 45
rect -2435 17 -2401 45
rect -2373 17 -2339 45
rect -2311 17 -2277 45
rect -2249 17 -2215 45
rect -2187 17 -2153 45
rect -2125 17 -2091 45
rect -2063 17 -2029 45
rect -2001 17 -1967 45
rect -1939 17 -1905 45
rect -1877 17 -1843 45
rect -1815 17 -1781 45
rect -1753 17 -1719 45
rect -1691 17 -1657 45
rect -1629 17 -1595 45
rect -1567 17 -1533 45
rect -1505 17 -1471 45
rect -1443 17 -1409 45
rect -1381 17 -1347 45
rect -1319 17 -1285 45
rect -1257 17 -1223 45
rect -1195 17 -1161 45
rect -1133 17 -1099 45
rect -1071 17 -1037 45
rect -1009 17 -975 45
rect -947 17 -913 45
rect -885 17 -851 45
rect -823 17 -789 45
rect -761 17 -727 45
rect -699 17 -665 45
rect -637 17 -603 45
rect -575 17 -541 45
rect -513 17 -479 45
rect -451 17 -417 45
rect -389 17 -355 45
rect -327 17 -293 45
rect -265 17 -231 45
rect -203 17 -169 45
rect -141 17 -107 45
rect -79 17 -45 45
rect -17 17 17 45
rect 45 17 79 45
rect 107 17 141 45
rect 169 17 203 45
rect 231 17 265 45
rect 293 17 327 45
rect 355 17 389 45
rect 417 17 451 45
rect 479 17 513 45
rect 541 17 575 45
rect 603 17 637 45
rect 665 17 699 45
rect 727 17 761 45
rect 789 17 823 45
rect 851 17 885 45
rect 913 17 947 45
rect 975 17 1009 45
rect 1037 17 1071 45
rect 1099 17 1133 45
rect 1161 17 1195 45
rect 1223 17 1257 45
rect 1285 17 1319 45
rect 1347 17 1381 45
rect 1409 17 1443 45
rect 1471 17 1505 45
rect 1533 17 1567 45
rect 1595 17 1629 45
rect 1657 17 1691 45
rect 1719 17 1753 45
rect 1781 17 1815 45
rect 1843 17 1877 45
rect 1905 17 1939 45
rect 1967 17 2001 45
rect 2029 17 2063 45
rect 2091 17 2125 45
rect 2153 17 2187 45
rect 2215 17 2249 45
rect 2277 17 2311 45
rect 2339 17 2373 45
rect 2401 17 2435 45
rect 2463 17 2497 45
rect 2525 17 2559 45
rect 2587 17 2621 45
rect 2649 17 2683 45
rect 2711 17 2745 45
rect 2773 17 2807 45
rect 2835 17 2869 45
rect 2897 17 2931 45
rect 2959 17 2993 45
rect 3021 17 3055 45
rect 3083 17 3117 45
rect 3145 17 3179 45
rect 3207 17 3241 45
rect 3269 17 3303 45
rect 3331 17 3336 45
rect -3336 -17 3336 17
rect -3336 -45 -3331 -17
rect -3303 -45 -3269 -17
rect -3241 -45 -3207 -17
rect -3179 -45 -3145 -17
rect -3117 -45 -3083 -17
rect -3055 -45 -3021 -17
rect -2993 -45 -2959 -17
rect -2931 -45 -2897 -17
rect -2869 -45 -2835 -17
rect -2807 -45 -2773 -17
rect -2745 -45 -2711 -17
rect -2683 -45 -2649 -17
rect -2621 -45 -2587 -17
rect -2559 -45 -2525 -17
rect -2497 -45 -2463 -17
rect -2435 -45 -2401 -17
rect -2373 -45 -2339 -17
rect -2311 -45 -2277 -17
rect -2249 -45 -2215 -17
rect -2187 -45 -2153 -17
rect -2125 -45 -2091 -17
rect -2063 -45 -2029 -17
rect -2001 -45 -1967 -17
rect -1939 -45 -1905 -17
rect -1877 -45 -1843 -17
rect -1815 -45 -1781 -17
rect -1753 -45 -1719 -17
rect -1691 -45 -1657 -17
rect -1629 -45 -1595 -17
rect -1567 -45 -1533 -17
rect -1505 -45 -1471 -17
rect -1443 -45 -1409 -17
rect -1381 -45 -1347 -17
rect -1319 -45 -1285 -17
rect -1257 -45 -1223 -17
rect -1195 -45 -1161 -17
rect -1133 -45 -1099 -17
rect -1071 -45 -1037 -17
rect -1009 -45 -975 -17
rect -947 -45 -913 -17
rect -885 -45 -851 -17
rect -823 -45 -789 -17
rect -761 -45 -727 -17
rect -699 -45 -665 -17
rect -637 -45 -603 -17
rect -575 -45 -541 -17
rect -513 -45 -479 -17
rect -451 -45 -417 -17
rect -389 -45 -355 -17
rect -327 -45 -293 -17
rect -265 -45 -231 -17
rect -203 -45 -169 -17
rect -141 -45 -107 -17
rect -79 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 79 -17
rect 107 -45 141 -17
rect 169 -45 203 -17
rect 231 -45 265 -17
rect 293 -45 327 -17
rect 355 -45 389 -17
rect 417 -45 451 -17
rect 479 -45 513 -17
rect 541 -45 575 -17
rect 603 -45 637 -17
rect 665 -45 699 -17
rect 727 -45 761 -17
rect 789 -45 823 -17
rect 851 -45 885 -17
rect 913 -45 947 -17
rect 975 -45 1009 -17
rect 1037 -45 1071 -17
rect 1099 -45 1133 -17
rect 1161 -45 1195 -17
rect 1223 -45 1257 -17
rect 1285 -45 1319 -17
rect 1347 -45 1381 -17
rect 1409 -45 1443 -17
rect 1471 -45 1505 -17
rect 1533 -45 1567 -17
rect 1595 -45 1629 -17
rect 1657 -45 1691 -17
rect 1719 -45 1753 -17
rect 1781 -45 1815 -17
rect 1843 -45 1877 -17
rect 1905 -45 1939 -17
rect 1967 -45 2001 -17
rect 2029 -45 2063 -17
rect 2091 -45 2125 -17
rect 2153 -45 2187 -17
rect 2215 -45 2249 -17
rect 2277 -45 2311 -17
rect 2339 -45 2373 -17
rect 2401 -45 2435 -17
rect 2463 -45 2497 -17
rect 2525 -45 2559 -17
rect 2587 -45 2621 -17
rect 2649 -45 2683 -17
rect 2711 -45 2745 -17
rect 2773 -45 2807 -17
rect 2835 -45 2869 -17
rect 2897 -45 2931 -17
rect 2959 -45 2993 -17
rect 3021 -45 3055 -17
rect 3083 -45 3117 -17
rect 3145 -45 3179 -17
rect 3207 -45 3241 -17
rect 3269 -45 3303 -17
rect 3331 -45 3336 -17
rect -3336 -79 3336 -45
rect -3336 -107 -3331 -79
rect -3303 -107 -3269 -79
rect -3241 -107 -3207 -79
rect -3179 -107 -3145 -79
rect -3117 -107 -3083 -79
rect -3055 -107 -3021 -79
rect -2993 -107 -2959 -79
rect -2931 -107 -2897 -79
rect -2869 -107 -2835 -79
rect -2807 -107 -2773 -79
rect -2745 -107 -2711 -79
rect -2683 -107 -2649 -79
rect -2621 -107 -2587 -79
rect -2559 -107 -2525 -79
rect -2497 -107 -2463 -79
rect -2435 -107 -2401 -79
rect -2373 -107 -2339 -79
rect -2311 -107 -2277 -79
rect -2249 -107 -2215 -79
rect -2187 -107 -2153 -79
rect -2125 -107 -2091 -79
rect -2063 -107 -2029 -79
rect -2001 -107 -1967 -79
rect -1939 -107 -1905 -79
rect -1877 -107 -1843 -79
rect -1815 -107 -1781 -79
rect -1753 -107 -1719 -79
rect -1691 -107 -1657 -79
rect -1629 -107 -1595 -79
rect -1567 -107 -1533 -79
rect -1505 -107 -1471 -79
rect -1443 -107 -1409 -79
rect -1381 -107 -1347 -79
rect -1319 -107 -1285 -79
rect -1257 -107 -1223 -79
rect -1195 -107 -1161 -79
rect -1133 -107 -1099 -79
rect -1071 -107 -1037 -79
rect -1009 -107 -975 -79
rect -947 -107 -913 -79
rect -885 -107 -851 -79
rect -823 -107 -789 -79
rect -761 -107 -727 -79
rect -699 -107 -665 -79
rect -637 -107 -603 -79
rect -575 -107 -541 -79
rect -513 -107 -479 -79
rect -451 -107 -417 -79
rect -389 -107 -355 -79
rect -327 -107 -293 -79
rect -265 -107 -231 -79
rect -203 -107 -169 -79
rect -141 -107 -107 -79
rect -79 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 79 -79
rect 107 -107 141 -79
rect 169 -107 203 -79
rect 231 -107 265 -79
rect 293 -107 327 -79
rect 355 -107 389 -79
rect 417 -107 451 -79
rect 479 -107 513 -79
rect 541 -107 575 -79
rect 603 -107 637 -79
rect 665 -107 699 -79
rect 727 -107 761 -79
rect 789 -107 823 -79
rect 851 -107 885 -79
rect 913 -107 947 -79
rect 975 -107 1009 -79
rect 1037 -107 1071 -79
rect 1099 -107 1133 -79
rect 1161 -107 1195 -79
rect 1223 -107 1257 -79
rect 1285 -107 1319 -79
rect 1347 -107 1381 -79
rect 1409 -107 1443 -79
rect 1471 -107 1505 -79
rect 1533 -107 1567 -79
rect 1595 -107 1629 -79
rect 1657 -107 1691 -79
rect 1719 -107 1753 -79
rect 1781 -107 1815 -79
rect 1843 -107 1877 -79
rect 1905 -107 1939 -79
rect 1967 -107 2001 -79
rect 2029 -107 2063 -79
rect 2091 -107 2125 -79
rect 2153 -107 2187 -79
rect 2215 -107 2249 -79
rect 2277 -107 2311 -79
rect 2339 -107 2373 -79
rect 2401 -107 2435 -79
rect 2463 -107 2497 -79
rect 2525 -107 2559 -79
rect 2587 -107 2621 -79
rect 2649 -107 2683 -79
rect 2711 -107 2745 -79
rect 2773 -107 2807 -79
rect 2835 -107 2869 -79
rect 2897 -107 2931 -79
rect 2959 -107 2993 -79
rect 3021 -107 3055 -79
rect 3083 -107 3117 -79
rect 3145 -107 3179 -79
rect 3207 -107 3241 -79
rect 3269 -107 3303 -79
rect 3331 -107 3336 -79
rect -3336 -112 3336 -107
<< via2 >>
rect -3331 79 -3303 107
rect -3269 79 -3241 107
rect -3207 79 -3179 107
rect -3145 79 -3117 107
rect -3083 79 -3055 107
rect -3021 79 -2993 107
rect -2959 79 -2931 107
rect -2897 79 -2869 107
rect -2835 79 -2807 107
rect -2773 79 -2745 107
rect -2711 79 -2683 107
rect -2649 79 -2621 107
rect -2587 79 -2559 107
rect -2525 79 -2497 107
rect -2463 79 -2435 107
rect -2401 79 -2373 107
rect -2339 79 -2311 107
rect -2277 79 -2249 107
rect -2215 79 -2187 107
rect -2153 79 -2125 107
rect -2091 79 -2063 107
rect -2029 79 -2001 107
rect -1967 79 -1939 107
rect -1905 79 -1877 107
rect -1843 79 -1815 107
rect -1781 79 -1753 107
rect -1719 79 -1691 107
rect -1657 79 -1629 107
rect -1595 79 -1567 107
rect -1533 79 -1505 107
rect -1471 79 -1443 107
rect -1409 79 -1381 107
rect -1347 79 -1319 107
rect -1285 79 -1257 107
rect -1223 79 -1195 107
rect -1161 79 -1133 107
rect -1099 79 -1071 107
rect -1037 79 -1009 107
rect -975 79 -947 107
rect -913 79 -885 107
rect -851 79 -823 107
rect -789 79 -761 107
rect -727 79 -699 107
rect -665 79 -637 107
rect -603 79 -575 107
rect -541 79 -513 107
rect -479 79 -451 107
rect -417 79 -389 107
rect -355 79 -327 107
rect -293 79 -265 107
rect -231 79 -203 107
rect -169 79 -141 107
rect -107 79 -79 107
rect -45 79 -17 107
rect 17 79 45 107
rect 79 79 107 107
rect 141 79 169 107
rect 203 79 231 107
rect 265 79 293 107
rect 327 79 355 107
rect 389 79 417 107
rect 451 79 479 107
rect 513 79 541 107
rect 575 79 603 107
rect 637 79 665 107
rect 699 79 727 107
rect 761 79 789 107
rect 823 79 851 107
rect 885 79 913 107
rect 947 79 975 107
rect 1009 79 1037 107
rect 1071 79 1099 107
rect 1133 79 1161 107
rect 1195 79 1223 107
rect 1257 79 1285 107
rect 1319 79 1347 107
rect 1381 79 1409 107
rect 1443 79 1471 107
rect 1505 79 1533 107
rect 1567 79 1595 107
rect 1629 79 1657 107
rect 1691 79 1719 107
rect 1753 79 1781 107
rect 1815 79 1843 107
rect 1877 79 1905 107
rect 1939 79 1967 107
rect 2001 79 2029 107
rect 2063 79 2091 107
rect 2125 79 2153 107
rect 2187 79 2215 107
rect 2249 79 2277 107
rect 2311 79 2339 107
rect 2373 79 2401 107
rect 2435 79 2463 107
rect 2497 79 2525 107
rect 2559 79 2587 107
rect 2621 79 2649 107
rect 2683 79 2711 107
rect 2745 79 2773 107
rect 2807 79 2835 107
rect 2869 79 2897 107
rect 2931 79 2959 107
rect 2993 79 3021 107
rect 3055 79 3083 107
rect 3117 79 3145 107
rect 3179 79 3207 107
rect 3241 79 3269 107
rect 3303 79 3331 107
rect -3331 17 -3303 45
rect -3269 17 -3241 45
rect -3207 17 -3179 45
rect -3145 17 -3117 45
rect -3083 17 -3055 45
rect -3021 17 -2993 45
rect -2959 17 -2931 45
rect -2897 17 -2869 45
rect -2835 17 -2807 45
rect -2773 17 -2745 45
rect -2711 17 -2683 45
rect -2649 17 -2621 45
rect -2587 17 -2559 45
rect -2525 17 -2497 45
rect -2463 17 -2435 45
rect -2401 17 -2373 45
rect -2339 17 -2311 45
rect -2277 17 -2249 45
rect -2215 17 -2187 45
rect -2153 17 -2125 45
rect -2091 17 -2063 45
rect -2029 17 -2001 45
rect -1967 17 -1939 45
rect -1905 17 -1877 45
rect -1843 17 -1815 45
rect -1781 17 -1753 45
rect -1719 17 -1691 45
rect -1657 17 -1629 45
rect -1595 17 -1567 45
rect -1533 17 -1505 45
rect -1471 17 -1443 45
rect -1409 17 -1381 45
rect -1347 17 -1319 45
rect -1285 17 -1257 45
rect -1223 17 -1195 45
rect -1161 17 -1133 45
rect -1099 17 -1071 45
rect -1037 17 -1009 45
rect -975 17 -947 45
rect -913 17 -885 45
rect -851 17 -823 45
rect -789 17 -761 45
rect -727 17 -699 45
rect -665 17 -637 45
rect -603 17 -575 45
rect -541 17 -513 45
rect -479 17 -451 45
rect -417 17 -389 45
rect -355 17 -327 45
rect -293 17 -265 45
rect -231 17 -203 45
rect -169 17 -141 45
rect -107 17 -79 45
rect -45 17 -17 45
rect 17 17 45 45
rect 79 17 107 45
rect 141 17 169 45
rect 203 17 231 45
rect 265 17 293 45
rect 327 17 355 45
rect 389 17 417 45
rect 451 17 479 45
rect 513 17 541 45
rect 575 17 603 45
rect 637 17 665 45
rect 699 17 727 45
rect 761 17 789 45
rect 823 17 851 45
rect 885 17 913 45
rect 947 17 975 45
rect 1009 17 1037 45
rect 1071 17 1099 45
rect 1133 17 1161 45
rect 1195 17 1223 45
rect 1257 17 1285 45
rect 1319 17 1347 45
rect 1381 17 1409 45
rect 1443 17 1471 45
rect 1505 17 1533 45
rect 1567 17 1595 45
rect 1629 17 1657 45
rect 1691 17 1719 45
rect 1753 17 1781 45
rect 1815 17 1843 45
rect 1877 17 1905 45
rect 1939 17 1967 45
rect 2001 17 2029 45
rect 2063 17 2091 45
rect 2125 17 2153 45
rect 2187 17 2215 45
rect 2249 17 2277 45
rect 2311 17 2339 45
rect 2373 17 2401 45
rect 2435 17 2463 45
rect 2497 17 2525 45
rect 2559 17 2587 45
rect 2621 17 2649 45
rect 2683 17 2711 45
rect 2745 17 2773 45
rect 2807 17 2835 45
rect 2869 17 2897 45
rect 2931 17 2959 45
rect 2993 17 3021 45
rect 3055 17 3083 45
rect 3117 17 3145 45
rect 3179 17 3207 45
rect 3241 17 3269 45
rect 3303 17 3331 45
rect -3331 -45 -3303 -17
rect -3269 -45 -3241 -17
rect -3207 -45 -3179 -17
rect -3145 -45 -3117 -17
rect -3083 -45 -3055 -17
rect -3021 -45 -2993 -17
rect -2959 -45 -2931 -17
rect -2897 -45 -2869 -17
rect -2835 -45 -2807 -17
rect -2773 -45 -2745 -17
rect -2711 -45 -2683 -17
rect -2649 -45 -2621 -17
rect -2587 -45 -2559 -17
rect -2525 -45 -2497 -17
rect -2463 -45 -2435 -17
rect -2401 -45 -2373 -17
rect -2339 -45 -2311 -17
rect -2277 -45 -2249 -17
rect -2215 -45 -2187 -17
rect -2153 -45 -2125 -17
rect -2091 -45 -2063 -17
rect -2029 -45 -2001 -17
rect -1967 -45 -1939 -17
rect -1905 -45 -1877 -17
rect -1843 -45 -1815 -17
rect -1781 -45 -1753 -17
rect -1719 -45 -1691 -17
rect -1657 -45 -1629 -17
rect -1595 -45 -1567 -17
rect -1533 -45 -1505 -17
rect -1471 -45 -1443 -17
rect -1409 -45 -1381 -17
rect -1347 -45 -1319 -17
rect -1285 -45 -1257 -17
rect -1223 -45 -1195 -17
rect -1161 -45 -1133 -17
rect -1099 -45 -1071 -17
rect -1037 -45 -1009 -17
rect -975 -45 -947 -17
rect -913 -45 -885 -17
rect -851 -45 -823 -17
rect -789 -45 -761 -17
rect -727 -45 -699 -17
rect -665 -45 -637 -17
rect -603 -45 -575 -17
rect -541 -45 -513 -17
rect -479 -45 -451 -17
rect -417 -45 -389 -17
rect -355 -45 -327 -17
rect -293 -45 -265 -17
rect -231 -45 -203 -17
rect -169 -45 -141 -17
rect -107 -45 -79 -17
rect -45 -45 -17 -17
rect 17 -45 45 -17
rect 79 -45 107 -17
rect 141 -45 169 -17
rect 203 -45 231 -17
rect 265 -45 293 -17
rect 327 -45 355 -17
rect 389 -45 417 -17
rect 451 -45 479 -17
rect 513 -45 541 -17
rect 575 -45 603 -17
rect 637 -45 665 -17
rect 699 -45 727 -17
rect 761 -45 789 -17
rect 823 -45 851 -17
rect 885 -45 913 -17
rect 947 -45 975 -17
rect 1009 -45 1037 -17
rect 1071 -45 1099 -17
rect 1133 -45 1161 -17
rect 1195 -45 1223 -17
rect 1257 -45 1285 -17
rect 1319 -45 1347 -17
rect 1381 -45 1409 -17
rect 1443 -45 1471 -17
rect 1505 -45 1533 -17
rect 1567 -45 1595 -17
rect 1629 -45 1657 -17
rect 1691 -45 1719 -17
rect 1753 -45 1781 -17
rect 1815 -45 1843 -17
rect 1877 -45 1905 -17
rect 1939 -45 1967 -17
rect 2001 -45 2029 -17
rect 2063 -45 2091 -17
rect 2125 -45 2153 -17
rect 2187 -45 2215 -17
rect 2249 -45 2277 -17
rect 2311 -45 2339 -17
rect 2373 -45 2401 -17
rect 2435 -45 2463 -17
rect 2497 -45 2525 -17
rect 2559 -45 2587 -17
rect 2621 -45 2649 -17
rect 2683 -45 2711 -17
rect 2745 -45 2773 -17
rect 2807 -45 2835 -17
rect 2869 -45 2897 -17
rect 2931 -45 2959 -17
rect 2993 -45 3021 -17
rect 3055 -45 3083 -17
rect 3117 -45 3145 -17
rect 3179 -45 3207 -17
rect 3241 -45 3269 -17
rect 3303 -45 3331 -17
rect -3331 -107 -3303 -79
rect -3269 -107 -3241 -79
rect -3207 -107 -3179 -79
rect -3145 -107 -3117 -79
rect -3083 -107 -3055 -79
rect -3021 -107 -2993 -79
rect -2959 -107 -2931 -79
rect -2897 -107 -2869 -79
rect -2835 -107 -2807 -79
rect -2773 -107 -2745 -79
rect -2711 -107 -2683 -79
rect -2649 -107 -2621 -79
rect -2587 -107 -2559 -79
rect -2525 -107 -2497 -79
rect -2463 -107 -2435 -79
rect -2401 -107 -2373 -79
rect -2339 -107 -2311 -79
rect -2277 -107 -2249 -79
rect -2215 -107 -2187 -79
rect -2153 -107 -2125 -79
rect -2091 -107 -2063 -79
rect -2029 -107 -2001 -79
rect -1967 -107 -1939 -79
rect -1905 -107 -1877 -79
rect -1843 -107 -1815 -79
rect -1781 -107 -1753 -79
rect -1719 -107 -1691 -79
rect -1657 -107 -1629 -79
rect -1595 -107 -1567 -79
rect -1533 -107 -1505 -79
rect -1471 -107 -1443 -79
rect -1409 -107 -1381 -79
rect -1347 -107 -1319 -79
rect -1285 -107 -1257 -79
rect -1223 -107 -1195 -79
rect -1161 -107 -1133 -79
rect -1099 -107 -1071 -79
rect -1037 -107 -1009 -79
rect -975 -107 -947 -79
rect -913 -107 -885 -79
rect -851 -107 -823 -79
rect -789 -107 -761 -79
rect -727 -107 -699 -79
rect -665 -107 -637 -79
rect -603 -107 -575 -79
rect -541 -107 -513 -79
rect -479 -107 -451 -79
rect -417 -107 -389 -79
rect -355 -107 -327 -79
rect -293 -107 -265 -79
rect -231 -107 -203 -79
rect -169 -107 -141 -79
rect -107 -107 -79 -79
rect -45 -107 -17 -79
rect 17 -107 45 -79
rect 79 -107 107 -79
rect 141 -107 169 -79
rect 203 -107 231 -79
rect 265 -107 293 -79
rect 327 -107 355 -79
rect 389 -107 417 -79
rect 451 -107 479 -79
rect 513 -107 541 -79
rect 575 -107 603 -79
rect 637 -107 665 -79
rect 699 -107 727 -79
rect 761 -107 789 -79
rect 823 -107 851 -79
rect 885 -107 913 -79
rect 947 -107 975 -79
rect 1009 -107 1037 -79
rect 1071 -107 1099 -79
rect 1133 -107 1161 -79
rect 1195 -107 1223 -79
rect 1257 -107 1285 -79
rect 1319 -107 1347 -79
rect 1381 -107 1409 -79
rect 1443 -107 1471 -79
rect 1505 -107 1533 -79
rect 1567 -107 1595 -79
rect 1629 -107 1657 -79
rect 1691 -107 1719 -79
rect 1753 -107 1781 -79
rect 1815 -107 1843 -79
rect 1877 -107 1905 -79
rect 1939 -107 1967 -79
rect 2001 -107 2029 -79
rect 2063 -107 2091 -79
rect 2125 -107 2153 -79
rect 2187 -107 2215 -79
rect 2249 -107 2277 -79
rect 2311 -107 2339 -79
rect 2373 -107 2401 -79
rect 2435 -107 2463 -79
rect 2497 -107 2525 -79
rect 2559 -107 2587 -79
rect 2621 -107 2649 -79
rect 2683 -107 2711 -79
rect 2745 -107 2773 -79
rect 2807 -107 2835 -79
rect 2869 -107 2897 -79
rect 2931 -107 2959 -79
rect 2993 -107 3021 -79
rect 3055 -107 3083 -79
rect 3117 -107 3145 -79
rect 3179 -107 3207 -79
rect 3241 -107 3269 -79
rect 3303 -107 3331 -79
<< metal3 >>
rect -3336 107 3336 112
rect -3336 79 -3331 107
rect -3303 79 -3269 107
rect -3241 79 -3207 107
rect -3179 79 -3145 107
rect -3117 79 -3083 107
rect -3055 79 -3021 107
rect -2993 79 -2959 107
rect -2931 79 -2897 107
rect -2869 79 -2835 107
rect -2807 79 -2773 107
rect -2745 79 -2711 107
rect -2683 79 -2649 107
rect -2621 79 -2587 107
rect -2559 79 -2525 107
rect -2497 79 -2463 107
rect -2435 79 -2401 107
rect -2373 79 -2339 107
rect -2311 79 -2277 107
rect -2249 79 -2215 107
rect -2187 79 -2153 107
rect -2125 79 -2091 107
rect -2063 79 -2029 107
rect -2001 79 -1967 107
rect -1939 79 -1905 107
rect -1877 79 -1843 107
rect -1815 79 -1781 107
rect -1753 79 -1719 107
rect -1691 79 -1657 107
rect -1629 79 -1595 107
rect -1567 79 -1533 107
rect -1505 79 -1471 107
rect -1443 79 -1409 107
rect -1381 79 -1347 107
rect -1319 79 -1285 107
rect -1257 79 -1223 107
rect -1195 79 -1161 107
rect -1133 79 -1099 107
rect -1071 79 -1037 107
rect -1009 79 -975 107
rect -947 79 -913 107
rect -885 79 -851 107
rect -823 79 -789 107
rect -761 79 -727 107
rect -699 79 -665 107
rect -637 79 -603 107
rect -575 79 -541 107
rect -513 79 -479 107
rect -451 79 -417 107
rect -389 79 -355 107
rect -327 79 -293 107
rect -265 79 -231 107
rect -203 79 -169 107
rect -141 79 -107 107
rect -79 79 -45 107
rect -17 79 17 107
rect 45 79 79 107
rect 107 79 141 107
rect 169 79 203 107
rect 231 79 265 107
rect 293 79 327 107
rect 355 79 389 107
rect 417 79 451 107
rect 479 79 513 107
rect 541 79 575 107
rect 603 79 637 107
rect 665 79 699 107
rect 727 79 761 107
rect 789 79 823 107
rect 851 79 885 107
rect 913 79 947 107
rect 975 79 1009 107
rect 1037 79 1071 107
rect 1099 79 1133 107
rect 1161 79 1195 107
rect 1223 79 1257 107
rect 1285 79 1319 107
rect 1347 79 1381 107
rect 1409 79 1443 107
rect 1471 79 1505 107
rect 1533 79 1567 107
rect 1595 79 1629 107
rect 1657 79 1691 107
rect 1719 79 1753 107
rect 1781 79 1815 107
rect 1843 79 1877 107
rect 1905 79 1939 107
rect 1967 79 2001 107
rect 2029 79 2063 107
rect 2091 79 2125 107
rect 2153 79 2187 107
rect 2215 79 2249 107
rect 2277 79 2311 107
rect 2339 79 2373 107
rect 2401 79 2435 107
rect 2463 79 2497 107
rect 2525 79 2559 107
rect 2587 79 2621 107
rect 2649 79 2683 107
rect 2711 79 2745 107
rect 2773 79 2807 107
rect 2835 79 2869 107
rect 2897 79 2931 107
rect 2959 79 2993 107
rect 3021 79 3055 107
rect 3083 79 3117 107
rect 3145 79 3179 107
rect 3207 79 3241 107
rect 3269 79 3303 107
rect 3331 79 3336 107
rect -3336 45 3336 79
rect -3336 17 -3331 45
rect -3303 17 -3269 45
rect -3241 17 -3207 45
rect -3179 17 -3145 45
rect -3117 17 -3083 45
rect -3055 17 -3021 45
rect -2993 17 -2959 45
rect -2931 17 -2897 45
rect -2869 17 -2835 45
rect -2807 17 -2773 45
rect -2745 17 -2711 45
rect -2683 17 -2649 45
rect -2621 17 -2587 45
rect -2559 17 -2525 45
rect -2497 17 -2463 45
rect -2435 17 -2401 45
rect -2373 17 -2339 45
rect -2311 17 -2277 45
rect -2249 17 -2215 45
rect -2187 17 -2153 45
rect -2125 17 -2091 45
rect -2063 17 -2029 45
rect -2001 17 -1967 45
rect -1939 17 -1905 45
rect -1877 17 -1843 45
rect -1815 17 -1781 45
rect -1753 17 -1719 45
rect -1691 17 -1657 45
rect -1629 17 -1595 45
rect -1567 17 -1533 45
rect -1505 17 -1471 45
rect -1443 17 -1409 45
rect -1381 17 -1347 45
rect -1319 17 -1285 45
rect -1257 17 -1223 45
rect -1195 17 -1161 45
rect -1133 17 -1099 45
rect -1071 17 -1037 45
rect -1009 17 -975 45
rect -947 17 -913 45
rect -885 17 -851 45
rect -823 17 -789 45
rect -761 17 -727 45
rect -699 17 -665 45
rect -637 17 -603 45
rect -575 17 -541 45
rect -513 17 -479 45
rect -451 17 -417 45
rect -389 17 -355 45
rect -327 17 -293 45
rect -265 17 -231 45
rect -203 17 -169 45
rect -141 17 -107 45
rect -79 17 -45 45
rect -17 17 17 45
rect 45 17 79 45
rect 107 17 141 45
rect 169 17 203 45
rect 231 17 265 45
rect 293 17 327 45
rect 355 17 389 45
rect 417 17 451 45
rect 479 17 513 45
rect 541 17 575 45
rect 603 17 637 45
rect 665 17 699 45
rect 727 17 761 45
rect 789 17 823 45
rect 851 17 885 45
rect 913 17 947 45
rect 975 17 1009 45
rect 1037 17 1071 45
rect 1099 17 1133 45
rect 1161 17 1195 45
rect 1223 17 1257 45
rect 1285 17 1319 45
rect 1347 17 1381 45
rect 1409 17 1443 45
rect 1471 17 1505 45
rect 1533 17 1567 45
rect 1595 17 1629 45
rect 1657 17 1691 45
rect 1719 17 1753 45
rect 1781 17 1815 45
rect 1843 17 1877 45
rect 1905 17 1939 45
rect 1967 17 2001 45
rect 2029 17 2063 45
rect 2091 17 2125 45
rect 2153 17 2187 45
rect 2215 17 2249 45
rect 2277 17 2311 45
rect 2339 17 2373 45
rect 2401 17 2435 45
rect 2463 17 2497 45
rect 2525 17 2559 45
rect 2587 17 2621 45
rect 2649 17 2683 45
rect 2711 17 2745 45
rect 2773 17 2807 45
rect 2835 17 2869 45
rect 2897 17 2931 45
rect 2959 17 2993 45
rect 3021 17 3055 45
rect 3083 17 3117 45
rect 3145 17 3179 45
rect 3207 17 3241 45
rect 3269 17 3303 45
rect 3331 17 3336 45
rect -3336 -17 3336 17
rect -3336 -45 -3331 -17
rect -3303 -45 -3269 -17
rect -3241 -45 -3207 -17
rect -3179 -45 -3145 -17
rect -3117 -45 -3083 -17
rect -3055 -45 -3021 -17
rect -2993 -45 -2959 -17
rect -2931 -45 -2897 -17
rect -2869 -45 -2835 -17
rect -2807 -45 -2773 -17
rect -2745 -45 -2711 -17
rect -2683 -45 -2649 -17
rect -2621 -45 -2587 -17
rect -2559 -45 -2525 -17
rect -2497 -45 -2463 -17
rect -2435 -45 -2401 -17
rect -2373 -45 -2339 -17
rect -2311 -45 -2277 -17
rect -2249 -45 -2215 -17
rect -2187 -45 -2153 -17
rect -2125 -45 -2091 -17
rect -2063 -45 -2029 -17
rect -2001 -45 -1967 -17
rect -1939 -45 -1905 -17
rect -1877 -45 -1843 -17
rect -1815 -45 -1781 -17
rect -1753 -45 -1719 -17
rect -1691 -45 -1657 -17
rect -1629 -45 -1595 -17
rect -1567 -45 -1533 -17
rect -1505 -45 -1471 -17
rect -1443 -45 -1409 -17
rect -1381 -45 -1347 -17
rect -1319 -45 -1285 -17
rect -1257 -45 -1223 -17
rect -1195 -45 -1161 -17
rect -1133 -45 -1099 -17
rect -1071 -45 -1037 -17
rect -1009 -45 -975 -17
rect -947 -45 -913 -17
rect -885 -45 -851 -17
rect -823 -45 -789 -17
rect -761 -45 -727 -17
rect -699 -45 -665 -17
rect -637 -45 -603 -17
rect -575 -45 -541 -17
rect -513 -45 -479 -17
rect -451 -45 -417 -17
rect -389 -45 -355 -17
rect -327 -45 -293 -17
rect -265 -45 -231 -17
rect -203 -45 -169 -17
rect -141 -45 -107 -17
rect -79 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 79 -17
rect 107 -45 141 -17
rect 169 -45 203 -17
rect 231 -45 265 -17
rect 293 -45 327 -17
rect 355 -45 389 -17
rect 417 -45 451 -17
rect 479 -45 513 -17
rect 541 -45 575 -17
rect 603 -45 637 -17
rect 665 -45 699 -17
rect 727 -45 761 -17
rect 789 -45 823 -17
rect 851 -45 885 -17
rect 913 -45 947 -17
rect 975 -45 1009 -17
rect 1037 -45 1071 -17
rect 1099 -45 1133 -17
rect 1161 -45 1195 -17
rect 1223 -45 1257 -17
rect 1285 -45 1319 -17
rect 1347 -45 1381 -17
rect 1409 -45 1443 -17
rect 1471 -45 1505 -17
rect 1533 -45 1567 -17
rect 1595 -45 1629 -17
rect 1657 -45 1691 -17
rect 1719 -45 1753 -17
rect 1781 -45 1815 -17
rect 1843 -45 1877 -17
rect 1905 -45 1939 -17
rect 1967 -45 2001 -17
rect 2029 -45 2063 -17
rect 2091 -45 2125 -17
rect 2153 -45 2187 -17
rect 2215 -45 2249 -17
rect 2277 -45 2311 -17
rect 2339 -45 2373 -17
rect 2401 -45 2435 -17
rect 2463 -45 2497 -17
rect 2525 -45 2559 -17
rect 2587 -45 2621 -17
rect 2649 -45 2683 -17
rect 2711 -45 2745 -17
rect 2773 -45 2807 -17
rect 2835 -45 2869 -17
rect 2897 -45 2931 -17
rect 2959 -45 2993 -17
rect 3021 -45 3055 -17
rect 3083 -45 3117 -17
rect 3145 -45 3179 -17
rect 3207 -45 3241 -17
rect 3269 -45 3303 -17
rect 3331 -45 3336 -17
rect -3336 -79 3336 -45
rect -3336 -107 -3331 -79
rect -3303 -107 -3269 -79
rect -3241 -107 -3207 -79
rect -3179 -107 -3145 -79
rect -3117 -107 -3083 -79
rect -3055 -107 -3021 -79
rect -2993 -107 -2959 -79
rect -2931 -107 -2897 -79
rect -2869 -107 -2835 -79
rect -2807 -107 -2773 -79
rect -2745 -107 -2711 -79
rect -2683 -107 -2649 -79
rect -2621 -107 -2587 -79
rect -2559 -107 -2525 -79
rect -2497 -107 -2463 -79
rect -2435 -107 -2401 -79
rect -2373 -107 -2339 -79
rect -2311 -107 -2277 -79
rect -2249 -107 -2215 -79
rect -2187 -107 -2153 -79
rect -2125 -107 -2091 -79
rect -2063 -107 -2029 -79
rect -2001 -107 -1967 -79
rect -1939 -107 -1905 -79
rect -1877 -107 -1843 -79
rect -1815 -107 -1781 -79
rect -1753 -107 -1719 -79
rect -1691 -107 -1657 -79
rect -1629 -107 -1595 -79
rect -1567 -107 -1533 -79
rect -1505 -107 -1471 -79
rect -1443 -107 -1409 -79
rect -1381 -107 -1347 -79
rect -1319 -107 -1285 -79
rect -1257 -107 -1223 -79
rect -1195 -107 -1161 -79
rect -1133 -107 -1099 -79
rect -1071 -107 -1037 -79
rect -1009 -107 -975 -79
rect -947 -107 -913 -79
rect -885 -107 -851 -79
rect -823 -107 -789 -79
rect -761 -107 -727 -79
rect -699 -107 -665 -79
rect -637 -107 -603 -79
rect -575 -107 -541 -79
rect -513 -107 -479 -79
rect -451 -107 -417 -79
rect -389 -107 -355 -79
rect -327 -107 -293 -79
rect -265 -107 -231 -79
rect -203 -107 -169 -79
rect -141 -107 -107 -79
rect -79 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 79 -79
rect 107 -107 141 -79
rect 169 -107 203 -79
rect 231 -107 265 -79
rect 293 -107 327 -79
rect 355 -107 389 -79
rect 417 -107 451 -79
rect 479 -107 513 -79
rect 541 -107 575 -79
rect 603 -107 637 -79
rect 665 -107 699 -79
rect 727 -107 761 -79
rect 789 -107 823 -79
rect 851 -107 885 -79
rect 913 -107 947 -79
rect 975 -107 1009 -79
rect 1037 -107 1071 -79
rect 1099 -107 1133 -79
rect 1161 -107 1195 -79
rect 1223 -107 1257 -79
rect 1285 -107 1319 -79
rect 1347 -107 1381 -79
rect 1409 -107 1443 -79
rect 1471 -107 1505 -79
rect 1533 -107 1567 -79
rect 1595 -107 1629 -79
rect 1657 -107 1691 -79
rect 1719 -107 1753 -79
rect 1781 -107 1815 -79
rect 1843 -107 1877 -79
rect 1905 -107 1939 -79
rect 1967 -107 2001 -79
rect 2029 -107 2063 -79
rect 2091 -107 2125 -79
rect 2153 -107 2187 -79
rect 2215 -107 2249 -79
rect 2277 -107 2311 -79
rect 2339 -107 2373 -79
rect 2401 -107 2435 -79
rect 2463 -107 2497 -79
rect 2525 -107 2559 -79
rect 2587 -107 2621 -79
rect 2649 -107 2683 -79
rect 2711 -107 2745 -79
rect 2773 -107 2807 -79
rect 2835 -107 2869 -79
rect 2897 -107 2931 -79
rect 2959 -107 2993 -79
rect 3021 -107 3055 -79
rect 3083 -107 3117 -79
rect 3145 -107 3179 -79
rect 3207 -107 3241 -79
rect 3269 -107 3303 -79
rect 3331 -107 3336 -79
rect -3336 -112 3336 -107
<< end >>
