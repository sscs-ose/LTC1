magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1090 -1729 1090 1729
<< metal2 >>
rect -90 724 90 729
rect -90 696 -85 724
rect -57 696 -14 724
rect 14 696 57 724
rect 85 696 90 724
rect -90 653 90 696
rect -90 625 -85 653
rect -57 625 -14 653
rect 14 625 57 653
rect 85 625 90 653
rect -90 582 90 625
rect -90 554 -85 582
rect -57 554 -14 582
rect 14 554 57 582
rect 85 554 90 582
rect -90 511 90 554
rect -90 483 -85 511
rect -57 483 -14 511
rect 14 483 57 511
rect 85 483 90 511
rect -90 440 90 483
rect -90 412 -85 440
rect -57 412 -14 440
rect 14 412 57 440
rect 85 412 90 440
rect -90 369 90 412
rect -90 341 -85 369
rect -57 341 -14 369
rect 14 341 57 369
rect 85 341 90 369
rect -90 298 90 341
rect -90 270 -85 298
rect -57 270 -14 298
rect 14 270 57 298
rect 85 270 90 298
rect -90 227 90 270
rect -90 199 -85 227
rect -57 199 -14 227
rect 14 199 57 227
rect 85 199 90 227
rect -90 156 90 199
rect -90 128 -85 156
rect -57 128 -14 156
rect 14 128 57 156
rect 85 128 90 156
rect -90 85 90 128
rect -90 57 -85 85
rect -57 57 -14 85
rect 14 57 57 85
rect 85 57 90 85
rect -90 14 90 57
rect -90 -14 -85 14
rect -57 -14 -14 14
rect 14 -14 57 14
rect 85 -14 90 14
rect -90 -57 90 -14
rect -90 -85 -85 -57
rect -57 -85 -14 -57
rect 14 -85 57 -57
rect 85 -85 90 -57
rect -90 -128 90 -85
rect -90 -156 -85 -128
rect -57 -156 -14 -128
rect 14 -156 57 -128
rect 85 -156 90 -128
rect -90 -199 90 -156
rect -90 -227 -85 -199
rect -57 -227 -14 -199
rect 14 -227 57 -199
rect 85 -227 90 -199
rect -90 -270 90 -227
rect -90 -298 -85 -270
rect -57 -298 -14 -270
rect 14 -298 57 -270
rect 85 -298 90 -270
rect -90 -341 90 -298
rect -90 -369 -85 -341
rect -57 -369 -14 -341
rect 14 -369 57 -341
rect 85 -369 90 -341
rect -90 -412 90 -369
rect -90 -440 -85 -412
rect -57 -440 -14 -412
rect 14 -440 57 -412
rect 85 -440 90 -412
rect -90 -483 90 -440
rect -90 -511 -85 -483
rect -57 -511 -14 -483
rect 14 -511 57 -483
rect 85 -511 90 -483
rect -90 -554 90 -511
rect -90 -582 -85 -554
rect -57 -582 -14 -554
rect 14 -582 57 -554
rect 85 -582 90 -554
rect -90 -625 90 -582
rect -90 -653 -85 -625
rect -57 -653 -14 -625
rect 14 -653 57 -625
rect 85 -653 90 -625
rect -90 -696 90 -653
rect -90 -724 -85 -696
rect -57 -724 -14 -696
rect 14 -724 57 -696
rect 85 -724 90 -696
rect -90 -729 90 -724
<< via2 >>
rect -85 696 -57 724
rect -14 696 14 724
rect 57 696 85 724
rect -85 625 -57 653
rect -14 625 14 653
rect 57 625 85 653
rect -85 554 -57 582
rect -14 554 14 582
rect 57 554 85 582
rect -85 483 -57 511
rect -14 483 14 511
rect 57 483 85 511
rect -85 412 -57 440
rect -14 412 14 440
rect 57 412 85 440
rect -85 341 -57 369
rect -14 341 14 369
rect 57 341 85 369
rect -85 270 -57 298
rect -14 270 14 298
rect 57 270 85 298
rect -85 199 -57 227
rect -14 199 14 227
rect 57 199 85 227
rect -85 128 -57 156
rect -14 128 14 156
rect 57 128 85 156
rect -85 57 -57 85
rect -14 57 14 85
rect 57 57 85 85
rect -85 -14 -57 14
rect -14 -14 14 14
rect 57 -14 85 14
rect -85 -85 -57 -57
rect -14 -85 14 -57
rect 57 -85 85 -57
rect -85 -156 -57 -128
rect -14 -156 14 -128
rect 57 -156 85 -128
rect -85 -227 -57 -199
rect -14 -227 14 -199
rect 57 -227 85 -199
rect -85 -298 -57 -270
rect -14 -298 14 -270
rect 57 -298 85 -270
rect -85 -369 -57 -341
rect -14 -369 14 -341
rect 57 -369 85 -341
rect -85 -440 -57 -412
rect -14 -440 14 -412
rect 57 -440 85 -412
rect -85 -511 -57 -483
rect -14 -511 14 -483
rect 57 -511 85 -483
rect -85 -582 -57 -554
rect -14 -582 14 -554
rect 57 -582 85 -554
rect -85 -653 -57 -625
rect -14 -653 14 -625
rect 57 -653 85 -625
rect -85 -724 -57 -696
rect -14 -724 14 -696
rect 57 -724 85 -696
<< metal3 >>
rect -90 724 90 729
rect -90 696 -85 724
rect -57 696 -14 724
rect 14 696 57 724
rect 85 696 90 724
rect -90 653 90 696
rect -90 625 -85 653
rect -57 625 -14 653
rect 14 625 57 653
rect 85 625 90 653
rect -90 582 90 625
rect -90 554 -85 582
rect -57 554 -14 582
rect 14 554 57 582
rect 85 554 90 582
rect -90 511 90 554
rect -90 483 -85 511
rect -57 483 -14 511
rect 14 483 57 511
rect 85 483 90 511
rect -90 440 90 483
rect -90 412 -85 440
rect -57 412 -14 440
rect 14 412 57 440
rect 85 412 90 440
rect -90 369 90 412
rect -90 341 -85 369
rect -57 341 -14 369
rect 14 341 57 369
rect 85 341 90 369
rect -90 298 90 341
rect -90 270 -85 298
rect -57 270 -14 298
rect 14 270 57 298
rect 85 270 90 298
rect -90 227 90 270
rect -90 199 -85 227
rect -57 199 -14 227
rect 14 199 57 227
rect 85 199 90 227
rect -90 156 90 199
rect -90 128 -85 156
rect -57 128 -14 156
rect 14 128 57 156
rect 85 128 90 156
rect -90 85 90 128
rect -90 57 -85 85
rect -57 57 -14 85
rect 14 57 57 85
rect 85 57 90 85
rect -90 14 90 57
rect -90 -14 -85 14
rect -57 -14 -14 14
rect 14 -14 57 14
rect 85 -14 90 14
rect -90 -57 90 -14
rect -90 -85 -85 -57
rect -57 -85 -14 -57
rect 14 -85 57 -57
rect 85 -85 90 -57
rect -90 -128 90 -85
rect -90 -156 -85 -128
rect -57 -156 -14 -128
rect 14 -156 57 -128
rect 85 -156 90 -128
rect -90 -199 90 -156
rect -90 -227 -85 -199
rect -57 -227 -14 -199
rect 14 -227 57 -199
rect 85 -227 90 -199
rect -90 -270 90 -227
rect -90 -298 -85 -270
rect -57 -298 -14 -270
rect 14 -298 57 -270
rect 85 -298 90 -270
rect -90 -341 90 -298
rect -90 -369 -85 -341
rect -57 -369 -14 -341
rect 14 -369 57 -341
rect 85 -369 90 -341
rect -90 -412 90 -369
rect -90 -440 -85 -412
rect -57 -440 -14 -412
rect 14 -440 57 -412
rect 85 -440 90 -412
rect -90 -483 90 -440
rect -90 -511 -85 -483
rect -57 -511 -14 -483
rect 14 -511 57 -483
rect 85 -511 90 -483
rect -90 -554 90 -511
rect -90 -582 -85 -554
rect -57 -582 -14 -554
rect 14 -582 57 -554
rect 85 -582 90 -554
rect -90 -625 90 -582
rect -90 -653 -85 -625
rect -57 -653 -14 -625
rect 14 -653 57 -625
rect 85 -653 90 -625
rect -90 -696 90 -653
rect -90 -724 -85 -696
rect -57 -724 -14 -696
rect 14 -724 57 -696
rect 85 -724 90 -696
rect -90 -729 90 -724
<< end >>
