magic
tech gf180mcuC
magscale 1 10
timestamp 1692078773
<< nwell >>
rect 153 589 557 1135
rect 1195 617 2079 1135
rect 3578 617 4462 1135
rect 153 -1121 557 -167
rect 1195 -1403 2079 -505
rect 3578 -885 4462 -505
rect 2913 -1023 4946 -885
rect 2913 -1476 4085 -1023
rect 4222 -1408 4946 -1023
<< pwell >>
rect 215 279 495 515
rect 777 307 2497 543
rect 3160 307 4880 543
rect 215 -93 495 143
rect 777 -431 2497 -195
rect 3160 -431 4880 -195
rect 215 -1431 495 -1195
rect 777 -1713 2497 -1477
rect 3135 -1786 3735 -1550
rect 4124 -1718 4884 -1482
rect 4902 -1718 5182 -1482
<< nmos >>
rect 327 347 383 447
rect 889 375 945 475
rect 1049 375 1105 475
rect 1209 375 1265 475
rect 1369 375 1425 475
rect 1529 375 1585 475
rect 1689 375 1745 475
rect 1849 375 1905 475
rect 2009 375 2065 475
rect 2169 375 2225 475
rect 2329 375 2385 475
rect 3272 375 3328 475
rect 3432 375 3488 475
rect 3592 375 3648 475
rect 3752 375 3808 475
rect 3912 375 3968 475
rect 4072 375 4128 475
rect 4232 375 4288 475
rect 4392 375 4448 475
rect 4552 375 4608 475
rect 4712 375 4768 475
rect 327 -25 383 75
rect 889 -363 945 -263
rect 1049 -363 1105 -263
rect 1209 -363 1265 -263
rect 1369 -363 1425 -263
rect 1529 -363 1585 -263
rect 1689 -363 1745 -263
rect 1849 -363 1905 -263
rect 2009 -363 2065 -263
rect 2169 -363 2225 -263
rect 2329 -363 2385 -263
rect 3272 -363 3328 -263
rect 3432 -363 3488 -263
rect 3592 -363 3648 -263
rect 3752 -363 3808 -263
rect 3912 -363 3968 -263
rect 4072 -363 4128 -263
rect 4232 -363 4288 -263
rect 4392 -363 4448 -263
rect 4552 -363 4608 -263
rect 4712 -363 4768 -263
rect 327 -1363 383 -1263
rect 889 -1645 945 -1545
rect 1049 -1645 1105 -1545
rect 1209 -1645 1265 -1545
rect 1369 -1645 1425 -1545
rect 1529 -1645 1585 -1545
rect 1689 -1645 1745 -1545
rect 1849 -1645 1905 -1545
rect 2009 -1645 2065 -1545
rect 2169 -1645 2225 -1545
rect 2329 -1645 2385 -1545
rect 3247 -1718 3303 -1618
rect 3407 -1718 3463 -1618
rect 3567 -1718 3623 -1618
rect 4236 -1650 4292 -1550
rect 4396 -1650 4452 -1550
rect 4556 -1650 4612 -1550
rect 4716 -1650 4772 -1550
rect 5014 -1650 5070 -1550
<< pmos >>
rect 327 719 383 919
rect 1369 747 1425 947
rect 1529 747 1585 947
rect 1689 747 1745 947
rect 1849 747 1905 947
rect 3752 747 3808 947
rect 3912 747 3968 947
rect 4072 747 4128 947
rect 4232 747 4288 947
rect 327 -497 383 -297
rect 327 -991 383 -791
rect 1369 -835 1425 -635
rect 1529 -835 1585 -635
rect 1689 -835 1745 -635
rect 1849 -835 1905 -635
rect 3752 -835 3808 -635
rect 3912 -835 3968 -635
rect 4072 -835 4128 -635
rect 4232 -835 4288 -635
rect 1369 -1273 1425 -1073
rect 1529 -1273 1585 -1073
rect 1689 -1273 1745 -1073
rect 1849 -1273 1905 -1073
rect 3087 -1346 3143 -1146
rect 3247 -1346 3303 -1146
rect 3407 -1346 3463 -1146
rect 3567 -1346 3623 -1146
rect 3855 -1346 3911 -1146
rect 4396 -1278 4452 -1078
rect 4556 -1278 4612 -1078
rect 4716 -1278 4772 -1078
<< ndiff >>
rect 801 462 889 475
rect 239 434 327 447
rect 239 360 252 434
rect 298 360 327 434
rect 239 347 327 360
rect 383 434 471 447
rect 383 360 412 434
rect 458 360 471 434
rect 801 388 814 462
rect 860 388 889 462
rect 801 375 889 388
rect 945 462 1049 475
rect 945 388 974 462
rect 1020 388 1049 462
rect 945 375 1049 388
rect 1105 462 1209 475
rect 1105 388 1134 462
rect 1180 388 1209 462
rect 1105 375 1209 388
rect 1265 462 1369 475
rect 1265 388 1294 462
rect 1340 388 1369 462
rect 1265 375 1369 388
rect 1425 462 1529 475
rect 1425 388 1454 462
rect 1500 388 1529 462
rect 1425 375 1529 388
rect 1585 462 1689 475
rect 1585 388 1614 462
rect 1660 388 1689 462
rect 1585 375 1689 388
rect 1745 462 1849 475
rect 1745 388 1774 462
rect 1820 388 1849 462
rect 1745 375 1849 388
rect 1905 462 2009 475
rect 1905 388 1934 462
rect 1980 388 2009 462
rect 1905 375 2009 388
rect 2065 462 2169 475
rect 2065 388 2094 462
rect 2140 388 2169 462
rect 2065 375 2169 388
rect 2225 462 2329 475
rect 2225 388 2254 462
rect 2300 388 2329 462
rect 2225 375 2329 388
rect 2385 462 2473 475
rect 2385 388 2414 462
rect 2460 388 2473 462
rect 2385 375 2473 388
rect 3184 462 3272 475
rect 3184 388 3197 462
rect 3243 388 3272 462
rect 3184 375 3272 388
rect 3328 462 3432 475
rect 3328 388 3357 462
rect 3403 388 3432 462
rect 3328 375 3432 388
rect 3488 462 3592 475
rect 3488 388 3517 462
rect 3563 388 3592 462
rect 3488 375 3592 388
rect 3648 462 3752 475
rect 3648 388 3677 462
rect 3723 388 3752 462
rect 3648 375 3752 388
rect 3808 462 3912 475
rect 3808 388 3837 462
rect 3883 388 3912 462
rect 3808 375 3912 388
rect 3968 462 4072 475
rect 3968 388 3997 462
rect 4043 388 4072 462
rect 3968 375 4072 388
rect 4128 462 4232 475
rect 4128 388 4157 462
rect 4203 388 4232 462
rect 4128 375 4232 388
rect 4288 462 4392 475
rect 4288 388 4317 462
rect 4363 388 4392 462
rect 4288 375 4392 388
rect 4448 462 4552 475
rect 4448 388 4477 462
rect 4523 388 4552 462
rect 4448 375 4552 388
rect 4608 462 4712 475
rect 4608 388 4637 462
rect 4683 388 4712 462
rect 4608 375 4712 388
rect 4768 462 4856 475
rect 4768 388 4797 462
rect 4843 388 4856 462
rect 4768 375 4856 388
rect 383 347 471 360
rect 239 62 327 75
rect 239 -12 252 62
rect 298 -12 327 62
rect 239 -25 327 -12
rect 383 62 471 75
rect 383 -12 412 62
rect 458 -12 471 62
rect 383 -25 471 -12
rect 801 -276 889 -263
rect 801 -350 814 -276
rect 860 -350 889 -276
rect 801 -363 889 -350
rect 945 -276 1049 -263
rect 945 -350 974 -276
rect 1020 -350 1049 -276
rect 945 -363 1049 -350
rect 1105 -276 1209 -263
rect 1105 -350 1134 -276
rect 1180 -350 1209 -276
rect 1105 -363 1209 -350
rect 1265 -276 1369 -263
rect 1265 -350 1294 -276
rect 1340 -350 1369 -276
rect 1265 -363 1369 -350
rect 1425 -276 1529 -263
rect 1425 -350 1454 -276
rect 1500 -350 1529 -276
rect 1425 -363 1529 -350
rect 1585 -276 1689 -263
rect 1585 -350 1614 -276
rect 1660 -350 1689 -276
rect 1585 -363 1689 -350
rect 1745 -276 1849 -263
rect 1745 -350 1774 -276
rect 1820 -350 1849 -276
rect 1745 -363 1849 -350
rect 1905 -276 2009 -263
rect 1905 -350 1934 -276
rect 1980 -350 2009 -276
rect 1905 -363 2009 -350
rect 2065 -276 2169 -263
rect 2065 -350 2094 -276
rect 2140 -350 2169 -276
rect 2065 -363 2169 -350
rect 2225 -276 2329 -263
rect 2225 -350 2254 -276
rect 2300 -350 2329 -276
rect 2225 -363 2329 -350
rect 2385 -276 2473 -263
rect 2385 -350 2414 -276
rect 2460 -350 2473 -276
rect 2385 -363 2473 -350
rect 3184 -276 3272 -263
rect 3184 -350 3197 -276
rect 3243 -350 3272 -276
rect 3184 -363 3272 -350
rect 3328 -276 3432 -263
rect 3328 -350 3357 -276
rect 3403 -350 3432 -276
rect 3328 -363 3432 -350
rect 3488 -276 3592 -263
rect 3488 -350 3517 -276
rect 3563 -350 3592 -276
rect 3488 -363 3592 -350
rect 3648 -276 3752 -263
rect 3648 -350 3677 -276
rect 3723 -350 3752 -276
rect 3648 -363 3752 -350
rect 3808 -276 3912 -263
rect 3808 -350 3837 -276
rect 3883 -350 3912 -276
rect 3808 -363 3912 -350
rect 3968 -276 4072 -263
rect 3968 -350 3997 -276
rect 4043 -350 4072 -276
rect 3968 -363 4072 -350
rect 4128 -276 4232 -263
rect 4128 -350 4157 -276
rect 4203 -350 4232 -276
rect 4128 -363 4232 -350
rect 4288 -276 4392 -263
rect 4288 -350 4317 -276
rect 4363 -350 4392 -276
rect 4288 -363 4392 -350
rect 4448 -276 4552 -263
rect 4448 -350 4477 -276
rect 4523 -350 4552 -276
rect 4448 -363 4552 -350
rect 4608 -276 4712 -263
rect 4608 -350 4637 -276
rect 4683 -350 4712 -276
rect 4608 -363 4712 -350
rect 4768 -276 4856 -263
rect 4768 -350 4797 -276
rect 4843 -350 4856 -276
rect 4768 -363 4856 -350
rect 239 -1276 327 -1263
rect 239 -1350 252 -1276
rect 298 -1350 327 -1276
rect 239 -1363 327 -1350
rect 383 -1276 471 -1263
rect 383 -1350 412 -1276
rect 458 -1350 471 -1276
rect 383 -1363 471 -1350
rect 801 -1558 889 -1545
rect 801 -1632 814 -1558
rect 860 -1632 889 -1558
rect 801 -1645 889 -1632
rect 945 -1558 1049 -1545
rect 945 -1632 974 -1558
rect 1020 -1632 1049 -1558
rect 945 -1645 1049 -1632
rect 1105 -1558 1209 -1545
rect 1105 -1632 1134 -1558
rect 1180 -1632 1209 -1558
rect 1105 -1645 1209 -1632
rect 1265 -1558 1369 -1545
rect 1265 -1632 1294 -1558
rect 1340 -1632 1369 -1558
rect 1265 -1645 1369 -1632
rect 1425 -1558 1529 -1545
rect 1425 -1632 1454 -1558
rect 1500 -1632 1529 -1558
rect 1425 -1645 1529 -1632
rect 1585 -1558 1689 -1545
rect 1585 -1632 1614 -1558
rect 1660 -1632 1689 -1558
rect 1585 -1645 1689 -1632
rect 1745 -1558 1849 -1545
rect 1745 -1632 1774 -1558
rect 1820 -1632 1849 -1558
rect 1745 -1645 1849 -1632
rect 1905 -1558 2009 -1545
rect 1905 -1632 1934 -1558
rect 1980 -1632 2009 -1558
rect 1905 -1645 2009 -1632
rect 2065 -1558 2169 -1545
rect 2065 -1632 2094 -1558
rect 2140 -1632 2169 -1558
rect 2065 -1645 2169 -1632
rect 2225 -1558 2329 -1545
rect 2225 -1632 2254 -1558
rect 2300 -1632 2329 -1558
rect 2225 -1645 2329 -1632
rect 2385 -1558 2473 -1545
rect 2385 -1632 2414 -1558
rect 2460 -1632 2473 -1558
rect 4148 -1563 4236 -1550
rect 2385 -1645 2473 -1632
rect 3159 -1631 3247 -1618
rect 3159 -1705 3172 -1631
rect 3218 -1705 3247 -1631
rect 3159 -1718 3247 -1705
rect 3303 -1631 3407 -1618
rect 3303 -1705 3332 -1631
rect 3378 -1705 3407 -1631
rect 3303 -1718 3407 -1705
rect 3463 -1631 3567 -1618
rect 3463 -1705 3492 -1631
rect 3538 -1705 3567 -1631
rect 3463 -1718 3567 -1705
rect 3623 -1631 3711 -1618
rect 3623 -1705 3652 -1631
rect 3698 -1705 3711 -1631
rect 4148 -1637 4161 -1563
rect 4207 -1637 4236 -1563
rect 4148 -1650 4236 -1637
rect 4292 -1563 4396 -1550
rect 4292 -1637 4321 -1563
rect 4367 -1637 4396 -1563
rect 4292 -1650 4396 -1637
rect 4452 -1563 4556 -1550
rect 4452 -1637 4481 -1563
rect 4527 -1637 4556 -1563
rect 4452 -1650 4556 -1637
rect 4612 -1563 4716 -1550
rect 4612 -1637 4641 -1563
rect 4687 -1637 4716 -1563
rect 4612 -1650 4716 -1637
rect 4772 -1563 4860 -1550
rect 4772 -1637 4801 -1563
rect 4847 -1637 4860 -1563
rect 4772 -1650 4860 -1637
rect 4926 -1563 5014 -1550
rect 4926 -1637 4939 -1563
rect 4985 -1637 5014 -1563
rect 4926 -1650 5014 -1637
rect 5070 -1563 5158 -1550
rect 5070 -1637 5099 -1563
rect 5145 -1637 5158 -1563
rect 5070 -1650 5158 -1637
rect 3623 -1718 3711 -1705
<< pdiff >>
rect 1281 934 1369 947
rect 239 906 327 919
rect 239 732 252 906
rect 298 732 327 906
rect 239 719 327 732
rect 383 906 471 919
rect 383 732 412 906
rect 458 732 471 906
rect 1281 760 1294 934
rect 1340 760 1369 934
rect 1281 747 1369 760
rect 1425 934 1529 947
rect 1425 760 1454 934
rect 1500 760 1529 934
rect 1425 747 1529 760
rect 1585 934 1689 947
rect 1585 760 1614 934
rect 1660 760 1689 934
rect 1585 747 1689 760
rect 1745 934 1849 947
rect 1745 760 1774 934
rect 1820 760 1849 934
rect 1745 747 1849 760
rect 1905 934 1993 947
rect 1905 760 1934 934
rect 1980 760 1993 934
rect 1905 747 1993 760
rect 3664 934 3752 947
rect 3664 760 3677 934
rect 3723 760 3752 934
rect 3664 747 3752 760
rect 3808 934 3912 947
rect 3808 760 3837 934
rect 3883 760 3912 934
rect 3808 747 3912 760
rect 3968 934 4072 947
rect 3968 760 3997 934
rect 4043 760 4072 934
rect 3968 747 4072 760
rect 4128 934 4232 947
rect 4128 760 4157 934
rect 4203 760 4232 934
rect 4128 747 4232 760
rect 4288 934 4376 947
rect 4288 760 4317 934
rect 4363 760 4376 934
rect 4288 747 4376 760
rect 383 719 471 732
rect 239 -310 327 -297
rect 239 -484 252 -310
rect 298 -484 327 -310
rect 239 -497 327 -484
rect 383 -310 471 -297
rect 383 -484 412 -310
rect 458 -484 471 -310
rect 383 -497 471 -484
rect 1281 -648 1369 -635
rect 239 -804 327 -791
rect 239 -978 252 -804
rect 298 -978 327 -804
rect 239 -991 327 -978
rect 383 -804 471 -791
rect 383 -978 412 -804
rect 458 -978 471 -804
rect 1281 -822 1294 -648
rect 1340 -822 1369 -648
rect 1281 -835 1369 -822
rect 1425 -648 1529 -635
rect 1425 -822 1454 -648
rect 1500 -822 1529 -648
rect 1425 -835 1529 -822
rect 1585 -648 1689 -635
rect 1585 -822 1614 -648
rect 1660 -822 1689 -648
rect 1585 -835 1689 -822
rect 1745 -648 1849 -635
rect 1745 -822 1774 -648
rect 1820 -822 1849 -648
rect 1745 -835 1849 -822
rect 1905 -648 1993 -635
rect 1905 -822 1934 -648
rect 1980 -822 1993 -648
rect 1905 -835 1993 -822
rect 3664 -648 3752 -635
rect 3664 -822 3677 -648
rect 3723 -822 3752 -648
rect 3664 -835 3752 -822
rect 3808 -648 3912 -635
rect 3808 -822 3837 -648
rect 3883 -822 3912 -648
rect 3808 -835 3912 -822
rect 3968 -648 4072 -635
rect 3968 -822 3997 -648
rect 4043 -822 4072 -648
rect 3968 -835 4072 -822
rect 4128 -648 4232 -635
rect 4128 -822 4157 -648
rect 4203 -822 4232 -648
rect 4128 -835 4232 -822
rect 4288 -648 4376 -635
rect 4288 -822 4317 -648
rect 4363 -822 4376 -648
rect 4288 -835 4376 -822
rect 383 -991 471 -978
rect 1281 -1086 1369 -1073
rect 1281 -1260 1294 -1086
rect 1340 -1260 1369 -1086
rect 1281 -1273 1369 -1260
rect 1425 -1086 1529 -1073
rect 1425 -1260 1454 -1086
rect 1500 -1260 1529 -1086
rect 1425 -1273 1529 -1260
rect 1585 -1086 1689 -1073
rect 1585 -1260 1614 -1086
rect 1660 -1260 1689 -1086
rect 1585 -1273 1689 -1260
rect 1745 -1086 1849 -1073
rect 1745 -1260 1774 -1086
rect 1820 -1260 1849 -1086
rect 1745 -1273 1849 -1260
rect 1905 -1086 1993 -1073
rect 1905 -1260 1934 -1086
rect 1980 -1260 1993 -1086
rect 4308 -1091 4396 -1078
rect 1905 -1273 1993 -1260
rect 2999 -1159 3087 -1146
rect 2999 -1333 3012 -1159
rect 3058 -1333 3087 -1159
rect 2999 -1346 3087 -1333
rect 3143 -1159 3247 -1146
rect 3143 -1333 3172 -1159
rect 3218 -1333 3247 -1159
rect 3143 -1346 3247 -1333
rect 3303 -1159 3407 -1146
rect 3303 -1333 3332 -1159
rect 3378 -1333 3407 -1159
rect 3303 -1346 3407 -1333
rect 3463 -1159 3567 -1146
rect 3463 -1333 3492 -1159
rect 3538 -1333 3567 -1159
rect 3463 -1346 3567 -1333
rect 3623 -1159 3711 -1146
rect 3623 -1333 3652 -1159
rect 3698 -1333 3711 -1159
rect 3623 -1346 3711 -1333
rect 3767 -1159 3855 -1146
rect 3767 -1333 3780 -1159
rect 3826 -1333 3855 -1159
rect 3767 -1346 3855 -1333
rect 3911 -1159 3999 -1146
rect 3911 -1333 3940 -1159
rect 3986 -1333 3999 -1159
rect 4308 -1265 4321 -1091
rect 4367 -1265 4396 -1091
rect 4308 -1278 4396 -1265
rect 4452 -1091 4556 -1078
rect 4452 -1265 4481 -1091
rect 4527 -1265 4556 -1091
rect 4452 -1278 4556 -1265
rect 4612 -1091 4716 -1078
rect 4612 -1265 4641 -1091
rect 4687 -1265 4716 -1091
rect 4612 -1278 4716 -1265
rect 4772 -1091 4860 -1078
rect 4772 -1265 4801 -1091
rect 4847 -1265 4860 -1091
rect 4772 -1278 4860 -1265
rect 3911 -1346 3999 -1333
<< ndiffc >>
rect 252 360 298 434
rect 412 360 458 434
rect 814 388 860 462
rect 974 388 1020 462
rect 1134 388 1180 462
rect 1294 388 1340 462
rect 1454 388 1500 462
rect 1614 388 1660 462
rect 1774 388 1820 462
rect 1934 388 1980 462
rect 2094 388 2140 462
rect 2254 388 2300 462
rect 2414 388 2460 462
rect 3197 388 3243 462
rect 3357 388 3403 462
rect 3517 388 3563 462
rect 3677 388 3723 462
rect 3837 388 3883 462
rect 3997 388 4043 462
rect 4157 388 4203 462
rect 4317 388 4363 462
rect 4477 388 4523 462
rect 4637 388 4683 462
rect 4797 388 4843 462
rect 252 -12 298 62
rect 412 -12 458 62
rect 814 -350 860 -276
rect 974 -350 1020 -276
rect 1134 -350 1180 -276
rect 1294 -350 1340 -276
rect 1454 -350 1500 -276
rect 1614 -350 1660 -276
rect 1774 -350 1820 -276
rect 1934 -350 1980 -276
rect 2094 -350 2140 -276
rect 2254 -350 2300 -276
rect 2414 -350 2460 -276
rect 3197 -350 3243 -276
rect 3357 -350 3403 -276
rect 3517 -350 3563 -276
rect 3677 -350 3723 -276
rect 3837 -350 3883 -276
rect 3997 -350 4043 -276
rect 4157 -350 4203 -276
rect 4317 -350 4363 -276
rect 4477 -350 4523 -276
rect 4637 -350 4683 -276
rect 4797 -350 4843 -276
rect 252 -1350 298 -1276
rect 412 -1350 458 -1276
rect 814 -1632 860 -1558
rect 974 -1632 1020 -1558
rect 1134 -1632 1180 -1558
rect 1294 -1632 1340 -1558
rect 1454 -1632 1500 -1558
rect 1614 -1632 1660 -1558
rect 1774 -1632 1820 -1558
rect 1934 -1632 1980 -1558
rect 2094 -1632 2140 -1558
rect 2254 -1632 2300 -1558
rect 2414 -1632 2460 -1558
rect 3172 -1705 3218 -1631
rect 3332 -1705 3378 -1631
rect 3492 -1705 3538 -1631
rect 3652 -1705 3698 -1631
rect 4161 -1637 4207 -1563
rect 4321 -1637 4367 -1563
rect 4481 -1637 4527 -1563
rect 4641 -1637 4687 -1563
rect 4801 -1637 4847 -1563
rect 4939 -1637 4985 -1563
rect 5099 -1637 5145 -1563
<< pdiffc >>
rect 252 732 298 906
rect 412 732 458 906
rect 1294 760 1340 934
rect 1454 760 1500 934
rect 1614 760 1660 934
rect 1774 760 1820 934
rect 1934 760 1980 934
rect 3677 760 3723 934
rect 3837 760 3883 934
rect 3997 760 4043 934
rect 4157 760 4203 934
rect 4317 760 4363 934
rect 252 -484 298 -310
rect 412 -484 458 -310
rect 252 -978 298 -804
rect 412 -978 458 -804
rect 1294 -822 1340 -648
rect 1454 -822 1500 -648
rect 1614 -822 1660 -648
rect 1774 -822 1820 -648
rect 1934 -822 1980 -648
rect 3677 -822 3723 -648
rect 3837 -822 3883 -648
rect 3997 -822 4043 -648
rect 4157 -822 4203 -648
rect 4317 -822 4363 -648
rect 1294 -1260 1340 -1086
rect 1454 -1260 1500 -1086
rect 1614 -1260 1660 -1086
rect 1774 -1260 1820 -1086
rect 1934 -1260 1980 -1086
rect 3012 -1333 3058 -1159
rect 3172 -1333 3218 -1159
rect 3332 -1333 3378 -1159
rect 3492 -1333 3538 -1159
rect 3652 -1333 3698 -1159
rect 3780 -1333 3826 -1159
rect 3940 -1333 3986 -1159
rect 4321 -1265 4367 -1091
rect 4481 -1265 4527 -1091
rect 4641 -1265 4687 -1091
rect 4801 -1265 4847 -1091
<< psubdiff >>
rect 225 234 485 247
rect 225 188 238 234
rect 284 188 332 234
rect 378 188 426 234
rect 472 188 485 234
rect 225 175 485 188
rect 801 79 2472 92
rect 801 33 814 79
rect 860 33 908 79
rect 954 33 1002 79
rect 1048 33 1096 79
rect 1142 33 1190 79
rect 1236 33 1284 79
rect 1330 33 1378 79
rect 1424 33 1472 79
rect 1518 33 1566 79
rect 1612 33 1660 79
rect 1706 33 1754 79
rect 1800 33 1848 79
rect 1894 33 1942 79
rect 1988 33 2036 79
rect 2082 33 2130 79
rect 2176 33 2224 79
rect 2270 33 2318 79
rect 2364 33 2412 79
rect 2458 33 2472 79
rect 801 20 2472 33
rect 3184 79 4855 92
rect 3184 33 3197 79
rect 3243 33 3291 79
rect 3337 33 3385 79
rect 3431 33 3479 79
rect 3525 33 3573 79
rect 3619 33 3667 79
rect 3713 33 3761 79
rect 3807 33 3855 79
rect 3901 33 3949 79
rect 3995 33 4043 79
rect 4089 33 4137 79
rect 4183 33 4231 79
rect 4277 33 4325 79
rect 4371 33 4419 79
rect 4465 33 4513 79
rect 4559 33 4607 79
rect 4653 33 4701 79
rect 4747 33 4795 79
rect 4841 33 4855 79
rect 3184 20 4855 33
rect 225 -1476 485 -1463
rect 225 -1522 238 -1476
rect 284 -1522 332 -1476
rect 378 -1522 426 -1476
rect 472 -1522 485 -1476
rect 225 -1535 485 -1522
rect 801 -1941 2472 -1928
rect 801 -1987 814 -1941
rect 860 -1987 908 -1941
rect 954 -1987 1002 -1941
rect 1048 -1987 1096 -1941
rect 1142 -1987 1190 -1941
rect 1236 -1987 1284 -1941
rect 1330 -1987 1378 -1941
rect 1424 -1987 1472 -1941
rect 1518 -1987 1566 -1941
rect 1612 -1987 1660 -1941
rect 1706 -1987 1754 -1941
rect 1800 -1987 1848 -1941
rect 1894 -1987 1942 -1941
rect 1988 -1987 2036 -1941
rect 2082 -1987 2130 -1941
rect 2176 -1987 2224 -1941
rect 2270 -1987 2318 -1941
rect 2364 -1987 2412 -1941
rect 2458 -1987 2472 -1941
rect 801 -2000 2472 -1987
rect 3164 -1947 3706 -1934
rect 3164 -1993 3177 -1947
rect 3223 -1993 3271 -1947
rect 3317 -1993 3365 -1947
rect 3411 -1993 3459 -1947
rect 3505 -1993 3553 -1947
rect 3599 -1993 3647 -1947
rect 3693 -1993 3706 -1947
rect 3164 -2006 3706 -1993
rect 4152 -1947 5165 -1934
rect 4152 -1993 4165 -1947
rect 4211 -1993 4259 -1947
rect 4305 -1993 4353 -1947
rect 4399 -1993 4447 -1947
rect 4493 -1993 4541 -1947
rect 4587 -1993 4635 -1947
rect 4681 -1993 4729 -1947
rect 4775 -1993 4823 -1947
rect 4869 -1993 4917 -1947
rect 4963 -1993 5011 -1947
rect 5057 -1993 5105 -1947
rect 5151 -1993 5165 -1947
rect 4152 -2006 5165 -1993
<< nsubdiff >>
rect 178 1089 532 1102
rect 178 1043 191 1089
rect 237 1043 285 1089
rect 331 1043 379 1089
rect 425 1043 473 1089
rect 519 1043 532 1089
rect 178 1030 532 1043
rect 1225 1089 2049 1102
rect 1225 1043 1238 1089
rect 1284 1043 1332 1089
rect 1378 1043 1426 1089
rect 1472 1043 1520 1089
rect 1566 1043 1614 1089
rect 1660 1043 1708 1089
rect 1754 1043 1802 1089
rect 1848 1043 1896 1089
rect 1942 1043 1990 1089
rect 2036 1043 2049 1089
rect 1225 1030 2049 1043
rect 3608 1089 4432 1102
rect 3608 1043 3621 1089
rect 3667 1043 3715 1089
rect 3761 1043 3809 1089
rect 3855 1043 3903 1089
rect 3949 1043 3997 1089
rect 4043 1043 4091 1089
rect 4137 1043 4185 1089
rect 4231 1043 4279 1089
rect 4325 1043 4373 1089
rect 4419 1043 4432 1089
rect 3608 1030 4432 1043
rect 178 -621 532 -608
rect 178 -667 191 -621
rect 237 -667 285 -621
rect 331 -667 379 -621
rect 425 -667 473 -621
rect 519 -667 532 -621
rect 178 -680 532 -667
rect 1225 -931 2049 -918
rect 1225 -977 1238 -931
rect 1284 -977 1332 -931
rect 1378 -977 1426 -931
rect 1472 -977 1520 -931
rect 1566 -977 1614 -931
rect 1660 -977 1708 -931
rect 1754 -977 1802 -931
rect 1848 -977 1896 -931
rect 1942 -977 1990 -931
rect 2036 -977 2049 -931
rect 1225 -990 2049 -977
rect 2937 -931 4902 -918
rect 2937 -977 2950 -931
rect 2996 -977 3044 -931
rect 3090 -977 3138 -931
rect 3184 -977 3232 -931
rect 3278 -977 3326 -931
rect 3372 -977 3420 -931
rect 3466 -977 3514 -931
rect 3560 -977 3621 -931
rect 3667 -977 3715 -931
rect 3761 -977 3809 -931
rect 3855 -977 3903 -931
rect 3949 -977 3997 -931
rect 4043 -977 4091 -931
rect 4137 -977 4185 -931
rect 4231 -977 4279 -931
rect 4325 -977 4373 -931
rect 4419 -977 4467 -931
rect 4513 -977 4561 -931
rect 4607 -977 4655 -931
rect 4701 -977 4749 -931
rect 4795 -977 4843 -931
rect 4889 -977 4902 -931
rect 2937 -990 4902 -977
<< psubdiffcont >>
rect 238 188 284 234
rect 332 188 378 234
rect 426 188 472 234
rect 814 33 860 79
rect 908 33 954 79
rect 1002 33 1048 79
rect 1096 33 1142 79
rect 1190 33 1236 79
rect 1284 33 1330 79
rect 1378 33 1424 79
rect 1472 33 1518 79
rect 1566 33 1612 79
rect 1660 33 1706 79
rect 1754 33 1800 79
rect 1848 33 1894 79
rect 1942 33 1988 79
rect 2036 33 2082 79
rect 2130 33 2176 79
rect 2224 33 2270 79
rect 2318 33 2364 79
rect 2412 33 2458 79
rect 3197 33 3243 79
rect 3291 33 3337 79
rect 3385 33 3431 79
rect 3479 33 3525 79
rect 3573 33 3619 79
rect 3667 33 3713 79
rect 3761 33 3807 79
rect 3855 33 3901 79
rect 3949 33 3995 79
rect 4043 33 4089 79
rect 4137 33 4183 79
rect 4231 33 4277 79
rect 4325 33 4371 79
rect 4419 33 4465 79
rect 4513 33 4559 79
rect 4607 33 4653 79
rect 4701 33 4747 79
rect 4795 33 4841 79
rect 238 -1522 284 -1476
rect 332 -1522 378 -1476
rect 426 -1522 472 -1476
rect 814 -1987 860 -1941
rect 908 -1987 954 -1941
rect 1002 -1987 1048 -1941
rect 1096 -1987 1142 -1941
rect 1190 -1987 1236 -1941
rect 1284 -1987 1330 -1941
rect 1378 -1987 1424 -1941
rect 1472 -1987 1518 -1941
rect 1566 -1987 1612 -1941
rect 1660 -1987 1706 -1941
rect 1754 -1987 1800 -1941
rect 1848 -1987 1894 -1941
rect 1942 -1987 1988 -1941
rect 2036 -1987 2082 -1941
rect 2130 -1987 2176 -1941
rect 2224 -1987 2270 -1941
rect 2318 -1987 2364 -1941
rect 2412 -1987 2458 -1941
rect 3177 -1993 3223 -1947
rect 3271 -1993 3317 -1947
rect 3365 -1993 3411 -1947
rect 3459 -1993 3505 -1947
rect 3553 -1993 3599 -1947
rect 3647 -1993 3693 -1947
rect 4165 -1993 4211 -1947
rect 4259 -1993 4305 -1947
rect 4353 -1993 4399 -1947
rect 4447 -1993 4493 -1947
rect 4541 -1993 4587 -1947
rect 4635 -1993 4681 -1947
rect 4729 -1993 4775 -1947
rect 4823 -1993 4869 -1947
rect 4917 -1993 4963 -1947
rect 5011 -1993 5057 -1947
rect 5105 -1993 5151 -1947
<< nsubdiffcont >>
rect 191 1043 237 1089
rect 285 1043 331 1089
rect 379 1043 425 1089
rect 473 1043 519 1089
rect 1238 1043 1284 1089
rect 1332 1043 1378 1089
rect 1426 1043 1472 1089
rect 1520 1043 1566 1089
rect 1614 1043 1660 1089
rect 1708 1043 1754 1089
rect 1802 1043 1848 1089
rect 1896 1043 1942 1089
rect 1990 1043 2036 1089
rect 3621 1043 3667 1089
rect 3715 1043 3761 1089
rect 3809 1043 3855 1089
rect 3903 1043 3949 1089
rect 3997 1043 4043 1089
rect 4091 1043 4137 1089
rect 4185 1043 4231 1089
rect 4279 1043 4325 1089
rect 4373 1043 4419 1089
rect 191 -667 237 -621
rect 285 -667 331 -621
rect 379 -667 425 -621
rect 473 -667 519 -621
rect 1238 -977 1284 -931
rect 1332 -977 1378 -931
rect 1426 -977 1472 -931
rect 1520 -977 1566 -931
rect 1614 -977 1660 -931
rect 1708 -977 1754 -931
rect 1802 -977 1848 -931
rect 1896 -977 1942 -931
rect 1990 -977 2036 -931
rect 2950 -977 2996 -931
rect 3044 -977 3090 -931
rect 3138 -977 3184 -931
rect 3232 -977 3278 -931
rect 3326 -977 3372 -931
rect 3420 -977 3466 -931
rect 3514 -977 3560 -931
rect 3621 -977 3667 -931
rect 3715 -977 3761 -931
rect 3809 -977 3855 -931
rect 3903 -977 3949 -931
rect 3997 -977 4043 -931
rect 4091 -977 4137 -931
rect 4185 -977 4231 -931
rect 4279 -977 4325 -931
rect 4373 -977 4419 -931
rect 4467 -977 4513 -931
rect 4561 -977 4607 -931
rect 4655 -977 4701 -931
rect 4749 -977 4795 -931
rect 4843 -977 4889 -931
<< polysilicon >>
rect 327 919 383 963
rect 1369 947 1425 991
rect 1529 947 1585 991
rect 1689 947 1745 991
rect 1849 947 1905 991
rect 3752 947 3808 991
rect 3912 947 3968 991
rect 4072 947 4128 991
rect 4232 947 4288 991
rect 327 553 383 719
rect 1056 703 1134 712
rect 1369 703 1425 747
rect 1056 699 1425 703
rect 1056 652 1069 699
rect 1116 652 1425 699
rect 1056 647 1425 652
rect 1056 639 1134 647
rect 431 553 503 561
rect 327 548 503 553
rect 327 502 444 548
rect 490 502 503 548
rect 327 497 503 502
rect 327 447 383 497
rect 431 489 503 497
rect 889 475 945 519
rect 1049 475 1105 519
rect 1209 475 1265 647
rect 1369 475 1425 519
rect 1529 475 1585 747
rect 1689 623 1745 747
rect 1849 727 1905 747
rect 1849 692 2385 727
rect 1849 671 2080 692
rect 2067 646 2080 671
rect 2126 671 2385 692
rect 2126 646 2139 671
rect 2067 633 2139 646
rect 1689 567 1905 623
rect 1689 475 1745 519
rect 1849 475 1905 567
rect 2009 475 2065 519
rect 2169 475 2225 519
rect 2329 475 2385 671
rect 3439 703 3517 712
rect 3752 703 3808 747
rect 3439 699 3808 703
rect 3439 652 3452 699
rect 3499 652 3808 699
rect 3439 647 3808 652
rect 3439 639 3517 647
rect 3272 475 3328 519
rect 3432 475 3488 519
rect 3592 475 3648 647
rect 3752 475 3808 519
rect 3912 475 3968 747
rect 4072 623 4128 747
rect 4232 727 4288 747
rect 4232 692 4768 727
rect 4232 671 4463 692
rect 4450 646 4463 671
rect 4509 671 4768 692
rect 4509 646 4522 671
rect 4450 633 4522 646
rect 4072 567 4288 623
rect 4072 475 4128 519
rect 4232 475 4288 567
rect 4392 475 4448 519
rect 4552 475 4608 519
rect 4712 475 4768 671
rect 889 355 945 375
rect 1049 355 1105 375
rect 1209 355 1265 375
rect 327 303 383 347
rect 889 299 1265 355
rect 1369 355 1425 375
rect 1529 355 1585 375
rect 1689 355 1745 375
rect 1369 299 1745 355
rect 1849 355 1905 375
rect 2009 355 2065 375
rect 2169 355 2225 375
rect 1849 299 2225 355
rect 2329 331 2385 375
rect 3272 355 3328 375
rect 3432 355 3488 375
rect 3592 355 3648 375
rect 3272 299 3648 355
rect 3752 355 3808 375
rect 3912 355 3968 375
rect 4072 355 4128 375
rect 3752 299 4128 355
rect 4232 355 4288 375
rect 4392 355 4448 375
rect 4552 355 4608 375
rect 4232 299 4608 355
rect 4712 331 4768 375
rect 1350 225 1424 234
rect 1472 225 1528 299
rect 1350 221 1528 225
rect 1350 169 1363 221
rect 1411 169 1528 221
rect 2169 252 2225 299
rect 2376 252 2449 261
rect 2169 248 2449 252
rect 2169 201 2389 248
rect 2436 201 2449 248
rect 2169 196 2449 201
rect 2376 188 2449 196
rect 3733 225 3807 234
rect 3855 225 3911 299
rect 3733 221 3911 225
rect 3733 169 3746 221
rect 3794 169 3911 221
rect 4552 252 4608 299
rect 4759 252 4832 261
rect 4552 248 4832 252
rect 4552 201 4772 248
rect 4819 201 4832 248
rect 4552 196 4832 201
rect 4759 188 4832 196
rect 1350 156 1424 169
rect 3733 156 3807 169
rect 327 75 383 119
rect 327 -75 383 -25
rect 1350 -57 1424 -44
rect 3733 -57 3807 -44
rect 431 -75 503 -67
rect 327 -80 503 -75
rect 327 -126 444 -80
rect 490 -126 503 -80
rect 1350 -109 1363 -57
rect 1411 -109 1528 -57
rect 2376 -84 2449 -76
rect 1350 -113 1528 -109
rect 1350 -122 1424 -113
rect 327 -131 503 -126
rect 327 -297 383 -131
rect 431 -139 503 -131
rect 1472 -187 1528 -113
rect 2169 -89 2449 -84
rect 2169 -136 2389 -89
rect 2436 -136 2449 -89
rect 3733 -109 3746 -57
rect 3794 -109 3911 -57
rect 4759 -84 4832 -76
rect 3733 -113 3911 -109
rect 3733 -122 3807 -113
rect 2169 -140 2449 -136
rect 2169 -187 2225 -140
rect 2376 -149 2449 -140
rect 3855 -187 3911 -113
rect 4552 -89 4832 -84
rect 4552 -136 4772 -89
rect 4819 -136 4832 -89
rect 4552 -140 4832 -136
rect 4552 -187 4608 -140
rect 4759 -149 4832 -140
rect 889 -243 1265 -187
rect 889 -263 945 -243
rect 1049 -263 1105 -243
rect 1209 -263 1265 -243
rect 1369 -243 1745 -187
rect 1369 -263 1425 -243
rect 1529 -263 1585 -243
rect 1689 -263 1745 -243
rect 1849 -243 2225 -187
rect 1849 -263 1905 -243
rect 2009 -263 2065 -243
rect 2169 -263 2225 -243
rect 2329 -263 2385 -219
rect 3272 -243 3648 -187
rect 3272 -263 3328 -243
rect 3432 -263 3488 -243
rect 3592 -263 3648 -243
rect 3752 -243 4128 -187
rect 3752 -263 3808 -243
rect 3912 -263 3968 -243
rect 4072 -263 4128 -243
rect 4232 -243 4608 -187
rect 4232 -263 4288 -243
rect 4392 -263 4448 -243
rect 4552 -263 4608 -243
rect 4712 -263 4768 -219
rect 889 -407 945 -363
rect 1049 -407 1105 -363
rect 327 -541 383 -497
rect 1056 -535 1134 -527
rect 1209 -535 1265 -363
rect 1369 -407 1425 -363
rect 1056 -540 1425 -535
rect 1056 -587 1069 -540
rect 1116 -587 1425 -540
rect 1056 -591 1425 -587
rect 1056 -600 1134 -591
rect 1369 -635 1425 -591
rect 1529 -635 1585 -363
rect 1689 -407 1745 -363
rect 1849 -455 1905 -363
rect 2009 -407 2065 -363
rect 2169 -407 2225 -363
rect 1689 -511 1905 -455
rect 1689 -635 1745 -511
rect 2067 -534 2139 -521
rect 2067 -559 2080 -534
rect 1849 -580 2080 -559
rect 2126 -559 2139 -534
rect 2329 -559 2385 -363
rect 3272 -407 3328 -363
rect 3432 -407 3488 -363
rect 2126 -580 2385 -559
rect 1849 -615 2385 -580
rect 3439 -535 3517 -527
rect 3592 -535 3648 -363
rect 3752 -407 3808 -363
rect 3439 -540 3808 -535
rect 3439 -587 3452 -540
rect 3499 -587 3808 -540
rect 3439 -591 3808 -587
rect 3439 -600 3517 -591
rect 1849 -635 1905 -615
rect 3752 -635 3808 -591
rect 3912 -635 3968 -363
rect 4072 -407 4128 -363
rect 4232 -455 4288 -363
rect 4392 -407 4448 -363
rect 4552 -407 4608 -363
rect 4072 -511 4288 -455
rect 4072 -635 4128 -511
rect 4450 -534 4522 -521
rect 4450 -559 4463 -534
rect 4232 -580 4463 -559
rect 4509 -559 4522 -534
rect 4712 -559 4768 -363
rect 4509 -580 4768 -559
rect 4232 -615 4768 -580
rect 4232 -635 4288 -615
rect 327 -791 383 -747
rect 1369 -879 1425 -835
rect 1529 -879 1585 -835
rect 1689 -879 1745 -835
rect 1849 -879 1905 -835
rect 3752 -879 3808 -835
rect 3912 -879 3968 -835
rect 4072 -879 4128 -835
rect 4232 -879 4288 -835
rect 327 -1157 383 -991
rect 1369 -1073 1425 -1029
rect 1529 -1073 1585 -1029
rect 1689 -1073 1745 -1029
rect 1849 -1073 1905 -1029
rect 431 -1157 503 -1149
rect 327 -1162 503 -1157
rect 327 -1208 444 -1162
rect 490 -1208 503 -1162
rect 327 -1213 503 -1208
rect 327 -1263 383 -1213
rect 431 -1221 503 -1213
rect 4396 -1078 4452 -1034
rect 4556 -1078 4612 -1034
rect 4716 -1078 4772 -1034
rect 3087 -1146 3143 -1102
rect 3247 -1146 3303 -1102
rect 3407 -1146 3463 -1102
rect 3567 -1146 3623 -1102
rect 3855 -1146 3911 -1102
rect 1056 -1317 1134 -1308
rect 1369 -1317 1425 -1273
rect 1056 -1321 1425 -1317
rect 327 -1407 383 -1363
rect 1056 -1368 1069 -1321
rect 1116 -1368 1425 -1321
rect 1056 -1373 1425 -1368
rect 1056 -1381 1134 -1373
rect 889 -1545 945 -1501
rect 1049 -1545 1105 -1501
rect 1209 -1545 1265 -1373
rect 1369 -1545 1425 -1501
rect 1529 -1545 1585 -1273
rect 1689 -1397 1745 -1273
rect 1849 -1293 1905 -1273
rect 1849 -1328 2385 -1293
rect 1849 -1349 2080 -1328
rect 2067 -1374 2080 -1349
rect 2126 -1349 2385 -1328
rect 2126 -1374 2139 -1349
rect 2067 -1387 2139 -1374
rect 1689 -1453 1905 -1397
rect 1689 -1545 1745 -1501
rect 1849 -1545 1905 -1453
rect 2009 -1545 2065 -1501
rect 2169 -1545 2225 -1501
rect 2329 -1545 2385 -1349
rect 3087 -1366 3143 -1346
rect 3247 -1366 3303 -1346
rect 3087 -1422 3303 -1366
rect 3091 -1489 3163 -1481
rect 3247 -1489 3303 -1422
rect 3091 -1494 3303 -1489
rect 3091 -1540 3104 -1494
rect 3150 -1540 3303 -1494
rect 3091 -1545 3303 -1540
rect 3091 -1553 3163 -1545
rect 3247 -1618 3303 -1545
rect 3407 -1366 3463 -1346
rect 3567 -1366 3623 -1346
rect 3407 -1422 3623 -1366
rect 3407 -1618 3463 -1422
rect 3535 -1510 3607 -1502
rect 3855 -1510 3911 -1346
rect 4203 -1437 4275 -1429
rect 4396 -1437 4452 -1278
rect 4203 -1442 4452 -1437
rect 4203 -1488 4216 -1442
rect 4262 -1488 4452 -1442
rect 4203 -1493 4452 -1488
rect 4203 -1501 4292 -1493
rect 3535 -1515 3911 -1510
rect 3535 -1561 3548 -1515
rect 3594 -1561 3911 -1515
rect 4236 -1550 4292 -1501
rect 4396 -1550 4452 -1493
rect 4556 -1550 4612 -1278
rect 4716 -1317 4772 -1278
rect 4713 -1325 4785 -1317
rect 4713 -1330 5070 -1325
rect 4713 -1376 4726 -1330
rect 4772 -1376 5070 -1330
rect 4713 -1381 5070 -1376
rect 4713 -1389 4785 -1381
rect 4716 -1550 4772 -1501
rect 5014 -1550 5070 -1381
rect 3535 -1566 3911 -1561
rect 3535 -1574 3623 -1566
rect 3567 -1618 3623 -1574
rect 889 -1665 945 -1645
rect 1049 -1665 1105 -1645
rect 1209 -1665 1265 -1645
rect 889 -1721 1265 -1665
rect 1369 -1665 1425 -1645
rect 1529 -1665 1585 -1645
rect 1689 -1665 1745 -1645
rect 1369 -1721 1745 -1665
rect 1849 -1665 1905 -1645
rect 2009 -1665 2065 -1645
rect 2169 -1665 2225 -1645
rect 1849 -1721 2225 -1665
rect 2329 -1689 2385 -1645
rect 4236 -1694 4292 -1650
rect 4396 -1694 4452 -1650
rect 4556 -1670 4612 -1650
rect 4716 -1670 4772 -1650
rect 1350 -1795 1424 -1786
rect 1472 -1795 1528 -1721
rect 1350 -1799 1528 -1795
rect 1350 -1851 1363 -1799
rect 1411 -1851 1528 -1799
rect 2169 -1768 2225 -1721
rect 2376 -1768 2449 -1759
rect 3247 -1762 3303 -1718
rect 2169 -1772 2449 -1768
rect 2169 -1819 2389 -1772
rect 2436 -1819 2449 -1772
rect 2169 -1824 2449 -1819
rect 2376 -1832 2449 -1824
rect 3045 -1810 3117 -1798
rect 3407 -1810 3463 -1718
rect 3567 -1762 3623 -1718
rect 4556 -1726 4772 -1670
rect 5014 -1694 5070 -1650
rect 3045 -1811 3463 -1810
rect 1350 -1864 1424 -1851
rect 3045 -1857 3058 -1811
rect 3104 -1857 3463 -1811
rect 4716 -1792 4772 -1726
rect 5057 -1792 5129 -1784
rect 4716 -1797 5129 -1792
rect 4716 -1843 5070 -1797
rect 5116 -1843 5129 -1797
rect 4716 -1848 5129 -1843
rect 5057 -1856 5129 -1848
rect 3045 -1866 3463 -1857
rect 3045 -1870 3117 -1866
<< polycontact >>
rect 1069 652 1116 699
rect 444 502 490 548
rect 2080 646 2126 692
rect 3452 652 3499 699
rect 4463 646 4509 692
rect 1363 169 1411 221
rect 2389 201 2436 248
rect 3746 169 3794 221
rect 4772 201 4819 248
rect 444 -126 490 -80
rect 1363 -109 1411 -57
rect 2389 -136 2436 -89
rect 3746 -109 3794 -57
rect 4772 -136 4819 -89
rect 1069 -587 1116 -540
rect 2080 -580 2126 -534
rect 3452 -587 3499 -540
rect 4463 -580 4509 -534
rect 444 -1208 490 -1162
rect 1069 -1368 1116 -1321
rect 2080 -1374 2126 -1328
rect 3104 -1540 3150 -1494
rect 4216 -1488 4262 -1442
rect 3548 -1561 3594 -1515
rect 4726 -1376 4772 -1330
rect 1363 -1851 1411 -1799
rect 2389 -1819 2436 -1772
rect 3058 -1857 3104 -1811
rect 5070 -1843 5116 -1797
<< metal1 >>
rect 2272 1553 2348 1565
rect 2272 1501 2284 1553
rect 2336 1550 2348 1553
rect 2336 1504 2799 1550
rect 2336 1501 2348 1504
rect 2272 1489 2348 1501
rect 690 1446 766 1458
rect 690 1443 702 1446
rect 377 1397 702 1443
rect 690 1394 702 1397
rect 754 1394 766 1446
rect 690 1382 766 1394
rect 2395 1446 2471 1458
rect 2395 1394 2407 1446
rect 2459 1443 2471 1446
rect 2459 1397 2799 1443
rect 2459 1394 2471 1397
rect 2395 1382 2471 1394
rect 554 1339 630 1351
rect 554 1336 566 1339
rect 377 1290 566 1336
rect 554 1287 566 1290
rect 618 1287 630 1339
rect 554 1275 630 1287
rect 2518 1339 2594 1351
rect 2518 1287 2530 1339
rect 2582 1336 2594 1339
rect 2582 1290 2799 1336
rect 2582 1287 2594 1290
rect 2518 1275 2594 1287
rect 2654 1232 2730 1244
rect 2654 1229 2666 1232
rect 377 1183 2666 1229
rect 2654 1180 2666 1183
rect 2718 1180 2730 1232
rect 2654 1168 2730 1180
rect 69 1092 4462 1122
rect 69 1040 99 1092
rect 151 1089 1611 1092
rect 1663 1089 4462 1092
rect 151 1043 191 1089
rect 237 1043 285 1089
rect 331 1043 379 1089
rect 425 1043 473 1089
rect 519 1043 1238 1089
rect 1284 1043 1332 1089
rect 1378 1043 1426 1089
rect 1472 1043 1520 1089
rect 1566 1043 1611 1089
rect 1663 1043 1708 1089
rect 1754 1043 1802 1089
rect 1848 1043 1896 1089
rect 1942 1043 1990 1089
rect 2036 1043 3621 1089
rect 3667 1043 3715 1089
rect 3761 1043 3809 1089
rect 3855 1043 3903 1089
rect 3949 1043 3997 1089
rect 4043 1043 4091 1089
rect 4137 1043 4185 1089
rect 4231 1043 4279 1089
rect 4325 1043 4373 1089
rect 4419 1043 4462 1089
rect 151 1040 1611 1043
rect 1663 1040 4462 1043
rect 69 1010 4462 1040
rect 252 906 298 917
rect 252 690 298 732
rect 412 906 458 1010
rect 1452 945 1498 1010
rect 412 721 458 732
rect 1294 934 1340 945
rect 1452 934 1500 945
rect 1452 916 1454 934
rect 1056 703 1127 710
rect 237 678 313 690
rect 237 675 249 678
rect 155 629 249 675
rect 237 626 249 629
rect 301 626 313 678
rect 688 647 700 703
rect 756 699 1127 703
rect 756 652 1069 699
rect 1116 652 1127 699
rect 756 647 1127 652
rect 688 635 768 647
rect 1056 641 1127 647
rect 1294 692 1340 760
rect 1454 749 1500 760
rect 1614 934 1660 945
rect 1614 692 1660 760
rect 1774 934 1820 1010
rect 3835 945 3881 1010
rect 1774 749 1820 760
rect 1934 934 1980 945
rect 3677 934 3723 945
rect 2272 798 2348 810
rect 2272 795 2284 798
rect 1980 760 2284 795
rect 1934 749 2284 760
rect 2272 746 2284 749
rect 2336 795 2348 798
rect 2336 749 2560 795
rect 3835 934 3883 945
rect 3835 916 3837 934
rect 2336 746 2348 749
rect 2272 734 2348 746
rect 2069 692 2137 703
rect 1294 646 2080 692
rect 2126 646 2137 692
rect 237 614 313 626
rect 252 434 298 614
rect 433 548 501 559
rect 682 558 762 570
rect 1294 565 1340 646
rect 2069 635 2137 646
rect 682 548 694 558
rect 414 502 444 548
rect 490 502 694 548
rect 750 502 762 558
rect 433 491 501 502
rect 682 490 762 502
rect 814 519 1340 565
rect 1454 519 2140 565
rect 814 462 860 519
rect 252 349 298 360
rect 412 434 458 445
rect 814 377 860 388
rect 974 462 1020 473
rect 412 267 458 360
rect 974 331 1020 388
rect 1134 462 1180 519
rect 1134 377 1180 388
rect 1294 462 1340 473
rect 1294 331 1340 388
rect 1454 462 1500 519
rect 1454 377 1500 388
rect 1614 462 1660 473
rect 1614 331 1660 388
rect 1774 462 1820 519
rect 1774 377 1820 388
rect 1934 462 1980 473
rect 974 285 1660 331
rect -99 237 505 267
rect -99 185 -69 237
rect -17 234 505 237
rect -17 188 238 234
rect 284 188 332 234
rect 378 188 426 234
rect 472 188 505 234
rect -17 185 505 188
rect -99 155 505 185
rect 552 222 632 234
rect 1082 222 1158 234
rect 1362 222 1422 232
rect 552 166 564 222
rect 620 170 1094 222
rect 1146 221 1422 222
rect 1146 170 1363 221
rect 620 169 1363 170
rect 1411 169 1422 221
rect 620 166 1422 169
rect 252 62 298 73
rect 252 -196 298 -12
rect 412 62 458 155
rect 552 154 632 166
rect 1082 158 1158 166
rect 1362 158 1422 166
rect 1934 112 1980 388
rect 2094 462 2140 519
rect 2094 377 2140 388
rect 2254 462 2300 473
rect 2254 112 2300 388
rect 2414 462 2460 749
rect 2652 703 2733 715
rect 3439 703 3510 710
rect 2652 647 2664 703
rect 2720 699 3510 703
rect 2720 652 3452 699
rect 3499 652 3510 699
rect 2720 647 3510 652
rect 2652 635 2733 647
rect 3439 641 3510 647
rect 3677 692 3723 760
rect 3837 749 3883 760
rect 3997 934 4043 945
rect 3997 692 4043 760
rect 4157 934 4203 1010
rect 4157 749 4203 760
rect 4317 934 4363 945
rect 4363 760 5362 795
rect 4317 749 5362 760
rect 4452 692 4520 703
rect 3677 646 4463 692
rect 4509 646 4520 692
rect 3677 565 3723 646
rect 4452 635 4520 646
rect 2414 377 2460 388
rect 3197 519 3723 565
rect 3837 519 4523 565
rect 3197 462 3243 519
rect 3197 377 3243 388
rect 3357 462 3403 473
rect 3357 331 3403 388
rect 3517 462 3563 519
rect 3517 377 3563 388
rect 3677 462 3723 473
rect 3677 331 3723 388
rect 3837 462 3883 519
rect 3837 377 3883 388
rect 3997 462 4043 473
rect 3997 331 4043 388
rect 4157 462 4203 519
rect 4157 377 4203 388
rect 4317 462 4363 473
rect 3357 285 4043 331
rect 2378 251 2436 259
rect 2651 251 2732 263
rect 2378 248 2663 251
rect 2378 201 2389 248
rect 2436 201 2663 248
rect 2378 195 2663 201
rect 2719 195 2732 251
rect 3745 222 3805 232
rect 2378 190 2436 195
rect 2651 183 2732 195
rect 3643 221 3805 222
rect 3643 169 3744 221
rect 3796 169 3805 221
rect 3643 166 3805 169
rect 3745 158 3805 166
rect 4317 112 4363 388
rect 4477 462 4523 519
rect 4477 377 4523 388
rect 4637 462 4683 473
rect 4637 112 4683 388
rect 4797 462 4843 749
rect 4797 377 4843 388
rect 4761 251 4819 259
rect 5056 251 5132 261
rect 4761 249 5132 251
rect 4761 248 5067 249
rect 4761 201 4772 248
rect 4819 201 5067 248
rect 4761 197 5067 201
rect 5119 197 5132 249
rect 4761 195 5132 197
rect 4761 190 4819 195
rect 5056 185 5132 195
rect 781 82 4875 112
rect 781 79 2033 82
rect 2085 79 4875 82
rect 781 33 814 79
rect 860 33 908 79
rect 954 33 1002 79
rect 1048 33 1096 79
rect 1142 33 1190 79
rect 1236 33 1284 79
rect 1330 33 1378 79
rect 1424 33 1472 79
rect 1518 33 1566 79
rect 1612 33 1660 79
rect 1706 33 1754 79
rect 1800 33 1848 79
rect 1894 33 1942 79
rect 1988 33 2033 79
rect 2085 33 2130 79
rect 2176 33 2224 79
rect 2270 33 2318 79
rect 2364 33 2412 79
rect 2458 33 3197 79
rect 3243 33 3291 79
rect 3337 33 3385 79
rect 3431 33 3479 79
rect 3525 33 3573 79
rect 3619 33 3667 79
rect 3713 33 3761 79
rect 3807 33 3855 79
rect 3901 33 3949 79
rect 3995 33 4043 79
rect 4089 33 4137 79
rect 4183 33 4231 79
rect 4277 33 4325 79
rect 4371 33 4419 79
rect 4465 33 4513 79
rect 4559 33 4607 79
rect 4653 33 4701 79
rect 4747 33 4795 79
rect 4841 33 4875 79
rect 781 30 2033 33
rect 2085 30 4875 33
rect 781 0 4875 30
rect 412 -23 458 -12
rect 552 -54 632 -42
rect 1362 -54 1422 -46
rect 433 -80 501 -69
rect 552 -80 564 -54
rect 414 -126 444 -80
rect 490 -110 564 -80
rect 620 -57 1422 -54
rect 620 -109 1363 -57
rect 1411 -109 1422 -57
rect 620 -110 1422 -109
rect 490 -122 632 -110
rect 1362 -120 1422 -110
rect 490 -126 582 -122
rect 433 -137 501 -126
rect 237 -207 313 -196
rect 155 -208 313 -207
rect 155 -253 249 -208
rect 237 -260 249 -253
rect 301 -260 313 -208
rect 237 -272 313 -260
rect 974 -219 1660 -173
rect 252 -310 298 -272
rect 814 -276 860 -265
rect 252 -495 298 -484
rect 412 -310 458 -299
rect 814 -407 860 -350
rect 974 -276 1020 -219
rect 974 -361 1020 -350
rect 1134 -276 1180 -265
rect 1134 -407 1180 -350
rect 1294 -276 1340 -219
rect 1294 -361 1340 -350
rect 1454 -276 1500 -265
rect 1454 -407 1500 -350
rect 1614 -276 1660 -219
rect 1614 -361 1660 -350
rect 1774 -276 1820 -265
rect 1774 -407 1820 -350
rect 1934 -276 1980 0
rect 1934 -361 1980 -350
rect 2094 -276 2140 -265
rect 2094 -407 2140 -350
rect 2254 -276 2300 0
rect 2914 -54 2990 -46
rect 3745 -54 3805 -46
rect 2914 -57 3805 -54
rect 2914 -58 3746 -57
rect 2378 -83 2436 -78
rect 2780 -83 2860 -71
rect 2378 -89 2792 -83
rect 2378 -136 2389 -89
rect 2436 -136 2792 -89
rect 2378 -139 2792 -136
rect 2848 -139 2860 -83
rect 2914 -110 2926 -58
rect 2978 -109 3746 -58
rect 3794 -109 3805 -57
rect 2978 -110 3805 -109
rect 2914 -122 2990 -110
rect 3745 -120 3805 -110
rect 2378 -147 2436 -139
rect 2780 -151 2860 -139
rect 3357 -219 4043 -173
rect 2254 -361 2300 -350
rect 2414 -276 2460 -265
rect 814 -453 1340 -407
rect 1454 -453 2140 -407
rect 412 -588 458 -484
rect 688 -535 768 -523
rect 1056 -535 1127 -529
rect 69 -618 557 -588
rect 688 -591 700 -535
rect 756 -540 1127 -535
rect 756 -587 1069 -540
rect 1116 -587 1127 -540
rect 756 -591 1127 -587
rect 688 -603 768 -591
rect 1056 -598 1127 -591
rect 1294 -534 1340 -453
rect 2069 -534 2137 -523
rect 1294 -580 2080 -534
rect 2126 -580 2137 -534
rect 69 -670 99 -618
rect 151 -621 557 -618
rect 151 -667 191 -621
rect 237 -667 285 -621
rect 331 -667 379 -621
rect 425 -667 473 -621
rect 519 -667 557 -621
rect 151 -670 557 -667
rect 69 -700 557 -670
rect 1294 -648 1340 -580
rect 252 -804 298 -793
rect 252 -1014 298 -978
rect 412 -804 458 -700
rect 1454 -648 1500 -637
rect 1294 -833 1340 -822
rect 1452 -822 1454 -804
rect 1452 -833 1500 -822
rect 1614 -648 1660 -580
rect 2069 -591 2137 -580
rect 2414 -622 2460 -350
rect 3197 -276 3243 -265
rect 3197 -407 3243 -350
rect 3357 -276 3403 -219
rect 3357 -361 3403 -350
rect 3517 -276 3563 -265
rect 3517 -407 3563 -350
rect 3677 -276 3723 -219
rect 3677 -361 3723 -350
rect 3837 -276 3883 -265
rect 3837 -407 3883 -350
rect 3997 -276 4043 -219
rect 3997 -361 4043 -350
rect 4157 -276 4203 -265
rect 4157 -407 4203 -350
rect 4317 -276 4363 0
rect 4317 -361 4363 -350
rect 4477 -276 4523 -265
rect 4477 -407 4523 -350
rect 4637 -276 4683 0
rect 4755 -83 4835 -72
rect 4755 -84 4940 -83
rect 4755 -140 4767 -84
rect 4823 -139 4940 -84
rect 4823 -140 4835 -139
rect 4755 -152 4835 -140
rect 4637 -361 4683 -350
rect 4797 -276 4843 -265
rect 3197 -453 3723 -407
rect 3837 -453 4523 -407
rect 2782 -532 2858 -520
rect 2782 -594 2794 -532
rect 2846 -535 2858 -532
rect 3439 -535 3510 -529
rect 2846 -540 3510 -535
rect 2846 -587 3452 -540
rect 3499 -587 3510 -540
rect 2846 -591 3510 -587
rect 2846 -594 2858 -591
rect 2782 -606 2858 -594
rect 3439 -598 3510 -591
rect 3677 -534 3723 -453
rect 4452 -534 4520 -523
rect 3677 -580 4463 -534
rect 4509 -580 4520 -534
rect 2395 -634 2471 -622
rect 2395 -637 2407 -634
rect 1614 -833 1660 -822
rect 1774 -648 1820 -637
rect 1452 -898 1498 -833
rect 1774 -898 1820 -822
rect 1934 -648 2407 -637
rect 1980 -683 2407 -648
rect 2395 -686 2407 -683
rect 2459 -637 2471 -634
rect 2459 -683 2560 -637
rect 3677 -648 3723 -580
rect 2459 -686 2471 -683
rect 2395 -698 2471 -686
rect 1934 -833 1980 -822
rect 3837 -648 3883 -637
rect 3677 -833 3723 -822
rect 3835 -822 3837 -804
rect 3835 -833 3883 -822
rect 3997 -648 4043 -580
rect 4452 -591 4520 -580
rect 4797 -637 4843 -350
rect 3997 -833 4043 -822
rect 4157 -648 4203 -637
rect 3835 -898 3881 -833
rect 4157 -898 4203 -822
rect 4317 -648 5362 -637
rect 4363 -683 5362 -648
rect 4317 -833 4363 -822
rect 412 -989 458 -978
rect 1195 -928 4946 -898
rect 1195 -931 1611 -928
rect 1663 -931 4946 -928
rect 1195 -977 1238 -931
rect 1284 -977 1332 -931
rect 1378 -977 1426 -931
rect 1472 -977 1520 -931
rect 1566 -977 1611 -931
rect 1663 -977 1708 -931
rect 1754 -977 1802 -931
rect 1848 -977 1896 -931
rect 1942 -977 1990 -931
rect 2036 -977 2950 -931
rect 2996 -977 3044 -931
rect 3090 -977 3138 -931
rect 3184 -977 3232 -931
rect 3278 -977 3326 -931
rect 3372 -977 3420 -931
rect 3466 -977 3514 -931
rect 3560 -977 3621 -931
rect 3667 -977 3715 -931
rect 3761 -977 3809 -931
rect 3855 -977 3903 -931
rect 3949 -977 3997 -931
rect 4043 -977 4091 -931
rect 4137 -977 4185 -931
rect 4231 -977 4279 -931
rect 4325 -977 4373 -931
rect 4419 -977 4467 -931
rect 4513 -977 4561 -931
rect 4607 -977 4655 -931
rect 4701 -977 4749 -931
rect 4795 -977 4843 -931
rect 4889 -977 4946 -931
rect 1195 -980 1611 -977
rect 1663 -980 4946 -977
rect 1195 -1010 4946 -980
rect 235 -1026 315 -1014
rect 235 -1035 247 -1026
rect 155 -1081 247 -1035
rect 235 -1082 247 -1081
rect 303 -1082 315 -1026
rect 1452 -1075 1498 -1010
rect 235 -1094 315 -1082
rect 1294 -1086 1340 -1075
rect 252 -1276 298 -1094
rect 427 -1151 507 -1139
rect 427 -1207 439 -1151
rect 495 -1162 507 -1151
rect 495 -1207 555 -1162
rect 427 -1208 444 -1207
rect 490 -1208 555 -1207
rect 427 -1219 507 -1208
rect 1452 -1086 1500 -1075
rect 1452 -1104 1454 -1086
rect 252 -1361 298 -1350
rect 412 -1276 458 -1265
rect 412 -1441 458 -1350
rect 688 -1317 768 -1305
rect 1056 -1317 1127 -1310
rect 688 -1373 700 -1317
rect 756 -1321 1127 -1317
rect 756 -1368 1069 -1321
rect 1116 -1368 1127 -1321
rect 756 -1373 1127 -1368
rect 688 -1385 768 -1373
rect 1056 -1379 1127 -1373
rect 1294 -1328 1340 -1260
rect 1454 -1271 1500 -1260
rect 1614 -1086 1660 -1075
rect 1614 -1328 1660 -1260
rect 1774 -1086 1820 -1010
rect 1774 -1271 1820 -1260
rect 1934 -1086 1980 -1075
rect 3012 -1159 3058 -1148
rect 2516 -1220 2596 -1208
rect 2516 -1225 2528 -1220
rect 1980 -1260 2528 -1225
rect 1934 -1271 2528 -1260
rect 2069 -1328 2137 -1317
rect 1294 -1374 2080 -1328
rect 2126 -1374 2137 -1328
rect -99 -1471 505 -1441
rect 1294 -1455 1340 -1374
rect 2069 -1385 2137 -1374
rect -99 -1523 -69 -1471
rect -17 -1476 505 -1471
rect -17 -1522 238 -1476
rect 284 -1522 332 -1476
rect 378 -1522 426 -1476
rect 472 -1522 505 -1476
rect -17 -1523 505 -1522
rect -99 -1553 505 -1523
rect 205 -1555 505 -1553
rect 393 -1908 505 -1555
rect 814 -1501 1340 -1455
rect 1454 -1501 2140 -1455
rect 814 -1558 860 -1501
rect 814 -1643 860 -1632
rect 974 -1558 1020 -1547
rect 974 -1689 1020 -1632
rect 1134 -1558 1180 -1501
rect 1134 -1643 1180 -1632
rect 1294 -1558 1340 -1547
rect 1294 -1689 1340 -1632
rect 1454 -1558 1500 -1501
rect 1454 -1643 1500 -1632
rect 1614 -1558 1660 -1547
rect 1614 -1689 1660 -1632
rect 1774 -1558 1820 -1501
rect 1774 -1643 1820 -1632
rect 1934 -1558 1980 -1547
rect 974 -1735 1660 -1689
rect 1362 -1798 1422 -1788
rect 1260 -1799 1422 -1798
rect 1260 -1851 1361 -1799
rect 1413 -1851 1422 -1799
rect 1260 -1854 1422 -1851
rect 1362 -1862 1422 -1854
rect 1934 -1908 1980 -1632
rect 2094 -1558 2140 -1501
rect 2094 -1643 2140 -1632
rect 2254 -1558 2300 -1547
rect 2254 -1908 2300 -1632
rect 2414 -1558 2460 -1271
rect 2516 -1276 2528 -1271
rect 2584 -1276 2596 -1220
rect 2516 -1288 2596 -1276
rect 3012 -1390 3058 -1333
rect 3172 -1159 3218 -1010
rect 3172 -1344 3218 -1333
rect 3332 -1102 3698 -1056
rect 3332 -1159 3378 -1102
rect 3332 -1390 3378 -1333
rect 3012 -1436 3378 -1390
rect 3492 -1159 3538 -1148
rect 2915 -1489 2993 -1478
rect 3093 -1489 3161 -1483
rect 2915 -1490 3161 -1489
rect 2915 -1544 2927 -1490
rect 2979 -1494 3161 -1490
rect 2979 -1540 3104 -1494
rect 3150 -1540 3161 -1494
rect 3492 -1504 3538 -1333
rect 3652 -1159 3698 -1102
rect 3652 -1344 3698 -1333
rect 3780 -1159 3826 -1148
rect 3780 -1442 3826 -1333
rect 3940 -1159 3986 -1010
rect 4321 -1091 4367 -1010
rect 4321 -1276 4367 -1265
rect 4481 -1091 4527 -1080
rect 4481 -1330 4527 -1265
rect 4641 -1091 4687 -1010
rect 4641 -1276 4687 -1265
rect 4801 -1091 4847 -1080
rect 4847 -1265 5362 -1230
rect 4801 -1276 5362 -1265
rect 4715 -1330 4783 -1319
rect 3940 -1344 3986 -1333
rect 4321 -1376 4726 -1330
rect 4772 -1376 4783 -1330
rect 4205 -1442 4273 -1431
rect 3780 -1488 4216 -1442
rect 4262 -1488 4273 -1442
rect 3492 -1515 3605 -1504
rect 3492 -1528 3548 -1515
rect 2979 -1544 3161 -1540
rect 2915 -1545 3161 -1544
rect 2915 -1556 2993 -1545
rect 3093 -1551 3161 -1545
rect 3332 -1561 3548 -1528
rect 3594 -1561 3605 -1515
rect 3780 -1558 3826 -1488
rect 4205 -1499 4273 -1488
rect 3332 -1572 3605 -1561
rect 3332 -1574 3538 -1572
rect 2414 -1643 2460 -1632
rect 3172 -1631 3218 -1620
rect 2378 -1769 2436 -1761
rect 2652 -1769 2732 -1757
rect 2378 -1772 2664 -1769
rect 2378 -1819 2389 -1772
rect 2436 -1819 2664 -1772
rect 2378 -1825 2664 -1819
rect 2720 -1825 2732 -1769
rect 2378 -1830 2436 -1825
rect 2652 -1837 2732 -1825
rect 2782 -1804 2858 -1792
rect 2782 -1856 2794 -1804
rect 2846 -1811 2858 -1804
rect 3047 -1811 3115 -1800
rect 2846 -1856 3058 -1811
rect 2782 -1857 3058 -1856
rect 3104 -1857 3115 -1811
rect 2782 -1868 2858 -1857
rect 3047 -1868 3115 -1857
rect 393 -1914 2492 -1908
rect 3172 -1914 3218 -1705
rect 3332 -1631 3378 -1574
rect 3652 -1604 3826 -1558
rect 4161 -1563 4207 -1552
rect 3332 -1716 3378 -1705
rect 3492 -1631 3538 -1620
rect 3492 -1914 3538 -1705
rect 3652 -1631 3698 -1604
rect 3652 -1716 3698 -1705
rect 4161 -1694 4207 -1637
rect 4321 -1563 4367 -1376
rect 4715 -1387 4783 -1376
rect 4321 -1648 4367 -1637
rect 4481 -1506 4847 -1460
rect 4481 -1563 4527 -1506
rect 4481 -1694 4527 -1637
rect 4161 -1740 4527 -1694
rect 4641 -1563 4687 -1552
rect 4641 -1914 4687 -1637
rect 4801 -1563 4847 -1506
rect 4801 -1648 4847 -1637
rect 4939 -1563 4985 -1552
rect 4939 -1914 4985 -1637
rect 5099 -1563 5145 -1276
rect 5099 -1648 5145 -1637
rect 5059 -1794 5127 -1786
rect 5059 -1846 5067 -1794
rect 5119 -1797 5127 -1794
rect 5119 -1843 5176 -1797
rect 5119 -1846 5127 -1843
rect 5059 -1854 5127 -1846
rect 393 -1938 5185 -1914
rect 393 -1941 2033 -1938
rect 2085 -1941 5185 -1938
rect 393 -1987 814 -1941
rect 860 -1987 908 -1941
rect 954 -1987 1002 -1941
rect 1048 -1987 1096 -1941
rect 1142 -1987 1190 -1941
rect 1236 -1987 1284 -1941
rect 1330 -1987 1378 -1941
rect 1424 -1987 1472 -1941
rect 1518 -1987 1566 -1941
rect 1612 -1987 1660 -1941
rect 1706 -1987 1754 -1941
rect 1800 -1987 1848 -1941
rect 1894 -1987 1942 -1941
rect 1988 -1987 2033 -1941
rect 2085 -1987 2130 -1941
rect 2176 -1987 2224 -1941
rect 2270 -1987 2318 -1941
rect 2364 -1987 2412 -1941
rect 2458 -1947 5185 -1941
rect 2458 -1987 3177 -1947
rect 393 -1990 2033 -1987
rect 2085 -1990 3177 -1987
rect 393 -1993 3177 -1990
rect 3223 -1993 3271 -1947
rect 3317 -1993 3365 -1947
rect 3411 -1993 3459 -1947
rect 3505 -1993 3553 -1947
rect 3599 -1993 3647 -1947
rect 3693 -1993 4165 -1947
rect 4211 -1993 4259 -1947
rect 4305 -1993 4353 -1947
rect 4399 -1993 4447 -1947
rect 4493 -1993 4541 -1947
rect 4587 -1993 4635 -1947
rect 4681 -1993 4729 -1947
rect 4775 -1993 4823 -1947
rect 4869 -1993 4917 -1947
rect 4963 -1993 5011 -1947
rect 5057 -1993 5105 -1947
rect 5151 -1993 5185 -1947
rect 393 -2020 5185 -1993
rect 3135 -2026 5185 -2020
<< via1 >>
rect 2284 1501 2336 1553
rect 702 1394 754 1446
rect 2407 1394 2459 1446
rect 566 1287 618 1339
rect 2530 1287 2582 1339
rect 2666 1180 2718 1232
rect 99 1040 151 1092
rect 1611 1089 1663 1092
rect 1611 1043 1614 1089
rect 1614 1043 1660 1089
rect 1660 1043 1663 1089
rect 1611 1040 1663 1043
rect 249 626 301 678
rect 700 647 756 703
rect 2284 746 2336 798
rect 694 502 750 558
rect -69 185 -17 237
rect 564 166 620 222
rect 1094 170 1146 222
rect 2664 647 2720 703
rect 2663 195 2719 251
rect 3744 169 3746 221
rect 3746 169 3794 221
rect 3794 169 3796 221
rect 5067 197 5119 249
rect 2033 79 2085 82
rect 2033 33 2036 79
rect 2036 33 2082 79
rect 2082 33 2085 79
rect 2033 30 2085 33
rect 564 -110 620 -54
rect 249 -260 301 -208
rect 2792 -139 2848 -83
rect 2926 -110 2978 -58
rect 700 -591 756 -535
rect 99 -670 151 -618
rect 4767 -89 4823 -84
rect 4767 -136 4772 -89
rect 4772 -136 4819 -89
rect 4819 -136 4823 -89
rect 4767 -140 4823 -136
rect 2794 -594 2846 -532
rect 2407 -686 2459 -634
rect 1611 -931 1663 -928
rect 1611 -977 1614 -931
rect 1614 -977 1660 -931
rect 1660 -977 1663 -931
rect 1611 -980 1663 -977
rect 247 -1082 303 -1026
rect 439 -1162 495 -1151
rect 439 -1207 444 -1162
rect 444 -1207 490 -1162
rect 490 -1207 495 -1162
rect 700 -1373 756 -1317
rect -69 -1523 -17 -1471
rect 1361 -1851 1363 -1799
rect 1363 -1851 1411 -1799
rect 1411 -1851 1413 -1799
rect 2528 -1276 2584 -1220
rect 2927 -1544 2979 -1490
rect 2664 -1825 2720 -1769
rect 2794 -1856 2846 -1804
rect 5067 -1797 5119 -1794
rect 5067 -1843 5070 -1797
rect 5070 -1843 5116 -1797
rect 5116 -1843 5119 -1797
rect 5067 -1846 5119 -1843
rect 2033 -1941 2085 -1938
rect 2033 -1987 2036 -1941
rect 2036 -1987 2082 -1941
rect 2082 -1987 2085 -1941
rect 2033 -1990 2085 -1987
<< metal2 >>
rect 2272 1553 2348 1565
rect 2272 1501 2284 1553
rect 2336 1501 2348 1553
rect 2272 1489 2348 1501
rect 690 1446 766 1458
rect 690 1394 702 1446
rect 754 1394 766 1446
rect 690 1382 766 1394
rect 554 1339 630 1351
rect 554 1287 566 1339
rect 618 1287 630 1339
rect 554 1275 630 1287
rect 69 1092 181 1122
rect 69 1040 99 1092
rect 151 1040 181 1092
rect -99 237 13 267
rect -99 185 -69 237
rect -17 185 13 237
rect -99 -1471 13 185
rect 69 -618 181 1040
rect 237 680 313 690
rect 237 624 247 680
rect 303 624 313 680
rect 237 614 313 624
rect 564 234 620 1275
rect 700 715 756 1382
rect 1581 1092 1693 1122
rect 1581 1040 1611 1092
rect 1663 1040 1693 1092
rect 688 703 768 715
rect 688 647 700 703
rect 756 647 768 703
rect 688 635 768 647
rect 700 570 756 635
rect 682 558 762 570
rect 682 502 694 558
rect 750 502 762 558
rect 682 490 762 502
rect 552 222 632 234
rect 552 166 564 222
rect 620 166 632 222
rect 552 154 632 166
rect 564 -42 620 154
rect 552 -54 632 -42
rect 552 -110 564 -54
rect 620 -110 632 -54
rect 700 -74 756 490
rect 1082 225 1158 234
rect 1082 169 1092 225
rect 1148 169 1158 225
rect 1082 158 1158 169
rect 552 -122 632 -110
rect 690 -84 766 -74
rect 690 -140 700 -84
rect 756 -140 766 -84
rect 690 -150 766 -140
rect 237 -206 313 -196
rect 237 -262 247 -206
rect 303 -262 313 -206
rect 237 -272 313 -262
rect 700 -523 756 -150
rect 688 -535 768 -523
rect 688 -591 700 -535
rect 756 -591 768 -535
rect 688 -603 768 -591
rect 69 -670 99 -618
rect 151 -670 181 -618
rect 69 -700 181 -670
rect 235 -1026 315 -1014
rect 235 -1082 247 -1026
rect 303 -1082 315 -1026
rect 235 -1094 315 -1082
rect 427 -1151 507 -1139
rect 427 -1207 439 -1151
rect 495 -1207 507 -1151
rect 427 -1219 507 -1207
rect 700 -1305 756 -603
rect 1581 -928 1693 1040
rect 2282 810 2338 1489
rect 2395 1446 2471 1458
rect 2395 1394 2407 1446
rect 2459 1394 2471 1446
rect 2395 1382 2471 1394
rect 2272 798 2348 810
rect 2272 746 2284 798
rect 2336 746 2348 798
rect 2272 734 2348 746
rect 1581 -980 1611 -928
rect 1663 -980 1693 -928
rect 1581 -1010 1693 -980
rect 2003 82 2115 112
rect 2003 30 2033 82
rect 2085 30 2115 82
rect 688 -1317 768 -1305
rect 688 -1373 700 -1317
rect 756 -1373 768 -1317
rect 688 -1385 768 -1373
rect -99 -1523 -69 -1471
rect -17 -1523 13 -1471
rect -99 -1553 13 -1523
rect 1349 -1797 1425 -1787
rect 1349 -1853 1359 -1797
rect 1415 -1853 1425 -1797
rect 1349 -1863 1425 -1853
rect 2003 -1938 2115 30
rect 2405 -622 2461 1382
rect 2518 1339 2594 1351
rect 2518 1287 2530 1339
rect 2582 1287 2594 1339
rect 2518 1275 2594 1287
rect 2395 -634 2471 -622
rect 2395 -686 2407 -634
rect 2459 -686 2471 -634
rect 2395 -698 2471 -686
rect 2528 -1208 2584 1275
rect 2654 1232 2730 1244
rect 2654 1180 2666 1232
rect 2718 1180 2730 1232
rect 2654 1168 2730 1180
rect 2664 715 2720 1168
rect 2652 703 2733 715
rect 2652 647 2664 703
rect 2720 647 2733 703
rect 2652 635 2733 647
rect 5065 680 5121 690
rect 2664 263 2720 635
rect 2651 251 2732 263
rect 2651 195 2663 251
rect 2719 195 2732 251
rect 5065 249 5121 624
rect 2651 183 2732 195
rect 3732 223 3808 233
rect 2664 -1141 2720 183
rect 3732 167 3742 223
rect 3798 167 3808 223
rect 3732 157 3808 167
rect 5065 197 5067 249
rect 5119 197 5121 249
rect 2924 -58 2980 -46
rect 2780 -83 2860 -71
rect 2780 -139 2792 -83
rect 2848 -139 2860 -83
rect 2780 -151 2860 -139
rect 2924 -110 2926 -58
rect 2978 -110 2980 -58
rect 2792 -532 2848 -151
rect 2924 -196 2980 -110
rect 4757 -84 4833 -74
rect 4757 -140 4767 -84
rect 4823 -140 4833 -84
rect 4757 -150 4833 -140
rect 2914 -206 2990 -196
rect 2914 -262 2924 -206
rect 2980 -262 2990 -206
rect 2914 -272 2990 -262
rect 2792 -594 2794 -532
rect 2846 -594 2848 -532
rect 2792 -1016 2848 -594
rect 2782 -1026 2858 -1016
rect 2782 -1082 2792 -1026
rect 2848 -1082 2858 -1026
rect 2782 -1092 2858 -1082
rect 2654 -1151 2730 -1141
rect 2654 -1207 2664 -1151
rect 2720 -1207 2730 -1151
rect 2516 -1220 2596 -1208
rect 2654 -1217 2730 -1207
rect 2516 -1276 2528 -1220
rect 2584 -1276 2596 -1220
rect 2516 -1288 2596 -1276
rect 2664 -1757 2720 -1217
rect 2652 -1769 2732 -1757
rect 2652 -1825 2664 -1769
rect 2720 -1825 2732 -1769
rect 2652 -1837 2732 -1825
rect 2792 -1804 2848 -1092
rect 2924 -1478 2980 -272
rect 2915 -1490 2993 -1478
rect 2915 -1544 2927 -1490
rect 2979 -1544 2993 -1490
rect 2915 -1556 2993 -1544
rect 2924 -1787 2980 -1556
rect 2792 -1856 2794 -1804
rect 2846 -1856 2848 -1804
rect 2792 -1868 2848 -1856
rect 2914 -1797 2990 -1787
rect 2914 -1853 2924 -1797
rect 2980 -1853 2990 -1797
rect 2914 -1863 2990 -1853
rect 5065 -1794 5121 197
rect 5065 -1846 5067 -1794
rect 5119 -1846 5121 -1794
rect 5065 -1858 5121 -1846
rect 2003 -1990 2033 -1938
rect 2085 -1990 2115 -1938
rect 2003 -2020 2115 -1990
<< via2 >>
rect 247 678 303 680
rect 247 626 249 678
rect 249 626 301 678
rect 301 626 303 678
rect 247 624 303 626
rect 1092 222 1148 225
rect 1092 170 1094 222
rect 1094 170 1146 222
rect 1146 170 1148 222
rect 1092 169 1148 170
rect 700 -140 756 -84
rect 247 -208 303 -206
rect 247 -260 249 -208
rect 249 -260 301 -208
rect 301 -260 303 -208
rect 247 -262 303 -260
rect 247 -1082 303 -1026
rect 439 -1207 495 -1151
rect 1359 -1799 1415 -1797
rect 1359 -1851 1361 -1799
rect 1361 -1851 1413 -1799
rect 1413 -1851 1415 -1799
rect 1359 -1853 1415 -1851
rect 5065 624 5121 680
rect 3742 221 3798 223
rect 3742 169 3744 221
rect 3744 169 3796 221
rect 3796 169 3798 221
rect 3742 167 3798 169
rect 4767 -140 4823 -84
rect 2924 -262 2980 -206
rect 2792 -1082 2848 -1026
rect 2664 -1207 2720 -1151
rect 2924 -1853 2980 -1797
<< metal3 >>
rect 237 680 313 690
rect 5055 680 5131 690
rect 237 624 247 680
rect 303 624 5065 680
rect 5121 624 5131 680
rect 237 614 313 624
rect 5055 614 5131 624
rect 1082 225 1158 234
rect 1082 169 1092 225
rect 1148 223 1158 225
rect 2234 223 2389 224
rect 3732 223 3808 233
rect 1148 169 3742 223
rect 1082 167 3742 169
rect 3798 167 3808 223
rect 1082 158 1158 167
rect 3732 157 3808 167
rect 690 -84 766 -74
rect 4757 -84 4833 -74
rect 690 -140 700 -84
rect 756 -140 4767 -84
rect 4823 -140 4833 -84
rect 690 -150 766 -140
rect 4757 -150 4833 -140
rect 237 -206 313 -196
rect 2914 -206 2990 -196
rect 237 -262 247 -206
rect 303 -262 2924 -206
rect 2980 -262 2990 -206
rect 237 -272 313 -262
rect 2914 -272 2990 -262
rect 237 -1026 313 -1016
rect 2782 -1026 2858 -1016
rect 237 -1082 247 -1026
rect 303 -1082 2792 -1026
rect 2848 -1082 2858 -1026
rect 237 -1092 313 -1082
rect 2782 -1092 2858 -1082
rect 427 -1151 507 -1139
rect 2654 -1151 2730 -1141
rect 427 -1207 439 -1151
rect 495 -1207 2664 -1151
rect 2720 -1207 2730 -1151
rect 427 -1219 507 -1207
rect 2654 -1217 2730 -1207
rect 1349 -1797 1425 -1787
rect 2914 -1797 2990 -1781
rect 1349 -1853 1359 -1797
rect 1415 -1853 2924 -1797
rect 2980 -1853 2990 -1797
rect 1349 -1863 1425 -1853
rect 2914 -1863 2990 -1853
<< labels >>
flabel metal1 400 1313 400 1313 0 FreeSans 320 0 0 0 B
port 1 nsew
flabel metal1 400 1206 400 1206 0 FreeSans 320 0 0 0 C
port 2 nsew
flabel metal1 400 1420 400 1420 0 FreeSans 320 0 0 0 A
port 0 nsew
flabel metal1 5339 -1253 5339 -1253 0 FreeSans 320 0 0 0 S1
port 4 nsew
flabel metal1 5339 -660 5339 -660 0 FreeSans 320 0 0 0 S3
port 5 nsew
flabel metal1 5339 772 5339 772 0 FreeSans 320 0 0 0 S2
port 6 nsew
flabel metal1 2776 1527 2776 1527 0 FreeSans 320 0 0 0 S6
port 7 nsew
flabel metal1 2776 1420 2776 1420 0 FreeSans 320 0 0 0 S5
port 8 nsew
flabel metal1 2776 1313 2776 1313 0 FreeSans 320 0 0 0 S4
port 9 nsew
flabel metal1 3209 1066 3209 1066 0 FreeSans 320 0 0 0 VDD
port 11 nsew
flabel metal1 3014 -1964 3014 -1964 0 FreeSans 320 0 0 0 VSS
port 12 nsew
flabel psubdiffcont 355 -1499 355 -1499 0 FreeSans 320 0 0 0 Inverter_Layout_0.VSS
flabel metal1 355 -641 355 -641 0 FreeSans 320 0 0 0 Inverter_Layout_0.VDD
flabel metal1 535 -1185 535 -1185 0 FreeSans 320 0 0 0 Inverter_Layout_0.IN
flabel metal1 216 -1058 216 -1058 0 FreeSans 320 0 0 0 Inverter_Layout_0.OUT
flabel metal1 1270 -1828 1270 -1828 0 FreeSans 320 0 0 0 AND_3_In_Layout_0.B
flabel metal1 2537 -1251 2537 -1251 0 FreeSans 320 0 0 0 AND_3_In_Layout_0.OUT
flabel nsubdiffcont 1637 -954 1637 -954 0 FreeSans 320 0 0 0 AND_3_In_Layout_0.VDD
flabel psubdiff 1635 -1964 1635 -1964 0 FreeSans 320 0 0 0 AND_3_In_Layout_0.VSS
flabel metal1 2547 -1799 2547 -1799 0 FreeSans 320 180 0 0 AND_3_In_Layout_0.C
flabel metal1 990 -1351 990 -1351 0 FreeSans 320 0 0 0 AND_3_In_Layout_0.A
flabel metal1 1270 -80 1270 -80 0 FreeSans 320 0 0 0 AND_3_In_Layout_4.B
flabel metal1 2537 -657 2537 -657 0 FreeSans 320 0 0 0 AND_3_In_Layout_4.OUT
flabel nsubdiffcont 1637 -954 1637 -954 0 FreeSans 320 0 0 0 AND_3_In_Layout_4.VDD
flabel psubdiff 1635 56 1635 56 0 FreeSans 320 0 0 0 AND_3_In_Layout_4.VSS
flabel metal1 2547 -109 2547 -109 0 FreeSans 320 180 0 0 AND_3_In_Layout_4.C
flabel metal1 990 -557 990 -557 0 FreeSans 320 0 0 0 AND_3_In_Layout_4.A
flabel metal1 3490 -954 3490 -954 0 FreeSans 320 0 0 0 OR_2_In_Layout_0.VDD
flabel metal1 3443 -1970 3443 -1970 0 FreeSans 320 0 0 0 OR_2_In_Layout_0.VSS
flabel polycontact 3127 -1517 3127 -1517 0 FreeSans 320 0 0 0 OR_2_In_Layout_0.A
flabel polycontact 3081 -1834 3081 -1834 0 FreeSans 320 0 0 0 OR_2_In_Layout_0.B
flabel metal1 3970 -1458 3970 -1458 0 FreeSans 320 0 0 0 OR_2_In_Layout_0.OUT
flabel metal1 3653 -80 3653 -80 0 FreeSans 320 0 0 0 AND_3_In_Layout_2.B
flabel metal1 4920 -657 4920 -657 0 FreeSans 320 0 0 0 AND_3_In_Layout_2.OUT
flabel nsubdiffcont 4020 -954 4020 -954 0 FreeSans 320 0 0 0 AND_3_In_Layout_2.VDD
flabel psubdiff 4018 56 4018 56 0 FreeSans 320 0 0 0 AND_3_In_Layout_2.VSS
flabel metal1 4930 -109 4930 -109 0 FreeSans 320 180 0 0 AND_3_In_Layout_2.C
flabel metal1 3373 -557 3373 -557 0 FreeSans 320 0 0 0 AND_3_In_Layout_2.A
flabel metal1 4195 -1465 4195 -1465 0 FreeSans 320 0 0 0 AND_2_In_Layout_0.A
flabel metal1 5149 -1253 5149 -1253 0 FreeSans 320 0 0 0 AND_2_In_Layout_0.OUT
flabel nsubdiffcont 4584 -954 4584 -954 0 FreeSans 320 0 0 0 AND_2_In_Layout_0.VDD
flabel metal1 5162 -1820 5162 -1820 0 FreeSans 320 180 0 0 AND_2_In_Layout_0.B
flabel psubdiffcont 4658 -1970 4658 -1970 0 FreeSans 320 0 0 0 AND_2_In_Layout_0.VSS
flabel psubdiffcont 355 211 355 211 0 FreeSans 320 0 0 0 Inverter_Layout_1.VSS
flabel metal1 355 1069 355 1069 0 FreeSans 320 0 0 0 Inverter_Layout_1.VDD
flabel metal1 535 525 535 525 0 FreeSans 320 0 0 0 Inverter_Layout_1.IN
flabel metal1 216 652 216 652 0 FreeSans 320 0 0 0 Inverter_Layout_1.OUT
flabel psubdiffcont 355 211 355 211 0 FreeSans 320 0 0 0 Inverter_Layout_2.VSS
flabel metal1 355 -647 355 -647 0 FreeSans 320 0 0 0 Inverter_Layout_2.VDD
flabel metal1 535 -103 535 -103 0 FreeSans 320 0 0 0 Inverter_Layout_2.IN
flabel metal1 216 -230 216 -230 0 FreeSans 320 0 0 0 Inverter_Layout_2.OUT
flabel metal1 1270 192 1270 192 0 FreeSans 320 0 0 0 AND_3_In_Layout_3.B
flabel metal1 2537 769 2537 769 0 FreeSans 320 0 0 0 AND_3_In_Layout_3.OUT
flabel nsubdiffcont 1637 1066 1637 1066 0 FreeSans 320 0 0 0 AND_3_In_Layout_3.VDD
flabel psubdiff 1635 56 1635 56 0 FreeSans 320 0 0 0 AND_3_In_Layout_3.VSS
flabel metal1 2547 221 2547 221 0 FreeSans 320 180 0 0 AND_3_In_Layout_3.C
flabel metal1 990 669 990 669 0 FreeSans 320 0 0 0 AND_3_In_Layout_3.A
flabel metal1 3653 192 3653 192 0 FreeSans 320 0 0 0 AND_3_In_Layout_1.B
flabel metal1 4920 769 4920 769 0 FreeSans 320 0 0 0 AND_3_In_Layout_1.OUT
flabel nsubdiffcont 4020 1066 4020 1066 0 FreeSans 320 0 0 0 AND_3_In_Layout_1.VDD
flabel psubdiff 4018 56 4018 56 0 FreeSans 320 0 0 0 AND_3_In_Layout_1.VSS
flabel metal1 4930 221 4930 221 0 FreeSans 320 180 0 0 AND_3_In_Layout_1.C
flabel metal1 3373 669 3373 669 0 FreeSans 320 0 0 0 AND_3_In_Layout_1.A
<< end >>
