magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -8888 2128 8888
<< nwell >>
rect -128 -6888 128 6888
<< nsubdiff >>
rect -45 6783 45 6805
rect -45 6737 -23 6783
rect 23 6737 45 6783
rect -45 6679 45 6737
rect -45 6633 -23 6679
rect 23 6633 45 6679
rect -45 6575 45 6633
rect -45 6529 -23 6575
rect 23 6529 45 6575
rect -45 6471 45 6529
rect -45 6425 -23 6471
rect 23 6425 45 6471
rect -45 6367 45 6425
rect -45 6321 -23 6367
rect 23 6321 45 6367
rect -45 6263 45 6321
rect -45 6217 -23 6263
rect 23 6217 45 6263
rect -45 6159 45 6217
rect -45 6113 -23 6159
rect 23 6113 45 6159
rect -45 6055 45 6113
rect -45 6009 -23 6055
rect 23 6009 45 6055
rect -45 5951 45 6009
rect -45 5905 -23 5951
rect 23 5905 45 5951
rect -45 5847 45 5905
rect -45 5801 -23 5847
rect 23 5801 45 5847
rect -45 5743 45 5801
rect -45 5697 -23 5743
rect 23 5697 45 5743
rect -45 5639 45 5697
rect -45 5593 -23 5639
rect 23 5593 45 5639
rect -45 5535 45 5593
rect -45 5489 -23 5535
rect 23 5489 45 5535
rect -45 5431 45 5489
rect -45 5385 -23 5431
rect 23 5385 45 5431
rect -45 5327 45 5385
rect -45 5281 -23 5327
rect 23 5281 45 5327
rect -45 5223 45 5281
rect -45 5177 -23 5223
rect 23 5177 45 5223
rect -45 5119 45 5177
rect -45 5073 -23 5119
rect 23 5073 45 5119
rect -45 5015 45 5073
rect -45 4969 -23 5015
rect 23 4969 45 5015
rect -45 4911 45 4969
rect -45 4865 -23 4911
rect 23 4865 45 4911
rect -45 4807 45 4865
rect -45 4761 -23 4807
rect 23 4761 45 4807
rect -45 4703 45 4761
rect -45 4657 -23 4703
rect 23 4657 45 4703
rect -45 4599 45 4657
rect -45 4553 -23 4599
rect 23 4553 45 4599
rect -45 4495 45 4553
rect -45 4449 -23 4495
rect 23 4449 45 4495
rect -45 4391 45 4449
rect -45 4345 -23 4391
rect 23 4345 45 4391
rect -45 4287 45 4345
rect -45 4241 -23 4287
rect 23 4241 45 4287
rect -45 4183 45 4241
rect -45 4137 -23 4183
rect 23 4137 45 4183
rect -45 4079 45 4137
rect -45 4033 -23 4079
rect 23 4033 45 4079
rect -45 3975 45 4033
rect -45 3929 -23 3975
rect 23 3929 45 3975
rect -45 3871 45 3929
rect -45 3825 -23 3871
rect 23 3825 45 3871
rect -45 3767 45 3825
rect -45 3721 -23 3767
rect 23 3721 45 3767
rect -45 3663 45 3721
rect -45 3617 -23 3663
rect 23 3617 45 3663
rect -45 3559 45 3617
rect -45 3513 -23 3559
rect 23 3513 45 3559
rect -45 3455 45 3513
rect -45 3409 -23 3455
rect 23 3409 45 3455
rect -45 3351 45 3409
rect -45 3305 -23 3351
rect 23 3305 45 3351
rect -45 3247 45 3305
rect -45 3201 -23 3247
rect 23 3201 45 3247
rect -45 3143 45 3201
rect -45 3097 -23 3143
rect 23 3097 45 3143
rect -45 3039 45 3097
rect -45 2993 -23 3039
rect 23 2993 45 3039
rect -45 2935 45 2993
rect -45 2889 -23 2935
rect 23 2889 45 2935
rect -45 2831 45 2889
rect -45 2785 -23 2831
rect 23 2785 45 2831
rect -45 2727 45 2785
rect -45 2681 -23 2727
rect 23 2681 45 2727
rect -45 2623 45 2681
rect -45 2577 -23 2623
rect 23 2577 45 2623
rect -45 2519 45 2577
rect -45 2473 -23 2519
rect 23 2473 45 2519
rect -45 2415 45 2473
rect -45 2369 -23 2415
rect 23 2369 45 2415
rect -45 2311 45 2369
rect -45 2265 -23 2311
rect 23 2265 45 2311
rect -45 2207 45 2265
rect -45 2161 -23 2207
rect 23 2161 45 2207
rect -45 2103 45 2161
rect -45 2057 -23 2103
rect 23 2057 45 2103
rect -45 1999 45 2057
rect -45 1953 -23 1999
rect 23 1953 45 1999
rect -45 1895 45 1953
rect -45 1849 -23 1895
rect 23 1849 45 1895
rect -45 1791 45 1849
rect -45 1745 -23 1791
rect 23 1745 45 1791
rect -45 1687 45 1745
rect -45 1641 -23 1687
rect 23 1641 45 1687
rect -45 1583 45 1641
rect -45 1537 -23 1583
rect 23 1537 45 1583
rect -45 1479 45 1537
rect -45 1433 -23 1479
rect 23 1433 45 1479
rect -45 1375 45 1433
rect -45 1329 -23 1375
rect 23 1329 45 1375
rect -45 1271 45 1329
rect -45 1225 -23 1271
rect 23 1225 45 1271
rect -45 1167 45 1225
rect -45 1121 -23 1167
rect 23 1121 45 1167
rect -45 1063 45 1121
rect -45 1017 -23 1063
rect 23 1017 45 1063
rect -45 959 45 1017
rect -45 913 -23 959
rect 23 913 45 959
rect -45 855 45 913
rect -45 809 -23 855
rect 23 809 45 855
rect -45 751 45 809
rect -45 705 -23 751
rect 23 705 45 751
rect -45 647 45 705
rect -45 601 -23 647
rect 23 601 45 647
rect -45 543 45 601
rect -45 497 -23 543
rect 23 497 45 543
rect -45 439 45 497
rect -45 393 -23 439
rect 23 393 45 439
rect -45 335 45 393
rect -45 289 -23 335
rect 23 289 45 335
rect -45 231 45 289
rect -45 185 -23 231
rect 23 185 45 231
rect -45 127 45 185
rect -45 81 -23 127
rect 23 81 45 127
rect -45 23 45 81
rect -45 -23 -23 23
rect 23 -23 45 23
rect -45 -81 45 -23
rect -45 -127 -23 -81
rect 23 -127 45 -81
rect -45 -185 45 -127
rect -45 -231 -23 -185
rect 23 -231 45 -185
rect -45 -289 45 -231
rect -45 -335 -23 -289
rect 23 -335 45 -289
rect -45 -393 45 -335
rect -45 -439 -23 -393
rect 23 -439 45 -393
rect -45 -497 45 -439
rect -45 -543 -23 -497
rect 23 -543 45 -497
rect -45 -601 45 -543
rect -45 -647 -23 -601
rect 23 -647 45 -601
rect -45 -705 45 -647
rect -45 -751 -23 -705
rect 23 -751 45 -705
rect -45 -809 45 -751
rect -45 -855 -23 -809
rect 23 -855 45 -809
rect -45 -913 45 -855
rect -45 -959 -23 -913
rect 23 -959 45 -913
rect -45 -1017 45 -959
rect -45 -1063 -23 -1017
rect 23 -1063 45 -1017
rect -45 -1121 45 -1063
rect -45 -1167 -23 -1121
rect 23 -1167 45 -1121
rect -45 -1225 45 -1167
rect -45 -1271 -23 -1225
rect 23 -1271 45 -1225
rect -45 -1329 45 -1271
rect -45 -1375 -23 -1329
rect 23 -1375 45 -1329
rect -45 -1433 45 -1375
rect -45 -1479 -23 -1433
rect 23 -1479 45 -1433
rect -45 -1537 45 -1479
rect -45 -1583 -23 -1537
rect 23 -1583 45 -1537
rect -45 -1641 45 -1583
rect -45 -1687 -23 -1641
rect 23 -1687 45 -1641
rect -45 -1745 45 -1687
rect -45 -1791 -23 -1745
rect 23 -1791 45 -1745
rect -45 -1849 45 -1791
rect -45 -1895 -23 -1849
rect 23 -1895 45 -1849
rect -45 -1953 45 -1895
rect -45 -1999 -23 -1953
rect 23 -1999 45 -1953
rect -45 -2057 45 -1999
rect -45 -2103 -23 -2057
rect 23 -2103 45 -2057
rect -45 -2161 45 -2103
rect -45 -2207 -23 -2161
rect 23 -2207 45 -2161
rect -45 -2265 45 -2207
rect -45 -2311 -23 -2265
rect 23 -2311 45 -2265
rect -45 -2369 45 -2311
rect -45 -2415 -23 -2369
rect 23 -2415 45 -2369
rect -45 -2473 45 -2415
rect -45 -2519 -23 -2473
rect 23 -2519 45 -2473
rect -45 -2577 45 -2519
rect -45 -2623 -23 -2577
rect 23 -2623 45 -2577
rect -45 -2681 45 -2623
rect -45 -2727 -23 -2681
rect 23 -2727 45 -2681
rect -45 -2785 45 -2727
rect -45 -2831 -23 -2785
rect 23 -2831 45 -2785
rect -45 -2889 45 -2831
rect -45 -2935 -23 -2889
rect 23 -2935 45 -2889
rect -45 -2993 45 -2935
rect -45 -3039 -23 -2993
rect 23 -3039 45 -2993
rect -45 -3097 45 -3039
rect -45 -3143 -23 -3097
rect 23 -3143 45 -3097
rect -45 -3201 45 -3143
rect -45 -3247 -23 -3201
rect 23 -3247 45 -3201
rect -45 -3305 45 -3247
rect -45 -3351 -23 -3305
rect 23 -3351 45 -3305
rect -45 -3409 45 -3351
rect -45 -3455 -23 -3409
rect 23 -3455 45 -3409
rect -45 -3513 45 -3455
rect -45 -3559 -23 -3513
rect 23 -3559 45 -3513
rect -45 -3617 45 -3559
rect -45 -3663 -23 -3617
rect 23 -3663 45 -3617
rect -45 -3721 45 -3663
rect -45 -3767 -23 -3721
rect 23 -3767 45 -3721
rect -45 -3825 45 -3767
rect -45 -3871 -23 -3825
rect 23 -3871 45 -3825
rect -45 -3929 45 -3871
rect -45 -3975 -23 -3929
rect 23 -3975 45 -3929
rect -45 -4033 45 -3975
rect -45 -4079 -23 -4033
rect 23 -4079 45 -4033
rect -45 -4137 45 -4079
rect -45 -4183 -23 -4137
rect 23 -4183 45 -4137
rect -45 -4241 45 -4183
rect -45 -4287 -23 -4241
rect 23 -4287 45 -4241
rect -45 -4345 45 -4287
rect -45 -4391 -23 -4345
rect 23 -4391 45 -4345
rect -45 -4449 45 -4391
rect -45 -4495 -23 -4449
rect 23 -4495 45 -4449
rect -45 -4553 45 -4495
rect -45 -4599 -23 -4553
rect 23 -4599 45 -4553
rect -45 -4657 45 -4599
rect -45 -4703 -23 -4657
rect 23 -4703 45 -4657
rect -45 -4761 45 -4703
rect -45 -4807 -23 -4761
rect 23 -4807 45 -4761
rect -45 -4865 45 -4807
rect -45 -4911 -23 -4865
rect 23 -4911 45 -4865
rect -45 -4969 45 -4911
rect -45 -5015 -23 -4969
rect 23 -5015 45 -4969
rect -45 -5073 45 -5015
rect -45 -5119 -23 -5073
rect 23 -5119 45 -5073
rect -45 -5177 45 -5119
rect -45 -5223 -23 -5177
rect 23 -5223 45 -5177
rect -45 -5281 45 -5223
rect -45 -5327 -23 -5281
rect 23 -5327 45 -5281
rect -45 -5385 45 -5327
rect -45 -5431 -23 -5385
rect 23 -5431 45 -5385
rect -45 -5489 45 -5431
rect -45 -5535 -23 -5489
rect 23 -5535 45 -5489
rect -45 -5593 45 -5535
rect -45 -5639 -23 -5593
rect 23 -5639 45 -5593
rect -45 -5697 45 -5639
rect -45 -5743 -23 -5697
rect 23 -5743 45 -5697
rect -45 -5801 45 -5743
rect -45 -5847 -23 -5801
rect 23 -5847 45 -5801
rect -45 -5905 45 -5847
rect -45 -5951 -23 -5905
rect 23 -5951 45 -5905
rect -45 -6009 45 -5951
rect -45 -6055 -23 -6009
rect 23 -6055 45 -6009
rect -45 -6113 45 -6055
rect -45 -6159 -23 -6113
rect 23 -6159 45 -6113
rect -45 -6217 45 -6159
rect -45 -6263 -23 -6217
rect 23 -6263 45 -6217
rect -45 -6321 45 -6263
rect -45 -6367 -23 -6321
rect 23 -6367 45 -6321
rect -45 -6425 45 -6367
rect -45 -6471 -23 -6425
rect 23 -6471 45 -6425
rect -45 -6529 45 -6471
rect -45 -6575 -23 -6529
rect 23 -6575 45 -6529
rect -45 -6633 45 -6575
rect -45 -6679 -23 -6633
rect 23 -6679 45 -6633
rect -45 -6737 45 -6679
rect -45 -6783 -23 -6737
rect 23 -6783 45 -6737
rect -45 -6805 45 -6783
<< nsubdiffcont >>
rect -23 6737 23 6783
rect -23 6633 23 6679
rect -23 6529 23 6575
rect -23 6425 23 6471
rect -23 6321 23 6367
rect -23 6217 23 6263
rect -23 6113 23 6159
rect -23 6009 23 6055
rect -23 5905 23 5951
rect -23 5801 23 5847
rect -23 5697 23 5743
rect -23 5593 23 5639
rect -23 5489 23 5535
rect -23 5385 23 5431
rect -23 5281 23 5327
rect -23 5177 23 5223
rect -23 5073 23 5119
rect -23 4969 23 5015
rect -23 4865 23 4911
rect -23 4761 23 4807
rect -23 4657 23 4703
rect -23 4553 23 4599
rect -23 4449 23 4495
rect -23 4345 23 4391
rect -23 4241 23 4287
rect -23 4137 23 4183
rect -23 4033 23 4079
rect -23 3929 23 3975
rect -23 3825 23 3871
rect -23 3721 23 3767
rect -23 3617 23 3663
rect -23 3513 23 3559
rect -23 3409 23 3455
rect -23 3305 23 3351
rect -23 3201 23 3247
rect -23 3097 23 3143
rect -23 2993 23 3039
rect -23 2889 23 2935
rect -23 2785 23 2831
rect -23 2681 23 2727
rect -23 2577 23 2623
rect -23 2473 23 2519
rect -23 2369 23 2415
rect -23 2265 23 2311
rect -23 2161 23 2207
rect -23 2057 23 2103
rect -23 1953 23 1999
rect -23 1849 23 1895
rect -23 1745 23 1791
rect -23 1641 23 1687
rect -23 1537 23 1583
rect -23 1433 23 1479
rect -23 1329 23 1375
rect -23 1225 23 1271
rect -23 1121 23 1167
rect -23 1017 23 1063
rect -23 913 23 959
rect -23 809 23 855
rect -23 705 23 751
rect -23 601 23 647
rect -23 497 23 543
rect -23 393 23 439
rect -23 289 23 335
rect -23 185 23 231
rect -23 81 23 127
rect -23 -23 23 23
rect -23 -127 23 -81
rect -23 -231 23 -185
rect -23 -335 23 -289
rect -23 -439 23 -393
rect -23 -543 23 -497
rect -23 -647 23 -601
rect -23 -751 23 -705
rect -23 -855 23 -809
rect -23 -959 23 -913
rect -23 -1063 23 -1017
rect -23 -1167 23 -1121
rect -23 -1271 23 -1225
rect -23 -1375 23 -1329
rect -23 -1479 23 -1433
rect -23 -1583 23 -1537
rect -23 -1687 23 -1641
rect -23 -1791 23 -1745
rect -23 -1895 23 -1849
rect -23 -1999 23 -1953
rect -23 -2103 23 -2057
rect -23 -2207 23 -2161
rect -23 -2311 23 -2265
rect -23 -2415 23 -2369
rect -23 -2519 23 -2473
rect -23 -2623 23 -2577
rect -23 -2727 23 -2681
rect -23 -2831 23 -2785
rect -23 -2935 23 -2889
rect -23 -3039 23 -2993
rect -23 -3143 23 -3097
rect -23 -3247 23 -3201
rect -23 -3351 23 -3305
rect -23 -3455 23 -3409
rect -23 -3559 23 -3513
rect -23 -3663 23 -3617
rect -23 -3767 23 -3721
rect -23 -3871 23 -3825
rect -23 -3975 23 -3929
rect -23 -4079 23 -4033
rect -23 -4183 23 -4137
rect -23 -4287 23 -4241
rect -23 -4391 23 -4345
rect -23 -4495 23 -4449
rect -23 -4599 23 -4553
rect -23 -4703 23 -4657
rect -23 -4807 23 -4761
rect -23 -4911 23 -4865
rect -23 -5015 23 -4969
rect -23 -5119 23 -5073
rect -23 -5223 23 -5177
rect -23 -5327 23 -5281
rect -23 -5431 23 -5385
rect -23 -5535 23 -5489
rect -23 -5639 23 -5593
rect -23 -5743 23 -5697
rect -23 -5847 23 -5801
rect -23 -5951 23 -5905
rect -23 -6055 23 -6009
rect -23 -6159 23 -6113
rect -23 -6263 23 -6217
rect -23 -6367 23 -6321
rect -23 -6471 23 -6425
rect -23 -6575 23 -6529
rect -23 -6679 23 -6633
rect -23 -6783 23 -6737
<< metal1 >>
rect -34 6783 34 6794
rect -34 6737 -23 6783
rect 23 6737 34 6783
rect -34 6679 34 6737
rect -34 6633 -23 6679
rect 23 6633 34 6679
rect -34 6575 34 6633
rect -34 6529 -23 6575
rect 23 6529 34 6575
rect -34 6471 34 6529
rect -34 6425 -23 6471
rect 23 6425 34 6471
rect -34 6367 34 6425
rect -34 6321 -23 6367
rect 23 6321 34 6367
rect -34 6263 34 6321
rect -34 6217 -23 6263
rect 23 6217 34 6263
rect -34 6159 34 6217
rect -34 6113 -23 6159
rect 23 6113 34 6159
rect -34 6055 34 6113
rect -34 6009 -23 6055
rect 23 6009 34 6055
rect -34 5951 34 6009
rect -34 5905 -23 5951
rect 23 5905 34 5951
rect -34 5847 34 5905
rect -34 5801 -23 5847
rect 23 5801 34 5847
rect -34 5743 34 5801
rect -34 5697 -23 5743
rect 23 5697 34 5743
rect -34 5639 34 5697
rect -34 5593 -23 5639
rect 23 5593 34 5639
rect -34 5535 34 5593
rect -34 5489 -23 5535
rect 23 5489 34 5535
rect -34 5431 34 5489
rect -34 5385 -23 5431
rect 23 5385 34 5431
rect -34 5327 34 5385
rect -34 5281 -23 5327
rect 23 5281 34 5327
rect -34 5223 34 5281
rect -34 5177 -23 5223
rect 23 5177 34 5223
rect -34 5119 34 5177
rect -34 5073 -23 5119
rect 23 5073 34 5119
rect -34 5015 34 5073
rect -34 4969 -23 5015
rect 23 4969 34 5015
rect -34 4911 34 4969
rect -34 4865 -23 4911
rect 23 4865 34 4911
rect -34 4807 34 4865
rect -34 4761 -23 4807
rect 23 4761 34 4807
rect -34 4703 34 4761
rect -34 4657 -23 4703
rect 23 4657 34 4703
rect -34 4599 34 4657
rect -34 4553 -23 4599
rect 23 4553 34 4599
rect -34 4495 34 4553
rect -34 4449 -23 4495
rect 23 4449 34 4495
rect -34 4391 34 4449
rect -34 4345 -23 4391
rect 23 4345 34 4391
rect -34 4287 34 4345
rect -34 4241 -23 4287
rect 23 4241 34 4287
rect -34 4183 34 4241
rect -34 4137 -23 4183
rect 23 4137 34 4183
rect -34 4079 34 4137
rect -34 4033 -23 4079
rect 23 4033 34 4079
rect -34 3975 34 4033
rect -34 3929 -23 3975
rect 23 3929 34 3975
rect -34 3871 34 3929
rect -34 3825 -23 3871
rect 23 3825 34 3871
rect -34 3767 34 3825
rect -34 3721 -23 3767
rect 23 3721 34 3767
rect -34 3663 34 3721
rect -34 3617 -23 3663
rect 23 3617 34 3663
rect -34 3559 34 3617
rect -34 3513 -23 3559
rect 23 3513 34 3559
rect -34 3455 34 3513
rect -34 3409 -23 3455
rect 23 3409 34 3455
rect -34 3351 34 3409
rect -34 3305 -23 3351
rect 23 3305 34 3351
rect -34 3247 34 3305
rect -34 3201 -23 3247
rect 23 3201 34 3247
rect -34 3143 34 3201
rect -34 3097 -23 3143
rect 23 3097 34 3143
rect -34 3039 34 3097
rect -34 2993 -23 3039
rect 23 2993 34 3039
rect -34 2935 34 2993
rect -34 2889 -23 2935
rect 23 2889 34 2935
rect -34 2831 34 2889
rect -34 2785 -23 2831
rect 23 2785 34 2831
rect -34 2727 34 2785
rect -34 2681 -23 2727
rect 23 2681 34 2727
rect -34 2623 34 2681
rect -34 2577 -23 2623
rect 23 2577 34 2623
rect -34 2519 34 2577
rect -34 2473 -23 2519
rect 23 2473 34 2519
rect -34 2415 34 2473
rect -34 2369 -23 2415
rect 23 2369 34 2415
rect -34 2311 34 2369
rect -34 2265 -23 2311
rect 23 2265 34 2311
rect -34 2207 34 2265
rect -34 2161 -23 2207
rect 23 2161 34 2207
rect -34 2103 34 2161
rect -34 2057 -23 2103
rect 23 2057 34 2103
rect -34 1999 34 2057
rect -34 1953 -23 1999
rect 23 1953 34 1999
rect -34 1895 34 1953
rect -34 1849 -23 1895
rect 23 1849 34 1895
rect -34 1791 34 1849
rect -34 1745 -23 1791
rect 23 1745 34 1791
rect -34 1687 34 1745
rect -34 1641 -23 1687
rect 23 1641 34 1687
rect -34 1583 34 1641
rect -34 1537 -23 1583
rect 23 1537 34 1583
rect -34 1479 34 1537
rect -34 1433 -23 1479
rect 23 1433 34 1479
rect -34 1375 34 1433
rect -34 1329 -23 1375
rect 23 1329 34 1375
rect -34 1271 34 1329
rect -34 1225 -23 1271
rect 23 1225 34 1271
rect -34 1167 34 1225
rect -34 1121 -23 1167
rect 23 1121 34 1167
rect -34 1063 34 1121
rect -34 1017 -23 1063
rect 23 1017 34 1063
rect -34 959 34 1017
rect -34 913 -23 959
rect 23 913 34 959
rect -34 855 34 913
rect -34 809 -23 855
rect 23 809 34 855
rect -34 751 34 809
rect -34 705 -23 751
rect 23 705 34 751
rect -34 647 34 705
rect -34 601 -23 647
rect 23 601 34 647
rect -34 543 34 601
rect -34 497 -23 543
rect 23 497 34 543
rect -34 439 34 497
rect -34 393 -23 439
rect 23 393 34 439
rect -34 335 34 393
rect -34 289 -23 335
rect 23 289 34 335
rect -34 231 34 289
rect -34 185 -23 231
rect 23 185 34 231
rect -34 127 34 185
rect -34 81 -23 127
rect 23 81 34 127
rect -34 23 34 81
rect -34 -23 -23 23
rect 23 -23 34 23
rect -34 -81 34 -23
rect -34 -127 -23 -81
rect 23 -127 34 -81
rect -34 -185 34 -127
rect -34 -231 -23 -185
rect 23 -231 34 -185
rect -34 -289 34 -231
rect -34 -335 -23 -289
rect 23 -335 34 -289
rect -34 -393 34 -335
rect -34 -439 -23 -393
rect 23 -439 34 -393
rect -34 -497 34 -439
rect -34 -543 -23 -497
rect 23 -543 34 -497
rect -34 -601 34 -543
rect -34 -647 -23 -601
rect 23 -647 34 -601
rect -34 -705 34 -647
rect -34 -751 -23 -705
rect 23 -751 34 -705
rect -34 -809 34 -751
rect -34 -855 -23 -809
rect 23 -855 34 -809
rect -34 -913 34 -855
rect -34 -959 -23 -913
rect 23 -959 34 -913
rect -34 -1017 34 -959
rect -34 -1063 -23 -1017
rect 23 -1063 34 -1017
rect -34 -1121 34 -1063
rect -34 -1167 -23 -1121
rect 23 -1167 34 -1121
rect -34 -1225 34 -1167
rect -34 -1271 -23 -1225
rect 23 -1271 34 -1225
rect -34 -1329 34 -1271
rect -34 -1375 -23 -1329
rect 23 -1375 34 -1329
rect -34 -1433 34 -1375
rect -34 -1479 -23 -1433
rect 23 -1479 34 -1433
rect -34 -1537 34 -1479
rect -34 -1583 -23 -1537
rect 23 -1583 34 -1537
rect -34 -1641 34 -1583
rect -34 -1687 -23 -1641
rect 23 -1687 34 -1641
rect -34 -1745 34 -1687
rect -34 -1791 -23 -1745
rect 23 -1791 34 -1745
rect -34 -1849 34 -1791
rect -34 -1895 -23 -1849
rect 23 -1895 34 -1849
rect -34 -1953 34 -1895
rect -34 -1999 -23 -1953
rect 23 -1999 34 -1953
rect -34 -2057 34 -1999
rect -34 -2103 -23 -2057
rect 23 -2103 34 -2057
rect -34 -2161 34 -2103
rect -34 -2207 -23 -2161
rect 23 -2207 34 -2161
rect -34 -2265 34 -2207
rect -34 -2311 -23 -2265
rect 23 -2311 34 -2265
rect -34 -2369 34 -2311
rect -34 -2415 -23 -2369
rect 23 -2415 34 -2369
rect -34 -2473 34 -2415
rect -34 -2519 -23 -2473
rect 23 -2519 34 -2473
rect -34 -2577 34 -2519
rect -34 -2623 -23 -2577
rect 23 -2623 34 -2577
rect -34 -2681 34 -2623
rect -34 -2727 -23 -2681
rect 23 -2727 34 -2681
rect -34 -2785 34 -2727
rect -34 -2831 -23 -2785
rect 23 -2831 34 -2785
rect -34 -2889 34 -2831
rect -34 -2935 -23 -2889
rect 23 -2935 34 -2889
rect -34 -2993 34 -2935
rect -34 -3039 -23 -2993
rect 23 -3039 34 -2993
rect -34 -3097 34 -3039
rect -34 -3143 -23 -3097
rect 23 -3143 34 -3097
rect -34 -3201 34 -3143
rect -34 -3247 -23 -3201
rect 23 -3247 34 -3201
rect -34 -3305 34 -3247
rect -34 -3351 -23 -3305
rect 23 -3351 34 -3305
rect -34 -3409 34 -3351
rect -34 -3455 -23 -3409
rect 23 -3455 34 -3409
rect -34 -3513 34 -3455
rect -34 -3559 -23 -3513
rect 23 -3559 34 -3513
rect -34 -3617 34 -3559
rect -34 -3663 -23 -3617
rect 23 -3663 34 -3617
rect -34 -3721 34 -3663
rect -34 -3767 -23 -3721
rect 23 -3767 34 -3721
rect -34 -3825 34 -3767
rect -34 -3871 -23 -3825
rect 23 -3871 34 -3825
rect -34 -3929 34 -3871
rect -34 -3975 -23 -3929
rect 23 -3975 34 -3929
rect -34 -4033 34 -3975
rect -34 -4079 -23 -4033
rect 23 -4079 34 -4033
rect -34 -4137 34 -4079
rect -34 -4183 -23 -4137
rect 23 -4183 34 -4137
rect -34 -4241 34 -4183
rect -34 -4287 -23 -4241
rect 23 -4287 34 -4241
rect -34 -4345 34 -4287
rect -34 -4391 -23 -4345
rect 23 -4391 34 -4345
rect -34 -4449 34 -4391
rect -34 -4495 -23 -4449
rect 23 -4495 34 -4449
rect -34 -4553 34 -4495
rect -34 -4599 -23 -4553
rect 23 -4599 34 -4553
rect -34 -4657 34 -4599
rect -34 -4703 -23 -4657
rect 23 -4703 34 -4657
rect -34 -4761 34 -4703
rect -34 -4807 -23 -4761
rect 23 -4807 34 -4761
rect -34 -4865 34 -4807
rect -34 -4911 -23 -4865
rect 23 -4911 34 -4865
rect -34 -4969 34 -4911
rect -34 -5015 -23 -4969
rect 23 -5015 34 -4969
rect -34 -5073 34 -5015
rect -34 -5119 -23 -5073
rect 23 -5119 34 -5073
rect -34 -5177 34 -5119
rect -34 -5223 -23 -5177
rect 23 -5223 34 -5177
rect -34 -5281 34 -5223
rect -34 -5327 -23 -5281
rect 23 -5327 34 -5281
rect -34 -5385 34 -5327
rect -34 -5431 -23 -5385
rect 23 -5431 34 -5385
rect -34 -5489 34 -5431
rect -34 -5535 -23 -5489
rect 23 -5535 34 -5489
rect -34 -5593 34 -5535
rect -34 -5639 -23 -5593
rect 23 -5639 34 -5593
rect -34 -5697 34 -5639
rect -34 -5743 -23 -5697
rect 23 -5743 34 -5697
rect -34 -5801 34 -5743
rect -34 -5847 -23 -5801
rect 23 -5847 34 -5801
rect -34 -5905 34 -5847
rect -34 -5951 -23 -5905
rect 23 -5951 34 -5905
rect -34 -6009 34 -5951
rect -34 -6055 -23 -6009
rect 23 -6055 34 -6009
rect -34 -6113 34 -6055
rect -34 -6159 -23 -6113
rect 23 -6159 34 -6113
rect -34 -6217 34 -6159
rect -34 -6263 -23 -6217
rect 23 -6263 34 -6217
rect -34 -6321 34 -6263
rect -34 -6367 -23 -6321
rect 23 -6367 34 -6321
rect -34 -6425 34 -6367
rect -34 -6471 -23 -6425
rect 23 -6471 34 -6425
rect -34 -6529 34 -6471
rect -34 -6575 -23 -6529
rect 23 -6575 34 -6529
rect -34 -6633 34 -6575
rect -34 -6679 -23 -6633
rect 23 -6679 34 -6633
rect -34 -6737 34 -6679
rect -34 -6783 -23 -6737
rect 23 -6783 34 -6737
rect -34 -6794 34 -6783
<< end >>
