magic
tech gf180mcuC
magscale 1 10
timestamp 1692171811
<< nwell >>
rect -762 -1220 762 1220
<< pmos >>
rect -588 840 -532 1090
rect -428 840 -372 1090
rect -268 840 -212 1090
rect -108 840 -52 1090
rect 52 840 108 1090
rect 212 840 268 1090
rect 372 840 428 1090
rect 532 840 588 1090
rect -588 454 -532 704
rect -428 454 -372 704
rect -268 454 -212 704
rect -108 454 -52 704
rect 52 454 108 704
rect 212 454 268 704
rect 372 454 428 704
rect 532 454 588 704
rect -588 68 -532 318
rect -428 68 -372 318
rect -268 68 -212 318
rect -108 68 -52 318
rect 52 68 108 318
rect 212 68 268 318
rect 372 68 428 318
rect 532 68 588 318
rect -588 -318 -532 -68
rect -428 -318 -372 -68
rect -268 -318 -212 -68
rect -108 -318 -52 -68
rect 52 -318 108 -68
rect 212 -318 268 -68
rect 372 -318 428 -68
rect 532 -318 588 -68
rect -588 -704 -532 -454
rect -428 -704 -372 -454
rect -268 -704 -212 -454
rect -108 -704 -52 -454
rect 52 -704 108 -454
rect 212 -704 268 -454
rect 372 -704 428 -454
rect 532 -704 588 -454
rect -588 -1090 -532 -840
rect -428 -1090 -372 -840
rect -268 -1090 -212 -840
rect -108 -1090 -52 -840
rect 52 -1090 108 -840
rect 212 -1090 268 -840
rect 372 -1090 428 -840
rect 532 -1090 588 -840
<< pdiff >>
rect -676 1077 -588 1090
rect -676 853 -663 1077
rect -617 853 -588 1077
rect -676 840 -588 853
rect -532 1077 -428 1090
rect -532 853 -503 1077
rect -457 853 -428 1077
rect -532 840 -428 853
rect -372 1077 -268 1090
rect -372 853 -343 1077
rect -297 853 -268 1077
rect -372 840 -268 853
rect -212 1077 -108 1090
rect -212 853 -183 1077
rect -137 853 -108 1077
rect -212 840 -108 853
rect -52 1077 52 1090
rect -52 853 -23 1077
rect 23 853 52 1077
rect -52 840 52 853
rect 108 1077 212 1090
rect 108 853 137 1077
rect 183 853 212 1077
rect 108 840 212 853
rect 268 1077 372 1090
rect 268 853 297 1077
rect 343 853 372 1077
rect 268 840 372 853
rect 428 1077 532 1090
rect 428 853 457 1077
rect 503 853 532 1077
rect 428 840 532 853
rect 588 1077 676 1090
rect 588 853 617 1077
rect 663 853 676 1077
rect 588 840 676 853
rect -676 691 -588 704
rect -676 467 -663 691
rect -617 467 -588 691
rect -676 454 -588 467
rect -532 691 -428 704
rect -532 467 -503 691
rect -457 467 -428 691
rect -532 454 -428 467
rect -372 691 -268 704
rect -372 467 -343 691
rect -297 467 -268 691
rect -372 454 -268 467
rect -212 691 -108 704
rect -212 467 -183 691
rect -137 467 -108 691
rect -212 454 -108 467
rect -52 691 52 704
rect -52 467 -23 691
rect 23 467 52 691
rect -52 454 52 467
rect 108 691 212 704
rect 108 467 137 691
rect 183 467 212 691
rect 108 454 212 467
rect 268 691 372 704
rect 268 467 297 691
rect 343 467 372 691
rect 268 454 372 467
rect 428 691 532 704
rect 428 467 457 691
rect 503 467 532 691
rect 428 454 532 467
rect 588 691 676 704
rect 588 467 617 691
rect 663 467 676 691
rect 588 454 676 467
rect -676 305 -588 318
rect -676 81 -663 305
rect -617 81 -588 305
rect -676 68 -588 81
rect -532 305 -428 318
rect -532 81 -503 305
rect -457 81 -428 305
rect -532 68 -428 81
rect -372 305 -268 318
rect -372 81 -343 305
rect -297 81 -268 305
rect -372 68 -268 81
rect -212 305 -108 318
rect -212 81 -183 305
rect -137 81 -108 305
rect -212 68 -108 81
rect -52 305 52 318
rect -52 81 -23 305
rect 23 81 52 305
rect -52 68 52 81
rect 108 305 212 318
rect 108 81 137 305
rect 183 81 212 305
rect 108 68 212 81
rect 268 305 372 318
rect 268 81 297 305
rect 343 81 372 305
rect 268 68 372 81
rect 428 305 532 318
rect 428 81 457 305
rect 503 81 532 305
rect 428 68 532 81
rect 588 305 676 318
rect 588 81 617 305
rect 663 81 676 305
rect 588 68 676 81
rect -676 -81 -588 -68
rect -676 -305 -663 -81
rect -617 -305 -588 -81
rect -676 -318 -588 -305
rect -532 -81 -428 -68
rect -532 -305 -503 -81
rect -457 -305 -428 -81
rect -532 -318 -428 -305
rect -372 -81 -268 -68
rect -372 -305 -343 -81
rect -297 -305 -268 -81
rect -372 -318 -268 -305
rect -212 -81 -108 -68
rect -212 -305 -183 -81
rect -137 -305 -108 -81
rect -212 -318 -108 -305
rect -52 -81 52 -68
rect -52 -305 -23 -81
rect 23 -305 52 -81
rect -52 -318 52 -305
rect 108 -81 212 -68
rect 108 -305 137 -81
rect 183 -305 212 -81
rect 108 -318 212 -305
rect 268 -81 372 -68
rect 268 -305 297 -81
rect 343 -305 372 -81
rect 268 -318 372 -305
rect 428 -81 532 -68
rect 428 -305 457 -81
rect 503 -305 532 -81
rect 428 -318 532 -305
rect 588 -81 676 -68
rect 588 -305 617 -81
rect 663 -305 676 -81
rect 588 -318 676 -305
rect -676 -467 -588 -454
rect -676 -691 -663 -467
rect -617 -691 -588 -467
rect -676 -704 -588 -691
rect -532 -467 -428 -454
rect -532 -691 -503 -467
rect -457 -691 -428 -467
rect -532 -704 -428 -691
rect -372 -467 -268 -454
rect -372 -691 -343 -467
rect -297 -691 -268 -467
rect -372 -704 -268 -691
rect -212 -467 -108 -454
rect -212 -691 -183 -467
rect -137 -691 -108 -467
rect -212 -704 -108 -691
rect -52 -467 52 -454
rect -52 -691 -23 -467
rect 23 -691 52 -467
rect -52 -704 52 -691
rect 108 -467 212 -454
rect 108 -691 137 -467
rect 183 -691 212 -467
rect 108 -704 212 -691
rect 268 -467 372 -454
rect 268 -691 297 -467
rect 343 -691 372 -467
rect 268 -704 372 -691
rect 428 -467 532 -454
rect 428 -691 457 -467
rect 503 -691 532 -467
rect 428 -704 532 -691
rect 588 -467 676 -454
rect 588 -691 617 -467
rect 663 -691 676 -467
rect 588 -704 676 -691
rect -676 -853 -588 -840
rect -676 -1077 -663 -853
rect -617 -1077 -588 -853
rect -676 -1090 -588 -1077
rect -532 -853 -428 -840
rect -532 -1077 -503 -853
rect -457 -1077 -428 -853
rect -532 -1090 -428 -1077
rect -372 -853 -268 -840
rect -372 -1077 -343 -853
rect -297 -1077 -268 -853
rect -372 -1090 -268 -1077
rect -212 -853 -108 -840
rect -212 -1077 -183 -853
rect -137 -1077 -108 -853
rect -212 -1090 -108 -1077
rect -52 -853 52 -840
rect -52 -1077 -23 -853
rect 23 -1077 52 -853
rect -52 -1090 52 -1077
rect 108 -853 212 -840
rect 108 -1077 137 -853
rect 183 -1077 212 -853
rect 108 -1090 212 -1077
rect 268 -853 372 -840
rect 268 -1077 297 -853
rect 343 -1077 372 -853
rect 268 -1090 372 -1077
rect 428 -853 532 -840
rect 428 -1077 457 -853
rect 503 -1077 532 -853
rect 428 -1090 532 -1077
rect 588 -853 676 -840
rect 588 -1077 617 -853
rect 663 -1077 676 -853
rect 588 -1090 676 -1077
<< pdiffc >>
rect -663 853 -617 1077
rect -503 853 -457 1077
rect -343 853 -297 1077
rect -183 853 -137 1077
rect -23 853 23 1077
rect 137 853 183 1077
rect 297 853 343 1077
rect 457 853 503 1077
rect 617 853 663 1077
rect -663 467 -617 691
rect -503 467 -457 691
rect -343 467 -297 691
rect -183 467 -137 691
rect -23 467 23 691
rect 137 467 183 691
rect 297 467 343 691
rect 457 467 503 691
rect 617 467 663 691
rect -663 81 -617 305
rect -503 81 -457 305
rect -343 81 -297 305
rect -183 81 -137 305
rect -23 81 23 305
rect 137 81 183 305
rect 297 81 343 305
rect 457 81 503 305
rect 617 81 663 305
rect -663 -305 -617 -81
rect -503 -305 -457 -81
rect -343 -305 -297 -81
rect -183 -305 -137 -81
rect -23 -305 23 -81
rect 137 -305 183 -81
rect 297 -305 343 -81
rect 457 -305 503 -81
rect 617 -305 663 -81
rect -663 -691 -617 -467
rect -503 -691 -457 -467
rect -343 -691 -297 -467
rect -183 -691 -137 -467
rect -23 -691 23 -467
rect 137 -691 183 -467
rect 297 -691 343 -467
rect 457 -691 503 -467
rect 617 -691 663 -467
rect -663 -1077 -617 -853
rect -503 -1077 -457 -853
rect -343 -1077 -297 -853
rect -183 -1077 -137 -853
rect -23 -1077 23 -853
rect 137 -1077 183 -853
rect 297 -1077 343 -853
rect 457 -1077 503 -853
rect 617 -1077 663 -853
<< polysilicon >>
rect -588 1090 -532 1134
rect -428 1090 -372 1134
rect -268 1090 -212 1134
rect -108 1090 -52 1134
rect 52 1090 108 1134
rect 212 1090 268 1134
rect 372 1090 428 1134
rect 532 1090 588 1134
rect -588 796 -532 840
rect -428 796 -372 840
rect -268 796 -212 840
rect -108 796 -52 840
rect 52 796 108 840
rect 212 796 268 840
rect 372 796 428 840
rect 532 796 588 840
rect -588 704 -532 748
rect -428 704 -372 748
rect -268 704 -212 748
rect -108 704 -52 748
rect 52 704 108 748
rect 212 704 268 748
rect 372 704 428 748
rect 532 704 588 748
rect -588 410 -532 454
rect -428 410 -372 454
rect -268 410 -212 454
rect -108 410 -52 454
rect 52 410 108 454
rect 212 410 268 454
rect 372 410 428 454
rect 532 410 588 454
rect -588 318 -532 362
rect -428 318 -372 362
rect -268 318 -212 362
rect -108 318 -52 362
rect 52 318 108 362
rect 212 318 268 362
rect 372 318 428 362
rect 532 318 588 362
rect -588 24 -532 68
rect -428 24 -372 68
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect 372 24 428 68
rect 532 24 588 68
rect -588 -68 -532 -24
rect -428 -68 -372 -24
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect 372 -68 428 -24
rect 532 -68 588 -24
rect -588 -362 -532 -318
rect -428 -362 -372 -318
rect -268 -362 -212 -318
rect -108 -362 -52 -318
rect 52 -362 108 -318
rect 212 -362 268 -318
rect 372 -362 428 -318
rect 532 -362 588 -318
rect -588 -454 -532 -410
rect -428 -454 -372 -410
rect -268 -454 -212 -410
rect -108 -454 -52 -410
rect 52 -454 108 -410
rect 212 -454 268 -410
rect 372 -454 428 -410
rect 532 -454 588 -410
rect -588 -748 -532 -704
rect -428 -748 -372 -704
rect -268 -748 -212 -704
rect -108 -748 -52 -704
rect 52 -748 108 -704
rect 212 -748 268 -704
rect 372 -748 428 -704
rect 532 -748 588 -704
rect -588 -840 -532 -796
rect -428 -840 -372 -796
rect -268 -840 -212 -796
rect -108 -840 -52 -796
rect 52 -840 108 -796
rect 212 -840 268 -796
rect 372 -840 428 -796
rect 532 -840 588 -796
rect -588 -1134 -532 -1090
rect -428 -1134 -372 -1090
rect -268 -1134 -212 -1090
rect -108 -1134 -52 -1090
rect 52 -1134 108 -1090
rect 212 -1134 268 -1090
rect 372 -1134 428 -1090
rect 532 -1134 588 -1090
<< metal1 >>
rect -663 1077 -617 1088
rect -663 842 -617 853
rect -503 1077 -457 1088
rect -503 842 -457 853
rect -343 1077 -297 1088
rect -343 842 -297 853
rect -183 1077 -137 1088
rect -183 842 -137 853
rect -23 1077 23 1088
rect -23 842 23 853
rect 137 1077 183 1088
rect 137 842 183 853
rect 297 1077 343 1088
rect 297 842 343 853
rect 457 1077 503 1088
rect 457 842 503 853
rect 617 1077 663 1088
rect 617 842 663 853
rect -663 691 -617 702
rect -663 456 -617 467
rect -503 691 -457 702
rect -503 456 -457 467
rect -343 691 -297 702
rect -343 456 -297 467
rect -183 691 -137 702
rect -183 456 -137 467
rect -23 691 23 702
rect -23 456 23 467
rect 137 691 183 702
rect 137 456 183 467
rect 297 691 343 702
rect 297 456 343 467
rect 457 691 503 702
rect 457 456 503 467
rect 617 691 663 702
rect 617 456 663 467
rect -663 305 -617 316
rect -663 70 -617 81
rect -503 305 -457 316
rect -503 70 -457 81
rect -343 305 -297 316
rect -343 70 -297 81
rect -183 305 -137 316
rect -183 70 -137 81
rect -23 305 23 316
rect -23 70 23 81
rect 137 305 183 316
rect 137 70 183 81
rect 297 305 343 316
rect 297 70 343 81
rect 457 305 503 316
rect 457 70 503 81
rect 617 305 663 316
rect 617 70 663 81
rect -663 -81 -617 -70
rect -663 -316 -617 -305
rect -503 -81 -457 -70
rect -503 -316 -457 -305
rect -343 -81 -297 -70
rect -343 -316 -297 -305
rect -183 -81 -137 -70
rect -183 -316 -137 -305
rect -23 -81 23 -70
rect -23 -316 23 -305
rect 137 -81 183 -70
rect 137 -316 183 -305
rect 297 -81 343 -70
rect 297 -316 343 -305
rect 457 -81 503 -70
rect 457 -316 503 -305
rect 617 -81 663 -70
rect 617 -316 663 -305
rect -663 -467 -617 -456
rect -663 -702 -617 -691
rect -503 -467 -457 -456
rect -503 -702 -457 -691
rect -343 -467 -297 -456
rect -343 -702 -297 -691
rect -183 -467 -137 -456
rect -183 -702 -137 -691
rect -23 -467 23 -456
rect -23 -702 23 -691
rect 137 -467 183 -456
rect 137 -702 183 -691
rect 297 -467 343 -456
rect 297 -702 343 -691
rect 457 -467 503 -456
rect 457 -702 503 -691
rect 617 -467 663 -456
rect 617 -702 663 -691
rect -663 -853 -617 -842
rect -663 -1088 -617 -1077
rect -503 -853 -457 -842
rect -503 -1088 -457 -1077
rect -343 -853 -297 -842
rect -343 -1088 -297 -1077
rect -183 -853 -137 -842
rect -183 -1088 -137 -1077
rect -23 -853 23 -842
rect -23 -1088 23 -1077
rect 137 -853 183 -842
rect 137 -1088 183 -1077
rect 297 -853 343 -842
rect 297 -1088 343 -1077
rect 457 -853 503 -842
rect 457 -1088 503 -1077
rect 617 -853 663 -842
rect 617 -1088 663 -1077
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 1.25 l 0.280 m 6 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
