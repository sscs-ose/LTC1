magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1045 1045 1045
<< metal1 >>
rect -45 39 45 45
rect -45 -39 -39 39
rect 39 -39 45 39
rect -45 -45 45 -39
<< via1 >>
rect -39 -39 39 39
<< metal2 >>
rect -45 39 45 45
rect -45 -39 -39 39
rect 39 -39 45 39
rect -45 -45 45 -39
<< end >>
