magic
tech gf180mcuC
magscale 1 10
timestamp 1714460654
<< nwell >>
rect -4713 20 -2077 2476
rect -4713 -160 -1992 20
<< nsubdiff >>
rect -3418 35 -3337 55
rect -3418 24 -3281 35
rect -3437 -34 -3281 24
rect -3437 -115 -3406 -34
rect -3325 -115 -3281 -34
rect -3437 -130 -3281 -115
<< nsubdiffcont >>
rect -3406 -115 -3325 -34
<< metal1 >>
rect -4496 2754 -4336 2772
rect -4496 2700 -4454 2754
rect -4387 2700 -4336 2754
rect -4496 2665 -4336 2700
rect -2336 2771 -2176 2782
rect -2336 2712 -2302 2771
rect -2222 2712 -2176 2771
rect -2336 2692 -2176 2712
rect -4497 2400 -4336 2408
rect -4497 2330 -4478 2400
rect -4352 2330 -4336 2400
rect -4497 2307 -4336 2330
rect -4257 2306 -3857 2409
rect -3777 2306 -3377 2409
rect -3297 2306 -2897 2409
rect -2817 2306 -2417 2409
rect -2337 2395 -2176 2408
rect -2337 2328 -2304 2395
rect -2202 2328 -2176 2395
rect -2337 2306 -2176 2328
rect -4497 204 -4097 307
rect -4017 204 -3617 307
rect -3537 204 -3137 307
rect -3057 204 -2657 307
rect -2577 205 -2177 308
rect -3488 -34 -3189 -23
rect -3488 -115 -3406 -34
rect -3325 -115 -3189 -34
rect -3488 -141 -3189 -115
<< via1 >>
rect -4454 2700 -4387 2754
rect -2302 2712 -2222 2771
rect -4478 2330 -4352 2400
rect -2304 2328 -2202 2395
<< metal2 >>
rect -4496 2754 -4336 2772
rect -4496 2700 -4454 2754
rect -4387 2700 -4336 2754
rect -4496 2408 -4336 2700
rect -2336 2771 -2176 2782
rect -2336 2712 -2302 2771
rect -2222 2712 -2176 2771
rect -2336 2408 -2176 2712
rect -4497 2400 -4336 2408
rect -4497 2330 -4478 2400
rect -4352 2330 -4336 2400
rect -4497 2307 -4336 2330
rect -4496 2306 -4336 2307
rect -2337 2395 -2176 2408
rect -2337 2328 -2304 2395
rect -2202 2328 -2176 2395
rect -2337 2306 -2176 2328
use ppolyf_u_3D7VPB  ppolyf_u_3D7VPB_0
timestamp 1714140926
transform 1 0 -3337 0 1 1306
box -1376 -1318 1376 1318
<< labels >>
flabel nsubdiffcont -3366 -71 -3366 -71 0 FreeSans 640 0 0 0 VDD
port 2 nsew
flabel via1 -2266 2743 -2266 2743 0 FreeSans 640 0 0 0 B
port 3 nsew
flabel via1 -4421 2728 -4421 2728 0 FreeSans 640 0 0 0 A
port 4 nsew
<< end >>
