magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2468 2045 2468
<< psubdiff >>
rect -45 446 45 468
rect -45 -446 -23 446
rect 23 -446 45 446
rect -45 -468 45 -446
<< psubdiffcont >>
rect -23 -446 23 446
<< metal1 >>
rect -34 446 34 457
rect -34 -446 -23 446
rect 23 -446 34 446
rect -34 -457 34 -446
<< end >>
