magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -6839 2045 6839
<< psubdiff >>
rect -45 4817 45 4839
rect -45 -4817 -23 4817
rect 23 -4817 45 4817
rect -45 -4839 45 -4817
<< psubdiffcont >>
rect -23 -4817 23 4817
<< metal1 >>
rect -34 4817 34 4828
rect -34 -4817 -23 4817
rect 23 -4817 34 4817
rect -34 -4828 34 -4817
<< end >>
