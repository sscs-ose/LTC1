* NGSPICE file created from CLK_div_96_mag_flat.ext - technology: gf180mcuC

.subckt CLK_div_96_mag_flat VDD VSS Vdiv96 RST CLK
X0 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_2.OUT VDD.t263 VDD.t262 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 JK_FF_mag_2.QB JK_FF_mag_2.nand2_mag_4.IN2 VDD.t171 VDD.t170 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 VDD JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_1.IN2 VDD.t356 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t362 VDD.t361 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X4 VDD JK_FF_mag_0.Q JK_FF_mag_2.nand3_mag_0.OUT VDD.t293 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X5 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t360 VDD.t359 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X6 VDD JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_1.IN2 VDD.t191 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X7 VDD JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t76 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X8 JK_FF_mag_4.nand3_mag_0.OUT CLK.t0 VDD.t299 VDD.t298 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X9 VDD CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t47 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X10 JK_FF_mag_4.nand2_mag_1.IN2 JK_FF_mag_4.nand2_mag_3.IN1 VDD.t221 VDD.t220 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 VDD JK_FF_mag_5.QB JK_FF_mag_5.nand3_mag_0.OUT VDD.t314 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X12 a_3934_1448# VDD.t368 VSS.t85 VSS.t84 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X13 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t144 VSS.t143 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X14 a_1426_417# JK_FF_mag_0.nand3_mag_2.OUT VSS.t39 VSS.t38 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X15 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT a_1432_1558# VSS.t5 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_4697_2604# VSS.t228 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X17 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.QB a_4094_1448# VSS.t213 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X18 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand3_mag_1.OUT VDD.t20 VDD.t19 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 VDD JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_0.OUT VDD.t157 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 a_3973_2604# JK_FF_mag_3.Q a_3813_2604# VSS.t55 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X21 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 VDD.t24 VDD.t23 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X22 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 VDD.t39 VDD.t38 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X23 a_7745_351# JK_FF_mag_3.nand3_mag_2.OUT VSS.t174 VSS.t173 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X24 a_5418_5266# CLK.t1 a_5258_5266# VSS.t13 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X25 a_4094_1448# JK_FF_mag_0.Q a_3934_1448# VSS.t188 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X26 JK_FF_mag_4.nand2_mag_4.IN2 JK_FF_mag_4.nand2_mag_3.IN1 VDD.t219 VDD.t218 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X27 a_4130_5266# JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand2_mag_1.IN2 VSS.t140 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X28 a_2147_3060# JK_FF_mag_5.QB JK_FF_mag_5.nand3_mag_0.OUT VSS.t205 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X29 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0 a_8842_2648# VSS.t120 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X30 VDD JK_FF_mag_0.QB JK_FF_mag_0.Q VDD.t174 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X31 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT VDD.t32 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X32 JK_FF_mag_4.nand3_mag_1.OUT RST.t0 VDD.t169 VDD.t168 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 JK_FF_mag_4.QB JK_FF_mag_4.Q.t3 VDD.t274 VDD.t273 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X34 JK_FF_mag_4.nand3_mag_2.OUT CLK.t2 VDD.t250 VDD.t249 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 a_5258_5266# JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_0.OUT VSS.t107 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X36 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB VDD.t173 VDD.t172 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X37 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t28 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X38 JK_FF_mag_3.nand3_mag_2.OUT VDD.t118 VDD.t120 VDD.t119 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X39 JK_FF_mag_0.Q JK_FF_mag_0.nand2_mag_1.IN2 VDD.t53 VDD.t52 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X40 JK_FF_mag_3.QB JK_FF_mag_3.Q a_9033_395# VSS.t54 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X41 VSS CLK.t3 JK_FF_mag_4.nand2_mag_3.IN1 VSS.t10 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X42 VDD JK_FF_mag_2.Q JK_FF_mag_2.QB VDD.t207 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X43 a_3976_6363# JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand2_mag_4.IN2 VSS.t139 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X44 VDD JK_FF_mag_4.Q.t4 JK_FF_mag_4.nand3_mag_2.OUT VDD.t275 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X45 VDD JK_FF_mag_5.Q.t3 JK_FF_mag_0.nand3_mag_0.OUT VDD.t130 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X46 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 a_4812_351# VSS.t22 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X47 VDD JK_FF_mag_0.Q JK_FF_mag_0.QB VDD.t290 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X48 a_4700_6363# RST.t1 a_4540_6363# VSS.t111 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X49 a_5107_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t227 VSS.t226 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X50 a_3412_6363# JK_FF_mag_4.Q.t5 JK_FF_mag_4.QB VSS.t191 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X51 a_5424_6363# CLK.t4 a_5264_6363# VSS.t9 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X52 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_5.Q.t4 VDD.t134 VDD.t133 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X53 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 a_5825_2648# VSS.t37 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X54 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t115 VDD.t117 VDD.t116 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X55 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t234 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X56 VDD JK_FF_mag_2.QB JK_FF_mag_2.Q VDD.t328 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X57 a_5940_395# JK_FF_mag_2.nand2_mag_4.IN2 VSS.t113 VSS.t112 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X58 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 VDD.t182 VDD.t181 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X59 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t248 VDD.t247 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X60 VDD JK_FF_mag_5.Q.t5 JK_FF_mag_0.nand3_mag_2.OUT VDD.t317 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X61 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t55 VDD.t54 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X62 JK_FF_mag_3.nand3_mag_0.OUT VDD.t112 VDD.t114 VDD.t113 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X63 a_7021_351# VDD.t369 VSS.t83 VSS.t82 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X64 VDD JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_4.IN2 VDD.t188 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X65 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_2.OUT VDD.t223 VDD.t222 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB a_868_1514# VSS.t115 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X67 VDD JK_FF_mag_3.QB JK_FF_mag_3.Q VDD.t270 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X68 a_5264_6363# JK_FF_mag_4.Q.t6 JK_FF_mag_4.nand3_mag_2.OUT VSS.t192 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X69 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X70 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.QB VDD.t269 VDD.t268 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X71 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_0.OUT VDD.t217 VDD.t216 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X72 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t141 VDD.t140 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X73 a_6830_2604# VDD.t370 VSS.t81 VSS.t80 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X74 JK_FF_mag_2.Q JK_FF_mag_2.nand2_mag_1.IN2 VDD.t297 VDD.t296 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X75 VDD VDD.t108 JK_FF_mag_5.nand3_mag_2.OUT VDD.t109 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X76 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 a_6990_2604# VSS.t119 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X77 a_7554_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t43 VSS.t42 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X78 a_868_1514# JK_FF_mag_5.Q.t6 a_708_1514# VSS.t206 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X79 JK_FF_mag_3.Q JK_FF_mag_3.nand2_mag_1.IN2 VDD.t143 VDD.t142 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X80 VDD JK_FF_mag_2.Q JK_FF_mag_3.nand3_mag_0.OUT VDD.t204 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 a_2714_461# JK_FF_mag_0.nand2_mag_4.IN2 VSS.t149 VSS.t148 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X82 VDD JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X83 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand3_mag_1.IN1 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X84 a_8469_395# JK_FF_mag_3.nand3_mag_1.OUT VSS.t19 VSS.t18 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X85 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t137 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X86 VDD RST.t2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t165 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X87 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand3_mag_1.IN1 VDD.t154 VDD.t153 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X88 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_3.Q VDD.t72 VDD.t71 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X89 VDD JK_FF_mag_2.Q JK_FF_mag_3.nand3_mag_2.OUT VDD.t201 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X90 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand3_mag_1.OUT VDD.t339 VDD.t338 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X91 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_0.Q VSS.t187 VSS.t186 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X92 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t105 VDD.t107 VDD.t106 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X93 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t127 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X94 a_862_417# JK_FF_mag_5.Q.t7 a_702_417# VSS.t14 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X95 a_1996_1558# JK_FF_mag_0.nand3_mag_1.IN1 VSS.t32 VSS.t31 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X96 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 VDD.t46 VDD.t45 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X97 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t238 VDD.t237 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X98 a_4652_351# JK_FF_mag_2.nand3_mag_2.OUT VSS.t142 VSS.t141 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X99 a_7027_1448# VDD.t372 VSS.t79 VSS.t78 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X100 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.Q VSS.t132 VSS.t131 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X101 VSS VDD.t373 a_2313_4157# VSS.t75 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X102 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VDD.t161 VDD.t160 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X103 a_6996_3701# JK_FF_mag_3.Q a_6836_3701# VSS.t53 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X104 a_2150_461# JK_FF_mag_0.nand3_mag_1.OUT VSS.t4 VSS.t3 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X105 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.QB a_7187_1448# VSS.t179 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X106 JK_FF_mag_0.Q JK_FF_mag_0.QB a_2560_1558# VSS.t114 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X107 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t136 VDD.t135 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X108 a_1432_1558# JK_FF_mag_0.nand3_mag_0.OUT VSS.t26 VSS.t25 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X109 a_4697_2604# RST.t3 a_4537_2604# VSS.t222 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X110 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t231 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X111 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t282 VDD.t281 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X112 a_3813_2604# VDD.t374 VSS.t74 VSS.t73 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X113 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_1996_1558# VSS.t24 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X114 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 a_3973_2604# VSS.t36 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X115 JK_FF_mag_2.nand3_mag_2.OUT VDD.t102 VDD.t104 VDD.t103 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X116 a_7187_1448# JK_FF_mag_2.Q a_7027_1448# VSS.t130 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X117 a_2560_1558# JK_FF_mag_0.nand2_mag_1.IN2 VSS.t41 VSS.t40 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X118 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t4 a_6996_3701# VSS.t223 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X119 VDD RST.t4 JK_FF_mag_0.nand3_mag_1.OUT VDD.t347 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X120 VDD JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t68 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X121 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_8278_2648# VSS.t151 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X122 JK_FF_mag_2.QB JK_FF_mag_2.Q a_5940_395# VSS.t129 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X123 a_8842_2648# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t163 VSS.t162 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X124 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.Q VDD.t289 VDD.t288 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X125 VDD JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand2_mag_4.IN2 VDD.t365 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X126 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t278 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X127 a_7181_351# JK_FF_mag_2.Q a_7021_351# VSS.t128 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X128 VDD JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand3_mag_1.OUT VDD.t259 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X129 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_3.Q VDD.t67 VDD.t66 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X130 VDD RST.t5 JK_FF_mag_3.nand3_mag_1.OUT VDD.t121 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X131 a_8278_2648# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t94 VSS.t93 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X132 a_3979_3701# JK_FF_mag_3.Q a_3819_3701# VSS.t52 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X133 VDD JK_FF_mag_5.nand3_mag_0.OUT JK_FF_mag_5.nand3_mag_1.IN1 VDD.t241 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X134 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand2_mag_3.IN1 a_8469_395# VSS.t125 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X135 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_1.OUT a_4658_1492# VSS.t219 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X136 VSS JK_FF_mag_4.nand3_mag_1.OUT a_3976_6363# VSS.t230 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X137 VDD VDD.t98 JK_FF_mag_5.nand3_mag_0.OUT VDD.t99 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X138 JK_FF_mag_0.nand3_mag_0.OUT VDD.t95 VDD.t97 VDD.t96 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X139 a_3928_351# VDD.t376 VSS.t72 VSS.t71 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X140 a_4540_6363# JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand3_mag_1.OUT VSS.t172 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X141 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_7560_3745# VSS.t92 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X142 VDD JK_FF_mag_4.Q.t7 JK_FF_mag_5.nand2_mag_3.IN1 VDD.t300 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X143 a_1586_417# RST.t6 a_1426_417# VSS.t86 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X144 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.Q VDD.t65 VDD.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X145 VDD JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_4.IN2 VDD.t353 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X146 VDD JK_FF_mag_5.nand3_mag_1.IN1 JK_FF_mag_5.nand2_mag_1.IN2 VDD.t309 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X147 JK_FF_mag_5.nand3_mag_1.IN1 JK_FF_mag_5.nand3_mag_1.OUT VDD.t150 VDD.t149 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X148 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_1.OUT a_7751_1492# VSS.t17 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X149 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.Q a_862_417# VSS.t185 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X150 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5261_2648# VSS.t88 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X151 a_5825_2648# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t153 VSS.t152 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X152 a_4658_1492# JK_FF_mag_2.nand3_mag_0.OUT VSS.t122 VSS.t121 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X153 VDD JK_FF_mag_5.nand3_mag_2.OUT JK_FF_mag_5.nand3_mag_1.OUT VDD.t244 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X154 VSS JK_FF_mag_5.nand3_mag_0.OUT a_1583_3060# VSS.t156 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X155 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_5.Q.t8 VSS.t16 VSS.t15 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X156 a_7560_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t90 VSS.t89 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X157 a_7905_351# RST.t7 a_7745_351# VSS.t133 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X158 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_3.IN1 a_5222_1492# VSS.t225 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X159 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_8124_3745# VSS.t150 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X160 VSS VDD.t377 a_2307_3060# VSS.t68 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X161 VDD JK_FF_mag_5.nand2_mag_1.IN2 JK_FF_mag_5.Q.t0 VDD.t226 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X162 a_5376_395# JK_FF_mag_2.nand3_mag_1.OUT VSS.t218 VSS.t217 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X163 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand2_mag_3.IN1 a_8315_1492# VSS.t124 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X164 VDD CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t42 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X165 VSS JK_FF_mag_5.nand3_mag_1.IN1 a_1019_3060# VSS.t201 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X166 VSS JK_FF_mag_4.Q.t8 JK_FF_mag_5.nand2_mag_3.IN1 VSS.t193 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X167 a_5261_2648# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t182 VSS.t181 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X168 JK_FF_mag_5.nand3_mag_1.OUT RST.t8 VDD.t211 VDD.t210 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X169 a_1583_3060# JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_5.nand3_mag_1.IN1 VSS.t102 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X170 VDD JK_FF_mag_0.Q JK_FF_mag_2.nand3_mag_2.OUT VDD.t285 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t37 VDD.t36 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X172 JK_FF_mag_5.nand3_mag_2.OUT JK_FF_mag_4.Q.t9 VDD.t265 VDD.t264 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X173 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_3.Q VSS.t51 VSS.t50 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X174 a_708_1514# VDD.t378 VSS.t67 VSS.t66 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X175 VSS JK_FF_mag_5.nand3_mag_2.OUT a_1589_4157# VSS.t159 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X176 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.Q a_7181_351# VSS.t49 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X177 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_3.Q VDD.t63 VDD.t62 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X178 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 VDD.t41 VDD.t40 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X179 VDD CLK_div_3_mag_0.JK_FF_mag_1.K.t5 CLK_div_3_mag_0.Q0 VDD.t350 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X180 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_4543_3745# VSS.t180 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X181 VSS JK_FF_mag_5.nand2_mag_1.IN2 a_455_3060# VSS.t145 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X182 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t323 VDD.t322 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X183 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 VDD.t152 VDD.t151 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X184 VDD JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_5.nand2_mag_4.IN2 VDD.t146 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X185 a_1589_4157# RST.t9 a_1429_4157# VSS.t8 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X186 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0 a_8245_5080# VDD.t180 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X187 a_2313_4157# JK_FF_mag_4.Q.t10 a_2153_4157# VSS.t175 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X188 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t321 VDD.t320 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X189 a_6836_3701# CLK_div_3_mag_0.Q1 VSS.t35 VSS.t34 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X190 VDD JK_FF_mag_5.nand2_mag_4.IN2 JK_FF_mag_5.QB VDD.t251 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X191 JK_FF_mag_5.nand2_mag_4.IN2 JK_FF_mag_5.nand2_mag_3.IN1 VDD.t343 VDD.t342 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X192 a_4537_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t210 VSS.t209 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X193 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 a_1586_417# VSS.t30 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X194 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t334 VDD.t333 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X195 a_4088_351# JK_FF_mag_0.Q a_3928_351# VSS.t184 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X196 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t332 VDD.t331 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X197 VDD RST.t10 JK_FF_mag_2.nand3_mag_1.OUT VDD.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X198 VSS JK_FF_mag_5.nand3_mag_1.OUT a_865_4157# VSS.t99 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X199 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_3.Q VSS.t48 VSS.t47 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X200 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VDD.t215 VDD.t214 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X201 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X202 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 a_7905_351# VSS.t105 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X203 VSS CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t116 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X204 VSS JK_FF_mag_5.nand2_mag_4.IN2 a_301_4157# VSS.t164 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X205 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t9 VDD.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X206 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t145 VDD.t144 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X207 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_7714_2604# VSS.t216 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X208 VDD JK_FF_mag_4.nand2_mag_1.IN2 JK_FF_mag_4.Q.t0 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X209 a_865_4157# JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.nand2_mag_4.IN2 VSS.t221 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X210 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_3.IN1 a_5376_395# VSS.t224 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X211 JK_FF_mag_0.QB JK_FF_mag_0.Q a_2714_461# VSS.t183 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X212 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q1 a_7272_4844# VSS.t33 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X213 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t124 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X214 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.Q VDD.t200 VDD.t199 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X215 VDD JK_FF_mag_4.nand3_mag_0.OUT JK_FF_mag_4.nand3_mag_1.IN1 VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X216 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t255 VDD.t254 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X217 a_3819_3701# CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS.t136 VSS.t135 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X218 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB a_3979_3701# VSS.t7 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X219 JK_FF_mag_4.Q JK_FF_mag_4.QB VDD.t156 VDD.t155 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X220 JK_FF_mag_2.Q JK_FF_mag_2.QB a_5786_1492# VSS.t212 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X221 VDD VDD.t91 JK_FF_mag_4.nand3_mag_0.OUT VDD.t92 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X222 a_7272_4844# JK_FF_mag_3.Q VSS.t46 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X223 a_4812_351# RST.t11 a_4652_351# VSS.t123 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X224 VDD JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand2_mag_1.IN2 VDD.t256 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X225 VDD CLK.t5 JK_FF_mag_4.nand2_mag_3.IN1 VDD.t344 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X226 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 a_8688_3745# VSS.t91 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X227 JK_FF_mag_5.nand3_mag_0.OUT JK_FF_mag_4.Q.t11 VDD.t325 VDD.t324 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X228 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_4.IN2 VDD.t267 VDD.t266 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X229 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_4.IN2 VDD.t230 VDD.t229 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X230 JK_FF_mag_3.Q JK_FF_mag_3.QB a_8879_1492# VSS.t178 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X231 VSS JK_FF_mag_4.nand2_mag_1.IN2 a_3566_5266# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X232 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand3_mag_1.OUT VDD.t364 VDD.t363 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X233 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t155 VSS.t154 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X234 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_2150_461# VSS.t23 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X235 a_7751_1492# JK_FF_mag_3.nand3_mag_0.OUT VSS.t138 VSS.t137 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X236 a_5786_1492# JK_FF_mag_2.nand2_mag_1.IN2 VSS.t190 VSS.t189 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X237 VSS JK_FF_mag_4.nand3_mag_0.OUT a_4694_5266# VSS.t27 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X238 a_8688_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t208 VSS.t207 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X239 JK_FF_mag_5.nand2_mag_1.IN2 JK_FF_mag_5.nand2_mag_3.IN1 VDD.t341 VDD.t340 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X240 a_8879_1492# JK_FF_mag_3.nand2_mag_1.IN2 VSS.t96 VSS.t95 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X241 a_3566_5266# JK_FF_mag_4.QB JK_FF_mag_4.Q.t1 VSS.t106 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X242 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t225 VDD.t224 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X243 JK_FF_mag_0.nand3_mag_2.OUT VDD.t88 VDD.t90 VDD.t89 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X244 a_5222_1492# JK_FF_mag_2.nand3_mag_1.IN1 VSS.t21 VSS.t20 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X245 VSS VDD.t380 a_5418_5266# VSS.t63 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X246 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.Q a_4088_351# VSS.t127 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X247 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t7 VDD.t6 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X248 VSS JK_FF_mag_4.nand3_mag_1.IN1 a_4130_5266# VSS.t169 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X249 a_4694_5266# JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_1.IN1 VSS.t229 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X250 a_8124_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t215 VSS.t214 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X251 a_2307_3060# JK_FF_mag_4.Q.t12 a_2147_3060# VSS.t211 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X252 JK_FF_mag_5.Q JK_FF_mag_5.QB VDD.t313 VDD.t312 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X253 a_8315_1492# JK_FF_mag_3.nand3_mag_1.IN1 VSS.t104 VSS.t103 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X254 VDD JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X255 VDD JK_FF_mag_4.nand3_mag_2.OUT JK_FF_mag_4.nand3_mag_1.OUT VDD.t162 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X256 VDD JK_FF_mag_5.nand3_mag_1.IN1 JK_FF_mag_5.nand3_mag_1.OUT VDD.t306 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X257 VDD JK_FF_mag_4.nand2_mag_4.IN2 JK_FF_mag_4.QB VDD.t303 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X258 VDD VDD.t84 JK_FF_mag_4.nand3_mag_2.OUT VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X259 VDD JK_FF_mag_5.Q.t9 JK_FF_mag_5.nand3_mag_2.OUT VDD.t194 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X260 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB a_5671_3745# VSS.t6 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X261 a_1019_3060# JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.nand2_mag_1.IN2 VSS.t220 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X262 a_4543_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t98 VSS.t97 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X263 a_455_3060# JK_FF_mag_5.QB JK_FF_mag_5.Q.t2 VSS.t204 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X264 Vdiv96 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t80 VDD.t79 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X265 VSS JK_FF_mag_4.nand3_mag_2.OUT a_4700_6363# VSS.t108 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X266 a_1429_4157# JK_FF_mag_5.nand3_mag_1.IN1 JK_FF_mag_5.nand3_mag_1.OUT VSS.t200 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X267 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_5107_3745# VSS.t87 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X268 a_5671_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t168 VSS.t167 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X269 a_702_417# VDD.t382 VSS.t61 VSS.t60 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X270 VSS JK_FF_mag_4.nand2_mag_4.IN2 a_3412_6363# VSS.t196 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X271 Vdiv96 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t57 VSS.t56 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X272 VSS VDD.t383 a_5424_6363# VSS.t58 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X273 a_8245_5080# CLK_div_3_mag_0.or_2_mag_0.IN2 VDD.t240 VDD.t239 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X274 a_2153_4157# JK_FF_mag_5.Q.t10 JK_FF_mag_5.nand3_mag_2.OUT VSS.t126 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X275 JK_FF_mag_5.QB JK_FF_mag_5.Q.t11 VDD.t213 VDD.t212 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X276 VDD JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t58 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X277 VDD JK_FF_mag_3.Q JK_FF_mag_3.QB VDD.t56 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X278 VDD CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VDD.t177 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X279 VDD RST.t12 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t185 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X280 VDD JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 VDD.t335 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X281 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_0.Q VDD.t284 VDD.t283 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X282 JK_FF_mag_2.nand3_mag_0.OUT VDD.t81 VDD.t83 VDD.t82 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X283 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT VDD.t51 VDD.t50 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X284 VDD JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 VDD.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X285 a_6990_2604# JK_FF_mag_3.Q a_6830_2604# VSS.t44 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X286 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.QB VDD.t327 VDD.t326 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X287 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.Q VDD.t198 VDD.t197 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X288 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_0.OUT VDD.t184 VDD.t183 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X289 a_9033_395# JK_FF_mag_3.nand2_mag_4.IN2 VSS.t177 VSS.t176 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X290 a_301_4157# JK_FF_mag_5.Q.t12 JK_FF_mag_5.QB VSS.t134 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X291 a_7714_2604# RST.t13 a_7554_2604# VSS.t199 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
R0 VDD.n113 VDD.n112 11185.2
R1 VDD.n307 VDD.n306 2201.41
R2 VDD.t356 VDD.t296 961.905
R3 VDD.t183 VDD.t326 961.905
R4 VDD.t234 VDD.t247 765.152
R5 VDD.t331 VDD.t140 765.152
R6 VDD.t181 VDD.t54 765.152
R7 VDD.t320 VDD.t231 765.152
R8 VDD.t137 VDD.t333 765.152
R9 VDD.t135 VDD.t160 765.152
R10 VDD.t127 VDD.t237 765.152
R11 VDD.t359 VDD.t281 765.152
R12 VDD.t45 VDD.t322 765.152
R13 VDD.t244 VDD.t194 765.152
R14 VDD.t306 VDD.t146 765.152
R15 VDD.t251 VDD.t342 765.152
R16 VDD.t25 VDD.t229 765.152
R17 VDD.t36 VDD.t6 765.152
R18 VDD.t288 VDD.t50 765.152
R19 VDD.t142 VDD.t191 765.152
R20 VDD.t16 VDD.t153 765.152
R21 VDD.t216 VDD.t268 765.152
R22 VDD.t188 VDD.t266 765.152
R23 VDD.t151 VDD.t19 765.152
R24 VDD.t64 VDD.t262 765.152
R25 VDD.t353 VDD.t170 765.152
R26 VDD.t23 VDD.t338 765.152
R27 VDD.t199 VDD.t222 765.152
R28 VDD.t162 VDD.t275 765.152
R29 VDD.t259 VDD.t365 765.152
R30 VDD.t303 VDD.t218 765.152
R31 VDD.n112 VDD.t21 676.191
R32 VDD.n113 VDD.t82 485.714
R33 VDD VDD.n98 429.187
R34 VDD VDD.n293 427.092
R35 VDD.t283 VDD.n113 426.44
R36 VDD.n297 VDD 420.935
R37 VDD.n98 VDD.t113 386.365
R38 VDD.t326 VDD.t293 380.952
R39 VDD.t42 VDD.n297 378.788
R40 VDD.n305 VDD.t40 329.546
R41 VDD.n306 VDD.n305 324.075
R42 VDD.n297 VDD.t239 322.223
R43 VDD.n293 VDD.t180 320.635
R44 VDD.t185 VDD.t331 303.031
R45 VDD.t58 VDD.t181 303.031
R46 VDD.t160 VDD.t73 303.031
R47 VDD.t165 VDD.t359 303.031
R48 VDD.t76 VDD.t45 303.031
R49 VDD.t194 VDD.t264 303.031
R50 VDD.t210 VDD.t306 303.031
R51 VDD.t347 VDD.t36 303.031
R52 VDD.t317 VDD.t288 303.031
R53 VDD.t268 VDD.t204 303.031
R54 VDD.t121 VDD.t151 303.031
R55 VDD.t201 VDD.t64 303.031
R56 VDD.t13 VDD.t23 303.031
R57 VDD.t285 VDD.t199 303.031
R58 VDD.t275 VDD.t249 303.031
R59 VDD.t168 VDD.t259 303.031
R60 VDD.n112 VDD.t335 285.714
R61 VDD.n104 VDD.t328 242.857
R62 VDD.n105 VDD.t356 242.857
R63 VDD.t335 VDD.n111 242.857
R64 VDD.t293 VDD.n20 242.857
R65 VDD.t241 VDD.t38 239.583
R66 VDD.t309 VDD.t31 239.583
R67 VDD.t33 VDD.t361 235.35
R68 VDD.t256 VDD.t144 235.35
R69 VDD.n258 VDD.t177 193.183
R70 VDD.n260 VDD.t234 193.183
R71 VDD.n263 VDD.t185 193.183
R72 VDD.n266 VDD.t58 193.183
R73 VDD.n279 VDD.t350 193.183
R74 VDD.n285 VDD.t231 193.183
R75 VDD.n286 VDD.t137 193.183
R76 VDD.n304 VDD.t73 193.183
R77 VDD.n298 VDD.t42 193.183
R78 VDD.n9 VDD.t47 193.183
R79 VDD.n11 VDD.t127 193.183
R80 VDD.n14 VDD.t165 193.183
R81 VDD.n17 VDD.t76 193.183
R82 VDD.n191 VDD.t290 193.183
R83 VDD.n193 VDD.t25 193.183
R84 VDD.n196 VDD.t347 193.183
R85 VDD.n199 VDD.t317 193.183
R86 VDD.n85 VDD.t270 193.183
R87 VDD.n91 VDD.t191 193.183
R88 VDD.n92 VDD.t16 193.183
R89 VDD.n97 VDD.t204 193.183
R90 VDD.n59 VDD.t56 193.183
R91 VDD.n61 VDD.t188 193.183
R92 VDD.n64 VDD.t121 193.183
R93 VDD.n67 VDD.t201 193.183
R94 VDD.n26 VDD.t207 193.183
R95 VDD.n28 VDD.t353 193.183
R96 VDD.n31 VDD.t13 193.183
R97 VDD.n34 VDD.t285 193.183
R98 VDD.t264 VDD.n151 191.288
R99 VDD.n152 VDD.t210 191.288
R100 VDD.t342 VDD.n160 191.288
R101 VDD.n161 VDD.t212 191.288
R102 VDD.t249 VDD.n359 191.288
R103 VDD.n360 VDD.t168 191.288
R104 VDD.t218 VDD.n368 191.288
R105 VDD.n369 VDD.t273 191.288
R106 VDD.t174 VDD.t300 142.993
R107 VDD.t28 VDD.t324 142.993
R108 VDD.t130 VDD.t340 142.993
R109 VDD.t133 VDD.t312 142.993
R110 VDD.n296 VDD.t180 142.857
R111 VDD.t344 VDD.t10 140.465
R112 VDD.t298 VDD.t124 140.465
R113 VDD.t220 VDD.t68 140.465
R114 VDD.t296 VDD.n104 138.095
R115 VDD.n105 VDD.t21 138.095
R116 VDD.n111 VDD.t183 138.095
R117 VDD.t82 VDD.n20 138.095
R118 VDD.n305 VDD.t71 125.001
R119 VDD.n151 VDD.t109 111.743
R120 VDD.n152 VDD.t244 111.743
R121 VDD.n160 VDD.t146 111.743
R122 VDD.n161 VDD.t251 111.743
R123 VDD.n359 VDD.t85 111.743
R124 VDD.n360 VDD.t162 111.743
R125 VDD.n368 VDD.t365 111.743
R126 VDD.n369 VDD.t303 111.743
R127 VDD.t239 VDD.n296 111.112
R128 VDD.t247 VDD.n258 109.849
R129 VDD.t140 VDD.n260 109.849
R130 VDD.t54 VDD.n263 109.849
R131 VDD.n266 VDD.t116 109.849
R132 VDD.n279 VDD.t320 109.849
R133 VDD.t333 VDD.n285 109.849
R134 VDD.n286 VDD.t135 109.849
R135 VDD.t40 VDD.n304 109.849
R136 VDD.n298 VDD.t62 109.849
R137 VDD.t237 VDD.n9 109.849
R138 VDD.t281 VDD.n11 109.849
R139 VDD.t322 VDD.n14 109.849
R140 VDD.n17 VDD.t106 109.849
R141 VDD.t229 VDD.n191 109.849
R142 VDD.t6 VDD.n193 109.849
R143 VDD.t50 VDD.n196 109.849
R144 VDD.n199 VDD.t89 109.849
R145 VDD.n85 VDD.t142 109.849
R146 VDD.t153 VDD.n91 109.849
R147 VDD.n92 VDD.t216 109.849
R148 VDD.t113 VDD.n97 109.849
R149 VDD.t266 VDD.n59 109.849
R150 VDD.t19 VDD.n61 109.849
R151 VDD.t262 VDD.n64 109.849
R152 VDD.n67 VDD.t119 109.849
R153 VDD.t170 VDD.n26 109.849
R154 VDD.t338 VDD.n28 109.849
R155 VDD.t222 VDD.n31 109.849
R156 VDD.n34 VDD.t103 109.849
R157 VDD.n116 VDD.t174 96.5914
R158 VDD.n131 VDD.t130 96.5914
R159 VDD.t324 VDD.n118 95.6444
R160 VDD.t312 VDD.n133 95.6444
R161 VDD.n314 VDD.t10 94.8842
R162 VDD.n341 VDD.t68 94.8842
R163 VDD.n315 VDD.t298 93.954
R164 VDD.n342 VDD.t155 93.954
R165 VDD.t99 VDD.t52 88.0687
R166 VDD.n122 VDD.t314 88.0687
R167 VDD.n126 VDD.t149 88.0687
R168 VDD.t226 VDD.t96 88.0687
R169 VDD.t3 VDD.n124 87.1217
R170 VDD.t172 VDD.n128 87.1217
R171 VDD.t92 VDD.t254 86.5121
R172 VDD.n323 VDD.t157 86.5121
R173 VDD.n332 VDD.t363 86.5121
R174 VDD.t0 VDD.t214 86.5121
R175 VDD.n333 VDD.t8 85.5819
R176 VDD.n98 VDD.t197 59.702
R177 VDD.n293 VDD.t79 59.4064
R178 VDD.n297 VDD.t224 58.5371
R179 VDD.n118 VDD.t99 55.8717
R180 VDD.n124 VDD.t241 55.8717
R181 VDD.n128 VDD.t309 55.8717
R182 VDD.n133 VDD.t226 55.8717
R183 VDD.t52 VDD.n116 54.9247
R184 VDD.t38 VDD.n122 54.9247
R185 VDD.t31 VDD.n126 54.9247
R186 VDD.t96 VDD.n131 54.9247
R187 VDD.n315 VDD.t92 54.8842
R188 VDD.n324 VDD.t33 54.8842
R189 VDD.n333 VDD.t256 54.8842
R190 VDD.n342 VDD.t0 54.8842
R191 VDD.t254 VDD.n314 53.954
R192 VDD.t361 VDD.n323 53.954
R193 VDD.t144 VDD.n332 53.954
R194 VDD.t214 VDD.n341 53.954
R195 VDD.n225 VDD.t115 30.9379
R196 VDD.n140 VDD.t108 30.9379
R197 VDD.n142 VDD.t98 30.9379
R198 VDD.n200 VDD.t95 30.9379
R199 VDD.n202 VDD.t88 30.9379
R200 VDD.n69 VDD.t118 30.9379
R201 VDD.n68 VDD.t112 30.9379
R202 VDD.n35 VDD.t81 30.9379
R203 VDD.n36 VDD.t102 30.9379
R204 VDD.n350 VDD.t84 30.9379
R205 VDD.n352 VDD.t91 30.9379
R206 VDD.n231 VDD.t105 30.0062
R207 VDD.n225 VDD.t370 24.5101
R208 VDD.n140 VDD.t373 24.5101
R209 VDD.n142 VDD.t377 24.5101
R210 VDD.n200 VDD.t378 24.5101
R211 VDD.n202 VDD.t382 24.5101
R212 VDD.n69 VDD.t369 24.5101
R213 VDD.n68 VDD.t372 24.5101
R214 VDD.n35 VDD.t368 24.5101
R215 VDD.n36 VDD.t376 24.5101
R216 VDD.n350 VDD.t383 24.5101
R217 VDD.n352 VDD.t380 24.5101
R218 VDD.n230 VDD.t374 24.4392
R219 VDD VDD.t283 10.5649
R220 VDD.t314 VDD.t28 8.52323
R221 VDD.t149 VDD.t3 8.52323
R222 VDD.t340 VDD.t172 8.52323
R223 VDD.t124 VDD.t157 8.37259
R224 VDD.t363 VDD.t278 8.37259
R225 VDD.t8 VDD.t220 8.37259
R226 VDD VDD.t133 8.19444
R227 VDD VDD.t300 8.19444
R228 VDD VDD.t66 8.16097
R229 VDD.n267 VDD.n266 6.3005
R230 VDD.n270 VDD.n263 6.3005
R231 VDD.n273 VDD.n260 6.3005
R232 VDD.n276 VDD.n258 6.3005
R233 VDD.n287 VDD.n286 6.3005
R234 VDD.n285 VDD.n284 6.3005
R235 VDD.n280 VDD.n279 6.3005
R236 VDD.n296 VDD.n295 6.3005
R237 VDD.n299 VDD.n298 6.3005
R238 VDD.n304 VDD.n303 6.3005
R239 VDD.n306 VDD 6.3005
R240 VDD.n151 VDD.n150 6.3005
R241 VDD.n153 VDD.n152 6.3005
R242 VDD.n160 VDD.n159 6.3005
R243 VDD.n162 VDD.n161 6.3005
R244 VDD.n184 VDD.n118 6.3005
R245 VDD.n178 VDD.n124 6.3005
R246 VDD.n172 VDD.n128 6.3005
R247 VDD.n166 VDD.n133 6.3005
R248 VDD.n169 VDD.n131 6.3005
R249 VDD.n175 VDD.n126 6.3005
R250 VDD.n181 VDD.n122 6.3005
R251 VDD.n187 VDD.n116 6.3005
R252 VDD.n208 VDD.n199 6.3005
R253 VDD.n211 VDD.n196 6.3005
R254 VDD.n214 VDD.n193 6.3005
R255 VDD.n217 VDD.n191 6.3005
R256 VDD.n73 VDD.n67 6.3005
R257 VDD.n76 VDD.n64 6.3005
R258 VDD.n79 VDD.n61 6.3005
R259 VDD.n82 VDD.n59 6.3005
R260 VDD.n86 VDD.n85 6.3005
R261 VDD.n91 VDD.n90 6.3005
R262 VDD.n93 VDD.n92 6.3005
R263 VDD.n97 VDD.n96 6.3005
R264 VDD.n40 VDD.n34 6.3005
R265 VDD.n43 VDD.n31 6.3005
R266 VDD.n46 VDD.n28 6.3005
R267 VDD.n49 VDD.n26 6.3005
R268 VDD.n222 VDD.n20 6.3005
R269 VDD.n104 VDD.n103 6.3005
R270 VDD.n106 VDD.n105 6.3005
R271 VDD.n111 VDD.n110 6.3005
R272 VDD.n238 VDD.n17 6.3005
R273 VDD.n241 VDD.n14 6.3005
R274 VDD.n244 VDD.n11 6.3005
R275 VDD.n247 VDD.n9 6.3005
R276 VDD VDD.n307 6.3005
R277 VDD.n316 VDD.n315 6.3005
R278 VDD.n325 VDD.n324 6.3005
R279 VDD.n334 VDD.n333 6.3005
R280 VDD.n343 VDD.n342 6.3005
R281 VDD.n341 VDD.n340 6.3005
R282 VDD.n332 VDD.n331 6.3005
R283 VDD.n323 VDD.n322 6.3005
R284 VDD.n314 VDD.n313 6.3005
R285 VDD.n359 VDD.n358 6.3005
R286 VDD.n361 VDD.n360 6.3005
R287 VDD.n368 VDD.n367 6.3005
R288 VDD.n370 VDD.n369 6.3005
R289 VDD.n227 VDD.n226 5.63356
R290 VDD.n267 VDD.t117 5.213
R291 VDD.n308 VDD.n7 5.19407
R292 VDD.n310 VDD.n309 5.19167
R293 VDD.n288 VDD.t136 5.13287
R294 VDD.n254 VDD.n253 5.13287
R295 VDD.n283 VDD.t334 5.13287
R296 VDD.n282 VDD.n255 5.13287
R297 VDD.n281 VDD.t321 5.13287
R298 VDD.n278 VDD.n256 5.13287
R299 VDD.n269 VDD.t55 5.13287
R300 VDD.n272 VDD.t141 5.13287
R301 VDD.n274 VDD.n259 5.13287
R302 VDD.n275 VDD.t248 5.13287
R303 VDD.n277 VDD.n257 5.13287
R304 VDD.n300 VDD.t63 5.13287
R305 VDD.n291 VDD.n290 5.13287
R306 VDD.n301 VDD.t41 5.13287
R307 VDD.n146 VDD.n139 5.13287
R308 VDD.n138 VDD.n137 5.13287
R309 VDD.n155 VDD.n134 5.13287
R310 VDD.n158 VDD.t343 5.13287
R311 VDD.n157 VDD.n156 5.13287
R312 VDD.n163 VDD.t213 5.13287
R313 VDD.n207 VDD.t90 5.13287
R314 VDD.n210 VDD.t51 5.13287
R315 VDD.n213 VDD.t7 5.13287
R316 VDD.n215 VDD.n192 5.13287
R317 VDD.n216 VDD.t230 5.13287
R318 VDD.n218 VDD.n190 5.13287
R319 VDD.n51 VDD.t114 5.13287
R320 VDD.n94 VDD.t217 5.13287
R321 VDD.n55 VDD.n54 5.13287
R322 VDD.n89 VDD.t154 5.13287
R323 VDD.n88 VDD.n56 5.13287
R324 VDD.n87 VDD.t143 5.13287
R325 VDD.n84 VDD.n57 5.13287
R326 VDD.n72 VDD.t120 5.13287
R327 VDD.n75 VDD.t263 5.13287
R328 VDD.n78 VDD.t20 5.13287
R329 VDD.n80 VDD.n60 5.13287
R330 VDD.n81 VDD.t267 5.13287
R331 VDD.n83 VDD.n58 5.13287
R332 VDD.n39 VDD.t104 5.13287
R333 VDD.n42 VDD.t223 5.13287
R334 VDD.n45 VDD.t339 5.13287
R335 VDD.n47 VDD.n27 5.13287
R336 VDD.n48 VDD.t171 5.13287
R337 VDD.n50 VDD.n25 5.13287
R338 VDD.n221 VDD.t83 5.13287
R339 VDD.n109 VDD.t184 5.13287
R340 VDD.n108 VDD.n21 5.13287
R341 VDD.n107 VDD.t22 5.13287
R342 VDD.n23 VDD.n22 5.13287
R343 VDD.n102 VDD.t297 5.13287
R344 VDD.n101 VDD.n24 5.13287
R345 VDD.n240 VDD.t323 5.13287
R346 VDD.n243 VDD.t282 5.13287
R347 VDD.n245 VDD.n10 5.13287
R348 VDD.n246 VDD.t238 5.13287
R349 VDD.n248 VDD.n8 5.13287
R350 VDD.n312 VDD.n311 5.13287
R351 VDD.n320 VDD.n319 5.13287
R352 VDD.n327 VDD.t364 5.13287
R353 VDD.n329 VDD.n328 5.13287
R354 VDD.n336 VDD.t221 5.13287
R355 VDD.n339 VDD.n337 5.13287
R356 VDD.n338 VDD.t215 5.13287
R357 VDD.n330 VDD.t145 5.13287
R358 VDD.n326 VDD.n2 5.13287
R359 VDD.n321 VDD.t362 5.13287
R360 VDD.n317 VDD.n5 5.13287
R361 VDD.n6 VDD.t255 5.13287
R362 VDD.n354 VDD.n349 5.13287
R363 VDD.n348 VDD.n347 5.13287
R364 VDD.n363 VDD.n344 5.13287
R365 VDD.n366 VDD.t219 5.13287
R366 VDD.n365 VDD.n364 5.13287
R367 VDD.n371 VDD.t274 5.13287
R368 VDD.n372 VDD.t156 5.13287
R369 VDD.n186 VDD.n117 5.11708
R370 VDD.n179 VDD.n123 5.11708
R371 VDD.n176 VDD.t150 5.11708
R372 VDD.n173 VDD.n127 5.11708
R373 VDD.n170 VDD.t341 5.11708
R374 VDD.n168 VDD.n132 5.11708
R375 VDD.n165 VDD.t313 5.11708
R376 VDD.n167 VDD.t97 5.1155
R377 VDD.n174 VDD.t32 5.1155
R378 VDD.n177 VDD.n125 5.1155
R379 VDD.n180 VDD.t39 5.1155
R380 VDD.n183 VDD.n119 5.1155
R381 VDD.n185 VDD.t53 5.1155
R382 VDD.n188 VDD.n115 5.1155
R383 VDD VDD.t80 5.10321
R384 VDD VDD.t67 5.10312
R385 VDD.n292 VDD.t225 5.09407
R386 VDD.n189 VDD.n114 5.09407
R387 VDD.n220 VDD.t284 5.09407
R388 VDD.n99 VDD.t198 5.09407
R389 VDD.n250 VDD.t72 5.09264
R390 VDD.n164 VDD.t134 5.09264
R391 VDD.n237 VDD.t107 4.8755
R392 VDD.n294 VDD.t240 4.12326
R393 VDD.n143 VDD.n142 4.08796
R394 VDD VDD.n35 4.08442
R395 VDD.n70 VDD.n69 4.08323
R396 VDD.n351 VDD.n350 4.07925
R397 VDD.n37 VDD.n36 4.07855
R398 VDD.n141 VDD.n140 4.07362
R399 VDD.n201 VDD.n200 4.04647
R400 VDD VDD.n352 4.04611
R401 VDD VDD.n68 4.04234
R402 VDD.n203 VDD.n202 4.041
R403 VDD.n232 VDD.n231 3.61662
R404 VDD.n145 VDD.n144 3.13455
R405 VDD.n206 VDD.n201 3.01689
R406 VDD.n353 VDD 3.01101
R407 VDD.n38 VDD 2.99823
R408 VDD.n71 VDD 2.9975
R409 VDD.n145 VDD.n141 2.95902
R410 VDD.n353 VDD.n351 2.91542
R411 VDD.n71 VDD.n70 2.87793
R412 VDD.n38 VDD.n37 2.86761
R413 VDD.n289 VDD.n252 2.85787
R414 VDD.n268 VDD.n265 2.85787
R415 VDD.n271 VDD.n262 2.85787
R416 VDD.n149 VDD.n148 2.85787
R417 VDD.n154 VDD.n136 2.85787
R418 VDD.n209 VDD.n198 2.85787
R419 VDD.n212 VDD.n195 2.85787
R420 VDD.n95 VDD.n53 2.85787
R421 VDD.n74 VDD.n66 2.85787
R422 VDD.n77 VDD.n63 2.85787
R423 VDD.n41 VDD.n33 2.85787
R424 VDD.n44 VDD.n30 2.85787
R425 VDD.n223 VDD.n19 2.85787
R426 VDD.n239 VDD.n16 2.85787
R427 VDD.n242 VDD.n13 2.85787
R428 VDD.n318 VDD.n4 2.85787
R429 VDD.n335 VDD.n1 2.85787
R430 VDD.n357 VDD.n356 2.85787
R431 VDD.n362 VDD.n346 2.85787
R432 VDD.n206 VDD.n205 2.84443
R433 VDD.n182 VDD.n121 2.84208
R434 VDD.n171 VDD.n130 2.8405
R435 VDD.n227 VDD.n224 2.65604
R436 VDD.n252 VDD.t161 2.2755
R437 VDD.n252 VDD.n251 2.2755
R438 VDD.n265 VDD.t182 2.2755
R439 VDD.n265 VDD.n264 2.2755
R440 VDD.n262 VDD.t332 2.2755
R441 VDD.n262 VDD.n261 2.2755
R442 VDD.n121 VDD.t325 2.2755
R443 VDD.n121 VDD.n120 2.2755
R444 VDD.n148 VDD.t265 2.2755
R445 VDD.n148 VDD.n147 2.2755
R446 VDD.n136 VDD.t211 2.2755
R447 VDD.n136 VDD.n135 2.2755
R448 VDD.n130 VDD.t173 2.2755
R449 VDD.n130 VDD.n129 2.2755
R450 VDD.n198 VDD.t289 2.2755
R451 VDD.n198 VDD.n197 2.2755
R452 VDD.n195 VDD.t37 2.2755
R453 VDD.n195 VDD.n194 2.2755
R454 VDD.n53 VDD.t269 2.2755
R455 VDD.n53 VDD.n52 2.2755
R456 VDD.n66 VDD.t65 2.2755
R457 VDD.n66 VDD.n65 2.2755
R458 VDD.n63 VDD.t152 2.2755
R459 VDD.n63 VDD.n62 2.2755
R460 VDD.n33 VDD.t200 2.2755
R461 VDD.n33 VDD.n32 2.2755
R462 VDD.n30 VDD.t24 2.2755
R463 VDD.n30 VDD.n29 2.2755
R464 VDD.n19 VDD.t327 2.2755
R465 VDD.n19 VDD.n18 2.2755
R466 VDD.n16 VDD.t46 2.2755
R467 VDD.n16 VDD.n15 2.2755
R468 VDD.n13 VDD.t360 2.2755
R469 VDD.n13 VDD.n12 2.2755
R470 VDD.n4 VDD.t299 2.2755
R471 VDD.n4 VDD.n3 2.2755
R472 VDD.n1 VDD.t9 2.2755
R473 VDD.n1 VDD.n0 2.2755
R474 VDD.n356 VDD.t250 2.2755
R475 VDD.n356 VDD.n355 2.2755
R476 VDD.n346 VDD.t169 2.2755
R477 VDD.n346 VDD.n345 2.2755
R478 VDD.n207 VDD.n206 2.26792
R479 VDD.n354 VDD.n353 2.26734
R480 VDD.n39 VDD.n38 2.26618
R481 VDD.n72 VDD.n71 2.2656
R482 VDD.n146 VDD.n145 2.26502
R483 VDD.n226 VDD.n225 2.11318
R484 VDD.n307 VDD.t344 1.86097
R485 VDD.n229 VDD.n228 1.54785
R486 VDD.n228 VDD.n227 1.35532
R487 VDD.n278 VDD.n277 1.16167
R488 VDD.n84 VDD.n83 1.16167
R489 VDD.n249 VDD.n248 1.06836
R490 VDD.n219 VDD.n218 1.04079
R491 VDD.n164 VDD.n163 1.03836
R492 VDD.n100 VDD.n50 1.02405
R493 VDD.n372 VDD.n371 0.993021
R494 VDD.n231 VDD.n230 0.840632
R495 VDD.n143 VDD 0.533317
R496 VDD.n302 VDD 0.468962
R497 VDD.n238 VDD.n237 0.337997
R498 VDD.n237 VDD.n236 0.328132
R499 VDD VDD.n300 0.243482
R500 VDD.n272 VDD.n271 0.233919
R501 VDD.n269 VDD.n268 0.233919
R502 VDD.n149 VDD.n138 0.233919
R503 VDD.n155 VDD.n154 0.233919
R504 VDD.n213 VDD.n212 0.233919
R505 VDD.n210 VDD.n209 0.233919
R506 VDD.n78 VDD.n77 0.233919
R507 VDD.n75 VDD.n74 0.233919
R508 VDD.n45 VDD.n44 0.233919
R509 VDD.n42 VDD.n41 0.233919
R510 VDD.n243 VDD.n242 0.233919
R511 VDD.n240 VDD.n239 0.233919
R512 VDD.n357 VDD.n348 0.233919
R513 VDD.n363 VDD.n362 0.233919
R514 VDD.n220 VDD.n219 0.211434
R515 VDD.n295 VDD 0.185839
R516 VDD.n221 VDD 0.182611
R517 VDD VDD.n51 0.179233
R518 VDD.n301 VDD 0.17738
R519 VDD.n219 VDD.n189 0.158852
R520 VDD.n100 VDD.n99 0.152441
R521 VDD.n294 VDD 0.147753
R522 VDD.n275 VDD.n274 0.141016
R523 VDD.n282 VDD.n281 0.141016
R524 VDD.n283 VDD.n254 0.141016
R525 VDD.n158 VDD.n157 0.141016
R526 VDD.n216 VDD.n215 0.141016
R527 VDD.n81 VDD.n80 0.141016
R528 VDD.n88 VDD.n87 0.141016
R529 VDD.n89 VDD.n55 0.141016
R530 VDD.n48 VDD.n47 0.141016
R531 VDD.n102 VDD.n23 0.141016
R532 VDD.n108 VDD.n107 0.141016
R533 VDD.n246 VDD.n245 0.141016
R534 VDD.n366 VDD.n365 0.141016
R535 VDD.n101 VDD.n100 0.131304
R536 VDD VDD.n288 0.122435
R537 VDD VDD.n94 0.122435
R538 VDD.n109 VDD 0.122435
R539 VDD.n289 VDD 0.111984
R540 VDD.n95 VDD 0.111984
R541 VDD.n277 VDD.n276 0.107339
R542 VDD.n274 VDD.n273 0.107339
R543 VDD.n280 VDD.n278 0.107339
R544 VDD.n284 VDD.n282 0.107339
R545 VDD.n287 VDD.n254 0.107339
R546 VDD.n159 VDD.n158 0.107339
R547 VDD.n163 VDD.n162 0.107339
R548 VDD.n218 VDD.n217 0.107339
R549 VDD.n215 VDD.n214 0.107339
R550 VDD.n83 VDD.n82 0.107339
R551 VDD.n80 VDD.n79 0.107339
R552 VDD.n86 VDD.n84 0.107339
R553 VDD.n90 VDD.n88 0.107339
R554 VDD.n93 VDD.n55 0.107339
R555 VDD.n50 VDD.n49 0.107339
R556 VDD.n47 VDD.n46 0.107339
R557 VDD.n103 VDD.n101 0.107339
R558 VDD.n106 VDD.n23 0.107339
R559 VDD.n110 VDD.n108 0.107339
R560 VDD.n248 VDD.n247 0.107339
R561 VDD.n245 VDD.n244 0.107339
R562 VDD.n367 VDD.n366 0.107339
R563 VDD.n371 VDD.n370 0.107339
R564 VDD.n292 VDD.n291 0.10725
R565 VDD.n226 VDD 0.106795
R566 VDD VDD.n149 0.106758
R567 VDD.n154 VDD 0.106758
R568 VDD VDD.n357 0.106758
R569 VDD.n362 VDD 0.106758
R570 VDD.n271 VDD 0.106177
R571 VDD.n268 VDD 0.106177
R572 VDD.n212 VDD 0.106177
R573 VDD.n209 VDD 0.106177
R574 VDD.n77 VDD 0.106177
R575 VDD.n74 VDD 0.106177
R576 VDD VDD.n95 0.106177
R577 VDD.n44 VDD 0.106177
R578 VDD.n41 VDD 0.106177
R579 VDD.n223 VDD 0.106177
R580 VDD.n242 VDD 0.106177
R581 VDD.n239 VDD 0.106177
R582 VDD.n203 VDD 0.102091
R583 VDD.n299 VDD.n291 0.0854231
R584 VDD.n250 VDD.n249 0.0852977
R585 VDD.n224 VDD.n223 0.0846936
R586 VDD.n270 VDD.n269 0.080629
R587 VDD.n150 VDD.n146 0.080629
R588 VDD.n153 VDD.n138 0.080629
R589 VDD.n211 VDD.n210 0.080629
R590 VDD.n208 VDD.n207 0.080629
R591 VDD.n76 VDD.n75 0.080629
R592 VDD.n73 VDD.n72 0.080629
R593 VDD.n96 VDD.n51 0.080629
R594 VDD.n43 VDD.n42 0.080629
R595 VDD.n40 VDD.n39 0.080629
R596 VDD.n222 VDD.n221 0.080629
R597 VDD.n241 VDD.n240 0.080629
R598 VDD.n358 VDD.n354 0.080629
R599 VDD.n361 VDD.n348 0.080629
R600 VDD VDD.n275 0.0794677
R601 VDD VDD.n272 0.0794677
R602 VDD.n281 VDD 0.0794677
R603 VDD VDD.n283 0.0794677
R604 VDD.n288 VDD 0.0794677
R605 VDD VDD.n216 0.0794677
R606 VDD VDD.n213 0.0794677
R607 VDD VDD.n81 0.0794677
R608 VDD VDD.n78 0.0794677
R609 VDD.n87 VDD 0.0794677
R610 VDD VDD.n89 0.0794677
R611 VDD.n94 VDD 0.0794677
R612 VDD VDD.n48 0.0794677
R613 VDD VDD.n45 0.0794677
R614 VDD VDD.n102 0.0794677
R615 VDD.n107 VDD 0.0794677
R616 VDD VDD.n109 0.0794677
R617 VDD VDD.n246 0.0794677
R618 VDD VDD.n243 0.0794677
R619 VDD VDD.n155 0.0788871
R620 VDD.n157 VDD 0.0788871
R621 VDD VDD.n363 0.0788871
R622 VDD.n365 VDD 0.0788871
R623 VDD.n235 VDD 0.0733571
R624 VDD VDD.n294 0.0674231
R625 VDD.n300 VDD 0.0605
R626 VDD.n302 VDD.n301 0.0562419
R627 VDD.n308 VDD.n249 0.0557941
R628 VDD.n188 VDD.n187 0.0505302
R629 VDD.n166 VDD.n165 0.0505302
R630 VDD.n327 VDD.n326 0.0480988
R631 VDD.n177 VDD.n176 0.0478112
R632 VDD.n236 VDD.n235 0.0471071
R633 VDD.n322 VDD.n318 0.0470046
R634 VDD.n335 VDD.n334 0.0470046
R635 VDD.n308 VDD 0.046755
R636 VDD.n317 VDD 0.046731
R637 VDD.n182 VDD.n181 0.0467236
R638 VDD.n172 VDD.n171 0.0467236
R639 VDD VDD.n336 0.0464574
R640 VDD VDD.n183 0.0464517
R641 VDD.n170 VDD 0.0461798
R642 VDD VDD.n220 0.0457727
R643 VDD.n99 VDD 0.0444412
R644 VDD VDD.n250 0.0438334
R645 VDD.n302 VDD.n289 0.0411452
R646 VDD VDD.n330 0.0377036
R647 VDD VDD.n174 0.0374789
R648 VDD.n320 VDD 0.0374301
R649 VDD.n179 VDD 0.0372069
R650 VDD VDD.n292 0.036939
R651 VDD.n234 VDD.n233 0.0358571
R652 VDD.n236 VDD.n234 0.03425
R653 VDD VDD.n372 0.0327059
R654 VDD VDD.n321 0.0325061
R655 VDD VDD.n180 0.0323127
R656 VDD.n329 VDD 0.0322325
R657 VDD.n173 VDD 0.0320408
R658 VDD VDD.n373 0.0298382
R659 VDD.n224 VDD 0.0277903
R660 VDD.n321 VDD.n320 0.0262143
R661 VDD.n330 VDD.n329 0.0262143
R662 VDD.n180 VDD.n179 0.0260589
R663 VDD.n174 VDD.n173 0.0260589
R664 VDD VDD.n164 0.023068
R665 VDD.n189 VDD 0.0227961
R666 VDD.n316 VDD.n6 0.020196
R667 VDD.n340 VDD.n339 0.020196
R668 VDD.n303 VDD.n302 0.0201154
R669 VDD.n185 VDD.n184 0.020077
R670 VDD.n169 VDD.n168 0.020077
R671 VDD VDD.n188 0.0198051
R672 VDD VDD.n312 0.0196489
R673 VDD VDD.n186 0.0195332
R674 VDD.n165 VDD 0.0195332
R675 VDD.n338 VDD 0.0193754
R676 VDD.n167 VDD 0.0192613
R677 VDD.n312 VDD.n6 0.0185547
R678 VDD.n339 VDD.n338 0.0185547
R679 VDD.n186 VDD.n185 0.0184456
R680 VDD.n168 VDD.n167 0.0184456
R681 VDD.n313 VDD.n310 0.0144514
R682 VDD.n373 VDD.n343 0.0141778
R683 VDD.n205 VDD.n204 0.0141364
R684 VDD.n141 VDD 0.012875
R685 VDD.n144 VDD 0.00810563
R686 VDD.n204 VDD.n203 0.00725
R687 VDD.n351 VDD 0.00725
R688 VDD.n205 VDD 0.00595455
R689 VDD.n204 VDD 0.00595455
R690 VDD.n70 VDD 0.00543151
R691 VDD.n235 VDD 0.00478571
R692 VDD.n373 VDD 0.00469118
R693 VDD.n318 VDD.n317 0.00432979
R694 VDD.n336 VDD.n335 0.00432979
R695 VDD.n183 VDD.n182 0.00430665
R696 VDD.n171 VDD.n170 0.00430665
R697 VDD VDD.n299 0.00419231
R698 VDD.n295 VDD 0.00373077
R699 VDD.n233 VDD.n232 0.00371429
R700 VDD.n326 VDD.n325 0.00323556
R701 VDD.n331 VDD.n327 0.00323556
R702 VDD.n178 VDD.n177 0.00321903
R703 VDD.n176 VDD.n175 0.00321903
R704 VDD.n37 VDD 0.00256897
R705 VDD.n310 VDD.n308 0.00229283
R706 VDD.n159 VDD 0.00224194
R707 VDD.n162 VDD 0.00224194
R708 VDD.n367 VDD 0.00224194
R709 VDD.n370 VDD 0.00224194
R710 VDD.n232 VDD.n229 0.00210714
R711 VDD.n144 VDD.n143 0.00176761
R712 VDD.n276 VDD 0.00166129
R713 VDD.n273 VDD 0.00166129
R714 VDD VDD.n270 0.00166129
R715 VDD VDD.n267 0.00166129
R716 VDD VDD.n280 0.00166129
R717 VDD.n284 VDD 0.00166129
R718 VDD VDD.n287 0.00166129
R719 VDD.n217 VDD 0.00166129
R720 VDD.n214 VDD 0.00166129
R721 VDD VDD.n211 0.00166129
R722 VDD VDD.n208 0.00166129
R723 VDD.n82 VDD 0.00166129
R724 VDD.n79 VDD 0.00166129
R725 VDD VDD.n76 0.00166129
R726 VDD VDD.n73 0.00166129
R727 VDD VDD.n86 0.00166129
R728 VDD.n90 VDD 0.00166129
R729 VDD VDD.n93 0.00166129
R730 VDD.n96 VDD 0.00166129
R731 VDD.n49 VDD 0.00166129
R732 VDD.n46 VDD 0.00166129
R733 VDD VDD.n43 0.00166129
R734 VDD VDD.n40 0.00166129
R735 VDD.n103 VDD 0.00166129
R736 VDD VDD.n106 0.00166129
R737 VDD.n110 VDD 0.00166129
R738 VDD VDD.n222 0.00166129
R739 VDD.n247 VDD 0.00166129
R740 VDD.n244 VDD 0.00166129
R741 VDD VDD.n241 0.00166129
R742 VDD VDD.n238 0.00166129
R743 VDD.n201 VDD 0.00152273
R744 VDD.n325 VDD 0.00132067
R745 VDD.n334 VDD 0.00132067
R746 VDD.n343 VDD 0.00132067
R747 VDD VDD.n178 0.00131571
R748 VDD VDD.n172 0.00131571
R749 VDD VDD.n166 0.00131571
R750 VDD.n150 VDD 0.00108064
R751 VDD VDD.n153 0.00108064
R752 VDD.n358 VDD 0.00108064
R753 VDD VDD.n361 0.00108064
R754 VDD.n303 VDD 0.00107692
R755 VDD.n313 VDD 0.00104711
R756 VDD.n322 VDD 0.00104711
R757 VDD.n331 VDD 0.00104711
R758 VDD.n340 VDD 0.00104711
R759 VDD.n187 VDD 0.00104381
R760 VDD.n181 VDD 0.00104381
R761 VDD.n175 VDD 0.00104381
R762 VDD VDD.n169 0.00104381
R763 VDD VDD.n316 0.000773556
R764 VDD.n184 VDD 0.000771903
R765 CLK.n1 CLK.t1 36.935
R766 CLK.n5 CLK.t4 36.935
R767 CLK.n14 CLK.t5 25.4742
R768 CLK.n1 CLK.t0 18.1962
R769 CLK.n5 CLK.t2 18.1962
R770 CLK.n14 CLK.t3 14.142
R771 CLK.n12 CLK.n4 2.25107
R772 CLK.n16 CLK.n13 2.24196
R773 CLK.n8 CLK.n5 2.12464
R774 CLK.n2 CLK.n1 2.12188
R775 CLK.n11 CLK.n10 1.71671
R776 CLK.n9 CLK.n8 1.50503
R777 CLK.n15 CLK.n14 1.42126
R778 CLK.n13 CLK.n12 0.969075
R779 CLK CLK.n17 0.1605
R780 CLK.n3 CLK 0.0457995
R781 CLK.n6 CLK 0.0457995
R782 CLK.n10 CLK.n9 0.0386356
R783 CLK.n4 CLK.n3 0.0377414
R784 CLK.n7 CLK.n6 0.0377414
R785 CLK.n17 CLK.n16 0.03175
R786 CLK.n13 CLK.n0 0.0238218
R787 CLK.n12 CLK.n11 0.0122182
R788 CLK.n4 CLK.n2 0.00360345
R789 CLK.n8 CLK.n7 0.00203726
R790 CLK.n16 CLK.n15 0.00175
R791 VSS.n168 VSS.n167 3.48725e+06
R792 VSS.t106 VSS.n71 1.74697e+06
R793 VSS.n22 VSS.n21 1.11109e+06
R794 VSS.n77 VSS.t58 285299
R795 VSS.n21 VSS.t75 284437
R796 VSS.n222 VSS.n221 110325
R797 VSS.n221 VSS.t134 89236.1
R798 VSS.n71 VSS.n22 22695.3
R799 VSS.n167 VSS.n22 15212.9
R800 VSS.n78 VSS.n77 13762.5
R801 VSS.n38 VSS.n37 8589.75
R802 VSS.n179 VSS.n169 8129.71
R803 VSS.n134 VSS.n133 7369.71
R804 VSS.n151 VSS.t80 5069.75
R805 VSS.n167 VSS.t47 4991.36
R806 VSS.n77 VSS.n76 4628.79
R807 VSS.n181 VSS.n180 4482.15
R808 VSS.n120 VSS.n104 3320.93
R809 VSS.t6 VSS.n151 3278.56
R810 VSS.t56 VSS.n78 3194.51
R811 VSS.n180 VSS.t183 2872.22
R812 VSS.t143 VSS.t154 2781.65
R813 VSS.n104 VSS.t82 2689.86
R814 VSS.n104 VSS.t129 2684.02
R815 VSS.n180 VSS.t71 2599.49
R816 VSS.t125 VSS.t176 2357.27
R817 VSS.t49 VSS.t173 2357.27
R818 VSS.t224 VSS.t112 2357.27
R819 VSS.t127 VSS.t141 2357.27
R820 VSS.t150 VSS.t207 2307.56
R821 VSS.t214 VSS.t92 2307.56
R822 VSS.t223 VSS.t89 2307.56
R823 VSS.t34 VSS.t50 2307.56
R824 VSS.t167 VSS.t87 2307.56
R825 VSS.t180 VSS.t226 2307.56
R826 VSS.t107 VSS.t27 2307.56
R827 VSS.t229 VSS.t169 2307.56
R828 VSS.t140 VSS.t0 2307.56
R829 VSS.t205 VSS.t156 2307.56
R830 VSS.t102 VSS.t201 2307.56
R831 VSS.t40 VSS.t24 2307.56
R832 VSS.t31 VSS.t5 2307.56
R833 VSS.t66 VSS.t15 2307.56
R834 VSS.t95 VSS.t124 2307.56
R835 VSS.t17 VSS.t103 2307.56
R836 VSS.t137 VSS.t179 2307.56
R837 VSS.t131 VSS.t78 2307.56
R838 VSS.t189 VSS.t225 2307.56
R839 VSS.t20 VSS.t219 2307.56
R840 VSS.t121 VSS.t213 2307.56
R841 VSS.n169 VSS.n168 2273.68
R842 VSS.t108 VSS.t192 2191.99
R843 VSS.t196 VSS.t139 2191.99
R844 VSS.t23 VSS.t148 2107.54
R845 VSS.t185 VSS.t38 2107.54
R846 VSS.t88 VSS.t152 2090.76
R847 VSS.t36 VSS.t209 2090.76
R848 VSS.t151 VSS.t162 2090.76
R849 VSS.t119 VSS.t42 2090.76
R850 VSS.n133 VSS.t212 1930.58
R851 VSS.n179 VSS.t114 1751.51
R852 VSS.n221 VSS.t204 1650.7
R853 VSS.t178 VSS.n105 1644.99
R854 VSS.t120 VSS.n38 1588.77
R855 VSS.n133 VSS.n120 1565.03
R856 VSS.n181 VSS.n179 1365.3
R857 VSS.n39 VSS.t10 1272.1
R858 VSS.n204 VSS.t193 1272.1
R859 VSS.n183 VSS.t186 1272.1
R860 VSS.n165 VSS.t135 1199.47
R861 VSS.n76 VSS.t63 1199.47
R862 VSS.n203 VSS.t68 1199.47
R863 VSS.t47 VSS.n166 941.59
R864 VSS.t133 VSS.t105 933.573
R865 VSS.t128 VSS.t49 933.573
R866 VSS.t123 VSS.t22 933.573
R867 VSS.t184 VSS.t127 933.573
R868 VSS.t53 VSS.t223 913.885
R869 VSS.t52 VSS.t7 913.885
R870 VSS.t13 VSS.t107 913.885
R871 VSS.t211 VSS.t205 913.885
R872 VSS.t206 VSS.t115 913.885
R873 VSS.t179 VSS.t130 913.885
R874 VSS.t213 VSS.t188 913.885
R875 VSS.t192 VSS.t9 868.115
R876 VSS.t111 VSS.t172 868.115
R877 VSS.t86 VSS.t30 834.672
R878 VSS.t14 VSS.t185 834.672
R879 VSS.t37 VSS.n134 833.202
R880 VSS.t222 VSS.t228 828.027
R881 VSS.t55 VSS.t36 828.027
R882 VSS.t199 VSS.t216 828.027
R883 VSS.t44 VSS.t119 828.027
R884 VSS.n81 VSS.t116 776.83
R885 VSS.n0 VSS.t54 560.144
R886 VSS.n1 VSS.t125 560.144
R887 VSS.n2 VSS.t133 560.144
R888 VSS.n3 VSS.t128 560.144
R889 VSS.t129 VSS.n5 560.144
R890 VSS.n6 VSS.t224 560.144
R891 VSS.n7 VSS.t123 560.144
R892 VSS.n8 VSS.t184 560.144
R893 VSS.t154 VSS.n81 554.879
R894 VSS.n26 VSS.t91 548.331
R895 VSS.n27 VSS.t150 548.331
R896 VSS.n32 VSS.t92 548.331
R897 VSS.n33 VSS.t53 548.331
R898 VSS.n152 VSS.t6 548.331
R899 VSS.n157 VSS.t87 548.331
R900 VSS.n158 VSS.t180 548.331
R901 VSS.n164 VSS.t52 548.331
R902 VSS.n75 VSS.t13 548.331
R903 VSS.n74 VSS.t229 548.331
R904 VSS.n73 VSS.t140 548.331
R905 VSS.n72 VSS.t106 548.331
R906 VSS.n202 VSS.t211 548.331
R907 VSS.n201 VSS.t102 548.331
R908 VSS.n200 VSS.t220 548.331
R909 VSS.n196 VSS.t204 548.331
R910 VSS.t114 VSS.n178 548.331
R911 VSS.t24 VSS.n177 548.331
R912 VSS.t5 VSS.n176 548.331
R913 VSS.n224 VSS.t206 548.331
R914 VSS.n106 VSS.t178 548.331
R915 VSS.n111 VSS.t124 548.331
R916 VSS.n112 VSS.t17 548.331
R917 VSS.n117 VSS.t130 548.331
R918 VSS.t212 VSS.n132 548.331
R919 VSS.t225 VSS.n131 548.331
R920 VSS.t219 VSS.n130 548.331
R921 VSS.t188 VSS.n129 548.331
R922 VSS.n85 VSS.t33 546.41
R923 VSS.t9 VSS.n42 520.869
R924 VSS.n44 VSS.t111 520.869
R925 VSS.t139 VSS.n46 520.869
R926 VSS.n48 VSS.t191 520.869
R927 VSS.t183 VSS.n10 500.803
R928 VSS.n11 VSS.t23 500.803
R929 VSS.n12 VSS.t86 500.803
R930 VSS.n13 VSS.t14 500.803
R931 VSS.n135 VSS.t37 496.815
R932 VSS.n136 VSS.t88 496.815
R933 VSS.n137 VSS.t222 496.815
R934 VSS.n139 VSS.t55 496.815
R935 VSS.n95 VSS.t120 496.815
R936 VSS.n96 VSS.t151 496.815
R937 VSS.n100 VSS.t199 496.815
R938 VSS.n101 VSS.t44 496.815
R939 VSS.t159 VSS.t126 468.094
R940 VSS.t221 VSS.t164 468.094
R941 VSS.t176 VSS.n0 373.43
R942 VSS.n1 VSS.t18 373.43
R943 VSS.t173 VSS.n2 373.43
R944 VSS.t82 VSS.n3 373.43
R945 VSS.t112 VSS.n5 373.43
R946 VSS.n6 VSS.t217 373.43
R947 VSS.t141 VSS.n7 373.43
R948 VSS.t71 VSS.n8 373.43
R949 VSS.t207 VSS.n26 365.555
R950 VSS.n27 VSS.t214 365.555
R951 VSS.t89 VSS.n32 365.555
R952 VSS.n33 VSS.t34 365.555
R953 VSS.n152 VSS.t167 365.555
R954 VSS.t226 VSS.n157 365.555
R955 VSS.n158 VSS.t97 365.555
R956 VSS.t135 VSS.n164 365.555
R957 VSS.t63 VSS.n75 365.555
R958 VSS.t27 VSS.n74 365.555
R959 VSS.t169 VSS.n73 365.555
R960 VSS.t0 VSS.n72 365.555
R961 VSS.t68 VSS.n202 365.555
R962 VSS.t156 VSS.n201 365.555
R963 VSS.t201 VSS.n200 365.555
R964 VSS.n196 VSS.t145 365.555
R965 VSS.n178 VSS.t40 365.555
R966 VSS.n177 VSS.t31 365.555
R967 VSS.n176 VSS.t25 365.555
R968 VSS.n224 VSS.t66 365.555
R969 VSS.n106 VSS.t95 365.555
R970 VSS.t103 VSS.n111 365.555
R971 VSS.n112 VSS.t137 365.555
R972 VSS.t78 VSS.n117 365.555
R973 VSS.n132 VSS.t189 365.555
R974 VSS.n131 VSS.t20 365.555
R975 VSS.n130 VSS.t121 365.555
R976 VSS.n129 VSS.t84 365.555
R977 VSS.n85 VSS.t45 364.274
R978 VSS.n42 VSS.t58 347.245
R979 VSS.n44 VSS.t108 347.245
R980 VSS.n46 VSS.t230 347.245
R981 VSS.n48 VSS.t196 347.245
R982 VSS.n120 VSS.n119 336.995
R983 VSS.t148 VSS.n10 333.868
R984 VSS.n11 VSS.t3 333.868
R985 VSS.t38 VSS.n12 333.868
R986 VSS.n13 VSS.t60 333.868
R987 VSS.t152 VSS.n135 331.211
R988 VSS.n136 VSS.t181 331.211
R989 VSS.t209 VSS.n137 331.211
R990 VSS.n139 VSS.t73 331.211
R991 VSS.t162 VSS.n95 331.211
R992 VSS.n96 VSS.t93 331.211
R993 VSS.t42 VSS.n100 331.211
R994 VSS.n101 VSS.t80 331.211
R995 VSS.t126 VSS.t175 185.383
R996 VSS.t8 VSS.t200 185.383
R997 VSS.n182 VSS.n181 172.349
R998 VSS.n151 VSS.n150 119.948
R999 VSS.t175 VSS.n212 111.231
R1000 VSS.n213 VSS.t8 111.231
R1001 VSS.n216 VSS.t221 111.231
R1002 VSS.t134 VSS.n220 111.231
R1003 VSS.n212 VSS.t75 74.1538
R1004 VSS.n213 VSS.t159 74.1538
R1005 VSS.n216 VSS.t99 74.1538
R1006 VSS.n220 VSS.t164 74.1538
R1007 VSS.n223 VSS.n222 51.4065
R1008 VSS.n79 VSS.t56 47.5615
R1009 VSS.n183 VSS.n182 41.0359
R1010 VSS.n150 VSS.t50 34.2711
R1011 VSS.t15 VSS.n223 34.2711
R1012 VSS.n119 VSS.t131 34.2711
R1013 VSS.n82 VSS.t143 34.1511
R1014 VSS.n76 VSS.n39 32.8288
R1015 VSS.n204 VSS.n203 32.8288
R1016 VSS.n134 VSS.t80 32.6553
R1017 VSS.n166 VSS.n165 30.3743
R1018 VSS.n118 VSS.t132 9.3736
R1019 VSS.n14 VSS.t16 9.3736
R1020 VSS.n149 VSS.t51 9.3736
R1021 VSS.n23 VSS.t48 9.3736
R1022 VSS.n58 VSS.n57 9.37275
R1023 VSS.n84 VSS.t144 9.36521
R1024 VSS.n188 VSS.n187 9.3508
R1025 VSS.n90 VSS.n80 9.3221
R1026 VSS.n88 VSS.t155 9.3221
R1027 VSS.n91 VSS.t57 9.30652
R1028 VSS.n185 VSS.t187 9.30652
R1029 VSS.n186 VSS.n185 9.19275
R1030 VSS VSS.t46 7.30633
R1031 VSS.n108 VSS.t96 7.19156
R1032 VSS.n109 VSS.t104 7.19156
R1033 VSS.n114 VSS.t138 7.19156
R1034 VSS.n234 VSS.t149 7.19156
R1035 VSS.n232 VSS.t4 7.19156
R1036 VSS.n171 VSS.t41 7.19156
R1037 VSS.n173 VSS.t32 7.19156
R1038 VSS.n174 VSS.t26 7.19156
R1039 VSS.n93 VSS.t163 7.19156
R1040 VSS.n98 VSS.t94 7.19156
R1041 VSS.n24 VSS.t208 7.19156
R1042 VSS.n29 VSS.t215 7.19156
R1043 VSS.n30 VSS.t90 7.19156
R1044 VSS.n145 VSS.t153 7.19156
R1045 VSS.n143 VSS.t182 7.19156
R1046 VSS.n154 VSS.t168 7.19156
R1047 VSS.n155 VSS.t227 7.19156
R1048 VSS.n160 VSS.t98 7.19156
R1049 VSS.n198 VSS.n195 7.19156
R1050 VSS.n194 VSS.n193 7.19156
R1051 VSS.n191 VSS.n190 7.19156
R1052 VSS.n69 VSS.n68 7.19156
R1053 VSS.n66 VSS.n65 7.19156
R1054 VSS.n63 VSS.n62 7.19156
R1055 VSS.n122 VSS.t190 7.19156
R1056 VSS.n124 VSS.t21 7.19156
R1057 VSS.n126 VSS.t122 7.19156
R1058 VSS.n218 VSS.n15 7.14989
R1059 VSS.n215 VSS.n16 7.14989
R1060 VSS.n50 VSS.n47 7.14489
R1061 VSS.n52 VSS.n45 7.14489
R1062 VSS.n252 VSS.t177 7.11489
R1063 VSS.n250 VSS.t19 7.11489
R1064 VSS.n243 VSS.t113 7.11489
R1065 VSS.n241 VSS.t218 7.11489
R1066 VSS.n115 VSS.t79 5.91399
R1067 VSS.n230 VSS.t39 5.91399
R1068 VSS.n228 VSS.t61 5.91399
R1069 VSS.n226 VSS.t67 5.91399
R1070 VSS.n36 VSS.t43 5.91399
R1071 VSS.n103 VSS.t81 5.91399
R1072 VSS.n35 VSS.t35 5.91399
R1073 VSS.n141 VSS.t210 5.91399
R1074 VSS.n138 VSS.t74 5.91399
R1075 VSS.n162 VSS.t136 5.91399
R1076 VSS.n19 VSS.n18 5.91399
R1077 VSS.n60 VSS.n40 5.91399
R1078 VSS.n127 VSS.t85 5.91399
R1079 VSS.n210 VSS.n209 5.87232
R1080 VSS.n208 VSS.n17 5.87232
R1081 VSS.n54 VSS.n43 5.86732
R1082 VSS.n56 VSS.n41 5.86732
R1083 VSS.n248 VSS.t174 5.83732
R1084 VSS.n246 VSS.t83 5.83732
R1085 VSS.n239 VSS.t142 5.83732
R1086 VSS.n237 VSS.t72 5.83732
R1087 VSS.n55 VSS.n42 5.2005
R1088 VSS.n53 VSS.n44 5.2005
R1089 VSS.n51 VSS.n46 5.2005
R1090 VSS.n49 VSS.n48 5.2005
R1091 VSS.n140 VSS.n139 5.2005
R1092 VSS.n142 VSS.n137 5.2005
R1093 VSS.n144 VSS.n136 5.2005
R1094 VSS.n146 VSS.n135 5.2005
R1095 VSS.n102 VSS.n101 5.2005
R1096 VSS.n100 VSS.n99 5.2005
R1097 VSS.n97 VSS.n96 5.2005
R1098 VSS.n95 VSS.n94 5.2005
R1099 VSS.n153 VSS.n152 5.2005
R1100 VSS.n157 VSS.n156 5.2005
R1101 VSS.n159 VSS.n158 5.2005
R1102 VSS.n164 VSS.n163 5.2005
R1103 VSS.n26 VSS.n25 5.2005
R1104 VSS.n28 VSS.n27 5.2005
R1105 VSS.n32 VSS.n31 5.2005
R1106 VSS.n34 VSS.n33 5.2005
R1107 VSS.n150 VSS.n149 5.2005
R1108 VSS.n89 VSS.n81 5.2005
R1109 VSS.n92 VSS.n79 5.2005
R1110 VSS.n86 VSS.n85 5.2005
R1111 VSS.n83 VSS.n82 5.2005
R1112 VSS.n58 VSS.n39 5.2005
R1113 VSS.n72 VSS.n70 5.2005
R1114 VSS.n73 VSS.n67 5.2005
R1115 VSS.n74 VSS.n64 5.2005
R1116 VSS.n75 VSS.n61 5.2005
R1117 VSS.n166 VSS.n23 5.2005
R1118 VSS.n205 VSS.n204 5.2005
R1119 VSS.n220 VSS.n219 5.2005
R1120 VSS.n217 VSS.n216 5.2005
R1121 VSS.n214 VSS.n213 5.2005
R1122 VSS.n212 VSS.n211 5.2005
R1123 VSS.n197 VSS.n196 5.2005
R1124 VSS.n200 VSS.n199 5.2005
R1125 VSS.n201 VSS.n192 5.2005
R1126 VSS.n202 VSS.n189 5.2005
R1127 VSS.n178 VSS.n170 5.2005
R1128 VSS.n177 VSS.n172 5.2005
R1129 VSS.n176 VSS.n175 5.2005
R1130 VSS.n225 VSS.n224 5.2005
R1131 VSS.n223 VSS.n14 5.2005
R1132 VSS.n229 VSS.n13 5.2005
R1133 VSS.n231 VSS.n12 5.2005
R1134 VSS.n233 VSS.n11 5.2005
R1135 VSS.n235 VSS.n10 5.2005
R1136 VSS.n184 VSS.n183 5.2005
R1137 VSS.n107 VSS.n106 5.2005
R1138 VSS.n111 VSS.n110 5.2005
R1139 VSS.n113 VSS.n112 5.2005
R1140 VSS.n117 VSS.n116 5.2005
R1141 VSS.n119 VSS.n118 5.2005
R1142 VSS.n129 VSS.n128 5.2005
R1143 VSS.n130 VSS.n125 5.2005
R1144 VSS.n131 VSS.n123 5.2005
R1145 VSS.n132 VSS.n121 5.2005
R1146 VSS.n238 VSS.n8 5.2005
R1147 VSS.n240 VSS.n7 5.2005
R1148 VSS.n242 VSS.n6 5.2005
R1149 VSS.n244 VSS.n5 5.2005
R1150 VSS.n247 VSS.n3 5.2005
R1151 VSS.n249 VSS.n2 5.2005
R1152 VSS.n251 VSS.n1 5.2005
R1153 VSS.n253 VSS.n0 5.2005
R1154 VSS.n207 VSS 1.98504
R1155 VSS.n228 VSS.n227 0.943665
R1156 VSS.n59 VSS.n56 0.918836
R1157 VSS.n148 VSS.n147 0.845914
R1158 VSS.n207 VSS.n206 0.825821
R1159 VSS.n245 VSS.n4 0.807932
R1160 VSS.n236 VSS.n9 0.807932
R1161 VSS.n138 VSS.n20 0.692427
R1162 VSS.n99 VSS.n98 0.480225
R1163 VSS.n102 VSS.n36 0.480225
R1164 VSS.n143 VSS.n142 0.480225
R1165 VSS.n141 VSS.n140 0.480225
R1166 VSS VSS.n108 0.343161
R1167 VSS.n109 VSS 0.343161
R1168 VSS VSS.n171 0.343161
R1169 VSS VSS.n173 0.343161
R1170 VSS.n24 VSS 0.343161
R1171 VSS VSS.n29 0.343161
R1172 VSS VSS.n154 0.343161
R1173 VSS.n155 VSS 0.343161
R1174 VSS.n194 VSS 0.343161
R1175 VSS VSS.n198 0.343161
R1176 VSS.n66 VSS 0.343161
R1177 VSS.n69 VSS 0.343161
R1178 VSS.n93 VSS 0.343161
R1179 VSS.n145 VSS 0.343161
R1180 VSS VSS.n122 0.343161
R1181 VSS VSS.n124 0.343161
R1182 VSS.n245 VSS 0.336214
R1183 VSS.n88 VSS.n87 0.309418
R1184 VSS.n211 VSS.n210 0.308088
R1185 VSS.n215 VSS.n214 0.308088
R1186 VSS.n116 VSS 0.289491
R1187 VSS.n225 VSS 0.289491
R1188 VSS.n34 VSS 0.289491
R1189 VSS.n163 VSS 0.289491
R1190 VSS VSS.n189 0.289491
R1191 VSS VSS.n61 0.289491
R1192 VSS.n128 VSS 0.289491
R1193 VSS.n250 VSS.n249 0.277167
R1194 VSS.n248 VSS.n247 0.277167
R1195 VSS.n241 VSS.n240 0.277167
R1196 VSS.n239 VSS.n238 0.277167
R1197 VSS.n87 VSS.n86 0.255008
R1198 VSS.n161 VSS.n20 0.251419
R1199 VSS.n232 VSS.n231 0.250691
R1200 VSS.n230 VSS.n229 0.250691
R1201 VSS.n188 VSS.n186 0.246335
R1202 VSS.n55 VSS.n54 0.245993
R1203 VSS.n53 VSS.n52 0.245993
R1204 VSS.n218 VSS 0.220206
R1205 VSS.n252 VSS 0.198119
R1206 VSS.n243 VSS 0.198119
R1207 VSS.n186 VSS.n20 0.194066
R1208 VSS VSS.n114 0.191234
R1209 VSS.n174 VSS 0.191234
R1210 VSS.n30 VSS 0.191234
R1211 VSS VSS.n160 0.191234
R1212 VSS.n191 VSS 0.191234
R1213 VSS.n63 VSS 0.191234
R1214 VSS VSS.n126 0.191234
R1215 VSS.n147 VSS.n103 0.187931
R1216 VSS.n147 VSS 0.183803
R1217 VSS.n234 VSS 0.179208
R1218 VSS VSS.n50 0.175852
R1219 VSS.n91 VSS.n90 0.168119
R1220 VSS.n87 VSS.n84 0.141461
R1221 VSS VSS.n4 0.137685
R1222 VSS.n227 VSS 0.137685
R1223 VSS VSS.n148 0.137685
R1224 VSS.n161 VSS 0.137685
R1225 VSS VSS.n9 0.137685
R1226 VSS.n59 VSS 0.137136
R1227 VSS.n206 VSS 0.137136
R1228 VSS.n90 VSS.n89 0.136634
R1229 VSS.n236 VSS 0.123833
R1230 VSS.n208 VSS.n207 0.120147
R1231 VSS.n108 VSS.n107 0.118573
R1232 VSS.n110 VSS.n109 0.118573
R1233 VSS.n114 VSS.n113 0.118573
R1234 VSS.n171 VSS.n170 0.118573
R1235 VSS.n173 VSS.n172 0.118573
R1236 VSS.n175 VSS.n174 0.118573
R1237 VSS.n25 VSS.n24 0.118573
R1238 VSS.n29 VSS.n28 0.118573
R1239 VSS.n31 VSS.n30 0.118573
R1240 VSS.n154 VSS.n153 0.118573
R1241 VSS.n156 VSS.n155 0.118573
R1242 VSS.n160 VSS.n159 0.118573
R1243 VSS.n192 VSS.n191 0.118573
R1244 VSS.n199 VSS.n194 0.118573
R1245 VSS.n198 VSS.n197 0.118573
R1246 VSS.n64 VSS.n63 0.118573
R1247 VSS.n67 VSS.n66 0.118573
R1248 VSS.n70 VSS.n69 0.118573
R1249 VSS.n94 VSS.n93 0.118573
R1250 VSS.n98 VSS.n97 0.118573
R1251 VSS.n146 VSS.n145 0.118573
R1252 VSS.n144 VSS.n143 0.118573
R1253 VSS.n122 VSS.n121 0.118573
R1254 VSS.n124 VSS.n123 0.118573
R1255 VSS.n126 VSS.n125 0.118573
R1256 VSS VSS.n88 0.115458
R1257 VSS VSS.n115 0.115271
R1258 VSS.n226 VSS 0.115271
R1259 VSS.n35 VSS 0.115271
R1260 VSS VSS.n162 0.115271
R1261 VSS VSS.n19 0.115271
R1262 VSS VSS.n60 0.115271
R1263 VSS VSS.n36 0.115271
R1264 VSS.n103 VSS 0.115271
R1265 VSS VSS.n141 0.115271
R1266 VSS VSS.n138 0.115271
R1267 VSS VSS.n127 0.115271
R1268 VSS.n246 VSS.n245 0.108595
R1269 VSS.n237 VSS.n236 0.108595
R1270 VSS.n115 VSS.n4 0.10206
R1271 VSS.n227 VSS.n226 0.10206
R1272 VSS.n148 VSS.n35 0.10206
R1273 VSS.n162 VSS.n161 0.10206
R1274 VSS.n206 VSS.n19 0.10206
R1275 VSS.n60 VSS.n59 0.10206
R1276 VSS.n127 VSS.n9 0.10206
R1277 VSS.n217 VSS.n215 0.0762059
R1278 VSS.n219 VSS.n218 0.0762059
R1279 VSS VSS.n208 0.0740882
R1280 VSS.n210 VSS 0.0740882
R1281 VSS.n253 VSS.n252 0.0685952
R1282 VSS.n251 VSS.n250 0.0685952
R1283 VSS.n244 VSS.n243 0.0685952
R1284 VSS.n242 VSS.n241 0.0685952
R1285 VSS.n185 VSS.n184 0.0675755
R1286 VSS VSS.n248 0.0666905
R1287 VSS VSS.n246 0.0666905
R1288 VSS VSS.n239 0.0666905
R1289 VSS VSS.n237 0.0666905
R1290 VSS.n205 VSS.n188 0.066226
R1291 VSS.n235 VSS.n234 0.0620789
R1292 VSS.n233 VSS.n232 0.0620789
R1293 VSS.n52 VSS.n51 0.0609225
R1294 VSS.n50 VSS.n49 0.0609225
R1295 VSS VSS.n230 0.0603565
R1296 VSS VSS.n228 0.0603565
R1297 VSS.n56 VSS 0.0592324
R1298 VSS.n54 VSS 0.0592324
R1299 VSS.n84 VSS.n83 0.0589274
R1300 VSS.n92 VSS.n91 0.0564843
R1301 VSS.n107 VSS 0.00545413
R1302 VSS.n110 VSS 0.00545413
R1303 VSS.n113 VSS 0.00545413
R1304 VSS.n170 VSS 0.00545413
R1305 VSS.n172 VSS 0.00545413
R1306 VSS.n175 VSS 0.00545413
R1307 VSS.n25 VSS 0.00545413
R1308 VSS.n28 VSS 0.00545413
R1309 VSS.n31 VSS 0.00545413
R1310 VSS.n153 VSS 0.00545413
R1311 VSS.n156 VSS 0.00545413
R1312 VSS.n159 VSS 0.00545413
R1313 VSS VSS.n192 0.00545413
R1314 VSS.n199 VSS 0.00545413
R1315 VSS.n197 VSS 0.00545413
R1316 VSS VSS.n64 0.00545413
R1317 VSS VSS.n67 0.00545413
R1318 VSS.n70 VSS 0.00545413
R1319 VSS.n94 VSS 0.00545413
R1320 VSS.n97 VSS 0.00545413
R1321 VSS VSS.n146 0.00545413
R1322 VSS VSS.n144 0.00545413
R1323 VSS.n121 VSS 0.00545413
R1324 VSS.n123 VSS 0.00545413
R1325 VSS.n125 VSS 0.00545413
R1326 VSS.n116 VSS 0.00380275
R1327 VSS VSS.n225 0.00380275
R1328 VSS.n86 VSS 0.00380275
R1329 VSS VSS.n34 0.00380275
R1330 VSS.n163 VSS 0.00380275
R1331 VSS.n189 VSS 0.00380275
R1332 VSS.n61 VSS 0.00380275
R1333 VSS.n99 VSS 0.00380275
R1334 VSS VSS.n102 0.00380275
R1335 VSS.n142 VSS 0.00380275
R1336 VSS.n140 VSS 0.00380275
R1337 VSS.n128 VSS 0.00380275
R1338 VSS VSS.n217 0.00367647
R1339 VSS.n219 VSS 0.00367647
R1340 VSS.n89 VSS 0.00352521
R1341 VSS VSS.n253 0.00335714
R1342 VSS VSS.n251 0.00335714
R1343 VSS VSS.n244 0.00335714
R1344 VSS VSS.n242 0.00335714
R1345 VSS VSS.n235 0.00308373
R1346 VSS VSS.n233 0.00308373
R1347 VSS.n51 VSS 0.00303521
R1348 VSS.n49 VSS 0.00303521
R1349 VSS.n211 VSS 0.00261765
R1350 VSS.n214 VSS 0.00261765
R1351 VSS.n249 VSS 0.00240476
R1352 VSS.n247 VSS 0.00240476
R1353 VSS.n240 VSS 0.00240476
R1354 VSS.n238 VSS 0.00240476
R1355 VSS.n231 VSS 0.00222249
R1356 VSS.n229 VSS 0.00222249
R1357 VSS.n118 VSS 0.00219811
R1358 VSS.n14 VSS 0.00219811
R1359 VSS.n83 VSS 0.00219811
R1360 VSS.n149 VSS 0.00219811
R1361 VSS VSS.n23 0.00219811
R1362 VSS.n184 VSS 0.00219811
R1363 VSS VSS.n58 0.00219811
R1364 VSS VSS.n205 0.00219811
R1365 VSS VSS.n55 0.00219014
R1366 VSS VSS.n53 0.00219014
R1367 VSS VSS.n92 0.00191732
R1368 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 37.1986
R1369 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 31.528
R1370 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 30.5184
R1371 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 24.7029
R1372 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 17.6614
R1373 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 15.3826
R1374 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 12.0843
R1375 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 9.86691
R1376 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R1377 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 2.99416
R1378 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 2.2755
R1379 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2755
R1380 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 2.2505
R1381 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.24173
R1382 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.93723
R1383 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n2 1.81225
R1384 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.43709
R1385 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n1 0.281955
R1386 RST.n8 RST.t13 37.1991
R1387 RST.n47 RST.t1 36.935
R1388 RST.n0 RST.t3 36.935
R1389 RST.n14 RST.t7 36.935
R1390 RST.n35 RST.t11 36.935
R1391 RST.n24 RST.t6 36.935
R1392 RST.n20 RST.t9 36.935
R1393 RST.n47 RST.t0 18.1962
R1394 RST.n0 RST.t2 18.1962
R1395 RST.n14 RST.t5 18.1962
R1396 RST.n35 RST.t10 18.1962
R1397 RST.n24 RST.t4 18.1962
R1398 RST.n20 RST.t8 18.1962
R1399 RST.n8 RST.t12 17.66
R1400 RST.n22 RST.n21 5.63344
R1401 RST.n45 RST.n5 4.84685
R1402 RST.n53 RST.n45 4.63847
R1403 RST.n5 RST.n4 4.5005
R1404 RST.n45 RST.n11 4.41239
R1405 RST.n32 RST.n31 2.96983
R1406 RST RST.n57 2.26757
R1407 RST.n2 RST.n1 2.25731
R1408 RST.n27 RST.n26 2.24515
R1409 RST.n11 RST.n10 2.24157
R1410 RST.n21 RST.n20 2.1497
R1411 RST.n2 RST.n0 2.12457
R1412 RST.n25 RST.n24 2.12403
R1413 RST.n48 RST.n47 2.12207
R1414 RST.n15 RST.n14 2.12188
R1415 RST.n36 RST.n35 2.12175
R1416 RST.n56 RST.n55 2.06978
R1417 RST.n45 RST.n44 1.97488
R1418 RST.n51 RST.n50 1.5005
R1419 RST.n30 RST.n29 1.5005
R1420 RST.n38 RST.n37 1.5005
R1421 RST.n41 RST.n40 1.5005
R1422 RST.n17 RST.n16 1.5005
R1423 RST.n53 RST.n52 1.49882
R1424 RST.n44 RST.n19 1.4372
R1425 RST.n44 RST.n43 1.42363
R1426 RST.n9 RST.n8 1.41552
R1427 RST.n57 RST.n56 1.12776
R1428 RST.n19 RST.n18 1.12389
R1429 RST.n3 RST 0.0593097
R1430 RST.n21 RST 0.0445432
R1431 RST.n7 RST 0.0410354
R1432 RST.n49 RST 0.0394837
R1433 RST.n13 RST 0.0394837
R1434 RST.n34 RST 0.0379319
R1435 RST.n50 RST.n49 0.0377414
R1436 RST.n10 RST.n7 0.0361897
R1437 RST.n16 RST.n13 0.0361897
R1438 RST.n37 RST.n34 0.0361897
R1439 RST.n41 RST.n32 0.0305
R1440 RST.n23 RST 0.0301733
R1441 RST.n43 RST.n42 0.0295625
R1442 RST.n5 RST 0.0293
R1443 RST.n51 RST.n46 0.0285519
R1444 RST.n55 RST.n54 0.02675
R1445 RST.n26 RST.n23 0.0253276
R1446 RST.n38 RST.n33 0.0237584
R1447 RST.n11 RST.n6 0.0230258
R1448 RST.n30 RST.n22 0.0221964
R1449 RST.n31 RST.n30 0.0221964
R1450 RST.n4 RST.n3 0.0187743
R1451 RST.n26 RST.n25 0.0160172
R1452 RST RST.n56 0.0130521
R1453 RST.n29 RST.n27 0.0127086
R1454 RST.n17 RST.n12 0.0125591
R1455 RST.n54 RST.n53 0.0115492
R1456 RST.n37 RST.n36 0.00825862
R1457 RST.n10 RST.n9 0.00515517
R1458 RST.n16 RST.n15 0.00515517
R1459 RST.n40 RST.n39 0.00454494
R1460 RST.n50 RST.n48 0.00360345
R1461 RST.n18 RST.n17 0.00353371
R1462 RST.n4 RST.n2 0.00333412
R1463 RST.n52 RST.n51 0.00283766
R1464 RST.n29 RST.n28 0.00245652
R1465 RST.n1 RST 0.0017
R1466 RST.n40 RST.n38 0.00151124
R1467 RST.n42 RST.n41 0.0014375
R1468 JK_FF_mag_4.Q.n7 JK_FF_mag_4.Q.t12 36.935
R1469 JK_FF_mag_4.Q.n6 JK_FF_mag_4.Q.t10 36.935
R1470 JK_FF_mag_4.Q.n3 JK_FF_mag_4.Q.t6 36.935
R1471 JK_FF_mag_4.Q.n4 JK_FF_mag_4.Q.t5 31.4332
R1472 JK_FF_mag_4.Q.n8 JK_FF_mag_4.Q.t7 25.4744
R1473 JK_FF_mag_4.Q.n7 JK_FF_mag_4.Q.t11 18.1962
R1474 JK_FF_mag_4.Q.n6 JK_FF_mag_4.Q.t9 18.1962
R1475 JK_FF_mag_4.Q.n3 JK_FF_mag_4.Q.t4 18.1962
R1476 JK_FF_mag_4.Q.n4 JK_FF_mag_4.Q.t3 15.3826
R1477 JK_FF_mag_4.Q.n8 JK_FF_mag_4.Q.t8 14.1417
R1478 JK_FF_mag_4.Q JK_FF_mag_4.Q.t1 7.09905
R1479 JK_FF_mag_4.Q JK_FF_mag_4.Q.n4 6.86029
R1480 JK_FF_mag_4.Q.n9 JK_FF_mag_4.Q 6.35399
R1481 JK_FF_mag_4.Q.n5 JK_FF_mag_4.Q 5.01077
R1482 JK_FF_mag_4.Q JK_FF_mag_4.Q.n2 3.25053
R1483 JK_FF_mag_4.Q.n2 JK_FF_mag_4.Q.t0 2.2755
R1484 JK_FF_mag_4.Q.n2 JK_FF_mag_4.Q.n1 2.2755
R1485 JK_FF_mag_4.Q JK_FF_mag_4.Q.n7 2.13265
R1486 JK_FF_mag_4.Q.n0 JK_FF_mag_4.Q 2.63776
R1487 JK_FF_mag_4.Q JK_FF_mag_4.Q.n9 2.3405
R1488 JK_FF_mag_4.Q JK_FF_mag_4.Q.n3 2.13459
R1489 JK_FF_mag_4.Q.n6 JK_FF_mag_4.Q 2.13261
R1490 JK_FF_mag_4.Q.n9 JK_FF_mag_4.Q.n5 1.54877
R1491 JK_FF_mag_4.Q.n0 JK_FF_mag_4.Q 2.1039
R1492 JK_FF_mag_4.Q JK_FF_mag_4.Q.n8 1.62425
R1493 JK_FF_mag_4.Q.n5 JK_FF_mag_4.Q 1.12067
R1494 JK_FF_mag_4.Q.n0 JK_FF_mag_4.Q 1.11863
R1495 JK_FF_mag_5.Q.n4 JK_FF_mag_5.Q.t6 36.935
R1496 JK_FF_mag_5.Q.n3 JK_FF_mag_5.Q.t7 36.935
R1497 JK_FF_mag_5.Q.n6 JK_FF_mag_5.Q.t10 36.935
R1498 JK_FF_mag_5.Q.n7 JK_FF_mag_5.Q.t12 31.4332
R1499 JK_FF_mag_5.Q.n5 JK_FF_mag_5.Q.t4 25.5361
R1500 JK_FF_mag_5.Q.n4 JK_FF_mag_5.Q.t3 18.1962
R1501 JK_FF_mag_5.Q.n3 JK_FF_mag_5.Q.t5 18.1962
R1502 JK_FF_mag_5.Q.n6 JK_FF_mag_5.Q.t9 18.1962
R1503 JK_FF_mag_5.Q.n7 JK_FF_mag_5.Q.t11 15.3826
R1504 JK_FF_mag_5.Q.n5 JK_FF_mag_5.Q.t8 14.0734
R1505 JK_FF_mag_5.Q JK_FF_mag_5.Q.t2 7.09905
R1506 JK_FF_mag_5.Q JK_FF_mag_5.Q.n7 6.86029
R1507 JK_FF_mag_5.Q.n8 JK_FF_mag_5.Q 5.01077
R1508 JK_FF_mag_5.Q.n9 JK_FF_mag_5.Q 4.16836
R1509 JK_FF_mag_5.Q JK_FF_mag_5.Q.n2 3.25053
R1510 JK_FF_mag_5.Q.n2 JK_FF_mag_5.Q.t0 2.2755
R1511 JK_FF_mag_5.Q.n2 JK_FF_mag_5.Q.n1 2.2755
R1512 JK_FF_mag_5.Q JK_FF_mag_5.Q.n4 2.13151
R1513 JK_FF_mag_5.Q.n0 JK_FF_mag_5.Q 2.63808
R1514 JK_FF_mag_5.Q JK_FF_mag_5.Q.n9 2.34284
R1515 JK_FF_mag_5.Q JK_FF_mag_5.Q.n6 2.13459
R1516 JK_FF_mag_5.Q JK_FF_mag_5.Q.n3 2.13042
R1517 JK_FF_mag_5.Q JK_FF_mag_5.Q.n0 2.10738
R1518 JK_FF_mag_5.Q.n9 JK_FF_mag_5.Q.n8 1.52539
R1519 JK_FF_mag_5.Q JK_FF_mag_5.Q.n5 1.43628
R1520 JK_FF_mag_5.Q.n8 JK_FF_mag_5.Q 1.12067
R1521 JK_FF_mag_5.Q JK_FF_mag_5.Q.n0 1.11863
R1522 Vdiv96.n2 Vdiv96.n1 9.33985
R1523 Vdiv96.n2 Vdiv96.n0 5.17836
R1524 Vdiv96 Vdiv96.n2 0.0749828
C0 VDD JK_FF_mag_0.Q 2.07f
C1 VDD a_8124_3745# 3.14e-19
C2 a_8842_2648# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C3 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C4 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_5.Q 0.235f
C5 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1 1.12e-19
C6 a_8278_2648# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C7 RST JK_FF_mag_4.nand2_mag_3.IN1 0.0768f
C8 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C9 JK_FF_mag_4.QB JK_FF_mag_3.Q 3.23e-19
C10 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C11 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.nand2_mag_1.IN2 0.36f
C12 RST CLK_div_3_mag_0.JK_FF_mag_1.K 0.305f
C13 JK_FF_mag_0.Q a_702_417# 0.00335f
C14 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.QB 0.199f
C15 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C16 VDD JK_FF_mag_3.nand3_mag_0.OUT 0.742f
C17 a_8469_395# JK_FF_mag_3.QB 0.00964f
C18 JK_FF_mag_4.Q a_2307_3060# 0.0101f
C19 JK_FF_mag_0.Q a_3928_351# 0.00143f
C20 a_3412_6363# JK_FF_mag_4.Q 0.0157f
C21 JK_FF_mag_4.Q JK_FF_mag_5.nand3_mag_0.OUT 0.267f
C22 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C23 JK_FF_mag_4.nand3_mag_1.OUT a_4130_5266# 4.52e-20
C24 CLK JK_FF_mag_3.Q 0.00936f
C25 JK_FF_mag_0.QB JK_FF_mag_5.nand2_mag_1.IN2 1.38e-19
C26 JK_FF_mag_5.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 5.51e-20
C27 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C28 RST a_1589_4157# 0.00103f
C29 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C30 VDD JK_FF_mag_4.nand2_mag_1.IN2 0.402f
C31 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 0.103f
C32 a_7021_351# JK_FF_mag_3.nand3_mag_1.OUT 1.17e-20
C33 JK_FF_mag_5.nand3_mag_1.OUT VDD 0.999f
C34 a_8278_2648# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C35 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_0.Q 0.235f
C36 RST JK_FF_mag_5.nand3_mag_1.IN1 0.218f
C37 JK_FF_mag_0.Q JK_FF_mag_2.nand2_mag_3.IN1 0.41f
C38 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.00167f
C39 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C40 a_3819_3701# CLK_div_3_mag_0.JK_FF_mag_1.K 8.64e-19
C41 VDD JK_FF_mag_5.Q 2.19f
C42 JK_FF_mag_4.Q a_2147_3060# 0.00939f
C43 CLK a_5418_5266# 0.0101f
C44 RST a_1429_4157# 0.00144f
C45 a_7554_2604# CLK_div_3_mag_0.Q1 3.6e-22
C46 JK_FF_mag_2.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 5.97e-20
C47 a_2153_4157# a_2313_4157# 0.0504f
C48 a_7751_1492# JK_FF_mag_3.nand3_mag_0.OUT 0.00378f
C49 a_702_417# JK_FF_mag_5.Q 0.00117f
C50 a_8124_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C51 VDD a_5424_6363# 0.00108f
C52 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C53 JK_FF_mag_3.Q CLK_div_3_mag_0.Q1 1.02f
C54 JK_FF_mag_4.Q CLK_div_3_mag_0.JK_FF_mag_1.QB 2.73e-21
C55 RST JK_FF_mag_2.nand3_mag_0.OUT 0.00571f
C56 RST a_7272_4844# 4.93e-19
C57 JK_FF_mag_4.QB a_5258_5266# 0.00392f
C58 JK_FF_mag_2.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 6.48e-19
C59 JK_FF_mag_4.nand3_mag_1.OUT a_4540_6363# 0.0733f
C60 RST JK_FF_mag_4.nand3_mag_2.OUT 0.0877f
C61 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.471f
C62 JK_FF_mag_4.Q a_1583_3060# 6.43e-21
C63 RST JK_FF_mag_0.nand3_mag_0.OUT 0.0134f
C64 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.Q 0.0343f
C65 CLK a_5258_5266# 0.00939f
C66 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_5.nand3_mag_0.OUT 0.0622f
C67 a_1583_3060# JK_FF_mag_0.nand3_mag_1.OUT 3.64e-20
C68 a_8245_5080# CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C69 JK_FF_mag_4.nand3_mag_1.OUT VDD 0.999f
C70 RST CLK_div_3_mag_0.Q0 0.044f
C71 a_6990_2604# CLK_div_3_mag_0.Q1 1.86e-20
C72 JK_FF_mag_3.nand2_mag_3.IN1 a_6830_2604# 9.14e-19
C73 JK_FF_mag_3.QB CLK_div_3_mag_0.JK_FF_mag_1.K 4.41e-19
C74 a_1432_1558# JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C75 VDD JK_FF_mag_0.nand3_mag_1.IN1 0.662f
C76 JK_FF_mag_3.nand3_mag_0.OUT a_7187_1448# 0.0732f
C77 JK_FF_mag_2.nand3_mag_1.OUT a_4652_351# 0.0203f
C78 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00205f
C79 a_1426_417# JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C80 JK_FF_mag_5.nand2_mag_3.IN1 a_455_3060# 0.00118f
C81 JK_FF_mag_5.nand2_mag_3.IN1 a_2560_1558# 2.73e-19
C82 JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.3e-19
C83 JK_FF_mag_3.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 3.12e-19
C84 JK_FF_mag_5.nand3_mag_0.OUT JK_FF_mag_5.Q 8.73e-19
C85 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.298f
C86 a_6990_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C87 JK_FF_mag_2.QB JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C88 JK_FF_mag_4.QB a_4694_5266# 3.08e-19
C89 JK_FF_mag_0.Q a_868_1514# 2.79e-20
C90 a_3934_1448# a_4094_1448# 0.0504f
C91 JK_FF_mag_4.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 1.34e-19
C92 JK_FF_mag_4.nand3_mag_1.OUT a_3976_6363# 0.00378f
C93 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C94 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand3_mag_0.OUT 0.122f
C95 JK_FF_mag_0.QB a_2560_1558# 0.0114f
C96 a_3973_2604# JK_FF_mag_3.Q 0.00164f
C97 JK_FF_mag_4.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 5.23e-20
C98 a_4540_6363# a_4700_6363# 0.0504f
C99 JK_FF_mag_0.Q JK_FF_mag_2.Q 0.155f
C100 CLK a_4694_5266# 6.43e-21
C101 JK_FF_mag_0.Q a_1426_417# 0.0102f
C102 VDD a_3566_5266# 3.56e-19
C103 a_2150_461# JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C104 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.Q 0.064f
C105 a_8245_5080# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00168f
C106 JK_FF_mag_3.nand3_mag_0.OUT a_7027_1448# 0.0203f
C107 JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 0.194f
C108 a_2147_3060# JK_FF_mag_5.Q 2.79e-20
C109 VDD a_4700_6363# 2.21e-19
C110 JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 6.33e-20
C111 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_2.Q 0.267f
C112 a_7021_351# JK_FF_mag_3.Q 0.00335f
C113 JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 1.32e-19
C114 JK_FF_mag_4.QB a_4130_5266# 2.96e-19
C115 JK_FF_mag_0.Q JK_FF_mag_2.QB 0.307f
C116 JK_FF_mag_5.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.00137f
C117 JK_FF_mag_2.nand3_mag_1.OUT a_5222_1492# 4.52e-20
C118 a_7745_351# JK_FF_mag_3.nand3_mag_1.OUT 0.0203f
C119 JK_FF_mag_0.QB a_1996_1558# 2.96e-19
C120 a_3813_2604# JK_FF_mag_3.Q 0.00117f
C121 a_4697_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C122 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C123 JK_FF_mag_5.nand3_mag_1.OUT a_1583_3060# 0.0202f
C124 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_2.QB 2.53e-20
C125 VDD a_6830_2604# 0.00743f
C126 JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00132f
C127 JK_FF_mag_5.QB VDD 0.914f
C128 a_5671_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C129 JK_FF_mag_5.nand2_mag_3.IN1 RST 0.0546f
C130 a_868_1514# JK_FF_mag_5.Q 0.00939f
C131 VDD CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.466f
C132 RST JK_FF_mag_5.nand3_mag_2.OUT 0.0544f
C133 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.Q1 0.00335f
C134 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C135 a_5940_395# JK_FF_mag_2.nand2_mag_4.IN2 0.00372f
C136 JK_FF_mag_0.nand3_mag_2.OUT a_1586_417# 2.88e-20
C137 RST JK_FF_mag_0.QB 0.227f
C138 JK_FF_mag_3.QB CLK_div_3_mag_0.Q0 0.0015f
C139 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C140 JK_FF_mag_2.nand3_mag_1.OUT a_4658_1492# 0.0202f
C141 JK_FF_mag_0.QB a_1432_1558# 3.33e-19
C142 JK_FF_mag_5.nand3_mag_1.OUT a_1019_3060# 4.52e-20
C143 VDD a_5825_2648# 0.00149f
C144 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_3.Q 1.07e-19
C145 a_5107_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C146 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00481f
C147 JK_FF_mag_4.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 4.46e-20
C148 JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand3_mag_2.OUT 0.00118f
C149 RST CLK_div_3_mag_0.or_2_mag_0.IN2 9.76e-19
C150 JK_FF_mag_4.nand2_mag_4.IN2 JK_FF_mag_4.Q 0.0635f
C151 JK_FF_mag_4.QB a_4540_6363# 0.00696f
C152 a_1429_4157# a_1589_4157# 0.0504f
C153 JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_3_mag_0.Q1 4.49e-20
C154 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C155 JK_FF_mag_4.nand3_mag_1.OUT a_4543_3745# 3.53e-20
C156 JK_FF_mag_4.Q JK_FF_mag_0.nand2_mag_1.IN2 1.87e-19
C157 JK_FF_mag_5.QB JK_FF_mag_5.nand3_mag_0.OUT 0.343f
C158 RST JK_FF_mag_3.nand3_mag_1.OUT 0.258f
C159 CLK_div_3_mag_0.Q0 a_8245_5080# 0.0134f
C160 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C161 a_1429_4157# JK_FF_mag_5.nand3_mag_1.IN1 8.64e-19
C162 JK_FF_mag_4.QB VDD 0.917f
C163 JK_FF_mag_0.Q a_4658_1492# 6.43e-21
C164 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C165 VDD JK_FF_mag_0.nand2_mag_3.IN1 1.28f
C166 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.37f
C167 VDD a_5261_2648# 0.00149f
C168 JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00126f
C169 a_4543_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.43e-19
C170 CLK VDD 1.12f
C171 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C172 JK_FF_mag_4.QB a_3976_6363# 0.00964f
C173 VDD a_5376_395# 3.14e-19
C174 a_7560_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C175 JK_FF_mag_5.nand2_mag_4.IN2 a_865_4157# 0.069f
C176 a_2313_4157# JK_FF_mag_5.nand3_mag_2.OUT 0.0202f
C177 RST JK_FF_mag_4.nand3_mag_0.OUT 0.00942f
C178 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_5.nand3_mag_1.IN1 0.00137f
C179 JK_FF_mag_0.Q JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C180 JK_FF_mag_5.QB a_2147_3060# 0.00392f
C181 VDD JK_FF_mag_2.nand2_mag_4.IN2 0.391f
C182 a_6830_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C183 a_7745_351# JK_FF_mag_3.Q 0.0102f
C184 JK_FF_mag_0.Q a_4094_1448# 0.00939f
C185 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.or_2_mag_0.IN2 4.52e-20
C186 VDD a_4697_2604# 9.82e-19
C187 JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.35e-19
C188 a_8469_395# JK_FF_mag_3.nand3_mag_1.OUT 0.00378f
C189 a_3979_3701# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00119f
C190 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.00206f
C191 a_6996_3701# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00119f
C192 JK_FF_mag_4.QB a_3412_6363# 0.0811f
C193 JK_FF_mag_5.nand2_mag_3.IN1 a_2153_4157# 1.46e-19
C194 JK_FF_mag_4.nand2_mag_4.IN2 JK_FF_mag_4.nand2_mag_1.IN2 8.16e-20
C195 JK_FF_mag_5.nand3_mag_0.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.0017f
C196 a_2153_4157# JK_FF_mag_5.nand3_mag_2.OUT 0.0731f
C197 a_7021_351# JK_FF_mag_3.nand3_mag_2.OUT 0.0202f
C198 JK_FF_mag_2.nand2_mag_3.IN1 a_5261_2648# 5.3e-20
C199 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C200 RST a_7714_2604# 0.00121f
C201 JK_FF_mag_3.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.08e-19
C202 JK_FF_mag_0.nand2_mag_4.IN2 a_2150_461# 0.069f
C203 VDD CLK_div_3_mag_0.Q1 2.48f
C204 JK_FF_mag_5.QB a_1583_3060# 2.25e-19
C205 a_5376_395# JK_FF_mag_2.nand2_mag_3.IN1 0.0036f
C206 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.or_2_mag_0.IN2 0.0445f
C207 Vdiv96 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1e-19
C208 JK_FF_mag_0.Q a_3934_1448# 0.0101f
C209 a_6836_3701# CLK_div_3_mag_0.Q1 0.00149f
C210 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C211 VDD a_4537_2604# 0.0012f
C212 CLK_div_3_mag_0.JK_FF_mag_1.K JK_FF_mag_5.nand3_mag_2.OUT 2.82e-21
C213 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C214 JK_FF_mag_4.nand3_mag_1.IN1 a_4694_5266# 0.0697f
C215 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_5.Q 1.48e-20
C216 a_5825_2648# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0811f
C217 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C218 JK_FF_mag_4.QB a_5107_3745# 2.05e-20
C219 a_4694_5266# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 3.53e-20
C220 a_8278_2648# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C221 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_1.OUT 0.25f
C222 JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 9.38e-20
C223 a_2147_3060# JK_FF_mag_0.nand2_mag_3.IN1 3.23e-20
C224 a_1589_4157# JK_FF_mag_5.nand3_mag_2.OUT 9.1e-19
C225 RST a_7554_2604# 0.00141f
C226 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C227 a_8315_1492# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.63e-20
C228 JK_FF_mag_5.QB a_1019_3060# 2.96e-19
C229 JK_FF_mag_5.nand3_mag_1.OUT a_865_4157# 0.00378f
C230 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.652f
C231 RST JK_FF_mag_3.Q 0.23f
C232 a_8245_5080# CLK_div_3_mag_0.or_2_mag_0.IN2 8.64e-19
C233 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.nand3_mag_1.IN1 0.233f
C234 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.394f
C235 JK_FF_mag_5.nand3_mag_1.IN1 JK_FF_mag_5.nand3_mag_2.OUT 0.00164f
C236 a_8879_1492# JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C237 a_5671_3745# CLK_div_3_mag_0.Q1 0.069f
C238 JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.Q1 1.1e-19
C239 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand2_mag_4.IN2 0.122f
C240 VDD a_3973_2604# 0.00888f
C241 JK_FF_mag_4.Q CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 5.69e-19
C242 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.or_2_mag_0.IN2 0.00761f
C243 JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00109f
C244 JK_FF_mag_4.nand3_mag_1.IN1 a_4130_5266# 0.0059f
C245 a_865_4157# JK_FF_mag_5.Q 0.00859f
C246 JK_FF_mag_0.QB JK_FF_mag_5.nand3_mag_1.IN1 1.4e-19
C247 a_5261_2648# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00964f
C248 a_868_1514# JK_FF_mag_0.nand2_mag_3.IN1 0.00119f
C249 VDD a_2714_461# 3.54e-19
C250 a_7714_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C251 a_8842_2648# CLK_div_3_mag_0.JK_FF_mag_1.K 0.0811f
C252 CLK CLK_div_3_mag_0.JK_FF_mag_1.QB 1.2e-19
C253 JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00105f
C254 VDD JK_FF_mag_3.nand2_mag_4.IN2 0.391f
C255 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C256 RST JK_FF_mag_3.nand3_mag_1.IN1 0.153f
C257 JK_FF_mag_2.QB a_5825_2648# 5.3e-20
C258 a_1429_4157# JK_FF_mag_5.nand3_mag_2.OUT 2.88e-20
C259 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C260 RST a_6990_2604# 0.00254f
C261 JK_FF_mag_3.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 6.87e-20
C262 a_1426_417# a_1586_417# 0.0504f
C263 VDD a_7021_351# 0.00108f
C264 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C265 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.Q1 6.7e-19
C266 RST a_5418_5266# 0.00173f
C267 a_3819_3701# JK_FF_mag_3.Q 0.0101f
C268 JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand3_mag_0.OUT 0.0884f
C269 JK_FF_mag_4.nand2_mag_4.IN2 a_3566_5266# 4.52e-20
C270 JK_FF_mag_0.Q CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 3.42e-20
C271 a_5376_395# JK_FF_mag_2.Q 0.00859f
C272 a_8469_395# JK_FF_mag_3.Q 0.00859f
C273 VDD a_3813_2604# 0.0133f
C274 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_0.OUT 0.0017f
C275 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C276 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_0.QB 1.7e-19
C277 VDD JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C278 a_4697_2604# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00696f
C279 JK_FF_mag_4.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.00392f
C280 a_7554_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C281 a_8278_2648# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00964f
C282 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 9.98e-19
C283 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C284 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C285 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00305f
C286 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.Q 0.0635f
C287 VDD JK_FF_mag_5.nand2_mag_1.IN2 0.408f
C288 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.0725f
C289 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C290 a_5376_395# JK_FF_mag_2.QB 0.00964f
C291 RST a_5258_5266# 0.0013f
C292 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 1.94f
C293 a_7021_351# a_7181_351# 0.0504f
C294 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_1.IN2 1.85e-19
C295 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_3.Q 5.57e-19
C296 a_7745_351# JK_FF_mag_3.nand3_mag_2.OUT 9.1e-19
C297 a_4540_6363# JK_FF_mag_4.nand3_mag_1.IN1 8.64e-19
C298 JK_FF_mag_0.nand3_mag_2.OUT a_862_417# 0.0731f
C299 JK_FF_mag_0.Q JK_FF_mag_2.nand3_mag_1.OUT 6.64e-19
C300 CLK_div_3_mag_0.or_2_mag_0.IN2 a_7272_4844# 7.48e-20
C301 JK_FF_mag_4.Q JK_FF_mag_0.Q 0.00927f
C302 JK_FF_mag_2.QB JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C303 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C304 JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00105f
C305 JK_FF_mag_3.QB JK_FF_mag_3.Q 1.98f
C306 a_4537_2604# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00695f
C307 Vdiv96 CLK_div_3_mag_0.Q1 2.53e-19
C308 a_6990_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C309 JK_FF_mag_0.Q JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C310 JK_FF_mag_2.nand2_mag_4.IN2 a_5786_1492# 4.52e-20
C311 a_7714_2604# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00696f
C312 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN JK_FF_mag_3.Q 7.03e-21
C313 JK_FF_mag_4.nand3_mag_1.IN1 VDD 0.656f
C314 JK_FF_mag_2.Q CLK_div_3_mag_0.Q1 4.57e-20
C315 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.01f
C316 JK_FF_mag_5.QB JK_FF_mag_0.nand2_mag_1.IN2 1.38e-19
C317 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.IN2 0.0655f
C318 a_8842_2648# CLK_div_3_mag_0.Q0 0.0157f
C319 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.196f
C320 RST a_4694_5266# 3.52e-19
C321 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C322 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C323 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_1.IN1 0.0387f
C324 VDD a_708_1514# 0.00534f
C325 JK_FF_mag_3.nand3_mag_1.OUT CLK_div_3_mag_0.Q0 4.55e-20
C326 JK_FF_mag_2.QB CLK_div_3_mag_0.Q1 0.00139f
C327 a_3979_3701# CLK_div_3_mag_0.Q1 2.79e-20
C328 JK_FF_mag_5.nand2_mag_4.IN2 JK_FF_mag_5.nand3_mag_1.OUT 0.122f
C329 a_4543_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00378f
C330 RST a_2150_461# 0.00112f
C331 JK_FF_mag_4.Q JK_FF_mag_4.nand2_mag_1.IN2 0.108f
C332 JK_FF_mag_4.nand3_mag_2.OUT JK_FF_mag_4.nand3_mag_0.OUT 0.00183f
C333 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_4.Q 6.64e-19
C334 a_7554_2604# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00695f
C335 JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_3.Q 0.00293f
C336 JK_FF_mag_5.QB a_865_4157# 0.00964f
C337 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.00162f
C338 JK_FF_mag_5.nand2_mag_4.IN2 JK_FF_mag_5.Q 0.0635f
C339 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.nand3_mag_2.OUT 0.00118f
C340 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.K 2.09f
C341 VDD JK_FF_mag_2.nand2_mag_1.IN2 0.402f
C342 RST JK_FF_mag_2.nand3_mag_1.IN1 0.195f
C343 JK_FF_mag_4.Q JK_FF_mag_5.Q 0.161f
C344 RST a_5940_395# 0.00101f
C345 JK_FF_mag_4.QB JK_FF_mag_4.nand2_mag_4.IN2 0.199f
C346 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_0.QB 0.00999f
C347 a_8278_2648# CLK_div_3_mag_0.Q0 0.00859f
C348 RST JK_FF_mag_3.nand3_mag_2.OUT 0.0884f
C349 RST a_4130_5266# 5.97e-19
C350 JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 2.89e-20
C351 a_702_417# a_862_417# 0.0504f
C352 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_5.Q 9.24e-19
C353 VDD a_7745_351# 2.21e-19
C354 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q0 0.107f
C355 RST JK_FF_mag_3.nand2_mag_3.IN1 0.0196f
C356 VDD a_455_3060# 3.6e-19
C357 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C358 a_3979_3701# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C359 a_3928_351# a_4088_351# 0.0504f
C360 JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 4.3e-20
C361 VDD a_2560_1558# 3.76e-19
C362 JK_FF_mag_4.Q a_5424_6363# 0.00335f
C363 RST a_7560_3745# 3.41e-19
C364 a_7021_351# JK_FF_mag_2.Q 0.00179f
C365 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C366 RST JK_FF_mag_0.nand3_mag_2.OUT 0.0585f
C367 JK_FF_mag_0.Q JK_FF_mag_5.Q 0.149f
C368 a_4812_351# JK_FF_mag_2.nand3_mag_1.IN1 8.64e-19
C369 a_7714_2604# CLK_div_3_mag_0.Q0 0.0101f
C370 JK_FF_mag_2.nand3_mag_2.OUT a_4088_351# 0.0731f
C371 a_5107_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C372 a_4088_351# JK_FF_mag_2.nand2_mag_3.IN1 1.46e-19
C373 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.Q 0.0343f
C374 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_1.IN2 0.36f
C375 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C376 JK_FF_mag_4.Q a_5264_6363# 0.00789f
C377 VDD a_1996_1558# 3.19e-19
C378 RST a_6996_3701# 0.00156f
C379 JK_FF_mag_4.nand2_mag_3.IN1 a_5258_5266# 0.00119f
C380 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_3.Q 2.57e-19
C381 JK_FF_mag_3.Q a_7272_4844# 0.0103f
C382 JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 1.34e-19
C383 a_8469_395# JK_FF_mag_3.nand2_mag_3.IN1 0.0036f
C384 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C385 a_4540_6363# RST 0.00189f
C386 JK_FF_mag_4.Q CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 9.6e-19
C387 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C388 a_7554_2604# CLK_div_3_mag_0.Q0 0.0102f
C389 a_4543_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0202f
C390 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_5.Q 0.0345f
C391 JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.08e-20
C392 JK_FF_mag_4.Q a_3566_5266# 0.069f
C393 JK_FF_mag_0.Q JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C394 RST VDD 3.15f
C395 CLK_div_3_mag_0.Q0 JK_FF_mag_3.Q 0.502f
C396 JK_FF_mag_4.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.32e-19
C397 JK_FF_mag_5.nand2_mag_1.IN2 a_1019_3060# 0.069f
C398 a_7560_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C399 a_4094_1448# CLK_div_3_mag_0.Q1 2.37e-20
C400 VDD a_1432_1558# 3.19e-19
C401 JK_FF_mag_4.Q a_4700_6363# 0.0102f
C402 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C403 a_708_1514# a_868_1514# 0.0504f
C404 JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 4.41e-20
C405 RST a_6836_3701# 0.00217f
C406 JK_FF_mag_4.nand2_mag_3.IN1 a_4694_5266# 1.43e-19
C407 CLK CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.8e-19
C408 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C409 a_3976_6363# RST 0.00101f
C410 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C411 RST a_3928_351# 0.00193f
C412 JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_3_mag_0.Q0 6.24e-20
C413 JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 6.43e-20
C414 JK_FF_mag_5.nand2_mag_4.IN2 JK_FF_mag_5.QB 0.199f
C415 a_6990_2604# CLK_div_3_mag_0.Q0 0.00707f
C416 JK_FF_mag_5.QB JK_FF_mag_4.Q 0.307f
C417 RST a_7181_351# 0.00193f
C418 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand2_mag_1.IN2 0.00975f
C419 VDD a_3819_3701# 5.99e-19
C420 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 2.62e-19
C421 JK_FF_mag_5.QB JK_FF_mag_0.nand3_mag_1.OUT 4.51e-20
C422 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.or_2_mag_0.IN2 3.81e-19
C423 RST JK_FF_mag_2.nand3_mag_2.OUT 0.0856f
C424 a_4088_351# JK_FF_mag_2.Q 0.00789f
C425 VDD a_8469_395# 3.14e-19
C426 RST a_5671_3745# 0.00155f
C427 RST JK_FF_mag_2.nand2_mag_3.IN1 0.0761f
C428 JK_FF_mag_4.nand2_mag_3.IN1 a_4130_5266# 0.011f
C429 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.Q 0.107f
C430 RST a_2307_3060# 9.45e-19
C431 a_3412_6363# RST 0.00101f
C432 RST JK_FF_mag_5.nand3_mag_0.OUT 0.0145f
C433 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_5.Q 3.64e-19
C434 JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.55e-20
C435 RST a_7751_1492# 3.83e-19
C436 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.998f
C437 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1 0.107f
C438 VDD a_301_4157# 3.14e-19
C439 JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 4.33e-20
C440 a_5222_1492# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.71e-20
C441 JK_FF_mag_4.nand2_mag_1.IN2 a_3566_5266# 0.00372f
C442 JK_FF_mag_2.QB JK_FF_mag_2.nand2_mag_1.IN2 0.0592f
C443 JK_FF_mag_4.nand3_mag_1.OUT a_5424_6363# 1.17e-20
C444 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.397f
C445 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.145f
C446 a_8879_1492# JK_FF_mag_3.QB 0.0114f
C447 JK_FF_mag_3.Q JK_FF_mag_5.nand3_mag_2.OUT 3.81e-20
C448 a_7560_3745# CLK_div_3_mag_0.JK_FF_mag_1.K 1.75e-19
C449 VDD a_2313_4157# 0.00108f
C450 JK_FF_mag_2.nand3_mag_2.OUT a_4812_351# 2.88e-20
C451 a_5786_1492# JK_FF_mag_2.nand2_mag_1.IN2 0.00372f
C452 a_5264_6363# a_5424_6363# 0.0504f
C453 RST a_5107_3745# 7.14e-19
C454 VDD JK_FF_mag_3.QB 0.902f
C455 a_7745_351# a_7905_351# 0.0504f
C456 RST a_7187_1448# 0.00182f
C457 RST a_2147_3060# 0.00102f
C458 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C459 VDD CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C460 JK_FF_mag_4.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 1.14e-20
C461 JK_FF_mag_4.QB JK_FF_mag_4.Q 1.96f
C462 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C463 JK_FF_mag_4.Q JK_FF_mag_0.nand2_mag_3.IN1 6.08e-19
C464 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C465 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C466 a_4697_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C467 a_1586_417# JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C468 CLK JK_FF_mag_4.Q 0.149f
C469 JK_FF_mag_4.nand3_mag_1.OUT a_5264_6363# 1.5e-20
C470 a_5376_395# JK_FF_mag_2.nand3_mag_1.OUT 0.00378f
C471 RST CLK_div_3_mag_0.JK_FF_mag_1.QB 0.602f
C472 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 0.101f
C473 a_8315_1492# JK_FF_mag_3.QB 2.96e-19
C474 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_5.QB 0.248f
C475 a_6996_3701# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00392f
C476 JK_FF_mag_3.Q CLK_div_3_mag_0.or_2_mag_0.IN2 6.62e-20
C477 a_5222_1492# JK_FF_mag_2.nand2_mag_1.IN2 0.069f
C478 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_5.nand3_mag_1.IN1 1.53e-20
C479 JK_FF_mag_4.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 2.19e-20
C480 RST a_868_1514# 9.48e-19
C481 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 0.338f
C482 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C483 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_5671_3745# 4.52e-20
C484 JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 9.28e-20
C485 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C486 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C487 JK_FF_mag_5.QB JK_FF_mag_5.Q 1.97f
C488 RST a_7027_1448# 0.00242f
C489 RST a_1583_3060# 0.00248f
C490 VDD a_8245_5080# 0.165f
C491 JK_FF_mag_4.nand2_mag_3.IN1 VDD 1.24f
C492 JK_FF_mag_0.Q JK_FF_mag_0.nand2_mag_3.IN1 0.0171f
C493 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.Q 0.0358f
C494 JK_FF_mag_0.Q a_1586_417# 0.0101f
C495 RST JK_FF_mag_2.Q 0.312f
C496 VDD CLK_div_3_mag_0.JK_FF_mag_1.K 2.58f
C497 JK_FF_mag_2.nand3_mag_1.OUT a_4697_2604# 3.87e-20
C498 RST a_1426_417# 8.64e-19
C499 a_4537_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C500 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C501 RST a_4652_351# 0.00172f
C502 JK_FF_mag_4.nand3_mag_1.OUT a_4700_6363# 0.0203f
C503 JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 2.45e-19
C504 a_7751_1492# JK_FF_mag_3.QB 3.33e-19
C505 a_3976_6363# JK_FF_mag_4.nand2_mag_3.IN1 0.0036f
C506 VDD a_1589_4157# 2.21e-19
C507 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C508 JK_FF_mag_4.nand3_mag_0.OUT JK_FF_mag_3.Q 1.45e-19
C509 JK_FF_mag_2.nand3_mag_1.OUT CLK_div_3_mag_0.Q1 6.72e-20
C510 RST JK_FF_mag_2.QB 0.255f
C511 JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.Q0 1.35e-19
C512 RST a_7905_351# 0.00157f
C513 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C514 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C515 RST a_5786_1492# 0.0019f
C516 JK_FF_mag_4.Q CLK_div_3_mag_0.Q1 9.66e-19
C517 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C518 RST a_1019_3060# 0.001f
C519 a_4812_351# JK_FF_mag_2.Q 0.0101f
C520 VDD JK_FF_mag_5.nand3_mag_1.IN1 0.661f
C521 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_3.Q 7.81e-19
C522 JK_FF_mag_3.nand2_mag_4.IN2 a_9033_395# 0.00372f
C523 JK_FF_mag_4.QB JK_FF_mag_4.nand2_mag_1.IN2 0.0592f
C524 a_8688_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C525 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_3.IN1 7.06e-19
C526 JK_FF_mag_5.QB JK_FF_mag_0.nand3_mag_1.IN1 1.4e-19
C527 a_4652_351# a_4812_351# 0.0504f
C528 a_3973_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C529 JK_FF_mag_3.QB a_7187_1448# 0.00392f
C530 JK_FF_mag_3.nand3_mag_1.IN1 a_8278_2648# 4.58e-20
C531 CLK JK_FF_mag_4.nand2_mag_1.IN2 1.48e-20
C532 a_7554_2604# a_7714_2604# 0.0504f
C533 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.175f
C534 JK_FF_mag_3.QB CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.06e-19
C535 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_5.Q 0.426f
C536 JK_FF_mag_2.QB a_4812_351# 0.00696f
C537 JK_FF_mag_4.nand3_mag_0.OUT a_5418_5266# 0.0203f
C538 a_4540_6363# JK_FF_mag_4.nand3_mag_2.OUT 2.88e-20
C539 JK_FF_mag_0.Q CLK_div_3_mag_0.Q1 0.00107f
C540 RST a_5222_1492# 0.00101f
C541 JK_FF_mag_4.Q CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 1.48e-20
C542 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C543 a_2560_1558# JK_FF_mag_0.nand2_mag_1.IN2 0.00372f
C544 a_3979_3701# a_3819_3701# 0.0504f
C545 a_6996_3701# CLK_div_3_mag_0.Q0 2.79e-20
C546 VDD JK_FF_mag_2.nand3_mag_0.OUT 0.746f
C547 VDD a_7272_4844# 5.92e-19
C548 a_8688_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C549 JK_FF_mag_2.Q CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 1.11e-19
C550 JK_FF_mag_4.nand3_mag_2.OUT VDD 0.752f
C551 a_8124_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C552 a_8879_1492# CLK_div_3_mag_0.Q0 1.63e-20
C553 JK_FF_mag_0.QB a_2150_461# 0.00964f
C554 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C555 a_3813_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C556 VDD JK_FF_mag_0.nand3_mag_0.OUT 0.765f
C557 CLK a_5424_6363# 0.00117f
C558 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN Vdiv96 0.127f
C559 VDD CLK_div_3_mag_0.Q0 1.23f
C560 JK_FF_mag_3.QB JK_FF_mag_2.Q 0.307f
C561 JK_FF_mag_5.nand3_mag_0.OUT JK_FF_mag_5.nand3_mag_1.IN1 0.122f
C562 JK_FF_mag_4.nand3_mag_0.OUT a_5258_5266# 0.0732f
C563 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.QB 0.25f
C564 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.0881f
C565 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C566 a_5786_1492# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 1.71e-20
C567 RST a_4658_1492# 3.73e-19
C568 a_1586_417# JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C569 a_1996_1558# JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C570 JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_3_mag_0.Q0 6.24e-20
C571 JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00182f
C572 JK_FF_mag_4.nand3_mag_1.OUT CLK 6.64e-19
C573 JK_FF_mag_3.QB JK_FF_mag_2.QB 2.36e-21
C574 JK_FF_mag_0.Q a_3973_2604# 3.87e-20
C575 a_7905_351# JK_FF_mag_3.QB 0.00696f
C576 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C577 RST JK_FF_mag_4.nand2_mag_4.IN2 0.0232f
C578 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C579 JK_FF_mag_4.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00182f
C580 JK_FF_mag_0.Q a_2714_461# 0.0157f
C581 JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 1.14e-20
C582 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.0889f
C583 CLK a_5264_6363# 0.00164f
C584 JK_FF_mag_5.nand2_mag_4.IN2 JK_FF_mag_5.nand2_mag_1.IN2 8.16e-20
C585 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.QB 0.103f
C586 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C587 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C588 a_5261_2648# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C589 JK_FF_mag_4.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00132f
C590 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.Q 0.00732f
C591 RST JK_FF_mag_0.nand2_mag_1.IN2 0.0112f
C592 JK_FF_mag_4.Q JK_FF_mag_5.nand2_mag_1.IN2 1.48e-20
C593 JK_FF_mag_4.nand3_mag_0.OUT a_4694_5266# 0.00378f
C594 Vdiv96 CLK_div_3_mag_0.JK_FF_mag_1.K 4.46e-19
C595 CLK CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.96e-19
C596 JK_FF_mag_4.QB a_3566_5266# 0.0114f
C597 a_6990_2604# JK_FF_mag_3.Q 0.0108f
C598 RST a_4094_1448# 7.66e-19
C599 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C600 JK_FF_mag_4.QB a_4700_6363# 0.00695f
C601 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C602 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.Q 0.0635f
C603 JK_FF_mag_4.nand2_mag_3.IN1 a_3979_3701# 3.13e-20
C604 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.Q 0.00358f
C605 JK_FF_mag_2.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.53e-20
C606 a_1583_3060# JK_FF_mag_5.nand3_mag_1.IN1 0.0697f
C607 JK_FF_mag_5.nand2_mag_3.IN1 VDD 1.28f
C608 VDD JK_FF_mag_5.nand3_mag_2.OUT 0.751f
C609 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C610 JK_FF_mag_5.QB JK_FF_mag_0.nand2_mag_3.IN1 0.00999f
C611 RST a_3934_1448# 9.2e-19
C612 VDD JK_FF_mag_0.QB 0.926f
C613 JK_FF_mag_2.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 6.61e-20
C614 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.Q1 0.0169f
C615 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 0.333f
C616 CLK CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.37e-20
C617 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00543f
C618 a_1019_3060# JK_FF_mag_5.nand3_mag_1.IN1 0.0059f
C619 a_868_1514# JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C620 JK_FF_mag_4.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 5.23e-20
C621 JK_FF_mag_2.nand3_mag_1.OUT a_4088_351# 1.5e-20
C622 VDD CLK_div_3_mag_0.or_2_mag_0.IN2 0.49f
C623 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.Q 7.24e-19
C624 a_862_417# JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C625 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C626 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_5.nand2_mag_1.IN2 0.00975f
C627 VDD a_8842_2648# 3.14e-19
C628 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.013f
C629 a_5258_5266# a_5418_5266# 0.0504f
C630 a_7027_1448# CLK_div_3_mag_0.Q0 1.01e-20
C631 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.nand3_mag_0.OUT 0.0888f
C632 JK_FF_mag_5.nand2_mag_4.IN2 a_455_3060# 4.52e-20
C633 CLK_div_3_mag_0.Q0 Vdiv96 0.00838f
C634 VDD JK_FF_mag_3.nand3_mag_1.OUT 0.994f
C635 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C636 JK_FF_mag_5.nand3_mag_0.OUT JK_FF_mag_5.nand3_mag_2.OUT 0.00183f
C637 JK_FF_mag_5.nand2_mag_1.IN2 JK_FF_mag_5.Q 0.109f
C638 a_8842_2648# JK_FF_mag_3.nand2_mag_1.IN2 4.58e-20
C639 JK_FF_mag_2.Q CLK_div_3_mag_0.Q0 0.00113f
C640 JK_FF_mag_0.QB JK_FF_mag_2.nand2_mag_3.IN1 5.83e-19
C641 JK_FF_mag_2.QB JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C642 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C643 JK_FF_mag_0.Q a_862_417# 0.00789f
C644 a_6830_2604# CLK_div_3_mag_0.Q1 2.55e-20
C645 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand2_mag_1.IN2 0.109f
C646 a_3973_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C647 JK_FF_mag_0.Q a_4088_351# 0.00185f
C648 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.305f
C649 a_8315_1492# JK_FF_mag_3.nand3_mag_1.OUT 4.52e-20
C650 JK_FF_mag_0.Q JK_FF_mag_2.nand2_mag_1.IN2 1.48e-20
C651 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00544f
C652 JK_FF_mag_4.nand2_mag_4.IN2 JK_FF_mag_4.nand2_mag_3.IN1 0.321f
C653 JK_FF_mag_4.QB CLK 0.307f
C654 VDD JK_FF_mag_4.nand3_mag_0.OUT 0.746f
C655 VDD a_8278_2648# 3.14e-19
C656 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.Q 0.338f
C657 JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 1.81e-19
C658 JK_FF_mag_5.nand2_mag_3.IN1 a_2147_3060# 0.00119f
C659 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0545f
C660 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C661 a_7181_351# JK_FF_mag_3.nand3_mag_1.OUT 1.5e-20
C662 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C663 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.Q 0.296f
C664 JK_FF_mag_0.Q a_2560_1558# 0.069f
C665 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C666 a_5825_2648# CLK_div_3_mag_0.Q1 0.0157f
C667 a_7560_3745# JK_FF_mag_3.Q 6.43e-21
C668 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_2.OUT 0.00167f
C669 a_1996_1558# JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C670 a_708_1514# JK_FF_mag_5.Q 0.0101f
C671 a_7751_1492# JK_FF_mag_3.nand3_mag_1.OUT 0.0202f
C672 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.or_2_mag_0.IN2 1.82e-19
C673 a_5376_395# JK_FF_mag_2.nand2_mag_4.IN2 0.069f
C674 JK_FF_mag_5.nand2_mag_4.IN2 RST 0.00125f
C675 JK_FF_mag_5.nand2_mag_3.IN1 a_868_1514# 3.23e-20
C676 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand2_mag_3.IN1 0.233f
C677 RST JK_FF_mag_2.nand3_mag_1.OUT 0.286f
C678 JK_FF_mag_5.nand2_mag_3.IN1 a_1583_3060# 1.43e-19
C679 a_862_417# JK_FF_mag_5.Q 0.00164f
C680 RST JK_FF_mag_4.Q 0.16f
C681 JK_FF_mag_0.QB a_868_1514# 0.00392f
C682 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_1.IN1 0.768f
C683 JK_FF_mag_3.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00104f
C684 RST JK_FF_mag_0.nand3_mag_1.OUT 0.39f
C685 JK_FF_mag_4.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00154f
C686 JK_FF_mag_0.Q a_1996_1558# 1.63e-20
C687 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C688 a_5261_2648# CLK_div_3_mag_0.Q1 0.00859f
C689 a_6996_3701# JK_FF_mag_3.Q 0.00959f
C690 JK_FF_mag_2.nand3_mag_0.OUT a_4658_1492# 0.00378f
C691 JK_FF_mag_0.QB JK_FF_mag_2.Q 7.83e-20
C692 a_1432_1558# JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C693 JK_FF_mag_0.QB a_1426_417# 0.00695f
C694 CLK CLK_div_3_mag_0.Q1 0.00215f
C695 a_8879_1492# JK_FF_mag_3.Q 0.0696f
C696 a_455_3060# JK_FF_mag_5.Q 0.069f
C697 JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 4.41e-20
C698 VDD a_7554_2604# 2.21e-19
C699 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C700 JK_FF_mag_2.nand3_mag_1.OUT a_4812_351# 0.0733f
C701 JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 3.55e-20
C702 RST JK_FF_mag_0.Q 0.141f
C703 JK_FF_mag_3.QB a_9033_395# 0.0811f
C704 JK_FF_mag_5.nand2_mag_3.IN1 a_1019_3060# 0.011f
C705 VDD JK_FF_mag_3.Q 4f
C706 JK_FF_mag_2.QB JK_FF_mag_0.QB 6.67e-20
C707 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C708 JK_FF_mag_4.Q a_3819_3701# 7.32e-19
C709 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C710 JK_FF_mag_0.QB a_1019_3060# 2.12e-20
C711 JK_FF_mag_5.QB JK_FF_mag_5.nand2_mag_1.IN2 0.0592f
C712 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.Q 0.118f
C713 a_6836_3701# JK_FF_mag_3.Q 0.0101f
C714 a_4697_2604# CLK_div_3_mag_0.Q1 0.0101f
C715 RST JK_FF_mag_3.nand3_mag_0.OUT 0.014f
C716 JK_FF_mag_2.nand3_mag_0.OUT a_4094_1448# 0.0732f
C717 VDD JK_FF_mag_3.nand3_mag_1.IN1 0.651f
C718 JK_FF_mag_5.nand2_mag_4.IN2 a_301_4157# 0.00372f
C719 JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.35e-20
C720 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_2.Q 6.64e-19
C721 VDD a_6990_2604# 3.1e-20
C722 a_7714_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C723 a_4537_2604# a_4697_2604# 0.0504f
C724 VDD a_5418_5266# 0.00533f
C725 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C726 RST JK_FF_mag_4.nand2_mag_1.IN2 0.00425f
C727 JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.27e-20
C728 a_7181_351# JK_FF_mag_3.Q 0.00789f
C729 JK_FF_mag_5.nand3_mag_1.OUT RST 0.376f
C730 JK_FF_mag_4.Q a_2313_4157# 0.0022f
C731 a_8315_1492# JK_FF_mag_3.nand3_mag_1.IN1 0.0059f
C732 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.Q1 0.104f
C733 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C734 JK_FF_mag_2.nand3_mag_0.OUT a_3934_1448# 0.0203f
C735 JK_FF_mag_5.nand3_mag_1.OUT a_1432_1558# 3.64e-20
C736 a_7905_351# JK_FF_mag_3.nand3_mag_1.OUT 0.0733f
C737 a_4537_2604# CLK_div_3_mag_0.Q1 0.0102f
C738 a_5671_3745# JK_FF_mag_3.Q 9.45e-19
C739 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_3.Q 2.33e-20
C740 a_8688_3745# CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C741 a_7714_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C742 RST JK_FF_mag_5.Q 0.0193f
C743 a_8124_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C744 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C745 a_1432_1558# JK_FF_mag_5.Q 6.43e-21
C746 JK_FF_mag_5.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.00352f
C747 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 7.24e-19
C748 RST a_5424_6363# 0.00195f
C749 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.nand3_mag_1.IN1 1.4e-21
C750 JK_FF_mag_3.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.66e-20
C751 a_1996_1558# JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C752 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00306f
C753 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C754 JK_FF_mag_4.Q a_2153_4157# 0.00239f
C755 a_7751_1492# JK_FF_mag_3.nand3_mag_1.IN1 0.0697f
C756 a_5107_3745# JK_FF_mag_3.Q 6.06e-21
C757 a_3973_2604# CLK_div_3_mag_0.Q1 0.00789f
C758 a_7187_1448# JK_FF_mag_3.Q 2.79e-20
C759 a_7554_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C760 JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.Q 0.0231f
C761 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C762 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_3.Q 0.257f
C763 a_8688_3745# CLK_div_3_mag_0.JK_FF_mag_1.K 0.012f
C764 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.00352f
C765 JK_FF_mag_4.Q CLK_div_3_mag_0.JK_FF_mag_1.K 0.16f
C766 JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.05e-19
C767 JK_FF_mag_4.nand3_mag_1.OUT RST 0.284f
C768 JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_1.IN1 0.0387f
C769 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C770 RST JK_FF_mag_0.nand3_mag_1.IN1 0.258f
C771 JK_FF_mag_4.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.46e-20
C772 JK_FF_mag_5.QB a_455_3060# 0.0114f
C773 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.66f
C774 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C775 VDD a_4694_5266# 3.14e-19
C776 RST a_5264_6363# 0.00195f
C777 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.QB 0.362f
C778 a_1432_1558# JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C779 a_5261_2648# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C780 JK_FF_mag_4.nand3_mag_1.IN1 CLK 9.71e-20
C781 JK_FF_mag_0.QB a_4094_1448# 1.09e-20
C782 JK_FF_mag_5.nand3_mag_1.OUT a_2313_4157# 1.17e-20
C783 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.136f
C784 a_301_4157# JK_FF_mag_5.Q 0.0157f
C785 a_3813_2604# CLK_div_3_mag_0.Q1 0.00335f
C786 a_4543_3745# JK_FF_mag_3.Q 6.43e-21
C787 VDD a_2150_461# 3.14e-19
C788 a_6990_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C789 JK_FF_mag_2.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 7.16e-20
C790 JK_FF_mag_4.Q JK_FF_mag_5.nand3_mag_1.IN1 1.2e-19
C791 JK_FF_mag_5.nand2_mag_3.IN1 a_865_4157# 0.0036f
C792 RST a_3566_5266# 5.97e-19
C793 JK_FF_mag_2.Q JK_FF_mag_3.Q 0.16f
C794 a_8124_3745# CLK_div_3_mag_0.JK_FF_mag_1.K 2.96e-19
C795 a_2313_4157# JK_FF_mag_5.Q 0.00335f
C796 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_5.nand3_mag_1.IN1 2.62e-19
C797 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C798 VDD JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C799 a_862_417# JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C800 VDD a_5940_395# 3.14e-19
C801 a_8879_1492# JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C802 VDD JK_FF_mag_3.nand3_mag_2.OUT 0.751f
C803 VDD a_4130_5266# 3.14e-19
C804 RST a_4700_6363# 0.00173f
C805 JK_FF_mag_5.QB a_1996_1558# 2.12e-20
C806 a_4697_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C807 JK_FF_mag_3.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 4.78e-20
C808 JK_FF_mag_0.QB a_3934_1448# 1.37e-20
C809 JK_FF_mag_5.nand3_mag_1.OUT a_2153_4157# 1.5e-20
C810 VDD JK_FF_mag_3.nand2_mag_3.IN1 1.21f
C811 a_7905_351# JK_FF_mag_3.Q 0.0101f
C812 JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 3.23e-20
C813 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_2.Q 9.71e-20
C814 JK_FF_mag_2.QB JK_FF_mag_3.Q 1.61e-19
C815 a_3979_3701# JK_FF_mag_3.Q 0.00939f
C816 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C817 VDD a_7560_3745# 3.14e-19
C818 a_455_3060# JK_FF_mag_0.nand2_mag_3.IN1 2.73e-19
C819 JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand2_mag_1.IN2 0.36f
C820 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.Q1 0.0343f
C821 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C822 RST a_6830_2604# 0.00359f
C823 a_2153_4157# JK_FF_mag_5.Q 0.00789f
C824 JK_FF_mag_5.QB RST 0.0683f
C825 a_2560_1558# JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C826 JK_FF_mag_4.nand3_mag_2.OUT JK_FF_mag_4.Q 0.338f
C827 VDD JK_FF_mag_0.nand3_mag_2.OUT 0.754f
C828 JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.00627f
C829 a_3813_2604# a_3973_2604# 0.0504f
C830 RST CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00347f
C831 a_8315_1492# JK_FF_mag_3.nand2_mag_3.IN1 0.011f
C832 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C833 a_7181_351# JK_FF_mag_3.nand3_mag_2.OUT 0.0731f
C834 a_7905_351# JK_FF_mag_3.nand3_mag_1.IN1 8.64e-19
C835 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C836 JK_FF_mag_0.nand2_mag_4.IN2 a_2714_461# 0.00372f
C837 a_8688_3745# CLK_div_3_mag_0.Q0 0.069f
C838 a_4537_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C839 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_1.IN1 0.00162f
C840 JK_FF_mag_0.nand3_mag_2.OUT a_702_417# 0.0202f
C841 JK_FF_mag_5.nand3_mag_1.OUT a_1589_4157# 0.0203f
C842 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C843 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C844 a_5107_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C845 a_7181_351# JK_FF_mag_3.nand2_mag_3.IN1 1.46e-19
C846 JK_FF_mag_0.Q JK_FF_mag_2.nand3_mag_0.OUT 0.267f
C847 JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00132f
C848 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.00219f
C849 RST a_5825_2648# 0.00186f
C850 a_1589_4157# JK_FF_mag_5.Q 0.0102f
C851 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C852 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_5.nand3_mag_1.IN1 0.768f
C853 VDD a_8879_1492# 3.56e-19
C854 a_1996_1558# JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C855 JK_FF_mag_0.Q JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C856 JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1 4.49e-20
C857 a_7751_1492# JK_FF_mag_3.nand2_mag_3.IN1 1.43e-19
C858 a_6836_3701# a_6996_3701# 0.0504f
C859 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C860 a_8879_1492# JK_FF_mag_3.nand2_mag_1.IN2 0.00372f
C861 JK_FF_mag_5.nand3_mag_1.IN1 JK_FF_mag_5.Q 0.00383f
C862 a_3973_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C863 JK_FF_mag_5.nand3_mag_1.OUT a_1429_4157# 0.0733f
C864 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand2_mag_3.IN1 0.16f
C865 a_4543_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0697f
C866 JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.62e-20
C867 a_6830_2604# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C868 JK_FF_mag_4.QB RST 0.242f
C869 RST a_1586_417# 0.00196f
C870 RST JK_FF_mag_0.nand2_mag_3.IN1 0.101f
C871 VDD JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C872 JK_FF_mag_4.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.00102f
C873 VDD a_6836_3701# 2.21e-19
C874 JK_FF_mag_3.nand3_mag_0.OUT CLK_div_3_mag_0.Q0 1.59e-19
C875 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C876 JK_FF_mag_5.QB a_301_4157# 0.0811f
C877 VDD a_702_417# 0.00108f
C878 JK_FF_mag_4.nand2_mag_3.IN1 a_5264_6363# 1.46e-19
C879 a_7560_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C880 RST a_5261_2648# 8.5e-19
C881 a_3976_6363# VDD 3.14e-19
C882 a_1429_4157# JK_FF_mag_5.Q 0.0101f
C883 a_1432_1558# JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C884 VDD a_8315_1492# 3.14e-19
C885 RST CLK 0.0771f
C886 JK_FF_mag_3.nand2_mag_3.IN1 a_7187_1448# 0.00119f
C887 VDD a_3928_351# 0.00108f
C888 JK_FF_mag_4.nand2_mag_4.IN2 JK_FF_mag_3.Q 1.86e-21
C889 JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 4.64e-20
C890 RST a_5376_395# 9.98e-19
C891 JK_FF_mag_5.nand2_mag_4.IN2 JK_FF_mag_5.nand2_mag_3.IN1 0.321f
C892 JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 6.43e-20
C893 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_0.OUT 5.51e-20
C894 JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.08e-19
C895 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C896 a_4130_5266# CLK_div_3_mag_0.JK_FF_mag_1.QB 2.05e-20
C897 a_8315_1492# JK_FF_mag_3.nand2_mag_1.IN2 0.069f
C898 a_3813_2604# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C899 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_4.Q 0.413f
C900 JK_FF_mag_4.nand2_mag_3.IN1 a_3566_5266# 0.00118f
C901 JK_FF_mag_4.Q JK_FF_mag_5.nand3_mag_2.OUT 0.235f
C902 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_1.OUT 7.06e-19
C903 RST JK_FF_mag_2.nand2_mag_4.IN2 0.0236f
C904 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C905 a_3566_5266# CLK_div_3_mag_0.JK_FF_mag_1.K 3.98e-19
C906 VDD JK_FF_mag_2.nand3_mag_2.OUT 0.751f
C907 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_5.Q 0.269f
C908 JK_FF_mag_4.Q JK_FF_mag_0.QB 2.26e-19
C909 VDD a_5671_3745# 3.56e-19
C910 VDD JK_FF_mag_2.nand2_mag_3.IN1 1.37f
C911 a_5940_395# JK_FF_mag_2.Q 0.0157f
C912 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.Q 0.00335f
C913 RST a_4697_2604# 0.00147f
C914 a_5825_2648# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00372f
C915 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_2.Q 0.235f
C916 VDD a_2307_3060# 0.00536f
C917 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C918 a_3412_6363# VDD 3.14e-19
C919 VDD JK_FF_mag_5.nand3_mag_0.OUT 0.762f
C920 JK_FF_mag_4.nand3_mag_2.OUT a_5424_6363# 0.0202f
C921 VDD a_7751_1492# 3.14e-19
C922 JK_FF_mag_2.nand3_mag_2.OUT a_3928_351# 0.0202f
C923 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.Q 0.41f
C924 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_0.Q 0.00211f
C925 RST CLK_div_3_mag_0.Q1 0.277f
C926 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.655f
C927 a_5940_395# JK_FF_mag_2.QB 0.0811f
C928 JK_FF_mag_2.QB JK_FF_mag_2.nand3_mag_1.IN1 0.0382f
C929 JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 2.51e-19
C930 a_7905_351# JK_FF_mag_3.nand3_mag_2.OUT 2.88e-20
C931 a_8245_5080# CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.25e-19
C932 JK_FF_mag_0.Q JK_FF_mag_0.QB 1.95f
C933 a_3934_1448# JK_FF_mag_3.Q 3.77e-20
C934 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_2.OUT 0.121f
C935 VDD a_5107_3745# 3.14e-19
C936 JK_FF_mag_0.nand3_mag_2.OUT a_1426_417# 9.1e-19
C937 RST CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0244f
C938 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C939 a_5261_2648# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.069f
C940 RST a_4537_2604# 8.64e-19
C941 a_6996_3701# CLK_div_3_mag_0.JK_FF_mag_1.QB 1.41e-20
C942 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.QB 3e-19
C943 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C944 JK_FF_mag_4.nand3_mag_2.OUT a_5264_6363# 0.0731f
C945 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C946 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.74f
C947 JK_FF_mag_5.QB a_1589_4157# 0.00695f
C948 JK_FF_mag_0.nand2_mag_4.IN2 a_2560_1558# 4.52e-20
C949 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0215f
C950 JK_FF_mag_5.nand2_mag_1.IN2 a_455_3060# 0.00372f
C951 a_8124_3745# CLK_div_3_mag_0.or_2_mag_0.IN2 4.9e-20
C952 JK_FF_mag_5.nand3_mag_0.OUT a_2307_3060# 0.0203f
C953 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.nand3_mag_1.OUT 0.16f
C954 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB 0.884f
C955 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_5.nand3_mag_2.OUT 0.121f
C956 JK_FF_mag_5.QB JK_FF_mag_5.nand3_mag_1.IN1 0.0385f
C957 a_5222_1492# JK_FF_mag_2.nand3_mag_1.IN1 0.0059f
C958 JK_FF_mag_4.Q JK_FF_mag_4.nand3_mag_0.OUT 7.24e-19
C959 RST CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00239f
C960 VDD a_4543_3745# 3.14e-19
C961 JK_FF_mag_5.nand3_mag_1.OUT JK_FF_mag_0.QB 4.51e-20
C962 a_6836_3701# CLK_div_3_mag_0.JK_FF_mag_1.QB 1.86e-20
C963 VDD a_7027_1448# 0.00535f
C964 VDD a_1583_3060# 3.18e-19
C965 JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.11e-19
C966 VDD Vdiv96 0.152f
C967 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.Q 0.0254f
C968 JK_FF_mag_4.nand3_mag_2.OUT a_4700_6363# 9.1e-19
C969 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_8688_3745# 0.00372f
C970 RST a_2714_461# 0.00111f
C971 JK_FF_mag_5.nand3_mag_2.OUT JK_FF_mag_5.Q 0.338f
C972 a_7751_1492# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.76e-20
C973 VDD JK_FF_mag_2.Q 2.13f
C974 VDD a_1426_417# 2.21e-19
C975 JK_FF_mag_5.QB a_1429_4157# 0.00696f
C976 JK_FF_mag_4.QB JK_FF_mag_4.nand2_mag_3.IN1 0.28f
C977 RST JK_FF_mag_3.nand2_mag_4.IN2 4.47e-19
C978 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.Q1 4.33e-19
C979 JK_FF_mag_0.QB JK_FF_mag_5.Q 0.308f
C980 VDD a_4652_351# 2.21e-19
C981 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C982 JK_FF_mag_4.QB CLK_div_3_mag_0.JK_FF_mag_1.K 0.0113f
C983 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_2.Q 1.48e-20
C984 a_2147_3060# a_2307_3060# 0.0504f
C985 JK_FF_mag_5.nand3_mag_0.OUT a_2147_3060# 0.0732f
C986 a_9033_395# JK_FF_mag_3.Q 0.0157f
C987 RST a_7021_351# 0.00193f
C988 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.Q1 0.0636f
C989 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C990 CLK JK_FF_mag_4.nand2_mag_3.IN1 0.41f
C991 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C992 a_4658_1492# JK_FF_mag_2.nand3_mag_1.IN1 0.0697f
C993 a_3928_351# JK_FF_mag_2.Q 0.00335f
C994 a_3819_3701# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C995 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_7272_4844# 0.069f
C996 VDD JK_FF_mag_2.QB 0.92f
C997 CLK CLK_div_3_mag_0.JK_FF_mag_1.K 0.014f
C998 VDD a_3979_3701# 2.65e-19
C999 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_3.Q 0.235f
C1000 VDD a_1019_3060# 3.18e-19
C1001 VDD a_5786_1492# 6.86e-19
C1002 a_5671_3745# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0112f
C1003 JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.QB 5.36e-20
C1004 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q1 0.00139f
C1005 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_8124_3745# 0.069f
C1006 RST JK_FF_mag_0.nand2_mag_4.IN2 0.0293f
C1007 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00169f
C1008 a_7181_351# JK_FF_mag_2.Q 0.00212f
C1009 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_1.IN1 0.0014f
C1010 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C1011 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_5.nand3_mag_2.OUT 1.53e-20
C1012 RST JK_FF_mag_5.nand2_mag_1.IN2 0.00682f
C1013 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_5.nand3_mag_1.IN1 0.0014f
C1014 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.Q 0.338f
C1015 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C1016 JK_FF_mag_5.nand3_mag_0.OUT a_1583_3060# 0.00378f
C1017 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.Q 0.0179f
C1018 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C1019 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_1.IN1 0.0388f
C1020 a_8469_395# JK_FF_mag_3.nand2_mag_4.IN2 0.069f
C1021 JK_FF_mag_2.nand3_mag_2.OUT a_4652_351# 9.1e-19
C1022 a_7751_1492# JK_FF_mag_2.Q 6.43e-21
C1023 VDD a_5222_1492# 3.14e-19
C1024 JK_FF_mag_4.Q JK_FF_mag_3.Q 0.0449f
C1025 JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_3_mag_0.Q1 1.02e-19
C1026 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.QB 0.103f
C1027 a_8245_5080# CLK_div_3_mag_0.Q1 6.83e-19
C1028 JK_FF_mag_3.nand3_mag_0.OUT a_7714_2604# 3.1e-20
C1029 JK_FF_mag_4.nand3_mag_1.IN1 RST 0.188f
C1030 JK_FF_mag_2.QB JK_FF_mag_2.nand2_mag_3.IN1 0.28f
C1031 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q1 0.36f
C1032 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.313f
C1033 a_5786_1492# JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C1034 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C1035 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C1036 a_7027_1448# a_7187_1448# 0.0504f
C1037 a_8245_5080# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C1038 JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_2.OUT 0.103f
C1039 a_7187_1448# JK_FF_mag_2.Q 0.00939f
C1040 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.0885f
C1041 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C1042 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C1043 RST a_708_1514# 8.86e-19
C1044 CLK JK_FF_mag_4.nand3_mag_2.OUT 0.235f
C1045 JK_FF_mag_2.Q CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.14e-19
C1046 VDD a_4658_1492# 3.14e-19
C1047 JK_FF_mag_0.Q JK_FF_mag_3.Q 2.64e-20
C1048 a_4543_3745# CLK_div_3_mag_0.JK_FF_mag_1.QB 3.33e-19
C1049 JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 1.49e-19
C1050 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_5.QB 0.28f
C1051 JK_FF_mag_5.QB JK_FF_mag_5.nand3_mag_2.OUT 0.103f
C1052 JK_FF_mag_2.QB a_7187_1448# 1.26e-20
C1053 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C1054 JK_FF_mag_4.nand2_mag_4.IN2 VDD 0.391f
C1055 a_5222_1492# JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C1056 RST a_4088_351# 0.00193f
C1057 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.Q 0.00864f
C1058 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_0.OUT 0.0622f
C1059 RST JK_FF_mag_2.nand2_mag_1.IN2 0.0123f
C1060 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.198f
C1061 a_7027_1448# JK_FF_mag_2.Q 0.0101f
C1062 VDD JK_FF_mag_0.nand2_mag_1.IN2 0.409f
C1063 RST a_7745_351# 0.00172f
C1064 a_3976_6363# JK_FF_mag_4.nand2_mag_4.IN2 0.069f
C1065 JK_FF_mag_2.QB CLK_div_3_mag_0.JK_FF_mag_1.QB 2.7e-19
C1066 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00166f
C1067 a_3979_3701# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00392f
C1068 RST a_455_3060# 4.11e-19
C1069 JK_FF_mag_4.Q a_5258_5266# 2.79e-20
C1070 JK_FF_mag_4.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.49e-19
C1071 a_4652_351# JK_FF_mag_2.Q 0.0102f
C1072 JK_FF_mag_4.nand2_mag_1.IN2 JK_FF_mag_3.Q 2.25e-19
C1073 RST a_2560_1558# 9.81e-19
C1074 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C1075 CLK_div_3_mag_0.Q1 a_7272_4844# 0.01f
C1076 JK_FF_mag_2.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 7.07e-20
C1077 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C1078 JK_FF_mag_2.QB a_7027_1448# 1.62e-20
C1079 a_4658_1492# JK_FF_mag_2.nand2_mag_3.IN1 1.43e-19
C1080 JK_FF_mag_2.QB JK_FF_mag_2.Q 1.96f
C1081 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.IN2 0.124f
C1082 JK_FF_mag_2.nand3_mag_0.OUT a_4537_2604# 9.78e-20
C1083 a_5786_1492# JK_FF_mag_2.Q 0.069f
C1084 VDD a_865_4157# 3.14e-19
C1085 JK_FF_mag_2.QB a_4652_351# 0.00695f
C1086 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.Q1 0.0276f
C1087 JK_FF_mag_2.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00129f
C1088 a_3412_6363# JK_FF_mag_4.nand2_mag_4.IN2 0.00372f
C1089 VDD a_3934_1448# 0.00533f
C1090 JK_FF_mag_5.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.0945f
C1091 RST a_1996_1558# 0.00163f
C1092 JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 1.47e-19
C1093 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C1094 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_3.IN1 0.28f
C1095 a_7560_3745# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C1096 JK_FF_mag_0.QB a_1586_417# 0.00696f
C1097 JK_FF_mag_2.QB a_5786_1492# 0.0114f
C1098 a_4094_1448# JK_FF_mag_2.nand2_mag_3.IN1 0.00119f
C1099 JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00109f
C1100 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.404f
C1101 a_5222_1492# JK_FF_mag_2.Q 5.39e-21
C1102 a_2150_461# JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C1103 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand2_mag_3.IN1 0.233f
C1104 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_3.Q 7.13e-20
C1105 JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 2.19e-20
C1106 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C1107 JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 0.00216f
C1108 JK_FF_mag_5.nand2_mag_1.IN2 JK_FF_mag_5.nand3_mag_1.IN1 0.109f
C1109 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C1110 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.Q0 0.0635f
C1111 RST a_1432_1558# 0.0013f
C1112 a_6996_3701# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C1113 JK_FF_mag_2.QB a_5222_1492# 2.96e-19
C1114 JK_FF_mag_3.Q CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.29f
C1115 a_7745_351# JK_FF_mag_3.QB 0.00695f
C1116 JK_FF_mag_0.Q a_2150_461# 0.00859f
C1117 VDD a_9033_395# 3.14e-19
C1118 RST a_4812_351# 0.00189f
C1119 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C1120 JK_FF_mag_0.Q JK_FF_mag_2.nand3_mag_1.IN1 9.71e-20
C1121 a_5671_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00372f
C1122 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C1123 JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_0.OUT 0.343f
C1124 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.806f
C1125 a_6836_3701# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C1126 JK_FF_mag_2.QB a_4658_1492# 3.33e-19
C1127 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C1128 CLK JK_FF_mag_4.nand3_mag_0.OUT 0.267f
C1129 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.279f
C1130 a_4094_1448# JK_FF_mag_2.Q 2.79e-20
C1131 a_6830_2604# JK_FF_mag_3.Q 0.00749f
C1132 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.nand2_mag_3.IN1 0.088f
C1133 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.Q 0.338f
C1134 a_4540_6363# JK_FF_mag_4.Q 0.0101f
C1135 JK_FF_mag_5.QB JK_FF_mag_3.Q 2.73e-21
C1136 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0592f
C1137 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.or_2_mag_0.IN2 0.0138f
C1138 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand3_mag_2.OUT 0.00167f
C1139 JK_FF_mag_3.Q CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0983f
C1140 JK_FF_mag_2.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 2.34e-19
C1141 a_5107_3745# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.069f
C1142 JK_FF_mag_5.nand2_mag_4.IN2 VDD 0.391f
C1143 VDD JK_FF_mag_2.nand3_mag_1.OUT 0.995f
C1144 JK_FF_mag_4.nand2_mag_1.IN2 a_4130_5266# 0.069f
C1145 VDD a_8688_3745# 3.56e-19
C1146 JK_FF_mag_4.Q VDD 2.21f
C1147 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.or_2_mag_0.IN2 5.32e-19
C1148 JK_FF_mag_2.QB a_4094_1448# 0.00392f
C1149 RST JK_FF_mag_3.QB 0.116f
C1150 a_5258_5266# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.13e-20
C1151 VDD JK_FF_mag_0.nand3_mag_1.OUT 0.999f
C1152 a_6990_2604# a_6830_2604# 0.0504f
C1153 JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 8.81e-20
C1154 JK_FF_mag_0.QB a_2714_461# 0.0811f
C1155 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C1156 a_708_1514# JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C1157 JK_FF_mag_2.nand3_mag_1.OUT a_3928_351# 1.17e-20
C1158 a_3976_6363# JK_FF_mag_4.Q 0.00859f
C1159 JK_FF_mag_4.nand3_mag_1.OUT a_4694_5266# 0.0202f
C1160 JK_FF_mag_4.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.51e-19
C1161 a_702_417# JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C1162 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C1163 a_9033_395# VSS 0.0765f
C1164 a_8469_395# VSS 0.0767f
C1165 a_7905_351# VSS 0.0522f
C1166 a_7745_351# VSS 0.106f
C1167 a_7181_351# VSS 0.0522f
C1168 a_7021_351# VSS 0.106f
C1169 a_5940_395# VSS 0.0765f
C1170 a_5376_395# VSS 0.0767f
C1171 a_4812_351# VSS 0.0522f
C1172 a_4652_351# VSS 0.106f
C1173 a_4088_351# VSS 0.0522f
C1174 a_3928_351# VSS 0.106f
C1175 a_2714_461# VSS 0.0675f
C1176 a_2150_461# VSS 0.0676f
C1177 a_1586_417# VSS 0.0343f
C1178 a_1426_417# VSS 0.0881f
C1179 a_862_417# VSS 0.0343f
C1180 a_702_417# VSS 0.0881f
C1181 JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.428f
C1182 JK_FF_mag_3.nand3_mag_2.OUT VSS 0.595f
C1183 JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.428f
C1184 JK_FF_mag_2.nand3_mag_2.OUT VSS 0.595f
C1185 JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C1186 JK_FF_mag_0.nand3_mag_2.OUT VSS 0.537f
C1187 a_8879_1492# VSS 0.0676f
C1188 a_8315_1492# VSS 0.0676f
C1189 a_7751_1492# VSS 0.0676f
C1190 a_7187_1448# VSS 0.0343f
C1191 a_7027_1448# VSS 0.0881f
C1192 a_5786_1492# VSS 0.0676f
C1193 a_5222_1492# VSS 0.0676f
C1194 a_4658_1492# VSS 0.0677f
C1195 a_4094_1448# VSS 0.0349f
C1196 a_3934_1448# VSS 0.0891f
C1197 a_2560_1558# VSS 0.0685f
C1198 a_1996_1558# VSS 0.068f
C1199 a_1432_1558# VSS 0.0676f
C1200 a_868_1514# VSS 0.0343f
C1201 a_708_1514# VSS 0.0881f
C1202 JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.414f
C1203 JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.711f
C1204 JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.726f
C1205 JK_FF_mag_3.nand3_mag_1.OUT VSS 0.865f
C1206 JK_FF_mag_3.nand3_mag_0.OUT VSS 0.507f
C1207 JK_FF_mag_3.QB VSS 0.906f
C1208 JK_FF_mag_2.Q VSS 2.24f
C1209 JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.414f
C1210 JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.774f
C1211 JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.727f
C1212 JK_FF_mag_2.nand3_mag_1.OUT VSS 0.866f
C1213 JK_FF_mag_2.nand3_mag_0.OUT VSS 0.514f
C1214 JK_FF_mag_2.QB VSS 0.907f
C1215 JK_FF_mag_0.Q VSS 2.39f
C1216 JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.416f
C1217 JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.742f
C1218 JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.723f
C1219 JK_FF_mag_0.nand3_mag_1.OUT VSS 0.805f
C1220 JK_FF_mag_0.nand3_mag_0.OUT VSS 0.505f
C1221 JK_FF_mag_0.QB VSS 0.894f
C1222 a_8842_2648# VSS 0.0675f
C1223 a_8278_2648# VSS 0.0676f
C1224 a_7714_2604# VSS 0.0343f
C1225 a_7554_2604# VSS 0.0881f
C1226 a_6990_2604# VSS 0.0343f
C1227 a_6830_2604# VSS 0.0881f
C1228 a_5825_2648# VSS 0.0675f
C1229 a_5261_2648# VSS 0.0676f
C1230 a_4697_2604# VSS 0.0344f
C1231 a_4537_2604# VSS 0.0883f
C1232 a_3973_2604# VSS 0.0352f
C1233 a_3813_2604# VSS 0.0893f
C1234 a_2307_3060# VSS 0.089f
C1235 a_2147_3060# VSS 0.0348f
C1236 a_1583_3060# VSS 0.0676f
C1237 a_1019_3060# VSS 0.0676f
C1238 a_455_3060# VSS 0.0676f
C1239 JK_FF_mag_5.nand3_mag_0.OUT VSS 0.509f
C1240 JK_FF_mag_5.nand2_mag_1.IN2 VSS 0.41f
C1241 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.412f
C1242 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.537f
C1243 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.413f
C1244 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.524f
C1245 a_8688_3745# VSS 0.0676f
C1246 a_8124_3745# VSS 0.0676f
C1247 a_7560_3745# VSS 0.0676f
C1248 a_6996_3701# VSS 0.0343f
C1249 a_6836_3701# VSS 0.0881f
C1250 a_5671_3745# VSS 0.0676f
C1251 a_5107_3745# VSS 0.0676f
C1252 a_4543_3745# VSS 0.0676f
C1253 a_3979_3701# VSS 0.0343f
C1254 a_3819_3701# VSS 0.0881f
C1255 a_2313_4157# VSS 0.0949f
C1256 a_2153_4157# VSS 0.041f
C1257 a_1589_4157# VSS 0.0948f
C1258 a_1429_4157# VSS 0.041f
C1259 a_865_4157# VSS 0.0715f
C1260 a_301_4157# VSS 0.0714f
C1261 JK_FF_mag_5.QB VSS 0.894f
C1262 JK_FF_mag_5.nand3_mag_1.OUT VSS 0.826f
C1263 JK_FF_mag_5.nand2_mag_3.IN1 VSS 0.746f
C1264 JK_FF_mag_5.nand2_mag_4.IN2 VSS 0.421f
C1265 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1266 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.687f
C1267 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.721f
C1268 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.806f
C1269 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1270 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.41f
C1271 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.699f
C1272 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.717f
C1273 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.802f
C1274 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.505f
C1275 CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.852f
C1276 CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.28f
C1277 JK_FF_mag_5.Q VSS 3.16f
C1278 JK_FF_mag_5.nand3_mag_2.OUT VSS 0.56f
C1279 JK_FF_mag_5.nand3_mag_1.IN1 VSS 0.722f
C1280 a_7272_4844# VSS 0.0676f
C1281 Vdiv96 VSS 0.247f
C1282 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C1283 a_8245_5080# VSS 0.0247f
C1284 CLK_div_3_mag_0.Q0 VSS 1.73f
C1285 CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.418f
C1286 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C1287 CLK_div_3_mag_0.Q1 VSS 1.73f
C1288 JK_FF_mag_3.Q VSS 4.14f
C1289 a_5418_5266# VSS 0.0881f
C1290 a_5258_5266# VSS 0.0343f
C1291 a_4694_5266# VSS 0.0676f
C1292 a_4130_5266# VSS 0.0676f
C1293 a_3566_5266# VSS 0.0676f
C1294 JK_FF_mag_4.nand3_mag_0.OUT VSS 0.505f
C1295 JK_FF_mag_4.nand2_mag_1.IN2 VSS 0.41f
C1296 a_5424_6363# VSS 0.0961f
C1297 a_5264_6363# VSS 0.0422f
C1298 a_4700_6363# VSS 0.096f
C1299 a_4540_6363# VSS 0.0422f
C1300 a_3976_6363# VSS 0.0721f
C1301 a_3412_6363# VSS 0.072f
C1302 JK_FF_mag_4.QB VSS 0.899f
C1303 JK_FF_mag_4.nand3_mag_1.OUT VSS 0.83f
C1304 JK_FF_mag_4.nand2_mag_3.IN1 VSS 0.706f
C1305 JK_FF_mag_4.nand2_mag_4.IN2 VSS 0.423f
C1306 CLK VSS 1.01f
C1307 JK_FF_mag_4.Q VSS 3.62f
C1308 JK_FF_mag_4.nand3_mag_2.OUT VSS 0.564f
C1309 RST VSS 6.49f
C1310 JK_FF_mag_4.nand3_mag_1.IN1 VSS 0.722f
C1311 VDD VSS 0.101p
C1312 JK_FF_mag_5.Q.n0 VSS 0.25f
C1313 JK_FF_mag_5.Q.t2 VSS 0.0172f
C1314 JK_FF_mag_5.Q.t0 VSS 0.0142f
C1315 JK_FF_mag_5.Q.n1 VSS 0.0142f
C1316 JK_FF_mag_5.Q.n2 VSS 0.0341f
C1317 JK_FF_mag_5.Q.t5 VSS 0.0208f
C1318 JK_FF_mag_5.Q.t7 VSS 0.0316f
C1319 JK_FF_mag_5.Q.n3 VSS 0.0559f
C1320 JK_FF_mag_5.Q.t3 VSS 0.0208f
C1321 JK_FF_mag_5.Q.t6 VSS 0.0316f
C1322 JK_FF_mag_5.Q.n4 VSS 0.0559f
C1323 JK_FF_mag_5.Q.t8 VSS 0.00668f
C1324 JK_FF_mag_5.Q.t4 VSS 0.0261f
C1325 JK_FF_mag_5.Q.n5 VSS 0.0433f
C1326 JK_FF_mag_5.Q.t10 VSS 0.0316f
C1327 JK_FF_mag_5.Q.t9 VSS 0.0208f
C1328 JK_FF_mag_5.Q.n6 VSS 0.0562f
C1329 JK_FF_mag_5.Q.t12 VSS 0.0227f
C1330 JK_FF_mag_5.Q.t11 VSS 0.0182f
C1331 JK_FF_mag_5.Q.n7 VSS 0.0527f
C1332 JK_FF_mag_5.Q.n8 VSS 0.419f
C1333 JK_FF_mag_5.Q.n9 VSS 0.295f
C1334 JK_FF_mag_4.Q.n0 VSS 0.225f
C1335 JK_FF_mag_4.Q.t1 VSS 0.0155f
C1336 JK_FF_mag_4.Q.t0 VSS 0.0128f
C1337 JK_FF_mag_4.Q.n1 VSS 0.0128f
C1338 JK_FF_mag_4.Q.n2 VSS 0.0307f
C1339 JK_FF_mag_4.Q.t6 VSS 0.0285f
C1340 JK_FF_mag_4.Q.t4 VSS 0.0187f
C1341 JK_FF_mag_4.Q.n3 VSS 0.0505f
C1342 JK_FF_mag_4.Q.t5 VSS 0.0204f
C1343 JK_FF_mag_4.Q.t3 VSS 0.0163f
C1344 JK_FF_mag_4.Q.n4 VSS 0.0474f
C1345 JK_FF_mag_4.Q.n5 VSS 0.378f
C1346 JK_FF_mag_4.Q.t10 VSS 0.0285f
C1347 JK_FF_mag_4.Q.t9 VSS 0.0187f
C1348 JK_FF_mag_4.Q.n6 VSS 0.0503f
C1349 JK_FF_mag_4.Q.t12 VSS 0.0285f
C1350 JK_FF_mag_4.Q.t11 VSS 0.0187f
C1351 JK_FF_mag_4.Q.n7 VSS 0.0503f
C1352 JK_FF_mag_4.Q.t7 VSS 0.0235f
C1353 JK_FF_mag_4.Q.t8 VSS 0.00607f
C1354 JK_FF_mag_4.Q.n8 VSS 0.039f
C1355 JK_FF_mag_4.Q.n9 VSS 0.39f
C1356 RST.t2 VSS 0.00813f
C1357 RST.t3 VSS 0.0123f
C1358 RST.n0 VSS 0.0218f
C1359 RST.n1 VSS 0.00383f
C1360 RST.n2 VSS 0.00281f
C1361 RST.n3 VSS 0.00131f
C1362 RST.n4 VSS 0.00102f
C1363 RST.n5 VSS 0.0812f
C1364 RST.n6 VSS 0.00366f
C1365 RST.n7 VSS 0.00189f
C1366 RST.t13 VSS 0.0125f
C1367 RST.t12 VSS 0.00793f
C1368 RST.n8 VSS 0.0219f
C1369 RST.n9 VSS 0.00281f
C1370 RST.n10 VSS 0.001f
C1371 RST.n11 VSS 0.0458f
C1372 RST.n12 VSS 0.00356f
C1373 RST.n13 VSS 0.00187f
C1374 RST.t5 VSS 0.00813f
C1375 RST.t7 VSS 0.0123f
C1376 RST.n14 VSS 0.0218f
C1377 RST.n15 VSS 0.00289f
C1378 RST.n16 VSS 0.001f
C1379 RST.n17 VSS 0.00154f
C1380 RST.n18 VSS 0.00572f
C1381 RST.n19 VSS 0.107f
C1382 RST.t9 VSS 0.0123f
C1383 RST.t8 VSS 0.00813f
C1384 RST.n20 VSS 0.0219f
C1385 RST.n21 VSS 0.126f
C1386 RST.n22 VSS 0.195f
C1387 RST.n23 VSS 0.00135f
C1388 RST.t4 VSS 0.00813f
C1389 RST.t6 VSS 0.0123f
C1390 RST.n24 VSS 0.0218f
C1391 RST.n25 VSS 0.00362f
C1392 RST.n26 VSS 0.001f
C1393 RST.n27 VSS 0.00281f
C1394 RST.n28 VSS 0.00379f
C1395 RST.n29 VSS 0.00159f
C1396 RST.n30 VSS 0.00386f
C1397 RST.n31 VSS 0.214f
C1398 RST.n32 VSS 0.205f
C1399 RST.n33 VSS 0.00385f
C1400 RST.n34 VSS 0.00182f
C1401 RST.t10 VSS 0.00813f
C1402 RST.t11 VSS 0.0123f
C1403 RST.n35 VSS 0.0218f
C1404 RST.n36 VSS 0.00289f
C1405 RST.n37 VSS 0.00108f
C1406 RST.n38 VSS 0.00142f
C1407 RST.n39 VSS 0.00519f
C1408 RST.n40 VSS 2.96e-19
C1409 RST.n41 VSS 0.00211f
C1410 RST.n42 VSS 0.00205f
C1411 RST.n43 VSS 0.099f
C1412 RST.n44 VSS 0.33f
C1413 RST.n45 VSS 0.583f
C1414 RST.n46 VSS 0.00307f
C1415 RST.t1 VSS 0.0123f
C1416 RST.t0 VSS 0.00813f
C1417 RST.n47 VSS 0.0218f
C1418 RST.n48 VSS 0.00285f
C1419 RST.n49 VSS 0.00189f
C1420 RST.n50 VSS 0.001f
C1421 RST.n51 VSS 0.00133f
C1422 RST.n52 VSS 0.00551f
C1423 RST.n53 VSS 0.32f
C1424 RST.n54 VSS 0.00351f
C1425 RST.n55 VSS 0.143f
C1426 RST.n56 VSS 0.151f
C1427 RST.n57 VSS 0.0754f
C1428 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.15f
C1429 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.208f
C1430 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0724f
C1431 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0562f
C1432 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.143f
C1433 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.0449f
C1434 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS 0.0563f
C1435 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.145f
C1436 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.079f
C1437 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0503f
C1438 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.14f
C1439 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 1.2f
C1440 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VSS 0.0351f
C1441 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 0.0351f
C1442 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.0828f
C1443 VDD.t68 VSS 0.08f
C1444 VDD.t221 VSS 0.00595f
C1445 VDD.t9 VSS 0.00245f
C1446 VDD.n0 VSS 0.00245f
C1447 VDD.n1 VSS 0.00534f
C1448 VDD.t278 VSS 0.0319f
C1449 VDD.t363 VSS 0.0323f
C1450 VDD.t364 VSS 0.00595f
C1451 VDD.n2 VSS 0.00595f
C1452 VDD.t157 VSS 0.0323f
C1453 VDD.t299 VSS 0.00245f
C1454 VDD.n3 VSS 0.00245f
C1455 VDD.n4 VSS 0.00534f
C1456 VDD.n5 VSS 0.00595f
C1457 VDD.t255 VSS 0.00595f
C1458 VDD.n6 VSS 0.0235f
C1459 VDD.t10 VSS 0.08f
C1460 VDD.n7 VSS 0.00629f
C1461 VDD.n8 VSS 0.00595f
C1462 VDD.t47 VSS 0.0775f
C1463 VDD.n9 VSS 0.0369f
C1464 VDD.t238 VSS 0.00595f
C1465 VDD.n10 VSS 0.00595f
C1466 VDD.t237 VSS 0.0718f
C1467 VDD.t127 VSS 0.0786f
C1468 VDD.n11 VSS 0.0369f
C1469 VDD.t282 VSS 0.00595f
C1470 VDD.t360 VSS 0.00245f
C1471 VDD.n12 VSS 0.00245f
C1472 VDD.n13 VSS 0.00534f
C1473 VDD.t281 VSS 0.0718f
C1474 VDD.t359 VSS 0.0876f
C1475 VDD.t165 VSS 0.0407f
C1476 VDD.n14 VSS 0.0369f
C1477 VDD.t323 VSS 0.00595f
C1478 VDD.t46 VSS 0.00245f
C1479 VDD.n15 VSS 0.00245f
C1480 VDD.n16 VSS 0.00534f
C1481 VDD.t322 VSS 0.0718f
C1482 VDD.t45 VSS 0.0876f
C1483 VDD.t76 VSS 0.0407f
C1484 VDD.t106 VSS 0.0716f
C1485 VDD.n17 VSS 0.0369f
C1486 VDD.t107 VSS 0.00556f
C1487 VDD.t327 VSS 0.00245f
C1488 VDD.n18 VSS 0.00245f
C1489 VDD.n19 VSS 0.00534f
C1490 VDD.n20 VSS 0.0319f
C1491 VDD.t83 VSS 0.00595f
C1492 VDD.t21 VSS 0.0423f
C1493 VDD.n21 VSS 0.00595f
C1494 VDD.t22 VSS 0.00595f
C1495 VDD.n22 VSS 0.00595f
C1496 VDD.n23 VSS 0.0295f
C1497 VDD.t328 VSS 0.0625f
C1498 VDD.n24 VSS 0.00595f
C1499 VDD.n25 VSS 0.00595f
C1500 VDD.t207 VSS 0.0775f
C1501 VDD.n26 VSS 0.0369f
C1502 VDD.t171 VSS 0.00595f
C1503 VDD.n27 VSS 0.00595f
C1504 VDD.t170 VSS 0.0718f
C1505 VDD.t353 VSS 0.0786f
C1506 VDD.n28 VSS 0.0369f
C1507 VDD.t339 VSS 0.00595f
C1508 VDD.t24 VSS 0.00245f
C1509 VDD.n29 VSS 0.00245f
C1510 VDD.n30 VSS 0.00534f
C1511 VDD.t338 VSS 0.0718f
C1512 VDD.t23 VSS 0.0876f
C1513 VDD.t13 VSS 0.0407f
C1514 VDD.n31 VSS 0.0369f
C1515 VDD.t223 VSS 0.00595f
C1516 VDD.t200 VSS 0.00245f
C1517 VDD.n32 VSS 0.00245f
C1518 VDD.n33 VSS 0.00534f
C1519 VDD.t222 VSS 0.0718f
C1520 VDD.t199 VSS 0.0876f
C1521 VDD.t285 VSS 0.0407f
C1522 VDD.t103 VSS 0.0716f
C1523 VDD.n34 VSS 0.0369f
C1524 VDD.t104 VSS 0.00595f
C1525 VDD.t81 VSS 0.00511f
C1526 VDD.t368 VSS 0.00387f
C1527 VDD.n35 VSS 0.01f
C1528 VDD.t102 VSS 0.00511f
C1529 VDD.t376 VSS 0.00387f
C1530 VDD.n36 VSS 0.01f
C1531 VDD.n37 VSS 0.00835f
C1532 VDD.n38 VSS 0.0437f
C1533 VDD.n39 VSS 0.0277f
C1534 VDD.n40 VSS 0.0185f
C1535 VDD.n41 VSS 0.0339f
C1536 VDD.n42 VSS 0.0348f
C1537 VDD.n43 VSS 0.0185f
C1538 VDD.n44 VSS 0.0339f
C1539 VDD.n45 VSS 0.0347f
C1540 VDD.n46 VSS 0.0206f
C1541 VDD.n47 VSS 0.0295f
C1542 VDD.n48 VSS 0.0274f
C1543 VDD.n49 VSS 0.0206f
C1544 VDD.n50 VSS 0.0515f
C1545 VDD.t198 VSS 0.00593f
C1546 VDD.t114 VSS 0.00595f
C1547 VDD.n51 VSS 0.0316f
C1548 VDD.t197 VSS 0.0525f
C1549 VDD.t204 VSS 0.0407f
C1550 VDD.t269 VSS 0.00245f
C1551 VDD.n52 VSS 0.00245f
C1552 VDD.n53 VSS 0.00534f
C1553 VDD.t217 VSS 0.00595f
C1554 VDD.n54 VSS 0.00595f
C1555 VDD.n55 VSS 0.0295f
C1556 VDD.t191 VSS 0.0786f
C1557 VDD.n56 VSS 0.00595f
C1558 VDD.t143 VSS 0.00595f
C1559 VDD.n57 VSS 0.00595f
C1560 VDD.n58 VSS 0.00595f
C1561 VDD.t56 VSS 0.0775f
C1562 VDD.n59 VSS 0.0369f
C1563 VDD.t267 VSS 0.00595f
C1564 VDD.n60 VSS 0.00595f
C1565 VDD.t266 VSS 0.0718f
C1566 VDD.t188 VSS 0.0786f
C1567 VDD.n61 VSS 0.0369f
C1568 VDD.t20 VSS 0.00595f
C1569 VDD.t152 VSS 0.00245f
C1570 VDD.n62 VSS 0.00245f
C1571 VDD.n63 VSS 0.00534f
C1572 VDD.t19 VSS 0.0718f
C1573 VDD.t151 VSS 0.0876f
C1574 VDD.t121 VSS 0.0407f
C1575 VDD.n64 VSS 0.0369f
C1576 VDD.t263 VSS 0.00595f
C1577 VDD.t65 VSS 0.00245f
C1578 VDD.n65 VSS 0.00245f
C1579 VDD.n66 VSS 0.00534f
C1580 VDD.t262 VSS 0.0718f
C1581 VDD.t64 VSS 0.0876f
C1582 VDD.t201 VSS 0.0407f
C1583 VDD.t119 VSS 0.0716f
C1584 VDD.n67 VSS 0.0369f
C1585 VDD.t120 VSS 0.00595f
C1586 VDD.t112 VSS 0.00511f
C1587 VDD.t372 VSS 0.00387f
C1588 VDD.n68 VSS 0.01f
C1589 VDD.t118 VSS 0.00511f
C1590 VDD.t369 VSS 0.00387f
C1591 VDD.n69 VSS 0.01f
C1592 VDD.n70 VSS 0.00762f
C1593 VDD.n71 VSS 0.0415f
C1594 VDD.n72 VSS 0.0277f
C1595 VDD.n73 VSS 0.0185f
C1596 VDD.n74 VSS 0.0339f
C1597 VDD.n75 VSS 0.0348f
C1598 VDD.n76 VSS 0.0185f
C1599 VDD.n77 VSS 0.0339f
C1600 VDD.n78 VSS 0.0347f
C1601 VDD.n79 VSS 0.0206f
C1602 VDD.n80 VSS 0.0295f
C1603 VDD.n81 VSS 0.0274f
C1604 VDD.n82 VSS 0.0206f
C1605 VDD.n83 VSS 0.0561f
C1606 VDD.n84 VSS 0.0638f
C1607 VDD.t270 VSS 0.0775f
C1608 VDD.t142 VSS 0.0718f
C1609 VDD.n85 VSS 0.0369f
C1610 VDD.n86 VSS 0.0206f
C1611 VDD.n87 VSS 0.0274f
C1612 VDD.n88 VSS 0.0295f
C1613 VDD.t154 VSS 0.00595f
C1614 VDD.n89 VSS 0.0274f
C1615 VDD.n90 VSS 0.0206f
C1616 VDD.n91 VSS 0.0369f
C1617 VDD.t153 VSS 0.0718f
C1618 VDD.t16 VSS 0.0786f
C1619 VDD.t268 VSS 0.0876f
C1620 VDD.t216 VSS 0.0718f
C1621 VDD.n92 VSS 0.0369f
C1622 VDD.n93 VSS 0.0206f
C1623 VDD.n94 VSS 0.026f
C1624 VDD.n95 VSS 0.0243f
C1625 VDD.n96 VSS 0.0185f
C1626 VDD.n97 VSS 0.0369f
C1627 VDD.t113 VSS 0.0407f
C1628 VDD.n98 VSS 0.0553f
C1629 VDD.n99 VSS 0.0292f
C1630 VDD.n100 VSS 0.0494f
C1631 VDD.n101 VSS 0.0288f
C1632 VDD.t297 VSS 0.00595f
C1633 VDD.n102 VSS 0.0274f
C1634 VDD.n103 VSS 0.0206f
C1635 VDD.n104 VSS 0.0319f
C1636 VDD.t296 VSS 0.0571f
C1637 VDD.t356 VSS 0.0625f
C1638 VDD.n105 VSS 0.0319f
C1639 VDD.n106 VSS 0.0206f
C1640 VDD.n107 VSS 0.0274f
C1641 VDD.n108 VSS 0.0295f
C1642 VDD.t184 VSS 0.00595f
C1643 VDD.n109 VSS 0.026f
C1644 VDD.n110 VSS 0.0206f
C1645 VDD.t293 VSS 0.0324f
C1646 VDD.t326 VSS 0.0697f
C1647 VDD.t183 VSS 0.0571f
C1648 VDD.n111 VSS 0.0319f
C1649 VDD.t335 VSS 0.0274f
C1650 VDD.n112 VSS 0.165f
C1651 VDD.t82 VSS 0.0324f
C1652 VDD.n113 VSS 0.0912f
C1653 VDD.t283 VSS 0.0656f
C1654 VDD.t284 VSS 0.00593f
C1655 VDD.n114 VSS 0.00593f
C1656 VDD.t300 VSS 0.03f
C1657 VDD.n115 VSS 0.00591f
C1658 VDD.t174 VSS 0.0786f
C1659 VDD.n116 VSS 0.0618f
C1660 VDD.n117 VSS 0.00592f
C1661 VDD.t53 VSS 0.00592f
C1662 VDD.t52 VSS 0.0469f
C1663 VDD.t99 VSS 0.0472f
C1664 VDD.n118 VSS 0.0618f
C1665 VDD.n119 VSS 0.00591f
C1666 VDD.t325 VSS 0.00245f
C1667 VDD.n120 VSS 0.00245f
C1668 VDD.n121 VSS 0.00531f
C1669 VDD.t324 VSS 0.0783f
C1670 VDD.t28 VSS 0.0497f
C1671 VDD.t314 VSS 0.0317f
C1672 VDD.n122 VSS 0.059f
C1673 VDD.t39 VSS 0.00592f
C1674 VDD.n123 VSS 0.00592f
C1675 VDD.t38 VSS 0.0966f
C1676 VDD.t241 VSS 0.0969f
C1677 VDD.n124 VSS 0.059f
C1678 VDD.n125 VSS 0.00591f
C1679 VDD.t150 VSS 0.00592f
C1680 VDD.t3 VSS 0.0314f
C1681 VDD.t149 VSS 0.0317f
C1682 VDD.n126 VSS 0.059f
C1683 VDD.t32 VSS 0.00592f
C1684 VDD.n127 VSS 0.00592f
C1685 VDD.t31 VSS 0.0966f
C1686 VDD.t309 VSS 0.0969f
C1687 VDD.n128 VSS 0.059f
C1688 VDD.t173 VSS 0.00245f
C1689 VDD.n129 VSS 0.00245f
C1690 VDD.n130 VSS 0.0053f
C1691 VDD.t341 VSS 0.00592f
C1692 VDD.t172 VSS 0.0314f
C1693 VDD.t340 VSS 0.0497f
C1694 VDD.t130 VSS 0.0786f
C1695 VDD.n131 VSS 0.0618f
C1696 VDD.n132 VSS 0.00592f
C1697 VDD.t97 VSS 0.00592f
C1698 VDD.t96 VSS 0.0469f
C1699 VDD.t226 VSS 0.0472f
C1700 VDD.n133 VSS 0.0618f
C1701 VDD.t313 VSS 0.00592f
C1702 VDD.t312 VSS 0.0783f
C1703 VDD.t133 VSS 0.0301f
C1704 VDD.t134 VSS 0.00592f
C1705 VDD.t213 VSS 0.00595f
C1706 VDD.t146 VSS 0.0719f
C1707 VDD.n134 VSS 0.00595f
C1708 VDD.t211 VSS 0.00245f
C1709 VDD.n135 VSS 0.00245f
C1710 VDD.n136 VSS 0.00534f
C1711 VDD.n137 VSS 0.00595f
C1712 VDD.n138 VSS 0.0348f
C1713 VDD.t109 VSS 0.0717f
C1714 VDD.n139 VSS 0.00595f
C1715 VDD.t373 VSS 0.00387f
C1716 VDD.t108 VSS 0.00511f
C1717 VDD.n140 VSS 0.01f
C1718 VDD.n141 VSS 0.00741f
C1719 VDD.t377 VSS 0.00387f
C1720 VDD.t98 VSS 0.00511f
C1721 VDD.n142 VSS 0.01f
C1722 VDD.n143 VSS 0.0045f
C1723 VDD.n144 VSS 0.0036f
C1724 VDD.n145 VSS 0.0365f
C1725 VDD.n146 VSS 0.0278f
C1726 VDD.t265 VSS 0.00245f
C1727 VDD.n147 VSS 0.00245f
C1728 VDD.n148 VSS 0.00534f
C1729 VDD.n149 VSS 0.0339f
C1730 VDD.n150 VSS 0.0184f
C1731 VDD.n151 VSS 0.0369f
C1732 VDD.t264 VSS 0.0405f
C1733 VDD.t194 VSS 0.0876f
C1734 VDD.t244 VSS 0.0719f
C1735 VDD.t306 VSS 0.0876f
C1736 VDD.t210 VSS 0.0405f
C1737 VDD.n152 VSS 0.0369f
C1738 VDD.n153 VSS 0.0184f
C1739 VDD.n154 VSS 0.0339f
C1740 VDD.n155 VSS 0.0347f
C1741 VDD.t343 VSS 0.00595f
C1742 VDD.n156 VSS 0.00595f
C1743 VDD.n157 VSS 0.0274f
C1744 VDD.n158 VSS 0.0295f
C1745 VDD.n159 VSS 0.0206f
C1746 VDD.n160 VSS 0.0369f
C1747 VDD.t342 VSS 0.0785f
C1748 VDD.t251 VSS 0.0719f
C1749 VDD.t212 VSS 0.0773f
C1750 VDD.n161 VSS 0.0369f
C1751 VDD.n162 VSS 0.0206f
C1752 VDD.n163 VSS 0.0521f
C1753 VDD.n164 VSS 0.0659f
C1754 VDD.n165 VSS 0.0345f
C1755 VDD.n166 VSS 0.0303f
C1756 VDD.n167 VSS 0.023f
C1757 VDD.n168 VSS 0.0233f
C1758 VDD.n169 VSS 0.0193f
C1759 VDD.n170 VSS 0.0275f
C1760 VDD.n171 VSS 0.0249f
C1761 VDD.n172 VSS 0.0289f
C1762 VDD.n173 VSS 0.0303f
C1763 VDD.n174 VSS 0.0322f
C1764 VDD.n175 VSS 0.0133f
C1765 VDD.n176 VSS 0.0277f
C1766 VDD.n177 VSS 0.0276f
C1767 VDD.n178 VSS 0.0133f
C1768 VDD.n179 VSS 0.0322f
C1769 VDD.n180 VSS 0.0304f
C1770 VDD.n181 VSS 0.0288f
C1771 VDD.n182 VSS 0.0249f
C1772 VDD.n183 VSS 0.0275f
C1773 VDD.n184 VSS 0.0192f
C1774 VDD.n185 VSS 0.0233f
C1775 VDD.n186 VSS 0.0231f
C1776 VDD.n187 VSS 0.0302f
C1777 VDD.n188 VSS 0.0346f
C1778 VDD.n189 VSS 0.0364f
C1779 VDD.n190 VSS 0.00595f
C1780 VDD.t290 VSS 0.0775f
C1781 VDD.n191 VSS 0.0369f
C1782 VDD.t230 VSS 0.00595f
C1783 VDD.n192 VSS 0.00595f
C1784 VDD.t229 VSS 0.0718f
C1785 VDD.t25 VSS 0.0786f
C1786 VDD.n193 VSS 0.0369f
C1787 VDD.t7 VSS 0.00595f
C1788 VDD.t37 VSS 0.00245f
C1789 VDD.n194 VSS 0.00245f
C1790 VDD.n195 VSS 0.00534f
C1791 VDD.t6 VSS 0.0718f
C1792 VDD.t36 VSS 0.0876f
C1793 VDD.t347 VSS 0.0407f
C1794 VDD.n196 VSS 0.0369f
C1795 VDD.t51 VSS 0.00595f
C1796 VDD.t289 VSS 0.00245f
C1797 VDD.n197 VSS 0.00245f
C1798 VDD.n198 VSS 0.00534f
C1799 VDD.t50 VSS 0.0718f
C1800 VDD.t288 VSS 0.0876f
C1801 VDD.t317 VSS 0.0407f
C1802 VDD.t89 VSS 0.0716f
C1803 VDD.n199 VSS 0.0369f
C1804 VDD.t90 VSS 0.00595f
C1805 VDD.t95 VSS 0.00511f
C1806 VDD.t378 VSS 0.00387f
C1807 VDD.n200 VSS 0.01f
C1808 VDD.n201 VSS 0.00924f
C1809 VDD.t88 VSS 0.00511f
C1810 VDD.t382 VSS 0.00387f
C1811 VDD.n202 VSS 0.01f
C1812 VDD.n203 VSS 0.00399f
C1813 VDD.n204 VSS 4.13e-19
C1814 VDD.n205 VSS 0.00266f
C1815 VDD.n206 VSS 0.0419f
C1816 VDD.n207 VSS 0.0277f
C1817 VDD.n208 VSS 0.0185f
C1818 VDD.n209 VSS 0.0339f
C1819 VDD.n210 VSS 0.0348f
C1820 VDD.n211 VSS 0.0185f
C1821 VDD.n212 VSS 0.0339f
C1822 VDD.n213 VSS 0.0347f
C1823 VDD.n214 VSS 0.0206f
C1824 VDD.n215 VSS 0.0295f
C1825 VDD.n216 VSS 0.0274f
C1826 VDD.n217 VSS 0.0206f
C1827 VDD.n218 VSS 0.0519f
C1828 VDD.n219 VSS 0.0468f
C1829 VDD.n220 VSS 0.0328f
C1830 VDD.n221 VSS 0.0315f
C1831 VDD.n222 VSS 0.0185f
C1832 VDD.n223 VSS 0.0222f
C1833 VDD.n224 VSS 0.0101f
C1834 VDD.t115 VSS 0.00511f
C1835 VDD.t370 VSS 0.00387f
C1836 VDD.n225 VSS 0.00997f
C1837 VDD.n226 VSS 0.0423f
C1838 VDD.n227 VSS 0.0817f
C1839 VDD.n228 VSS 0.0165f
C1840 VDD.n229 VSS 0.00131f
C1841 VDD.t374 VSS 0.00386f
C1842 VDD.n230 VSS 0.00523f
C1843 VDD.t105 VSS 0.00496f
C1844 VDD.n231 VSS 0.0049f
C1845 VDD.n232 VSS 4.94e-20
C1846 VDD.n233 VSS 0.00154f
C1847 VDD.n234 VSS 7.08e-19
C1848 VDD.n235 VSS 5.88e-19
C1849 VDD.n236 VSS 0.00443f
C1850 VDD.n237 VSS 0.0139f
C1851 VDD.n238 VSS 0.034f
C1852 VDD.n239 VSS 0.0339f
C1853 VDD.n240 VSS 0.0348f
C1854 VDD.n241 VSS 0.0185f
C1855 VDD.n242 VSS 0.0339f
C1856 VDD.n243 VSS 0.0347f
C1857 VDD.n244 VSS 0.0206f
C1858 VDD.n245 VSS 0.0295f
C1859 VDD.n246 VSS 0.0274f
C1860 VDD.n247 VSS 0.0206f
C1861 VDD.n248 VSS 0.0527f
C1862 VDD.n249 VSS 0.0438f
C1863 VDD.t72 VSS 0.00592f
C1864 VDD.n250 VSS 0.0235f
C1865 VDD.t71 VSS 0.0602f
C1866 VDD.t73 VSS 0.0407f
C1867 VDD.t161 VSS 0.00245f
C1868 VDD.n251 VSS 0.00245f
C1869 VDD.n252 VSS 0.00534f
C1870 VDD.t136 VSS 0.00595f
C1871 VDD.n253 VSS 0.00595f
C1872 VDD.n254 VSS 0.0295f
C1873 VDD.t231 VSS 0.0786f
C1874 VDD.n255 VSS 0.00595f
C1875 VDD.t321 VSS 0.00595f
C1876 VDD.n256 VSS 0.00595f
C1877 VDD.n257 VSS 0.00595f
C1878 VDD.t177 VSS 0.0775f
C1879 VDD.n258 VSS 0.0369f
C1880 VDD.t248 VSS 0.00595f
C1881 VDD.n259 VSS 0.00595f
C1882 VDD.t247 VSS 0.0718f
C1883 VDD.t234 VSS 0.0786f
C1884 VDD.n260 VSS 0.0369f
C1885 VDD.t141 VSS 0.00595f
C1886 VDD.t332 VSS 0.00245f
C1887 VDD.n261 VSS 0.00245f
C1888 VDD.n262 VSS 0.00534f
C1889 VDD.t140 VSS 0.0718f
C1890 VDD.t331 VSS 0.0876f
C1891 VDD.t185 VSS 0.0407f
C1892 VDD.n263 VSS 0.0369f
C1893 VDD.t55 VSS 0.00595f
C1894 VDD.t182 VSS 0.00245f
C1895 VDD.n264 VSS 0.00245f
C1896 VDD.n265 VSS 0.00534f
C1897 VDD.t54 VSS 0.0718f
C1898 VDD.t181 VSS 0.0876f
C1899 VDD.t58 VSS 0.0407f
C1900 VDD.t116 VSS 0.0716f
C1901 VDD.n266 VSS 0.0369f
C1902 VDD.t117 VSS 0.00638f
C1903 VDD.n267 VSS 0.0458f
C1904 VDD.n268 VSS 0.0339f
C1905 VDD.n269 VSS 0.0348f
C1906 VDD.n270 VSS 0.0185f
C1907 VDD.n271 VSS 0.0339f
C1908 VDD.n272 VSS 0.0347f
C1909 VDD.n273 VSS 0.0206f
C1910 VDD.n274 VSS 0.0295f
C1911 VDD.n275 VSS 0.0274f
C1912 VDD.n276 VSS 0.0206f
C1913 VDD.n277 VSS 0.0561f
C1914 VDD.n278 VSS 0.0638f
C1915 VDD.t350 VSS 0.0775f
C1916 VDD.t320 VSS 0.0718f
C1917 VDD.n279 VSS 0.0369f
C1918 VDD.n280 VSS 0.0206f
C1919 VDD.n281 VSS 0.0274f
C1920 VDD.n282 VSS 0.0295f
C1921 VDD.t334 VSS 0.00595f
C1922 VDD.n283 VSS 0.0274f
C1923 VDD.n284 VSS 0.0206f
C1924 VDD.n285 VSS 0.0369f
C1925 VDD.t333 VSS 0.0718f
C1926 VDD.t137 VSS 0.0786f
C1927 VDD.t160 VSS 0.0876f
C1928 VDD.t135 VSS 0.0718f
C1929 VDD.n286 VSS 0.0369f
C1930 VDD.n287 VSS 0.0206f
C1931 VDD.n288 VSS 0.026f
C1932 VDD.n289 VSS 0.0192f
C1933 VDD.t63 VSS 0.00595f
C1934 VDD.n290 VSS 0.00595f
C1935 VDD.n291 VSS 0.0342f
C1936 VDD.t225 VSS 0.00593f
C1937 VDD.n292 VSS 0.0303f
C1938 VDD.t224 VSS 0.0536f
C1939 VDD.t180 VSS 0.0533f
C1940 VDD.t79 VSS 0.0528f
C1941 VDD.n293 VSS 0.0611f
C1942 VDD.t80 VSS 0.00596f
C1943 VDD.t240 VSS 0.0142f
C1944 VDD.n294 VSS 0.0432f
C1945 VDD.n295 VSS 0.0485f
C1946 VDD.n296 VSS 0.0359f
C1947 VDD.t239 VSS 0.0506f
C1948 VDD.n297 VSS 0.0928f
C1949 VDD.t42 VSS 0.0469f
C1950 VDD.t62 VSS 0.0716f
C1951 VDD.n298 VSS 0.0369f
C1952 VDD.n299 VSS 0.0231f
C1953 VDD.n300 VSS 0.0495f
C1954 VDD.t41 VSS 0.00595f
C1955 VDD.n301 VSS 0.0298f
C1956 VDD.n302 VSS 0.0464f
C1957 VDD.n303 VSS 0.0137f
C1958 VDD.n304 VSS 0.0369f
C1959 VDD.t40 VSS 0.036f
C1960 VDD.n305 VSS 0.0517f
C1961 VDD.n306 VSS 0.0794f
C1962 VDD.t344 VSS 0.0484f
C1963 VDD.n307 VSS 0.087f
C1964 VDD.n308 VSS 0.0401f
C1965 VDD.n309 VSS 0.0062f
C1966 VDD.n310 VSS 0.0393f
C1967 VDD.n311 VSS 0.00595f
C1968 VDD.n312 VSS 0.0233f
C1969 VDD.n313 VSS 0.0172f
C1970 VDD.n314 VSS 0.0627f
C1971 VDD.t254 VSS 0.0478f
C1972 VDD.t92 VSS 0.0481f
C1973 VDD.t124 VSS 0.0506f
C1974 VDD.t298 VSS 0.0797f
C1975 VDD.n315 VSS 0.0627f
C1976 VDD.n316 VSS 0.0191f
C1977 VDD.n317 VSS 0.0278f
C1978 VDD.n318 VSS 0.0251f
C1979 VDD.t362 VSS 0.00595f
C1980 VDD.n319 VSS 0.00595f
C1981 VDD.n320 VSS 0.0323f
C1982 VDD.n321 VSS 0.0306f
C1983 VDD.n322 VSS 0.0287f
C1984 VDD.n323 VSS 0.0598f
C1985 VDD.t361 VSS 0.0984f
C1986 VDD.t33 VSS 0.0987f
C1987 VDD.n324 VSS 0.0598f
C1988 VDD.n325 VSS 0.0133f
C1989 VDD.n326 VSS 0.0279f
C1990 VDD.n327 VSS 0.0279f
C1991 VDD.t145 VSS 0.00595f
C1992 VDD.n328 VSS 0.00595f
C1993 VDD.n329 VSS 0.0305f
C1994 VDD.n330 VSS 0.0324f
C1995 VDD.n331 VSS 0.0132f
C1996 VDD.n332 VSS 0.0598f
C1997 VDD.t144 VSS 0.0984f
C1998 VDD.t256 VSS 0.0987f
C1999 VDD.t220 VSS 0.0506f
C2000 VDD.t8 VSS 0.0319f
C2001 VDD.n333 VSS 0.0598f
C2002 VDD.n334 VSS 0.0288f
C2003 VDD.n335 VSS 0.0251f
C2004 VDD.n336 VSS 0.0277f
C2005 VDD.n337 VSS 0.00595f
C2006 VDD.t215 VSS 0.00595f
C2007 VDD.n338 VSS 0.0232f
C2008 VDD.n339 VSS 0.0235f
C2009 VDD.n340 VSS 0.0192f
C2010 VDD.n341 VSS 0.0627f
C2011 VDD.t214 VSS 0.0478f
C2012 VDD.t0 VSS 0.0481f
C2013 VDD.t155 VSS 0.0797f
C2014 VDD.n342 VSS 0.0627f
C2015 VDD.n343 VSS 0.0172f
C2016 VDD.t156 VSS 0.00595f
C2017 VDD.t274 VSS 0.00595f
C2018 VDD.t365 VSS 0.0719f
C2019 VDD.n344 VSS 0.00595f
C2020 VDD.t169 VSS 0.00245f
C2021 VDD.n345 VSS 0.00245f
C2022 VDD.n346 VSS 0.00534f
C2023 VDD.n347 VSS 0.00595f
C2024 VDD.n348 VSS 0.0348f
C2025 VDD.t85 VSS 0.0717f
C2026 VDD.n349 VSS 0.00595f
C2027 VDD.t383 VSS 0.00387f
C2028 VDD.t84 VSS 0.00511f
C2029 VDD.n350 VSS 0.01f
C2030 VDD.n351 VSS 0.00775f
C2031 VDD.t380 VSS 0.00387f
C2032 VDD.t91 VSS 0.00511f
C2033 VDD.n352 VSS 0.01f
C2034 VDD.n353 VSS 0.0412f
C2035 VDD.n354 VSS 0.0278f
C2036 VDD.t250 VSS 0.00245f
C2037 VDD.n355 VSS 0.00245f
C2038 VDD.n356 VSS 0.00534f
C2039 VDD.n357 VSS 0.0339f
C2040 VDD.n358 VSS 0.0184f
C2041 VDD.n359 VSS 0.0369f
C2042 VDD.t249 VSS 0.0405f
C2043 VDD.t275 VSS 0.0876f
C2044 VDD.t162 VSS 0.0719f
C2045 VDD.t259 VSS 0.0876f
C2046 VDD.t168 VSS 0.0405f
C2047 VDD.n360 VSS 0.0369f
C2048 VDD.n361 VSS 0.0184f
C2049 VDD.n362 VSS 0.0339f
C2050 VDD.n363 VSS 0.0347f
C2051 VDD.t219 VSS 0.00595f
C2052 VDD.n364 VSS 0.00595f
C2053 VDD.n365 VSS 0.0274f
C2054 VDD.n366 VSS 0.0295f
C2055 VDD.n367 VSS 0.0206f
C2056 VDD.n368 VSS 0.0369f
C2057 VDD.t218 VSS 0.0785f
C2058 VDD.t303 VSS 0.0719f
C2059 VDD.t273 VSS 0.0773f
C2060 VDD.n369 VSS 0.0369f
C2061 VDD.n370 VSS 0.0206f
C2062 VDD.n371 VSS 0.0508f
C2063 VDD.n372 VSS 0.0569f
C2064 VDD.n373 VSS 0.0231f
C2065 VDD.t66 VSS 0.132f
C2066 VDD.t67 VSS 0.00596f
.ends

