magic
tech gf180mcuC
magscale 1 10
timestamp 1691493873
<< nwell >>
rect -107 407 1332 953
<< pwell >>
rect -45 97 235 333
rect 350 97 1430 333
<< nmos >>
rect 67 165 123 265
rect 462 165 518 265
rect 622 165 678 265
rect 782 165 838 265
rect 942 165 998 265
rect 1102 165 1158 265
rect 1262 165 1318 265
<< pmos >>
rect 67 537 123 737
rect 462 537 518 737
rect 622 537 678 737
rect 782 537 838 737
rect 942 537 998 737
rect 1102 537 1158 737
<< ndiff >>
rect -21 252 67 265
rect -21 178 -8 252
rect 38 178 67 252
rect -21 165 67 178
rect 123 252 211 265
rect 123 178 152 252
rect 198 178 211 252
rect 123 165 211 178
rect 374 252 462 265
rect 374 178 387 252
rect 433 178 462 252
rect 374 165 462 178
rect 518 252 622 265
rect 518 178 547 252
rect 593 178 622 252
rect 518 165 622 178
rect 678 252 782 265
rect 678 178 707 252
rect 753 178 782 252
rect 678 165 782 178
rect 838 252 942 265
rect 838 178 867 252
rect 913 178 942 252
rect 838 165 942 178
rect 998 252 1102 265
rect 998 178 1027 252
rect 1073 178 1102 252
rect 998 165 1102 178
rect 1158 252 1262 265
rect 1158 178 1187 252
rect 1233 178 1262 252
rect 1158 165 1262 178
rect 1318 252 1406 265
rect 1318 178 1347 252
rect 1393 178 1406 252
rect 1318 165 1406 178
<< pdiff >>
rect -21 724 67 737
rect -21 550 -8 724
rect 38 550 67 724
rect -21 537 67 550
rect 123 724 211 737
rect 123 550 152 724
rect 198 550 211 724
rect 123 537 211 550
rect 374 724 462 737
rect 374 550 387 724
rect 433 550 462 724
rect 374 537 462 550
rect 518 724 622 737
rect 518 550 547 724
rect 593 550 622 724
rect 518 537 622 550
rect 678 724 782 737
rect 678 550 707 724
rect 753 550 782 724
rect 678 537 782 550
rect 838 724 942 737
rect 838 550 867 724
rect 913 550 942 724
rect 838 537 942 550
rect 998 724 1102 737
rect 998 550 1027 724
rect 1073 550 1102 724
rect 998 537 1102 550
rect 1158 724 1246 737
rect 1158 550 1187 724
rect 1233 550 1246 724
rect 1158 537 1246 550
<< ndiffc >>
rect -8 178 38 252
rect 152 178 198 252
rect 387 178 433 252
rect 547 178 593 252
rect 707 178 753 252
rect 867 178 913 252
rect 1027 178 1073 252
rect 1187 178 1233 252
rect 1347 178 1393 252
<< pdiffc >>
rect -8 550 38 724
rect 152 550 198 724
rect 387 550 433 724
rect 547 550 593 724
rect 707 550 753 724
rect 867 550 913 724
rect 1027 550 1073 724
rect 1187 550 1233 724
<< psubdiff >>
rect -35 52 225 65
rect -35 6 -22 52
rect 24 6 72 52
rect 118 6 166 52
rect 212 6 225 52
rect -35 -7 225 6
<< nsubdiff >>
rect -82 907 272 920
rect -82 861 -69 907
rect -23 861 25 907
rect 71 861 119 907
rect 165 861 213 907
rect 259 861 272 907
rect -82 848 272 861
<< psubdiffcont >>
rect -22 6 24 52
rect 72 6 118 52
rect 166 6 212 52
<< nsubdiffcont >>
rect -69 861 -23 907
rect 25 861 71 907
rect 119 861 165 907
rect 213 861 259 907
<< polysilicon >>
rect 67 737 123 781
rect 462 757 1158 801
rect 462 737 518 757
rect 622 737 678 757
rect 782 737 838 757
rect 942 737 998 757
rect 1102 737 1158 757
rect 67 371 123 537
rect 227 498 299 506
rect 462 498 518 537
rect 227 493 518 498
rect 622 493 678 537
rect 782 493 838 537
rect 942 493 998 537
rect 1102 493 1158 537
rect 227 447 240 493
rect 286 447 518 493
rect 227 442 518 447
rect 227 434 299 442
rect 171 371 243 379
rect 67 366 518 371
rect 67 320 184 366
rect 230 320 518 366
rect 67 315 518 320
rect 67 265 123 315
rect 171 307 243 315
rect 462 265 518 315
rect 622 265 678 309
rect 782 265 838 309
rect 942 265 998 309
rect 1102 265 1158 309
rect 1262 265 1318 309
rect 67 121 123 165
rect 462 145 518 165
rect 622 145 678 165
rect 782 145 838 165
rect 942 145 998 165
rect 1102 145 1158 165
rect 1262 145 1318 165
rect 462 101 1318 145
<< polycontact >>
rect 240 447 286 493
rect 184 320 230 366
<< metal1 >>
rect -107 907 297 940
rect -107 861 -69 907
rect -23 861 25 907
rect 71 861 119 907
rect 165 861 213 907
rect 259 861 297 907
rect -107 828 297 861
rect -8 724 38 735
rect -8 493 38 550
rect 152 724 198 828
rect 152 539 198 550
rect 387 781 1073 827
rect 387 724 433 781
rect 229 493 297 504
rect -105 447 240 493
rect 286 447 297 493
rect -8 252 38 447
rect 229 436 297 447
rect 173 366 241 377
rect 173 320 184 366
rect 230 320 295 366
rect 173 309 241 320
rect -8 167 38 178
rect 152 252 198 263
rect 152 85 198 178
rect 387 252 433 550
rect 547 724 593 735
rect 547 493 593 550
rect 707 724 753 781
rect 707 539 753 550
rect 867 724 913 735
rect 867 493 913 550
rect 1027 724 1073 781
rect 1027 539 1073 550
rect 1187 724 1233 735
rect 1187 493 1233 550
rect 547 447 1337 493
rect 1187 355 1233 447
rect 387 121 433 178
rect 547 309 1233 355
rect 547 252 593 309
rect 547 167 593 178
rect 707 252 753 263
rect 707 121 753 178
rect 867 252 913 309
rect 867 167 913 178
rect 1027 252 1073 263
rect 1027 121 1073 178
rect 1187 252 1233 309
rect 1187 167 1233 178
rect 1347 304 1482 350
rect 1347 252 1393 304
rect 1347 121 1393 178
rect -55 52 245 85
rect 387 75 1393 121
rect -55 6 -22 52
rect 24 6 72 52
rect 118 6 166 52
rect 212 6 245 52
rect -55 -27 245 6
<< labels >>
flabel metal1 1436 326 1436 326 0 FreeSans 320 0 0 0 VOUT
port 3 nsew
flabel metal1 1296 470 1296 470 0 FreeSans 320 0 0 0 VIN
port 2 nsew
flabel metal1 95 29 95 29 0 FreeSans 320 0 0 0 VSS
port 4 nsew
flabel polysilicon 207 343 207 343 0 FreeSans 320 0 0 0 CLK
port 6 nsew
flabel metal1 95 887 95 887 0 FreeSans 320 0 0 0 VDD
port 5 nsew
flabel psubdiffcont 95 29 95 29 0 FreeSans 320 0 0 0 Inverter_Layout_0.VSS
flabel metal1 95 887 95 887 0 FreeSans 320 0 0 0 Inverter_Layout_0.VDD
flabel metal1 275 343 275 343 0 FreeSans 320 0 0 0 Inverter_Layout_0.IN
flabel metal1 -44 470 -44 470 0 FreeSans 320 0 0 0 Inverter_Layout_0.OUT
<< end >>
