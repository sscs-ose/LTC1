magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2496 -2083 6434 4575
<< isosubstrate >>
rect -496 -83 693 2575
<< nwell >>
rect -247 1551 693 2575
rect 1033 1281 4434 2575
<< polysilicon >>
rect -92 1107 48 1431
rect 152 1034 292 1867
rect 1411 1106 1551 1478
rect 1655 514 1795 1478
rect 1899 514 2039 1478
rect 2143 1106 2283 1478
rect 2559 614 2699 1478
rect 2803 614 2943 1478
rect 3047 614 3187 1478
rect 3291 614 3431 1478
rect 3535 614 3675 1478
rect 3779 614 3919 1478
<< metal1 >>
rect -85 2413 1 2481
rect 62 1811 138 2481
rect 445 2413 531 2481
rect 1195 2413 1281 2481
rect 306 1441 382 2211
rect 1321 1522 1397 2481
rect 1565 1442 1641 1958
rect 1809 1522 1885 2465
rect 2053 1442 2129 1958
rect 2297 1522 2373 2465
rect 2469 1522 2545 2465
rect 2713 1442 2789 2222
rect 2957 1522 3033 2465
rect 3201 1442 3277 2222
rect 3445 1522 3521 2465
rect 3588 2413 4272 2481
rect 3689 1442 3765 2222
rect 3933 1522 4009 2413
rect 306 1341 937 1441
rect 1565 1366 2667 1442
rect 2713 1366 4066 1442
rect -385 11 -332 79
rect -85 11 1 79
rect 62 11 138 990
rect 306 263 382 1341
rect 837 1276 937 1341
rect 2591 1276 2667 1366
rect 837 1114 2247 1276
rect 2591 1114 3859 1276
rect 2591 819 2667 1114
rect 3990 819 4066 1366
rect 1809 743 2667 819
rect 2713 743 4066 819
rect 440 11 540 79
rect 1195 11 1281 79
rect 1565 14 1641 470
rect 1809 270 1885 743
rect 2053 14 2129 470
rect 2469 14 2545 570
rect 2713 270 2789 743
rect 2957 14 3033 570
rect 3201 270 3277 743
rect 3445 14 3521 570
rect 3689 270 3765 743
rect 3931 79 4007 570
rect 3605 11 4255 79
<< metal2 >>
rect -135 435 314 573
use M1_NWELL_CDNS_40661953145273  M1_NWELL_CDNS_40661953145273_0
timestamp 1713338890
transform 1 0 223 0 1 2447
box -316 -128 316 128
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_0
timestamp 1713338890
transform 1 0 1161 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_1
timestamp 1713338890
transform 1 0 4255 0 1 1977
box -128 -598 128 598
use M1_NWELL_CDNS_40661953145325  M1_NWELL_CDNS_40661953145325_0
timestamp 1713338890
transform 1 0 2693 0 1 2447
box -1538 -128 1538 128
use M1_NWELL_CDNS_40661953145328  M1_NWELL_CDNS_40661953145328_0
timestamp 1713338890
transform 1 0 -119 0 1 2118
box -128 -457 128 457
use M1_NWELL_CDNS_40661953145328  M1_NWELL_CDNS_40661953145328_1
timestamp 1713338890
transform 1 0 565 0 1 2118
box -128 -457 128 457
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform 1 0 1969 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform 1 0 1481 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_2
timestamp 1713338890
transform 1 0 1725 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_3
timestamp 1713338890
transform 1 0 3117 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_4
timestamp 1713338890
transform 1 0 3361 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_5
timestamp 1713338890
transform 1 0 2213 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_6
timestamp 1713338890
transform 1 0 2873 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_7
timestamp 1713338890
transform 1 0 2629 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_8
timestamp 1713338890
transform 1 0 3605 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_9
timestamp 1713338890
transform 1 0 3849 0 1 1195
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_10
timestamp 1713338890
transform 1 0 222 0 1 1342
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_11
timestamp 1713338890
transform 1 0 -24 0 1 1342
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 1 0 1161 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 1 0 4289 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165612  M1_PSUB_CDNS_69033583165612_0
timestamp 1713338890
transform 1 0 72 0 -1 45
box -421 -45 421 45
use M1_PSUB_CDNS_69033583165618  M1_PSUB_CDNS_69033583165618_0
timestamp 1713338890
transform 1 0 2725 0 -1 45
box -1455 -45 1455 45
use M1_PSUB_CDNS_69033583165619  M1_PSUB_CDNS_69033583165619_0
timestamp 1713338890
transform 1 0 -398 0 -1 609
box -45 -609 45 609
use M1_PSUB_CDNS_69033583165619  M1_PSUB_CDNS_69033583165619_1
timestamp 1713338890
transform 1 0 565 0 -1 609
box -45 -609 45 609
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_0
timestamp 1713338890
transform 1 0 -144 0 1 514
box -38 -194 38 194
use M2_M1_CDNS_69033583165588  M2_M1_CDNS_69033583165588_1
timestamp 1713338890
transform 1 0 344 0 1 514
box -38 -194 38 194
use nmos_6p0_CDNS_4066195314547  nmos_6p0_CDNS_4066195314547_0
timestamp 1713338890
transform 1 0 -92 0 1 263
box -88 -44 472 844
use nmos_6p0_CDNS_4066195314549  nmos_6p0_CDNS_4066195314549_0
timestamp 1713338890
transform 1 0 2559 0 1 270
box -88 -44 1448 344
use nmos_6p0_CDNS_4066195314550  nmos_6p0_CDNS_4066195314550_0
timestamp 1713338890
transform 1 0 1655 0 1 270
box -88 -44 472 294
use pmos_6p0_CDNS_4066195314539  pmos_6p0_CDNS_4066195314539_0
timestamp 1713338890
transform 1 0 152 0 1 1811
box -208 -120 348 520
use pmos_6p0_CDNS_4066195314546  pmos_6p0_CDNS_4066195314546_0
timestamp 1713338890
transform 1 0 1411 0 1 1522
box -208 -120 1080 620
use pmos_6p0_CDNS_4066195314548  pmos_6p0_CDNS_4066195314548_0
timestamp 1713338890
transform 1 0 2559 0 1 1522
box -208 -120 1568 820
<< labels >>
rlabel metal1 s 225 1326 225 1326 4 A
port 1 nsew
rlabel metal1 s -21 1326 -21 1326 4 A
port 1 nsew
rlabel metal1 s 3512 1200 3512 1200 4 Z
port 2 nsew
rlabel metal1 s 1482 45 1482 45 4 VSS
port 3 nsew
rlabel metal1 s 1852 2452 1852 2452 4 VDD
port 4 nsew
rlabel metal1 s 80 45 80 45 4 DVSS
port 5 nsew
rlabel metal1 s 2 2452 2 2452 4 DVDD
port 6 nsew
<< end >>
