* NGSPICE file created from dec_2x4_ibr_mag_flat.ext - technology: gf180mcuC

.subckt pex_dec_2x4_ibr_mag IN1 VSS VDD D0 D1 D2 D3 IN2
X0 D0 nand2_0.OUT VDD.t14 VDD.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 nand2_1.OUT IN1.t0 VDD.t6 VDD.t5 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 a_2170_257# nand2_2.IN2 VSS.t15 VSS.t14 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3 nand2_3.OUT IN2.t0 a_3136_257# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X4 D2 nand2_2.OUT VDD.t26 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X5 nand2_0.OUT nand2_1.IN1 a_238_256# VSS.t1 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X6 a_1204_257# IN1.t1 VSS.t7 VSS.t6 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X7 nand2_2.OUT IN2.t1 a_2170_257# VSS.t20 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X8 D3 nand2_3.OUT VSS.t19 VSS.t18 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X9 nand2_1.IN1 IN2.t2 VSS.t23 VSS.t22 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X10 D0 nand2_0.OUT VSS.t9 VSS.t8 nfet_03v3 ad=0.168p pd=1.77u as=0.152p ps=1.64u w=0.22u l=0.28u
X11 nand2_3.OUT IN1.t2 VDD.t18 VDD.t17 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X12 D2 nand2_2.OUT VSS.t17 VSS.t16 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X13 VDD nand2_1.IN1 nand2_1.OUT VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X14 nand2_0.OUT nand2_2.IN2 VDD.t24 VDD.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 D1 nand2_1.OUT VDD.t20 VDD.t19 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X16 nand2_2.IN2 IN1.t3 VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X17 a_3136_257# IN1.t4 VSS.t5 VSS.t4 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X18 nand2_1.OUT nand2_1.IN1 a_1204_257# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X19 a_238_256# nand2_2.IN2 VSS.t13 VSS.t12 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X20 VDD IN2.t3 nand2_3.OUT VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X21 nand2_2.OUT nand2_2.IN2 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X22 D1 nand2_1.OUT VSS.t11 VSS.t10 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X23 nand2_2.IN2 IN1.t5 VSS.t3 VSS.t2 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X24 D3 nand2_3.OUT VDD.t28 VDD.t27 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X25 VDD nand2_1.IN1 nand2_0.OUT VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X26 VDD IN2.t4 nand2_2.OUT VDD.t29 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X27 nand2_1.IN1 IN2.t5 VDD.t16 VDD.t15 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 VDD.n21 VDD.t5 882.577
R1 VDD.t23 VDD.n26 763.259
R2 VDD.n15 VDD.t17 763.259
R3 VDD.n17 VDD.t21 763.259
R4 VDD.t29 VDD.t25 761.365
R5 VDD.t10 VDD.t19 761.365
R6 VDD.n28 VDD.t7 759.471
R7 VDD.t2 VDD.t27 746.062
R8 VDD.n29 VDD.n21 376.894
R9 VDD.t7 VDD.n27 193.183
R10 VDD.n9 VDD.t2 193.183
R11 VDD.n16 VDD.t29 193.183
R12 VDD.n19 VDD.t10 193.183
R13 VDD.n27 VDD.t23 109.849
R14 VDD.n9 VDD.t17 109.849
R15 VDD.t21 VDD.n16 109.849
R16 VDD.t5 VDD.n19 109.849
R17 VDD.n7 VDD.n0 35.263
R18 VDD.n30 VDD.n29 6.3005
R19 VDD.n27 VDD 6.3005
R20 VDD.n26 VDD.n25 6.3005
R21 VDD.n34 VDD.n17 6.3005
R22 VDD VDD.n19 6.3005
R23 VDD VDD.n9 6.3005
R24 VDD.n15 VDD.n14 6.3005
R25 VDD VDD.n16 6.3005
R26 VDD.n25 VDD.t1 5.19258
R27 VDD.n33 VDD.t20 5.14703
R28 VDD.n20 VDD.t14 5.14703
R29 VDD.n5 VDD.t28 5.14703
R30 VDD.n2 VDD.t16 5.14703
R31 VDD.n13 VDD.t26 5.14703
R32 VDD.n24 VDD.t24 5.13746
R33 VDD.n31 VDD.t6 5.13746
R34 VDD.n10 VDD.t18 5.13746
R35 VDD.n35 VDD.t22 5.13746
R36 VDD.n23 VDD.n22 5.13287
R37 VDD.n32 VDD.n18 5.13287
R38 VDD.n4 VDD.n3 5.13287
R39 VDD.n12 VDD.n11 5.13287
R40 VDD.n0 VDD.t15 4.96868
R41 VDD.n1 VDD.n0 3.1505
R42 VDD.n7 VDD.n6 3.1505
R43 VDD.n8 VDD.n7 3.1505
R44 VDD.n29 VDD.t13 1.89444
R45 VDD.t13 VDD.n28 1.89444
R46 VDD.n26 VDD.t0 1.89444
R47 VDD.t25 VDD.n15 1.89444
R48 VDD.t19 VDD.n17 1.89444
R49 VDD.t27 VDD.n8 1.81868
R50 VDD.n31 VDD 0.5425
R51 VDD VDD.n24 0.183056
R52 VDD VDD.n10 0.183056
R53 VDD VDD.n2 0.178278
R54 VDD.n23 VDD.n20 0.136194
R55 VDD.n33 VDD.n32 0.136194
R56 VDD.n5 VDD.n4 0.136194
R57 VDD.n13 VDD.n12 0.136194
R58 VDD VDD.n23 0.106177
R59 VDD.n32 VDD 0.106177
R60 VDD.n4 VDD 0.106177
R61 VDD.n12 VDD 0.106177
R62 VDD.n24 VDD 0.0800484
R63 VDD VDD.n31 0.0800484
R64 VDD.n10 VDD 0.0800484
R65 VDD VDD.n35 0.0800484
R66 VDD.n35 VDD 0.0498548
R67 VDD.n34 VDD.n33 0.0460556
R68 VDD.n30 VDD.n20 0.0460556
R69 VDD.n2 VDD.n1 0.0460556
R70 VDD.n6 VDD.n5 0.0460556
R71 VDD.n14 VDD.n13 0.0460556
R72 VDD.n25 VDD 0.00105556
R73 VDD VDD.n34 0.00105556
R74 VDD VDD.n30 0.00105556
R75 VDD.n1 VDD 0.00105556
R76 VDD.n6 VDD 0.00105556
R77 VDD.n14 VDD 0.00105556
R78 D0 D0.n0 5.13104
R79 D0.n2 D0.n1 4.5882
R80 D0 D0.n3 2.25244
R81 D0 D0.n2 1.5388
R82 D0.n2 D0 0.253082
R83 IN1.n0 IN1.t0 30.9379
R84 IN1.n1 IN1.t2 30.9379
R85 IN1.n5 IN1.t3 25.7638
R86 IN1.n0 IN1.t1 21.6422
R87 IN1.n1 IN1.t4 21.6422
R88 IN1.n5 IN1.t5 13.2969
R89 IN1.n4 IN1.n3 7.96122
R90 IN1.n6 IN1.n4 5.39718
R91 IN1.n3 IN1 4.52412
R92 IN1 IN1.n0 4.00388
R93 IN1 IN1.n5 4.00252
R94 IN1.n4 IN1 2.96831
R95 IN1.n2 IN1.n1 2.8805
R96 IN1.n6 IN1 2.373
R97 IN1.n8 IN1.n7 2.25347
R98 IN1.n3 IN1.n2 1.16475
R99 IN1.n8 IN1.n6 0.551491
R100 IN1 IN1.n2 0.003875
R101 IN1 IN1.n8 0.00346703
R102 VSS.t21 VSS.t18 2523.61
R103 VSS.n15 VSS.t12 1243.37
R104 VSS.n9 VSS.t4 1241.02
R105 VSS.n13 VSS.t6 1241.02
R106 VSS.t1 VSS.n13 1231.06
R107 VSS.t20 VSS.n9 1228.73
R108 VSS.t0 VSS.n11 1228.73
R109 VSS.n9 VSS.t16 1061.88
R110 VSS.n11 VSS.t10 1061.88
R111 VSS.n13 VSS.t8 1053.84
R112 VSS.n15 VSS.t2 1053.84
R113 VSS.n14 VSS.t1 590.909
R114 VSS.n5 VSS.t21 589.793
R115 VSS.n10 VSS.t20 589.793
R116 VSS.n12 VSS.t0 589.793
R117 VSS.t12 VSS.n14 393.94
R118 VSS.n5 VSS.t4 393.195
R119 VSS.n10 VSS.t14 393.195
R120 VSS.t6 VSS.n12 393.195
R121 VSS.n19 VSS.n13 375.25
R122 VSS.n16 VSS.n15 375.25
R123 VSS.n9 VSS.n8 367.205
R124 VSS.n22 VSS.n11 367.205
R125 VSS.n4 VSS.n0 35.7094
R126 VSS VSS.t3 9.40995
R127 VSS.n21 VSS.t11 9.34566
R128 VSS.n18 VSS.t9 9.34566
R129 VSS.n1 VSS.t23 9.34566
R130 VSS.n2 VSS.t19 9.34566
R131 VSS.n7 VSS.t17 9.34566
R132 VSS.n23 VSS.t15 7.19156
R133 VSS.n20 VSS.t7 7.19156
R134 VSS.n17 VSS.t13 7.19156
R135 VSS.n6 VSS.t5 7.19156
R136 VSS VSS.n5 5.2005
R137 VSS VSS.n14 5.2005
R138 VSS VSS.n12 5.2005
R139 VSS VSS.n10 5.2005
R140 VSS VSS.n0 2.60126
R141 VSS.n0 VSS.t22 2.6005
R142 VSS.t18 VSS.n4 2.6005
R143 VSS.n4 VSS.n3 2.6005
R144 VSS.n2 VSS 0.375997
R145 VSS.n18 VSS 0.375997
R146 VSS.n21 VSS 0.375997
R147 VSS.n23 VSS.n22 0.341085
R148 VSS.n8 VSS.n6 0.338957
R149 VSS.n17 VSS.n16 0.312136
R150 VSS.n20 VSS.n19 0.310702
R151 VSS.n3 VSS.n1 0.240248
R152 VSS.n7 VSS 0.189392
R153 VSS.n6 VSS 0.118573
R154 VSS VSS.n17 0.118573
R155 VSS VSS.n20 0.118573
R156 VSS VSS.n23 0.118573
R157 VSS.n1 VSS 0.0647857
R158 VSS VSS.n2 0.0647857
R159 VSS VSS.n7 0.0647857
R160 VSS VSS.n18 0.0647857
R161 VSS VSS.n21 0.0647857
R162 VSS.n3 VSS 0.0012563
R163 VSS.n8 VSS 0.0012563
R164 VSS.n16 VSS 0.0012563
R165 VSS.n19 VSS 0.0012563
R166 VSS.n22 VSS 0.0012563
R167 IN2.n0 IN2.t0 31.528
R168 IN2.n1 IN2.t1 31.528
R169 IN2.n3 IN2.t5 25.7638
R170 IN2.n0 IN2.t3 15.3826
R171 IN2.n1 IN2.t4 15.3826
R172 IN2.n3 IN2.t2 13.2969
R173 IN2 IN2.n1 8.85842
R174 IN2 IN2.n0 8.85606
R175 IN2.n2 IN2 6.02672
R176 IN2.n2 IN2 2.58284
R177 IN2.n7 IN2.n6 2.25518
R178 IN2.n4 IN2.n3 2.12228
R179 IN2.n5 IN2.n4 1.13447
R180 IN2.n7 IN2.n5 1.09227
R181 IN2.n5 IN2.n2 0.907343
R182 IN2 IN2.n7 0.00391772
R183 IN2.n4 IN2 0.00125099
R184 D2.n2 D2.n1 6.40201
R185 D2 D2.n0 5.13104
R186 D2.n4 D2.n3 2.25277
R187 D2.n4 D2.n2 1.53231
R188 D2.n2 D2 0.247244
R189 D2 D2.n4 0.00276891
R190 D3.n2 D3.n0 6.53652
R191 D3 D3.n1 5.13104
R192 D3.n4 D3.n3 2.25428
R193 D3.n4 D3.n2 1.577
R194 D3.n2 D3 0.261217
R195 D3 D3.n4 0.00428151
R196 D1.n2 D1.n1 7.86708
R197 D1 D1.n0 5.13104
R198 D1.n4 D1.n3 2.25819
R199 D1.n4 D1.n2 1.31873
R200 D1.n2 D1 0.243273
R201 D1 D1.n4 0.00819231
C0 IN1 nand2_3.OUT 0.107f
C1 VDD D3 0.122f
C2 VDD nand2_1.OUT 0.395f
C3 nand2_1.IN1 a_1204_257# 0.00352f
C4 nand2_1.OUT nand2_0.OUT 7.53e-19
C5 VDD a_2170_257# 3.14e-19
C6 nand2_2.IN2 D3 6.22e-21
C7 nand2_1.OUT nand2_2.IN2 0.0784f
C8 a_2170_257# nand2_0.OUT 3.72e-22
C9 D0 nand2_1.OUT 0.00978f
C10 a_2170_257# nand2_2.IN2 0.00347f
C11 D2 D1 0.0188f
C12 IN2 a_3136_257# 0.00556f
C13 nand2_2.OUT IN2 0.359f
C14 nand2_2.OUT a_3136_257# 9.69e-20
C15 VDD a_1204_257# 3.14e-19
C16 D2 nand2_3.OUT 0.0257f
C17 IN1 IN2 0.454f
C18 IN1 a_238_256# 8.25e-19
C19 IN1 a_3136_257# 0.0035f
C20 nand2_0.OUT a_1204_257# 1e-19
C21 nand2_2.OUT IN1 0.106f
C22 nand2_2.IN2 a_1204_257# 0.00375f
C23 D0 a_1204_257# 0.00173f
C24 nand2_1.OUT D1 0.129f
C25 D3 nand2_3.OUT 0.143f
C26 a_2170_257# D1 0.00171f
C27 D1 a_1204_257# 8.39e-19
C28 D2 IN2 0.0475f
C29 D2 a_3136_257# 0.00171f
C30 D2 nand2_2.OUT 0.129f
C31 VDD nand2_1.IN1 1.72f
C32 D2 IN1 0.0997f
C33 nand2_1.IN1 nand2_0.OUT 0.361f
C34 nand2_2.IN2 nand2_1.IN1 0.699f
C35 IN2 D3 0.123f
C36 D3 a_3136_257# 9.03e-19
C37 nand2_2.OUT D3 1.82e-20
C38 nand2_1.OUT nand2_2.OUT 7.49e-19
C39 D0 nand2_1.IN1 0.0457f
C40 VDD nand2_0.OUT 0.397f
C41 a_2170_257# IN2 0.00348f
C42 IN1 D3 0.00153f
C43 a_2170_257# nand2_2.OUT 0.0705f
C44 VDD nand2_2.IN2 0.546f
C45 nand2_1.OUT IN1 0.146f
C46 VDD D0 0.124f
C47 nand2_2.IN2 nand2_0.OUT 0.195f
C48 a_2170_257# IN1 0.00307f
C49 D0 nand2_0.OUT 0.128f
C50 D0 nand2_2.IN2 0.0719f
C51 nand2_1.IN1 D1 0.046f
C52 IN1 a_1204_257# 0.00347f
C53 nand2_1.IN1 nand2_3.OUT 0.0256f
C54 VDD D1 0.169f
C55 D2 D3 0.019f
C56 VDD nand2_3.OUT 0.401f
C57 D1 nand2_0.OUT 1.18e-21
C58 nand2_2.IN2 D1 0.0992f
C59 D2 a_2170_257# 8.5e-19
C60 D0 D1 0.0193f
C61 nand2_1.IN1 IN2 0.827f
C62 nand2_1.IN1 a_238_256# 0.00348f
C63 nand2_2.OUT nand2_1.IN1 0.0122f
C64 nand2_1.OUT a_2170_257# 9.69e-20
C65 IN1 nand2_1.IN1 0.874f
C66 VDD IN2 0.82f
C67 VDD a_238_256# 3.14e-19
C68 VDD a_3136_257# 3.14e-19
C69 VDD nand2_2.OUT 0.407f
C70 nand2_1.OUT a_1204_257# 0.0691f
C71 D1 nand2_3.OUT 1.96e-21
C72 a_238_256# nand2_0.OUT 0.0691f
C73 nand2_2.OUT nand2_0.OUT 4.89e-22
C74 VDD IN1 1.46f
C75 nand2_2.IN2 IN2 0.0465f
C76 nand2_2.IN2 a_238_256# 0.00719f
C77 nand2_2.OUT nand2_2.IN2 0.101f
C78 D0 IN2 6.05e-21
C79 D0 a_238_256# 8.3e-19
C80 D0 nand2_2.OUT 2.62e-21
C81 IN1 nand2_0.OUT 0.0355f
C82 IN1 nand2_2.IN2 0.341f
C83 D0 IN1 0.271f
C84 D2 nand2_1.IN1 0.00879f
C85 IN2 D1 0.00201f
C86 nand2_2.OUT D1 0.0258f
C87 VDD D2 0.17f
C88 IN2 nand2_3.OUT 0.415f
C89 nand2_3.OUT a_3136_257# 0.0691f
C90 nand2_2.OUT nand2_3.OUT 7.49e-19
C91 IN1 D1 0.0238f
C92 nand2_1.IN1 D3 0.385f
C93 nand2_1.OUT nand2_1.IN1 0.377f
C94 D2 nand2_2.IN2 9.49e-19
C95 a_3136_257# VSS 0.0676f
C96 a_2170_257# VSS 0.0675f
C97 D3 VSS 0.572f
C98 a_1204_257# VSS 0.0676f
C99 nand2_3.OUT VSS 0.433f
C100 D2 VSS 0.633f
C101 a_238_256# VSS 0.0678f
C102 nand2_2.OUT VSS 0.442f
C103 D1 VSS 0.599f
C104 IN2 VSS 1.14f
C105 nand2_1.OUT VSS 0.442f
C106 D0 VSS 0.592f
C107 nand2_0.OUT VSS 0.443f
C108 nand2_1.IN1 VSS 1.19f
C109 nand2_2.IN2 VSS 1.01f
C110 IN1 VSS 1.95f
C111 VDD VSS 8.49f
.ends

