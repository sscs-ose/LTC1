magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 4032 71968
<< psubdiff >>
rect 0 69778 2000 69968
rect 0 13287 93 69778
rect 1907 13287 2000 69778
rect 0 13097 2000 13287
<< metal1 >>
rect -32 69789 2032 69957
rect -32 13276 14 69789
rect 1986 13276 2032 69789
rect -32 13108 2032 13276
<< metal2 >>
rect 81 65000 282 69518
rect 0 63600 282 65000
rect 81 50600 282 63600
rect 0 49200 282 50600
rect 81 13611 282 49200
rect 418 23563 694 68152
rect 1349 14031 1591 69620
rect 1717 65000 1918 69518
rect 1717 63600 2000 65000
rect 1717 50600 1918 63600
rect 1717 49200 2000 50600
rect 1717 13611 1918 49200
<< metal3 >>
rect 0 68400 2000 69678
rect 0 66800 2000 68200
rect 0 65200 2000 66600
rect 0 63600 2000 65000
rect 0 62000 2000 63400
rect 0 60400 2000 61800
rect 0 58800 2000 60200
rect 0 57200 2000 58600
rect 0 55600 2000 57000
rect 0 54000 2000 55400
rect 0 52400 2000 53800
rect 0 50800 2000 52200
rect 0 49200 2000 50600
rect 0 46000 2000 49000
rect 0 42800 2000 45800
rect 0 41200 2000 42600
rect 0 39600 2000 41000
rect 0 36400 2000 39400
rect 0 33200 2000 36200
rect 0 30000 2000 33000
rect 0 26800 2000 29800
rect 0 25200 2000 26600
rect 0 23600 2000 25000
rect 0 20400 2000 23400
rect 0 17200 2000 20200
rect 0 14000 2000 17000
use M1_PSUB_CDNS_690335831656  M1_PSUB_CDNS_690335831656_0
timestamp 1713338890
transform 1 0 1952 0 1 41524
box -45 -28395 45 28395
use M1_PSUB_CDNS_690335831656  M1_PSUB_CDNS_690335831656_1
timestamp 1713338890
transform -1 0 48 0 1 41524
box -45 -28395 45 28395
use M1_PSUB_CDNS_6903358316568  M1_PSUB_CDNS_6903358316568_0
timestamp 1713338890
transform 1 0 1001 0 -1 13192
box -845 -95 845 95
use M1_PSUB_CDNS_6903358316568  M1_PSUB_CDNS_6903358316568_1
timestamp 1713338890
transform 1 0 1001 0 1 69873
box -845 -95 845 95
use M2_M1_CDNS_6903358316571  M2_M1_CDNS_6903358316571_0
timestamp 1713338890
transform 1 0 1818 0 1 49901
box -100 -596 100 596
use M2_M1_CDNS_6903358316571  M2_M1_CDNS_6903358316571_1
timestamp 1713338890
transform 1 0 182 0 1 49901
box -100 -596 100 596
use M2_M1_CDNS_6903358316571  M2_M1_CDNS_6903358316571_2
timestamp 1713338890
transform 1 0 1818 0 1 64300
box -100 -596 100 596
use M2_M1_CDNS_6903358316571  M2_M1_CDNS_6903358316571_3
timestamp 1713338890
transform 1 0 182 0 1 64300
box -100 -596 100 596
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_0
timestamp 1713338890
transform 1 0 1475 0 1 15532
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_1
timestamp 1713338890
transform 1 0 1475 0 1 18722
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_2
timestamp 1713338890
transform 1 0 1475 0 1 21869
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_3
timestamp 1713338890
transform 1 0 552 0 1 28350
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_4
timestamp 1713338890
transform 1 0 552 0 1 31492
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_5
timestamp 1713338890
transform 1 0 552 0 1 34717
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_6
timestamp 1713338890
transform 1 0 552 0 1 37938
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_7
timestamp 1713338890
transform 1 0 552 0 1 44259
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_8
timestamp 1713338890
transform 1 0 1475 0 1 47483
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_0
timestamp 1713338890
transform 1 0 552 0 1 24301
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_1
timestamp 1713338890
transform 1 0 1475 0 1 25934
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_2
timestamp 1713338890
transform 1 0 552 0 1 41900
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_3
timestamp 1713338890
transform 1 0 1475 0 1 40328
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_4
timestamp 1713338890
transform 1 0 552 0 1 53091
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_5
timestamp 1713338890
transform 1 0 552 0 1 54705
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_6
timestamp 1713338890
transform 1 0 552 0 1 56328
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_7
timestamp 1713338890
transform 1 0 552 0 1 59480
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_8
timestamp 1713338890
transform 1 0 1475 0 1 57883
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_9
timestamp 1713338890
transform 1 0 1475 0 1 61121
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_10
timestamp 1713338890
transform 1 0 1475 0 1 65917
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_11
timestamp 1713338890
transform 1 0 552 0 1 67457
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_12
timestamp 1713338890
transform 1 0 1475 0 1 69054
box -38 -566 38 566
use M3_M2_CDNS_6903358316569  M3_M2_CDNS_6903358316569_0
timestamp 1713338890
transform 1 0 1025 0 1 51517
box -104 -632 104 632
use M3_M2_CDNS_6903358316569  M3_M2_CDNS_6903358316569_1
timestamp 1713338890
transform 1 0 1026 0 1 62699
box -104 -632 104 632
use M3_M2_CDNS_6903358316570  M3_M2_CDNS_6903358316570_0
timestamp 1713338890
transform 1 0 1818 0 1 49901
box -100 -596 100 596
use M3_M2_CDNS_6903358316570  M3_M2_CDNS_6903358316570_1
timestamp 1713338890
transform 1 0 182 0 1 49901
box -100 -596 100 596
use M3_M2_CDNS_6903358316570  M3_M2_CDNS_6903358316570_2
timestamp 1713338890
transform 1 0 182 0 1 64300
box -100 -596 100 596
use M3_M2_CDNS_6903358316570  M3_M2_CDNS_6903358316570_3
timestamp 1713338890
transform 1 0 1818 0 1 64300
box -100 -596 100 596
use POLY_SUB_FILL_1  POLY_SUB_FILL_1_0
array 0 0 0 0 15 3412
timestamp 1713338890
transform -1 0 2287 0 1 14392
box 310 -127 2260 3485
<< labels >>
rlabel metal3 s 1011 67458 1011 67458 4 DVDD
port 1 nsew
rlabel metal3 s 1011 59623 1011 59623 4 DVDD
port 1 nsew
rlabel metal3 s 1011 56423 1011 56423 4 DVDD
port 1 nsew
rlabel metal3 s 1011 54658 1011 54658 4 DVDD
port 1 nsew
rlabel metal3 s 1011 53223 1011 53223 4 DVDD
port 1 nsew
rlabel metal3 s 1011 44368 1011 44368 4 DVDD
port 1 nsew
rlabel metal3 s 1011 41977 1011 41977 4 DVDD
port 1 nsew
rlabel metal3 s 1011 37959 1011 37959 4 DVDD
port 1 nsew
rlabel metal3 s 1011 34723 1011 34723 4 DVDD
port 1 nsew
rlabel metal3 s 1011 31609 1011 31609 4 DVDD
port 1 nsew
rlabel metal3 s 1011 28394 1011 28394 4 DVDD
port 1 nsew
rlabel metal3 s 1011 24284 1011 24284 4 DVDD
port 1 nsew
rlabel metal3 s 1011 18921 1011 18921 4 DVSS
port 2 nsew
rlabel metal3 s 1011 15750 1011 15750 4 DVSS
port 2 nsew
rlabel metal3 s 1011 21907 1011 21907 4 DVSS
port 2 nsew
rlabel metal3 s 1011 26100 1011 26100 4 DVSS
port 2 nsew
rlabel metal3 s 1011 40342 1011 40342 4 DVSS
port 2 nsew
rlabel metal3 s 1011 47595 1011 47595 4 DVSS
port 2 nsew
rlabel metal3 s 1011 57858 1011 57858 4 DVSS
port 2 nsew
rlabel metal3 s 1011 61058 1011 61058 4 DVSS
port 2 nsew
rlabel metal3 s 1011 66023 1011 66023 4 DVSS
port 2 nsew
rlabel metal3 s 1011 69049 1011 69049 4 DVSS
port 2 nsew
rlabel metal3 s 1011 51458 1011 51458 4 VDD
port 3 nsew
rlabel metal3 s 1011 62823 1011 62823 4 VDD
port 3 nsew
rlabel metal3 s 1011 64258 1011 64258 4 VSS
port 4 nsew
rlabel metal3 s 1011 50023 1011 50023 4 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2000 70000
<< end >>
