magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1097 -1019 1097 1019
<< metal1 >>
rect -97 13 97 19
rect -97 -13 -91 13
rect 91 -13 97 13
rect -97 -19 97 -13
<< via1 >>
rect -91 -13 91 13
<< metal2 >>
rect -97 13 97 19
rect -97 -13 -91 13
rect 91 -13 97 13
rect -97 -19 97 -13
<< end >>
