magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6087 -2045 6087 2045
<< psubdiff >>
rect -4087 23 4087 45
rect -4087 -23 -4065 23
rect 4065 -23 4087 23
rect -4087 -45 4087 -23
<< psubdiffcont >>
rect -4065 -23 4065 23
<< metal1 >>
rect -4076 23 4076 34
rect -4076 -23 -4065 23
rect 4065 -23 4076 23
rect -4076 -34 4076 -23
<< end >>
