* NGSPICE file created from PLL_TOP_MUX_2_flat.ext - technology: gf180mcuC

.subckt pex_PLL_TOP_MUX_2 UP_INPUT VDD DN_INPUT VSS PRE_SCALAR UP F_IN DN ITAIL DIV_OUT S1 ITAIL1 VCTRL_IN S6 VCTRL2 S2 OUT
+ S3 S4 OUTB LF_OFFCHIP S5
X0 a_42928_8770.t1 a_43228_8148.t1 VDD.t376 ppolyf_u r_width=1.1u r_length=2.6u
X1 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.IN.t17 VSS.t577 VSS.t576 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.5u
X2 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t18 VDD.t344 VDD.t343 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X3 PFD_T2_0.FDIV a_20903_8375.t6 DIV_OUT.t4 VDD.t430 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X4 OUTB a_50528_5246.t24 VDD.t648 VDD.t603 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X5 CP_1_0.VCTRL ITAIL.t16 a_32731_10265.t7 VDD.t428 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X6 VSS.t516 VSS.t515 VSS.t516 VSS.t211 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X7 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t31 VSS.t307 VSS.t306 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X8 ITAIL ITAIL.t14 VDD.t427 VDD.t426 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X9 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t32 VDD.t614 VDD.t402 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X10 VSS VCTRL2.t1 a_25706_n567.t53 VSS.t724 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X11 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t31 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t3 VSS.t536 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X12 VSS a_50630_6066.t6 a_50528_5246.t7 VSS.t258 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X13 VSS a_50708_569.t24 OUT.t31 VSS.t298 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X14 VDD S1.t0 A_MUX_1.Tr_Gate_1.CLK.t11 VDD.t769 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X15 a_43528_12082.t0 a_43828_11460.t0 VDD.t133 ppolyf_u r_width=1.1u r_length=2.6u
X16 VDD a_32467_10269.t6 a_32731_10265.t2 VDD.t1 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X17 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t31 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t10 VDD.t383 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X18 RES_74k_1.M.t1 VSS.t705 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X19 VDD S2.t0 A_MUX_3.Tr_Gate_1.CLK.t11 VDD.t763 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X20 VSS PFD_T2_0.Buffer_V_2_0.IN.t11 a_25557_8739.t0 VSS.t325 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X21 VSS a_50528_5246.t25 OUTB.t31 VSS.t33 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X22 VSS.t514 VSS.t513 VSS.t514 VSS.t214 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X23 VSS.t512 VSS.t510 VSS.t512 VSS.t511 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X24 RES_74k_1.P.t45 RES_74k_1.P.t46 VDD.t272 ppolyf_u r_width=1.1u r_length=2.6u
X25 OUTB a_50528_5246.t26 VDD.t649 VDD.t213 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X26 CP_1_0.VCTRL A_MUX_0.Tr_Gate_1.CLK.t12 VCO_DFF_C_0.VCTRL.t15 VSS.t765 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X27 RES_74k_1.M.t1 VSS.t704 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X28 VDD a_22967_8787.t4 PFD_T2_0.INV_mag_1.IN.t4 VDD.t182 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X29 RES_74k_1.P.t81 RES_74k_1.P.t82 VDD.t376 ppolyf_u r_width=1.1u r_length=2.6u
X30 VSS VCTRL2.t3 a_34443_2598.t49 VSS.t729 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X31 VSS a_50810_1389.t6 a_50708_569.t5 VSS.t50 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X32 PRE_SCALAR A_MUX_1.Tr_Gate_1.CLK.t12 PFD_T2_0.FIN.t10 VSS.t343 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X33 VSS S6.t0 A_MUX_2.Tr_Gate_1.CLK.t3 VSS.t85 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X34 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t12 VCO_DFF_C_0.VCO_C_0.OUTB.t3 VSS.t912 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X35 RES_74k_1.M.t1 VSS.t703 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X36 VSS a_18508_8715.t6 PFD_T2_0.FDIV.t1 VDD.t68 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X37 RES_74k_1.M.t2 VSS.t778 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X38 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.OUT.t6 VSS.t144 VSS.t143 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X39 VDD a_22967_8787.t5 PFD_T2_0.INV_mag_1.IN.t10 VDD.t832 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X40 A_MUX_2.Tr_Gate_1.CLK S6.t1 VDD.t207 VDD.t206 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X41 a_43828_11254.t1 a_43528_10632.t0 VDD.t133 ppolyf_u r_width=1.1u r_length=2.6u
X42 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL.t16 VDD.t859 VDD.t672 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X43 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t16 VCO_DFF_C_0.OUT VSS.t249 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X44 VSS PFD_T2_0.INV_mag_1.OUT.t3 a_22879_10704.t1 VSS.t528 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X45 VDD a_32467_10269.t7 a_32731_10265.t1 VDD.t1 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X46 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.IN.t19 VDD.t342 VDD.t341 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X47 OUTB a_50528_5246.t27 VDD.t650 VDD.t598 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X48 VDD.t996 VDD.t994 VDD.t996 VDD.t995 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X49 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t31 VDD.t152 VDD.t93 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X50 VDD.t993 VDD.t992 VDD.t993 VDD.t934 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X51 RES_74k_1.M.t1 VSS.t702 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X52 RES_74k_1.M.t1 VSS.t701 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X53 OUTB a_50528_5246.t28 VDD.t651 VDD.t482 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X54 VSS.t509 VSS.t508 VSS.t509 VSS.t424 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X55 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t12 a_34443_2598.t10 VSS.t172 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X56 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t32 VDD.t510 VDD.t402 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X57 VDD a_50810_1389.t8 a_50708_569.t1 VDD.t32 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X58 RES_74k_1.M.t1 VSS.t700 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X59 OUT a_50708_569.t25 VDD.t607 VDD.t74 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X60 RES_74k_1.M.t2 VSS.t777 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X61 VSS UP_OUT.t16 a_32939_9624.t4 VSS.t918 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X62 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCTRL.t17 VDD.t860 VDD.t666 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X63 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t33 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t20 VDD.t383 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X64 VDD.t991 VDD.t989 VDD.t991 VDD.t990 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X65 OUT a_50708_569.t26 VDD.t608 VDD.t38 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X66 RES_74k_1.M.t1 VSS.t699 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X67 VSS a_50528_5246.t29 OUTB.t30 VSS.t292 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X68 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t12 a_34443_2598.t0 VSS.t5 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X69 OUT a_50708_569.t27 VDD.t609 VDD.t76 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X70 UP_OUT A_MUX_3.Tr_Gate_1.CLK.t12 UP1.t3 VSS.t245 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X71 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t34 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t19 VDD.t519 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X72 VSS VCTRL2.t6 a_34443_2598.t47 VSS.t736 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X73 VSS.t507 VSS.t506 VSS.t507 VSS.t499 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X74 RES_74k_1.M.t1 VSS.t698 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X75 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t12 a_44716_n517.t1 VSS.t148 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X76 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t12 VSS.t223 VSS.t222 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X77 VSS a_50708_569.t28 OUT.t30 VSS.t301 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X78 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t13 VCO_DFF_C_0.VCO_C_0.OUT.t11 VDD.t503 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X79 RES_74k_1.M.t1 VSS.t697 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X80 RES_74k_1.P.t59 RES_74k_1.P.t60 VDD.t31 ppolyf_u r_width=1.1u r_length=2.6u
X81 VSS.t505 VSS.t503 VSS.t505 VSS.t504 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X82 A_MUX_2.Tr_Gate_1.CLK S6.t2 VSS.t946 VSS.t945 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X83 VSS.t502 VSS.t501 VSS.t502 VSS.t435 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X84 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t32 VDD.t713 VDD.t180 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X85 RES_74k_1.M.t1 VSS.t696 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X86 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCTRL.t18 VDD.t861 VDD.t669 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X87 RES_74k_1.M.t1 VSS.t695 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X88 a_44728_10426.t1 a_44428_9804.t1 VDD.t31 ppolyf_u r_width=1.1u r_length=2.6u
X89 VDD a_50528_5246.t30 OUTB.t91 VDD.t464 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X90 OUTB a_50528_5246.t31 VDD.t654 VDD.t603 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X91 VSS A_MUX_3.Tr_Gate_1.CLK.t13 a_27480_10186.t1 VSS.t71 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X92 VDD S4.t0 A_MUX_0.Tr_Gate_1.CLK.t4 VDD.t281 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X93 a_42628_9598.t1 a_42928_8976.t1 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X94 VSS.t500 VSS.t498 VSS.t500 VSS.t499 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X95 a_44728_12082.t0 a_44428_11460.t0 VDD.t31 ppolyf_u r_width=1.1u r_length=2.6u
X96 OUTB a_50528_5246.t32 VDD.t655 VDD.t605 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X97 VDD VCO_DFF_C_0.OUTB.t21 a_50630_6066.t2 VDD.t467 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X98 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t33 VSS.t228 VSS.t227 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X99 RES_74k_1.M.t3 VSS.t336 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X100 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB.t12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t15 VSS.t28 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X101 VDD a_50708_569.t29 OUT.t92 VDD.t223 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X102 OUTB a_50528_5246.t33 VSS.t322 VSS.t169 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X103 RES_74k_1.M.t1 VSS.t694 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X104 OUTB a_50528_5246.t34 VDD.t656 VDD.t488 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X105 RES_74k_1.M.t1 VSS.t693 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X106 RES_74k_1.M.t1 VSS.t692 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X107 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.IN.t18 VDD.t1088 VDD.t341 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X108 VDD a_50810_1389.t10 a_50708_569.t3 VDD.t35 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X109 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t13 a_25706_n567.t11 VSS.t17 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X110 a_44428_11254.t1 a_44728_10632.t0 VDD.t31 ppolyf_u r_width=1.1u r_length=2.6u
X111 VSS VCO_DFF_C_0.OUT.t7 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t6 VSS.t249 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X112 VSS VCTRL2.t8 a_25706_n567.t50 VSS.t740 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X113 RES_74k_1.M.t3 VSS.t335 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X114 VSS PFD_T2_0.INV_mag_0.IN.t19 a_23836_10693.t2 VSS.t989 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X115 a_45928_10426.t1 a_46228_9804.t0 VDD.t131 ppolyf_u r_width=1.1u r_length=2.6u
X116 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t33 VDD.t714 VDD.t319 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X117 RES_74k_1.M.t1 VSS.t691 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X118 VDD a_50528_5246.t35 OUTB.t87 VDD.t494 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X119 A_MUX_1.Tr_Gate_1.CLK S1.t1 VSS.t988 VSS.t987 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X120 a_44428_9598.t0 a_44128_8976.t0 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X121 VDD S4.t1 a_42763_5679.t5 VDD.t367 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X122 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t13 VDD.t778 VDD.t753 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X123 RES_74k_1.M.t2 VSS.t776 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X124 VSS.t497 VSS.t496 VSS.t497 VSS.t46 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X125 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t13 VSS.t30 VSS.t29 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X126 VDD a_50708_569.t30 OUT.t91 VDD.t32 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X127 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t35 VDD.t619 VDD.t386 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X128 RES_74k_1.M.t1 VSS.t690 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X129 a_45928_8770.t1 a_45628_8148.t0 VDD.t243 ppolyf_u r_width=1.1u r_length=2.6u
X130 RES_74k_1.M.t1 VSS.t689 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X131 VCO_DFF_C_0.OUTB a_41879_1284.t6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t9 VDD.t49 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X132 a_42628_8770.t1 a_42628_8148.t1 VDD.t269 ppolyf_u r_width=1.1u r_length=2.6u
X133 OUTB a_50528_5246.t36 VSS.t324 VSS.t323 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X134 CP_1_0.VCTRL ITAIL.t19 a_32731_10265.t6 VDD.t426 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X135 VSS.t495 VSS.t494 VSS.t495 VSS.t173 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X136 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t14 a_25706_n567.t12 VSS.t78 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X137 RES_74k_1.P.t17 RES_74k_1.P.t18 VDD.t22 ppolyf_u r_width=1.1u r_length=2.6u
X138 RES_74k_1.M.t1 VSS.t688 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X139 OUT a_50708_569.t31 VSS.t305 VSS.t304 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X140 VSS VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t14 VCO_DFF_C_0.VCO_C_0.OUT.t2 VSS.t224 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X141 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t34 VDD.t715 VDD.t93 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X142 VDD A_MUX_2.Tr_Gate_1.CLK.t12 a_20903_8375.t4 VDD.t709 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X143 VDD.t988 VDD.t987 VDD.t988 VDD.t958 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X144 VSS VCTRL2.t9 a_25706_n567.t49 VSS.t740 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X145 RES_74k_1.M.t1 VSS.t687 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X146 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t20 VDD.t328 VDD.t327 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X147 RES_74k_1.P.t79 RES_74k_1.P.t80 VDD.t243 ppolyf_u r_width=1.1u r_length=2.6u
X148 VSS VCO_DFF_C_0.OUT.t8 VCO_DFF_C_0.OUTB.t8 VSS.t252 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X149 A_MUX_6.Tr_Gate_1.CLK S5.t0 VDD.t271 VDD.t270 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X150 DN_OUT A_MUX_4.Tr_Gate_1.CLK.t14 DN1.t3 VSS.t121 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X151 RES_74k_1.P.t85 RES_74k_1.P.t86 VDD.t269 ppolyf_u r_width=1.1u r_length=2.6u
X152 VDD.t986 VDD.t985 VDD.t986 VDD.t666 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X153 PFD_T2_0.INV_mag_1.IN a_22967_8787.t6 VDD.t24 VDD.t23 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X154 A_MUX_1.Tr_Gate_1.CLK S1.t2 VDD.t774 VDD.t773 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X155 VDD a_50528_5246.t37 OUTB.t86 VDD.t464 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X156 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t35 VDD.t716 VDD.t174 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X157 VDD S2.t1 A_MUX_3.Tr_Gate_1.CLK.t10 VDD.t69 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X158 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t36 VDD.t717 VDD.t301 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X159 VDD A_MUX_0.Tr_Gate_1.CLK.t13 a_45158_5339.t5 VDD.t333 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X160 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t34 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t12 VDD.t398 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X161 a_45328_12082.t1 a_45628_11460.t0 VDD.t22 ppolyf_u r_width=1.1u r_length=2.6u
X162 VDD a_50528_5246.t38 OUTB.t85 VDD.t431 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X163 PRE_SCALAR A_MUX_1.Tr_Gate_1.CLK.t13 PFD_T2_0.FIN.t9 VSS.t344 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X164 VDD a_50528_5246.t39 OUTB.t84 VDD.t467 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X165 F_IN S1.t3 PFD_T2_0.FIN.t15 VSS.t562 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X166 A_MUX_4.Tr_Gate_1.CLK S3.t0 VDD.t841 VDD.t284 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X167 VDD a_50708_569.t32 OUT.t90 VDD.t223 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X168 A_MUX_4.Tr_Gate_1.CLK S3.t1 VSS.t761 VSS.t760 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X169 a_44128_8770.t1 a_43828_8148.t1 VDD.t242 ppolyf_u r_width=1.1u r_length=2.6u
X170 VDD.t984 VDD.t982 VDD.t984 VDD.t983 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X171 VDD a_50708_569.t33 OUT.t89 VDD.t807 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X172 VDD S1.t4 A_MUX_1.Tr_Gate_1.CLK.t9 VDD.t775 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X173 PFD_T2_0.FIN a_20945_11785.t6 PRE_SCALAR.t1 VDD.t163 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X174 VDD a_50528_5246.t40 OUTB.t83 VDD.t434 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X175 VSS VCTRL2.t10 a_25706_n567.t48 VSS.t745 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X176 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t32 VSS.t55 VSS.t54 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X177 RES_74k_1.P.t97 VSS.t281 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X178 RES_74k_1.M.t1 VSS.t686 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X179 CP_1_0.VCTRL ITAIL1.t8 a_32939_9624.t5 VSS.t330 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X180 VDD A_MUX_4.Tr_Gate_1.CLK.t15 a_27423_7180.t4 VDD.t540 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X181 RES_74k_1.M.t1 VSS.t685 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X182 VDD a_50708_569.t34 OUT.t88 VDD.t35 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X183 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t36 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t11 VDD.t390 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X184 a_45628_11254.t0 a_45328_10632.t0 VDD.t22 ppolyf_u r_width=1.1u r_length=2.6u
X185 VDD A_MUX_0.Tr_Gate_1.CLK.t14 a_45158_5339.t4 VDD.t334 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X186 VSS.t493 VSS.t492 VSS.t493 VSS.t103 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X187 PFD_T2_0.FIN a_20945_11785.t7 PRE_SCALAR.t2 VDD.t164 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X188 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t13 a_34443_2598.t9 VSS.t931 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X189 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB.t15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t14 VSS.t15 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X190 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t16 a_41879_1284.t3 VDD.t49 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X191 VDD a_50708_569.t35 OUT.t87 VDD.t208 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X192 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t33 VDD.t89 VDD.t88 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X193 VDD.t981 VDD.t980 VDD.t981 VDD.t934 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X194 RES_74k_1.M.t1 VSS.t684 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X195 VDD VCO_DFF_C_0.OUT.t9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t15 VDD.t9 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X196 VDD a_22966_11778.t4 PFD_T2_0.INV_mag_0.IN.t6 VDD.t897 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X197 RES_74k_1.P.t75 RES_74k_1.P.t76 VDD.t242 ppolyf_u r_width=1.1u r_length=2.6u
X198 VSS VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t34 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t2 VSS.t56 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X199 RES_74k_1.M.t1 VSS.t683 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X200 VSS S1.t5 A_MUX_1.Tr_Gate_1.CLK.t2 VSS.t563 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X201 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t37 VDD.t622 VDD.t396 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X202 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t35 VDD.t514 VDD.t513 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X203 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t37 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t9 VDD.t322 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X204 RES_74k_1.M.t1 VSS.t682 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X205 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t38 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t17 VDD.t398 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X206 OUT a_50708_569.t36 VDD.t852 VDD.t211 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X207 VSS a_50528_5246.t41 OUTB.t27 VSS.t205 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X208 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t38 VSS.t540 VSS.t539 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X209 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t11 VDD.t185 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X210 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t16 VDD.t576 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X211 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t14 VSS.t579 VSS.t578 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X212 RES_74k_1.M.t1 VSS.t681 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X213 VSS.t491 VSS.t489 VSS.t491 VSS.t490 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X214 VSS.t488 VSS.t487 VSS.t488 VSS.t178 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X215 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t15 VCO_DFF_C_0.VCO_C_0.OUTB.t10 VDD.t755 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X216 RES_74k_1.M.t1 VSS.t680 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X217 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t17 VCO_DFF_C_0.OUT VDD.t750 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X218 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t17 VDD.t200 VDD.t188 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X219 VSS ITAIL1.t6 ITAIL1.t7 VSS.t899 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X220 VSS VCTRL2.t12 a_25706_n567.t47 VSS.t724 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X221 VSS a_50528_5246.t42 OUTB.t26 VSS.t208 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X222 VDD.t979 VDD.t977 VDD.t979 VDD.t978 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X223 RES_74k_1.P.t93 RES_74k_1.P.t94 VDD.t269 ppolyf_u r_width=1.1u r_length=2.6u
X224 VSS VCTRL2.t13 a_25706_n567.t46 VSS.t724 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X225 UP_OUT a_27480_10186.t6 UP1.t4 VDD.t40 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X226 RES_74k_1.P.t77 RES_74k_1.P.t78 VDD.t272 ppolyf_u r_width=1.1u r_length=2.6u
X227 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t35 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t0 VDD.t90 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X228 VSS VCO_DFF_C_0.OUT.t10 a_50810_1389.t3 VSS.t580 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X229 DN_OUT a_29818_7696.t6 DN_INPUT.t7 VDD.t562 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X230 VSS a_50708_569.t37 OUT.t28 VSS.t464 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X231 RES_74k_1.P A_MUX_6.Tr_Gate_1.CLK.t13 CP_1_0.VCTRL.t26 VSS.t278 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X232 VDD S5.t2 A_MUX_6.Tr_Gate_1.CLK.t10 VDD.t273 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X233 VDD S6.t3 a_18508_8715.t5 VDD.t68 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X234 RES_74k_1.M.t1 VSS.t679 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X235 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t36 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t13 VDD.t393 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X236 RES_74k_1.M.t1 VSS.t678 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X237 VSS a_22967_8787.t7 a_22881_9554.t1 VSS.t6 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X238 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t39 VDD.t720 VDD.t180 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X239 VDD S5.t3 A_MUX_6.Tr_Gate_1.CLK.t9 VDD.t276 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X240 VDD a_25557_8739.t3 DN1.t10 VDD.t1079 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X241 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t37 VDD.t518 VDD.t517 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X242 RES_74k_1.M.t0 a_42628_11460.t1 VDD.t269 ppolyf_u r_width=1.1u r_length=2.6u
X243 VDD VCO_DFF_C_0.OUT.t11 VCO_DFF_C_0.OUTB.t10 VDD.t6 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X244 a_46528_12082.t1 a_46228_11460.t1 VDD.t272 ppolyf_u r_width=1.1u r_length=2.6u
X245 OUTB a_50528_5246.t43 VDD.t479 VDD.t442 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X246 VSS.t486 VSS.t485 VSS.t486 VSS.t368 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X247 UP_OUT a_29875_10702.t6 UP_INPUT.t3 VDD.t72 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X248 PFD_T2_0.INV_mag_0.IN a_22966_11778.t6 VDD.t901 VDD.t900 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X249 DN1 a_27423_7180.t6 DN_OUT.t1 VDD.t130 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X250 RES_74k_1.M.t1 VSS.t677 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X251 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t16 VDD.t674 VDD.t52 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X252 a_45328_10426.t0 a_45628_9804.t1 VDD.t22 ppolyf_u r_width=1.1u r_length=2.6u
X253 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t15 VDD.t123 VDD.t122 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X254 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t36 VDD.t94 VDD.t93 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X255 RES_74k_1.P.t65 RES_74k_1.P.t66 VDD.t21 ppolyf_u r_width=1.1u r_length=2.6u
X256 OUTB a_50528_5246.t44 VDD.t480 VDD.t444 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X257 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t20 VDD.t1089 VDD.t900 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X258 VDD a_22967_8787.t8 PFD_T2_0.INV_mag_1.IN.t15 VDD.t294 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X259 a_43828_9598.t1 a_43528_8976.t1 VDD.t133 ppolyf_u r_width=1.1u r_length=2.6u
X260 VCO_DFF_C_0.VCTRL S4.t3 VCTRL_IN.t7 VSS.t150 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X261 VSS a_50630_6066.t9 a_50528_5246.t16 VSS.t197 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X262 VCTRL_IN a_42763_5679.t6 VCO_DFF_C_0.VCTRL.t8 VDD.t367 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X263 OUT a_50708_569.t38 VDD.t853 VDD.t38 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X264 A_MUX_4.Tr_Gate_1.CLK S3.t2 VDD.t842 VDD.t286 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X265 VSS VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t37 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t1 VSS.t59 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X266 a_42628_11254.t1 a_42628_10426.t1 VDD.t269 ppolyf_u r_width=1.1u r_length=2.6u
X267 a_46228_11254.t1 a_46528_10632.t1 VDD.t272 ppolyf_u r_width=1.1u r_length=2.6u
X268 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t38 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t2 VDD.t95 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X269 RES_74k_1.M.t1 VSS.t676 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X270 OUT a_50708_569.t39 VDD.t855 VDD.t854 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X271 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t14 a_34443_2598.t52 VSS.t931 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X272 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t39 VDD.t99 VDD.t98 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X273 RES_74k_1.M.t1 VSS.t675 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X274 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t5 VSS.t142 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X275 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_0.OUT.t6 VSS.t938 VSS.t556 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X276 VSS A_MUX_4.Tr_Gate_1.CLK.t16 a_27423_7180.t0 VSS.t948 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X277 VSS a_50528_5246.t45 OUTB.t25 VSS.t211 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X278 VSS.t484 VSS.t482 VSS.t484 VSS.t483 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X279 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t39 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t16 VDD.t519 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X280 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t16 VDD.t125 VDD.t124 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X281 A_MUX_3.Tr_Gate_1.CLK S2.t3 VSS.t42 VSS.t41 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X282 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t40 VSS.t308 VSS.t227 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X283 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t18 a_25706_n567.t8 VSS.t78 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X284 OUT a_50708_569.t40 VDD.t856 VDD.t810 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X285 A_MUX_6.Tr_Gate_1.CLK S5.t4 VSS.t274 VSS.t273 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X286 VSS a_50630_6066.t10 a_50528_5246.t0 VSS.t33 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X287 OUTB a_50528_5246.t46 VSS.t215 VSS.t214 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X288 RES_74k_1.M.t1 VSS.t674 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X289 OUTB a_50528_5246.t47 VDD.t481 VDD.t213 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X290 DIV_OUT a_20903_8375.t7 PFD_T2_0.FDIV.t9 VDD.t709 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X291 RES_74k_1.P.t73 RES_74k_1.P.t74 VDD.t361 ppolyf_u r_width=1.1u r_length=2.6u
X292 VSS.t481 VSS.t479 VSS.t481 VSS.t480 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X293 RES_74k_1.M.t1 VSS.t673 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X294 VSS.t478 VSS.t477 VSS.t478 VSS.t181 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X295 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t40 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t10 VDD.t100 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X296 A_MUX_6.Tr_Gate_1.CLK S5.t5 VDD.t584 VDD.t555 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X297 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_n517.t6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t18 VDD.t192 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X298 OUT a_50708_569.t41 VSS.t764 VSS.t365 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X299 CP_1_0.VCTRL a_39080_11413.t6 RES_74k_1.P.t25 VDD.t411 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X300 a_45028_9598.t1 a_45328_8976.t1 VDD.t217 ppolyf_u r_width=1.1u r_length=2.6u
X301 VSS VCTRL2.t16 a_34443_2598.t44 VSS.t757 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X302 RES_74k_1.P.t95 RES_74k_1.P.t96 VDD.t262 ppolyf_u r_width=1.1u r_length=2.6u
X303 CP_1_0.VCTRL a_45158_5339.t6 VCO_DFF_C_0.VCTRL.t1 VDD.t333 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X304 OUTB a_50528_5246.t48 VSS.t217 VSS.t216 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X305 VSS VCTRL2.t18 a_34443_2598.t43 VSS.t729 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X306 CP_1_0.VCTRL a_39080_11413.t7 RES_74k_1.P.t26 VDD.t412 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X307 RES_74k_1.M.t1 VSS.t672 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X308 VDD PFD_T2_0.FDIV.t17 a_22967_8787.t0 VDD.t294 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X309 DIV_OUT A_MUX_2.Tr_Gate_1.CLK.t14 PFD_T2_0.FDIV.t3 VSS.t95 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X310 a_46528_8770.t1 RES_74k_1.P.t90 VDD.t109 ppolyf_u r_width=1.1u r_length=2.6u
X311 VDD a_50630_6066.t11 a_50528_5246.t18 VDD.t494 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X312 OUTB a_50528_5246.t49 VDD.t483 VDD.t482 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X313 VDD VCO_DFF_C_0.OUT.t12 a_50810_1389.t4 VDD.t807 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X314 OUT a_50708_569.t42 VSS.t843 VSS.t456 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X315 PFD_T2_0.FDIV a_18508_8715.t7 VSS.t39 VDD.t67 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X316 a_43528_8770.t1 a_43228_8148.t0 VDD.t262 ppolyf_u r_width=1.1u r_length=2.6u
X317 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t38 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t14 VDD.t519 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X318 RES_74k_1.M.t1 VSS.t671 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X319 RES_74k_1.M.t1 VSS.t670 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X320 VDD S4.t4 A_MUX_0.Tr_Gate_1.CLK.t5 VDD.t281 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X321 VDD S6.t4 A_MUX_2.Tr_Gate_1.CLK.t10 VDD.t891 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X322 RES_74k_1.M.t1 VSS.t669 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X323 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t19 a_44716_1837.t5 VDD.t201 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X324 VDD a_50810_1389.t13 a_50708_569.t12 VDD.t208 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X325 VDD.t976 VDD.t975 VDD.t976 VDD.t949 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X326 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.OUT.t5 VSS.t559 VSS.t558 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X327 VDD ITAIL.t12 ITAIL.t13 VDD.t423 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X328 a_43528_12082.t1 a_43228_11460.t1 VDD.t262 ppolyf_u r_width=1.1u r_length=2.6u
X329 CP_1_0.VCTRL a_45158_5339.t7 VCO_DFF_C_0.VCTRL.t2 VDD.t334 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X330 VSS.t476 VSS.t474 VSS.t476 VSS.t475 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X331 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t15 a_34443_2598.t53 VSS.t932 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X332 LF_OFFCHIP a_36685_10901.t6 CP_1_0.VCTRL.t10 VDD.t422 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X333 DN_OUT S3.t4 DN_INPUT.t3 VSS.t131 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X334 VDD a_50528_5246.t50 OUTB.t78 VDD.t449 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X335 RES_74k_1.M.t1 VSS.t668 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X336 OUT a_50708_569.t43 VDD.t922 VDD.t244 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X337 RES_74k_1.P.t61 RES_74k_1.P.t62 VDD.t109 ppolyf_u r_width=1.1u r_length=2.6u
X338 VSS VCTRL2.t21 a_34443_2598.t41 VSS.t729 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X339 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t40 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t12 VDD.t90 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X340 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t21 a_23836_10693.t4 VSS.t992 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X341 RES_74k_1.P.t19 RES_74k_1.P.t20 VDD.t262 ppolyf_u r_width=1.1u r_length=2.6u
X342 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t41 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t11 VDD.t171 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X343 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_n196.t6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t3 VDD.t44 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X344 RES_74k_1.M.t1 VSS.t667 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X345 CP_1_0.VCTRL A_MUX_0.Tr_Gate_1.CLK.t16 VCO_DFF_C_0.VCTRL.t14 VSS.t911 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X346 VSS.t473 VSS.t472 VSS.t473 VSS.t350 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X347 VSS S4.t5 A_MUX_0.Tr_Gate_1.CLK.t6 VSS.t65 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X348 VSS.t471 VSS.t470 VSS.t471 VSS.t304 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X349 a_43228_11254.t1 a_43528_10632.t1 VDD.t262 ppolyf_u r_width=1.1u r_length=2.6u
X350 RES_74k_1.M.t1 VSS.t666 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X351 VSS PFD_T2_0.INV_mag_1.IN.t22 a_23837_9553.t5 VSS.t568 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X352 a_44728_8770.t1 a_45028_8148.t1 VDD.t154 ppolyf_u r_width=1.1u r_length=2.6u
X353 OUTB a_50528_5246.t51 VSS.t218 VSS.t185 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X354 RES_74k_1.M.t1 VSS.t665 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X355 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t20 a_44716_n517.t3 VDD.t194 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X356 DN_INPUT S3.t5 DN_OUT.t4 VSS.t133 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X357 VSS.t469 VSS.t468 VSS.t469 VSS.t360 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X358 PFD_T2_0.FIN a_18550_11273.t6 F_IN.t0 VDD.t329 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X359 VDD a_50528_5246.t52 OUTB.t77 VDD.t431 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X360 VDD S4.t6 A_MUX_0.Tr_Gate_1.CLK.t7 VDD.t110 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X361 RES_74k_1.M.t1 VSS.t664 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X362 VCO_DFF_C_0.VCTRL a_42763_5679.t7 VCTRL_IN.t2 VDD.t370 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X363 VDD.t974 VDD.t972 VDD.t974 VDD.t973 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X364 A_MUX_3.Tr_Gate_1.CLK S2.t4 VDD.t889 VDD.t888 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X365 VDD a_50630_6066.t13 a_50528_5246.t10 VDD.t434 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X366 OUTB a_50528_5246.t53 VDD.t489 VDD.t488 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X367 VDD VCO_DFF_C_0.VCTRL.t19 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t25 VDD.t666 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X368 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t42 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t10 VDD.t90 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X369 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t19 VSS.t20 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X370 VSS S3.t6 A_MUX_4.Tr_Gate_1.CLK.t2 VSS.t155 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X371 RES_74k_1.P.t63 RES_74k_1.P.t64 VDD.t154 ppolyf_u r_width=1.1u r_length=2.6u
X372 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t41 VDD.t104 VDD.t103 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X373 OUTB a_50528_5246.t54 VSS.t219 VSS.t187 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X374 VSS.t467 VSS.t466 VSS.t467 VSS.t189 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X375 VDD a_50528_5246.t55 OUTB.t75 VDD.t446 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X376 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN a_44716_n517.t7 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t15 VDD.t194 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X377 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t16 a_34443_2598.t54 VSS.t847 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X378 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t42 VDD.t228 VDD.t174 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X379 VSS VCTRL2.t22 a_25706_n567.t42 VSS.t797 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X380 VSS a_50708_569.t44 OUT.t25 VSS.t357 nfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X381 OUT a_50708_569.t45 VSS.t846 VSS.t99 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X382 VDD.t971 VDD.t969 VDD.t971 VDD.t970 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X383 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t13 VSS.t22 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X384 RES_74k_1.P.t71 RES_74k_1.P.t72 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X385 VSS VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t39 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t2 VSS.t161 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X386 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t15 a_25706_n567.t13 VSS.t78 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X387 VDD a_50528_5246.t56 OUTB.t74 VDD.t106 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X388 RES_74k_1.M.t1 VSS.t663 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X389 VSS A_MUX_2.Tr_Gate_1.CLK.t16 a_20903_8375.t3 VSS.t96 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X390 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t43 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t8 VDD.t100 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X391 VSS a_50810_1389.t15 a_50708_569.t14 VSS.t90 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X392 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t21 a_41879_1284.t0 VSS.t110 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X393 PFD_T2_0.INV_mag_0.IN a_22966_11778.t7 VDD.t903 VDD.t902 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X394 VDD a_50528_5246.t57 OUTB.t73 VDD.t494 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X395 VDD a_50708_569.t46 OUT.t81 VDD.t807 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X396 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t40 VDD.t522 VDD.t388 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X397 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t43 VDD.t302 VDD.t301 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X398 VDD a_50528_5246.t58 OUTB.t72 VDD.t497 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X399 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t44 VSS.t107 VSS.t106 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X400 RES_74k_1.M.t1 VSS.t662 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X401 VDD a_50708_569.t47 OUT.t80 VDD.t246 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X402 PFD_T2_0.INV_mag_0.IN a_22966_11778.t8 VDD.t905 VDD.t904 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X403 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t22 VDD.t1090 VDD.t902 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X404 VSS VCTRL2.t24 a_34443_2598.t39 VSS.t779 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X405 OUT a_50708_569.t48 VDD.t927 VDD.t854 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X406 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t16 VDD.t781 VDD.t761 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X407 VDD a_50708_569.t49 OUT.t78 VDD.t208 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X408 a_44128_12082.t0 a_44428_11460.t1 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X409 VDD VCO_DFF_C_0.VCTRL.t20 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t30 VDD.t672 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X410 RES_74k_1.M.t1 VSS.t661 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X411 VSS.t465 VSS.t463 VSS.t465 VSS.t464 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X412 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t23 VDD.t1091 VDD.t904 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X413 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t23 a_25706_n567.t9 VSS.t78 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X414 RES_74k_1.M.t1 VSS.t660 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X415 VDD a_50708_569.t50 OUT.t77 VDD.t249 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X416 VDD A_MUX_3.Tr_Gate_1.CLK.t17 a_27480_10186.t3 VDD.t41 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X417 VSS.t462 VSS.t461 VSS.t462 VSS.t447 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X418 VDD a_32467_10269.t8 a_32731_10265.t0 VDD.t1 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X419 OUTB a_50528_5246.t59 VSS.t174 VSS.t173 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X420 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t44 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t9 VDD.t95 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X421 VSS VCO_DFF_C_0.VCO_C_0.OUTB.t24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t2 VSS.t82 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X422 OUT a_50708_569.t51 VDD.t932 VDD.t211 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X423 A_MUX_3.Tr_Gate_1.CLK S2.t6 VSS.t823 VSS.t822 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X424 VSS.t460 VSS.t458 VSS.t460 VSS.t459 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X425 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t22 a_44716_n517.t2 VDD.t201 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X426 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_1284.t7 VCO_DFF_C_0.OUTB.t14 VDD.t132 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X427 VSS S1.t6 a_18550_11273.t1 VSS.t562 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X428 UP1 a_25556_11637.t3 VDD.t156 VDD.t155 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X429 A_MUX_6.Tr_Gate_1.CLK S5.t6 VSS.t276 VSS.t275 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X430 a_44428_11254.t0 a_44128_10632.t1 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X431 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL.t21 VDD.t785 VDD.t784 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X432 RES_74k_1.M.t1 VSS.t659 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X433 VDD A_MUX_2.Tr_Gate_1.CLK.t17 a_20903_8375.t0 VDD.t85 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X434 a_46528_10426.t1 a_46228_9804.t1 VDD.t272 ppolyf_u r_width=1.1u r_length=2.6u
X435 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t45 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t8 VDD.t176 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X436 a_42928_10426.t0 a_43228_9804.t0 VDD.t376 ppolyf_u r_width=1.1u r_length=2.6u
X437 VSS VCO_DFF_C_0.OUT.t14 VCO_DFF_C_0.OUTB.t11 VSS.t583 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X438 VDD.t968 VDD.t967 VDD.t968 VDD.t672 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X439 a_44428_9598.t1 a_44728_8976.t1 VDD.t31 ppolyf_u r_width=1.1u r_length=2.6u
X440 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT a_41879_n196.t7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t4 VDD.t105 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X441 DN1 a_25557_8739.t4 VDD.t419 VDD.t418 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X442 DN_INPUT S3.t7 DN_OUT.t5 VSS.t158 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X443 VDD a_50528_5246.t60 OUTB.t71 VDD.t431 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X444 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t17 VDD.t543 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X445 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t41 VDD.t523 VDD.t386 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X446 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t46 VDD.t307 VDD.t98 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X447 VSS VCTRL2.t27 a_25706_n567.t40 VSS.t745 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X448 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t17 VSS.t340 VSS.t339 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X449 a_42928_8770.t0 a_42628_8148.t0 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X450 VDD a_50528_5246.t61 OUTB.t70 VDD.t434 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X451 RES_74k_1.M.t1 VSS.t658 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X452 VDD a_32467_10269.t9 a_32731_10265.t11 VDD.t1 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X453 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t7 VDD.t308 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X454 VSS a_50528_5246.t62 OUTB.t19 VSS.t175 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X455 VDD VCO_DFF_C_0.VCTRL.t22 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t22 VDD.t669 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X456 RES_74k_1.M.t1 VSS.t657 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X457 VDD a_50528_5246.t63 OUTB.t69 VDD.t437 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X458 CP_1_0.VCTRL S5.t7 LF_OFFCHIP.t7 VSS.t124 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X459 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t45 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t7 VDD.t166 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X460 VSS a_50708_569.t52 OUT.t23 VSS.t543 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X461 VDD S3.t8 A_MUX_4.Tr_Gate_1.CLK.t3 VDD.t377 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X462 RES_74k_1.P.t41 RES_74k_1.P.t42 VDD.t217 ppolyf_u r_width=1.1u r_length=2.6u
X463 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t15 a_34443_2598.t7 VSS.t847 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X464 VDD S5.t8 a_36685_10901.t5 VDD.t422 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X465 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t41 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t9 VDD.t404 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X466 RES_74k_1.M.t1 VSS.t656 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X467 LF_OFFCHIP a_36685_10901.t7 CP_1_0.VCTRL.t17 VDD.t548 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X468 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_44716_1837.t6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t0 VDD.t201 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X469 PFD_T2_0.FIN S1.t8 F_IN.t6 VSS.t561 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X470 RES_74k_1.P.t33 RES_74k_1.P.t34 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X471 RES_74k_1.M.t1 VSS.t655 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X472 VSS.t457 VSS.t455 VSS.t457 VSS.t456 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X473 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN.t24 a_23836_10693.t3 VSS.t989 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X474 VSS S2.t7 a_29875_10702.t0 VSS.t167 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X475 a_46228_9598.t1 a_45928_8976.t1 VDD.t131 ppolyf_u r_width=1.1u r_length=2.6u
X476 RES_74k_1.P A_MUX_6.Tr_Gate_1.CLK.t16 CP_1_0.VCTRL.t23 VSS.t68 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X477 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t42 VDD.t629 VDD.t407 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X478 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t42 VDD.t524 VDD.t517 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X479 VSS.t454 VSS.t453 VSS.t454 VSS.t368 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X480 VSS.t452 VSS.t451 VSS.t452 VSS.t350 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X481 OUTB a_50528_5246.t64 VDD.t441 VDD.t440 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X482 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t17 VCO_DFF_C_0.VCO_C_0.OUTB.t8 VDD.t758 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X483 RES_74k_1.M.t1 VSS.t654 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X484 VDD VCO_DFF_C_0.OUT.t15 VCO_DFF_C_0.OUTB.t12 VDD.t750 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X485 OUT a_50708_569.t53 VDD.t1016 VDD.t141 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X486 UP_INPUT S2.t8 UP_OUT.t11 VSS.t168 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X487 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t23 a_23837_9553.t1 VSS.t569 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X488 VSS.t450 VSS.t449 VSS.t450 VSS.t427 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X489 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t48 VDD.t311 VDD.t174 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X490 RES_74k_1.M.t1 VSS.t653 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X491 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.OUT.t16 VDD.t1107 VDD.t743 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X492 a_45328_12082.t0 a_45028_11460.t0 VDD.t217 ppolyf_u r_width=1.1u r_length=2.6u
X493 VSS a_50528_5246.t65 OUTB.t18 VSS.t178 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X494 OUT a_50708_569.t54 VDD.t1017 VDD.t854 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X495 PFD_T2_0.FDIV a_20903_8375.t8 DIV_OUT.t3 VDD.t215 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X496 a_44128_8770.t0 a_44428_8148.t0 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X497 RES_74k_1.M.t1 VSS.t652 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X498 VSS VCO_DFF_C_0.OUTB.t23 a_50630_6066.t4 VSS.t208 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X499 VSS.t448 VSS.t446 VSS.t448 VSS.t447 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X500 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t1 VSS.t136 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X501 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.OUT.t17 VDD.t1108 VDD.t748 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X502 VDD VCO_DFF_C_0.OUT.t18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t12 VDD.t745 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X503 OUT a_50708_569.t55 VSS.t893 VSS.t10 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X504 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t18 VCO_DFF_C_0.OUT VDD.t6 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X505 OUT a_50708_569.t56 VDD.t1018 VDD.t810 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X506 RES_74k_1.M.t1 VSS.t651 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X507 VSS.t445 VSS.t444 VSS.t445 VSS.t101 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X508 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t19 VDD.t1008 VDD.t19 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X509 VDD.t966 VDD.t964 VDD.t966 VDD.t965 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X510 VDD VCO_DFF_C_0.VCTRL.t23 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t27 VDD.t784 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X511 RES_74k_1.M.t1 VSS.t650 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X512 RES_74k_1.M.t1 VSS.t649 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X513 a_45028_11254.t1 a_45328_10632.t1 VDD.t217 ppolyf_u r_width=1.1u r_length=2.6u
X514 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t43 VDD.t630 VDD.t409 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X515 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t9 VDD.t46 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X516 VSS.t443 VSS.t441 VSS.t443 VSS.t442 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X517 VSS a_50708_569.t57 OUT.t21 VSS.t410 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X518 A_MUX_3.Tr_Gate_1.CLK S2.t9 VDD.t882 VDD.t881 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X519 RES_74k_1.P.t0 RES_74k_1.P.t1 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X520 CP_1_0.VCTRL ITAIL1.t9 a_32939_9624.t6 VSS.t328 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X521 VSS.t440 VSS.t439 VSS.t440 VSS.t350 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X522 RES_74k_1.M.t1 VSS.t648 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X523 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t46 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t11 VDD.t176 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X524 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t23 VCO_DFF_C_0.OUTB.t4 VSS.t113 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X525 A_MUX_1.Tr_Gate_1.CLK S1.t9 VDD.t768 VDD.t767 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X526 VSS A_MUX_0.Tr_Gate_1.CLK.t18 a_45158_5339.t0 VSS.t765 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X527 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t16 a_34443_2598.t6 VSS.t172 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X528 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t28 VDD.t56 VDD.t52 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X529 VDD a_22967_8787.t9 PFD_T2_0.INV_mag_1.IN.t16 VDD.t351 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X530 VDD a_50630_6066.t16 a_50528_5246.t20 VDD.t449 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X531 OUTB a_50528_5246.t66 VDD.t443 VDD.t442 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X532 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t23 VDD.t1042 VDD.t541 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X533 OUT a_50708_569.t58 VSS.t896 VSS.t0 nfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X534 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t12 VDD.t95 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X535 VSS.t438 VSS.t437 VSS.t438 VSS.t316 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X536 VSS VCTRL2.t32 a_34443_2598.t35 VSS.t757 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X537 UP1 a_27480_10186.t7 UP_OUT.t5 VDD.t41 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X538 RES_74k_1.M.t1 VSS.t647 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X539 OUTB a_50528_5246.t67 VDD.t445 VDD.t444 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X540 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t43 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t8 VDD.t525 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X541 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t18 VDD.t675 VDD.t188 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X542 VDD S2.t10 a_29875_10702.t4 VDD.t1035 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X543 VDD a_50810_1389.t17 a_50708_569.t16 VDD.t246 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X544 RES_74k_1.M.t1 VSS.t646 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X545 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUT.t19 VDD.t1111 VDD.t17 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X546 OUT a_50708_569.t59 VDD.t1019 VDD.t143 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X547 VDD a_22967_8787.t10 PFD_T2_0.INV_mag_1.IN.t11 VDD.t348 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X548 PFD_T2_0.INV_mag_0.IN a_22966_11778.t9 VDD.t906 VDD.t57 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X549 RES_74k_1.P.t67 RES_74k_1.P.t68 VDD.t21 ppolyf_u r_width=1.1u r_length=2.6u
X550 RES_74k_1.P.t35 RES_74k_1.P.t36 VDD.t131 ppolyf_u r_width=1.1u r_length=2.6u
X551 VDD a_50810_1389.t18 a_50708_569.t17 VDD.t249 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X552 RES_74k_1.M.t1 VSS.t645 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X553 OUT a_50708_569.t60 VDD.t1020 VDD.t244 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X554 RES_74k_1.M.t1 VSS.t644 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X555 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUT.t20 VDD.t1112 VDD.t19 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X556 VSS.t436 VSS.t434 VSS.t436 VSS.t435 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X557 VSS VCTRL2.t33 a_25706_n567.t37 VSS.t797 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X558 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t48 VDD.t237 VDD.t98 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X559 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t44 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t14 VDD.t393 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X560 OUT a_50708_569.t61 VDD.t1021 VDD.t825 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X561 VSS VCTRL2.t34 a_34443_2598.t34 VSS.t802 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X562 VDD S3.t9 A_MUX_4.Tr_Gate_1.CLK.t4 VDD.t380 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X563 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCTRL.t24 VDD.t790 VDD.t669 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X564 RES_74k_1.M.t1 VSS.t643 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X565 VSS.t433 VSS.t431 VSS.t433 VSS.t432 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X566 VDD S6.t6 A_MUX_2.Tr_Gate_1.CLK.t9 VDD.t564 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X567 RES_74k_1.M.t1 VSS.t642 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X568 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t24 VSS.t934 VSS.t339 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X569 OUT a_50708_569.t62 VDD.t814 VDD.t145 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X570 RES_74k_1.P.t29 RES_74k_1.P.t30 VDD.t21 ppolyf_u r_width=1.1u r_length=2.6u
X571 VCTRL_IN S4.t8 VCO_DFF_C_0.VCTRL.t0 VSS.t64 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X572 VDD.t963 VDD.t962 VDD.t963 VDD.t958 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X573 VSS.t430 VSS.t429 VSS.t430 VSS.t360 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X574 VDD a_50708_569.t63 OUT.t68 VDD.t679 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X575 VSS PFD_T2_0.INV_mag_0.OUT.t8 PFD_T2_0.Buffer_V_2_0.IN.t9 VSS.t940 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X576 a_45928_12082.t0 a_46228_11460.t0 VDD.t131 ppolyf_u r_width=1.1u r_length=2.6u
X577 OUTB a_50528_5246.t68 VSS.t182 VSS.t181 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X578 VSS.t428 VSS.t426 VSS.t428 VSS.t427 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X579 VSS VCTRL2.t35 a_34443_2598.t33 VSS.t978 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X580 VSS VCTRL2.t36 a_25706_n567.t36 VSS.t745 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X581 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t29 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t13 VSS.t18 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X582 VDD PFD_T2_0.INV_mag_1.IN.t24 PFD_T2_0.Buffer_V_2_0.IN.t6 VDD.t351 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X583 DIV_OUT a_20903_8375.t9 PFD_T2_0.FDIV.t7 VDD.t85 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X584 a_45928_10426.t0 a_45628_9804.t0 VDD.t243 ppolyf_u r_width=1.1u r_length=2.6u
X585 VDD a_50528_5246.t69 OUTB.t65 VDD.t446 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X586 VSS.t425 VSS.t423 VSS.t425 VSS.t424 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X587 A_MUX_2.Tr_Gate_1.CLK S6.t7 VDD.t1062 VDD.t567 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X588 a_42628_10426.t0 a_42628_9804.t0 VDD.t269 ppolyf_u r_width=1.1u r_length=2.6u
X589 VSS VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t45 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t1 VSS.t161 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X590 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_1837.t7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t1 VDD.t204 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X591 VSS.t422 VSS.t421 VSS.t422 VSS.t288 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X592 DN_OUT A_MUX_4.Tr_Gate_1.CLK.t18 DN1.t2 VSS.t119 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X593 VDD VCO_DFF_C_0.OUTB.t24 a_50630_6066.t0 VDD.t106 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X594 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t4 VSS.t269 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X595 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t20 VSS.t880 VSS.t879 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X596 DN1 a_25557_8739.t5 VSS.t338 VSS.t337 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X597 RES_74k_1.P.t5 RES_74k_1.P.t6 VDD.t21 ppolyf_u r_width=1.1u r_length=2.6u
X598 OUTB a_50528_5246.t70 VSS.t184 VSS.t183 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X599 VSS a_50708_569.t64 OUT.t19 VSS.t706 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X600 a_46228_11254.t0 a_45928_10632.t0 VDD.t131 ppolyf_u r_width=1.1u r_length=2.6u
X601 VSS.t420 VSS.t419 VSS.t420 VSS.t413 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X602 VSS.t418 VSS.t417 VSS.t418 VSS.t360 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X603 VDD S1.t10 A_MUX_1.Tr_Gate_1.CLK.t7 VDD.t769 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X604 VDD PFD_T2_0.INV_mag_1.IN.t25 PFD_T2_0.Buffer_V_2_0.IN.t5 VDD.t348 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X605 VDD a_50630_6066.t18 a_50528_5246.t15 VDD.t497 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X606 VSS.t416 VSS.t415 VSS.t416 VSS.t371 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X607 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t30 a_25706_n567.t3 VSS.t17 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X608 VDD PFD_T2_0.INV_mag_0.IN.t25 a_24437_9224.t0 VDD.t1092 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X609 PFD_T2_0.FDIV a_18508_8715.t8 VSS.t145 VDD.t364 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X610 VSS.t414 VSS.t412 VSS.t414 VSS.t413 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X611 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t49 VDD.t238 VDD.t88 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X612 VDD S4.t9 A_MUX_0.Tr_Gate_1.CLK.t0 VDD.t110 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X613 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t50 VDD.t239 VDD.t180 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X614 VDD PFD_T2_0.INV_mag_1.IN.t26 PFD_T2_0.INV_mag_1.OUT.t1 VDD.t345 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X615 VDD a_50528_5246.t71 OUTB.t64 VDD.t449 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X616 RES_74k_1.M.t1 VSS.t641 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X617 A_MUX_3.Tr_Gate_1.CLK S2.t11 VDD.t1077 VDD.t888 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X618 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCTRL.t25 VDD.t791 VDD.t784 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X619 VDD S5.t9 a_36685_10901.t4 VDD.t548 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X620 VDD a_50528_5246.t72 OUTB.t63 VDD.t452 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X621 RES_74k_1.M.t1 VSS.t640 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X622 PFD_T2_0.INV_mag_1.IN a_22967_8787.t11 VDD.t838 VDD.t837 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X623 A_MUX_2.Tr_Gate_1.CLK S6.t9 VDD.t1063 VDD.t206 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X624 a_44128_10426.t1 a_43828_9804.t1 VDD.t242 ppolyf_u r_width=1.1u r_length=2.6u
X625 A_MUX_2.Tr_Gate_1.CLK S6.t10 VSS.t825 VSS.t824 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X626 a_45628_9598.t0 a_45328_8976.t0 VDD.t22 ppolyf_u r_width=1.1u r_length=2.6u
X627 VDD a_50708_569.t65 OUT.t67 VDD.t246 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X628 RES_74k_1.P.t15 RES_74k_1.P.t16 VDD.t21 ppolyf_u r_width=1.1u r_length=2.6u
X629 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t18 a_25706_n567.t56 VSS.t17 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X630 RES_74k_1.M.t1 VSS.t639 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X631 VCO_DFF_C_0.VCTRL a_45158_5339.t8 CP_1_0.VCTRL.t4 VDD.t335 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X632 PRE_SCALAR A_MUX_1.Tr_Gate_1.CLK.t17 PFD_T2_0.FIN.t8 VSS.t343 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X633 UP1 a_25556_11637.t4 VSS.t75 VSS.t74 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X634 VSS S5.t10 a_36685_10901.t0 VSS.t246 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X635 PFD_T2_0.INV_mag_1.IN a_22967_8787.t12 VDD.t26 VDD.t25 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X636 RES_74k_1.P.t69 RES_74k_1.P.t70 VDD.t376 ppolyf_u r_width=1.1u r_length=2.6u
X637 VDD ITAIL.t10 ITAIL.t11 VDD.t423 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X638 RES_74k_1.P.t43 RES_74k_1.P.t44 VDD.t361 ppolyf_u r_width=1.1u r_length=2.6u
X639 OUTB a_50528_5246.t73 VSS.t186 VSS.t185 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X640 VSS S4.t10 A_MUX_0.Tr_Gate_1.CLK.t1 VSS.t65 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X641 VDD a_50708_569.t66 OUT.t66 VDD.t249 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X642 a_43528_8770.t0 a_43828_8148.t0 VDD.t133 ppolyf_u r_width=1.1u r_length=2.6u
X643 VSS VCTRL2.t39 a_34443_2598.t31 VSS.t779 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X644 RES_74k_1.M.t1 VSS.t638 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X645 VSS ITAIL1.t4 ITAIL1.t5 VSS.t332 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X646 VSS.t411 VSS.t409 VSS.t411 VSS.t410 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X647 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t44 VDD.t528 VDD.t402 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X648 RES_74k_1.M.t1 VSS.t637 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X649 VDD a_50708_569.t67 OUT.t65 VDD.t686 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X650 PFD_T2_0.INV_mag_0.IN a_22966_11778.t10 VDD.t1049 VDD.t1048 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X651 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t51 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t15 VDD.t171 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X652 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t46 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t13 VDD.t383 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X653 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t20 VDD.t676 VDD.t52 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X654 PFD_T2_0.FIN a_18550_11273.t7 F_IN.t1 VDD.t330 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X655 UP1 A_MUX_3.Tr_Gate_1.CLK.t18 UP_OUT.t3 VSS.t71 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X656 a_42928_12082.t1 a_43228_11460.t0 VDD.t376 ppolyf_u r_width=1.1u r_length=2.6u
X657 VDD VCO_DFF_C_0.VCTRL.t26 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t27 VDD.t666 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X658 VDD a_50708_569.t68 OUT.t64 VDD.t147 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X659 RES_74k_1.P.t55 RES_74k_1.P.t56 VDD.t361 ppolyf_u r_width=1.1u r_length=2.6u
X660 OUTB a_50528_5246.t74 VSS.t188 VSS.t187 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X661 VSS a_50528_5246.t75 OUTB.t13 VSS.t189 nfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X662 RES_74k_1.P.t88 RES_74k_1.P.t89 VDD.t133 ppolyf_u r_width=1.1u r_length=2.6u
X663 VDD a_50630_6066.t19 a_50528_5246.t14 VDD.t437 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X664 VDD a_50528_5246.t76 OUTB.t62 VDD.t446 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X665 RES_74k_1.M.t1 VSS.t636 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X666 RES_74k_1.P.t47 RES_74k_1.P.t48 VDD.t361 ppolyf_u r_width=1.1u r_length=2.6u
X667 A_MUX_0.Tr_Gate_1.CLK S4.t11 VDD.t114 VDD.t113 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X668 VSS a_50708_569.t69 OUT.t18 VSS.t580 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X669 PFD_T2_0.FDIV S6.t11 VSS.t826 VSS.t261 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X670 RES_74k_1.M.t1 VSS.t635 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X671 UP_OUT A_MUX_3.Tr_Gate_1.CLK.t19 UP1.t1 VSS.t245 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X672 DN_OUT A_MUX_4.Tr_Gate_1.CLK.t19 DN1.t1 VSS.t121 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X673 CP_1_0.VCTRL A_MUX_6.Tr_Gate_1.CLK.t17 RES_74k_1.P.t54 VSS.t277 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X674 VDD a_50528_5246.t77 OUTB.t61 VDD.t106 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X675 A_MUX_4.Tr_Gate_1.CLK S3.t10 VSS.t160 VSS.t159 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X676 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t45 VDD.t529 VDD.t386 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X677 VSS VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t46 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t1 VSS.t164 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X678 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.OUT.t21 VSS.t1001 VSS.t879 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X679 a_43228_11254.t0 a_42928_10632.t1 VDD.t376 ppolyf_u r_width=1.1u r_length=2.6u
X680 RES_74k_1.P.t21 RES_74k_1.P.t22 VDD.t361 ppolyf_u r_width=1.1u r_length=2.6u
X681 a_45328_8770.t0 a_45028_8148.t0 VDD.t217 ppolyf_u r_width=1.1u r_length=2.6u
X682 VSS a_50528_5246.t78 OUTB.t12 VSS.t309 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X683 UP1 a_27480_10186.t8 UP_OUT.t6 VDD.t42 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X684 VSS VCTRL2.t43 a_34443_2598.t29 VSS.t786 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X685 VSS VCTRL2.t44 a_25706_n567.t32 VSS.t745 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X686 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t21 VSS.t115 VSS.t114 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X687 VDD A_MUX_4.Tr_Gate_1.CLK.t20 a_27423_7180.t2 VDD.t130 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X688 VSS a_50810_1389.t21 a_50708_569.t7 VSS.t43 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X689 A_MUX_6.Tr_Gate_1.CLK S5.t11 VDD.t554 VDD.t270 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X690 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t28 VDD.t356 VDD.t25 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X691 OUTB a_50528_5246.t79 VDD.t637 VDD.t440 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X692 VDD a_50528_5246.t80 OUTB.t59 VDD.t497 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X693 RES_74k_1.M.t1 VSS.t634 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X694 A_MUX_0.Tr_Gate_1.CLK S4.t12 VDD.t116 VDD.t115 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X695 RES_74k_1.M.t1 VSS.t633 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X696 ITAIL ITAIL.t8 VDD.t695 VDD.t428 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X697 RES_74k_1.M.t1 VSS.t632 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X698 CP_1_0.VCTRL S5.t12 LF_OFFCHIP.t6 VSS.t122 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X699 OUT a_50708_569.t70 VDD.t826 VDD.t825 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X700 RES_74k_1.M.t1 VSS.t631 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X701 RES_74k_1.P.t49 RES_74k_1.P.t50 VDD.t217 ppolyf_u r_width=1.1u r_length=2.6u
X702 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t50 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t6 VDD.t308 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X703 OUTB a_50528_5246.t81 VDD.t640 VDD.t506 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X704 RES_74k_1.M.t4 VSS.t721 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X705 RES_74k_1.M.t1 VSS.t630 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X706 VDD a_50708_569.t71 OUT.t62 VDD.t679 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X707 VSS VCO_DFF_C_0.VCO_C_0.OUTB.t33 a_41879_n196.t0 VSS.t22 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X708 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t25 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t8 VSS.t269 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X709 VSS VCO_DFF_C_0.VCO_C_0.OUTB.t34 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t1 VSS.t25 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X710 OUT a_50708_569.t72 VDD.t682 VDD.t141 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X711 VSS a_18508_8715.t9 PFD_T2_0.FDIV.t15 VDD.t894 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X712 RES_74k_1.M.t1 VSS.t629 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X713 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t47 VDD.t387 VDD.t386 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X714 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL.t27 VDD.t794 VDD.t784 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X715 RES_74k_1.P.t11 RES_74k_1.P.t12 VDD.t242 ppolyf_u r_width=1.1u r_length=2.6u
X716 VSS.t408 VSS.t407 VSS.t408 VSS.t368 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X717 VSS.t406 VSS.t405 VSS.t406 VSS.t350 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X718 RES_74k_1.M.t5 VSS.t718 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X719 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t1 VSS.t146 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X720 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t48 VDD.t389 VDD.t388 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X721 VSS.t404 VSS.t403 VSS.t404 VSS.t295 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X722 RES_74k_1.M.t4 VSS.t720 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X723 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT a_41879_n196.t8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t1 VDD.t49 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X724 RES_74k_1.M.t1 VSS.t628 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X725 OUT a_50708_569.t73 VSS.t518 VSS.t88 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X726 a_44128_12082.t1 a_43828_11460.t1 VDD.t242 ppolyf_u r_width=1.1u r_length=2.6u
X727 VSS VCTRL2.t46 a_25706_n567.t31 VSS.t740 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X728 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t9 VDD.t576 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X729 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUT.t22 VSS.t1003 VSS.t1002 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X730 RES_74k_1.M.t5 VSS.t717 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X731 RES_74k_1.P a_39080_11413.t8 CP_1_0.VCTRL.t8 VDD.t413 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X732 PFD_T2_0.INV_mag_1.IN PFD_T2_0.FDIV.t18 a_22881_9554.t3 VSS.t907 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X733 VSS a_50528_5246.t82 OUTB.t11 VSS.t175 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X734 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t25 VCO_DFF_C_0.OUTB.t6 VSS.t147 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X735 VDD a_50528_5246.t83 OUTB.t57 VDD.t437 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X736 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCTRL.t28 VDD.t795 VDD.t666 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X737 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.IN.t2 a_24436_11277.t0 VDD.t1029 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X738 VSS.t402 VSS.t401 VSS.t402 VSS.t192 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X739 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUT.t23 VSS.t1005 VSS.t1004 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X740 OUTB a_50528_5246.t84 VDD.t643 VDD.t455 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X741 RES_74k_1.P a_39080_11413.t9 CP_1_0.VCTRL.t9 VDD.t414 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X742 VSS a_50708_569.t74 OUT.t16 VSS.t490 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X743 A_MUX_1.Tr_Gate_1.CLK S1.t13 VDD.t1024 VDD.t773 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X744 VSS.t400 VSS.t398 VSS.t400 VSS.t399 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X745 VDD PFD_T2_0.INV_mag_1.IN.t29 a_24436_11277.t2 VDD.t358 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X746 A_MUX_3.Tr_Gate_1.CLK S2.t12 VDD.t1078 VDD.t881 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X747 a_43828_11254.t0 a_44128_10632.t0 VDD.t242 ppolyf_u r_width=1.1u r_length=2.6u
X748 a_46528_10426.t0 a_46828_9598.t1 VDD.t109 ppolyf_u r_width=1.1u r_length=2.6u
X749 a_43528_10426.t1 a_43228_9804.t1 VDD.t262 ppolyf_u r_width=1.1u r_length=2.6u
X750 OUTB a_50528_5246.t85 VDD.t644 VDD.t134 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X751 PFD_T2_0.FIN S1.t14 F_IN.t5 VSS.t903 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X752 OUT a_50708_569.t75 VSS.t521 VSS.t48 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X753 A_MUX_4.Tr_Gate_1.CLK S3.t11 VDD.t285 VDD.t284 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X754 OUTB a_50528_5246.t86 VDD.t645 VDD.t440 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X755 OUT a_50708_569.t76 VDD.t683 VDD.t143 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X756 RES_74k_1.M.t1 VSS.t627 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X757 VDD S1.t15 A_MUX_1.Tr_Gate_1.CLK.t5 VDD.t775 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X758 OUTB a_50528_5246.t87 VDD.t646 VDD.t461 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X759 VDD VCO_DFF_C_0.OUT.t24 VCO_DFF_C_0.OUTB.t0 VDD.t6 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X760 OUT a_50708_569.t77 VDD.t685 VDD.t684 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X761 VSS PFD_T2_0.INV_mag_1.OUT.t7 a_22880_9797.t2 VSS.t525 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X762 VSS UP_OUT.t20 a_32939_9624.t0 VSS.t918 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X763 VDD a_50708_569.t78 OUT.t58 VDD.t686 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X764 RES_74k_1.P.t98 VSS.t282 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X765 OUT a_50708_569.t79 VDD.t1009 VDD.t825 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X766 VSS S6.t12 a_18508_8715.t0 VSS.t263 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X767 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t7 VDD.t390 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X768 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t7 VDD.t525 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X769 CP_1_0.VCTRL a_36685_10901.t8 LF_OFFCHIP.t1 VDD.t279 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X770 OUTB a_50528_5246.t88 VDD.t647 VDD.t136 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X771 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t50 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t10 VDD.t393 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X772 VDD.t961 VDD.t960 VDD.t961 VDD.t940 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X773 VSS VCTRL2.t49 a_25706_n567.t30 VSS.t797 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X774 OUT a_50708_569.t80 VDD.t1010 VDD.t12 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X775 VSS A_MUX_1.Tr_Gate_1.CLK.t18 a_20945_11785.t0 VSS.t344 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X776 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t18 VDD.t754 VDD.t753 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X777 RES_74k_1.M.t1 VSS.t626 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X778 VDD VCO_DFF_C_0.OUT.t25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t11 VDD.t9 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X779 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t10 VDD.t46 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X780 OUT a_50708_569.t81 VDD.t1011 VDD.t145 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X781 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t51 VDD.t397 VDD.t396 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X782 VSS VCTRL2.t51 a_34443_2598.t24 VSS.t802 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X783 VDD a_50810_1389.t24 a_50708_569.t10 VDD.t147 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X784 RES_74k_1.M.t1 VSS.t625 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X785 VDD a_50708_569.t82 OUT.t54 VDD.t679 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X786 DN1 A_MUX_4.Tr_Gate_1.CLK.t21 DN_OUT.t15 VSS.t948 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X787 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t51 VDD.t314 VDD.t93 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X788 RES_74k_1.P.t99 VSS.t283 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X789 RES_74k_1.P.t7 RES_74k_1.P.t8 VDD.t154 ppolyf_u r_width=1.1u r_length=2.6u
X790 VDD.t959 VDD.t957 VDD.t959 VDD.t958 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X791 VSS a_50708_569.t83 OUT.t14 VSS.t90 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X792 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t35 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t12 VSS.t14 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X793 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t5 VDD.t166 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X794 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t27 VSS.t272 VSS.t114 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X795 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t21 VDD.t999 VDD.t17 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X796 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t36 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t7 VDD.t185 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X797 PFD_T2_0.INV_mag_0.IN a_22966_11778.t11 VDD.t1051 VDD.t1050 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X798 a_44728_10426.t0 a_45028_9804.t0 VDD.t154 ppolyf_u r_width=1.1u r_length=2.6u
X799 VSS VCTRL2.t53 a_25706_n567.t28 VSS.t724 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X800 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT.t20 a_25706_n567.t58 VSS.t17 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X801 a_46228_9598.t0 a_46528_8976.t1 VDD.t272 ppolyf_u r_width=1.1u r_length=2.6u
X802 a_43228_9598.t1 a_42928_8976.t0 VDD.t376 ppolyf_u r_width=1.1u r_length=2.6u
X803 OUTB a_50528_5246.t89 VSS.t315 VSS.t314 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X804 RES_74k_1.M.t1 VSS.t624 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X805 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t9 VDD.t398 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X806 OUTB a_50528_5246.t90 VSS.t317 VSS.t316 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X807 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t22 VDD.t1000 VDD.t19 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X808 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t37 VDD.t189 VDD.t188 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X809 DN_INPUT a_29818_7696.t7 DN_OUT.t12 VDD.t288 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X810 VDD a_50630_6066.t20 a_50528_5246.t13 VDD.t452 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X811 VDD S4.t14 a_42763_5679.t2 VDD.t119 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X812 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t28 VDD.t579 VDD.t327 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X813 a_44728_12082.t1 a_45028_11460.t1 VDD.t154 ppolyf_u r_width=1.1u r_length=2.6u
X814 VSS.t397 VSS.t395 VSS.t397 VSS.t396 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X815 VSS VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t19 VCO_DFF_C_0.VCO_C_0.OUTB.t1 VSS.t547 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X816 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t2 VSS.t116 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X817 a_44728_8770.t0 a_44428_8148.t1 VDD.t31 ppolyf_u r_width=1.1u r_length=2.6u
X818 VSS.t394 VSS.t393 VSS.t394 VSS.t195 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X819 VSS a_50708_569.t84 OUT.t13 VSS.t50 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X820 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t48 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t19 VDD.t393 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X821 RES_74k_1.M.t1 VSS.t623 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X822 ITAIL ITAIL.t6 VDD.t694 VDD.t426 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X823 VSS.t392 VSS.t390 VSS.t392 VSS.t391 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X824 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t6 VDD.t534 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X825 RES_74k_1.M.t1 VSS.t622 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X826 A_MUX_6.Tr_Gate_1.CLK S5.t13 VDD.t556 VDD.t555 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X827 VDD S2.t13 a_29875_10702.t3 VDD.t62 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X828 VSS VCTRL2.t54 a_34443_2598.t23 VSS.t757 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X829 OUTB a_50528_5246.t91 VSS.t287 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X830 VDD a_50528_5246.t92 OUTB.t51 VDD.t138 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X831 VSS VCTRL2.t55 a_34443_2598.t22 VSS.t810 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X832 VDD.t956 VDD.t954 VDD.t956 VDD.t955 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X833 RES_74k_1.M.t1 VSS.t621 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X834 DN_INPUT a_29818_7696.t8 DN_OUT.t0 VDD.t0 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X835 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t9 VDD.t46 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X836 OUT a_50708_569.t85 VSS.t889 VSS.t483 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X837 a_45028_11254.t0 a_44728_10632.t1 VDD.t154 ppolyf_u r_width=1.1u r_length=2.6u
X838 RES_74k_1.P.t13 RES_74k_1.P.t14 VDD.t31 ppolyf_u r_width=1.1u r_length=2.6u
X839 VDD.t953 VDD.t951 VDD.t953 VDD.t952 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X840 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t50 VDD.t537 VDD.t409 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X841 VSS VCO_DFF_C_0.VCO_C_0.OUTB.t39 a_44716_1837.t0 VSS.t18 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X842 VDD PFD_T2_0.INV_mag_0.IN.t28 PFD_T2_0.INV_mag_0.OUT.t1 VDD.t345 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X843 VSS.t389 VSS.t387 VSS.t389 VSS.t388 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X844 VSS.t386 VSS.t384 VSS.t386 VSS.t385 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X845 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.IN.t29 VSS.t996 VSS.t995 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.5u
X846 PFD_T2_0.INV_mag_1.IN a_22967_8787.t13 VDD.t28 VDD.t27 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X847 VDD a_22966_11778.t12 PFD_T2_0.INV_mag_0.IN.t16 VDD.t1052 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X848 VSS VCTRL2.t56 a_34443_2598.t21 VSS.t757 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X849 VDD PFD_T2_0.INV_mag_0.IN.t30 PFD_T2_0.Buffer_V_2_1.IN.t4 VDD.t1052 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X850 VSS PFD_T2_0.INV_mag_1.IN.t30 a_23837_9553.t3 VSS.t569 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X851 VDD a_50528_5246.t93 OUTB.t50 VDD.t472 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X852 RES_74k_1.M.t1 VSS.t620 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X853 VDD a_22966_11778.t13 PFD_T2_0.INV_mag_0.IN.t11 VDD.t59 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X854 a_45928_8770.t0 a_46228_8148.t1 VDD.t131 ppolyf_u r_width=1.1u r_length=2.6u
X855 VDD a_50528_5246.t94 OUTB.t49 VDD.t458 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X856 VDD a_50708_569.t86 OUT.t53 VDD.t80 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X857 VSS PFD_T2_0.INV_mag_0.OUT.t9 PFD_T2_0.Buffer_V_2_0.IN.t10 VSS.t525 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X858 DN_OUT a_27423_7180.t7 DN1.t6 VDD.t267 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X859 A_MUX_4.Tr_Gate_1.CLK S3.t12 VDD.t287 VDD.t286 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X860 OUTB a_50528_5246.t95 VSS.t289 VSS.t288 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X861 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t17 VCO_DFF_C_0.VCO_C_0.OUT.t8 VDD.t126 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X862 VDD a_50708_569.t87 OUT.t52 VDD.t686 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X863 VSS S2.t14 A_MUX_3.Tr_Gate_1.CLK.t1 VSS.t36 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X864 DN_OUT a_29818_7696.t9 DN_INPUT.t4 VDD.t549 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X865 VDD PFD_T2_0.FIN.t18 a_22966_11778.t2 VDD.t59 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X866 PFD_T2_0.FDIV A_MUX_2.Tr_Gate_1.CLK.t18 DIV_OUT.t0 VSS.t53 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X867 VSS VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t53 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t0 VSS.t164 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X868 VDD a_50708_569.t88 OUT.t51 VDD.t14 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X869 RES_74k_1.M.t1 VSS.t619 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X870 VCO_DFF_C_0.VCTRL a_42763_5679.t8 VCTRL_IN.t1 VDD.t117 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X871 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t5 VDD.t90 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X872 VDD a_50708_569.t89 OUT.t50 VDD.t147 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X873 VDD ITAIL.t4 ITAIL.t5 VDD.t429 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X874 RES_74k_1.P.t31 RES_74k_1.P.t32 VDD.t131 ppolyf_u r_width=1.1u r_length=2.6u
X875 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t20 VCO_DFF_C_0.VCO_C_0.OUTB.t6 VDD.t755 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X876 VSS.t383 VSS.t381 VSS.t383 VSS.t382 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X877 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t25 VDD.t257 VDD.t188 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X878 VDD PFD_T2_0.Buffer_V_2_1.IN.t12 a_25556_11637.t1 VDD.t573 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X879 VDD A_MUX_6.Tr_Gate_1.CLK.t18 a_39080_11413.t3 VDD.t413 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X880 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t4 VDD.t171 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X881 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN a_44716_n517.t8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t8 VDD.t201 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X882 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t40 a_41879_n196.t5 VDD.t105 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X883 OUT a_50708_569.t90 VSS.t522 VSS.t12 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X884 CP_1_0.VCTRL ITAIL.t24 a_32731_10265.t5 VDD.t428 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X885 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.IN.t6 a_24437_9224.t2 VDD.t340 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X886 VDD S3.t14 a_29818_7696.t4 VDD.t288 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X887 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t18 VDD.t129 VDD.t124 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X888 RES_74k_1.M.t1 VSS.t618 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X889 RES_74k_1.M.t1 VSS.t617 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X890 VDD VCO_DFF_C_0.VCTRL.t29 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t28 VDD.t669 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X891 VDD S5.t14 A_MUX_6.Tr_Gate_1.CLK.t5 VDD.t273 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X892 VDD A_MUX_6.Tr_Gate_1.CLK.t19 a_39080_11413.t2 VDD.t414 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X893 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t32 VDD.t357 VDD.t27 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X894 VDD a_50528_5246.t96 OUTB.t48 VDD.t452 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X895 VSS.t380 VSS.t379 VSS.t380 VSS.t200 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X896 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t23 VCO_DFF_C_0.OUT VDD.t750 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X897 VDD S5.t15 A_MUX_6.Tr_Gate_1.CLK.t4 VDD.t276 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X898 a_42928_10426.t1 a_42628_9804.t1 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X899 A_MUX_0.Tr_Gate_1.CLK S4.t15 VDD.t538 VDD.t113 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X900 VCO_DFF_C_0.VCTRL A_MUX_0.Tr_Gate_1.CLK.t20 CP_1_0.VCTRL.t32 VSS.t909 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X901 VSS A_MUX_6.Tr_Gate_1.CLK.t20 a_39080_11413.t0 VSS.t278 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X902 VSS S3.t15 a_29818_7696.t0 VSS.t133 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X903 RES_74k_1.M.t1 VSS.t616 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X904 VSS a_50708_569.t91 OUT.t10 VSS.t382 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X905 PFD_T2_0.FIN A_MUX_1.Tr_Gate_1.CLK.t19 PRE_SCALAR.t4 VSS.t266 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X906 PFD_T2_0.FDIV S6.t14 VSS.t830 VSS.t829 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X907 VDD S3.t16 a_29818_7696.t3 VDD.t0 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X908 OUT a_50708_569.t92 VDD.t706 VDD.t684 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X909 VDD.t950 VDD.t948 VDD.t950 VDD.t949 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X910 RES_74k_1.M.t1 VSS.t615 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X911 VCO_DFF_C_0.VCTRL a_45158_5339.t9 CP_1_0.VCTRL.t5 VDD.t336 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X912 VSS a_50528_5246.t97 OUTB.t6 VSS.t258 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X913 RES_74k_1.P.t100 VSS.t284 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X914 RES_74k_1.M.t1 VSS.t614 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X915 ITAIL1 ITAIL1.t2 VSS.t331 VSS.t330 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X916 VDD a_50708_569.t93 OUT.t48 VDD.t220 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X917 PRE_SCALAR a_20945_11785.t8 PFD_T2_0.FIN.t3 VDD.t165 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X918 VDD S6.t15 A_MUX_2.Tr_Gate_1.CLK.t6 VDD.t891 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X919 RES_74k_1.M.t1 VSS.t613 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X920 VSS a_50810_1389.t25 a_50708_569.t19 VSS.t706 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X921 VDD A_MUX_3.Tr_Gate_1.CLK.t20 a_27480_10186.t2 VDD.t42 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X922 VDD S6.t16 a_18508_8715.t2 VDD.t894 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X923 VDD.t947 VDD.t945 VDD.t947 VDD.t946 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X924 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t51 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t22 VDD.t519 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X925 RES_74k_1.M.t1 VSS.t612 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X926 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t4 VSS.t148 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X927 CP_1_0.VCTRL a_36685_10901.t9 LF_OFFCHIP.t0 VDD.t563 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X928 A_MUX_0.Tr_Gate_1.CLK S4.t16 VDD.t539 VDD.t115 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X929 RES_74k_1.M.t1 VSS.t611 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X930 RES_74k_1.M.t1 VSS.t610 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X931 PRE_SCALAR a_20945_11785.t9 PFD_T2_0.FIN.t0 VDD.t153 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X932 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_1284.t8 VCO_DFF_C_0.OUTB.t15 VDD.t44 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X933 A_MUX_0.Tr_Gate_1.CLK S4.t17 VSS.t233 VSS.t65 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X934 VSS VCTRL2.t61 a_34443_2598.t19 VSS.t779 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X935 VSS VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t5 VSS.t116 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X936 VCO_DFF_C_0.VCTRL S4.t18 VCTRL_IN.t5 VSS.t234 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X937 OUTB a_50528_5246.t98 VDD.t599 VDD.t598 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X938 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL.t30 VDD.t798 VDD.t672 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X939 VDD a_50708_569.t94 OUT.t47 VDD.t723 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X940 OUT a_50708_569.t95 VDD.t875 VDD.t78 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X941 DN1 a_27423_7180.t8 DN_OUT.t6 VDD.t540 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X942 a_44128_10426.t0 a_44428_9804.t0 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X943 VSS VCTRL2.t62 a_25706_n567.t24 VSS.t740 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X944 VSS.t378 VSS.t376 VSS.t378 VSS.t377 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X945 A_MUX_1.Tr_Gate_1.CLK S1.t16 VSS.t905 VSS.t904 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X946 a_45628_9598.t1 a_45928_8976.t0 VDD.t243 ppolyf_u r_width=1.1u r_length=2.6u
X947 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t54 VDD.t401 VDD.t388 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X948 VSS a_22966_11778.t14 a_22880_10947.t2 VSS.t836 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X949 a_42628_9598.t0 a_42628_8770.t0 VDD.t269 ppolyf_u r_width=1.1u r_length=2.6u
X950 OUTB a_50528_5246.t99 VDD.t600 VDD.t455 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X951 RES_74k_1.M.t1 VSS.t609 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X952 RES_74k_1.M.t1 VSS.t608 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X953 A_MUX_0.Tr_Gate_1.CLK S4.t19 VSS.t235 VSS.t65 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X954 VDD.t944 VDD.t942 VDD.t944 VDD.t943 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X955 VSS a_50630_6066.t23 a_50528_5246.t21 VSS.t309 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X956 VCTRL_IN a_42763_5679.t9 VCO_DFF_C_0.VCTRL.t6 VDD.t119 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X957 OUT a_50708_569.t96 VSS.t768 VSS.t108 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X958 UP_OUT A_MUX_3.Tr_Gate_1.CLK.t21 UP1.t0 VSS.t9 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X959 VDD S2.t16 A_MUX_3.Tr_Gate_1.CLK.t5 VDD.t763 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X960 VSS VCTRL2.t64 a_34443_2598.t17 VSS.t779 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X961 F_IN a_18550_11273.t8 PFD_T2_0.FIN.t6 VDD.t331 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X962 VSS S6.t17 A_MUX_2.Tr_Gate_1.CLK.t0 VSS.t831 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X963 VSS a_50528_5246.t100 OUTB.t5 VSS.t292 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X964 VSS VCTRL2.t65 a_25706_n567.t23 VSS.t797 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X965 VSS S1.t17 A_MUX_1.Tr_Gate_1.CLK.t0 VSS.t915 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X966 VSS a_50708_569.t97 OUT.t8 VSS.t301 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X967 OUTB a_50528_5246.t101 VDD.t601 VDD.t461 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X968 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t55 VDD.t403 VDD.t402 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X969 VSS.t375 VSS.t373 VSS.t375 VSS.t374 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X970 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t23 VDD.t383 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X971 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t19 VSS.t241 VSS.t240 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X972 ITAIL1 ITAIL1.t0 VSS.t329 VSS.t328 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X973 VSS VCTRL2.t67 a_34443_2598.t15 VSS.t729 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X974 UP_OUT S2.t17 UP_INPUT.t6 VSS.t550 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X975 RES_74k_1.M.t1 VSS.t607 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X976 CP_1_0.VCTRL S5.t17 LF_OFFCHIP.t5 VSS.t124 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X977 OUTB a_50528_5246.t102 VDD.t602 VDD.t506 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X978 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t53 VDD.t734 VDD.t388 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X979 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t42 a_25706_n567.t7 VSS.t78 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X980 RES_74k_1.M.t1 VSS.t606 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X981 a_43828_9598.t0 a_44128_8976.t1 VDD.t242 ppolyf_u r_width=1.1u r_length=2.6u
X982 OUTB a_50528_5246.t103 VDD.t604 VDD.t603 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X983 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_n517.t9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t17 VDD.t204 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X984 VSS VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t24 VCO_DFF_C_0.OUT VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X985 UP_INPUT a_29875_10702.t7 UP_OUT.t13 VDD.t62 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X986 PFD_T2_0.FDIV S6.t18 VSS.t262 VSS.t261 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X987 DIV_OUT A_MUX_2.Tr_Gate_1.CLK.t19 PFD_T2_0.FDIV.t11 VSS.t766 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X988 DN_INPUT S3.t18 DN_OUT.t10 VSS.t158 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X989 OUT a_50708_569.t98 VSS.t771 VSS.t377 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X990 VDD a_22966_11778.t15 PFD_T2_0.INV_mag_0.IN.t12 VDD.t909 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X991 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t54 VSS.t546 VSS.t306 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X992 VDD a_50708_569.t99 OUT.t45 VDD.t80 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X993 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t54 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t6 VDD.t171 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X994 RES_74k_1.M.t1 VSS.t605 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X995 RES_74k_1.M.t1 VSS.t604 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X996 OUT a_50708_569.t100 VDD.t878 VDD.t684 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X997 RES_74k_1.M.t1 VSS.t603 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X998 OUTB a_50528_5246.t104 VDD.t606 VDD.t605 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X999 VSS.t372 VSS.t370 VSS.t372 VSS.t371 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X1000 UP_INPUT a_29875_10702.t8 UP_OUT.t14 VDD.t1035 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1001 a_45328_8770.t1 a_45628_8148.t1 VDD.t22 ppolyf_u r_width=1.1u r_length=2.6u
X1002 PFD_T2_0.INV_mag_1.IN a_22967_8787.t14 VDD.t30 VDD.t29 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1003 RES_74k_1.P.t39 RES_74k_1.P.t40 VDD.t21 ppolyf_u r_width=1.1u r_length=2.6u
X1004 OUT a_50708_569.t101 VDD.t879 VDD.t12 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.5u
X1005 VSS a_50528_5246.t105 OUTB.t4 VSS.t295 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1006 VDD VCO_DFF_C_0.OUT.t28 a_50810_1389.t2 VDD.t14 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1007 RES_74k_1.M.t1 VSS.t602 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1008 VSS.t369 VSS.t367 VSS.t369 VSS.t368 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X1009 RES_74k_1.P.t91 RES_74k_1.P.t92 VDD.t243 ppolyf_u r_width=1.1u r_length=2.6u
X1010 VSS VCTRL2.t69 a_25706_n567.t21 VSS.t724 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1011 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t43 a_44716_1837.t2 VDD.t194 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1012 OUT a_50708_569.t102 VDD.t75 VDD.t74 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1013 RES_74k_1.M.t1 VSS.t601 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1014 CP_1_0.VCTRL A_MUX_0.Tr_Gate_1.CLK.t21 VCO_DFF_C_0.VCTRL.t12 VSS.t911 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1015 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t21 VCO_DFF_C_0.VCO_C_0.OUTB.t5 VDD.t758 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1016 VSS.t366 VSS.t364 VSS.t366 VSS.t365 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X1017 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t7 VDD.t185 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1018 VSS S2.t18 A_MUX_3.Tr_Gate_1.CLK.t0 VSS.t551 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1019 RES_74k_1.P.t9 RES_74k_1.P.t10 VDD.t22 ppolyf_u r_width=1.1u r_length=2.6u
X1020 VSS a_50708_569.t103 OUT.t6 VSS.t43 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1021 RES_74k_1.P.t2 RES_74k_1.P.t3 VDD.t21 ppolyf_u r_width=1.1u r_length=2.6u
X1022 OUT a_50708_569.t104 VDD.t77 VDD.t76 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1023 PFD_T2_0.FIN S1.t18 F_IN.t4 VSS.t903 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1024 CP_1_0.VCTRL ITAIL.t25 a_32731_10265.t4 VDD.t426 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X1025 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t20 VCO_DFF_C_0.VCO_C_0.OUT.t6 VDD.t126 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1026 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN a_41879_n196.t9 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t1 VDD.t132 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1027 VSS a_50528_5246.t106 OUTB.t3 VSS.t192 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1028 VDD.t941 VDD.t939 VDD.t941 VDD.t940 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X1029 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t55 VDD.t175 VDD.t174 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X1030 VDD VCO_DFF_C_0.VCTRL.t31 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t18 VDD.t672 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.84u
X1031 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t45 VSS.t80 VSS.t79 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1032 VSS S5.t18 A_MUX_6.Tr_Gate_1.CLK.t1 VSS.t125 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1033 VDD a_50630_6066.t26 a_50528_5246.t3 VDD.t138 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1034 OUTB a_50528_5246.t107 VDD.t456 VDD.t455 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1035 RES_74k_1.M.t1 VSS.t600 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1036 VDD S1.t19 a_18550_11273.t3 VDD.t331 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1037 a_45928_12082.t1 a_45628_11460.t1 VDD.t243 ppolyf_u r_width=1.1u r_length=2.6u
X1038 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t19 a_34443_2598.t57 VSS.t932 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1039 VDD a_25556_11637.t5 UP1.t10 VDD.t157 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1040 VCO_DFF_C_0.OUTB a_41879_1284.t9 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t0 VDD.t105 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1041 VSS S5.t19 A_MUX_6.Tr_Gate_1.CLK.t0 VSS.t128 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1042 RES_74k_1.P.t23 RES_74k_1.P.t24 VDD.t361 ppolyf_u r_width=1.1u r_length=2.6u
X1043 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t25 VDD.t1003 VDD.t17 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1044 VCO_DFF_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t6 VSS.t110 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1045 OUTB a_50528_5246.t108 VDD.t457 VDD.t134 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1046 VSS.t363 VSS.t362 VSS.t363 VSS.t323 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X1047 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t21 a_34443_2598.t1 VSS.t171 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1048 RES_74k_1.M.t6 VSS.t719 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1049 ITAIL ITAIL.t2 VDD.t691 VDD.t428 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X1050 VDD PFD_T2_0.Buffer_V_2_0.IN.t13 a_25557_8739.t1 VDD.t160 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1051 VDD a_50630_6066.t27 a_50528_5246.t12 VDD.t472 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1052 OUT a_50708_569.t105 VSS.t47 VSS.t46 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1053 VDD a_50528_5246.t109 OUTB.t39 VDD.t458 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X1054 OUTB a_50528_5246.t110 VDD.t462 VDD.t461 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1055 VDD a_50810_1389.t26 a_50708_569.t20 VDD.t220 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1056 UP_INPUT S2.t19 UP_OUT.t10 VSS.t167 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1057 a_45628_11254.t1 a_45928_10632.t1 VDD.t243 ppolyf_u r_width=1.1u r_length=2.6u
X1058 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t30 VDD.t542 VDD.t541 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1059 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.VCO_C_0.OUTB.t46 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t11 VSS.t14 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1060 RES_74k_1.M.t1 VSS.t599 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1061 VDD A_MUX_1.Tr_Gate_1.CLK.t20 a_20945_11785.t3 VDD.t165 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1062 RES_74k_1.P.t57 RES_74k_1.P.t58 VDD.t361 ppolyf_u r_width=1.1u r_length=2.6u
X1063 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t55 VDD.t735 VDD.t409 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1064 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.VCO_C_0.OUTB.t47 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t13 VSS.t15 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1065 OUTB a_50528_5246.t111 VDD.t463 VDD.t136 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1066 VSS S3.t19 A_MUX_4.Tr_Gate_1.CLK.t6 VSS.t711 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1067 VDD S3.t20 A_MUX_4.Tr_Gate_1.CLK.t7 VDD.t377 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1068 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t53 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t3 VDD.t95 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1069 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t54 VDD.t320 VDD.t319 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1070 VSS PFD_T2_0.INV_mag_1.OUT.t8 PFD_T2_0.Buffer_V_2_1.IN.t9 VSS.t528 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1071 VDD VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t56 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t5 VDD.t404 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1072 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t56 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t5 VDD.t534 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1073 VDD VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t56 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t8 VDD.t176 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1074 VSS.t361 VSS.t359 VSS.t361 VSS.t360 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X1075 RES_74k_1.M.t1 VSS.t598 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1076 VDD A_MUX_1.Tr_Gate_1.CLK.t21 a_20945_11785.t2 VDD.t153 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1077 DIV_OUT A_MUX_2.Tr_Gate_1.CLK.t21 PFD_T2_0.FDIV.t12 VSS.t767 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1078 VDD a_50528_5246.t112 OUTB.t36 VDD.t464 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1079 VDD.t938 VDD.t936 VDD.t938 VDD.t937 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X1080 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t22 VDD.t762 VDD.t761 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1081 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUT.t29 VDD.t18 VDD.t17 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1082 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t29 VCO_DFF_C_0.OUTB.t5 VSS.t141 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1083 VSS VCTRL2.t73 a_25706_n567.t19 VSS.t740 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1084 VSS VCO_DFF_C_0.OUT.t30 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t4 VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1085 VSS PFD_T2_0.INV_mag_1.OUT.t9 PFD_T2_0.Buffer_V_2_1.IN.t8 VSS.t531 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1086 UP_OUT a_29875_10702.t9 UP_INPUT.t0 VDD.t65 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1087 VDD a_50810_1389.t27 a_50708_569.t21 VDD.t723 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1088 OUT a_50708_569.t106 VDD.t79 VDD.t78 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1089 VDD a_50708_569.t107 OUT.t39 VDD.t80 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1090 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t57 VDD.t408 VDD.t407 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1091 VDD a_50528_5246.t113 OUTB.t35 VDD.t467 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1092 RES_74k_1.M.t1 VSS.t597 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1093 VSS.t358 VSS.t356 VSS.t358 VSS.t357 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X1094 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT a_44716_1837.t8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t14 VDD.t192 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1095 VSS PFD_T2_0.Buffer_V_2_1.IN.t13 a_25556_11637.t0 VSS.t74 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1096 RES_74k_1.M.t1 VSS.t596 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1097 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUT.t31 VDD.t20 VDD.t19 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1098 a_43528_10426.t0 a_43828_9804.t0 VDD.t133 ppolyf_u r_width=1.1u r_length=2.6u
X1099 VSS S4.t20 a_42763_5679.t0 VSS.t64 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1100 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.OUT.t32 VDD.t744 VDD.t743 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1101 OUT a_50708_569.t108 VSS.t49 VSS.t48 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1102 VDD a_50708_569.t109 OUT.t38 VDD.t14 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1103 VSS VCTRL2.t74 a_34443_2598.t12 VSS.t802 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X1104 RES_74k_1.P.t83 RES_74k_1.P.t84 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X1105 RES_74k_1.M.t1 VSS.t595 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1106 PFD_T2_0.INV_mag_0.IN PFD_T2_0.FIN.t19 a_22880_10947.t0 VSS.t32 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1107 RES_74k_1.P.t37 RES_74k_1.P.t38 VDD.t109 ppolyf_u r_width=1.1u r_length=2.6u
X1108 VDD a_50708_569.t110 OUT.t37 VDD.t32 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1109 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t55 VDD.t321 VDD.t98 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1110 OUTB a_50528_5246.t114 VSS.t196 VSS.t195 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1111 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t57 VDD.t179 VDD.t103 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1112 VDD VCO_DFF_C_0.OUT.t33 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t9 VDD.t745 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1113 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.OUT.t34 VDD.t749 VDD.t748 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1114 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t58 VDD.t410 VDD.t409 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1115 VDD VCO_DFF_C_0.VCTRL.t32 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t17 VDD.t784 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1116 RES_74k_1.M.t1 VSS.t594 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1117 VSS S6.t19 PFD_T2_0.FDIV.t6 VSS.t263 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1118 F_IN a_18550_11273.t9 PFD_T2_0.FIN.t7 VDD.t332 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1119 VSS.t355 VSS.t354 VSS.t355 VSS.t298 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X1120 UP_INPUT S2.t20 UP_OUT.t9 VSS.t168 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1121 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t56 VSS.t140 VSS.t139 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1122 VDD.t935 VDD.t933 VDD.t935 VDD.t934 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X1123 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t49 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t5 VDD.t46 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1124 VDD a_50528_5246.t115 OUTB.t34 VDD.t138 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1125 VSS VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t21 VCO_DFF_C_0.VCO_C_0.OUT.t0 VSS.t242 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1126 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t7 VDD.t543 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1127 VDD VCO_DFF_C_0.VCO_C_0.OUTB.t51 a_41879_n196.t2 VDD.t49 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1128 OUT a_50708_569.t111 VSS.t100 VSS.t99 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1129 VDD S2.t21 A_MUX_3.Tr_Gate_1.CLK.t4 VDD.t69 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1130 a_42928_12082.t0 a_42628_11460.t0 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X1131 a_46528_12082.t0 a_46828_11254.t1 VDD.t109 ppolyf_u r_width=1.1u r_length=2.6u
X1132 VSS VCTRL2.t77 a_34443_2598.t11 VSS.t802 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X1133 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t23 VSS.t348 VSS.t347 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1134 VSS.t353 VSS.t352 VSS.t353 VSS.t205 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.5u
X1135 RES_74k_1.M.t1 VSS.t593 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1136 RES_74k_1.M.t1 VSS.t592 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1137 RES_74k_1.M.t7 VSS.t542 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1138 A_MUX_1.Tr_Gate_1.CLK S1.t20 VDD.t1032 VDD.t767 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1139 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.VCO_C_0.OUTB.t52 VDD.t53 VDD.t52 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1140 OUT a_50708_569.t112 VSS.t102 VSS.t101 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1141 a_45328_10426.t1 a_45028_9804.t1 VDD.t217 ppolyf_u r_width=1.1u r_length=2.6u
X1142 RES_74k_1.P.t101 VSS.t285 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X1143 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t26 VSS.t878 VSS.t143 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1144 VDD VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t6 VDD.t185 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1145 a_46828_9598.t0 a_46528_8976.t0 VDD.t109 ppolyf_u r_width=1.1u r_length=2.6u
X1146 RES_74k_1.P.t102 VSS.t286 cap_mim_2f0_m4m5_noshield c_width=30u c_length=30u
X1147 UP_OUT a_27480_10186.t9 UP1.t7 VDD.t43 pfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1148 a_43228_9598.t0 a_43528_8976.t0 VDD.t262 ppolyf_u r_width=1.1u r_length=2.6u
X1149 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t27 VCO_DFF_C_0.OUT VDD.t6 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1150 VDD VCO_DFF_C_0.VCTRL.t33 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t21 VDD.t666 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1151 VDD VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t57 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t26 VDD.t398 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1152 RES_74k_1.M.t1 VSS.t591 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1153 RES_74k_1.M.t1 VSS.t590 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1154 PFD_T2_0.INV_mag_1.IN a_22967_8787.t16 VDD.t712 VDD.t343 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1155 a_42628_11254.t0 a_42928_10632.t0 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X1156 VDD a_50528_5246.t116 OUTB.t33 VDD.t472 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1157 VSS.t351 VSS.t349 VSS.t351 VSS.t350 nfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.84u
X1158 VSS a_50708_569.t113 OUT.t1 VSS.t103 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1159 VDD a_22966_11778.t16 PFD_T2_0.INV_mag_0.IN.t13 VDD.t912 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1160 a_46828_11254.t0 a_46528_10632.t0 VDD.t109 ppolyf_u r_width=1.1u r_length=2.6u
X1161 VDD a_50528_5246.t117 OUTB.t32 VDD.t458 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.5u
X1162 RES_74k_1.M.t7 VSS.t541 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1163 VDD a_50708_569.t114 OUT.t36 VDD.t220 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1164 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t30 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t2 VSS.t142 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1165 VDD a_50708_569.t115 OUT.t35 VDD.t223 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1166 LF_OFFCHIP S5.t21 CP_1_0.VCTRL.t22 VSS.t246 nfet_03v3 ad=0.218p pd=1.36u as=0.37p ps=2.56u w=0.84u l=0.5u
X1167 VDD PFD_T2_0.INV_mag_0.IN.t32 PFD_T2_0.Buffer_V_2_1.IN.t3 VDD.t912 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1168 DN_OUT a_27423_7180.t9 DN1.t4 VDD.t665 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1169 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t58 VDD.t740 VDD.t513 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1170 VDD VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t22 VCO_DFF_C_0.VCO_C_0.OUT.t5 VDD.t503 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1171 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB.t53 a_25706_n567.t1 VSS.t17 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1172 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t57 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t4 VDD.t322 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1173 VDD VCO_DFF_C_0.OUT.t35 VCO_DFF_C_0.OUTB.t9 VDD.t750 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1174 RES_74k_1.M.t1 VSS.t589 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1175 VDD VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t31 a_41879_1284.t2 VDD.t105 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1176 VDD a_50708_569.t116 OUT.t34 VDD.t35 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1177 VCO_DFF_C_0.VCTRL S4.t21 VCTRL_IN.t4 VSS.t153 nfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1178 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t58 VDD.t181 VDD.t180 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1179 RES_74k_1.P A_MUX_6.Tr_Gate_1.CLK.t21 CP_1_0.VCTRL.t0 VSS.t68 nfet_03v3 ad=0.37p pd=2.56u as=0.37p ps=2.56u w=0.84u l=0.5u
X1180 VDD S3.t21 A_MUX_4.Tr_Gate_1.CLK.t8 VDD.t380 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1181 VSS VCTRL2.t78 a_25706_n567.t16 VSS.t745 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.84u
X1182 VDD a_50708_569.t117 OUT.t33 VDD.t723 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1183 OUT a_50708_569.t118 VDD.t726 VDD.t78 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1184 VSS PFD_T2_0.INV_mag_0.IN.t33 a_23836_10693.t0 VSS.t992 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1185 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t23 VDD.t885 VDD.t122 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1186 VDD S6.t20 A_MUX_2.Tr_Gate_1.CLK.t5 VDD.t564 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X1187 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT a_44716_1837.t9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t7 VDD.t194 pfet_03v3 ad=0.37p pd=2.56u as=0.218p ps=1.36u w=0.84u l=0.5u
X1188 RES_74k_1.M.t1 VSS.t588 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1189 a_45028_9598.t0 a_44728_8976.t0 VDD.t154 ppolyf_u r_width=1.1u r_length=2.6u
X1190 VDD VCO_DFF_C_0.VCTRL.t34 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t5 VDD.t669 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.84u
X1191 RES_74k_1.P.t51 RES_74k_1.P.t52 VDD.t133 ppolyf_u r_width=1.1u r_length=2.6u
X1192 RES_74k_1.M.t1 VSS.t587 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1193 VDD S1.t21 a_18550_11273.t2 VDD.t332 pfet_03v3 ad=0.218p pd=1.36u as=0.218p ps=1.36u w=0.84u l=0.5u
X1194 VDD ITAIL.t0 ITAIL.t1 VDD.t429 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X1195 A_MUX_2.Tr_Gate_1.CLK S6.t21 VDD.t568 VDD.t567 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1196 VSS a_50528_5246.t118 OUTB.t1 VSS.t197 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1197 VSS VCTRL2.t79 a_25706_n567.t15 VSS.t797 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1198 VDD VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t58 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t1 VDD.t176 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1199 VSS a_50708_569.t119 OUT.t0 VSS.t543 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1200 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.INV_mag_1.IN.t33 a_23837_9553.t0 VSS.t568 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X1201 a_46528_8770.t0 a_46228_8148.t0 VDD.t272 ppolyf_u r_width=1.1u r_length=2.6u
X1202 VSS a_50528_5246.t119 OUTB.t0 VSS.t200 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.5u
X1203 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCTRL.t35 VDD.t673 VDD.t672 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.84u
X1204 RES_74k_1.M.t1 VSS.t586 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
R0 a_42928_8770.t0 a_42928_8770.t1 12.9675
R1 a_43228_8148.t0 a_43228_8148.t1 12.9675
R2 VDD.n1520 VDD.n322 130000
R3 VDD.n1301 VDD.n471 129000
R4 VDD.n1521 VDD.n1520 65000
R5 VDD.n1256 VDD.n471 64500
R6 VDD.n1710 VDD.n1709 6501.29
R7 VDD.n1468 VDD.n1467 947.995
R8 VDD.n1522 VDD.n314 947.995
R9 VDD.n1273 VDD.n1249 947.995
R10 VDD.n1264 VDD.n1257 947.995
R11 VDD.n1467 VDD.n1458 944.883
R12 VDD.n1458 VDD.n321 944.883
R13 VDD.n1266 VDD.n1265 944.883
R14 VDD.n1265 VDD.n1264 944.883
R15 VDD.n1522 VDD.n1521 842.52
R16 VDD.n1256 VDD.n1249 842.52
R17 VDD.n1710 VDD.n1649 447.029
R18 VDD.t339 VDD.t337 432.243
R19 VDD.n1519 VDD.n280 371.986
R20 VDD.n1289 VDD.n478 371.986
R21 VDD.n1507 VDD.n1506 353.928
R22 VDD.n1304 VDD.n468 353.928
R23 VDD.n1508 VDD.n1507 350.877
R24 VDD.n1512 VDD.n323 350.877
R25 VDD.n1300 VDD.n473 350.877
R26 VDD.n1304 VDD.n1303 350.877
R27 VDD.t571 VDD.t1085 339.613
R28 VDD.t418 VDD.t1079 316.279
R29 VDD.t337 VDD.t160 316.279
R30 VDD.n1512 VDD.n322 312.866
R31 VDD.n1301 VDD.n1300 312.866
R32 VDD.n1674 VDD.n1673 310.428
R33 VDD.n1675 VDD.n1674 307.495
R34 VDD.n1675 VDD.n1658 307.495
R35 VDD.n1660 VDD.n1659 307.495
R36 VDD.n1684 VDD.n1660 307.495
R37 VDD.n1707 VDD.n1651 307.495
R38 VDD.n1700 VDD.n1651 307.495
R39 VDD.n1698 VDD.n1697 307.495
R40 VDD.n1697 VDD.n1685 307.495
R41 VDD.n1690 VDD.n1649 307.495
R42 VDD.n1708 VDD.n1650 304.911
R43 VDD.t973 VDD.n1519 283.627
R44 VDD.n1289 VDD.t978 283.627
R45 VDD.t155 VDD.t157 282.159
R46 VDD.t573 VDD.t571 282.159
R47 VDD.n1510 VDD.t666 279.885
R48 VDD.t672 VDD.n1302 279.885
R49 VDD.t958 VDD.n1698 263.567
R50 VDD.t958 VDD.n1659 235.143
R51 VDD.t958 VDD.n1684 209.303
R52 VDD.t909 VDD.t900 188.018
R53 VDD.t900 VDD.t912 188.018
R54 VDD.t912 VDD.t902 188.018
R55 VDD.t902 VDD.t1052 188.018
R56 VDD.t1052 VDD.t904 188.018
R57 VDD.t904 VDD.t59 188.018
R58 VDD.t59 VDD.t57 188.018
R59 VDD.t160 VDD.n1785 184.496
R60 VDD.n1685 VDD.t946 180.88
R61 VDD.t25 VDD.t832 180.213
R62 VDD.t351 VDD.t25 180.213
R63 VDD.t343 VDD.t348 180.213
R64 VDD.t348 VDD.t27 180.213
R65 VDD.t27 VDD.t294 180.213
R66 VDD.t294 VDD.t23 180.213
R67 VDD.n1976 VDD.t573 164.593
R68 VDD.n1786 VDD.t343 161.661
R69 VDD.n1337 VDD.t943 160.7
R70 VDD.n1496 VDD.t970 160.284
R71 VDD.n1937 VDD.n1815 132.696
R72 VDD.n1898 VDD.n1897 132.696
R73 VDD.n134 VDD.n133 132.696
R74 VDD.n74 VDD.n73 132.696
R75 VDD.n1437 VDD.n1436 132.696
R76 VDD.n1428 VDD.n1427 132.696
R77 VDD.n1362 VDD.n1361 132.696
R78 VDD.n446 VDD.n403 132.696
R79 VDD.n428 VDD.n427 132.696
R80 VDD.n867 VDD.n866 132.696
R81 VDD.n957 VDD.n956 132.696
R82 VDD.n1376 VDD.n1373 132.696
R83 VDD.n1785 VDD.t418 131.784
R84 VDD.n1937 VDD.n1936 128.591
R85 VDD.t567 VDD.n1935 128.591
R86 VDD.n1935 VDD.n1816 128.591
R87 VDD.n1930 VDD.n1929 128.591
R88 VDD.n1899 VDD.n1898 128.591
R89 VDD.t767 VDD.n1884 128.591
R90 VDD.n1904 VDD.n1884 128.591
R91 VDD.n1909 VDD.n1905 128.591
R92 VDD.n143 VDD.n142 128.591
R93 VDD.n141 VDD.n123 128.591
R94 VDD.t377 VDD.n123 128.591
R95 VDD.n135 VDD.n134 128.591
R96 VDD.n64 VDD.n63 128.591
R97 VDD.n66 VDD.n65 128.591
R98 VDD.n65 VDD.t763 128.591
R99 VDD.n73 VDD.n72 128.591
R100 VDD.n1438 VDD.n1437 128.591
R101 VDD.t517 VDD.n347 128.591
R102 VDD.n1444 VDD.n347 128.591
R103 VDD.n1446 VDD.n1445 128.591
R104 VDD.n1427 VDD.n1400 128.591
R105 VDD.n1410 VDD.t407 128.591
R106 VDD.n1420 VDD.n1410 128.591
R107 VDD.n1419 VDD.n1418 128.591
R108 VDD.n1354 VDD.n374 128.591
R109 VDD.n1356 VDD.n1355 128.591
R110 VDD.n1356 VDD.t166 128.591
R111 VDD.n1361 VDD.n365 128.591
R112 VDD.n460 VDD.n394 128.591
R113 VDD.n454 VDD.n453 128.591
R114 VDD.n453 VDD.t308 128.591
R115 VDD.n452 VDD.n403 128.591
R116 VDD.n437 VDD.n436 128.591
R117 VDD.n435 VDD.n412 128.591
R118 VDD.t758 VDD.n412 128.591
R119 VDD.n428 VDD.n423 128.591
R120 VDD.n858 VDD.n857 128.591
R121 VDD.n864 VDD.n841 128.591
R122 VDD.t745 VDD.n864 128.591
R123 VDD.n867 VDD.n865 128.591
R124 VDD.n964 VDD.n942 128.591
R125 VDD.t543 VDD.n942 128.591
R126 VDD.n957 VDD.n950 128.591
R127 VDD.n1372 VDD.n1371 128.591
R128 VDD.n1385 VDD.n1384 128.591
R129 VDD.n1384 VDD.t126 128.591
R130 VDD.n1383 VDD.n1373 128.591
R131 VDD.n1690 VDD.t946 126.615
R132 VDD.n1839 VDD.t67 124.386
R133 VDD.n1869 VDD.t329 124.386
R134 VDD.n162 VDD.t267 124.386
R135 VDD.n102 VDD.t43 124.386
R136 VDD.t85 VDD.n1798 123.376
R137 VDD.t165 VDD.n1853 123.376
R138 VDD.t288 VDD.n27 123.376
R139 VDD.t62 VDD.n84 123.376
R140 VDD.n1833 VDD.t68 122.1
R141 VDD.n1863 VDD.t332 122.1
R142 VDD.n156 VDD.t130 122.1
R143 VDD.n96 VDD.t42 122.1
R144 VDD.n2085 VDD.t548 122.1
R145 VDD.n2595 VDD.t367 122.1
R146 VDD.n1799 VDD.t430 121.091
R147 VDD.n1854 VDD.t163 121.091
R148 VDD.n28 VDD.t562 121.091
R149 VDD.n85 VDD.t72 121.091
R150 VDD.t411 VDD.n2113 121.091
R151 VDD.t336 VDD.n2657 121.091
R152 VDD.n1969 VDD.t345 120.213
R153 VDD.n1804 VDD.t215 119.317
R154 VDD.n1859 VDD.t164 119.317
R155 VDD.n33 VDD.t549 119.317
R156 VDD.n90 VDD.t65 119.317
R157 VDD.n1842 VDD.t894 118.308
R158 VDD.n1872 VDD.t331 118.308
R159 VDD.n165 VDD.t540 118.308
R160 VDD.n105 VDD.t41 118.308
R161 VDD.t1085 VDD.t1050 118.191
R162 VDD.t1029 VDD.t897 118.191
R163 VDD.t354 VDD.t1048 118.191
R164 VDD.t564 VDD.n1814 118.061
R165 VDD.n1887 VDD.t775 118.061
R166 VDD.n128 VDD.t284 118.061
R167 VDD.t881 VDD.n43 118.061
R168 VDD.n1391 VDD.t534 118.061
R169 VDD.n1429 VDD.t404 118.061
R170 VDD.n1363 VDD.t103 118.061
R171 VDD.t319 VDD.n445 118.061
R172 VDD.t753 VDD.n426 118.061
R173 VDD.t541 VDD.n955 118.061
R174 VDD.n1377 VDD.t124 118.061
R175 VDD.n1976 VDD.t155 117.567
R176 VDD.n1803 VDD.t709 117.053
R177 VDD.n1858 VDD.t153 117.053
R178 VDD.n32 VDD.t0 117.053
R179 VDD.n89 VDD.t1035 117.053
R180 VDD.t364 VDD.n1831 116.044
R181 VDD.t330 VDD.n1861 116.044
R182 VDD.t665 VDD.n154 116.044
R183 VDD.t40 VDD.n94 116.044
R184 VDD.t279 VDD.n2083 116.044
R185 VDD.t370 VDD.n2593 116.044
R186 VDD.t29 VDD.t339 113.275
R187 VDD.t182 VDD.t340 113.275
R188 VDD.t837 VDD.t1086 113.275
R189 VDD.n1930 VDD.t891 110.808
R190 VDD.n1905 VDD.t769 110.808
R191 VDD.n142 VDD.t286 110.808
R192 VDD.t888 VDD.n64 110.808
R193 VDD.n1445 VDD.t525 110.808
R194 VDD.t390 VDD.n1419 110.808
R195 VDD.t88 VDD.n1354 110.808
R196 VDD.t301 VDD.n394 110.808
R197 VDD.n436 VDD.t761 110.808
R198 VDD.n858 VDD.t743 110.808
R199 VDD.t122 VDD.n1372 110.808
R200 VDD.n965 VDD.t327 109.439
R201 VDD.t358 VDD.t909 108.948
R202 VDD.n1832 VDD.t364 105.954
R203 VDD.n1862 VDD.t330 105.954
R204 VDD.n155 VDD.t665 105.954
R205 VDD.n95 VDD.t40 105.954
R206 VDD.n2084 VDD.t279 105.954
R207 VDD.n2594 VDD.t370 105.954
R208 VDD.t709 VDD.n1802 104.945
R209 VDD.t153 VDD.n1857 104.945
R210 VDD.t0 VDD.n31 104.945
R211 VDD.t1035 VDD.n88 104.945
R212 VDD.n2114 VDD.t414 104.945
R213 VDD.n2658 VDD.t334 104.945
R214 VDD.t832 VDD.t1092 104.418
R215 VDD.n1521 VDD.n321 102.362
R216 VDD.n1266 VDD.n1256 102.362
R217 VDD.n1802 VDD.t430 100.909
R218 VDD.n1857 VDD.t163 100.909
R219 VDD.n31 VDD.t562 100.909
R220 VDD.n88 VDD.t72 100.909
R221 VDD.n2114 VDD.t411 100.909
R222 VDD.n2658 VDD.t336 100.909
R223 VDD.t68 VDD.n1832 99.8996
R224 VDD.t332 VDD.n1862 99.8996
R225 VDD.t130 VDD.n155 99.8996
R226 VDD.t42 VDD.n95 99.8996
R227 VDD.t548 VDD.n2084 99.8996
R228 VDD.t367 VDD.n2594 99.8996
R229 VDD.n1520 VDD.t666 99.5009
R230 VDD.t672 VDD.n471 99.0846
R231 VDD.n873 VDD.t748 98.4957
R232 VDD.t958 VDD.n1650 98.1917
R233 VDD.n1448 VDD.t513 97.5562
R234 VDD.n1969 VDD.t341 96.809
R235 VDD.t206 VDD.n1928 95.9239
R236 VDD.t380 VDD.n111 95.9239
R237 VDD.n48 VDD.t69 95.9239
R238 VDD.t9 VDD.n856 95.9239
R239 VDD.t773 VDD.n1908 95.9239
R240 VDD.n1413 VDD.t396 95.9239
R241 VDD.n1347 VDD.t100 95.9239
R242 VDD.n461 VDD.t322 95.9239
R243 VDD.n440 VDD.t755 95.9239
R244 VDD.n1368 VDD.t503 95.9239
R245 VDD.t965 VDD.n282 92.4235
R246 VDD.t955 VDD.n1288 92.4235
R247 VDD.n1831 VDD.t894 89.8088
R248 VDD.n1861 VDD.t331 89.8088
R249 VDD.n154 VDD.t540 89.8088
R250 VDD.n94 VDD.t41 89.8088
R251 VDD.n2083 VDD.t422 89.8088
R252 VDD.n2593 VDD.t119 89.8088
R253 VDD.t215 VDD.n1803 88.7997
R254 VDD.t164 VDD.n1858 88.7997
R255 VDD.t549 VDD.n32 88.7997
R256 VDD.t65 VDD.n89 88.7997
R257 VDD.n2116 VDD.t412 88.7997
R258 VDD.n2660 VDD.t335 88.7997
R259 VDD.n564 VDD.n563 86.1787
R260 VDD.t461 VDD.t464 85.5351
R261 VDD.t482 VDD.t452 85.5351
R262 VDD.t106 VDD.t605 85.5351
R263 VDD.t825 VDD.t80 85.5351
R264 VDD.t807 VDD.t12 85.5351
R265 VDD.t576 VDD.n931 84.8158
R266 VDD.n1799 VDD.t85 84.7634
R267 VDD.n1854 VDD.t165 84.7634
R268 VDD.n28 VDD.t288 84.7634
R269 VDD.n85 VDD.t62 84.7634
R270 VDD.n2113 VDD.t413 84.7634
R271 VDD.n2657 VDD.t333 84.7634
R272 VDD.t67 VDD.n1833 83.7543
R273 VDD.t329 VDD.n1863 83.7543
R274 VDD.t267 VDD.n156 83.7543
R275 VDD.t43 VDD.n96 83.7543
R276 VDD.n2085 VDD.t563 83.7543
R277 VDD.n2595 VDD.t117 83.7543
R278 VDD.n2288 VDD.t431 75.0529
R279 VDD.n2504 VDD.t223 75.0529
R280 VDD.n976 VDD.n932 73.8719
R281 VDD.t958 VDD.n1658 72.3519
R282 VDD.t1050 VDD.t1029 70.1759
R283 VDD.t897 VDD.t354 70.1759
R284 VDD.t1048 VDD.t358 70.1759
R285 VDD.n1508 VDD.t666 70.1759
R286 VDD.n1303 VDD.t672 70.1759
R287 VDD.n2291 VDD.t446 67.925
R288 VDD.n2507 VDD.t679 67.925
R289 VDD.t340 VDD.t29 67.2571
R290 VDD.t1086 VDD.t182 67.2571
R291 VDD.t1092 VDD.t837 67.2571
R292 VDD.t973 VDD.n323 67.252
R293 VDD.t978 VDD.n473 67.252
R294 VDD.n795 VDD.n779 66.348
R295 VDD.n796 VDD.n795 64.296
R296 VDD.t17 VDD.n775 64.296
R297 VDD.n812 VDD.n775 64.296
R298 VDD.n816 VDD.n815 64.296
R299 VDD.n822 VDD.n821 64.296
R300 VDD.n2294 VDD.t497 62.055
R301 VDD.n2510 VDD.t208 62.055
R302 VDD.n683 VDD.t44 61.8854
R303 VDD.n895 VDD.t194 60.8721
R304 VDD.n682 VDD.t105 60.7435
R305 VDD.t204 VDD.n897 59.702
R306 VDD.t132 VDD.n679 59.0509
R307 VDD.t192 VDD.n899 58.9084
R308 VDD.t201 VDD.n900 57.7119
R309 VDD.n789 VDD.t6 57.456
R310 VDD.n602 VDD.n601 56.5021
R311 VDD.n664 VDD.n663 56.5021
R312 VDD.n2297 VDD.t494 56.185
R313 VDD.n2513 VDD.t32 56.185
R314 VDD.n815 VDD.t750 55.4041
R315 VDD.n1717 VDD.n1643 54.5384
R316 VDD.n1034 VDD.n1033 54.5384
R317 VDD.n734 VDD.n593 53.3521
R318 VDD.n720 VDD.n641 53.3521
R319 VDD.n717 VDD.n716 53.3521
R320 VDD.n662 VDD.n658 53.3521
R321 VDD.n680 VDD.t132 52.7113
R322 VDD.n1573 VDD.n1572 52.4568
R323 VDD.n1188 VDD.n493 52.0405
R324 VDD.n901 VDD.t201 51.7418
R325 VDD.t452 VDD.n2300 51.1535
R326 VDD.n2539 VDD.t246 51.1535
R327 VDD.t978 VDD.n471 50.3542
R328 VDD.n1520 VDD.t973 49.9381
R329 VDD.n901 VDD.t204 49.7517
R330 VDD.n680 VDD.t105 49.6993
R331 VDD.t361 VDD.t109 49.5054
R332 VDD.t109 VDD.t272 49.5054
R333 VDD.t272 VDD.t131 49.5054
R334 VDD.t22 VDD.t243 49.5054
R335 VDD.t217 VDD.t22 49.5054
R336 VDD.t154 VDD.t217 49.5054
R337 VDD.t31 VDD.t154 49.5054
R338 VDD.t31 VDD.t4 49.5054
R339 VDD.t4 VDD.t242 49.5054
R340 VDD.t242 VDD.t133 49.5054
R341 VDD.t133 VDD.t262 49.5054
R342 VDD.t5 VDD.t376 49.5054
R343 VDD.t269 VDD.t5 49.5054
R344 VDD.t21 VDD.t269 49.5054
R345 VDD.n2028 VDD.t423 47.9334
R346 VDD.n2285 VDD.t458 46.9607
R347 VDD.n2315 VDD.t444 46.9607
R348 VDD.n2501 VDD.t686 46.9607
R349 VDD.n2558 VDD.t38 46.9607
R350 VDD.n2326 VDD.t488 46.5414
R351 VDD.n2569 VDD.t810 46.5414
R352 VDD.t52 VDD.n708 46.5121
R353 VDD.n821 VDD.t19 46.5121
R354 VDD.n1580 VDD.n270 45.7957
R355 VDD.n1579 VDD.n271 45.7957
R356 VDD.n1586 VDD.n266 45.7957
R357 VDD.t386 VDD.n1587 45.7957
R358 VDD.n1606 VDD.n242 45.7957
R359 VDD.n1597 VDD.n1594 45.7957
R360 VDD.n1762 VDD.n176 45.7957
R361 VDD.n184 VDD.n183 45.7957
R362 VDD.n1755 VDD.n1754 45.7957
R363 VDD.n191 VDD.n185 45.7957
R364 VDD.n1748 VDD.n192 45.7957
R365 VDD.n203 VDD.n202 45.7957
R366 VDD.n211 VDD.n204 45.7957
R367 VDD.n1732 VDD.n210 45.7957
R368 VDD.n1633 VDD.n1632 45.7957
R369 VDD.n1641 VDD.n1634 45.7957
R370 VDD.n1718 VDD.n1642 45.7957
R371 VDD.n1041 VDD.n554 45.7957
R372 VDD.n1040 VDD.n556 45.7957
R373 VDD.n1049 VDD.n1048 45.7957
R374 VDD.n1058 VDD.n542 45.7957
R375 VDD.n547 VDD.n546 45.7957
R376 VDD.n1122 VDD.n533 45.7957
R377 VDD.n1132 VDD.n1131 45.7957
R378 VDD.n1139 VDD.n521 45.7957
R379 VDD.n1138 VDD.n522 45.7957
R380 VDD.n1146 VDD.n517 45.7957
R381 VDD.n1156 VDD.n511 45.7957
R382 VDD.n1163 VDD.n507 45.7957
R383 VDD.n1173 VDD.n501 45.7957
R384 VDD.n1179 VDD.n497 45.7957
R385 VDD.n1181 VDD.n1180 45.7957
R386 VDD.n1189 VDD.n492 45.7957
R387 VDD.n2025 VDD.t426 45.5368
R388 VDD.n1172 VDD.t171 45.3794
R389 VDD.n721 VDD.n640 45.1441
R390 VDD.n2343 VDD.t482 44.0257
R391 VDD.n2586 VDD.t74 44.0257
R392 VDD.n1700 VDD.t958 43.9281
R393 VDD.n900 VDD.t192 43.7816
R394 VDD.t519 VDD.n1724 43.2978
R395 VDD.n555 VDD.t174 42.8814
R396 VDD.t93 VDD.n1147 42.8814
R397 VDD.n1761 VDD.t383 42.4651
R398 VDD.n897 VDD.t194 41.7915
R399 VDD.n0 VDD.t361 41.7644
R400 VDD.n2173 VDD.t21 41.7644
R401 VDD.t44 VDD.n682 41.6672
R402 VDD.n2343 VDD.t449 41.5099
R403 VDD.n2586 VDD.t249 41.5099
R404 VDD.n1929 VDD.t206 39.6722
R405 VDD.n1909 VDD.t773 39.6722
R406 VDD.n143 VDD.t380 39.6722
R407 VDD.n63 VDD.t69 39.6722
R408 VDD.n1446 VDD.t513 39.6722
R409 VDD.n1418 VDD.t396 39.6722
R410 VDD.t100 VDD.n374 39.6722
R411 VDD.t322 VDD.n460 39.6722
R412 VDD.n437 VDD.t755 39.6722
R413 VDD.n647 VDD.n646 39.6722
R414 VDD.n857 VDD.t9 39.6722
R415 VDD.n1371 VDD.t503 39.6722
R416 VDD.n2156 VDD.t555 39.6722
R417 VDD.n2619 VDD.t115 39.6722
R418 VDD.n1571 VDD.n275 39.5509
R419 VDD.n1279 VDD.n487 39.5509
R420 VDD.n2326 VDD.t106 38.9942
R421 VDD.n2569 VDD.t807 38.9942
R422 VDD.n2285 VDD.t455 38.5749
R423 VDD.n2315 VDD.t437 38.5749
R424 VDD.n2501 VDD.t78 38.5749
R425 VDD.n2558 VDD.t147 38.5749
R426 VDD.n1559 VDD.n282 38.3019
R427 VDD.n544 VDD.t95 38.3019
R428 VDD.n1288 VDD.n479 38.3019
R429 VDD.n1510 VDD.n322 37.9019
R430 VDD.n1302 VDD.n1301 37.9019
R431 VDD.n212 VDD.t409 37.8856
R432 VDD.n201 VDD.t388 36.2203
R433 VDD.n1498 VDD.n330 35.8675
R434 VDD.n1310 VDD.n1309 35.8675
R435 VDD.n532 VDD.t90 35.804
R436 VDD.n619 VDD.t185 35.5682
R437 VDD.n2300 VDD.t213 34.382
R438 VDD.n2539 VDD.t211 34.382
R439 VDD.n2032 VDD.t429 33.5535
R440 VDD.n978 VDD.t576 32.8322
R441 VDD.n1470 VDD.n1469 32.7175
R442 VDD.n1339 VDD.n378 32.7175
R443 VDD.n1559 VDD.n283 32.0571
R444 VDD.n1280 VDD.n479 32.0571
R445 VDD.n562 VDD.t983 31.6415
R446 VDD.n1593 VDD.t393 31.6408
R447 VDD.n1165 VDD.t180 31.2245
R448 VDD.n2071 VDD.t915 31.1569
R449 VDD.n283 VDD.n275 30.8082
R450 VDD.n1280 VDD.n1279 30.8082
R451 VDD.n2312 VDD.t472 30.1892
R452 VDD.n2555 VDD.t723 30.1892
R453 VDD.n966 VDD.n932 30.0963
R454 VDD.n2323 VDD.t467 29.7699
R455 VDD.n2566 VDD.t14 29.7699
R456 VDD.n2297 VDD.t506 29.3506
R457 VDD.n2513 VDD.t141 29.3506
R458 VDD.n930 VDD.n921 28.8809
R459 VDD.t176 VDD.n512 28.7266
R460 VDD.n1599 VDD.t402 28.3102
R461 VDD.n1529 VDD.n1528 28.1746
R462 VDD.n1274 VDD.n489 28.1746
R463 VDD.n679 VDD.t49 24.6667
R464 VDD.n977 VDD.n976 24.6243
R465 VDD.n1123 VDD.t98 24.147
R466 VDD.n1740 VDD.t398 23.7307
R467 VDD.n2294 VDD.t603 23.4806
R468 VDD.n2510 VDD.t684 23.4806
R469 VDD.n1828 VDD.n1826 23.2342
R470 VDD.n1912 VDD.n1879 23.2342
R471 VDD.n1454 VDD.n1453 23.2342
R472 VDD.n2159 VDD.n2154 23.2342
R473 VDD.n2622 VDD.n2617 23.2342
R474 VDD.n120 VDD.n119 23.1442
R475 VDD.n60 VDD.n58 23.1442
R476 VDD.t398 VDD.n1739 22.0654
R477 VDD.t891 VDD.n1816 21.8883
R478 VDD.t769 VDD.n1904 21.8883
R479 VDD.t286 VDD.n141 21.8883
R480 VDD.n66 VDD.t888 21.8883
R481 VDD.t525 VDD.n1444 21.8883
R482 VDD.n1420 VDD.t390 21.8883
R483 VDD.n1355 VDD.t88 21.8883
R484 VDD.n454 VDD.t301 21.8883
R485 VDD.t761 VDD.n435 21.8883
R486 VDD.t743 VDD.n841 21.8883
R487 VDD.t327 VDD.n964 21.8883
R488 VDD.n1385 VDD.t122 21.8883
R489 VDD.n2144 VDD.t276 21.8883
R490 VDD.n2635 VDD.t281 21.8883
R491 VDD.n545 VDD.t98 21.6491
R492 VDD.n2316 VDD.t134 21.3841
R493 VDD.n2559 VDD.t143 21.3841
R494 VDD.n1032 VDD.t934 21.2328
R495 VDD.n2305 VDD.t598 20.9649
R496 VDD.n2548 VDD.t76 20.9649
R497 VDD.t958 VDD.n1699 20.8165
R498 VDD.n120 VDD.n114 20.4798
R499 VDD.n60 VDD.n53 20.4798
R500 VDD.n1455 VDD.n1454 20.395
R501 VDD.n1828 VDD.n1827 20.3898
R502 VDD.n1912 VDD.n1880 20.3898
R503 VDD.n2159 VDD.n2155 20.3898
R504 VDD.n2622 VDD.n2618 20.3898
R505 VDD.n816 VDD.t19 19.8363
R506 VDD.t995 VDD.n1571 19.5675
R507 VDD.t937 VDD.n487 19.5675
R508 VDD.n874 VDD.n873 19.0194
R509 VDD.n1786 VDD.t351 18.5517
R510 VDD.n2291 VDD.t440 17.6106
R511 VDD.n2507 VDD.t854 17.6106
R512 VDD.n995 VDD.n559 17.5593
R513 VDD.t402 VDD.n1598 17.4859
R514 VDD.n1155 VDD.t176 17.0696
R515 VDD.n1673 VDD.n1666 16.2393
R516 VDD.t180 VDD.n1164 14.5717
R517 VDD.n1605 VDD.t393 14.1554
R518 VDD.n1815 VDD.t564 13.6804
R519 VDD.n1897 VDD.t775 13.6804
R520 VDD.n133 VDD.t284 13.6804
R521 VDD.n74 VDD.t881 13.6804
R522 VDD.n1436 VDD.t534 13.6804
R523 VDD.t404 VDD.n1428 13.6804
R524 VDD.t103 VDD.n1362 13.6804
R525 VDD.n446 VDD.t319 13.6804
R526 VDD.n427 VDD.t753 13.6804
R527 VDD.n646 VDD.n594 13.6804
R528 VDD.n866 VDD.t748 13.6804
R529 VDD.n956 VDD.t541 13.6804
R530 VDD.t124 VDD.n1376 13.6804
R531 VDD.n2125 VDD.t273 13.6804
R532 VDD.n2646 VDD.t110 13.6804
R533 VDD.n1570 VDD.n269 13.33
R534 VDD.n1187 VDD.n486 13.2637
R535 VDD.n2309 VDD.t442 12.9984
R536 VDD.n2552 VDD.t244 12.9984
R537 VDD.n618 VDD.n593 12.9964
R538 VDD.n709 VDD.n662 12.9964
R539 VDD.n2320 VDD.t136 12.5791
R540 VDD.n2563 VDD.t145 12.5791
R541 VDD.n1574 VDD.n274 11.6418
R542 VDD.n1278 VDD.n488 11.6418
R543 VDD.n1518 VDD.n325 11.2373
R544 VDD.n1570 VDD.n276 11.2079
R545 VDD.n1281 VDD.n486 11.2079
R546 VDD.n1290 VDD.n477 11.1709
R547 VDD.n1027 VDD.n560 11.094
R548 VDD.n619 VDD.n617 10.9444
R549 VDD.n721 VDD.n720 10.9444
R550 VDD.t46 VDD.n641 10.9444
R551 VDD.n716 VDD.n658 10.9444
R552 VDD.n708 VDD.n663 10.9444
R553 VDD.n812 VDD.t750 10.9444
R554 VDD.n1928 VDD.n1927 10.7369
R555 VDD.n147 VDD.n111 10.7369
R556 VDD.n49 VDD.n48 10.7369
R557 VDD.n1908 VDD.n1907 10.7362
R558 VDD.n856 VDD.n855 10.723
R559 VDD.n1414 VDD.n1413 10.7223
R560 VDD.n1347 VDD.n1346 10.7223
R561 VDD.n462 VDD.n461 10.7223
R562 VDD.n441 VDD.n440 10.7223
R563 VDD.n1368 VDD.n1367 10.7223
R564 VDD.n2288 VDD.t461 10.4827
R565 VDD.n2504 VDD.t825 10.4827
R566 VDD.n1666 VDD.n1640 10.4784
R567 VDD.n1035 VDD.n559 10.4784
R568 VDD.n1716 VDD.n1645 10.3407
R569 VDD.n1031 VDD.n553 10.3407
R570 VDD.n1539 VDD.n1538 10.2548
R571 VDD.n1239 VDD.n1238 10.2548
R572 VDD.n1027 VDD.n564 10.2279
R573 VDD.n1689 VDD.n1648 10.1865
R574 VDD.n1027 VDD.n1026 10.1865
R575 VDD.n1573 VDD.t940 9.99217
R576 VDD.n1130 VDD.t90 9.99217
R577 VDD.n493 VDD.t949 9.99217
R578 VDD.n1712 VDD.n1645 9.86137
R579 VDD.n1031 VDD.n560 9.86137
R580 VDD.n1529 VDD.n274 9.78981
R581 VDD.n1278 VDD.n489 9.78981
R582 VDD.n2175 VDD.n2174 9.6468
R583 VDD.n1747 VDD.t388 9.57585
R584 VDD.n578 VDD.t933 9.55982
R585 VDD.n574 VDD.t992 9.55982
R586 VDD.n570 VDD.t980 9.55982
R587 VDD.n566 VDD.t982 9.55982
R588 VDD.n1668 VDD.t987 9.51591
R589 VDD.n1662 VDD.t957 9.51591
R590 VDD.n1655 VDD.t962 9.51591
R591 VDD.n1687 VDD.t945 9.51591
R592 VDD.n2049 VDD.n2048 9.4133
R593 VDD.n1719 VDD.n1640 9.28471
R594 VDD.n1035 VDD.n557 9.28471
R595 VDD.n1574 VDD.n272 9.24507
R596 VDD.n1190 VDD.n488 9.17659
R597 VDD.n924 VDD.n921 9.16567
R598 VDD.n2 VDD.n1 9.09976
R599 VDD.n481 VDD.n480 9.08576
R600 VDD.n2073 VDD.t916 9.02932
R601 VDD.n1564 VDD.n1563 9.01945
R602 VDD.n734 VDD.n733 8.89243
R603 VDD.n2051 VDD.n2050 8.82188
R604 VDD.n1472 VDD.n334 8.80618
R605 VDD.n2049 VDD.t695 8.79795
R606 VDD.n1557 VDD.n290 8.78029
R607 VDD.n1552 VDD.n1551 8.78029
R608 VDD.n1226 VDD.n1225 8.78029
R609 VDD.n1223 VDD.n1212 8.78029
R610 VDD.n1547 VDD.n1546 8.71327
R611 VDD.n1534 VDD.n1533 8.71327
R612 VDD.n1244 VDD.n1243 8.71327
R613 VDD.n1231 VDD.n1230 8.71327
R614 VDD.n2073 VDD.t917 8.6005
R615 VDD.n2074 VDD.t918 8.6005
R616 VDD.n2075 VDD.t919 8.6005
R617 VDD.n1505 VDD.n328 8.59141
R618 VDD.n1509 VDD.n328 8.59141
R619 VDD.n1511 VDD.n1509 8.59141
R620 VDD.n1513 VDD.n1511 8.59141
R621 VDD.n1513 VDD.n324 8.59141
R622 VDD.n1518 VDD.n324 8.59141
R623 VDD.n1466 VDD.n1457 8.59141
R624 VDD.n1466 VDD.n1459 8.59141
R625 VDD.n1459 VDD.n319 8.59141
R626 VDD.n1523 VDD.n319 8.59141
R627 VDD.n1524 VDD.n1523 8.59141
R628 VDD.n1272 VDD.n1250 8.59141
R629 VDD.n1267 VDD.n1250 8.59141
R630 VDD.n1267 VDD.n1255 8.59141
R631 VDD.n1263 VDD.n1255 8.59141
R632 VDD.n1263 VDD.n1258 8.59141
R633 VDD.n1290 VDD.n474 8.59141
R634 VDD.n1299 VDD.n474 8.59141
R635 VDD.n1299 VDD.n472 8.59141
R636 VDD.n472 VDD.n470 8.59141
R637 VDD.n1305 VDD.n470 8.59141
R638 VDD.n1306 VDD.n1305 8.59141
R639 VDD.n1938 VDD.n1808 8.488
R640 VDD.n1934 VDD.n1809 8.488
R641 VDD.n1931 VDD.n1817 8.488
R642 VDD.n1821 VDD.n1820 8.488
R643 VDD.n1896 VDD.n1885 8.488
R644 VDD.n1901 VDD.n1900 8.488
R645 VDD.n1903 VDD.n1882 8.488
R646 VDD.n1910 VDD.n1883 8.488
R647 VDD.n145 VDD.n144 8.488
R648 VDD.n140 VDD.n122 8.488
R649 VDD.n136 VDD.n124 8.488
R650 VDD.n132 VDD.n127 8.488
R651 VDD.n62 VDD.n47 8.488
R652 VDD.n67 VDD.n46 8.488
R653 VDD.n71 VDD.n44 8.488
R654 VDD.n75 VDD.n42 8.488
R655 VDD.n1435 VDD.n1390 8.488
R656 VDD.n1439 VDD.n348 8.488
R657 VDD.n1443 VDD.n346 8.488
R658 VDD.n1426 VDD.n1399 8.488
R659 VDD.n1402 VDD.n1401 8.488
R660 VDD.n1421 VDD.n1409 8.488
R661 VDD.n1417 VDD.n1411 8.488
R662 VDD.n1348 VDD.n375 8.488
R663 VDD.n1353 VDD.n373 8.488
R664 VDD.n1357 VDD.n366 8.488
R665 VDD.n1360 VDD.n364 8.488
R666 VDD.n459 VDD.n393 8.488
R667 VDD.n455 VDD.n395 8.488
R668 VDD.n451 VDD.n402 8.488
R669 VDD.n447 VDD.n404 8.488
R670 VDD.n439 VDD.n438 8.488
R671 VDD.n434 VDD.n410 8.488
R672 VDD.n420 VDD.n413 8.488
R673 VDD.n429 VDD.n422 8.488
R674 VDD.n719 VDD.n718 8.488
R675 VDD.n710 VDD.n656 8.488
R676 VDD.n735 VDD.n591 8.488
R677 VDD.n722 VDD.n592 8.488
R678 VDD.n715 VDD.n639 8.488
R679 VDD.n707 VDD.n659 8.488
R680 VDD.n850 VDD.n849 8.488
R681 VDD.n859 VDD.n842 8.488
R682 VDD.n863 VDD.n840 8.488
R683 VDD.n868 VDD.n838 8.488
R684 VDD.n794 VDD.n793 8.488
R685 VDD.n810 VDD.n776 8.488
R686 VDD.n811 VDD.n772 8.488
R687 VDD.n817 VDD.n769 8.488
R688 VDD.n791 VDD.n778 8.488
R689 VDD.n797 VDD.n773 8.488
R690 VDD.n814 VDD.n813 8.488
R691 VDD.n820 VDD.n770 8.488
R692 VDD.n959 VDD.n943 8.488
R693 VDD.n958 VDD.n951 8.488
R694 VDD.n1370 VDD.n1369 8.488
R695 VDD.n1382 VDD.n357 8.488
R696 VDD.n1381 VDD.n1374 8.488
R697 VDD.n1469 VDD.n1468 8.48682
R698 VDD.n1528 VDD.n314 8.48682
R699 VDD.n1274 VDD.n1273 8.48682
R700 VDD.n1257 VDD.n378 8.48682
R701 VDD.n963 VDD.n941 8.4005
R702 VDD.n1475 VDD.n334 8.37664
R703 VDD.n1699 VDD.n1643 8.32689
R704 VDD.n1034 VDD.n1032 8.32689
R705 VDD.n1506 VDD.n330 8.31689
R706 VDD.n1309 VDD.n468 8.31615
R707 VDD.n1814 VDD.n1808 8.2255
R708 VDD.n1938 VDD.n1809 8.2255
R709 VDD.n1934 VDD.n1817 8.2255
R710 VDD.n1931 VDD.n1820 8.2255
R711 VDD.n1896 VDD.n1887 8.2255
R712 VDD.n1900 VDD.n1885 8.2255
R713 VDD.n1903 VDD.n1901 8.2255
R714 VDD.n1910 VDD.n1882 8.2255
R715 VDD.n144 VDD.n122 8.2255
R716 VDD.n140 VDD.n124 8.2255
R717 VDD.n136 VDD.n127 8.2255
R718 VDD.n132 VDD.n128 8.2255
R719 VDD.n62 VDD.n46 8.2255
R720 VDD.n67 VDD.n44 8.2255
R721 VDD.n71 VDD.n42 8.2255
R722 VDD.n75 VDD.n43 8.2255
R723 VDD.n1435 VDD.n1391 8.2255
R724 VDD.n1439 VDD.n1390 8.2255
R725 VDD.n1443 VDD.n348 8.2255
R726 VDD.n1447 VDD.n346 8.2255
R727 VDD.n1429 VDD.n1399 8.2255
R728 VDD.n1426 VDD.n1401 8.2255
R729 VDD.n1421 VDD.n1402 8.2255
R730 VDD.n1417 VDD.n1409 8.2255
R731 VDD.n1353 VDD.n375 8.2255
R732 VDD.n1357 VDD.n373 8.2255
R733 VDD.n1360 VDD.n366 8.2255
R734 VDD.n1363 VDD.n364 8.2255
R735 VDD.n459 VDD.n395 8.2255
R736 VDD.n455 VDD.n402 8.2255
R737 VDD.n451 VDD.n404 8.2255
R738 VDD.n447 VDD.n445 8.2255
R739 VDD.n438 VDD.n410 8.2255
R740 VDD.n434 VDD.n413 8.2255
R741 VDD.n429 VDD.n420 8.2255
R742 VDD.n426 VDD.n422 8.2255
R743 VDD.n718 VDD.n656 8.2255
R744 VDD.n710 VDD.n661 8.2255
R745 VDD.n611 VDD.n591 8.2255
R746 VDD.n735 VDD.n592 8.2255
R747 VDD.n722 VDD.n639 8.2255
R748 VDD.n715 VDD.n659 8.2255
R749 VDD.n707 VDD.n664 8.2255
R750 VDD.n859 VDD.n849 8.2255
R751 VDD.n863 VDD.n842 8.2255
R752 VDD.n868 VDD.n840 8.2255
R753 VDD.n793 VDD.n780 8.2255
R754 VDD.n794 VDD.n776 8.2255
R755 VDD.n811 VDD.n810 8.2255
R756 VDD.n817 VDD.n772 8.2255
R757 VDD.n823 VDD.n769 8.2255
R758 VDD.n791 VDD.n790 8.2255
R759 VDD.n797 VDD.n778 8.2255
R760 VDD.n813 VDD.n773 8.2255
R761 VDD.n814 VDD.n770 8.2255
R762 VDD.n820 VDD.n768 8.2255
R763 VDD.n963 VDD.n943 8.2255
R764 VDD.n959 VDD.n958 8.2255
R765 VDD.n955 VDD.n951 8.2255
R766 VDD.n1370 VDD.n356 8.2255
R767 VDD.n1386 VDD.n357 8.2255
R768 VDD.n1382 VDD.n1381 8.2255
R769 VDD.n1377 VDD.n1374 8.2255
R770 VDD.n2145 VDD.n2143 8.2255
R771 VDD.n2638 VDD.n2636 8.2255
R772 VDD.n648 VDD.n640 8.20843
R773 VDD.n931 VDD.n930 8.20843
R774 VDD.n1578 VDD.n272 8.14941
R775 VDD.n1578 VDD.n265 8.14941
R776 VDD.n1588 VDD.n265 8.14941
R777 VDD.n1588 VDD.n243 8.14941
R778 VDD.n1604 VDD.n243 8.14941
R779 VDD.n1604 VDD.n244 8.14941
R780 VDD.n1600 VDD.n244 8.14941
R781 VDD.n1600 VDD.n177 8.14941
R782 VDD.n1760 VDD.n177 8.14941
R783 VDD.n1760 VDD.n178 8.14941
R784 VDD.n1756 VDD.n178 8.14941
R785 VDD.n1756 VDD.n181 8.14941
R786 VDD.n193 VDD.n181 8.14941
R787 VDD.n1746 VDD.n193 8.14941
R788 VDD.n1746 VDD.n194 8.14941
R789 VDD.n1741 VDD.n194 8.14941
R790 VDD.n1741 VDD.n200 8.14941
R791 VDD.n213 VDD.n200 8.14941
R792 VDD.n1731 VDD.n213 8.14941
R793 VDD.n1731 VDD.n214 8.14941
R794 VDD.n1726 VDD.n214 8.14941
R795 VDD.n1726 VDD.n1631 8.14941
R796 VDD.n1644 VDD.n1631 8.14941
R797 VDD.n1716 VDD.n1644 8.14941
R798 VDD.n1042 VDD.n553 8.14941
R799 VDD.n1042 VDD.n551 8.14941
R800 VDD.n1046 VDD.n551 8.14941
R801 VDD.n1046 VDD.n540 8.14941
R802 VDD.n1059 VDD.n540 8.14941
R803 VDD.n1059 VDD.n541 8.14941
R804 VDD.n541 VDD.n531 8.14941
R805 VDD.n1124 VDD.n531 8.14941
R806 VDD.n1124 VDD.n526 8.14941
R807 VDD.n1129 VDD.n526 8.14941
R808 VDD.n1129 VDD.n520 8.14941
R809 VDD.n1140 VDD.n520 8.14941
R810 VDD.n1140 VDD.n518 8.14941
R811 VDD.n1145 VDD.n518 8.14941
R812 VDD.n1145 VDD.n510 8.14941
R813 VDD.n1157 VDD.n510 8.14941
R814 VDD.n1157 VDD.n508 8.14941
R815 VDD.n1162 VDD.n508 8.14941
R816 VDD.n1162 VDD.n500 8.14941
R817 VDD.n1174 VDD.n500 8.14941
R818 VDD.n1174 VDD.n498 8.14941
R819 VDD.n1178 VDD.n498 8.14941
R820 VDD.n1178 VDD.n491 8.14941
R821 VDD.n1190 VDD.n491 8.14941
R822 VDD.n732 VDD.n621 7.963
R823 VDD.n1733 VDD.t409 7.91057
R824 VDD.n1581 VDD.n269 7.89208
R825 VDD.n1581 VDD.n267 7.89208
R826 VDD.n1585 VDD.n267 7.89208
R827 VDD.n1585 VDD.n240 7.89208
R828 VDD.n1607 VDD.n240 7.89208
R829 VDD.n1607 VDD.n241 7.89208
R830 VDD.n1596 VDD.n241 7.89208
R831 VDD.n1596 VDD.n174 7.89208
R832 VDD.n1763 VDD.n174 7.89208
R833 VDD.n1763 VDD.n175 7.89208
R834 VDD.n186 VDD.n175 7.89208
R835 VDD.n1753 VDD.n186 7.89208
R836 VDD.n1753 VDD.n187 7.89208
R837 VDD.n1749 VDD.n187 7.89208
R838 VDD.n1749 VDD.n190 7.89208
R839 VDD.n205 VDD.n190 7.89208
R840 VDD.n1738 VDD.n205 7.89208
R841 VDD.n1738 VDD.n206 7.89208
R842 VDD.n1734 VDD.n206 7.89208
R843 VDD.n1734 VDD.n209 7.89208
R844 VDD.n1635 VDD.n209 7.89208
R845 VDD.n1723 VDD.n1635 7.89208
R846 VDD.n1723 VDD.n1636 7.89208
R847 VDD.n1719 VDD.n1636 7.89208
R848 VDD.n1039 VDD.n557 7.89208
R849 VDD.n1039 VDD.n550 7.89208
R850 VDD.n1050 VDD.n550 7.89208
R851 VDD.n1050 VDD.n543 7.89208
R852 VDD.n1056 VDD.n543 7.89208
R853 VDD.n1056 VDD.n548 7.89208
R854 VDD.n548 VDD.n534 7.89208
R855 VDD.n1121 VDD.n534 7.89208
R856 VDD.n1121 VDD.n525 7.89208
R857 VDD.n1133 VDD.n525 7.89208
R858 VDD.n1133 VDD.n523 7.89208
R859 VDD.n1137 VDD.n523 7.89208
R860 VDD.n1137 VDD.n516 7.89208
R861 VDD.n1149 VDD.n516 7.89208
R862 VDD.n1149 VDD.n513 7.89208
R863 VDD.n1154 VDD.n513 7.89208
R864 VDD.n1154 VDD.n506 7.89208
R865 VDD.n1166 VDD.n506 7.89208
R866 VDD.n1166 VDD.n503 7.89208
R867 VDD.n1171 VDD.n503 7.89208
R868 VDD.n1171 VDD.n496 7.89208
R869 VDD.n1182 VDD.n496 7.89208
R870 VDD.n1182 VDD.n494 7.89208
R871 VDD.n1187 VDD.n494 7.89208
R872 VDD.n615 VDD.n602 7.613
R873 VDD.n2061 VDD.t427 7.58462
R874 VDD.n2062 VDD.t694 7.58462
R875 VDD.n2043 VDD.n2027 7.58109
R876 VDD.n979 VDD.n919 7.5255
R877 VDD.n649 VDD.n648 7.52444
R878 VDD.n1057 VDD.t95 7.49426
R879 VDD.n1543 VDD.n1542 7.30582
R880 VDD.n1235 VDD.n1234 7.30582
R881 VDD.n1283 VDD.n485 7.30582
R882 VDD.n2030 VDD.t428 7.19043
R883 VDD.n2067 VDD.t1 7.19043
R884 VDD.n719 VDD.n655 7.1755
R885 VDD.n872 VDD.n838 7.1755
R886 VDD.n621 VDD.n620 7.088
R887 VDD.n1672 VDD.n1664 7.00704
R888 VDD.n1676 VDD.n1664 7.00704
R889 VDD.n1677 VDD.n1676 7.00704
R890 VDD.n1678 VDD.n1677 7.00704
R891 VDD.n1678 VDD.n1661 7.00704
R892 VDD.n1683 VDD.n1661 7.00704
R893 VDD.n1683 VDD.n1652 7.00704
R894 VDD.n1706 VDD.n1652 7.00704
R895 VDD.n1706 VDD.n1653 7.00704
R896 VDD.n1701 VDD.n1653 7.00704
R897 VDD.n1701 VDD.n1657 7.00704
R898 VDD.n1696 VDD.n1657 7.00704
R899 VDD.n1696 VDD.n1686 7.00704
R900 VDD.n1691 VDD.n1686 7.00704
R901 VDD.n1691 VDD.n1689 7.00704
R902 VDD.n1024 VDD.n565 7.00704
R903 VDD.n1019 VDD.n1018 7.00704
R904 VDD.n1016 VDD.n569 7.00704
R905 VDD.n1011 VDD.n1010 7.00704
R906 VDD.n1008 VDD.n573 7.00704
R907 VDD.n1003 VDD.n1002 7.00704
R908 VDD.n1000 VDD.n577 7.00704
R909 VDD.n2000 VDD.t58 6.94485
R910 VDD.n310 VDD.n308 6.94485
R911 VDD.n1196 VDD.t798 6.94485
R912 VDD.n1957 VDD.t293 6.94485
R913 VDD.t185 VDD.n618 6.84045
R914 VDD.n709 VDD.t52 6.84045
R915 VDD.t6 VDD.n779 6.84045
R916 VDD.n978 VDD.n977 6.84045
R917 VDD.n1812 VDD.n1811 6.70224
R918 VDD.n1890 VDD.n1888 6.70224
R919 VDD.n129 VDD.t285 6.70224
R920 VDD.n40 VDD.t882 6.70224
R921 VDD.n1397 VDD.n1396 6.70224
R922 VDD.n1394 VDD.n1392 6.70224
R923 VDD.n424 VDD.t778 6.70224
R924 VDD.n405 VDD.t714 6.70224
R925 VDD.n666 VDD.t53 6.70224
R926 VDD.n605 VDD.n604 6.70224
R927 VDD.n835 VDD.t749 6.70224
R928 VDD.n783 VDD.n781 6.70224
R929 VDD.n786 VDD.n785 6.70224
R930 VDD.n953 VDD.t542 6.70224
R931 VDD.n362 VDD.t104 6.70224
R932 VDD.n1375 VDD.t129 6.70224
R933 VDD.n2122 VDD.n2120 6.70224
R934 VDD.n2643 VDD.n2642 6.70224
R935 VDD.n344 VDD.t740 6.68489
R936 VDD.n465 VDD.n463 6.68371
R937 VDD.n2009 VDD.t572 6.68267
R938 VDD.n1827 VDD.t1063 6.65503
R939 VDD.n1880 VDD.t1024 6.65503
R940 VDD.n114 VDD.n112 6.65503
R941 VDD.n53 VDD.n51 6.65503
R942 VDD.n1412 VDD.t622 6.65503
R943 VDD.n408 VDD.n406 6.65503
R944 VDD.n694 VDD.t676 6.65503
R945 VDD.n608 VDD.n606 6.65503
R946 VDD.n853 VDD.n851 6.65503
R947 VDD.n750 VDD.t1112 6.65503
R948 VDD.n927 VDD.n925 6.65503
R949 VDD.n1345 VDD.n1344 6.65503
R950 VDD.n361 VDD.n360 6.65503
R951 VDD.n2155 VDD.t584 6.65503
R952 VDD.n2618 VDD.t539 6.65503
R953 VDD.n828 VDD.t1008 6.64521
R954 VDD.n1562 VDD.n1561 6.63561
R955 VDD.n1972 VDD.n1971 6.61305
R956 VDD.n2013 VDD.n2012 6.58706
R957 VDD.n1283 VDD.n1282 6.56859
R958 VDD.n1970 VDD.t1088 6.54616
R959 VDD.n1970 VDD.t342 6.54616
R960 VDD.n1782 VDD.t338 6.52811
R961 VDD.n5 VDD.n4 6.52199
R962 VDD.n1973 VDD.n1968 6.51831
R963 VDD.t956 VDD.n1251 6.50716
R964 VDD.n316 VDD.t966 6.50716
R965 VDD.n2057 VDD.n2056 6.44895
R966 VDD.n1209 VDD.t936 6.43191
R967 VDD.n1195 VDD.t975 6.43124
R968 VDD.n1218 VDD.t948 6.4298
R969 VDD.n291 VDD.t939 6.42961
R970 VDD.n299 VDD.t994 6.37351
R971 VDD.n1199 VDD.t989 6.37275
R972 VDD.n306 VDD.t951 6.37256
R973 VDD.n312 VDD.t960 6.37217
R974 VDD.n326 VDD.t972 6.36486
R975 VDD.n1501 VDD.t985 6.36262
R976 VDD.n1461 VDD.t969 6.36128
R977 VDD.n1294 VDD.t967 6.30795
R978 VDD.n475 VDD.t977 6.30193
R979 VDD.n2016 VDD.n1976 6.3005
R980 VDD.n1841 VDD.n1831 6.3005
R981 VDD VDD.n1832 6.3005
R982 VDD.n1840 VDD.n1833 6.3005
R983 VDD.n1800 VDD.n1799 6.3005
R984 VDD.n1802 VDD.n1801 6.3005
R985 VDD.n1803 VDD.n1792 6.3005
R986 VDD.n1870 VDD.n1863 6.3005
R987 VDD VDD.n1862 6.3005
R988 VDD.n1871 VDD.n1861 6.3005
R989 VDD.n1858 VDD.n1847 6.3005
R990 VDD.n1857 VDD.n1856 6.3005
R991 VDD.n1855 VDD.n1854 6.3005
R992 VDD.n164 VDD.n154 6.3005
R993 VDD VDD.n155 6.3005
R994 VDD.n163 VDD.n156 6.3005
R995 VDD.n32 VDD.n21 6.3005
R996 VDD.n31 VDD.n30 6.3005
R997 VDD.n29 VDD.n28 6.3005
R998 VDD.n104 VDD.n94 6.3005
R999 VDD VDD.n95 6.3005
R1000 VDD.n103 VDD.n96 6.3005
R1001 VDD.n89 VDD.n78 6.3005
R1002 VDD.n88 VDD.n87 6.3005
R1003 VDD.n86 VDD.n85 6.3005
R1004 VDD.n645 VDD.n644 6.3005
R1005 VDD.n646 VDD.n645 6.3005
R1006 VDD.n651 VDD.n650 6.3005
R1007 VDD.n650 VDD.n649 6.3005
R1008 VDD.n615 VDD.n614 6.3005
R1009 VDD.n616 VDD.n615 6.3005
R1010 VDD.n872 VDD.n871 6.3005
R1011 VDD.n873 VDD.n872 6.3005
R1012 VDD.n923 VDD.n922 6.3005
R1013 VDD.n941 VDD.n940 6.3005
R1014 VDD.n965 VDD.n941 6.3005
R1015 VDD.n980 VDD.n979 6.3005
R1016 VDD.n979 VDD.n978 6.3005
R1017 VDD.n920 VDD.n918 6.3005
R1018 VDD.n977 VDD.n920 6.3005
R1019 VDD.n968 VDD.n967 6.3005
R1020 VDD.n967 VDD.n966 6.3005
R1021 VDD.n1785 VDD.n1784 6.3005
R1022 VDD VDD.n1786 6.3005
R1023 VDD.n2072 VDD.n2071 6.3005
R1024 VDD.n2070 VDD.n2069 6.3005
R1025 VDD.n2068 VDD.n2067 6.3005
R1026 VDD.n2065 VDD.n2064 6.3005
R1027 VDD.n2026 VDD.n2025 6.3005
R1028 VDD.n2035 VDD.n2034 6.3005
R1029 VDD.n2036 VDD.n2033 6.3005
R1030 VDD.n2037 VDD.n2032 6.3005
R1031 VDD.n2038 VDD.n2031 6.3005
R1032 VDD.n2039 VDD.n2030 6.3005
R1033 VDD.n2040 VDD.n2029 6.3005
R1034 VDD.n2041 VDD.n2028 6.3005
R1035 VDD.n2092 VDD.n2085 6.3005
R1036 VDD VDD.n2084 6.3005
R1037 VDD.n2093 VDD.n2083 6.3005
R1038 VDD.n2117 VDD.n2116 6.3005
R1039 VDD.n2115 VDD.n2114 6.3005
R1040 VDD.n2113 VDD.n2112 6.3005
R1041 VDD.n2603 VDD.n2593 6.3005
R1042 VDD VDD.n2594 6.3005
R1043 VDD.n2602 VDD.n2595 6.3005
R1044 VDD.n2657 VDD.n2656 6.3005
R1045 VDD.n2659 VDD.n2658 6.3005
R1046 VDD.n2661 VDD.n2660 6.3005
R1047 VDD.n2344 VDD.n2343 6.3005
R1048 VDD.n2347 VDD.n2300 6.3005
R1049 VDD.n2342 VDD.n2305 6.3005
R1050 VDD.n2340 VDD.n2308 6.3005
R1051 VDD.n2339 VDD.n2309 6.3005
R1052 VDD.n2337 VDD.n2312 6.3005
R1053 VDD.n2335 VDD.n2315 6.3005
R1054 VDD.n2334 VDD.n2316 6.3005
R1055 VDD.n2332 VDD.n2319 6.3005
R1056 VDD.n2331 VDD.n2320 6.3005
R1057 VDD.n2329 VDD.n2323 6.3005
R1058 VDD.n2327 VDD.n2326 6.3005
R1059 VDD.n2292 VDD.n2291 6.3005
R1060 VDD.n2289 VDD.n2288 6.3005
R1061 VDD.n2286 VDD.n2285 6.3005
R1062 VDD.n2354 VDD.n2297 6.3005
R1063 VDD.n2295 VDD.n2294 6.3005
R1064 VDD.n2587 VDD.n2586 6.3005
R1065 VDD.n2585 VDD.n2548 6.3005
R1066 VDD.n2583 VDD.n2551 6.3005
R1067 VDD.n2582 VDD.n2552 6.3005
R1068 VDD.n2580 VDD.n2555 6.3005
R1069 VDD.n2578 VDD.n2558 6.3005
R1070 VDD.n2577 VDD.n2559 6.3005
R1071 VDD.n2575 VDD.n2562 6.3005
R1072 VDD.n2574 VDD.n2563 6.3005
R1073 VDD.n2572 VDD.n2566 6.3005
R1074 VDD.n2570 VDD.n2569 6.3005
R1075 VDD.n2511 VDD.n2510 6.3005
R1076 VDD.n2508 VDD.n2507 6.3005
R1077 VDD.n2505 VDD.n2504 6.3005
R1078 VDD.n2502 VDD.n2501 6.3005
R1079 VDD.n2540 VDD.n2539 6.3005
R1080 VDD.n2514 VDD.n2513 6.3005
R1081 VDD.n1259 VDD.t942 6.29942
R1082 VDD.n316 VDD.t964 6.29685
R1083 VDD.n2052 VDD.t691 6.27989
R1084 VDD.n828 VDD.t1000 6.26273
R1085 VDD.n465 VDD.n464 6.24167
R1086 VDD.n2000 VDD.t906 6.2405
R1087 VDD.n1827 VDD.t207 6.2405
R1088 VDD.n1812 VDD.n1810 6.2405
R1089 VDD.n1890 VDD.n1889 6.2405
R1090 VDD.n1880 VDD.t774 6.2405
R1091 VDD.n114 VDD.n113 6.2405
R1092 VDD.n129 VDD.t841 6.2405
R1093 VDD.n53 VDD.n52 6.2405
R1094 VDD.n40 VDD.t1078 6.2405
R1095 VDD.n310 VDD.n309 6.2405
R1096 VDD.n344 VDD.t514 6.2405
R1097 VDD.n1412 VDD.t397 6.2405
R1098 VDD.n1397 VDD.n1395 6.2405
R1099 VDD.n1394 VDD.n1393 6.2405
R1100 VDD.n1252 VDD.t956 6.2405
R1101 VDD.n1196 VDD.t785 6.2405
R1102 VDD.n424 VDD.t754 6.2405
R1103 VDD.n408 VDD.n407 6.2405
R1104 VDD.n405 VDD.t320 6.2405
R1105 VDD.n666 VDD.t56 6.2405
R1106 VDD.n694 VDD.t674 6.2405
R1107 VDD.n608 VDD.n607 6.2405
R1108 VDD.n605 VDD.n603 6.2405
R1109 VDD.n853 VDD.n852 6.2405
R1110 VDD.n835 VDD.t1108 6.2405
R1111 VDD.n786 VDD.n784 6.2405
R1112 VDD.n783 VDD.n782 6.2405
R1113 VDD.n750 VDD.t20 6.2405
R1114 VDD.n953 VDD.t1042 6.2405
R1115 VDD.n927 VDD.n926 6.2405
R1116 VDD.n1345 VDD.n1343 6.2405
R1117 VDD.n362 VDD.t179 6.2405
R1118 VDD.n361 VDD.n359 6.2405
R1119 VDD.n1375 VDD.t125 6.2405
R1120 VDD.t966 VDD.n315 6.2405
R1121 VDD.n1957 VDD.t24 6.2405
R1122 VDD.n2122 VDD.n2121 6.2405
R1123 VDD.n2155 VDD.t556 6.2405
R1124 VDD.n2618 VDD.t116 6.2405
R1125 VDD.n2643 VDD.n2641 6.2405
R1126 VDD.n1251 VDD.t954 6.23498
R1127 VDD.n616 VDD.n601 6.15645
R1128 VDD.n1282 VDD.n480 6.03524
R1129 VDD.n1563 VDD.n1562 5.96892
R1130 VDD.n1837 VDD.n1836 5.77744
R1131 VDD.n1795 VDD.t216 5.77744
R1132 VDD.n1867 VDD.n1866 5.77744
R1133 VDD.n1850 VDD.t1043 5.77744
R1134 VDD.n160 VDD.n159 5.77744
R1135 VDD.n24 VDD.t827 5.77744
R1136 VDD.n100 VDD.n99 5.77744
R1137 VDD.n81 VDD.t66 5.77744
R1138 VDD.n687 VDD.n686 5.77744
R1139 VDD.n676 VDD.n675 5.77744
R1140 VDD.n892 VDD.t252 5.77744
R1141 VDD.n887 VDD.t193 5.77744
R1142 VDD.n2089 VDD.n2088 5.77744
R1143 VDD.n2108 VDD.t1023 5.77744
R1144 VDD.n2599 VDD.n2598 5.77744
R1145 VDD.n2652 VDD.t1105 5.77744
R1146 VDD.n650 VDD.n645 5.7755
R1147 VDD.n2022 VDD.n2021 5.7405
R1148 VDD.n875 VDD.n874 5.2962
R1149 VDD.n2024 VDD.n2018 5.2005
R1150 VDD.n2023 VDD.n2019 5.2005
R1151 VDD.n2022 VDD.n2020 5.2005
R1152 VDD.n1562 VDD.n276 5.10682
R1153 VDD.n1282 VDD.n1281 5.10682
R1154 VDD.n1838 VDD.t1059 5.07264
R1155 VDD.n1797 VDD.n1796 5.07264
R1156 VDD.n1868 VDD.t766 5.07264
R1157 VDD.n1852 VDD.n1851 5.07264
R1158 VDD.n161 VDD.t268 5.07264
R1159 VDD.n26 VDD.n25 5.07264
R1160 VDD.n101 VDD.t417 5.07264
R1161 VDD.n83 VDD.n82 5.07264
R1162 VDD.n677 VDD.t45 5.07264
R1163 VDD.n894 VDD.n893 5.07264
R1164 VDD.n889 VDD.n888 5.07264
R1165 VDD.n2090 VDD.t585 5.07264
R1166 VDD.n2110 VDD.n2109 5.07264
R1167 VDD.n2600 VDD.t118 5.07264
R1168 VDD.n2654 VDD.n2653 5.07264
R1169 VDD.n1709 VDD.t946 4.99634
R1170 VDD.n691 VDD.t558 4.79075
R1171 VDD.n617 VDD.n616 4.78846
R1172 VDD.n975 VDD.n933 4.7255
R1173 VDD.n108 VDD.n107 4.57581
R1174 VDD.n702 VDD.n669 4.52789
R1175 VDD.n971 VDD.n970 4.52785
R1176 VDD.n600 VDD.n585 4.51855
R1177 VDD.n875 VDD.n834 4.5152
R1178 VDD.n726 VDD.n725 4.5084
R1179 VDD.n764 VDD.n763 4.50489
R1180 VDD.n1926 VDD.n1925 4.50248
R1181 VDD.n1918 VDD.n1917 4.50129
R1182 VDD.n1892 VDD.n1791 4.50129
R1183 VDD.n1914 VDD.n1845 4.5005
R1184 VDD.n1906 VDD.n1844 4.5005
R1185 VDD.n1924 VDD.n1923 4.5005
R1186 VDD.n1920 VDD.n1919 4.5005
R1187 VDD.n1942 VDD.n1941 4.5005
R1188 VDD.n151 VDD.n150 4.5005
R1189 VDD.n109 VDD.n37 4.5005
R1190 VDD.n110 VDD.n36 4.5005
R1191 VDD.n108 VDD.n38 4.5005
R1192 VDD.n149 VDD.n148 4.5005
R1193 VDD.n20 VDD.n18 4.5005
R1194 VDD.n168 VDD.n167 4.5005
R1195 VDD.n701 VDD.n700 4.5005
R1196 VDD.n699 VDD.n670 4.5005
R1197 VDD.n695 VDD.n668 4.5005
R1198 VDD.n669 VDD.n660 4.5005
R1199 VDD.n705 VDD.n665 4.5005
R1200 VDD.n654 VDD.n653 4.5005
R1201 VDD.n655 VDD.n654 4.5005
R1202 VDD.n655 VDD.n640 4.5005
R1203 VDD.n738 VDD.n737 4.5005
R1204 VDD.n731 VDD.n730 4.5005
R1205 VDD.n732 VDD.n731 4.5005
R1206 VDD.n733 VDD.n732 4.5005
R1207 VDD.n620 VDD.n600 4.5005
R1208 VDD.n620 VDD.n619 4.5005
R1209 VDD.n597 VDD.n587 4.5005
R1210 VDD.n741 VDD.n740 4.5005
R1211 VDD.n727 VDD.n624 4.5005
R1212 VDD.n729 VDD.n728 4.5005
R1213 VDD.n739 VDD.n586 4.5005
R1214 VDD.n879 VDD.n833 4.5005
R1215 VDD.n880 VDD.n832 4.5005
R1216 VDD.n764 VDD.n753 4.5005
R1217 VDD.n767 VDD.n754 4.5005
R1218 VDD.n825 VDD.n824 4.5005
R1219 VDD.n826 VDD.n825 4.5005
R1220 VDD.n767 VDD.n766 4.5005
R1221 VDD.n760 VDD.n755 4.5005
R1222 VDD.n757 VDD.n756 4.5005
R1223 VDD.n748 VDD.n747 4.5005
R1224 VDD.n762 VDD.n761 4.5005
R1225 VDD.n912 VDD.n911 4.5005
R1226 VDD.n906 VDD.n905 4.5005
R1227 VDD.n907 VDD.n745 4.5005
R1228 VDD.n910 VDD.n744 4.5005
R1229 VDD.n970 VDD.n969 4.5005
R1230 VDD.n969 VDD.n933 4.5005
R1231 VDD.n933 VDD.n932 4.5005
R1232 VDD.n939 VDD.n936 4.5005
R1233 VDD.n974 VDD.n973 4.5005
R1234 VDD.n975 VDD.n974 4.5005
R1235 VDD.n976 VDD.n975 4.5005
R1236 VDD.n938 VDD.n935 4.5005
R1237 VDD.n937 VDD.n916 4.5005
R1238 VDD.n982 VDD.n981 4.5005
R1239 VDD.n986 VDD.n985 4.5005
R1240 VDD.n923 VDD.n583 4.5005
R1241 VDD.n923 VDD.n919 4.5005
R1242 VDD.n931 VDD.n919 4.5005
R1243 VDD.n584 VDD.n582 4.5005
R1244 VDD.n1770 VDD.n1769 4.5005
R1245 VDD.n1962 VDD.n1774 4.5005
R1246 VDD.n1963 VDD.n1773 4.5005
R1247 VDD.n1960 VDD.n1789 4.5005
R1248 VDD.n1959 VDD.n1944 4.5005
R1249 VDD.n2060 VDD.n2059 4.5005
R1250 VDD.n2327 VDD.t729 4.21354
R1251 VDD.n2570 VDD.t13 4.21354
R1252 VDD.n2308 VDD.t138 4.19337
R1253 VDD.n2319 VDD.t434 4.19337
R1254 VDD.n2551 VDD.t220 4.19337
R1255 VDD.n2562 VDD.t35 4.19337
R1256 VDD.n1936 VDD.t567 4.10447
R1257 VDD.n1899 VDD.t767 4.10447
R1258 VDD.n135 VDD.t377 4.10447
R1259 VDD.n72 VDD.t763 4.10447
R1260 VDD.n1438 VDD.t517 4.10447
R1261 VDD.t407 VDD.n1400 4.10447
R1262 VDD.t166 VDD.n365 4.10447
R1263 VDD.t308 VDD.n452 4.10447
R1264 VDD.n423 VDD.t758 4.10447
R1265 VDD.n865 VDD.t745 4.10447
R1266 VDD.n950 VDD.t543 4.10447
R1267 VDD.t126 VDD.n1383 4.10447
R1268 VDD.n2138 VDD.t270 4.10447
R1269 VDD.n2628 VDD.t113 4.10447
R1270 VDD.n14 VDD.n13 3.99669
R1271 VDD.n1981 VDD.n1980 3.99665
R1272 VDD.n13 VDD.t1087 3.80383
R1273 VDD.n1980 VDD.t355 3.80304
R1274 VDD.n1572 VDD.n270 3.74738
R1275 VDD.n1580 VDD.n1579 3.74738
R1276 VDD.n271 VDD.n266 3.74738
R1277 VDD.t386 VDD.n1586 3.74738
R1278 VDD.n1587 VDD.n242 3.74738
R1279 VDD.n1606 VDD.n1605 3.74738
R1280 VDD.n1594 VDD.n1593 3.74738
R1281 VDD.n1599 VDD.n1597 3.74738
R1282 VDD.n1598 VDD.n176 3.74738
R1283 VDD.n1762 VDD.n1761 3.74738
R1284 VDD.n183 VDD.n182 3.74738
R1285 VDD.n1755 VDD.n184 3.74738
R1286 VDD.n1754 VDD.n185 3.74738
R1287 VDD.n192 VDD.n191 3.74738
R1288 VDD.n1748 VDD.n1747 3.74738
R1289 VDD.n202 VDD.n201 3.74738
R1290 VDD.n1740 VDD.n203 3.74738
R1291 VDD.n1739 VDD.n204 3.74738
R1292 VDD.n212 VDD.n211 3.74738
R1293 VDD.n1733 VDD.n1732 3.74738
R1294 VDD.n1632 VDD.n210 3.74738
R1295 VDD.n1725 VDD.n1633 3.74738
R1296 VDD.n1724 VDD.n1634 3.74738
R1297 VDD.n1642 VDD.n1641 3.74738
R1298 VDD.n1718 VDD.n1717 3.74738
R1299 VDD.n1033 VDD.n554 3.74738
R1300 VDD.n1041 VDD.n1040 3.74738
R1301 VDD.n556 VDD.n555 3.74738
R1302 VDD.n1049 VDD.n1047 3.74738
R1303 VDD.n1048 VDD.n542 3.74738
R1304 VDD.n1058 VDD.n1057 3.74738
R1305 VDD.n547 VDD.n544 3.74738
R1306 VDD.n546 VDD.n545 3.74738
R1307 VDD.n1123 VDD.n1122 3.74738
R1308 VDD.n533 VDD.n532 3.74738
R1309 VDD.n1132 VDD.n1130 3.74738
R1310 VDD.n1131 VDD.n521 3.74738
R1311 VDD.n1139 VDD.n1138 3.74738
R1312 VDD.n522 VDD.n517 3.74738
R1313 VDD.n1148 VDD.n1146 3.74738
R1314 VDD.n1147 VDD.n511 3.74738
R1315 VDD.n1156 VDD.n1155 3.74738
R1316 VDD.n512 VDD.n507 3.74738
R1317 VDD.n1165 VDD.n1163 3.74738
R1318 VDD.n1164 VDD.n501 3.74738
R1319 VDD.n1173 VDD.n1172 3.74738
R1320 VDD.n502 VDD.n497 3.74738
R1321 VDD.n1181 VDD.n1179 3.74738
R1322 VDD.n1180 VDD.n492 3.74738
R1323 VDD.n1189 VDD.n1188 3.74738
R1324 VDD.n1990 VDD.t905 3.6405
R1325 VDD.n1990 VDD.n1989 3.6405
R1326 VDD.n1992 VDD.t1091 3.6405
R1327 VDD.n1992 VDD.n1991 3.6405
R1328 VDD.n1994 VDD.t1090 3.6405
R1329 VDD.n1994 VDD.n1993 3.6405
R1330 VDD.n1996 VDD.t1089 3.6405
R1331 VDD.n1996 VDD.n1995 3.6405
R1332 VDD.n1988 VDD.t903 3.6405
R1333 VDD.n1988 VDD.n1987 3.6405
R1334 VDD.n1985 VDD.t901 3.6405
R1335 VDD.n1985 VDD.n1984 3.6405
R1336 VDD.n1983 VDD.t1049 3.6405
R1337 VDD.n1983 VDD.n1982 3.6405
R1338 VDD.n1978 VDD.t1051 3.6405
R1339 VDD.n1978 VDD.n1977 3.6405
R1340 VDD.n2011 VDD.t156 3.6405
R1341 VDD.n2011 VDD.n2010 3.6405
R1342 VDD.n1823 VDD.t1062 3.6405
R1343 VDD.n1823 VDD.n1822 3.6405
R1344 VDD.n1825 VDD.t568 3.6405
R1345 VDD.n1825 VDD.n1824 3.6405
R1346 VDD.n1878 VDD.t768 3.6405
R1347 VDD.n1878 VDD.n1877 3.6405
R1348 VDD.n1876 VDD.t1032 3.6405
R1349 VDD.n1876 VDD.n1875 3.6405
R1350 VDD.n118 VDD.t287 3.6405
R1351 VDD.n118 VDD.n117 3.6405
R1352 VDD.n116 VDD.t842 3.6405
R1353 VDD.n116 VDD.n115 3.6405
R1354 VDD.n57 VDD.t1077 3.6405
R1355 VDD.n57 VDD.n56 3.6405
R1356 VDD.n55 VDD.t889 3.6405
R1357 VDD.n55 VDD.n54 3.6405
R1358 VDD.n1612 VDD.t529 3.6405
R1359 VDD.n1612 VDD.n1611 3.6405
R1360 VDD.n249 VDD.t510 3.6405
R1361 VDD.n249 VDD.n248 3.6405
R1362 VDD.n233 VDD.t528 3.6405
R1363 VDD.n233 VDD.n232 3.6405
R1364 VDD.n230 VDD.t614 3.6405
R1365 VDD.n230 VDD.n229 3.6405
R1366 VDD.n227 VDD.t522 3.6405
R1367 VDD.n227 VDD.n226 3.6405
R1368 VDD.n255 VDD.t734 3.6405
R1369 VDD.n255 VDD.n254 3.6405
R1370 VDD.n1624 VDD.t410 3.6405
R1371 VDD.n1624 VDD.n1623 3.6405
R1372 VDD.n1621 VDD.t630 3.6405
R1373 VDD.n1621 VDD.n1620 3.6405
R1374 VDD.n218 VDD.t735 3.6405
R1375 VDD.n218 VDD.n217 3.6405
R1376 VDD.n297 VDD.t861 3.6405
R1377 VDD.n297 VDD.n296 3.6405
R1378 VDD.n295 VDD.t795 3.6405
R1379 VDD.n295 VDD.n294 3.6405
R1380 VDD.n303 VDD.t790 3.6405
R1381 VDD.n303 VDD.n302 3.6405
R1382 VDD.n301 VDD.t860 3.6405
R1383 VDD.n301 VDD.n300 3.6405
R1384 VDD.n1452 VDD.t524 3.6405
R1385 VDD.n1452 VDD.n1451 3.6405
R1386 VDD.n1450 VDD.t518 3.6405
R1387 VDD.n1450 VDD.n1449 3.6405
R1388 VDD.n1404 VDD.t408 3.6405
R1389 VDD.n1404 VDD.n1403 3.6405
R1390 VDD.n1406 VDD.t629 3.6405
R1391 VDD.n1406 VDD.n1405 3.6405
R1392 VDD.n1214 VDD.t791 3.6405
R1393 VDD.n1214 VDD.n1213 3.6405
R1394 VDD.n1216 VDD.t673 3.6405
R1395 VDD.n1216 VDD.n1215 3.6405
R1396 VDD.n1203 VDD.t794 3.6405
R1397 VDD.n1203 VDD.n1202 3.6405
R1398 VDD.n1205 VDD.t859 3.6405
R1399 VDD.n1205 VDD.n1204 3.6405
R1400 VDD.n1093 VDD.t713 3.6405
R1401 VDD.n1093 VDD.n1092 3.6405
R1402 VDD.n1079 VDD.t715 3.6405
R1403 VDD.n1079 VDD.n1078 3.6405
R1404 VDD.n1081 VDD.t314 3.6405
R1405 VDD.n1081 VDD.n1080 3.6405
R1406 VDD.n1087 VDD.t181 3.6405
R1407 VDD.n1087 VDD.n1086 3.6405
R1408 VDD.n1090 VDD.t239 3.6405
R1409 VDD.n1090 VDD.n1089 3.6405
R1410 VDD.n1075 VDD.t720 3.6405
R1411 VDD.n1075 VDD.n1074 3.6405
R1412 VDD.n418 VDD.t762 3.6405
R1413 VDD.n418 VDD.n417 3.6405
R1414 VDD.n416 VDD.t781 3.6405
R1415 VDD.n416 VDD.n415 3.6405
R1416 VDD.n399 VDD.t717 3.6405
R1417 VDD.n399 VDD.n398 3.6405
R1418 VDD.n397 VDD.t302 3.6405
R1419 VDD.n397 VDD.n396 3.6405
R1420 VDD.n1083 VDD.t94 3.6405
R1421 VDD.n1083 VDD.n1082 3.6405
R1422 VDD.n1116 VDD.t237 3.6405
R1423 VDD.n1116 VDD.n1115 3.6405
R1424 VDD.n1111 VDD.t311 3.6405
R1425 VDD.n1111 VDD.n1110 3.6405
R1426 VDD.n1105 VDD.t228 3.6405
R1427 VDD.n1105 VDD.n1104 3.6405
R1428 VDD.n1108 VDD.t175 3.6405
R1429 VDD.n1108 VDD.n1107 3.6405
R1430 VDD.n1063 VDD.t716 3.6405
R1431 VDD.n1063 VDD.n1062 3.6405
R1432 VDD.n1068 VDD.t321 3.6405
R1433 VDD.n1068 VDD.n1067 3.6405
R1434 VDD.n1066 VDD.t307 3.6405
R1435 VDD.n1066 VDD.n1065 3.6405
R1436 VDD.n1072 VDD.t152 3.6405
R1437 VDD.n1072 VDD.n1071 3.6405
R1438 VDD.n528 VDD.t99 3.6405
R1439 VDD.n528 VDD.n527 3.6405
R1440 VDD.n631 VDD.t189 3.6405
R1441 VDD.n631 VDD.n630 3.6405
R1442 VDD.n629 VDD.t200 3.6405
R1443 VDD.n629 VDD.n628 3.6405
R1444 VDD.n635 VDD.t675 3.6405
R1445 VDD.n635 VDD.n634 3.6405
R1446 VDD.n637 VDD.t257 3.6405
R1447 VDD.n637 VDD.n636 3.6405
R1448 VDD.n846 VDD.t1107 3.6405
R1449 VDD.n846 VDD.n845 3.6405
R1450 VDD.n844 VDD.t744 3.6405
R1451 VDD.n844 VDD.n843 3.6405
R1452 VDD.n805 VDD.t999 3.6405
R1453 VDD.n805 VDD.n804 3.6405
R1454 VDD.n807 VDD.t1003 3.6405
R1455 VDD.n807 VDD.n806 3.6405
R1456 VDD.n802 VDD.t18 3.6405
R1457 VDD.n802 VDD.n801 3.6405
R1458 VDD.n800 VDD.t1111 3.6405
R1459 VDD.n800 VDD.n799 3.6405
R1460 VDD.n947 VDD.t579 3.6405
R1461 VDD.n947 VDD.n946 3.6405
R1462 VDD.n945 VDD.t328 3.6405
R1463 VDD.n945 VDD.n944 3.6405
R1464 VDD.n368 VDD.t89 3.6405
R1465 VDD.n368 VDD.n367 3.6405
R1466 VDD.n370 VDD.t238 3.6405
R1467 VDD.n370 VDD.n369 3.6405
R1468 VDD.n351 VDD.t123 3.6405
R1469 VDD.n351 VDD.n350 3.6405
R1470 VDD.n353 VDD.t885 3.6405
R1471 VDD.n353 VDD.n352 3.6405
R1472 VDD.n1628 VDD.t537 3.6405
R1473 VDD.n1628 VDD.n1627 3.6405
R1474 VDD.n197 VDD.t389 3.6405
R1475 VDD.n197 VDD.n196 3.6405
R1476 VDD.n252 VDD.t403 3.6405
R1477 VDD.n252 VDD.n251 3.6405
R1478 VDD.n262 VDD.t523 3.6405
R1479 VDD.n262 VDD.n261 3.6405
R1480 VDD.n236 VDD.t619 3.6405
R1481 VDD.n236 VDD.n235 3.6405
R1482 VDD.n246 VDD.t387 3.6405
R1483 VDD.n246 VDD.n245 3.6405
R1484 VDD.n224 VDD.t401 3.6405
R1485 VDD.n224 VDD.n223 3.6405
R1486 VDD.n1781 VDD.t419 3.6405
R1487 VDD.n1781 VDD.n1780 3.6405
R1488 VDD.n11 VDD.t30 3.6405
R1489 VDD.n11 VDD.n10 3.6405
R1490 VDD.n9 VDD.t838 3.6405
R1491 VDD.n9 VDD.n8 3.6405
R1492 VDD.n1778 VDD.t26 3.6405
R1493 VDD.n1778 VDD.n1777 3.6405
R1494 VDD.n1776 VDD.t712 3.6405
R1495 VDD.n1776 VDD.n1775 3.6405
R1496 VDD.n1954 VDD.t28 3.6405
R1497 VDD.n1954 VDD.n1953 3.6405
R1498 VDD.n1946 VDD.t357 3.6405
R1499 VDD.n1946 VDD.n1945 3.6405
R1500 VDD.n1950 VDD.t356 3.6405
R1501 VDD.n1950 VDD.n1949 3.6405
R1502 VDD.n1948 VDD.t344 3.6405
R1503 VDD.n1948 VDD.n1947 3.6405
R1504 VDD.n2153 VDD.t554 3.6405
R1505 VDD.n2153 VDD.n2152 3.6405
R1506 VDD.n2151 VDD.t271 3.6405
R1507 VDD.n2151 VDD.n2150 3.6405
R1508 VDD.n2614 VDD.t114 3.6405
R1509 VDD.n2614 VDD.n2613 3.6405
R1510 VDD.n2616 VDD.t538 3.6405
R1511 VDD.n2616 VDD.n2615 3.6405
R1512 VDD.n1997 VDD.n1996 3.54622
R1513 VDD.n1951 VDD.n1950 3.54622
R1514 VDD.n649 VDD.t188 3.42047
R1515 VDD.n182 VDD.t383 3.33106
R1516 VDD.n991 VDD.n989 3.32815
R1517 VDD.n298 VDD.n295 3.30485
R1518 VDD.n304 VDD.n301 3.30485
R1519 VDD.n1217 VDD.n1216 3.30485
R1520 VDD.n1206 VDD.n1205 3.30485
R1521 VDD.n2202 VDD.t606 3.28543
R1522 VDD.n2418 VDD.t1010 3.28543
R1523 VDD.n1246 VDD.n489 3.28454
R1524 VDD.n2243 VDD.t655 3.27944
R1525 VDD.n2459 VDD.t879 3.27944
R1526 VDD.n2328 VDD.n2325 3.27159
R1527 VDD.n2333 VDD.n2318 3.27159
R1528 VDD.n2336 VDD.n2314 3.27159
R1529 VDD.n2338 VDD.n2311 3.27159
R1530 VDD.n2341 VDD.n2307 3.27159
R1531 VDD.n2345 VDD.n2304 3.27159
R1532 VDD.n2346 VDD.n2302 3.27159
R1533 VDD.n2293 VDD.n2193 3.27159
R1534 VDD.n2290 VDD.n2195 3.27159
R1535 VDD.n2287 VDD.n2197 3.27159
R1536 VDD.n2352 VDD.n2299 3.27159
R1537 VDD.n2571 VDD.n2568 3.27159
R1538 VDD.n2576 VDD.n2561 3.27159
R1539 VDD.n2579 VDD.n2557 3.27159
R1540 VDD.n2581 VDD.n2554 3.27159
R1541 VDD.n2584 VDD.n2550 3.27159
R1542 VDD.n2588 VDD.n2547 3.27159
R1543 VDD.n2509 VDD.n2409 3.27159
R1544 VDD.n2506 VDD.n2411 3.27159
R1545 VDD.n2503 VDD.n2413 3.27159
R1546 VDD.n2542 VDD.n2394 3.27159
R1547 VDD.n2515 VDD.n2405 3.27159
R1548 VDD.n2330 VDD.n2322 3.26834
R1549 VDD.n2573 VDD.n2565 3.26834
R1550 VDD.n2296 VDD.n2191 3.26449
R1551 VDD.n2512 VDD.n2407 3.26449
R1552 VDD.n2284 VDD.n2198 3.2505
R1553 VDD.n2500 VDD.n2414 3.2505
R1554 VDD.n1511 VDD.n1510 3.2486
R1555 VDD.n1302 VDD.n472 3.2486
R1556 VDD.n1668 VDD.t988 3.22394
R1557 VDD.n1662 VDD.t959 3.22394
R1558 VDD.n1655 VDD.t963 3.22394
R1559 VDD.n1687 VDD.t947 3.22394
R1560 VDD.n578 VDD.t935 3.22347
R1561 VDD.n574 VDD.t993 3.22347
R1562 VDD.n570 VDD.t981 3.22347
R1563 VDD.n566 VDD.t984 3.22347
R1564 VDD.n1199 VDD.t991 3.21802
R1565 VDD.n306 VDD.t953 3.21788
R1566 VDD.n291 VDD.t941 3.21785
R1567 VDD.n1195 VDD.t976 3.21781
R1568 VDD.n312 VDD.t961 3.21767
R1569 VDD.n1218 VDD.t950 3.21766
R1570 VDD.n1530 VDD.n1529 3.21752
R1571 VDD.n1209 VDD.t938 3.21671
R1572 VDD.n299 VDD.t996 3.21657
R1573 VDD.n2061 VDD.n2060 3.21512
R1574 VDD.n13 VDD.n12 3.20353
R1575 VDD.n1980 VDD.n1979 3.20342
R1576 VDD.n1294 VDD.t968 3.19864
R1577 VDD.n1259 VDD.t944 3.19113
R1578 VDD.n1461 VDD.t971 3.19113
R1579 VDD.n1501 VDD.t986 3.18927
R1580 VDD.n326 VDD.t974 3.1878
R1581 VDD.n475 VDD.t979 3.1878
R1582 VDD.n1028 VDD.n1027 3.16769
R1583 VDD.n1648 VDD.n1647 3.16769
R1584 VDD.n2063 VDD.n2062 3.16326
R1585 VDD.n2053 VDD.n2052 3.15744
R1586 VDD.n682 VDD.n681 3.15287
R1587 VDD VDD.n680 3.15287
R1588 VDD.n900 VDD.n898 3.15287
R1589 VDD.n902 VDD.n901 3.15287
R1590 VDD.n897 VDD.n896 3.15287
R1591 VDD VDD.n1969 3.15269
R1592 VDD.n1566 VDD.n278 3.15151
R1593 VDD.n1808 VDD.n1806 3.1505
R1594 VDD.n1815 VDD.n1808 3.1505
R1595 VDD.n1939 VDD.n1938 3.1505
R1596 VDD.n1938 VDD.n1937 3.1505
R1597 VDD.n1809 VDD.n1807 3.1505
R1598 VDD.n1936 VDD.n1809 3.1505
R1599 VDD.n1934 VDD 3.1505
R1600 VDD.n1935 VDD.n1934 3.1505
R1601 VDD.n1933 VDD.n1817 3.1505
R1602 VDD.n1817 VDD.n1816 3.1505
R1603 VDD.n1932 VDD.n1931 3.1505
R1604 VDD.n1931 VDD.n1930 3.1505
R1605 VDD.n1829 VDD.n1820 3.1505
R1606 VDD.n1929 VDD.n1820 3.1505
R1607 VDD.n1830 VDD.n1821 3.1505
R1608 VDD.n1814 VDD.n1813 3.1505
R1609 VDD.n1891 VDD.n1887 3.1505
R1610 VDD.n1896 VDD.n1895 3.1505
R1611 VDD.n1897 VDD.n1896 3.1505
R1612 VDD.n1893 VDD.n1885 3.1505
R1613 VDD.n1898 VDD.n1885 3.1505
R1614 VDD.n1900 VDD.n1886 3.1505
R1615 VDD.n1900 VDD.n1899 3.1505
R1616 VDD VDD.n1901 3.1505
R1617 VDD.n1901 VDD.n1884 3.1505
R1618 VDD.n1903 VDD.n1902 3.1505
R1619 VDD.n1904 VDD.n1903 3.1505
R1620 VDD.n1882 VDD.n1874 3.1505
R1621 VDD.n1905 VDD.n1882 3.1505
R1622 VDD.n1911 VDD.n1910 3.1505
R1623 VDD.n1910 VDD.n1909 3.1505
R1624 VDD.n1883 VDD.n1881 3.1505
R1625 VDD.n146 VDD.n145 3.1505
R1626 VDD.n144 VDD.n121 3.1505
R1627 VDD.n144 VDD.n143 3.1505
R1628 VDD.n125 VDD.n122 3.1505
R1629 VDD.n142 VDD.n122 3.1505
R1630 VDD.n140 VDD.n139 3.1505
R1631 VDD.n141 VDD.n140 3.1505
R1632 VDD VDD.n124 3.1505
R1633 VDD.n124 VDD.n123 3.1505
R1634 VDD.n137 VDD.n136 3.1505
R1635 VDD.n136 VDD.n135 3.1505
R1636 VDD.n127 VDD.n126 3.1505
R1637 VDD.n134 VDD.n127 3.1505
R1638 VDD.n132 VDD.n131 3.1505
R1639 VDD.n133 VDD.n132 3.1505
R1640 VDD.n130 VDD.n128 3.1505
R1641 VDD.n50 VDD.n47 3.1505
R1642 VDD.n62 VDD.n61 3.1505
R1643 VDD.n63 VDD.n62 3.1505
R1644 VDD.n46 VDD.n45 3.1505
R1645 VDD.n64 VDD.n46 3.1505
R1646 VDD.n68 VDD.n67 3.1505
R1647 VDD.n67 VDD.n66 3.1505
R1648 VDD VDD.n44 3.1505
R1649 VDD.n65 VDD.n44 3.1505
R1650 VDD.n71 VDD.n70 3.1505
R1651 VDD.n72 VDD.n71 3.1505
R1652 VDD.n42 VDD.n39 3.1505
R1653 VDD.n73 VDD.n42 3.1505
R1654 VDD.n76 VDD.n75 3.1505
R1655 VDD.n75 VDD.n74 3.1505
R1656 VDD.n43 VDD.n41 3.1505
R1657 VDD.n1500 VDD.n330 3.1505
R1658 VDD.n1505 VDD.n1504 3.1505
R1659 VDD.n1503 VDD.n328 3.1505
R1660 VDD.n1507 VDD.n328 3.1505
R1661 VDD.n1509 VDD.n329 3.1505
R1662 VDD.n1509 VDD.n1508 3.1505
R1663 VDD.n1511 VDD.n327 3.1505
R1664 VDD.n1514 VDD.n1513 3.1505
R1665 VDD.n1513 VDD.n1512 3.1505
R1666 VDD.n1516 VDD.n324 3.1505
R1667 VDD.n324 VDD.n323 3.1505
R1668 VDD.n1518 VDD.n1517 3.1505
R1669 VDD.n1519 VDD.n1518 3.1505
R1670 VDD.n325 VDD.n279 3.1505
R1671 VDD.n1565 VDD.n1564 3.1505
R1672 VDD.n282 VDD.n278 3.1505
R1673 VDD.n1568 VDD.n276 3.1505
R1674 VDD.n283 VDD.n276 3.1505
R1675 VDD.n1570 VDD.n1569 3.1505
R1676 VDD.n1571 VDD.n1570 3.1505
R1677 VDD.n269 VDD.n268 3.1505
R1678 VDD.n1572 VDD.n269 3.1505
R1679 VDD.n1582 VDD.n1581 3.1505
R1680 VDD.n1581 VDD.n1580 3.1505
R1681 VDD.n1583 VDD.n267 3.1505
R1682 VDD.n271 VDD.n267 3.1505
R1683 VDD.n1585 VDD.n1584 3.1505
R1684 VDD.n1586 VDD.n1585 3.1505
R1685 VDD.n240 VDD.n238 3.1505
R1686 VDD.n1587 VDD.n240 3.1505
R1687 VDD.n1608 VDD.n1607 3.1505
R1688 VDD.n1607 VDD.n1606 3.1505
R1689 VDD.n241 VDD.n239 3.1505
R1690 VDD.n1593 VDD.n241 3.1505
R1691 VDD.n1596 VDD.n1595 3.1505
R1692 VDD.n1597 VDD.n1596 3.1505
R1693 VDD.n174 VDD.n171 3.1505
R1694 VDD.n1598 VDD.n174 3.1505
R1695 VDD.n1561 VDD.n277 3.1505
R1696 VDD.n292 VDD.n281 3.1505
R1697 VDD.n1557 VDD.n1556 3.1505
R1698 VDD.n1554 VDD.n290 3.1505
R1699 VDD.n1553 VDD.n1552 3.1505
R1700 VDD.n1551 VDD.n1550 3.1505
R1701 VDD.n1548 VDD.n1547 3.1505
R1702 VDD.n1546 VDD.n1545 3.1505
R1703 VDD.n1544 VDD.n1543 3.1505
R1704 VDD.n1542 VDD.n1541 3.1505
R1705 VDD.n1540 VDD.n1539 3.1505
R1706 VDD.n1538 VDD.n1537 3.1505
R1707 VDD.n1535 VDD.n1534 3.1505
R1708 VDD.n1533 VDD.n1532 3.1505
R1709 VDD.n1531 VDD.n1530 3.1505
R1710 VDD.n1476 VDD.n1475 3.1505
R1711 VDD.n1478 VDD.n1477 3.1505
R1712 VDD.n1480 VDD.n1479 3.1505
R1713 VDD.n1482 VDD.n1481 3.1505
R1714 VDD.n1484 VDD.n1483 3.1505
R1715 VDD.n1486 VDD.n1485 3.1505
R1716 VDD.n1488 VDD.n1487 3.1505
R1717 VDD.n1490 VDD.n1489 3.1505
R1718 VDD.n1492 VDD.n1491 3.1505
R1719 VDD.n1494 VDD.n1493 3.1505
R1720 VDD.n332 VDD.n331 3.1505
R1721 VDD.n1499 VDD.n1498 3.1505
R1722 VDD VDD.n1402 3.1505
R1723 VDD.n1410 VDD.n1402 3.1505
R1724 VDD.n1422 VDD.n1421 3.1505
R1725 VDD.n1421 VDD.n1420 3.1505
R1726 VDD.n1409 VDD.n1408 3.1505
R1727 VDD.n1419 VDD.n1409 3.1505
R1728 VDD.n1417 VDD.n1416 3.1505
R1729 VDD.n1418 VDD.n1417 3.1505
R1730 VDD.n1415 VDD.n1411 3.1505
R1731 VDD.n1430 VDD.n1429 3.1505
R1732 VDD.n1399 VDD.n1398 3.1505
R1733 VDD.n1428 VDD.n1399 3.1505
R1734 VDD.n1426 VDD.n1425 3.1505
R1735 VDD.n1427 VDD.n1426 3.1505
R1736 VDD.n1424 VDD.n1401 3.1505
R1737 VDD.n1401 VDD.n1400 3.1505
R1738 VDD.n1390 VDD.n1389 3.1505
R1739 VDD.n1437 VDD.n1390 3.1505
R1740 VDD.n1435 VDD.n1434 3.1505
R1741 VDD.n1436 VDD.n1435 3.1505
R1742 VDD.n1433 VDD.n1391 3.1505
R1743 VDD.n431 VDD.n420 3.1505
R1744 VDD.n423 VDD.n420 3.1505
R1745 VDD.n430 VDD.n429 3.1505
R1746 VDD.n429 VDD.n428 3.1505
R1747 VDD.n422 VDD.n421 3.1505
R1748 VDD.n427 VDD.n422 3.1505
R1749 VDD.n426 VDD.n425 3.1505
R1750 VDD.n439 VDD.n409 3.1505
R1751 VDD.n438 VDD.n411 3.1505
R1752 VDD.n438 VDD.n437 3.1505
R1753 VDD.n414 VDD.n410 3.1505
R1754 VDD.n436 VDD.n410 3.1505
R1755 VDD.n434 VDD.n433 3.1505
R1756 VDD.n435 VDD.n434 3.1505
R1757 VDD VDD.n413 3.1505
R1758 VDD.n413 VDD.n412 3.1505
R1759 VDD.n445 VDD.n444 3.1505
R1760 VDD.n451 VDD.n450 3.1505
R1761 VDD.n452 VDD.n451 3.1505
R1762 VDD.n449 VDD.n404 3.1505
R1763 VDD.n404 VDD.n403 3.1505
R1764 VDD.n448 VDD.n447 3.1505
R1765 VDD.n447 VDD.n446 3.1505
R1766 VDD.n393 VDD.n392 3.1505
R1767 VDD.n459 VDD.n458 3.1505
R1768 VDD.n460 VDD.n459 3.1505
R1769 VDD.n457 VDD.n395 3.1505
R1770 VDD.n395 VDD.n394 3.1505
R1771 VDD.n456 VDD.n455 3.1505
R1772 VDD.n455 VDD.n454 3.1505
R1773 VDD VDD.n402 3.1505
R1774 VDD.n453 VDD.n402 3.1505
R1775 VDD.n1309 VDD.n1308 3.1505
R1776 VDD.n1292 VDD.n474 3.1505
R1777 VDD.n474 VDD.n473 3.1505
R1778 VDD.n1299 VDD.n1298 3.1505
R1779 VDD.n1300 VDD.n1299 3.1505
R1780 VDD.n1297 VDD.n472 3.1505
R1781 VDD.n1296 VDD.n470 3.1505
R1782 VDD.n1303 VDD.n470 3.1505
R1783 VDD.n1305 VDD.n469 3.1505
R1784 VDD.n1305 VDD.n1304 3.1505
R1785 VDD.n1307 VDD.n1306 3.1505
R1786 VDD.n1291 VDD.n1290 3.1505
R1787 VDD.n1290 VDD.n1289 3.1505
R1788 VDD.n482 VDD.n481 3.1505
R1789 VDD.n477 VDD.n476 3.1505
R1790 VDD.n1036 VDD.n1035 3.1505
R1791 VDD.n1035 VDD.n1034 3.1505
R1792 VDD.n1037 VDD.n557 3.1505
R1793 VDD.n557 VDD.n554 3.1505
R1794 VDD.n1039 VDD.n1038 3.1505
R1795 VDD.n1040 VDD.n1039 3.1505
R1796 VDD.n550 VDD.n549 3.1505
R1797 VDD.n555 VDD.n550 3.1505
R1798 VDD.n1051 VDD.n1050 3.1505
R1799 VDD.n1050 VDD.n1049 3.1505
R1800 VDD.n1052 VDD.n543 3.1505
R1801 VDD.n543 VDD.n542 3.1505
R1802 VDD.n1056 VDD.n1055 3.1505
R1803 VDD.n1057 VDD.n1056 3.1505
R1804 VDD.n1054 VDD.n548 3.1505
R1805 VDD.n548 VDD.n547 3.1505
R1806 VDD.n535 VDD.n534 3.1505
R1807 VDD.n545 VDD.n534 3.1505
R1808 VDD.n1121 VDD.n1120 3.1505
R1809 VDD.n1122 VDD.n1121 3.1505
R1810 VDD.n525 VDD.n524 3.1505
R1811 VDD.n532 VDD.n525 3.1505
R1812 VDD.n1134 VDD.n1133 3.1505
R1813 VDD.n1133 VDD.n1132 3.1505
R1814 VDD.n1135 VDD.n523 3.1505
R1815 VDD.n523 VDD.n521 3.1505
R1816 VDD.n1137 VDD.n1136 3.1505
R1817 VDD.n1138 VDD.n1137 3.1505
R1818 VDD.n516 VDD.n515 3.1505
R1819 VDD.n517 VDD.n516 3.1505
R1820 VDD.n1150 VDD.n1149 3.1505
R1821 VDD.n1149 VDD.n1148 3.1505
R1822 VDD.n1151 VDD.n513 3.1505
R1823 VDD.n513 VDD.n511 3.1505
R1824 VDD.n1154 VDD.n1153 3.1505
R1825 VDD.n1155 VDD.n1154 3.1505
R1826 VDD.n506 VDD.n505 3.1505
R1827 VDD.n507 VDD.n506 3.1505
R1828 VDD.n1167 VDD.n1166 3.1505
R1829 VDD.n1166 VDD.n1165 3.1505
R1830 VDD.n1168 VDD.n503 3.1505
R1831 VDD.n503 VDD.n501 3.1505
R1832 VDD.n559 VDD.n558 3.1505
R1833 VDD.n562 VDD.n559 3.1505
R1834 VDD.n696 VDD.n664 3.1505
R1835 VDD.n639 VDD.n633 3.1505
R1836 VDD.n641 VDD.n639 3.1505
R1837 VDD.n715 VDD.n714 3.1505
R1838 VDD.n716 VDD.n715 3.1505
R1839 VDD.n712 VDD.n659 3.1505
R1840 VDD.n662 VDD.n659 3.1505
R1841 VDD.n707 VDD.n706 3.1505
R1842 VDD.n708 VDD.n707 3.1505
R1843 VDD.n718 VDD.n657 3.1505
R1844 VDD.n718 VDD.n717 3.1505
R1845 VDD.n713 VDD.n656 3.1505
R1846 VDD.n658 VDD.n656 3.1505
R1847 VDD.n711 VDD.n710 3.1505
R1848 VDD.n710 VDD.n709 3.1505
R1849 VDD VDD.n722 3.1505
R1850 VDD.n722 VDD.n721 3.1505
R1851 VDD.n719 VDD 3.1505
R1852 VDD.n720 VDD.n719 3.1505
R1853 VDD.n596 VDD.n591 3.1505
R1854 VDD.n618 VDD.n591 3.1505
R1855 VDD.n736 VDD.n735 3.1505
R1856 VDD.n735 VDD.n734 3.1505
R1857 VDD.n643 VDD.n592 3.1505
R1858 VDD.n647 VDD.n592 3.1505
R1859 VDD.n612 VDD.n611 3.1505
R1860 VDD.n611 VDD.n601 3.1505
R1861 VDD.n622 VDD.n594 3.1505
R1862 VDD.n623 VDD.n622 3.1505
R1863 VDD.n652 VDD.n642 3.1505
R1864 VDD.n648 VDD.n642 3.1505
R1865 VDD.n617 VDD.n595 3.1505
R1866 VDD.n609 VDD.n602 3.1505
R1867 VDD.n613 VDD.n595 3.1505
R1868 VDD.n621 VDD.n589 3.1505
R1869 VDD.n621 VDD.n593 3.1505
R1870 VDD.n854 VDD.n850 3.1505
R1871 VDD.n849 VDD.n848 3.1505
R1872 VDD.n857 VDD.n849 3.1505
R1873 VDD.n860 VDD.n859 3.1505
R1874 VDD.n859 VDD.n858 3.1505
R1875 VDD.n861 VDD.n842 3.1505
R1876 VDD.n842 VDD.n841 3.1505
R1877 VDD.n863 VDD 3.1505
R1878 VDD.n864 VDD.n863 3.1505
R1879 VDD.n840 VDD.n839 3.1505
R1880 VDD.n865 VDD.n840 3.1505
R1881 VDD.n869 VDD.n868 3.1505
R1882 VDD.n868 VDD.n867 3.1505
R1883 VDD.n870 VDD.n838 3.1505
R1884 VDD.n866 VDD.n838 3.1505
R1885 VDD.n837 VDD.n836 3.1505
R1886 VDD.n790 VDD.n788 3.1505
R1887 VDD.n790 VDD.n789 3.1505
R1888 VDD.n792 VDD.n791 3.1505
R1889 VDD.n791 VDD.n779 3.1505
R1890 VDD.n778 VDD.n777 3.1505
R1891 VDD.n795 VDD.n778 3.1505
R1892 VDD.n798 VDD.n797 3.1505
R1893 VDD.n797 VDD.n796 3.1505
R1894 VDD.n788 VDD.n780 3.1505
R1895 VDD.n789 VDD.n780 3.1505
R1896 VDD.n793 VDD.n792 3.1505
R1897 VDD.n793 VDD.n779 3.1505
R1898 VDD.n794 VDD.n777 3.1505
R1899 VDD.n795 VDD.n794 3.1505
R1900 VDD.n798 VDD.n776 3.1505
R1901 VDD.n796 VDD.n776 3.1505
R1902 VDD VDD.n773 3.1505
R1903 VDD.n775 VDD.n773 3.1505
R1904 VDD.n813 VDD.n774 3.1505
R1905 VDD.n813 VDD.n812 3.1505
R1906 VDD.n814 VDD.n771 3.1505
R1907 VDD.n815 VDD.n814 3.1505
R1908 VDD.n818 VDD.n770 3.1505
R1909 VDD.n816 VDD.n770 3.1505
R1910 VDD.n820 VDD.n819 3.1505
R1911 VDD.n821 VDD.n820 3.1505
R1912 VDD.n824 VDD.n768 3.1505
R1913 VDD.n822 VDD.n768 3.1505
R1914 VDD.n810 VDD 3.1505
R1915 VDD.n810 VDD.n775 3.1505
R1916 VDD.n811 VDD.n774 3.1505
R1917 VDD.n812 VDD.n811 3.1505
R1918 VDD.n772 VDD.n771 3.1505
R1919 VDD.n815 VDD.n772 3.1505
R1920 VDD.n818 VDD.n817 3.1505
R1921 VDD.n817 VDD.n816 3.1505
R1922 VDD.n819 VDD.n769 3.1505
R1923 VDD.n821 VDD.n769 3.1505
R1924 VDD.n960 VDD.n959 3.1505
R1925 VDD.n959 VDD.n950 3.1505
R1926 VDD.n958 VDD.n949 3.1505
R1927 VDD.n958 VDD.n957 3.1505
R1928 VDD.n952 VDD.n951 3.1505
R1929 VDD.n956 VDD.n951 3.1505
R1930 VDD.n955 VDD.n954 3.1505
R1931 VDD.n930 VDD.n929 3.1505
R1932 VDD.n963 VDD.n962 3.1505
R1933 VDD.n964 VDD.n963 3.1505
R1934 VDD VDD.n943 3.1505
R1935 VDD.n943 VDD.n942 3.1505
R1936 VDD.n1026 VDD.n561 3.1505
R1937 VDD.n1024 VDD.n1023 3.1505
R1938 VDD.n1022 VDD.n565 3.1505
R1939 VDD.n1020 VDD.n1019 3.1505
R1940 VDD.n1018 VDD.n567 3.1505
R1941 VDD.n1016 VDD.n1015 3.1505
R1942 VDD.n1014 VDD.n569 3.1505
R1943 VDD.n1012 VDD.n1011 3.1505
R1944 VDD.n1010 VDD.n571 3.1505
R1945 VDD.n1008 VDD.n1007 3.1505
R1946 VDD.n1005 VDD.n573 3.1505
R1947 VDD.n1004 VDD.n1003 3.1505
R1948 VDD.n1002 VDD.n575 3.1505
R1949 VDD.n1000 VDD.n999 3.1505
R1950 VDD.n997 VDD.n577 3.1505
R1951 VDD.n996 VDD.n995 3.1505
R1952 VDD.n1029 VDD.n560 3.1505
R1953 VDD.n563 VDD.n560 3.1505
R1954 VDD.n1031 VDD.n1030 3.1505
R1955 VDD.n1032 VDD.n1031 3.1505
R1956 VDD.n553 VDD.n552 3.1505
R1957 VDD.n1033 VDD.n553 3.1505
R1958 VDD.n1043 VDD.n1042 3.1505
R1959 VDD.n1042 VDD.n1041 3.1505
R1960 VDD.n1044 VDD.n551 3.1505
R1961 VDD.n556 VDD.n551 3.1505
R1962 VDD.n1046 VDD.n1045 3.1505
R1963 VDD.n1047 VDD.n1046 3.1505
R1964 VDD.n540 VDD.n538 3.1505
R1965 VDD.n1048 VDD.n540 3.1505
R1966 VDD.n1060 VDD.n1059 3.1505
R1967 VDD.n1059 VDD.n1058 3.1505
R1968 VDD.n541 VDD.n539 3.1505
R1969 VDD.n544 VDD.n541 3.1505
R1970 VDD.n531 VDD.n530 3.1505
R1971 VDD.n546 VDD.n531 3.1505
R1972 VDD.n1125 VDD.n1124 3.1505
R1973 VDD.n1124 VDD.n1123 3.1505
R1974 VDD.n1127 VDD.n526 3.1505
R1975 VDD.n533 VDD.n526 3.1505
R1976 VDD.n1129 VDD.n1128 3.1505
R1977 VDD.n1130 VDD.n1129 3.1505
R1978 VDD.n520 VDD.n519 3.1505
R1979 VDD.n1131 VDD.n520 3.1505
R1980 VDD.n1141 VDD.n1140 3.1505
R1981 VDD.n1140 VDD.n1139 3.1505
R1982 VDD.n1142 VDD.n518 3.1505
R1983 VDD.n522 VDD.n518 3.1505
R1984 VDD.n1145 VDD.n1144 3.1505
R1985 VDD.n1146 VDD.n1145 3.1505
R1986 VDD.n1143 VDD.n510 3.1505
R1987 VDD.n1147 VDD.n510 3.1505
R1988 VDD.n1158 VDD.n1157 3.1505
R1989 VDD.n1157 VDD.n1156 3.1505
R1990 VDD.n1159 VDD.n508 3.1505
R1991 VDD.n512 VDD.n508 3.1505
R1992 VDD.n1162 VDD.n1161 3.1505
R1993 VDD.n1163 VDD.n1162 3.1505
R1994 VDD.n1160 VDD.n500 3.1505
R1995 VDD.n1164 VDD.n500 3.1505
R1996 VDD.n1175 VDD.n1174 3.1505
R1997 VDD.n1174 VDD.n1173 3.1505
R1998 VDD.n1176 VDD.n498 3.1505
R1999 VDD.n502 VDD.n498 3.1505
R2000 VDD.n1178 VDD.n1177 3.1505
R2001 VDD.n1179 VDD.n1178 3.1505
R2002 VDD.n491 VDD.n490 3.1505
R2003 VDD.n1180 VDD.n491 3.1505
R2004 VDD.n1191 VDD.n1190 3.1505
R2005 VDD.n1190 VDD.n1189 3.1505
R2006 VDD.n1192 VDD.n488 3.1505
R2007 VDD.n493 VDD.n488 3.1505
R2008 VDD.n1278 VDD.n1277 3.1505
R2009 VDD.n1279 VDD.n1278 3.1505
R2010 VDD.n1171 VDD.n1170 3.1505
R2011 VDD.n1172 VDD.n1171 3.1505
R2012 VDD.n496 VDD.n495 3.1505
R2013 VDD.n497 VDD.n496 3.1505
R2014 VDD.n1183 VDD.n1182 3.1505
R2015 VDD.n1182 VDD.n1181 3.1505
R2016 VDD.n1184 VDD.n494 3.1505
R2017 VDD.n494 VDD.n492 3.1505
R2018 VDD.n1187 VDD.n1186 3.1505
R2019 VDD.n1188 VDD.n1187 3.1505
R2020 VDD.n1185 VDD.n486 3.1505
R2021 VDD.n487 VDD.n486 3.1505
R2022 VDD.n1281 VDD.n483 3.1505
R2023 VDD.n1281 VDD.n1280 3.1505
R2024 VDD.n1287 VDD.n1286 3.1505
R2025 VDD.n1288 VDD.n1287 3.1505
R2026 VDD.n1244 VDD.n1193 3.1505
R2027 VDD.n1243 VDD.n1242 3.1505
R2028 VDD.n1240 VDD.n1239 3.1505
R2029 VDD.n1238 VDD.n1237 3.1505
R2030 VDD.n1236 VDD.n1235 3.1505
R2031 VDD.n1234 VDD.n1233 3.1505
R2032 VDD.n1232 VDD.n1231 3.1505
R2033 VDD.n1230 VDD.n1229 3.1505
R2034 VDD.n1227 VDD.n1226 3.1505
R2035 VDD.n1225 VDD.n1210 3.1505
R2036 VDD.n1223 VDD.n1222 3.1505
R2037 VDD.n1220 VDD.n1212 3.1505
R2038 VDD.n485 VDD.n484 3.1505
R2039 VDD.n1284 VDD.n1283 3.1505
R2040 VDD.n1283 VDD.n479 3.1505
R2041 VDD.n1247 VDD.n1246 3.1505
R2042 VDD.n1275 VDD.n1274 3.1505
R2043 VDD.n1272 VDD.n1271 3.1505
R2044 VDD.n1269 VDD.n1250 3.1505
R2045 VDD.n1250 VDD.n1249 3.1505
R2046 VDD.n1268 VDD.n1267 3.1505
R2047 VDD.n1267 VDD.n1266 3.1505
R2048 VDD.n1255 VDD.n1254 3.1505
R2049 VDD.n1265 VDD.n1255 3.1505
R2050 VDD.n1263 VDD.n1262 3.1505
R2051 VDD.n1264 VDD.n1263 3.1505
R2052 VDD.n1261 VDD.n1258 3.1505
R2053 VDD.n378 VDD.n376 3.1505
R2054 VDD.n1311 VDD.n1310 3.1505
R2055 VDD.n1313 VDD.n1312 3.1505
R2056 VDD.n1315 VDD.n1314 3.1505
R2057 VDD.n1317 VDD.n1316 3.1505
R2058 VDD.n1319 VDD.n1318 3.1505
R2059 VDD.n1321 VDD.n1320 3.1505
R2060 VDD.n1323 VDD.n1322 3.1505
R2061 VDD.n1325 VDD.n1324 3.1505
R2062 VDD.n1327 VDD.n1326 3.1505
R2063 VDD.n1329 VDD.n1328 3.1505
R2064 VDD.n1331 VDD.n1330 3.1505
R2065 VDD.n1333 VDD.n1332 3.1505
R2066 VDD.n1335 VDD.n1334 3.1505
R2067 VDD.n379 VDD.n377 3.1505
R2068 VDD.n1340 VDD.n1339 3.1505
R2069 VDD VDD.n1357 3.1505
R2070 VDD.n1357 VDD.n1356 3.1505
R2071 VDD.n1349 VDD.n1348 3.1505
R2072 VDD.n1350 VDD.n375 3.1505
R2073 VDD.n375 VDD.n374 3.1505
R2074 VDD.n1353 VDD.n1352 3.1505
R2075 VDD.n1354 VDD.n1353 3.1505
R2076 VDD.n1351 VDD.n373 3.1505
R2077 VDD.n1355 VDD.n373 3.1505
R2078 VDD.n1358 VDD.n366 3.1505
R2079 VDD.n366 VDD.n365 3.1505
R2080 VDD.n1360 VDD.n1359 3.1505
R2081 VDD.n1361 VDD.n1360 3.1505
R2082 VDD.n364 VDD.n363 3.1505
R2083 VDD.n1362 VDD.n364 3.1505
R2084 VDD.n1364 VDD.n1363 3.1505
R2085 VDD.n1378 VDD.n1377 3.1505
R2086 VDD.n1382 VDD.n349 3.1505
R2087 VDD.n1383 VDD.n1382 3.1505
R2088 VDD.n1381 VDD.n1380 3.1505
R2089 VDD.n1381 VDD.n1373 3.1505
R2090 VDD.n1379 VDD.n1374 3.1505
R2091 VDD.n1376 VDD.n1374 3.1505
R2092 VDD.n357 VDD 3.1505
R2093 VDD.n1384 VDD.n357 3.1505
R2094 VDD.n1369 VDD.n358 3.1505
R2095 VDD.n1370 VDD.n355 3.1505
R2096 VDD.n1371 VDD.n1370 3.1505
R2097 VDD.n1372 VDD.n356 3.1505
R2098 VDD.n1386 VDD.n1385 3.1505
R2099 VDD.n1440 VDD.n1439 3.1505
R2100 VDD.n1439 VDD.n1438 3.1505
R2101 VDD VDD.n348 3.1505
R2102 VDD.n348 VDD.n347 3.1505
R2103 VDD.n1443 VDD.n1442 3.1505
R2104 VDD.n1444 VDD.n1443 3.1505
R2105 VDD.n346 VDD.n345 3.1505
R2106 VDD.n1445 VDD.n346 3.1505
R2107 VDD.n1447 VDD.n1446 3.1505
R2108 VDD.n1474 VDD.n334 3.1505
R2109 VDD.n1496 VDD.n334 3.1505
R2110 VDD.n1473 VDD.n1472 3.1505
R2111 VDD.n1471 VDD.n1470 3.1505
R2112 VDD.n1460 VDD.n1457 3.1505
R2113 VDD.n1466 VDD.n1465 3.1505
R2114 VDD.n1467 VDD.n1466 3.1505
R2115 VDD.n1463 VDD.n1459 3.1505
R2116 VDD.n1459 VDD.n1458 3.1505
R2117 VDD.n1462 VDD.n319 3.1505
R2118 VDD.n321 VDD.n319 3.1505
R2119 VDD.n1523 VDD.n320 3.1505
R2120 VDD.n1523 VDD.n1522 3.1505
R2121 VDD.n1525 VDD.n1524 3.1505
R2122 VDD.n1528 VDD.n1527 3.1505
R2123 VDD.n1469 VDD.n1456 3.1505
R2124 VDD.n274 VDD.n273 3.1505
R2125 VDD.n275 VDD.n274 3.1505
R2126 VDD.n1575 VDD.n1574 3.1505
R2127 VDD.n1574 VDD.n1573 3.1505
R2128 VDD.n1576 VDD.n272 3.1505
R2129 VDD.n272 VDD.n270 3.1505
R2130 VDD.n1578 VDD.n1577 3.1505
R2131 VDD.n1579 VDD.n1578 3.1505
R2132 VDD.n265 VDD.n264 3.1505
R2133 VDD.n266 VDD.n265 3.1505
R2134 VDD.n1589 VDD.n1588 3.1505
R2135 VDD.n1588 VDD.t386 3.1505
R2136 VDD.n1590 VDD.n243 3.1505
R2137 VDD.n243 VDD.n242 3.1505
R2138 VDD.n1604 VDD.n1603 3.1505
R2139 VDD.n1605 VDD.n1604 3.1505
R2140 VDD.n1602 VDD.n244 3.1505
R2141 VDD.n1594 VDD.n244 3.1505
R2142 VDD.n1601 VDD.n1600 3.1505
R2143 VDD.n1600 VDD.n1599 3.1505
R2144 VDD.n1592 VDD.n177 3.1505
R2145 VDD.n177 VDD.n176 3.1505
R2146 VDD.n1760 VDD.n1759 3.1505
R2147 VDD.n1761 VDD.n1760 3.1505
R2148 VDD.n1758 VDD.n178 3.1505
R2149 VDD.n183 VDD.n178 3.1505
R2150 VDD.n1757 VDD.n1756 3.1505
R2151 VDD.n1756 VDD.n1755 3.1505
R2152 VDD.n181 VDD.n180 3.1505
R2153 VDD.n185 VDD.n181 3.1505
R2154 VDD.n195 VDD.n193 3.1505
R2155 VDD.n193 VDD.n192 3.1505
R2156 VDD.n1746 VDD.n1745 3.1505
R2157 VDD.n1747 VDD.n1746 3.1505
R2158 VDD.n1744 VDD.n194 3.1505
R2159 VDD.n202 VDD.n194 3.1505
R2160 VDD.n1742 VDD.n1741 3.1505
R2161 VDD.n1741 VDD.n1740 3.1505
R2162 VDD.n200 VDD.n199 3.1505
R2163 VDD.n204 VDD.n200 3.1505
R2164 VDD.n215 VDD.n213 3.1505
R2165 VDD.n213 VDD.n212 3.1505
R2166 VDD.n1731 VDD.n1730 3.1505
R2167 VDD.n1732 VDD.n1731 3.1505
R2168 VDD.n1728 VDD.n214 3.1505
R2169 VDD.n1632 VDD.n214 3.1505
R2170 VDD.n1727 VDD.n1726 3.1505
R2171 VDD.n1726 VDD.n1725 3.1505
R2172 VDD.n1631 VDD.n1630 3.1505
R2173 VDD.n1634 VDD.n1631 3.1505
R2174 VDD.n1646 VDD.n1644 3.1505
R2175 VDD.n1644 VDD.n1642 3.1505
R2176 VDD.n1716 VDD.n1715 3.1505
R2177 VDD.n1717 VDD.n1716 3.1505
R2178 VDD.n1714 VDD.n1645 3.1505
R2179 VDD.n1699 VDD.n1645 3.1505
R2180 VDD.n1713 VDD.n1712 3.1505
R2181 VDD.n1670 VDD.n1664 3.1505
R2182 VDD.n1674 VDD.n1664 3.1505
R2183 VDD.n1676 VDD.n1665 3.1505
R2184 VDD.n1676 VDD.n1675 3.1505
R2185 VDD.n1677 VDD.n1663 3.1505
R2186 VDD.n1677 VDD.n1658 3.1505
R2187 VDD.n1679 VDD.n1678 3.1505
R2188 VDD.n1678 VDD.n1659 3.1505
R2189 VDD.n1680 VDD.n1661 3.1505
R2190 VDD.n1661 VDD.n1660 3.1505
R2191 VDD.n1683 VDD.n1682 3.1505
R2192 VDD.n1684 VDD.n1683 3.1505
R2193 VDD.n1654 VDD.n1652 3.1505
R2194 VDD.n1652 VDD.n1650 3.1505
R2195 VDD.n1706 VDD.n1705 3.1505
R2196 VDD.n1707 VDD.n1706 3.1505
R2197 VDD.n1703 VDD.n1653 3.1505
R2198 VDD.n1653 VDD.n1651 3.1505
R2199 VDD.n1702 VDD.n1701 3.1505
R2200 VDD.n1701 VDD.n1700 3.1505
R2201 VDD.n1657 VDD.n1656 3.1505
R2202 VDD.n1698 VDD.n1657 3.1505
R2203 VDD.n1696 VDD.n1695 3.1505
R2204 VDD.n1697 VDD.n1696 3.1505
R2205 VDD.n1693 VDD.n1686 3.1505
R2206 VDD.n1686 VDD.n1685 3.1505
R2207 VDD.n1692 VDD.n1691 3.1505
R2208 VDD.n1691 VDD.n1690 3.1505
R2209 VDD.n1689 VDD.n1688 3.1505
R2210 VDD.n1689 VDD.n1649 3.1505
R2211 VDD.n1672 VDD.n1671 3.1505
R2212 VDD.n1667 VDD.n1666 3.1505
R2213 VDD.n1640 VDD.n1639 3.1505
R2214 VDD.n1643 VDD.n1640 3.1505
R2215 VDD.n175 VDD.n172 3.1505
R2216 VDD.n182 VDD.n175 3.1505
R2217 VDD.n188 VDD.n186 3.1505
R2218 VDD.n186 VDD.n184 3.1505
R2219 VDD.n1753 VDD.n1752 3.1505
R2220 VDD.n1754 VDD.n1753 3.1505
R2221 VDD.n1751 VDD.n187 3.1505
R2222 VDD.n191 VDD.n187 3.1505
R2223 VDD.n1750 VDD.n1749 3.1505
R2224 VDD.n1749 VDD.n1748 3.1505
R2225 VDD.n190 VDD.n189 3.1505
R2226 VDD.n201 VDD.n190 3.1505
R2227 VDD.n207 VDD.n205 3.1505
R2228 VDD.n205 VDD.n203 3.1505
R2229 VDD.n1738 VDD.n1737 3.1505
R2230 VDD.n1739 VDD.n1738 3.1505
R2231 VDD.n1736 VDD.n206 3.1505
R2232 VDD.n211 VDD.n206 3.1505
R2233 VDD.n1735 VDD.n1734 3.1505
R2234 VDD.n1734 VDD.n1733 3.1505
R2235 VDD.n1637 VDD.n209 3.1505
R2236 VDD.n210 VDD.n209 3.1505
R2237 VDD.n1638 VDD.n1635 3.1505
R2238 VDD.n1635 VDD.n1633 3.1505
R2239 VDD.n1723 VDD.n1722 3.1505
R2240 VDD.n1724 VDD.n1723 3.1505
R2241 VDD.n1721 VDD.n1636 3.1505
R2242 VDD.n1641 VDD.n1636 3.1505
R2243 VDD.n1720 VDD.n1719 3.1505
R2244 VDD.n1719 VDD.n1718 3.1505
R2245 VDD.n1764 VDD.n1763 3.1505
R2246 VDD.n1763 VDD.n1762 3.1505
R2247 VDD.n2124 VDD.n2123 3.1505
R2248 VDD.n2127 VDD.n2126 3.1505
R2249 VDD.n2126 VDD.n2125 3.1505
R2250 VDD.n2130 VDD.n2129 3.1505
R2251 VDD.n2129 VDD.n2128 3.1505
R2252 VDD.n2140 VDD.n2139 3.1505
R2253 VDD.n2139 VDD.n2138 3.1505
R2254 VDD.n2143 VDD 3.1505
R2255 VDD.n2143 VDD.n2142 3.1505
R2256 VDD.n2146 VDD.n2145 3.1505
R2257 VDD.n2145 VDD.n2144 3.1505
R2258 VDD.n2149 VDD.n2148 3.1505
R2259 VDD.n2148 VDD.n2147 3.1505
R2260 VDD.n2158 VDD.n2157 3.1505
R2261 VDD.n2157 VDD.n2156 3.1505
R2262 VDD.n2081 VDD.n2080 3.1505
R2263 VDD.n2648 VDD.n2647 3.1505
R2264 VDD.n2647 VDD.n2646 3.1505
R2265 VDD.n2627 VDD.n2626 3.1505
R2266 VDD.n2626 VDD.n2625 3.1505
R2267 VDD.n2630 VDD.n2629 3.1505
R2268 VDD.n2629 VDD.n2628 3.1505
R2269 VDD VDD.n2638 3.1505
R2270 VDD.n2638 VDD.n2637 3.1505
R2271 VDD.n2636 VDD.n2634 3.1505
R2272 VDD.n2636 VDD.n2635 3.1505
R2273 VDD.n2633 VDD.n2632 3.1505
R2274 VDD.n2632 VDD.n2631 3.1505
R2275 VDD.n2621 VDD.n2620 3.1505
R2276 VDD.n2620 VDD.n2619 3.1505
R2277 VDD.n2608 VDD.n2607 3.1505
R2278 VDD.n2645 VDD.n2644 3.1505
R2279 VDD.n2682 VDD.n2681 3.1505
R2280 VDD.n2681 VDD.t31 3.1505
R2281 VDD.n2174 VDD.n2173 3.1505
R2282 VDD.n2680 VDD.n2679 3.1505
R2283 VDD.t31 VDD.n2680 3.1505
R2284 VDD.n1 VDD.n0 3.1505
R2285 VDD.n929 VDD.n928 3.14819
R2286 VDD.n2004 VDD.n1988 3.13854
R2287 VDD.n2006 VDD.n1985 3.13854
R2288 VDD.n2007 VDD.n1983 3.13854
R2289 VDD.n16 VDD.n9 3.13659
R2290 VDD.n1779 VDD.n1778 3.13659
R2291 VDD.n1787 VDD.n1776 3.13659
R2292 VDD.n1338 VDD.n379 3.09085
R2293 VDD.n1826 VDD.n1825 3.06224
R2294 VDD.n1879 VDD.n1876 3.06224
R2295 VDD.n119 VDD.n116 3.06224
R2296 VDD.n58 VDD.n55 3.06224
R2297 VDD.n1453 VDD.n1450 3.06224
R2298 VDD.n1407 VDD.n1406 3.06224
R2299 VDD.n419 VDD.n416 3.06224
R2300 VDD.n400 VDD.n397 3.06224
R2301 VDD.n638 VDD.n637 3.06224
R2302 VDD.n632 VDD.n629 3.06224
R2303 VDD.n847 VDD.n844 3.06224
R2304 VDD.n803 VDD.n800 3.06224
R2305 VDD.n808 VDD.n807 3.06224
R2306 VDD.n948 VDD.n945 3.06224
R2307 VDD.n371 VDD.n370 3.06224
R2308 VDD.n354 VDD.n353 3.06224
R2309 VDD.n2154 VDD.n2151 3.06224
R2310 VDD.n2617 VDD.n2616 3.06224
R2311 VDD.n2592 VDD.n2384 3.04367
R2312 VDD.n1497 VDD.n332 3.04049
R2313 VDD.n1477 VDD.n335 3.03982
R2314 VDD.n1312 VDD.n380 3.03982
R2315 VDD.n1047 VDD.t174 2.91474
R2316 VDD.n1148 VDD.t93 2.91474
R2317 VDD.n1783 VDD.n1781 2.88811
R2318 VDD.n1837 VDD.n1835 2.87637
R2319 VDD.n1795 VDD.n1794 2.87637
R2320 VDD.n1867 VDD.n1865 2.87637
R2321 VDD.n1850 VDD.n1849 2.87637
R2322 VDD.n160 VDD.n158 2.87637
R2323 VDD.n24 VDD.n23 2.87637
R2324 VDD.n100 VDD.n98 2.87637
R2325 VDD.n81 VDD.n80 2.87637
R2326 VDD.n687 VDD.n685 2.87637
R2327 VDD.n676 VDD.n674 2.87637
R2328 VDD.n892 VDD.n891 2.87637
R2329 VDD.n887 VDD.n886 2.87637
R2330 VDD.n2089 VDD.n2087 2.87637
R2331 VDD.n2108 VDD.n2107 2.87637
R2332 VDD.n2599 VDD.n2597 2.87637
R2333 VDD.n2652 VDD.n2651 2.87637
R2334 VDD.n2014 VDD.n2011 2.87577
R2335 VDD.n149 VDD.n110 2.83323
R2336 VDD.n2043 VDD.n2042 2.82741
R2337 VDD.n1998 VDD.n1992 2.78441
R2338 VDD.n1997 VDD.n1994 2.78441
R2339 VDD.n1952 VDD.n1946 2.78441
R2340 VDD.n1951 VDD.n1948 2.78441
R2341 VDD.n1560 VDD.n281 2.7478
R2342 VDD.n1558 VDD.n281 2.7478
R2343 VDD.n2679 VDD.n2678 2.60854
R2344 VDD.n1999 VDD.n1990 2.6005
R2345 VDD.n1826 VDD.n1823 2.6005
R2346 VDD.n1879 VDD.n1878 2.6005
R2347 VDD.n119 VDD.n118 2.6005
R2348 VDD.n58 VDD.n57 2.6005
R2349 VDD.n231 VDD.n230 2.6005
R2350 VDD.n298 VDD.n297 2.6005
R2351 VDD.n304 VDD.n303 2.6005
R2352 VDD.n1453 VDD.n1452 2.6005
R2353 VDD.n1407 VDD.n1404 2.6005
R2354 VDD.n1217 VDD.n1214 2.6005
R2355 VDD.n1206 VDD.n1203 2.6005
R2356 VDD.n419 VDD.n418 2.6005
R2357 VDD.n400 VDD.n399 2.6005
R2358 VDD.n1084 VDD.n1083 2.6005
R2359 VDD.n1064 VDD.n1063 2.6005
R2360 VDD.n1070 VDD.n1066 2.6005
R2361 VDD.n1069 VDD.n1068 2.6005
R2362 VDD.n1073 VDD.n1072 2.6005
R2363 VDD.n529 VDD.n528 2.6005
R2364 VDD.n1109 VDD.n1108 2.6005
R2365 VDD.n1106 VDD.n1105 2.6005
R2366 VDD.n1112 VDD.n1111 2.6005
R2367 VDD.n1117 VDD.n1116 2.6005
R2368 VDD.n638 VDD.n635 2.6005
R2369 VDD.n632 VDD.n631 2.6005
R2370 VDD.n847 VDD.n846 2.6005
R2371 VDD.n803 VDD.n802 2.6005
R2372 VDD.n808 VDD.n805 2.6005
R2373 VDD.n948 VDD.n947 2.6005
R2374 VDD.n1076 VDD.n1075 2.6005
R2375 VDD.n1091 VDD.n1090 2.6005
R2376 VDD.n1088 VDD.n1087 2.6005
R2377 VDD.n1097 VDD.n1081 2.6005
R2378 VDD.n1098 VDD.n1079 2.6005
R2379 VDD.n1094 VDD.n1093 2.6005
R2380 VDD.n371 VDD.n368 2.6005
R2381 VDD.n354 VDD.n351 2.6005
R2382 VDD.n247 VDD.n246 2.6005
R2383 VDD.n237 VDD.n236 2.6005
R2384 VDD.n263 VDD.n262 2.6005
R2385 VDD.n253 VDD.n252 2.6005
R2386 VDD.n198 VDD.n197 2.6005
R2387 VDD.n1629 VDD.n1628 2.6005
R2388 VDD.n225 VDD.n224 2.6005
R2389 VDD.n219 VDD.n218 2.6005
R2390 VDD.n1622 VDD.n1621 2.6005
R2391 VDD.n1625 VDD.n1624 2.6005
R2392 VDD.n256 VDD.n255 2.6005
R2393 VDD.n228 VDD.n227 2.6005
R2394 VDD.n234 VDD.n233 2.6005
R2395 VDD.n250 VDD.n249 2.6005
R2396 VDD.n1613 VDD.n1612 2.6005
R2397 VDD.n1955 VDD.n1954 2.6005
R2398 VDD.n2154 VDD.n2153 2.6005
R2399 VDD.n2617 VDD.n2614 2.6005
R2400 VDD.n1491 VDD.n343 2.59264
R2401 VDD.n1487 VDD.n341 2.59264
R2402 VDD.n1483 VDD.n339 2.59264
R2403 VDD.n1479 VDD.n337 2.59264
R2404 VDD.n1494 VDD.n343 2.59264
R2405 VDD.n1489 VDD.n341 2.59264
R2406 VDD.n1485 VDD.n339 2.59264
R2407 VDD.n1481 VDD.n337 2.59264
R2408 VDD.n1336 VDD.n1335 2.59264
R2409 VDD.n1330 VDD.n390 2.59264
R2410 VDD.n1326 VDD.n388 2.59264
R2411 VDD.n1322 VDD.n386 2.59264
R2412 VDD.n1318 VDD.n384 2.59264
R2413 VDD.n1314 VDD.n382 2.59264
R2414 VDD.n1336 VDD.n379 2.59264
R2415 VDD.n1332 VDD.n390 2.59264
R2416 VDD.n1328 VDD.n388 2.59264
R2417 VDD.n1324 VDD.n386 2.59264
R2418 VDD.n1320 VDD.n384 2.59264
R2419 VDD.n1316 VDD.n382 2.59264
R2420 VDD.n1708 VDD.n1707 2.58448
R2421 VDD.n1489 VDD.n342 2.5167
R2422 VDD.n1485 VDD.n340 2.5167
R2423 VDD.n1481 VDD.n338 2.5167
R2424 VDD.n1477 VDD.n336 2.5167
R2425 VDD.n1491 VDD.n342 2.5167
R2426 VDD.n1487 VDD.n340 2.5167
R2427 VDD.n1483 VDD.n338 2.5167
R2428 VDD.n1479 VDD.n336 2.5167
R2429 VDD.n1332 VDD.n391 2.5167
R2430 VDD.n1328 VDD.n389 2.5167
R2431 VDD.n1324 VDD.n387 2.5167
R2432 VDD.n1320 VDD.n385 2.5167
R2433 VDD.n1316 VDD.n383 2.5167
R2434 VDD.n1335 VDD.n391 2.5167
R2435 VDD.n1330 VDD.n389 2.5167
R2436 VDD.n1326 VDD.n387 2.5167
R2437 VDD.n1322 VDD.n385 2.5167
R2438 VDD.n1318 VDD.n383 2.5167
R2439 VDD.n1725 VDD.t519 2.49842
R2440 VDD.n1709 VDD.n1708 2.49842
R2441 VDD.n563 VDD.n562 2.49842
R2442 VDD.n1495 VDD.n1494 2.47755
R2443 VDD.n1495 VDD.n332 2.47755
R2444 VDD.n1312 VDD.n381 2.47755
R2445 VDD.n1314 VDD.n381 2.47755
R2446 VDD.n2279 VDD.n2278 2.42419
R2447 VDD.n2495 VDD.n2494 2.42419
R2448 VDD.n2267 VDD.n2266 2.42339
R2449 VDD.n2483 VDD.n2482 2.42339
R2450 VDD.n2264 VDD.n2263 2.42315
R2451 VDD.n2480 VDD.n2479 2.42315
R2452 VDD.n2270 VDD.n2269 2.42282
R2453 VDD.n2486 VDD.n2485 2.42282
R2454 VDD.n2276 VDD.n2275 2.42265
R2455 VDD.n2492 VDD.n2491 2.42265
R2456 VDD.n2273 VDD.n2272 2.42222
R2457 VDD.n2489 VDD.n2488 2.42222
R2458 VDD.n2261 VDD.n2260 2.42152
R2459 VDD.n2477 VDD.n2476 2.42152
R2460 VDD.n2258 VDD.n2257 2.41849
R2461 VDD.n2474 VDD.n2473 2.41849
R2462 VDD.n2255 VDD.n2254 2.41843
R2463 VDD.n2471 VDD.n2470 2.41843
R2464 VDD.n2252 VDD.n2251 2.41556
R2465 VDD.n2468 VDD.n2467 2.41556
R2466 VDD.n2249 VDD.n2248 2.41444
R2467 VDD.n2465 VDD.n2464 2.41444
R2468 VDD.n2238 VDD.n2237 2.41251
R2469 VDD.n2454 VDD.n2453 2.41251
R2470 VDD.n2246 VDD.n2245 2.41018
R2471 VDD.n2462 VDD.n2461 2.41018
R2472 VDD.n2235 VDD.n2234 2.41016
R2473 VDD.n2451 VDD.n2450 2.41016
R2474 VDD.n2243 VDD.n2242 2.40994
R2475 VDD.n2459 VDD.n2458 2.40994
R2476 VDD.n2202 VDD.n2201 2.40758
R2477 VDD.n2418 VDD.n2417 2.40758
R2478 VDD.n2208 VDD.n2207 2.40707
R2479 VDD.n2424 VDD.n2423 2.40707
R2480 VDD.n2232 VDD.n2231 2.40667
R2481 VDD.n2448 VDD.n2447 2.40667
R2482 VDD.n2205 VDD.n2204 2.40626
R2483 VDD.n2421 VDD.n2420 2.40626
R2484 VDD.n2211 VDD.n2210 2.40299
R2485 VDD.n2427 VDD.n2426 2.40299
R2486 VDD.n2214 VDD.n2213 2.40275
R2487 VDD.n2430 VDD.n2429 2.40275
R2488 VDD.n2226 VDD.n2225 2.4026
R2489 VDD.n2442 VDD.n2441 2.4026
R2490 VDD.n2229 VDD.n2228 2.40255
R2491 VDD.n2445 VDD.n2444 2.40255
R2492 VDD.n2223 VDD.n2222 2.40212
R2493 VDD.n2439 VDD.n2438 2.40212
R2494 VDD.n2217 VDD.n2216 2.40139
R2495 VDD.n2433 VDD.n2432 2.40139
R2496 VDD.n2220 VDD.n2219 2.40019
R2497 VDD.n2436 VDD.n2435 2.40019
R2498 VDD.n2283 VDD.n2282 2.38241
R2499 VDD.n2499 VDD.n2498 2.38241
R2500 VDD.n992 VDD.n991 2.37611
R2501 VDD.n2671 VDD.n2610 2.35567
R2502 VDD.n2099 VDD.n2098 2.34775
R2503 VDD.n2135 VDD.n3 2.34754
R2504 VDD.n989 VDD.n988 2.34319
R2505 VDD.n988 VDD.n580 2.33916
R2506 VDD.n2592 VDD.n2591 2.33309
R2507 VDD.n2166 VDD.n2165 2.33218
R2508 VDD.n2677 VDD.n2676 2.32106
R2509 VDD.n830 VDD.n829 2.31932
R2510 VDD.n692 VDD.n691 2.29638
R2511 VDD.n692 VDD.n671 2.29115
R2512 VDD.n988 VDD.n987 2.28732
R2513 VDD.n698 VDD.n697 2.2804
R2514 VDD.n1768 VDD.n1767 2.27396
R2515 VDD.n1432 VDD.n1431 2.25904
R2516 VDD.n2179 VDD.n2178 2.25144
R2517 VDD.n1766 VDD.n170 2.25144
R2518 VDD.n704 VDD.n703 2.2505
R2519 VDD.n590 VDD.n588 2.2505
R2520 VDD.n599 VDD.n598 2.2505
R2521 VDD.n627 VDD.n626 2.2505
R2522 VDD.n909 VDD.n746 2.2505
R2523 VDD.n878 VDD.n877 2.2505
R2524 VDD.n759 VDD.n749 2.2505
R2525 VDD.n899 VDD.n743 2.2505
R2526 VDD.n904 VDD.n903 2.2505
R2527 VDD.n2054 VDD.n2053 2.2505
R2528 VDD.n2670 VDD.n2669 2.2505
R2529 VDD.n983 VDD.n581 2.24806
R2530 VDD.n1835 VDD.t890 2.16717
R2531 VDD.n1835 VDD.n1834 2.16717
R2532 VDD.n1794 VDD.t870 2.16717
R2533 VDD.n1794 VDD.n1793 2.16717
R2534 VDD.n1865 VDD.t772 2.16717
R2535 VDD.n1865 VDD.n1864 2.16717
R2536 VDD.n1849 VDD.t1046 2.16717
R2537 VDD.n1849 VDD.n1848 2.16717
R2538 VDD.n158 VDD.t1066 2.16717
R2539 VDD.n158 VDD.n157 2.16717
R2540 VDD.n23 VDD.t843 2.16717
R2541 VDD.n23 VDD.n22 2.16717
R2542 VDD.n98 VDD.t678 2.16717
R2543 VDD.n98 VDD.n97 2.16717
R2544 VDD.n80 VDD.t73 2.16717
R2545 VDD.n80 VDD.n79 2.16717
R2546 VDD.n685 VDD.t557 2.16717
R2547 VDD.n685 VDD.n684 2.16717
R2548 VDD.n674 VDD.t197 2.16717
R2549 VDD.n674 VDD.n673 2.16717
R2550 VDD.n891 VDD.t561 2.16717
R2551 VDD.n891 VDD.n890 2.16717
R2552 VDD.n886 VDD.t205 2.16717
R2553 VDD.n886 VDD.n885 2.16717
R2554 VDD.n2087 VDD.t280 2.16717
R2555 VDD.n2087 VDD.n2086 2.16717
R2556 VDD.n2107 VDD.t1022 2.16717
R2557 VDD.n2107 VDD.n2106 2.16717
R2558 VDD.n2597 VDD.t371 2.16717
R2559 VDD.n2597 VDD.n2596 2.16717
R2560 VDD.n2651 VDD.t1106 2.16717
R2561 VDD.n2651 VDD.n2650 2.16717
R2562 VDD.n733 VDD.n594 2.05248
R2563 VDD.t188 VDD.n647 2.05248
R2564 VDD.n717 VDD.t46 2.05248
R2565 VDD.n796 VDD.t17 2.05248
R2566 VDD.n1243 VDD.n1194 2.04683
R2567 VDD.n1239 VDD.n1194 2.04625
R2568 VDD.n1534 VDD.n285 2.04615
R2569 VDD.n1538 VDD.n285 2.04615
R2570 VDD.n1712 VDD.n1711 2.00622
R2571 VDD.n1711 VDD.n1648 2.00565
R2572 VDD.n1238 VDD.n1198 1.94801
R2573 VDD.n1235 VDD.n1198 1.94746
R2574 VDD.n1539 VDD.n286 1.94734
R2575 VDD.n1542 VDD.n286 1.94734
R2576 VDD.n693 VDD.n692 1.94241
R2577 VDD.n967 VDD.n933 1.9255
R2578 VDD.n1496 VDD.n1495 1.91272
R2579 VDD.n1337 VDD.n381 1.91272
R2580 VDD.n2239 VDD.n2199 1.91067
R2581 VDD.n2455 VDD.n2415 1.91067
R2582 VDD.n1448 VDD.n1447 1.8985
R2583 VDD.n1496 VDD.n336 1.89315
R2584 VDD.n1496 VDD.n338 1.89315
R2585 VDD.n1496 VDD.n340 1.89315
R2586 VDD.n1496 VDD.n342 1.89315
R2587 VDD.n1337 VDD.n383 1.89315
R2588 VDD.n1337 VDD.n385 1.89315
R2589 VDD.n1337 VDD.n387 1.89315
R2590 VDD.n1337 VDD.n389 1.89315
R2591 VDD.n1337 VDD.n391 1.89315
R2592 VDD.n325 VDD.n280 1.87282
R2593 VDD.n481 VDD.n478 1.87282
R2594 VDD.n1564 VDD.n280 1.87228
R2595 VDD.n478 VDD.n477 1.87228
R2596 VDD.n1470 VDD.n333 1.8617
R2597 VDD.n1472 VDD.n333 1.8617
R2598 VDD.n1496 VDD.n337 1.85518
R2599 VDD.n1496 VDD.n339 1.85518
R2600 VDD.n1496 VDD.n341 1.85518
R2601 VDD.n1496 VDD.n343 1.85518
R2602 VDD.n1337 VDD.n382 1.85518
R2603 VDD.n1337 VDD.n384 1.85518
R2604 VDD.n1337 VDD.n386 1.85518
R2605 VDD.n1337 VDD.n388 1.85518
R2606 VDD.n1337 VDD.n390 1.85518
R2607 VDD.n1337 VDD.n1336 1.85518
R2608 VDD.n663 VDD.n661 1.85344
R2609 VDD.n705 VDD.n661 1.85344
R2610 VDD.n823 VDD.n822 1.85344
R2611 VDD.n824 VDD.n823 1.85344
R2612 VDD.n1230 VDD.n1208 1.83567
R2613 VDD.n1226 VDD.n1208 1.83513
R2614 VDD.n1547 VDD.n288 1.835
R2615 VDD.n1551 VDD.n288 1.835
R2616 VDD.n1225 VDD.n1224 1.82979
R2617 VDD.n1224 VDD.n1223 1.82925
R2618 VDD.n1552 VDD.n289 1.82912
R2619 VDD.n290 VDD.n289 1.82912
R2620 VDD VDD.n679 1.82452
R2621 VDD.n1387 VDD.n356 1.80965
R2622 VDD.n1387 VDD.n1386 1.80912
R2623 VDD.n645 VDD.n622 1.7505
R2624 VDD.n1245 VDD.n1244 1.69304
R2625 VDD.n1234 VDD.n1201 1.69304
R2626 VDD.n1212 VDD.n1211 1.69304
R2627 VDD.n1211 VDD.n485 1.69252
R2628 VDD.n1231 VDD.n1201 1.69252
R2629 VDD.n1246 VDD.n1245 1.69252
R2630 VDD.n1543 VDD.n287 1.69238
R2631 VDD.n1530 VDD.n284 1.69238
R2632 VDD.n1546 VDD.n287 1.69238
R2633 VDD.n1533 VDD.n284 1.69238
R2634 VDD.n1773 VDD.n1772 1.68275
R2635 VDD.n1026 VDD.n1025 1.66029
R2636 VDD.n1025 VDD.n1024 1.65977
R2637 VDD.n1019 VDD.n568 1.65963
R2638 VDD.n1017 VDD.n1016 1.65963
R2639 VDD.n1011 VDD.n572 1.65963
R2640 VDD.n1009 VDD.n1008 1.65963
R2641 VDD.n1003 VDD.n576 1.65963
R2642 VDD.n1001 VDD.n1000 1.65963
R2643 VDD.n995 VDD.n994 1.65963
R2644 VDD.n568 VDD.n565 1.65963
R2645 VDD.n1018 VDD.n1017 1.65963
R2646 VDD.n572 VDD.n569 1.65963
R2647 VDD.n1010 VDD.n1009 1.65963
R2648 VDD.n576 VDD.n573 1.65963
R2649 VDD.n1002 VDD.n1001 1.65963
R2650 VDD.n994 VDD.n577 1.65963
R2651 VDD.n1981 VDD.n1978 1.64018
R2652 VDD.n14 VDD.n11 1.64018
R2653 VDD.n1085 VDD.n537 1.5755
R2654 VDD.n975 VDD.n920 1.5755
R2655 VDD.n1617 VDD.n1616 1.5755
R2656 VDD.n1101 VDD.n1100 1.57159
R2657 VDD.n258 VDD.n257 1.57159
R2658 VDD.n1339 VDD.n1338 1.54574
R2659 VDD.n1498 VDD.n1497 1.52056
R2660 VDD.n1475 VDD.n335 1.52041
R2661 VDD.n1310 VDD.n380 1.52041
R2662 VDD.n972 VDD.n934 1.5005
R2663 VDD.n1118 VDD.n514 1.49724
R2664 VDD.n222 VDD.n173 1.49724
R2665 VDD.n929 VDD.n922 1.488
R2666 VDD.n1944 VDD.n1943 1.48015
R2667 VDD.n915 VDD.n914 1.42211
R2668 VDD.n883 VDD.n882 1.42018
R2669 VDD.n620 VDD.n595 1.4005
R2670 VDD.n2239 VDD.n2238 1.38687
R2671 VDD.n2455 VDD.n2454 1.38687
R2672 VDD.n1561 VDD.n1560 1.3744
R2673 VDD.n1558 VDD.n1557 1.3744
R2674 VDD.n966 VDD.n965 1.36849
R2675 VDD.n1474 VDD.n1455 1.35142
R2676 VDD.n2280 VDD.n2279 1.34148
R2677 VDD.n2496 VDD.n2495 1.34148
R2678 VDD.n2672 VDD.n2671 1.25782
R2679 VDD.n2284 VDD.n2283 1.25144
R2680 VDD.n2500 VDD.n2499 1.25144
R2681 VDD.t970 VDD.t666 1.24946
R2682 VDD.t672 VDD.t943 1.24946
R2683 VDD.n881 VDD.n833 1.2474
R2684 VDD.n2676 VDD.n2675 1.19777
R2685 VDD.n1560 VDD.n1559 1.1854
R2686 VDD.n1559 VDD.n1558 1.1854
R2687 VDD.n2674 VDD.n2673 1.17139
R2688 VDD.n991 VDD.n990 1.14837
R2689 VDD.n2172 VDD.n2171 1.13742
R2690 VDD.n2100 VDD.n2078 1.13054
R2691 VDD.n2171 VDD.n3 1.12799
R2692 VDD.n2098 VDD.n2097 1.12796
R2693 VDD.n703 VDD.n702 1.1255
R2694 VDD.n625 VDD.n588 1.1255
R2695 VDD.n759 VDD.n758 1.1255
R2696 VDD.n909 VDD.n908 1.1255
R2697 VDD.n972 VDD.n971 1.1255
R2698 VDD.n984 VDD.n983 1.1255
R2699 VDD.n2134 VDD.n2133 1.1255
R2700 VDD.n2164 VDD.n2163 1.1255
R2701 VDD.n2136 VDD.n2135 1.1255
R2702 VDD.n2384 VDD.n2383 1.1255
R2703 VDD.n2591 VDD.n2590 1.1255
R2704 VDD.n2170 VDD.n2169 1.1255
R2705 VDD.n2168 VDD.n2167 1.1255
R2706 VDD.n2102 VDD.n2101 1.1255
R2707 VDD.n2100 VDD.n2099 1.1255
R2708 VDD.n763 VDD.n752 1.12549
R2709 VDD.n1767 VDD.n169 1.11762
R2710 VDD.n1497 VDD.n1496 1.08825
R2711 VDD.n1496 VDD.n335 1.08806
R2712 VDD.n1337 VDD.n380 1.08806
R2713 VDD.n1338 VDD.n1337 1.07146
R2714 VDD.n1103 VDD.n1102 1.06485
R2715 VDD.n1114 VDD.n1113 1.06485
R2716 VDD.n1099 VDD.n1077 1.06485
R2717 VDD.n1096 VDD.n1095 1.06485
R2718 VDD.n260 VDD.n259 1.06485
R2719 VDD.n1626 VDD.n216 1.06485
R2720 VDD.n1619 VDD.n1618 1.06485
R2721 VDD.n1615 VDD.n1614 1.06485
R2722 VDD.n1974 VDD.n1967 1.06047
R2723 VDD.n2014 VDD.n2013 1.05511
R2724 VDD.n655 VDD.n642 1.0505
R2725 VDD.n872 VDD.n837 1.0505
R2726 VDD.n2674 VDD.n2592 1.04546
R2727 VDD.n1975 VDD.n1974 1.03869
R2728 VDD VDD.n2017 1.02937
R2729 VDD.n1118 VDD.n536 1.01789
R2730 VDD.n514 VDD.n504 1.01789
R2731 VDD.n222 VDD.n221 1.01789
R2732 VDD.n1610 VDD.n173 1.01789
R2733 VDD.n2240 VDD.n2239 0.996686
R2734 VDD.n2456 VDD.n2455 0.996686
R2735 VDD.n1342 VDD.n1341 0.984049
R2736 VDD.n650 VDD.n642 0.963
R2737 VDD.n884 VDD.n883 0.950899
R2738 VDD.n2044 VDD.n2043 0.93487
R2739 VDD.n993 VDD.n992 0.931466
R2740 VDD.n727 VDD.n726 0.927241
R2741 VDD.n584 VDD.n579 0.92659
R2742 VDD.n834 VDD.n832 0.925561
R2743 VDD.n742 VDD.n585 0.904541
R2744 VDD.n2535 VDD.n2534 0.9005
R2745 VDD.n2524 VDD.n2523 0.9005
R2746 VDD.n2590 VDD.n2589 0.9005
R2747 VDD.n831 VDD.n830 0.899617
R2748 VDD.n698 VDD.n693 0.898206
R2749 VDD.n904 VDD.n884 0.897926
R2750 VDD.n913 VDD.n743 0.897926
R2751 VDD.n1772 VDD.n1771 0.872556
R2752 VDD.n2066 VDD.n2024 0.867239
R2753 VDD.n2062 VDD.n2061 0.847535
R2754 VDD.t952 VDD.t995 0.833139
R2755 VDD.t940 VDD.t952 0.833139
R2756 VDD.t958 VDD.t946 0.833139
R2757 VDD.t949 VDD.t990 0.833139
R2758 VDD.t990 VDD.t937 0.833139
R2759 VDD.n990 VDD 0.830218
R2760 VDD.n2286 VDD.n2284 0.828172
R2761 VDD.n2502 VDD.n2500 0.828172
R2762 VDD.n1919 VDD.n1918 0.810896
R2763 VDD.n1942 VDD.n1791 0.810896
R2764 VDD.n1925 VDD.n1844 0.809707
R2765 VDD.n1070 VDD.n1069 0.802674
R2766 VDD.n1109 VDD.n1106 0.802674
R2767 VDD.n1091 VDD.n1088 0.802674
R2768 VDD.n1098 VDD.n1097 0.802674
R2769 VDD.n247 VDD.n237 0.802674
R2770 VDD.n1625 VDD.n1622 0.802674
R2771 VDD.n256 VDD.n228 0.802674
R2772 VDD.n250 VDD.n234 0.802674
R2773 VDD.n1998 VDD.n1997 0.798761
R2774 VDD.n1952 VDD.n1951 0.798761
R2775 VDD.n467 VDD.n466 0.795217
R2776 VDD.n914 VDD.n913 0.792748
R2777 VDD.n2078 VDD.n2077 0.776876
R2778 VDD.n1025 VDD.n564 0.746922
R2779 VDD.n568 VDD.n564 0.746686
R2780 VDD.n1017 VDD.n564 0.746686
R2781 VDD.n572 VDD.n564 0.746686
R2782 VDD.n1009 VDD.n564 0.746686
R2783 VDD.n576 VDD.n564 0.746686
R2784 VDD.n1001 VDD.n564 0.746686
R2785 VDD.n994 VDD.n564 0.746686
R2786 VDD.n2052 VDD.n2051 0.735716
R2787 VDD.n1201 VDD.n479 0.730547
R2788 VDD.n1211 VDD.n479 0.730547
R2789 VDD.n1245 VDD.n479 0.730547
R2790 VDD.n1559 VDD.n287 0.73031
R2791 VDD.n1559 VDD.n284 0.73031
R2792 VDD.n688 VDD.n687 0.7187
R2793 VDD.n1388 VDD.n1387 0.674731
R2794 VDD.n1224 VDD.n479 0.662176
R2795 VDD.n1559 VDD.n289 0.661938
R2796 VDD.n1770 VDD.n170 0.660673
R2797 VDD.n1208 VDD.n479 0.659239
R2798 VDD.n1559 VDD.n288 0.659
R2799 VDD.n2325 VDD.t502 0.6505
R2800 VDD.n2325 VDD.n2324 0.6505
R2801 VDD.n2322 VDD.t137 0.6505
R2802 VDD.n2322 VDD.n2321 0.6505
R2803 VDD.n2318 VDD.t135 0.6505
R2804 VDD.n2318 VDD.n2317 0.6505
R2805 VDD.n2314 VDD.t1047 0.6505
R2806 VDD.n2314 VDD.n2313 0.6505
R2807 VDD.n2311 VDD.t1084 0.6505
R2808 VDD.n2311 VDD.n2310 0.6505
R2809 VDD.n2307 VDD.t677 0.6505
R2810 VDD.n2307 VDD.n2306 0.6505
R2811 VDD.n2304 VDD.t880 0.6505
R2812 VDD.n2304 VDD.n2303 0.6505
R2813 VDD.n2302 VDD.t214 0.6505
R2814 VDD.n2302 VDD.n2301 0.6505
R2815 VDD.n2193 VDD.t637 0.6505
R2816 VDD.n2193 VDD.n2192 0.6505
R2817 VDD.n2195 VDD.t601 0.6505
R2818 VDD.n2195 VDD.n2194 0.6505
R2819 VDD.n2197 VDD.t600 0.6505
R2820 VDD.n2197 VDD.n2196 0.6505
R2821 VDD.n2266 VDD.t602 0.6505
R2822 VDD.n2266 VDD.n2265 0.6505
R2823 VDD.n2242 VDD.t489 0.6505
R2824 VDD.n2242 VDD.n2241 0.6505
R2825 VDD.n2245 VDD.t463 0.6505
R2826 VDD.n2245 VDD.n2244 0.6505
R2827 VDD.n2248 VDD.t457 0.6505
R2828 VDD.n2248 VDD.n2247 0.6505
R2829 VDD.n2251 VDD.t445 0.6505
R2830 VDD.n2251 VDD.n2250 0.6505
R2831 VDD.n2254 VDD.t443 0.6505
R2832 VDD.n2254 VDD.n2253 0.6505
R2833 VDD.n2257 VDD.t650 0.6505
R2834 VDD.n2257 VDD.n2256 0.6505
R2835 VDD.n2260 VDD.t483 0.6505
R2836 VDD.n2260 VDD.n2259 0.6505
R2837 VDD.n2263 VDD.t481 0.6505
R2838 VDD.n2263 VDD.n2262 0.6505
R2839 VDD.n2269 VDD.t654 0.6505
R2840 VDD.n2269 VDD.n2268 0.6505
R2841 VDD.n2272 VDD.t645 0.6505
R2842 VDD.n2272 VDD.n2271 0.6505
R2843 VDD.n2275 VDD.t462 0.6505
R2844 VDD.n2275 VDD.n2274 0.6505
R2845 VDD.n2278 VDD.t456 0.6505
R2846 VDD.n2278 VDD.n2277 0.6505
R2847 VDD.n2282 VDD.n2281 0.6505
R2848 VDD.n2201 VDD.t656 0.6505
R2849 VDD.n2201 VDD.n2200 0.6505
R2850 VDD.n2204 VDD.t647 0.6505
R2851 VDD.n2204 VDD.n2203 0.6505
R2852 VDD.n2207 VDD.t644 0.6505
R2853 VDD.n2207 VDD.n2206 0.6505
R2854 VDD.n2210 VDD.t480 0.6505
R2855 VDD.n2210 VDD.n2209 0.6505
R2856 VDD.n2213 VDD.t479 0.6505
R2857 VDD.n2213 VDD.n2212 0.6505
R2858 VDD.n2216 VDD.t599 0.6505
R2859 VDD.n2216 VDD.n2215 0.6505
R2860 VDD.n2219 VDD.t651 0.6505
R2861 VDD.n2219 VDD.n2218 0.6505
R2862 VDD.n2222 VDD.t649 0.6505
R2863 VDD.n2222 VDD.n2221 0.6505
R2864 VDD.n2225 VDD.t640 0.6505
R2865 VDD.n2225 VDD.n2224 0.6505
R2866 VDD.n2228 VDD.t604 0.6505
R2867 VDD.n2228 VDD.n2227 0.6505
R2868 VDD.n2231 VDD.t441 0.6505
R2869 VDD.n2231 VDD.n2230 0.6505
R2870 VDD.n2234 VDD.t646 0.6505
R2871 VDD.n2234 VDD.n2233 0.6505
R2872 VDD.n2237 VDD.t643 0.6505
R2873 VDD.n2237 VDD.n2236 0.6505
R2874 VDD.n2299 VDD.t507 0.6505
R2875 VDD.n2299 VDD.n2298 0.6505
R2876 VDD.n2191 VDD.t648 0.6505
R2877 VDD.n2191 VDD.n2190 0.6505
R2878 VDD.n2568 VDD.t811 0.6505
R2879 VDD.n2568 VDD.n2567 0.6505
R2880 VDD.n2565 VDD.t146 0.6505
R2881 VDD.n2565 VDD.n2564 0.6505
R2882 VDD.n2561 VDD.t144 0.6505
R2883 VDD.n2561 VDD.n2560 0.6505
R2884 VDD.n2557 VDD.t39 0.6505
R2885 VDD.n2557 VDD.n2556 0.6505
R2886 VDD.n2554 VDD.t245 0.6505
R2887 VDD.n2554 VDD.n2553 0.6505
R2888 VDD.n2550 VDD.t1074 0.6505
R2889 VDD.n2550 VDD.n2549 0.6505
R2890 VDD.n2547 VDD.t1073 0.6505
R2891 VDD.n2547 VDD.n2546 0.6505
R2892 VDD.n2407 VDD.t706 0.6505
R2893 VDD.n2407 VDD.n2406 0.6505
R2894 VDD.n2409 VDD.t927 0.6505
R2895 VDD.n2409 VDD.n2408 0.6505
R2896 VDD.n2411 VDD.t826 0.6505
R2897 VDD.n2411 VDD.n2410 0.6505
R2898 VDD.n2413 VDD.t79 0.6505
R2899 VDD.n2413 VDD.n2412 0.6505
R2900 VDD.n2482 VDD.t682 0.6505
R2901 VDD.n2482 VDD.n2481 0.6505
R2902 VDD.n2458 VDD.t1018 0.6505
R2903 VDD.n2458 VDD.n2457 0.6505
R2904 VDD.n2461 VDD.t1011 0.6505
R2905 VDD.n2461 VDD.n2460 0.6505
R2906 VDD.n2464 VDD.t683 0.6505
R2907 VDD.n2464 VDD.n2463 0.6505
R2908 VDD.n2467 VDD.t853 0.6505
R2909 VDD.n2467 VDD.n2466 0.6505
R2910 VDD.n2470 VDD.t1020 0.6505
R2911 VDD.n2470 VDD.n2469 0.6505
R2912 VDD.n2473 VDD.t609 0.6505
R2913 VDD.n2473 VDD.n2472 0.6505
R2914 VDD.n2476 VDD.t607 0.6505
R2915 VDD.n2476 VDD.n2475 0.6505
R2916 VDD.n2479 VDD.t932 0.6505
R2917 VDD.n2479 VDD.n2478 0.6505
R2918 VDD.n2485 VDD.t878 0.6505
R2919 VDD.n2485 VDD.n2484 0.6505
R2920 VDD.n2488 VDD.t1017 0.6505
R2921 VDD.n2488 VDD.n2487 0.6505
R2922 VDD.n2491 VDD.t1009 0.6505
R2923 VDD.n2491 VDD.n2490 0.6505
R2924 VDD.n2494 VDD.t726 0.6505
R2925 VDD.n2494 VDD.n2493 0.6505
R2926 VDD.n2498 VDD.n2497 0.6505
R2927 VDD.n2417 VDD.t856 0.6505
R2928 VDD.n2417 VDD.n2416 0.6505
R2929 VDD.n2420 VDD.t814 0.6505
R2930 VDD.n2420 VDD.n2419 0.6505
R2931 VDD.n2423 VDD.t1019 0.6505
R2932 VDD.n2423 VDD.n2422 0.6505
R2933 VDD.n2426 VDD.t608 0.6505
R2934 VDD.n2426 VDD.n2425 0.6505
R2935 VDD.n2429 VDD.t922 0.6505
R2936 VDD.n2429 VDD.n2428 0.6505
R2937 VDD.n2432 VDD.t77 0.6505
R2938 VDD.n2432 VDD.n2431 0.6505
R2939 VDD.n2435 VDD.t75 0.6505
R2940 VDD.n2435 VDD.n2434 0.6505
R2941 VDD.n2438 VDD.t852 0.6505
R2942 VDD.n2438 VDD.n2437 0.6505
R2943 VDD.n2441 VDD.t1016 0.6505
R2944 VDD.n2441 VDD.n2440 0.6505
R2945 VDD.n2444 VDD.t685 0.6505
R2946 VDD.n2444 VDD.n2443 0.6505
R2947 VDD.n2447 VDD.t855 0.6505
R2948 VDD.n2447 VDD.n2446 0.6505
R2949 VDD.n2450 VDD.t1021 0.6505
R2950 VDD.n2450 VDD.n2449 0.6505
R2951 VDD.n2453 VDD.t875 0.6505
R2952 VDD.n2453 VDD.n2452 0.6505
R2953 VDD.n2394 VDD.t212 0.6505
R2954 VDD.n2394 VDD.n2393 0.6505
R2955 VDD.n2405 VDD.t142 0.6505
R2956 VDD.n2405 VDD.n2404 0.6505
R2957 VDD.n1496 VDD.n333 0.645651
R2958 VDD VDD.n2 0.642616
R2959 VDD.n1838 VDD.n1837 0.6395
R2960 VDD.n1797 VDD.n1795 0.6395
R2961 VDD.n1868 VDD.n1867 0.6395
R2962 VDD.n1852 VDD.n1850 0.6395
R2963 VDD.n161 VDD.n160 0.6395
R2964 VDD.n26 VDD.n24 0.6395
R2965 VDD.n101 VDD.n100 0.6395
R2966 VDD.n83 VDD.n81 0.6395
R2967 VDD.n677 VDD.n676 0.6395
R2968 VDD.n894 VDD.n892 0.6395
R2969 VDD.n889 VDD.n887 0.6395
R2970 VDD.n2090 VDD.n2089 0.6395
R2971 VDD.n2110 VDD.n2108 0.6395
R2972 VDD.n2600 VDD.n2599 0.6395
R2973 VDD.n2654 VDD.n2652 0.6395
R2974 VDD.n1965 VDD.n1964 0.626871
R2975 VDD.n615 VDD.n595 0.613
R2976 VDD.n1198 VDD.n479 0.60307
R2977 VDD.n1559 VDD.n286 0.602829
R2978 VDD.n166 VDD.n165 0.598557
R2979 VDD.n106 VDD.n105 0.598557
R2980 VDD.n1805 VDD.n1804 0.597767
R2981 VDD.n1860 VDD.n1859 0.597767
R2982 VDD.n2119 VDD.n2118 0.597767
R2983 VDD.n2663 VDD.n2662 0.597767
R2984 VDD.n1500 VDD.n1499 0.593699
R2985 VDD.n1771 VDD.n169 0.587674
R2986 VDD.n1964 VDD.n1963 0.586952
R2987 VDD.n1064 VDD.n1061 0.581587
R2988 VDD.n1073 VDD.n509 0.581587
R2989 VDD.n1126 VDD.n529 0.581587
R2990 VDD.n1076 VDD.n499 0.581587
R2991 VDD.n1591 VDD.n263 0.581587
R2992 VDD.n253 VDD.n179 0.581587
R2993 VDD.n1743 VDD.n198 0.581587
R2994 VDD.n1729 VDD.n1629 0.581587
R2995 VDD.n2001 VDD.n2000 0.577192
R2996 VDD.n2051 VDD.n2049 0.576883
R2997 VDD.n1711 VDD.n1710 0.573969
R2998 VDD.n1454 VDD.n1448 0.569476
R2999 VDD.n1194 VDD.n479 0.553668
R3000 VDD.n1559 VDD.n285 0.553425
R3001 VDD.n2024 VDD.n2023 0.5405
R3002 VDD.n2023 VDD.n2022 0.5405
R3003 VDD.n914 VDD.n742 0.539532
R3004 VDD.n1958 VDD.n1957 0.539417
R3005 VDD.n2002 VDD.n1999 0.538543
R3006 VDD.n1555 VDD.n298 0.536587
R3007 VDD.n305 VDD.n304 0.536587
R3008 VDD.n311 VDD.n310 0.536587
R3009 VDD.n1221 VDD.n1217 0.536587
R3010 VDD.n1207 VDD.n1206 0.536587
R3011 VDD.n1197 VDD.n1196 0.536587
R3012 VDD.n1956 VDD.n1955 0.536587
R3013 VDD.n1772 VDD.n168 0.531381
R3014 VDD.n929 VDD.n919 0.5255
R3015 VDD.n1967 VDD.n1966 0.514462
R3016 VDD.n1966 VDD.n1965 0.50421
R3017 VDD.n2008 VDD.n1981 0.502171
R3018 VDD.n2367 VDD.n2366 0.500448
R3019 VDD.n15 VDD.n14 0.500214
R3020 VDD.n2076 VDD.n2075 0.497736
R3021 VDD.n2675 VDD.n2674 0.496915
R3022 VDD.n1471 VDD.n1456 0.495796
R3023 VDD.n2682 VDD.n2175 0.489544
R3024 VDD VDD.n632 0.485717
R3025 VDD VDD.n638 0.485717
R3026 VDD.n107 VDD.n77 0.484683
R3027 VDD.n49 VDD.n36 0.475256
R3028 VDD VDD.n354 0.474784
R3029 VDD.n1926 VDD.n1843 0.470115
R3030 VDD.n167 VDD.n19 0.469543
R3031 VDD.n1118 VDD.n1117 0.467817
R3032 VDD.n225 VDD.n222 0.467817
R3033 VDD.n69 VDD.n38 0.46684
R3034 VDD.n1094 VDD.n504 0.466777
R3035 VDD.n1613 VDD.n1610 0.466777
R3036 VDD.n59 VDD.n37 0.464904
R3037 VDD.n1923 VDD.n1922 0.464346
R3038 VDD.n882 VDD.n881 0.462817
R3039 VDD.n1921 VDD.n1920 0.462038
R3040 VDD.n1941 VDD.n1805 0.461509
R3041 VDD.n148 VDD.n147 0.460249
R3042 VDD.n138 VDD.n20 0.452047
R3043 VDD.n151 VDD.n35 0.450132
R3044 VDD.n1106 VDD.n1103 0.440717
R3045 VDD.n1626 VDD.n1625 0.440717
R3046 VDD.n979 VDD.n920 0.438
R3047 VDD.n1999 VDD.n1998 0.430935
R3048 VDD.n231 VDD.n173 0.430935
R3049 VDD.n1084 VDD.n514 0.430935
R3050 VDD.n1112 VDD.n536 0.430935
R3051 VDD.n221 VDD.n219 0.430935
R3052 VDD.n1955 VDD.n1952 0.430935
R3053 VDD.n2075 VDD.n2074 0.429324
R3054 VDD.n2074 VDD.n2073 0.429324
R3055 VDD.n1113 VDD.n1109 0.421152
R3056 VDD.n1095 VDD.n1094 0.421152
R3057 VDD.n1622 VDD.n1619 0.421152
R3058 VDD.n1614 VDD.n1613 0.421152
R3059 VDD.n1917 VDD.n1916 0.420582
R3060 VDD.n1892 VDD.n1860 0.420066
R3061 VDD.n2668 VDD.n2624 0.419346
R3062 VDD.n2666 VDD.n2640 0.419346
R3063 VDD.n2664 VDD.n2663 0.419346
R3064 VDD.n2610 VDD.n2605 0.419346
R3065 VDD.n1915 VDD.n1914 0.418275
R3066 VDD.t973 VDD.t669 0.41682
R3067 VDD.t669 VDD.t965 0.41682
R3068 VDD.t983 VDD.t934 0.41682
R3069 VDD.t171 VDD.n502 0.41682
R3070 VDD.t784 VDD.t955 0.41682
R3071 VDD.t978 VDD.t784 0.41682
R3072 VDD.n1906 VDD.n1873 0.412505
R3073 VDD.n1276 VDD.n1275 0.405977
R3074 VDD.n1527 VDD.n313 0.405977
R3075 VDD.n2078 VDD 0.405532
R3076 VDD.n1119 VDD.n1118 0.394968
R3077 VDD.n1169 VDD.n504 0.394968
R3078 VDD.n222 VDD.n220 0.394968
R3079 VDD.n1610 VDD.n1609 0.394968
R3080 VDD.n1764 VDD.n173 0.39039
R3081 VDD.n1077 VDD.n1076 0.389848
R3082 VDD.n263 VDD.n260 0.389848
R3083 VDD.n1813 VDD.n1812 0.389323
R3084 VDD.n1891 VDD.n1890 0.389323
R3085 VDD.n130 VDD.n129 0.389323
R3086 VDD.n41 VDD.n40 0.389323
R3087 VDD.n425 VDD.n424 0.389323
R3088 VDD.n954 VDD.n953 0.389323
R3089 VDD.n1378 VDD.n1375 0.389323
R3090 VDD.n2124 VDD.n2122 0.389323
R3091 VDD.n2645 VDD.n2643 0.389323
R3092 VDD.n1843 VDD.n1842 0.388557
R3093 VDD.n1873 VDD.n1872 0.388557
R3094 VDD.n2095 VDD.n2094 0.388557
R3095 VDD.n2605 VDD.n2604 0.388557
R3096 VDD.n34 VDD.n33 0.387767
R3097 VDD.n91 VDD.n90 0.387767
R3098 VDD.n1431 VDD.n1397 0.376152
R3099 VDD.n1432 VDD.n1394 0.376152
R3100 VDD.n443 VDD.n405 0.376152
R3101 VDD.n667 VDD.n666 0.376152
R3102 VDD.n610 VDD.n605 0.376152
R3103 VDD.n876 VDD.n835 0.376152
R3104 VDD.n787 VDD.n783 0.376152
R3105 VDD.n787 VDD.n786 0.376152
R3106 VDD.n1365 VDD.n362 0.376152
R3107 VDD.n1423 VDD.n1407 0.374196
R3108 VDD.n432 VDD.n419 0.374196
R3109 VDD.n401 VDD.n400 0.374196
R3110 VDD.n862 VDD.n847 0.374196
R3111 VDD.n809 VDD.n803 0.374196
R3112 VDD.n809 VDD.n808 0.374196
R3113 VDD.n961 VDD.n948 0.374196
R3114 VDD.n372 VDD.n371 0.374196
R3115 VDD.n1441 VDD.n1388 0.372931
R3116 VDD.n1311 VDD.n467 0.359918
R3117 VDD.n1053 VDD.n536 0.358543
R3118 VDD.n1152 VDD.n514 0.358543
R3119 VDD.n221 VDD.n208 0.358543
R3120 VDD.n922 VDD.n921 0.350287
R3121 VDD.n1101 VDD.n1070 0.327239
R3122 VDD.n257 VDD.n256 0.327239
R3123 VDD.n1088 VDD.n1077 0.323326
R3124 VDD.n1099 VDD.n1098 0.323326
R3125 VDD.n260 VDD.n247 0.323326
R3126 VDD.n259 VDD.n250 0.323326
R3127 VDD.n1959 VDD.n1958 0.319855
R3128 VDD.n443 VDD.n442 0.312794
R3129 VDD.n1616 VDD.n231 0.311587
R3130 VDD.n1085 VDD.n1084 0.311587
R3131 VDD.n1366 VDD.n1365 0.306039
R3132 VDD.n2346 VDD.n2345 0.299037
R3133 VDD.n1961 VDD.n1788 0.292274
R3134 VDD.n1964 VDD.n17 0.292274
R3135 VDD.n1965 VDD.n7 0.292274
R3136 VDD.n1966 VDD.n6 0.292274
R3137 VDD.n998 VDD.n578 0.292144
R3138 VDD.n1006 VDD.n574 0.292144
R3139 VDD.n1013 VDD.n570 0.292144
R3140 VDD.n1113 VDD.n1112 0.292022
R3141 VDD.n1117 VDD.n1114 0.292022
R3142 VDD.n1095 VDD.n1091 0.292022
R3143 VDD.n1097 VDD.n1096 0.292022
R3144 VDD.n1614 VDD.n237 0.292022
R3145 VDD.n1618 VDD.n225 0.292022
R3146 VDD.n1619 VDD.n219 0.292022
R3147 VDD.n1615 VDD.n234 0.292022
R3148 VDD.n1669 VDD.n1668 0.291683
R3149 VDD.n1681 VDD.n1662 0.291683
R3150 VDD.n1704 VDD.n1655 0.291683
R3151 VDD.n1021 VDD.n566 0.288544
R3152 VDD.n1694 VDD.n1687 0.288083
R3153 VDD.n1671 VDD.n1667 0.284207
R3154 VDD.n1069 VDD.n537 0.278326
R3155 VDD.n1617 VDD.n228 0.278326
R3156 VDD.n1922 VDD.n1843 0.276269
R3157 VDD.n1915 VDD.n1873 0.276269
R3158 VDD.n152 VDD.n34 0.276269
R3159 VDD.n92 VDD.n91 0.276269
R3160 VDD.n1103 VDD.n1064 0.272457
R3161 VDD.n1102 VDD.n529 0.272457
R3162 VDD.n216 VDD.n198 0.272457
R3163 VDD.n1629 VDD.n1626 0.272457
R3164 VDD.n1100 VDD.n1073 0.266587
R3165 VDD.n258 VDD.n253 0.266587
R3166 VDD.n1536 VDD.n312 0.266523
R3167 VDD.n2280 VDD.n2240 0.265556
R3168 VDD.n2496 VDD.n2456 0.265556
R3169 VDD.n2511 VDD.n2509 0.265378
R3170 VDD.n1241 VDD.n1195 0.26536
R3171 VDD.n293 VDD.n291 0.264528
R3172 VDD.n1219 VDD.n1218 0.263373
R3173 VDD.n732 VDD.n622 0.263
R3174 VDD.n307 VDD.n306 0.262011
R3175 VDD.n1921 VDD.n1805 0.261269
R3176 VDD.n1916 VDD.n1860 0.261269
R3177 VDD.n166 VDD.n153 0.261269
R3178 VDD.n106 VDD.n93 0.261269
R3179 VDD.n1200 VDD.n1199 0.260887
R3180 VDD.n1549 VDD.n299 0.257984
R3181 VDD.n1228 VDD.n1209 0.257526
R3182 VDD.n2292 VDD.n2290 0.255134
R3183 VDD.n2508 VDD.n2506 0.255134
R3184 VDD.n1502 VDD.n1501 0.25389
R3185 VDD.n928 VDD.n927 0.253803
R3186 VDD.n993 VDD.n558 0.252505
R3187 VDD.n690 VDD.n689 0.252091
R3188 VDD.n1341 VDD.n376 0.248505
R3189 VDD.n1907 VDD.n1906 0.243962
R3190 VDD.n2001 VDD.n1986 0.238747
R3191 VDD.n1515 VDD.n326 0.238241
R3192 VDD.n1914 VDD.n1913 0.238192
R3193 VDD.n1295 VDD.n1294 0.238069
R3194 VDD.n1293 VDD.n475 0.237294
R3195 VDD.n1414 VDD.n1412 0.237044
R3196 VDD.n855 VDD.n853 0.237044
R3197 VDD.n1346 VDD.n1345 0.237044
R3198 VDD.n1917 VDD.n1846 0.235885
R3199 VDD.n2235 VDD.n2232 0.235837
R3200 VDD.n2451 VDD.n2448 0.235837
R3201 VDD.n2220 VDD.n2217 0.23543
R3202 VDD.n2436 VDD.n2433 0.23543
R3203 VDD.n1894 VDD.n1892 0.235355
R3204 VDD.n2223 VDD.n2220 0.235271
R3205 VDD.n2439 VDD.n2436 0.235271
R3206 VDD.n2211 VDD.n2208 0.234863
R3207 VDD.n2427 VDD.n2424 0.234863
R3208 VDD.n2217 VDD.n2214 0.234297
R3209 VDD.n2214 VDD.n2211 0.234297
R3210 VDD.n2433 VDD.n2430 0.234297
R3211 VDD.n2430 VDD.n2427 0.234297
R3212 VDD.n2205 VDD.n2202 0.234293
R3213 VDD.n2421 VDD.n2418 0.234293
R3214 VDD.n2238 VDD.n2235 0.234291
R3215 VDD.n2454 VDD.n2451 0.234291
R3216 VDD.n2226 VDD.n2223 0.233514
R3217 VDD.n2442 VDD.n2439 0.233514
R3218 VDD.n2232 VDD.n2229 0.233447
R3219 VDD.n2448 VDD.n2445 0.233447
R3220 VDD.n2208 VDD.n2205 0.233445
R3221 VDD.n2424 VDD.n2421 0.233445
R3222 VDD.n609 VDD.n608 0.233429
R3223 VDD.n2229 VDD.n2226 0.233389
R3224 VDD.n2445 VDD.n2442 0.233389
R3225 VDD.n442 VDD.n408 0.229786
R3226 VDD.n697 VDD.n694 0.229786
R3227 VDD.n751 VDD.n750 0.229786
R3228 VDD.n1366 VDD.n361 0.229786
R3229 VDD.n2005 VDD.n1986 0.228829
R3230 VDD.n2279 VDD.n2276 0.226747
R3231 VDD.n2495 VDD.n2492 0.226747
R3232 VDD.n2267 VDD.n2264 0.225529
R3233 VDD.n2483 VDD.n2480 0.225529
R3234 VDD.n2258 VDD.n2255 0.225387
R3235 VDD.n2474 VDD.n2471 0.225387
R3236 VDD.n2273 VDD.n2270 0.225121
R3237 VDD.n2489 VDD.n2486 0.225121
R3238 VDD.n2255 VDD.n2252 0.225121
R3239 VDD.n2471 VDD.n2468 0.225121
R3240 VDD.n2264 VDD.n2261 0.22512
R3241 VDD.n2480 VDD.n2477 0.22512
R3242 VDD.n2249 VDD.n2246 0.22512
R3243 VDD.n2465 VDD.n2462 0.22512
R3244 VDD.n2252 VDD.n2249 0.224578
R3245 VDD.n2468 VDD.n2465 0.224578
R3246 VDD.n2246 VDD.n2243 0.223901
R3247 VDD.n2462 VDD.n2459 0.223901
R3248 VDD.n2270 VDD.n2267 0.22363
R3249 VDD.n2486 VDD.n2483 0.22363
R3250 VDD.n2276 VDD.n2273 0.222816
R3251 VDD.n2492 VDD.n2489 0.222816
R3252 VDD.n2261 VDD.n2258 0.22281
R3253 VDD.n2477 VDD.n2474 0.22281
R3254 VDD.n1260 VDD.n1259 0.221442
R3255 VDD.n1464 VDD.n1461 0.220495
R3256 VDD VDD.n2682 0.218882
R3257 VDD.n883 VDD.n831 0.217222
R3258 VDD VDD.n1921 0.215115
R3259 VDD.n1916 VDD 0.215115
R3260 VDD.n153 VDD 0.215115
R3261 VDD.n93 VDD 0.215115
R3262 VDD.n2105 VDD 0.215115
R3263 VDD.n2640 VDD 0.215115
R3264 VDD.n1029 VDD.n1028 0.209826
R3265 VDD.n1713 VDD.n1647 0.209826
R3266 VDD.n2289 VDD.n2287 0.20611
R3267 VDD.n2505 VDD.n2503 0.20611
R3268 VDD.n1920 VDD.n1818 0.194429
R3269 VDD.n1941 VDD.n1940 0.193912
R3270 VDD.n1923 VDD.n1819 0.192121
R3271 VDD.n2162 VDD.n2160 0.189731
R3272 VDD.n2141 VDD.n2137 0.189731
R3273 VDD.n2132 VDD.n2131 0.189731
R3274 VDD.n2096 VDD.n2082 0.189731
R3275 VDD.n2015 VDD.n2014 0.189249
R3276 VDD.n148 VDD.n34 0.188457
R3277 VDD.n2295 VDD.n2293 0.186866
R3278 VDD.n2514 VDD.n2512 0.186802
R3279 VDD.n1927 VDD.n1926 0.186352
R3280 VDD.n2344 VDD.n2342 0.185622
R3281 VDD.n2587 VDD.n2585 0.185622
R3282 VDD.n1673 VDD.n1672 0.183919
R3283 VDD.n1928 VDD.n1821 0.182274
R3284 VDD.n145 VDD.n111 0.182274
R3285 VDD.n48 VDD.n47 0.182274
R3286 VDD.n856 VDD.n850 0.182274
R3287 VDD.n2607 VDD.n2606 0.182274
R3288 VDD.n167 VDD.n166 0.18216
R3289 VDD.n1908 VDD.n1883 0.182033
R3290 VDD.n1413 VDD.n1411 0.182033
R3291 VDD.n440 VDD.n439 0.182033
R3292 VDD.n461 VDD.n393 0.182033
R3293 VDD.n1348 VDD.n1347 0.182033
R3294 VDD.n1369 VDD.n1368 0.182033
R3295 VDD.n2080 VDD.n2079 0.182033
R3296 VDD.n152 VDD.n151 0.179788
R3297 VDD.n2340 VDD.n2339 0.179768
R3298 VDD.n2335 VDD.n2334 0.179768
R3299 VDD.n2583 VDD.n2582 0.179768
R3300 VDD.n2578 VDD.n2577 0.179768
R3301 VDD.n2332 VDD.n2331 0.179037
R3302 VDD.n2575 VDD.n2574 0.179037
R3303 VDD.n1526 VDD.n315 0.178585
R3304 VDD.n153 VDD.n20 0.177873
R3305 VDD.n1252 VDD.n1248 0.17667
R3306 VDD.n1517 VDD.n279 0.176655
R3307 VDD.n1291 VDD.n476 0.176655
R3308 VDD.n91 VDD.n36 0.175635
R3309 VDD.n1960 VDD.n1959 0.175419
R3310 VDD.n1841 VDD 0.174184
R3311 VDD VDD.n1840 0.174184
R3312 VDD.n1801 VDD.n1792 0.174184
R3313 VDD.n1871 VDD 0.174184
R3314 VDD VDD.n1870 0.174184
R3315 VDD.n1856 VDD.n1847 0.174184
R3316 VDD.n164 VDD 0.174184
R3317 VDD VDD.n163 0.174184
R3318 VDD.n30 VDD.n21 0.174184
R3319 VDD.n104 VDD 0.174184
R3320 VDD VDD.n103 0.174184
R3321 VDD.n87 VDD.n78 0.174184
R3322 VDD.n2093 VDD 0.174184
R3323 VDD VDD.n2092 0.174184
R3324 VDD.n2117 VDD.n2115 0.174184
R3325 VDD.n2603 VDD 0.174184
R3326 VDD VDD.n2602 0.174184
R3327 VDD.n2661 VDD.n2659 0.174184
R3328 VDD.n466 VDD.n462 0.174122
R3329 VDD VDD.n1800 0.173395
R3330 VDD VDD.n1855 0.173395
R3331 VDD VDD.n29 0.173395
R3332 VDD VDD.n86 0.173395
R3333 VDD.n2112 VDD 0.173395
R3334 VDD.n2656 VDD 0.173395
R3335 VDD.n2329 VDD.n2328 0.172451
R3336 VDD.n2572 VDD.n2571 0.172451
R3337 VDD.n1277 VDD.n1192 0.17241
R3338 VDD.n1575 VDD.n273 0.17241
R3339 VDD.n2337 VDD.n2336 0.17172
R3340 VDD.n2580 VDD.n2579 0.17172
R3341 VDD.n1569 VDD.n1568 0.171399
R3342 VDD.n1185 VDD.n483 0.171399
R3343 VDD.n107 VDD.n106 0.169275
R3344 VDD.n92 VDD.n37 0.166766
R3345 VDD.n1963 VDD.n1962 0.165258
R3346 VDD.n93 VDD.n38 0.16483
R3347 VDD.n1541 VDD.n1540 0.163357
R3348 VDD.n1237 VDD.n1236 0.163357
R3349 VDD.n1842 VDD.n1841 0.158395
R3350 VDD.n1804 VDD.n1792 0.158395
R3351 VDD.n1872 VDD.n1871 0.158395
R3352 VDD.n1859 VDD.n1847 0.158395
R3353 VDD.n165 VDD.n164 0.158395
R3354 VDD.n33 VDD.n21 0.158395
R3355 VDD.n105 VDD.n104 0.158395
R3356 VDD.n90 VDD.n78 0.158395
R3357 VDD.n2094 VDD.n2093 0.158395
R3358 VDD.n2118 VDD.n2117 0.158395
R3359 VDD.n2604 VDD.n2603 0.158395
R3360 VDD.n2662 VDD.n2661 0.158395
R3361 VDD.n1569 VDD.n268 0.157434
R3362 VDD.n1186 VDD.n1185 0.15672
R3363 VDD.n1030 VDD.n552 0.153197
R3364 VDD.n1715 VDD.n1714 0.153197
R3365 VDD.n1667 VDD.n1639 0.146319
R3366 VDD.n1536 VDD.n1535 0.146214
R3367 VDD.n1242 VDD.n1241 0.146214
R3368 VDD.n1030 VDD.n1029 0.146118
R3369 VDD.n1714 VDD.n1713 0.146118
R3370 VDD.n1036 VDD.n558 0.146022
R3371 VDD.n829 VDD.n827 0.143441
R3372 VDD.n1286 VDD.n482 0.143084
R3373 VDD.n1537 VDD.n311 0.143
R3374 VDD.n1277 VDD.n1276 0.142944
R3375 VDD.n313 VDD.n273 0.142944
R3376 VDD.n2287 VDD.n2286 0.142451
R3377 VDD.n2503 VDD.n2502 0.142451
R3378 VDD.n1253 VDD.n1252 0.142202
R3379 VDD.n317 VDD.n315 0.142202
R3380 VDD.n1566 VDD.n1565 0.142073
R3381 VDD.n1240 VDD.n1197 0.141929
R3382 VDD.n1565 VDD.n279 0.141062
R3383 VDD.n482 VDD.n476 0.141062
R3384 VDD.n1553 VDD.n1550 0.140857
R3385 VDD.n1227 VDD.n1210 0.140857
R3386 VDD.n2677 VDD.n2181 0.140627
R3387 VDD.n1028 VDD.n561 0.14038
R3388 VDD.n1688 VDD.n1647 0.14038
R3389 VDD.n1554 VDD.n1553 0.139786
R3390 VDD.n1535 VDD.n1532 0.139786
R3391 VDD.n1242 VDD.n1193 0.139786
R3392 VDD.n1222 VDD.n1210 0.139786
R3393 VDD VDD.n688 0.139763
R3394 VDD.n1341 VDD.n1340 0.139295
R3395 VDD.n1974 VDD.n1973 0.1385
R3396 VDD.n1340 VDD.n377 0.138211
R3397 VDD.n1473 VDD.n1471 0.138211
R3398 VDD.n1549 VDD.n1548 0.137643
R3399 VDD.n1229 VDD.n1228 0.137643
R3400 VDD.n1576 VDD.n1575 0.137017
R3401 VDD.n1192 VDD.n1191 0.136006
R3402 VDD.n1800 VDD.n1798 0.1355
R3403 VDD.n1855 VDD.n1853 0.1355
R3404 VDD.n29 VDD.n27 0.1355
R3405 VDD.n86 VDD.n84 0.1355
R3406 VDD.n2112 VDD.n2111 0.1355
R3407 VDD.n2132 VDD.n2119 0.1355
R3408 VDD.n2137 VDD.n2105 0.1355
R3409 VDD.n2162 VDD.n2104 0.1355
R3410 VDD.n2096 VDD.n2095 0.1355
R3411 VDD.n2656 VDD.n2655 0.1355
R3412 VDD.n2670 VDD.n2612 0.1355
R3413 VDD.n1840 VDD.n1839 0.134711
R3414 VDD.n1870 VDD.n1869 0.134711
R3415 VDD.n163 VDD.n162 0.134711
R3416 VDD.n103 VDD.n102 0.134711
R3417 VDD.n2092 VDD.n2091 0.134711
R3418 VDD.n2602 VDD.n2601 0.134711
R3419 VDD.n1499 VDD.n331 0.133873
R3420 VDD.n1493 VDD.n1492 0.133873
R3421 VDD.n1490 VDD.n1488 0.133873
R3422 VDD.n1486 VDD.n1484 0.133873
R3423 VDD.n1482 VDD.n1480 0.133873
R3424 VDD.n1478 VDD.n1476 0.133873
R3425 VDD.n1334 VDD.n377 0.133873
R3426 VDD.n1333 VDD.n1331 0.133873
R3427 VDD.n1329 VDD.n1327 0.133873
R3428 VDD.n1325 VDD.n1323 0.133873
R3429 VDD.n1321 VDD.n1319 0.133873
R3430 VDD.n1317 VDD.n1315 0.133873
R3431 VDD.n1313 VDD.n1311 0.133873
R3432 VDD.n1504 VDD.n1503 0.133833
R3433 VDD.n329 VDD.n327 0.133833
R3434 VDD.n1514 VDD.n327 0.133833
R3435 VDD.n1517 VDD.n1516 0.133833
R3436 VDD.n1292 VDD.n1291 0.133833
R3437 VDD.n1298 VDD.n1297 0.133833
R3438 VDD.n1297 VDD.n1296 0.133833
R3439 VDD.n1307 VDD.n469 0.133833
R3440 VDD.n2589 VDD.n2588 0.133683
R3441 VDD.n1563 VDD.n278 0.133132
R3442 VDD.n724 VDD 0.131587
R3443 VDD.n1270 VDD.n1253 0.131498
R3444 VDD.n318 VDD.n317 0.13055
R3445 VDD.n1961 VDD.n1960 0.130419
R3446 VDD.n1229 VDD.n1207 0.130143
R3447 VDD.n723 VDD 0.12963
R3448 VDD.n1023 VDD.n561 0.129536
R3449 VDD.n1023 VDD.n1022 0.129536
R3450 VDD.n1020 VDD.n567 0.129536
R3451 VDD.n1015 VDD.n567 0.129536
R3452 VDD.n1015 VDD.n1014 0.129536
R3453 VDD.n1012 VDD.n571 0.129536
R3454 VDD.n1007 VDD.n571 0.129536
R3455 VDD.n1005 VDD.n1004 0.129536
R3456 VDD.n1004 VDD.n575 0.129536
R3457 VDD.n999 VDD.n575 0.129536
R3458 VDD.n997 VDD.n996 0.129536
R3459 VDD.n1671 VDD.n1670 0.129536
R3460 VDD.n1665 VDD.n1663 0.129536
R3461 VDD.n1679 VDD.n1663 0.129536
R3462 VDD.n1680 VDD.n1679 0.129536
R3463 VDD.n1682 VDD.n1654 0.129536
R3464 VDD.n1705 VDD.n1654 0.129536
R3465 VDD.n1703 VDD.n1702 0.129536
R3466 VDD.n1702 VDD.n1656 0.129536
R3467 VDD.n1695 VDD.n1656 0.129536
R3468 VDD.n1693 VDD.n1692 0.129536
R3469 VDD.n1692 VDD.n1688 0.129536
R3470 VDD.n874 VDD.n837 0.129141
R3471 VDD.n1548 VDD.n305 0.129071
R3472 VDD.n2612 VDD.n2611 0.128577
R3473 VDD.n1253 VDD.n1251 0.128395
R3474 VDD.n317 VDD.n316 0.128395
R3475 VDD.n2338 VDD.n2337 0.127817
R3476 VDD.n2581 VDD.n2580 0.127817
R3477 VDD.n1492 VDD.n1490 0.127367
R3478 VDD.n1488 VDD.n1486 0.127367
R3479 VDD.n1484 VDD.n1482 0.127367
R3480 VDD.n1480 VDD.n1478 0.127367
R3481 VDD.n998 VDD.n997 0.127367
R3482 VDD.n1334 VDD.n1333 0.127367
R3483 VDD.n1331 VDD.n1329 0.127367
R3484 VDD.n1327 VDD.n1325 0.127367
R3485 VDD.n1323 VDD.n1321 0.127367
R3486 VDD.n1319 VDD.n1317 0.127367
R3487 VDD.n1670 VDD.n1669 0.127367
R3488 VDD.n2330 VDD.n2329 0.126354
R3489 VDD.n2573 VDD.n2572 0.126354
R3490 VDD.n2673 VDD.n2672 0.12616
R3491 VDD.n826 VDD.n749 0.126143
R3492 VDD.n1493 VDD.n331 0.124114
R3493 VDD.n1315 VDD.n1313 0.124114
R3494 VDD.n1269 VDD.n1268 0.123227
R3495 VDD.n1268 VDD.n1254 0.123227
R3496 VDD.n1262 VDD.n1261 0.123227
R3497 VDD.n1261 VDD.n376 0.123227
R3498 VDD.n1460 VDD.n1456 0.123227
R3499 VDD.n1465 VDD.n1460 0.123227
R3500 VDD.n1463 VDD.n1462 0.123227
R3501 VDD.n1462 VDD.n320 0.123227
R3502 VDD.n1013 VDD.n1012 0.12303
R3503 VDD.n1705 VDD.n1704 0.12303
R3504 VDD.n1260 VDD.n1254 0.122205
R3505 VDD.n1464 VDD.n1463 0.122205
R3506 VDD.n1043 VDD.n552 0.120837
R3507 VDD.n1044 VDD.n1043 0.120837
R3508 VDD.n1045 VDD.n1044 0.120837
R3509 VDD.n1045 VDD.n538 0.120837
R3510 VDD.n1060 VDD.n539 0.120837
R3511 VDD.n539 VDD.n530 0.120837
R3512 VDD.n1125 VDD.n530 0.120837
R3513 VDD.n1128 VDD.n1127 0.120837
R3514 VDD.n1128 VDD.n519 0.120837
R3515 VDD.n1141 VDD.n519 0.120837
R3516 VDD.n1142 VDD.n1141 0.120837
R3517 VDD.n1144 VDD.n1142 0.120837
R3518 VDD.n1144 VDD.n1143 0.120837
R3519 VDD.n1159 VDD.n1158 0.120837
R3520 VDD.n1161 VDD.n1159 0.120837
R3521 VDD.n1161 VDD.n1160 0.120837
R3522 VDD.n1176 VDD.n1175 0.120837
R3523 VDD.n1177 VDD.n1176 0.120837
R3524 VDD.n1177 VDD.n490 0.120837
R3525 VDD.n1191 VDD.n490 0.120837
R3526 VDD.n1577 VDD.n1576 0.120837
R3527 VDD.n1577 VDD.n264 0.120837
R3528 VDD.n1589 VDD.n264 0.120837
R3529 VDD.n1590 VDD.n1589 0.120837
R3530 VDD.n1603 VDD.n1602 0.120837
R3531 VDD.n1602 VDD.n1601 0.120837
R3532 VDD.n1601 VDD.n1592 0.120837
R3533 VDD.n1759 VDD.n1758 0.120837
R3534 VDD.n1758 VDD.n1757 0.120837
R3535 VDD.n1757 VDD.n180 0.120837
R3536 VDD.n195 VDD.n180 0.120837
R3537 VDD.n1745 VDD.n195 0.120837
R3538 VDD.n1745 VDD.n1744 0.120837
R3539 VDD.n1742 VDD.n199 0.120837
R3540 VDD.n215 VDD.n199 0.120837
R3541 VDD.n1730 VDD.n215 0.120837
R3542 VDD.n1728 VDD.n1727 0.120837
R3543 VDD.n1727 VDD.n1630 0.120837
R3544 VDD.n1646 VDD.n1630 0.120837
R3545 VDD.n1715 VDD.n1646 0.120837
R3546 VDD.n2348 VDD.n2347 0.119146
R3547 VDD.n1308 VDD.n467 0.119037
R3548 VDD.n292 VDD.n277 0.117286
R3549 VDD.n1545 VDD.n1544 0.117286
R3550 VDD.n1532 VDD.n1531 0.117286
R3551 VDD.n1247 VDD.n1193 0.117286
R3552 VDD.n1233 VDD.n1232 0.117286
R3553 VDD.n1284 VDD.n484 0.117286
R3554 VDD.n1783 VDD.n1782 0.115972
R3555 VDD.n16 VDD.n15 0.115972
R3556 VDD.n2180 VDD.n2179 0.115087
R3557 VDD.n1958 VDD.n1956 0.113142
R3558 VDD.n1271 VDD.n1270 0.113
R3559 VDD.n2334 VDD.n2333 0.112451
R3560 VDD.n2577 VDD.n2576 0.112451
R3561 VDD.n1525 VDD.n318 0.111977
R3562 VDD.n2342 VDD.n2341 0.11172
R3563 VDD.n2585 VDD.n2584 0.11172
R3564 VDD.n1061 VDD.n1060 0.110725
R3565 VDD.n15 VDD.n7 0.109745
R3566 VDD.n1730 VDD.n1729 0.109713
R3567 VDD.n1567 VDD.n277 0.108714
R3568 VDD.n2668 VDD.n2667 0.108385
R3569 VDD.n2678 VDD.n2677 0.108044
R3570 VDD.n1221 VDD.n1220 0.107643
R3571 VDD.n1285 VDD.n1284 0.107643
R3572 VDD.n881 VDD.n880 0.106797
R3573 VDD.n1556 VDD.n1555 0.106571
R3574 VDD.n1603 VDD.n1591 0.103646
R3575 VDD.n1160 VDD.n499 0.102635
R3576 VDD.n1766 VDD.n1765 0.101533
R3577 VDD.n985 VDD.n584 0.101088
R3578 VDD.n1037 VDD.n1036 0.1005
R3579 VDD.n1720 VDD.n1639 0.1005
R3580 VDD.n1788 VDD.n1787 0.0989906
R3581 VDD.n2666 VDD.n2665 0.0985769
R3582 VDD.n1516 VDD.n1515 0.0971667
R3583 VDD.n1293 VDD.n1292 0.0971667
R3584 VDD.n1779 VDD.n17 0.0964434
R3585 VDD.n168 VDD.n18 0.0960507
R3586 VDD.n1944 VDD.n1789 0.0960507
R3587 VDD.n150 VDD.n18 0.0952577
R3588 VDD.n1789 VDD.n1774 0.0952577
R3589 VDD.n293 VDD.n292 0.0947857
R3590 VDD.n1219 VDD.n484 0.0947857
R3591 VDD.n1286 VDD.n1285 0.0945449
R3592 VDD.n1504 VDD.n1500 0.0938198
R3593 VDD.n1308 VDD.n1307 0.0938198
R3594 VDD.n1567 VDD.n1566 0.0935337
R3595 VDD.n2290 VDD.n2289 0.0934268
R3596 VDD.n2506 VDD.n2505 0.0934268
R3597 VDD.n2042 VDD.n2041 0.0914091
R3598 VDD.n2041 VDD.n2040 0.0914091
R3599 VDD.n2040 VDD.n2039 0.0914091
R3600 VDD.n2039 VDD.n2038 0.0914091
R3601 VDD.n2038 VDD.n2037 0.0914091
R3602 VDD.n2037 VDD.n2036 0.0914091
R3603 VDD.n2035 VDD.n2026 0.0914091
R3604 VDD.n2070 VDD.n2068 0.0914091
R3605 VDD.n2072 VDD.n2070 0.0914091
R3606 VDD.n150 VDD.n149 0.0905
R3607 VDD.n1774 VDD.n1773 0.0905
R3608 VDD VDD.n2035 0.0900455
R3609 VDD.n1839 VDD.n1838 0.0893158
R3610 VDD.n1798 VDD.n1797 0.0893158
R3611 VDD.n1869 VDD.n1868 0.0893158
R3612 VDD.n1853 VDD.n1852 0.0893158
R3613 VDD.n162 VDD.n161 0.0893158
R3614 VDD.n27 VDD.n26 0.0893158
R3615 VDD.n102 VDD.n101 0.0893158
R3616 VDD.n84 VDD.n83 0.0893158
R3617 VDD.n678 VDD.n677 0.0893158
R3618 VDD.n895 VDD.n889 0.0893158
R3619 VDD.n895 VDD.n894 0.0893158
R3620 VDD.n2091 VDD.n2090 0.0893158
R3621 VDD.n2111 VDD.n2110 0.0893158
R3622 VDD.n2601 VDD.n2600 0.0893158
R3623 VDD.n2655 VDD.n2654 0.0893158
R3624 VDD.n1275 VDD.n1248 0.0884545
R3625 VDD.n967 VDD.n941 0.088
R3626 VDD.n1158 VDD.n509 0.0874663
R3627 VDD.n1527 VDD.n1526 0.0874318
R3628 VDD.n2179 VDD.n2176 0.0865195
R3629 VDD.n1592 VDD.n179 0.0864551
R3630 VDD.n1502 VDD.n329 0.0860556
R3631 VDD.n1296 VDD.n1295 0.0860556
R3632 VDD.n1582 VDD.n268 0.0855
R3633 VDD.n1583 VDD.n1582 0.0855
R3634 VDD.n1584 VDD.n1583 0.0855
R3635 VDD.n1584 VDD.n238 0.0855
R3636 VDD.n1608 VDD.n239 0.0855
R3637 VDD.n1595 VDD.n239 0.0855
R3638 VDD.n1595 VDD.n171 0.0855
R3639 VDD.n1038 VDD.n1037 0.0855
R3640 VDD.n1038 VDD.n549 0.0855
R3641 VDD.n1051 VDD.n549 0.0855
R3642 VDD.n1052 VDD.n1051 0.0855
R3643 VDD.n1055 VDD.n1054 0.0855
R3644 VDD.n1054 VDD.n535 0.0855
R3645 VDD.n1120 VDD.n535 0.0855
R3646 VDD.n1134 VDD.n524 0.0855
R3647 VDD.n1135 VDD.n1134 0.0855
R3648 VDD.n1136 VDD.n515 0.0855
R3649 VDD.n1150 VDD.n515 0.0855
R3650 VDD.n1151 VDD.n1150 0.0855
R3651 VDD.n1153 VDD.n505 0.0855
R3652 VDD.n1167 VDD.n505 0.0855
R3653 VDD.n1168 VDD.n1167 0.0855
R3654 VDD.n1170 VDD.n495 0.0855
R3655 VDD.n1183 VDD.n495 0.0855
R3656 VDD.n1184 VDD.n1183 0.0855
R3657 VDD.n1186 VDD.n1184 0.0855
R3658 VDD.n188 VDD.n172 0.0855
R3659 VDD.n1752 VDD.n188 0.0855
R3660 VDD.n1751 VDD.n1750 0.0855
R3661 VDD.n1750 VDD.n189 0.0855
R3662 VDD.n1737 VDD.n207 0.0855
R3663 VDD.n1737 VDD.n1736 0.0855
R3664 VDD.n1736 VDD.n1735 0.0855
R3665 VDD.n1638 VDD.n1637 0.0855
R3666 VDD.n1722 VDD.n1638 0.0855
R3667 VDD.n1722 VDD.n1721 0.0855
R3668 VDD.n1721 VDD.n1720 0.0855
R3669 VDD.n2009 VDD.n2008 0.0853962
R3670 VDD.n1022 VDD.n1021 0.0850783
R3671 VDD.n1694 VDD.n1693 0.0850783
R3672 VDD.n1055 VDD.n1053 0.0847857
R3673 VDD.n1735 VDD.n208 0.0840714
R3674 VDD.n681 VDD 0.0836933
R3675 VDD.n1476 VDD.n1474 0.0818253
R3676 VDD.n2008 VDD.n2007 0.0817389
R3677 VDD.n2007 VDD.n2006 0.0817389
R3678 VDD.n1787 VDD 0.0811604
R3679 VDD.n1743 VDD.n1742 0.0803876
R3680 VDD VDD.n1970 0.0798636
R3681 VDD.n1126 VDD.n1125 0.0793764
R3682 VDD.n905 VDD.n745 0.0790106
R3683 VDD.n1972 VDD 0.0778182
R3684 VDD.n896 VDD 0.0774922
R3685 VDD.n1568 VDD.n1567 0.0773539
R3686 VDD.n1285 VDD.n483 0.0773539
R3687 VDD.n1541 VDD.n307 0.0765714
R3688 VDD.n1236 VDD.n1200 0.0765714
R3689 VDD.n1506 VDD.n1505 0.0752312
R3690 VDD.n109 VDD.n108 0.0751875
R3691 VDD.n1306 VDD.n468 0.074985
R3692 VDD.n1007 VDD.n1006 0.0742349
R3693 VDD.n1682 VDD.n1681 0.0742349
R3694 VDD.n829 VDD.n828 0.07388
R3695 VDD.n1474 VDD.n1473 0.0731506
R3696 VDD.n701 VDD.n670 0.0717174
R3697 VDD.n700 VDD.n699 0.0717174
R3698 VDD.n1933 VDD.n1932 0.0714756
R3699 VDD.n1830 VDD.n1829 0.0714756
R3700 VDD.n1902 VDD.n1874 0.0714756
R3701 VDD.n1911 VDD.n1881 0.0714756
R3702 VDD.n146 VDD.n121 0.0714756
R3703 VDD.n139 VDD.n125 0.0714756
R3704 VDD.n61 VDD.n50 0.0714756
R3705 VDD.n68 VDD.n45 0.0714756
R3706 VDD.n1425 VDD.n1398 0.0714756
R3707 VDD.n1434 VDD.n1389 0.0714756
R3708 VDD.n430 VDD.n421 0.0714756
R3709 VDD.n449 VDD.n448 0.0714756
R3710 VDD.n870 VDD.n869 0.0714756
R3711 VDD.n952 VDD.n949 0.0714756
R3712 VDD.n1359 VDD.n363 0.0714756
R3713 VDD.n1380 VDD.n1379 0.0714756
R3714 VDD.n1442 VDD.n345 0.0714756
R3715 VDD.n2149 VDD.n2146 0.0714756
R3716 VDD.n2634 VDD.n2633 0.0714756
R3717 VDD.n907 VDD.n906 0.0714615
R3718 VDD.n110 VDD.n109 0.0714375
R3719 VDD.n1424 VDD 0.0713871
R3720 VDD VDD.n431 0.0713871
R3721 VDD.n450 VDD 0.0713871
R3722 VDD VDD.n839 0.0713871
R3723 VDD VDD.n960 0.0713871
R3724 VDD.n1358 VDD 0.0713871
R3725 VDD.n1422 VDD.n1408 0.0709032
R3726 VDD.n1416 VDD.n1415 0.0709032
R3727 VDD.n411 VDD.n409 0.0709032
R3728 VDD.n433 VDD.n414 0.0709032
R3729 VDD.n458 VDD.n392 0.0709032
R3730 VDD.n457 VDD.n456 0.0709032
R3731 VDD.n854 VDD.n848 0.0709032
R3732 VDD.n861 VDD.n860 0.0709032
R3733 VDD.n1350 VDD.n1349 0.0709032
R3734 VDD.n1352 VDD.n1351 0.0709032
R3735 VDD.n358 VDD.n355 0.0709032
R3736 VDD.n962 VDD.n940 0.0701774
R3737 VDD.n1813 VDD.n1806 0.0692805
R3738 VDD.n1939 VDD.n1807 0.0692805
R3739 VDD VDD.n1933 0.0692805
R3740 VDD.n1895 VDD.n1891 0.0692805
R3741 VDD.n1893 VDD.n1886 0.0692805
R3742 VDD.n1902 VDD 0.0692805
R3743 VDD.n139 VDD 0.0692805
R3744 VDD.n137 VDD.n126 0.0692805
R3745 VDD.n131 VDD.n130 0.0692805
R3746 VDD VDD.n68 0.0692805
R3747 VDD.n70 VDD.n39 0.0692805
R3748 VDD.n76 VDD.n41 0.0692805
R3749 VDD.n1430 VDD.n1398 0.0692805
R3750 VDD.n1425 VDD.n1424 0.0692805
R3751 VDD.n1434 VDD.n1433 0.0692805
R3752 VDD.n1440 VDD.n1389 0.0692805
R3753 VDD.n431 VDD.n430 0.0692805
R3754 VDD.n425 VDD.n421 0.0692805
R3755 VDD.n450 VDD.n449 0.0692805
R3756 VDD.n448 VDD.n444 0.0692805
R3757 VDD.n869 VDD.n839 0.0692805
R3758 VDD.n960 VDD.n949 0.0692805
R3759 VDD.n954 VDD.n952 0.0692805
R3760 VDD.n1359 VDD.n1358 0.0692805
R3761 VDD.n1364 VDD.n363 0.0692805
R3762 VDD.n1380 VDD.n349 0.0692805
R3763 VDD.n1379 VDD.n1378 0.0692805
R3764 VDD.n1442 VDD 0.0692805
R3765 VDD.n2127 VDD.n2124 0.0692805
R3766 VDD.n2146 VDD 0.0692805
R3767 VDD.n2648 VDD.n2645 0.0692805
R3768 VDD.n2630 VDD.n2627 0.0692805
R3769 VDD VDD.n2634 0.0692805
R3770 VDD.n2175 VDD.n2172 0.0692083
R3771 VDD.n1416 VDD.n1408 0.0687258
R3772 VDD.n1415 VDD.n1414 0.0687258
R3773 VDD.n441 VDD.n409 0.0687258
R3774 VDD.n414 VDD.n411 0.0687258
R3775 VDD.n462 VDD.n392 0.0687258
R3776 VDD.n458 VDD.n457 0.0687258
R3777 VDD.n855 VDD.n854 0.0687258
R3778 VDD.n860 VDD.n848 0.0687258
R3779 VDD.n1352 VDD.n1350 0.0687258
R3780 VDD.n1367 VDD.n358 0.0687258
R3781 VDD.n2671 VDD.n2670 0.0685545
R3782 VDD.n1153 VDD.n1152 0.0683571
R3783 VDD.n2065 VDD.n2063 0.0682273
R3784 VDD.n2341 VDD.n2340 0.0678171
R3785 VDD.n2333 VDD.n2332 0.0678171
R3786 VDD.n2584 VDD.n2583 0.0678171
R3787 VDD.n2576 VDD.n2575 0.0678171
R3788 VDD.n2015 VDD.n2009 0.0676691
R3789 VDD.n2676 VDD.n2182 0.0669557
R3790 VDD.n729 VDD.n624 0.0669486
R3791 VDD.n728 VDD.n727 0.0669486
R3792 VDD.n1287 VDD.n480 0.0668158
R3793 VDD.n1609 VDD.n1608 0.0662143
R3794 VDD.n1169 VDD.n1168 0.0662143
R3795 VDD.n740 VDD.n739 0.0661075
R3796 VDD.n741 VDD.n586 0.0661075
R3797 VDD.n681 VDD.n678 0.0647857
R3798 VDD.n911 VDD.n910 0.0646489
R3799 VDD.n2006 VDD.n2005 0.0643765
R3800 VDD.n2664 VDD.n2649 0.0639615
R3801 VDD.n2666 VDD.n2639 0.0639615
R3802 VDD.n2668 VDD.n2623 0.0639615
R3803 VDD.n2610 VDD.n2609 0.0639615
R3804 VDD.n1423 VDD.n1422 0.0629194
R3805 VDD.n433 VDD.n432 0.0629194
R3806 VDD.n456 VDD.n401 0.0629194
R3807 VDD.n862 VDD.n861 0.0629194
R3808 VDD.n962 VDD.n961 0.0629194
R3809 VDD.n1351 VDD.n372 0.0629194
R3810 VDD.n1922 VDD 0.0616538
R3811 VDD VDD.n1915 0.0616538
R3812 VDD VDD.n152 0.0616538
R3813 VDD VDD.n92 0.0616538
R3814 VDD VDD.n2104 0.0616538
R3815 VDD VDD.n2624 0.0616538
R3816 VDD.n896 VDD.n895 0.0606172
R3817 VDD.n871 VDD.n870 0.0605
R3818 VDD.n1388 VDD.n349 0.0605
R3819 VDD.n2178 VDD.n2177 0.0593952
R3820 VDD.n2283 VDD.n2280 0.0587571
R3821 VDD.n2499 VDD.n2496 0.0587571
R3822 VDD.n912 VDD.n744 0.0584808
R3823 VDD VDD.n6 0.0582358
R3824 VDD.n1818 VDD.n1807 0.0561098
R3825 VDD.n1886 VDD.n1846 0.0561098
R3826 VDD.n138 VDD.n137 0.0561098
R3827 VDD.n70 VDD.n69 0.0561098
R3828 VDD.n2141 VDD.n2140 0.0561098
R3829 VDD.n2639 VDD.n2630 0.0561098
R3830 VDD.n1006 VDD.n1005 0.0558012
R3831 VDD.n1681 VDD.n1680 0.0558012
R3832 VDD.n1927 VDD.n1830 0.055378
R3833 VDD.n1907 VDD.n1881 0.055378
R3834 VDD.n147 VDD.n146 0.055378
R3835 VDD.n50 VDD.n49 0.055378
R3836 VDD VDD.n1441 0.055378
R3837 VDD.n2082 VDD.n2081 0.055378
R3838 VDD.n2609 VDD.n2608 0.055378
R3839 VDD.n2068 VDD.n2066 0.0550455
R3840 VDD.n2003 VDD.n1986 0.0549355
R3841 VDD.n2331 VDD.n2330 0.0539146
R3842 VDD.n2574 VDD.n2573 0.0539146
R3843 VDD.n938 VDD.n937 0.0534412
R3844 VDD.n935 VDD.n916 0.0534412
R3845 VDD.n1114 VDD.n537 0.0533261
R3846 VDD.n1618 VDD.n1617 0.0533261
R3847 VDD.n2004 VDD.n2003 0.0530664
R3848 VDD.n1276 VDD.n1247 0.053
R3849 VDD.n1454 VDD.n345 0.0524512
R3850 VDD.n2339 VDD.n2338 0.0524512
R3851 VDD.n2582 VDD.n2581 0.0524512
R3852 VDD.n6 VDD.n5 0.0522925
R3853 VDD.n1531 VDD.n313 0.0519286
R3854 VDD.n2076 VDD.n2072 0.0514091
R3855 VDD.n672 VDD.n671 0.0509
R3856 VDD.n903 VDD.n746 0.0504219
R3857 VDD.n1388 VDD.n355 0.0498548
R3858 VDD.n1120 VDD.n1119 0.0497857
R3859 VDD.n220 VDD.n207 0.0497857
R3860 VDD.n1924 VDD.n1790 0.0495909
R3861 VDD.n1752 VDD 0.0483571
R3862 VDD.n1503 VDD.n1502 0.0482778
R3863 VDD.n1295 VDD.n469 0.0482778
R3864 VDD.n1943 VDD.n1790 0.0472532
R3865 VDD.n1918 VDD.n1791 0.0472532
R3866 VDD.n1845 VDD.n1844 0.046898
R3867 VDD.n2136 VDD.n2132 0.0468823
R3868 VDD.n1136 VDD 0.0462143
R3869 VDD.n690 VDD.n672 0.0458103
R3870 VDD.n1021 VDD.n1020 0.0449578
R3871 VDD.n1695 VDD.n1694 0.0449578
R3872 VDD.n2293 VDD.n2292 0.0444024
R3873 VDD.n2509 VDD.n2508 0.0444024
R3874 VDD.n1962 VDD.n1961 0.0440484
R3875 VDD.n1127 VDD.n1126 0.0419607
R3876 VDD.n1940 VDD.n1939 0.0414756
R3877 VDD.n1894 VDD.n1893 0.0414756
R3878 VDD.n126 VDD.n19 0.0414756
R3879 VDD.n77 VDD.n39 0.0414756
R3880 VDD.n2131 VDD.n2130 0.0414756
R3881 VDD.n1769 VDD.n169 0.0414381
R3882 VDD.n1765 VDD.n171 0.0412143
R3883 VDD.n1544 VDD.n307 0.0412143
R3884 VDD.n1537 VDD.n1536 0.0412143
R3885 VDD.n1241 VDD.n1240 0.0412143
R3886 VDD.n1233 VDD.n1200 0.0412143
R3887 VDD.n981 VDD.n980 0.0411452
R3888 VDD.n1744 VDD.n1743 0.0409494
R3889 VDD.n987 VDD.n582 0.0408043
R3890 VDD VDD.n1135 0.0397857
R3891 VDD.n996 VDD.n993 0.0395361
R3892 VDD.n992 VDD 0.0393983
R3893 VDD VDD.n1751 0.0376429
R3894 VDD.n829 VDD.n749 0.0375588
R3895 VDD.n1346 VDD.n1342 0.0375161
R3896 VDD.n2186 VDD.n2185 0.037431
R3897 VDD.n2135 VDD.n2134 0.0373601
R3898 VDD.n2164 VDD.n2103 0.0373601
R3899 VDD.n2383 VDD.n2382 0.0372474
R3900 VDD.n1515 VDD.n1514 0.0371667
R3901 VDD.n1298 VDD.n1293 0.0371667
R3902 VDD.n2384 VDD.n2189 0.0371207
R3903 VDD.n1765 VDD.n172 0.0369286
R3904 VDD.n466 VDD.n465 0.0369005
R3905 VDD.n2066 VDD.n2065 0.0368636
R3906 VDD.n2188 VDD.n2187 0.0368103
R3907 VDD.n899 VDD.n898 0.0367109
R3908 VDD.n2370 VDD.n2369 0.0366246
R3909 VDD.n2002 VDD.n2001 0.0365077
R3910 VDD.n2400 VDD.n2399 0.0365
R3911 VDD.n1973 VDD.n1972 0.0363784
R3912 VDD.n1526 VDD.n1525 0.0362955
R3913 VDD.n1119 VDD.n524 0.0362143
R3914 VDD.n220 VDD.n189 0.0362143
R3915 VDD.n792 VDD.n777 0.0359878
R3916 VDD VDD.n798 0.0359436
R3917 VDD.n774 VDD.n771 0.0357016
R3918 VDD.n819 VDD.n818 0.0357016
R3919 VDD.n1967 VDD.n5 0.0353113
R3920 VDD VDD.n1779 0.0353113
R3921 VDD.n1271 VDD.n1248 0.0352727
R3922 VDD.n792 VDD.n788 0.0348902
R3923 VDD.n798 VDD.n777 0.0348902
R3924 VDD.n1759 VDD.n179 0.034882
R3925 VDD.n1555 VDD.n1554 0.0347857
R3926 VDD.n818 VDD.n771 0.0346129
R3927 VDD.n2512 VDD.n2511 0.0341585
R3928 VDD.n761 VDD.n760 0.0340503
R3929 VDD.n1143 VDD.n509 0.0338708
R3930 VDD.n1100 VDD.n1099 0.0337609
R3931 VDD.n259 VDD.n258 0.0337609
R3932 VDD.n1222 VDD.n1221 0.0337143
R3933 VDD.n756 VDD.n748 0.0335178
R3934 VDD.n913 VDD.n912 0.0331389
R3935 VDD.n2665 VDD.n2664 0.0328077
R3936 VDD.n1828 VDD.n1819 0.0326951
R3937 VDD.n1913 VDD.n1912 0.0326951
R3938 VDD.n2160 VDD.n2159 0.0326951
R3939 VDD.n2623 VDD.n2622 0.0326951
R3940 VDD.n906 VDD.n884 0.0322736
R3941 VDD.n120 VDD.n35 0.0319634
R3942 VDD.n60 VDD.n59 0.0319634
R3943 VDD.n809 VDD.n774 0.0317097
R3944 VDD.n1349 VDD.n1342 0.0317097
R3945 VDD.n1940 VDD.n1806 0.0305
R3946 VDD.n1895 VDD.n1894 0.0305
R3947 VDD.n131 VDD.n19 0.0305
R3948 VDD.n77 VDD.n76 0.0305
R3949 VDD.n2131 VDD.n2127 0.0305
R3950 VDD.n2649 VDD.n2648 0.0305
R3951 VDD.n2667 VDD.n2666 0.0305
R3952 VDD.n911 VDD.n743 0.0301809
R3953 VDD.n693 VDD.n670 0.0299176
R3954 VDD.n905 VDD.n904 0.0292234
R3955 VDD.n909 VDD.n745 0.0292234
R3956 VDD.n910 VDD.n909 0.0292234
R3957 VDD.n1273 VDD.n1272 0.0291956
R3958 VDD.n1258 VDD.n1257 0.0291956
R3959 VDD.n1468 VDD.n1457 0.0291956
R3960 VDD.n1524 VDD.n314 0.0291956
R3961 VDD.n2003 VDD.n2002 0.0291726
R3962 VDD.n714 VDD.n657 0.0289211
R3963 VDD.n713 VDD.n712 0.0289211
R3964 VDD.n2045 VDD.n2044 0.028625
R3965 VDD.n985 VDD.n984 0.0278529
R3966 VDD.n971 VDD.n938 0.0278529
R3967 VDD.n762 VDD.n755 0.0277596
R3968 VDD.n2669 VDD.n2668 0.0276154
R3969 VDD.n2349 VDD.n2348 0.0274543
R3970 VDD.n757 VDD.n747 0.0273269
R3971 VDD.n1455 VDD.n344 0.0270909
R3972 VDD.n2364 VDD.n2363 0.0269975
R3973 VDD.n2388 VDD.n2387 0.0269444
R3974 VDD.n2591 VDD.n2391 0.0267222
R3975 VDD.n625 VDD.n586 0.0265748
R3976 VDD.n2390 VDD.n2389 0.0265
R3977 VDD.n908 VDD.n907 0.0264615
R3978 VDD.n908 VDD.n744 0.0264615
R3979 VDD.n2590 VDD.n2392 0.0264024
R3980 VDD.n2060 VDD.n2054 0.026375
R3981 VDD.n2386 VDD.n2385 0.0262778
R3982 VDD.n2589 VDD.n2545 0.0259067
R3983 VDD.n728 VDD.n625 0.0257336
R3984 VDD.n711 VDD.n660 0.0256417
R3985 VDD.n2522 VDD.n2521 0.0254761
R3986 VDD.n819 VDD.n753 0.0251774
R3987 VDD.n1918 VDD.n1845 0.0250455
R3988 VDD.n988 VDD.n581 0.0247707
R3989 VDD.n699 VDD.n698 0.0247609
R3990 VDD.n1102 VDD.n1101 0.0239783
R3991 VDD.n702 VDD.n701 0.0239783
R3992 VDD.n257 VDD.n216 0.0239783
R3993 VDD.n2171 VDD.n2170 0.0237258
R3994 VDD.n2170 VDD.n2168 0.0237258
R3995 VDD.n2168 VDD.n2102 0.0237258
R3996 VDD.n2102 VDD.n2100 0.0237258
R3997 VDD.n1767 VDD.n1766 0.0237036
R3998 VDD.n2063 VDD.n2026 0.0236818
R3999 VDD.n765 VDD.n764 0.0235488
R4000 VDD.n2137 VDD.n2136 0.0235375
R4001 VDD.n723 VDD.n633 0.0234555
R4002 VDD.n984 VDD.n915 0.0234412
R4003 VDD.n2163 VDD.n2162 0.0232304
R4004 VDD.n1556 VDD.n293 0.023
R4005 VDD.n1237 VDD.n1197 0.023
R4006 VDD.n1220 VDD.n1219 0.023
R4007 VDD.n2097 VDD.n2096 0.0229232
R4008 VDD.n737 VDD.n589 0.0227267
R4009 VDD.n973 VDD.n972 0.0225588
R4010 VDD.n970 VDD.n936 0.0225588
R4011 VDD.n610 VDD.n609 0.0223623
R4012 VDD.n1540 VDD.n311 0.0219286
R4013 VDD.n644 VDD.n643 0.0216336
R4014 VDD VDD.n1975 0.0214589
R4015 VDD.n742 VDD.n741 0.0206869
R4016 VDD.n1925 VDD.n1924 0.0203701
R4017 VDD.n1932 VDD.n1819 0.0202561
R4018 VDD.n1913 VDD.n1874 0.0202561
R4019 VDD.n125 VDD.n35 0.0202561
R4020 VDD.n59 VDD.n45 0.0202561
R4021 VDD.n2160 VDD.n2149 0.0202561
R4022 VDD.n2633 VDD.n2623 0.0202561
R4023 VDD.n669 VDD.n665 0.0200652
R4024 VDD.n703 VDD.n668 0.0200652
R4025 VDD.n1096 VDD.n1085 0.0200652
R4026 VDD.n1616 VDD.n1615 0.0200652
R4027 VDD.n2184 VDD.n2183 0.0200517
R4028 VDD.n17 VDD.n16 0.0200283
R4029 VDD.n740 VDD.n587 0.0198458
R4030 VDD.n2373 VDD.n2372 0.019808
R4031 VDD.n1609 VDD.n238 0.0197857
R4032 VDD.n1170 VDD.n1169 0.0197857
R4033 VDD.n2379 VDD.n2378 0.0194965
R4034 VDD.n903 VDD.n902 0.0191328
R4035 VDD.n691 VDD.n690 0.0191207
R4036 VDD.n696 VDD.n695 0.019083
R4037 VDD.n882 VDD.n832 0.0190047
R4038 VDD.n1175 VDD.n499 0.0187022
R4039 VDD.n974 VDD.n934 0.0186452
R4040 VDD.n969 VDD.n939 0.0186452
R4041 VDD.n2399 VDD.n2398 0.0185
R4042 VDD.n121 VDD.n120 0.018061
R4043 VDD.n61 VDD.n60 0.018061
R4044 VDD.n1782 VDD.n7 0.0180472
R4045 VDD.n1591 VDD.n1590 0.017691
R4046 VDD.n1152 VDD.n1151 0.0176429
R4047 VDD.n2366 VDD.n2296 0.0176235
R4048 VDD.n1956 VDD.n1788 0.0174811
R4049 VDD.n1829 VDD.n1828 0.0173293
R4050 VDD.n1912 VDD.n1911 0.0173293
R4051 VDD.n2159 VDD.n2158 0.0173293
R4052 VDD.n2622 VDD.n2621 0.0173293
R4053 VDD.n738 VDD.n588 0.0173224
R4054 VDD.n730 VDD.n729 0.0173224
R4055 VDD.n1769 VDD.n1768 0.0167254
R4056 VDD.n1441 VDD.n1440 0.0165976
R4057 VDD.n969 VDD.n968 0.0164677
R4058 VDD.n2402 VDD.n2400 0.0161
R4059 VDD.n831 VDD.n747 0.0160453
R4060 VDD.n760 VDD.n759 0.0159438
R4061 VDD.n759 VDD.n756 0.0159438
R4062 VDD.n830 VDD.n748 0.0159438
R4063 VDD VDD.n1818 0.0158659
R4064 VDD VDD.n1846 0.0158659
R4065 VDD VDD.n138 0.0158659
R4066 VDD.n69 VDD 0.0158659
R4067 VDD VDD.n2141 0.0158659
R4068 VDD.n2639 VDD 0.0158659
R4069 VDD.n989 VDD.n579 0.0157992
R4070 VDD.n653 VDD.n626 0.0156402
R4071 VDD.n880 VDD.n879 0.0156402
R4072 VDD.n983 VDD.n982 0.015009
R4073 VDD.n689 VDD.n671 0.0149
R4074 VDD.n2013 VDD 0.0147661
R4075 VDD.n2361 VDD.n2360 0.0146624
R4076 VDD.n2162 VDD.n2161 0.0146297
R4077 VDD.n2526 VDD.n2525 0.0141098
R4078 VDD.n688 VDD.n672 0.014
R4079 VDD.n2531 VDD.n2530 0.0138902
R4080 VDD.n2396 VDD.n2395 0.0138493
R4081 VDD.n1771 VDD.n1770 0.0136831
R4082 VDD.n1431 VDD.n1430 0.0136707
R4083 VDD.n1433 VDD.n1432 0.0136707
R4084 VDD.n444 VDD.n443 0.0136707
R4085 VDD.n1365 VDD.n1364 0.0136707
R4086 VDD VDD.n2346 0.0136707
R4087 VDD.n974 VDD.n918 0.0135645
R4088 VDD.n763 VDD.n762 0.0130481
R4089 VDD.n758 VDD.n755 0.0130481
R4090 VDD.n758 VDD.n757 0.0130481
R4091 VDD.n1765 VDD.n1764 0.0122692
R4092 VDD.n582 VDD.n580 0.0122391
R4093 VDD.n597 VDD.n596 0.0121599
R4094 VDD.n981 VDD.n917 0.0121129
R4095 VDD.n982 VDD.n916 0.0119706
R4096 VDD.n683 VDD.n678 0.0118445
R4097 VDD.n320 VDD.n318 0.01175
R4098 VDD.n1729 VDD.n1728 0.0116236
R4099 VDD.n653 VDD.n624 0.0114346
R4100 VDD.n1545 VDD.n305 0.0112143
R4101 VDD.n2167 VDD.n2166 0.0110882
R4102 VDD.n2296 VDD.n2295 0.0110076
R4103 VDD.n2540 VDD.n2538 0.0108349
R4104 VDD.n1270 VDD.n1269 0.0107273
R4105 VDD.n1061 VDD.n538 0.0106124
R4106 VDD.n879 VDD.n878 0.0105935
R4107 VDD.n2005 VDD.n2004 0.0104739
R4108 VDD.n2017 VDD.n1975 0.0103769
R4109 VDD.n2058 VDD.n2057 0.0103544
R4110 VDD.n1232 VDD.n1207 0.0101429
R4111 VDD.n761 VDD.n754 0.0100858
R4112 VDD.n824 VDD.n753 0.00993548
R4113 VDD.n2372 VDD.n2371 0.00984256
R4114 VDD.n739 VDD.n738 0.00975234
R4115 VDD.n2380 VDD.n2379 0.00953114
R4116 VDD.n2516 VDD.n2515 0.00932775
R4117 VDD.n1388 VDD 0.00932353
R4118 VDD.n898 VDD.n746 0.00928906
R4119 VDD.n871 VDD.n836 0.00928049
R4120 VDD.n877 VDD.n833 0.00928049
R4121 VDD.n730 VDD.n588 0.00891121
R4122 VDD.n2374 VDD.n2373 0.0089083
R4123 VDD.n600 VDD.n599 0.00888057
R4124 VDD.n2378 VDD.n2377 0.00859689
R4125 VDD.n875 VDD.n836 0.00854878
R4126 VDD.n877 VDD.n876 0.00854878
R4127 VDD.n825 VDD.n752 0.00853674
R4128 VDD.n725 VDD.n724 0.00851619
R4129 VDD.n2355 VDD.n2354 0.0082665
R4130 VDD.n688 VDD.n683 0.00806303
R4131 VDD.n2165 VDD.n2164 0.00787201
R4132 VDD.n2336 VDD.n2335 0.00781707
R4133 VDD.n2579 VDD.n2578 0.00781707
R4134 VDD.n644 VDD.n623 0.00778745
R4135 VDD.n442 VDD.n441 0.00775806
R4136 VDD.n1367 VDD.n1366 0.00775806
R4137 VDD.n986 VDD.n583 0.00754348
R4138 VDD.n657 VDD.n633 0.00742308
R4139 VDD.n712 VDD.n711 0.00742308
R4140 VDD.n596 VDD.n589 0.00742308
R4141 VDD.n2515 VDD.n2514 0.00738995
R4142 VDD.n917 VDD.n581 0.00738437
R4143 VDD.n2362 VDD.n2361 0.00735279
R4144 VDD.n2059 VDD.n2055 0.00725
R4145 VDD.n2059 VDD.n2058 0.00725
R4146 VDD.n788 VDD.n787 0.00708537
R4147 VDD.n2328 VDD.n2327 0.00708537
R4148 VDD.n2571 VDD.n2570 0.00708537
R4149 VDD.n2525 VDD.n2524 0.00708537
R4150 VDD.n612 VDD.n610 0.0070587
R4151 VDD.n654 VDD.n627 0.0070587
R4152 VDD.n1014 VDD.n1013 0.00700602
R4153 VDD.n1704 VDD.n1703 0.00700602
R4154 VDD.n2530 VDD.n2529 0.00686585
R4155 VDD.n737 VDD.n736 0.00669433
R4156 VDD.n2360 VDD.n2359 0.00666751
R4157 VDD.n2354 VDD.n2353 0.00666751
R4158 VDD.n928 VDD.n924 0.00661998
R4159 VDD.n2356 VDD.n2355 0.00643909
R4160 VDD.n2527 VDD.n2526 0.00642683
R4161 VDD.n598 VDD.n587 0.00638785
R4162 VDD.n714 VDD.n713 0.00632996
R4163 VDD.n706 VDD.n705 0.00632996
R4164 VDD.n704 VDD.n667 0.00632996
R4165 VDD.n613 VDD.n600 0.00632996
R4166 VDD.n2397 VDD.n2396 0.0063134
R4167 VDD VDD.n1423 0.00630645
R4168 VDD.n432 VDD 0.00630645
R4169 VDD VDD.n401 0.00630645
R4170 VDD VDD.n862 0.00630645
R4171 VDD.n961 VDD 0.00630645
R4172 VDD VDD.n372 0.00630645
R4173 VDD.n2532 VDD.n2531 0.00620732
R4174 VDD.n2538 VDD.n2537 0.00609809
R4175 VDD.n2352 VDD.n2351 0.00598223
R4176 VDD.n765 VDD.n754 0.00582544
R4177 VDD.n973 VDD.n935 0.00579412
R4178 VDD.n598 VDD.n585 0.00572908
R4179 VDD.n2181 VDD.n2180 0.00562658
R4180 VDD.n876 VDD.n875 0.00562195
R4181 VDD.n983 VDD.n583 0.00558696
R4182 VDD.n1784 VDD.n1783 0.00531132
R4183 VDD.n2543 VDD.n2542 0.00523684
R4184 VDD.n2517 VDD.n2516 0.00522019
R4185 VDD.n2017 VDD.n2016 0.0050197
R4186 VDD.n878 VDD.n834 0.00489628
R4187 VDD.n654 VDD.n652 0.00487247
R4188 VDD.n987 VDD.n986 0.00480435
R4189 VDD.n2403 VDD.n2402 0.00467073
R4190 VDD.n652 VDD.n651 0.0045081
R4191 VDD.n725 VDD.n627 0.0045081
R4192 VDD.n700 VDD.n668 0.00441304
R4193 VDD.n697 VDD.n696 0.00414372
R4194 VDD.n731 VDD.n590 0.00414372
R4195 VDD.n827 VDD.n751 0.00412903
R4196 VDD.n980 VDD.n918 0.00412903
R4197 VDD.n937 VDD.n915 0.00402941
R4198 VDD.n972 VDD.n936 0.00402941
R4199 VDD.n2046 VDD.n2045 0.003875
R4200 VDD.n2016 VDD.n2015 0.00380882
R4201 VDD.n706 VDD.n660 0.00377935
R4202 VDD.n695 VDD.n667 0.00377935
R4203 VDD.n614 VDD.n612 0.00377935
R4204 VDD.n767 VDD.n751 0.00376613
R4205 VDD.n1550 VDD.n1549 0.00371429
R4206 VDD.n1228 VDD.n1227 0.00371429
R4207 VDD.n580 VDD.n579 0.00360796
R4208 VDD.n766 VDD.n752 0.00350186
R4209 VDD.n651 VDD.n643 0.00341498
R4210 VDD VDD.n809 0.00340323
R4211 VDD.n939 VDD.n934 0.00340323
R4212 VDD.n2366 VDD.n2365 0.00326137
R4213 VDD.n614 VDD.n613 0.00305061
R4214 VDD.n599 VDD.n597 0.00305061
R4215 VDD.n827 VDD.n826 0.00304032
R4216 VDD.n2518 VDD.n2517 0.00301846
R4217 VDD.n2402 VDD.n2401 0.0029
R4218 VDD.n2541 VDD 0.00286842
R4219 VDD.n2053 VDD.n2047 0.00283766
R4220 VDD.n726 VDD.n626 0.00283401
R4221 VDD.n2054 VDD.n2046 0.00275
R4222 VDD.n2345 VDD.n2344 0.00269512
R4223 VDD.n2588 VDD.n2587 0.00269512
R4224 VDD.n999 VDD.n998 0.00266867
R4225 VDD.n1669 VDD.n1665 0.00266867
R4226 VDD.n689 VDD 0.00254545
R4227 VDD.n923 VDD.n917 0.00254545
R4228 VDD.n724 VDD.n723 0.00245652
R4229 VDD.n703 VDD.n665 0.00206522
R4230 VDD.n2187 VDD.n2186 0.00205172
R4231 VDD.n2542 VDD.n2541 0.00200718
R4232 VDD.n2347 VDD 0.00196341
R4233 VDD.n1637 VDD.n208 0.00192857
R4234 VDD.n2036 VDD 0.00186364
R4235 VDD.n2353 VDD.n2352 0.00164213
R4236 VDD.n2389 VDD.n2388 0.00161111
R4237 VDD.n736 VDD.n590 0.00159312
R4238 VDD.n731 VDD.n623 0.00159312
R4239 VDD.n1262 VDD.n1260 0.00152273
R4240 VDD.n1465 VDD.n1464 0.00152273
R4241 VDD.n990 VDD 0.00151695
R4242 VDD.n1784 VDD 0.00134906
R4243 VDD.n1768 VDD.n170 0.00132534
R4244 VDD.n2520 VDD.n2519 0.00132296
R4245 VDD.n1919 VDD.n1790 0.00129295
R4246 VDD.n1943 VDD.n1942 0.00129295
R4247 VDD.n1801 VDD 0.00128947
R4248 VDD.n1856 VDD 0.00128947
R4249 VDD.n30 VDD 0.00128947
R4250 VDD.n87 VDD 0.00128947
R4251 VDD.n2115 VDD 0.00128947
R4252 VDD.n2659 VDD 0.00128947
R4253 VDD.n705 VDD.n704 0.00122874
R4254 VDD.n968 VDD.n940 0.00122581
R4255 VDD.n1053 VDD.n1052 0.00121429
R4256 VDD.n2376 VDD.n2375 0.00112284
R4257 VDD.n2377 VDD.n2376 0.00112284
R4258 VDD.n2521 VDD.n2520 0.00110765
R4259 VDD.n766 VDD.n765 0.00103254
R4260 VDD.n2077 VDD.n2076 0.00101724
R4261 VDD.n924 VDD.n923 0.00101136
R4262 VDD.n2358 VDD.n2357 0.000956853
R4263 VDD.n2357 VDD.n2356 0.000956853
R4264 VDD.n2534 VDD.n2533 0.000939024
R4265 VDD.n2533 VDD.n2532 0.000939024
R4266 VDD.n2536 VDD.n2535 0.000930622
R4267 VDD.n2537 VDD.n2536 0.000930622
R4268 VDD VDD.n2540 0.000930622
R4269 VDD.n824 VDD.n767 0.000862903
R4270 VDD.n902 VDD 0.000851563
R4271 VDD.n2368 VDD.n2367 0.000811419
R4272 VDD.n2369 VDD.n2368 0.000811419
R4273 VDD.n2371 VDD.n2370 0.000811419
R4274 VDD.n2375 VDD.n2374 0.000811419
R4275 VDD.n2381 VDD.n2380 0.000811419
R4276 VDD.n2382 VDD.n2381 0.000811419
R4277 VDD.n2185 VDD.n2184 0.000810345
R4278 VDD.n2189 VDD.n2188 0.000810345
R4279 VDD.n2365 VDD.n2364 0.000728426
R4280 VDD.n2363 VDD.n2362 0.000728426
R4281 VDD.n2359 VDD.n2358 0.000728426
R4282 VDD.n2351 VDD.n2350 0.000728426
R4283 VDD.n2350 VDD.n2349 0.000728426
R4284 VDD.n2387 VDD.n2386 0.000722222
R4285 VDD.n2391 VDD.n2390 0.000722222
R4286 VDD.n2524 VDD.n2403 0.000719512
R4287 VDD.n2534 VDD.n2527 0.000719512
R4288 VDD.n2529 VDD.n2528 0.000719512
R4289 VDD.n2528 VDD.n2392 0.000719512
R4290 VDD.n2519 VDD.n2518 0.000715311
R4291 VDD.n2523 VDD.n2522 0.000715311
R4292 VDD.n2535 VDD.n2397 0.000715311
R4293 VDD.n2544 VDD.n2543 0.000715311
R4294 VDD.n2545 VDD.n2544 0.000715311
R4295 PFD_T2_0.INV_mag_1.IN.n9 PFD_T2_0.INV_mag_1.IN.t6 226.316
R4296 PFD_T2_0.INV_mag_1.IN.n6 PFD_T2_0.INV_mag_1.IN.t26 116.993
R4297 PFD_T2_0.INV_mag_1.IN.n30 PFD_T2_0.INV_mag_1.IN.t32 33.8279
R4298 PFD_T2_0.INV_mag_1.IN.n31 PFD_T2_0.INV_mag_1.IN.n30 30.2144
R4299 PFD_T2_0.INV_mag_1.IN.t28 PFD_T2_0.INV_mag_1.IN.n3 25.0458
R4300 PFD_T2_0.INV_mag_1.IN.n28 PFD_T2_0.INV_mag_1.IN.n27 16.5048
R4301 PFD_T2_0.INV_mag_1.IN.n29 PFD_T2_0.INV_mag_1.IN.n28 16.5048
R4302 PFD_T2_0.INV_mag_1.IN.n3 PFD_T2_0.INV_mag_1.IN.t23 15.3305
R4303 PFD_T2_0.INV_mag_1.IN.n4 PFD_T2_0.INV_mag_1.IN.t29 15.1914
R4304 PFD_T2_0.INV_mag_1.IN.n3 PFD_T2_0.INV_mag_1.IN.n31 12.8616
R4305 PFD_T2_0.INV_mag_1.IN.n4 PFD_T2_0.INV_mag_1.IN.t21 12.6987
R4306 PFD_T2_0.INV_mag_1.IN.n5 PFD_T2_0.INV_mag_1.IN.t28 12.1515
R4307 PFD_T2_0.INV_mag_1.IN.t19 PFD_T2_0.INV_mag_1.IN.n6 11.3159
R4308 PFD_T2_0.INV_mag_1.IN.n9 PFD_T2_0.INV_mag_1.IN.t8 10.9468
R4309 PFD_T2_0.INV_mag_1.IN.n6 PFD_T2_0.INV_mag_1.IN.t17 10.2935
R4310 PFD_T2_0.INV_mag_1.IN.n0 PFD_T2_0.INV_mag_1.IN.n4 10.261
R4311 PFD_T2_0.INV_mag_1.IN.n27 PFD_T2_0.INV_mag_1.IN.t33 9.4175
R4312 PFD_T2_0.INV_mag_1.IN.n28 PFD_T2_0.INV_mag_1.IN.t20 9.4175
R4313 PFD_T2_0.INV_mag_1.IN.t23 PFD_T2_0.INV_mag_1.IN.n29 9.4175
R4314 PFD_T2_0.INV_mag_1.IN.n27 PFD_T2_0.INV_mag_1.IN.t22 9.1985
R4315 PFD_T2_0.INV_mag_1.IN.n28 PFD_T2_0.INV_mag_1.IN.t27 9.1985
R4316 PFD_T2_0.INV_mag_1.IN.n29 PFD_T2_0.INV_mag_1.IN.t30 9.1985
R4317 PFD_T2_0.INV_mag_1.IN.n3 PFD_T2_0.INV_mag_1.IN.t24 8.05323
R4318 PFD_T2_0.INV_mag_1.IN.n21 PFD_T2_0.INV_mag_1.IN.n18 6.76657
R4319 PFD_T2_0.INV_mag_1.IN.n1 PFD_T2_0.INV_mag_1.IN.n10 6.46231
R4320 PFD_T2_0.INV_mag_1.IN.n21 PFD_T2_0.INV_mag_1.IN.n20 5.58741
R4321 PFD_T2_0.INV_mag_1.IN.n26 PFD_T2_0.INV_mag_1.IN.n14 5.17308
R4322 PFD_T2_0.INV_mag_1.IN.n1 PFD_T2_0.INV_mag_1.IN.n9 4.73858
R4323 PFD_T2_0.INV_mag_1.IN.n30 PFD_T2_0.INV_mag_1.IN.t25 3.6505
R4324 PFD_T2_0.INV_mag_1.IN.n31 PFD_T2_0.INV_mag_1.IN.t18 3.6505
R4325 PFD_T2_0.INV_mag_1.IN.n24 PFD_T2_0.INV_mag_1.IN.t16 3.6405
R4326 PFD_T2_0.INV_mag_1.IN.n24 PFD_T2_0.INV_mag_1.IN.n23 3.6405
R4327 PFD_T2_0.INV_mag_1.IN.n14 PFD_T2_0.INV_mag_1.IN.t10 3.6405
R4328 PFD_T2_0.INV_mag_1.IN.n14 PFD_T2_0.INV_mag_1.IN.n13 3.6405
R4329 PFD_T2_0.INV_mag_1.IN.n12 PFD_T2_0.INV_mag_1.IN.t4 3.6405
R4330 PFD_T2_0.INV_mag_1.IN.n12 PFD_T2_0.INV_mag_1.IN.n11 3.6405
R4331 PFD_T2_0.INV_mag_1.IN.n8 PFD_T2_0.INV_mag_1.IN.t9 3.6405
R4332 PFD_T2_0.INV_mag_1.IN.n8 PFD_T2_0.INV_mag_1.IN.n7 3.6405
R4333 PFD_T2_0.INV_mag_1.IN.n16 PFD_T2_0.INV_mag_1.IN.t11 3.6405
R4334 PFD_T2_0.INV_mag_1.IN.n16 PFD_T2_0.INV_mag_1.IN.n15 3.6405
R4335 PFD_T2_0.INV_mag_1.IN.n20 PFD_T2_0.INV_mag_1.IN.t15 3.6405
R4336 PFD_T2_0.INV_mag_1.IN.n20 PFD_T2_0.INV_mag_1.IN.n19 3.6405
R4337 PFD_T2_0.INV_mag_1.IN.n18 PFD_T2_0.INV_mag_1.IN.t14 3.2765
R4338 PFD_T2_0.INV_mag_1.IN.n18 PFD_T2_0.INV_mag_1.IN.n17 3.2765
R4339 PFD_T2_0.INV_mag_1.IN.n2 PFD_T2_0.INV_mag_1.IN.n26 3.17603
R4340 PFD_T2_0.INV_mag_1.IN.n26 PFD_T2_0.INV_mag_1.IN.n25 3.15378
R4341 PFD_T2_0.INV_mag_1.IN.n1 PFD_T2_0.INV_mag_1.IN.n8 2.94791
R4342 PFD_T2_0.INV_mag_1.IN.n22 PFD_T2_0.INV_mag_1.IN.n16 2.92863
R4343 PFD_T2_0.INV_mag_1.IN.n2 PFD_T2_0.INV_mag_1.IN.n12 2.6005
R4344 PFD_T2_0.INV_mag_1.IN.n25 PFD_T2_0.INV_mag_1.IN.n24 2.6005
R4345 PFD_T2_0.INV_mag_1.IN.n22 PFD_T2_0.INV_mag_1.IN.n21 2.26925
R4346 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.IN.n0 6.76224
R4347 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.IN.t19 4.69745
R4348 PFD_T2_0.INV_mag_1.IN.n0 PFD_T2_0.INV_mag_1.IN.n5 2.6584
R4349 PFD_T2_0.INV_mag_1.IN.n2 PFD_T2_0.INV_mag_1.IN.n1 1.0806
R4350 PFD_T2_0.INV_mag_1.IN.n5 PFD_T2_0.INV_mag_1.IN.n2 1.06506
R4351 PFD_T2_0.INV_mag_1.IN.n25 PFD_T2_0.INV_mag_1.IN.n22 1.00114
R4352 VSS.n4692 VSS.n4691 5.941e+06
R4353 VSS.n5384 VSS.n5383 5.93775e+06
R4354 VSS.n6985 VSS.t531 529014
R4355 VSS.n6717 VSS.n6709 19252.4
R4356 VSS.n4693 VSS.n4692 15212.8
R4357 VSS.t122 VSS.n1102 11524.5
R4358 VSS.n1731 VSS.n1730 11359.2
R4359 VSS.t337 VSS.n6971 9017.72
R4360 VSS.t122 VSS.t275 8844.94
R4361 VSS.n5961 VSS.n5960 7554.82
R4362 VSS.n1085 VSS.n1084 6960.92
R4363 VSS.t278 VSS.n831 6723.04
R4364 VSS.n6718 VSS.n6717 5785.45
R4365 VSS.n5960 VSS.n5959 4779.81
R4366 VSS.n1103 VSS.t124 4264.65
R4367 VSS.n7709 VSS.n7708 4047.38
R4368 VSS.n832 VSS.t68 3914.93
R4369 VSS.n6696 VSS.n6695 3820.73
R4370 VSS.t95 VSS.t93 3546.42
R4371 VSS.n1730 VSS.n1729 3501.04
R4372 VSS.n1003 VSS.n1002 3439.15
R4373 VSS.n4691 VSS.n4690 3301.18
R4374 VSS.n7710 VSS.n7709 3049.35
R4375 VSS.t275 VSS.t128 2797.47
R4376 VSS.n830 VSS.t273 2454.64
R4377 VSS.n5385 VSS.n5384 2225.75
R4378 VSS.t93 VSS.t96 2159.61
R4379 VSS.t234 VSS.t150 1822.88
R4380 VSS.t427 VSS.t715 1805.06
R4381 VSS.t839 VSS.n7297 1796.6
R4382 VSS.t447 VSS.t847 1778.39
R4383 VSS.n765 VSS.t234 1720.94
R4384 VSS.n1729 VSS.n1728 1678.53
R4385 VSS.t459 VSS.t203 1657.99
R4386 VSS.t435 VSS.t172 1649.75
R4387 VSS.n4636 VSS.t141 1557.29
R4388 VSS.t124 VSS.t246 1524.86
R4389 VSS.t68 VSS.t277 1520.6
R4390 VSS.n5506 VSS.n5505 1514.17
R4391 VSS.t836 VSS.t834 1510.25
R4392 VSS.t31 VSS.t836 1510.25
R4393 VSS.n7251 VSS.t95 1407.98
R4394 VSS.n5118 VSS.t447 1404.92
R4395 VSS.n7793 VSS.n7792 1377.01
R4396 VSS.n7868 VSS.t427 1316.01
R4397 VSS.n5101 VSS.t435 1303.3
R4398 VSS.n4770 VSS.t480 1229.06
R4399 VSS.n7851 VSS.t475 1229.06
R4400 VSS.n5101 VSS.t368 1224.94
R4401 VSS.t847 VSS.t204 1209.3
R4402 VSS.t715 VSS.t931 1209.3
R4403 VSS.n7799 VSS.n7798 1196.37
R4404 VSS.t172 VSS.t933 1121.83
R4405 VSS.t203 VSS.t932 1121.83
R4406 VSS.n804 VSS.n803 1110.55
R4407 VSS.n6716 VSS.t74 1061.73
R4408 VSS.n6710 VSS.t995 967.024
R4409 VSS.n668 VSS.n667 953.981
R4410 VSS.n238 VSS.n237 944.048
R4411 VSS.n1563 VSS.n1562 929.726
R4412 VSS.n4356 VSS.n4355 928.664
R4413 VSS.t246 VSS.t122 928.572
R4414 VSS.t277 VSS.t278 925.979
R4415 VSS.n7299 VSS.t534 878.801
R4416 VSS.t391 VSS.t802 855.827
R4417 VSS.n6390 VSS.n6389 804.534
R4418 VSS.n4983 VSS.t432 617.99
R4419 VSS.t729 VSS.t727 581.962
R4420 VSS.t748 VSS.t729 581.962
R4421 VSS.t757 VSS.t748 581.962
R4422 VSS.t819 VSS.t779 581.962
R4423 VSS.t779 VSS.t795 581.962
R4424 VSS.n7269 VSS.n7268 571.124
R4425 VSS.n745 VSS.t65 561.086
R4426 VSS.t534 VSS.t6 530.4
R4427 VSS.t6 VSS.t908 530.4
R4428 VSS.n6974 VSS.t325 490.178
R4429 VSS.n333 VSS.n332 477.231
R4430 VSS.n7394 VSS.n7393 431.716
R4431 VSS.n5962 VSS.n5961 431.19
R4432 VSS.n7298 VSS.t907 426.401
R4433 VSS.n4837 VSS.t757 421.495
R4434 VSS.n418 VSS.n417 407.524
R4435 VSS.n6987 VSS.t993 390.616
R4436 VSS.n6986 VSS.t992 390.616
R4437 VSS.t556 VSS.t528 389.693
R4438 VSS.t940 VSS.t558 389.693
R4439 VSS.n6972 VSS.t337 321.293
R4440 VSS.n5041 VSS.t800 297.88
R4441 VSS.t185 VSS.t175 289.267
R4442 VSS.t208 VSS.t62 289.267
R4443 VSS.n4993 VSS.t734 288.988
R4444 VSS.n6717 VSS.n6716 279.142
R4445 VSS.n5066 VSS.t374 266.759
R4446 VSS.n831 VSS.n830 265.524
R4447 VSS.n6809 VSS.t550 261.829
R4448 VSS.n4996 VSS.t736 253.421
R4449 VSS.n5038 VSS.t786 244.529
R4450 VSS.n6763 VSS.t9 236.893
R4451 VSS.n6554 VSS.t562 211.958
R4452 VSS.n4317 VSS.t33 211.279
R4453 VSS.n4336 VSS.t314 197.1
R4454 VSS.n6697 VSS.n6696 195.54
R4455 VSS.n4312 VSS.t169 194.263
R4456 VSS.n6509 VSS.t344 191.77
R4457 VSS.n5179 VSS.t930 191.177
R4458 VSS.n5054 VSS.t399 186.731
R4459 VSS.n5060 VSS.t5 182.286
R4460 VSS.t48 VSS.t543 180.655
R4461 VSS.n4291 VSS.t181 180.083
R4462 VSS.n4307 VSS.t292 177.248
R4463 VSS.t46 VSS.n1725 165.6
R4464 VSS.n4980 VSS.t810 164.501
R4465 VSS.n4295 VSS.t178 163.067
R4466 VSS.n6756 VSS.t71 162.084
R4467 VSS.n4837 VSS.t819 160.468
R4468 VSS.n4304 VSS.t323 160.232
R4469 VSS.n7321 VSS.n7320 159.956
R4470 VSS.n4285 VSS.t189 157.395
R4471 VSS.n76 VSS.t146 154.649
R4472 VSS.n4299 VSS.t316 146.052
R4473 VSS.n4357 VSS.n4356 145.571
R4474 VSS.n4299 VSS.t295 143.216
R4475 VSS.n5963 VSS.n5962 137.738
R4476 VSS.n279 VSS.t28 137.732
R4477 VSS.n6644 VSS.t167 137.149
R4478 VSS.t18 VSS.t25 134.906
R4479 VSS.n270 VSS.n269 132.9
R4480 VSS.n1712 VSS.t50 131.948
R4481 VSS.n6502 VSS.t266 131.212
R4482 VSS.n833 VSS.n832 130.123
R4483 VSS.n4304 VSS.t192 129.036
R4484 VSS.n5019 VSS.t967 128.934
R4485 VSS.n1286 VSS.n1285 127.87
R4486 VSS.n7828 VSS.t164 127.856
R4487 VSS.n4295 VSS.t195 126.201
R4488 VSS.n7488 VSS.n7487 125.534
R4489 VSS.n1629 VSS.t10 123.094
R4490 VSS.n6997 VSS.n6996 122.472
R4491 VSS.n1695 VSS.t12 121.323
R4492 VSS.n4947 VSS.t783 120.041
R4493 VSS.n395 VSS.n394 116.502
R4494 VSS.n4599 VSS.t113 115.596
R4495 VSS.n6502 VSS.n6501 114.389
R4496 VSS.n1748 VSS.t365 112.466
R4497 VSS.n6625 VSS.t168 112.213
R4498 VSS.n4307 VSS.t185 112.02
R4499 VSS.n6547 VSS.t561 111.025
R4500 VSS.n1693 VSS.t301 110.695
R4501 VSS.n118 VSS.n117 109.445
R4502 VSS.n4291 VSS.t200 109.184
R4503 VSS.t245 VSS.n6749 108.056
R4504 VSS.n7395 VSS.n7394 104.55
R4505 VSS.n1754 VSS.t410 101.84
R4506 VSS.n1726 VSS.t46 100.069
R4507 VSS.n6672 VSS.t822 99.7447
R4508 VSS.n1731 VSS.t357 98.2975
R4509 VSS.n4312 VSS.t309 95.0049
R4510 VSS.n4286 VSS.t288 92.1689
R4511 VSS.n4336 VSS.t208 92.1689
R4512 VSS.n1687 VSS.t483 91.213
R4513 VSS.t343 VSS.n6494 90.839
R4514 VSS.n1687 VSS.t103 89.4419
R4515 VSS.t139 VSS.t54 88.6679
R4516 VSS.n6401 VSS.t903 87.4746
R4517 VSS.n7742 VSS.n7741 87.2286
R4518 VSS.n7378 VSS.n7376 86.7869
R4519 VSS.n5605 VSS.t240 81.8473
R4520 VSS.n6522 VSS.t915 80.7458
R4521 VSS.n1726 VSS.t490 80.5863
R4522 VSS.n4170 VSS.n4169 79.7008
R4523 VSS.n1754 VSS.t101 78.8152
R4524 VSS.n4317 VSS.t183 77.9892
R4525 VSS.n4320 VSS.t216 75.1532
R4526 VSS.n831 VSS.t125 74.368
R4527 VSS.t939 VSS.n7298 73.1207
R4528 VSS.n396 VSS.n395 71.3171
R4529 VSS.n7807 VSS.t306 70.1147
R4530 VSS.n1693 VSS.t48 69.9596
R4531 VSS.n7746 VSS.n7745 69.1814
R4532 VSS.n614 VSS.t116 68.7194
R4533 VSS.n664 VSS.t339 68.7194
R4534 VSS.n1516 VSS.t249 68.7194
R4535 VSS.n1573 VSS.t879 68.7194
R4536 VSS.n1748 VSS.t382 68.1885
R4537 VSS.n5173 VSS.t171 66.69
R4538 VSS.n81 VSS.t142 64.2392
R4539 VSS.n7783 VSS.n7782 63.1657
R4540 VSS.n6785 VSS.t36 62.3407
R4541 VSS.n4171 VSS.n4170 61.9333
R4542 VSS.n5229 VSS.t227 61.866
R4543 VSS.n4334 VSS.t258 60.9734
R4544 VSS.n288 VSS.t22 60.4094
R4545 VSS.n1695 VSS.t43 59.3329
R4546 VSS.n7297 VSS.n7296 58.9653
R4547 VSS.n4315 VSS.t197 58.1375
R4548 VSS.n5512 VSS.t536 57.9753
R4549 VSS.n5587 VSS.t912 57.9753
R4550 VSS.n5546 VSS.t224 57.9753
R4551 VSS.n5167 VSS.t714 57.798
R4552 VSS.n5188 VSS.t385 57.798
R4553 VSS.n1732 VSS.t377 57.5618
R4554 VSS.n1629 VSS.t580 57.5618
R4555 VSS.n6933 VSS.t948 56.4521
R4556 VSS.n5323 VSS.t133 53.2263
R4557 VSS.n6147 VSS.t360 51.6521
R4558 VSS.n5483 VSS.t59 51.1548
R4559 VSS.n5596 VSS.t547 51.1548
R4560 VSS.n6446 VSS.t987 50.4663
R4561 VSS.n6656 VSS.t551 49.8726
R4562 VSS.n6219 VSS.t504 49.6265
R4563 VSS.n4637 VSS.n4636 49.1159
R4564 VSS.n1712 VSS.t108 48.7062
R4565 VSS.n6971 VSS.n6970 47.1997
R4566 VSS.n1622 VSS.t88 46.9351
R4567 VSS.n4358 VSS.n4357 45.2213
R4568 VSS.n7623 VSS.t158 45.1618
R4569 VSS.n5330 VSS.n5329 45.1618
R4570 VSS.n7217 VSS.t767 43.9924
R4571 VSS.n4288 VSS.t211 43.9577
R4572 VSS.n6421 VSS.n6420 43.7376
R4573 VSS.n1311 VSS.n1310 42.6234
R4574 VSS.n5696 VSS.t19 41.5243
R4575 VSS.n5798 VSS.t350 41.5243
R4576 VSS.n4310 VSS.t187 41.1218
R4577 VSS.n5557 VSS.n5556 40.9239
R4578 VSS.n6535 VSS.t904 40.3732
R4579 VSS.n5282 VSS.n5281 39.8468
R4580 VSS.n7378 VSS.n7377 38.9047
R4581 VSS.n1625 VSS.t706 38.0795
R4582 VSS.n5483 VSS.t136 37.5136
R4583 VSS.n7556 VSS.n7555 37.1434
R4584 VSS.n7522 VSS.n7521 37.1241
R4585 VSS.n1631 VSS.t90 36.3084
R4586 VSS.n4237 VSS.t466 36.0467
R4587 VSS.n4248 VSS.t362 36.0467
R4588 VSS.n1641 VSS.t356 36.0467
R4589 VSS.n1652 VSS.t496 36.0467
R4590 VSS.n6123 VSS.t78 35.4477
R4591 VSS.n7565 VSS.t159 34.2862
R4592 VSS.n6047 VSS.n6046 33.4221
R4593 VSS.n4494 VSS.n4493 32.9568
R4594 VSS.n5512 VSS.t56 30.6931
R4595 VSS.n6922 VSS.n6920 30.6457
R4596 VSS.n6929 VSS.t119 30.6457
R4597 VSS.n7236 VSS.t53 30.1002
R4598 VSS.n1375 VSS.n1374 29.9489
R4599 VSS.n6734 VSS.n6733 29.0926
R4600 VSS.n780 VSS.t110 28.751
R4601 VSS.n1473 VSS.n1472 28.7316
R4602 VSS.n6066 VSS.t722 28.3582
R4603 VSS.n1734 VSS.t298 27.4528
R4604 VSS.n1628 VSS.t0 27.4528
R4605 VSS.n5563 VSS.t347 27.2828
R4606 VSS.n4293 VSS.t214 26.942
R4607 VSS.n5838 VSS.t797 26.3327
R4608 VSS.n7236 VSS.n7235 26.2413
R4609 VSS.n4502 VSS.n4501 26.1965
R4610 VSS.n228 VSS.t148 26.1718
R4611 VSS.n309 VSS.n308 26.0884
R4612 VSS.n1694 VSS.t99 25.6817
R4613 VSS.n4493 VSS.t18 25.3911
R4614 VSS.n759 VSS.t79 25.3179
R4615 VSS.n294 VSS.t15 24.1641
R4616 VSS.t175 VSS.n4306 24.1061
R4617 VSS.n5256 VSS.t921 23.0103
R4618 VSS.n4237 VSS.t421 22.6305
R4619 VSS.n4238 VSS.t515 22.6305
R4620 VSS.n4239 VSS.t477 22.6305
R4621 VSS.n4240 VSS.t379 22.6305
R4622 VSS.n4241 VSS.t513 22.6305
R4623 VSS.n4242 VSS.t487 22.6305
R4624 VSS.n4243 VSS.t393 22.6305
R4625 VSS.n4244 VSS.t352 22.6305
R4626 VSS.n4245 VSS.t437 22.6305
R4627 VSS.n4246 VSS.t403 22.6305
R4628 VSS.n4247 VSS.t494 22.6305
R4629 VSS.n4248 VSS.t401 22.6305
R4630 VSS.n1641 VSS.t376 22.6305
R4631 VSS.n1642 VSS.t354 22.6305
R4632 VSS.n1643 VSS.t364 22.6305
R4633 VSS.n1644 VSS.t381 22.6305
R4634 VSS.n1645 VSS.t455 22.6305
R4635 VSS.n1646 VSS.t409 22.6305
R4636 VSS.n1647 VSS.t444 22.6305
R4637 VSS.n1648 VSS.t463 22.6305
R4638 VSS.n1649 VSS.t482 22.6305
R4639 VSS.n1650 VSS.t492 22.6305
R4640 VSS.n1651 VSS.t470 22.6305
R4641 VSS.n1652 VSS.t489 22.6305
R4642 VSS.n7079 VSS.n7078 22.1116
R4643 VSS.n4466 VSS.t909 21.9714
R4644 VSS.n7588 VSS.t155 21.4291
R4645 VSS.n6885 VSS.t131 20.9682
R4646 VSS.t766 VSS.n7247 20.8388
R4647 VSS.n7129 VSS.t263 20.7915
R4648 VSS.n4694 VSS.n4693 20.5962
R4649 VSS.n4147 VSS.n4146 19.6617
R4650 VSS.n719 VSS.t765 19.4363
R4651 VSS.n6898 VSS.n6897 19.3553
R4652 VSS.n239 VSS.n238 19.0342
R4653 VSS.n6026 VSS.t745 18.2305
R4654 VSS.n1084 VSS.n1083 17.1963
R4655 VSS.n5337 VSS.t711 17.1434
R4656 VSS.n5489 VSS.t139 17.0519
R4657 VSS.n11 VSS.t328 16.837
R4658 VSS.n7669 VSS.n7668 16.837
R4659 VSS.n1750 VSS.t456 16.8261
R4660 VSS.n6823 VSS.n6822 16.6245
R4661 VSS.n7252 VSS.n7251 16.2081
R4662 VSS.n6922 VSS.n6921 16.1295
R4663 VSS.n4475 VSS.n4474 15.2111
R4664 VSS.n4491 VSS.t20 15.2111
R4665 VSS.n6196 VSS.t740 15.1921
R4666 VSS.n7473 VSS.n7472 14.6645
R4667 VSS.n6953 VSS.n6952 14.5166
R4668 VSS.n4359 VSS.n4358 13.7634
R4669 VSS.n6495 VSS.t343 13.4581
R4670 VSS.n4238 VSS.n4237 13.4167
R4671 VSS.n4239 VSS.n4238 13.4167
R4672 VSS.n4240 VSS.n4239 13.4167
R4673 VSS.n4241 VSS.n4240 13.4167
R4674 VSS.n4242 VSS.n4241 13.4167
R4675 VSS.n4243 VSS.n4242 13.4167
R4676 VSS.n4244 VSS.n4243 13.4167
R4677 VSS.n4245 VSS.n4244 13.4167
R4678 VSS.n4246 VSS.n4245 13.4167
R4679 VSS.n4247 VSS.n4246 13.4167
R4680 VSS.n1642 VSS.n1641 13.4167
R4681 VSS.n1643 VSS.n1642 13.4167
R4682 VSS.n1644 VSS.n1643 13.4167
R4683 VSS.n1645 VSS.n1644 13.4167
R4684 VSS.n1646 VSS.n1645 13.4167
R4685 VSS.n1647 VSS.n1646 13.4167
R4686 VSS.n1648 VSS.n1647 13.4167
R4687 VSS.n1649 VSS.n1648 13.4167
R4688 VSS.n1650 VSS.n1649 13.4167
R4689 VSS.n1651 VSS.n1650 13.4167
R4690 VSS.n4249 VSS.n4247 13.2852
R4691 VSS.n1653 VSS.n1651 13.2852
R4692 VSS.n5669 VSS.t424 13.1666
R4693 VSS.n5690 VSS.t17 13.1666
R4694 VSS.n6202 VSS.t754 13.1666
R4695 VSS.n7299 VSS.t989 13.0005
R4696 VSS.n6978 VSS.n6610 12.9101
R4697 VSS.n1135 VSS.t329 11.3982
R4698 VSS.n4380 VSS.t1004 11.0483
R4699 VSS.n6750 VSS.t245 10.907
R4700 VSS.n7113 VSS.t829 10.891
R4701 VSS.n4440 VSS.t583 10.3984
R4702 VSS.n4577 VSS.t153 10.315
R4703 VSS.n5556 VSS.t242 10.2313
R4704 VSS.n6100 VSS.t815 10.1283
R4705 VSS.n5240 VSS.t918 10.1024
R4706 VSS.n4297 VSS.t205 9.92633
R4707 VSS.n4406 VSS.t1002 9.74855
R4708 VSS.n322 VSS.n321 9.61182
R4709 VSS.n5720 VSS.t417 9.55913
R4710 VSS.n22 VSS.t446 9.55885
R4711 VSS.n4936 VSS.t501 9.54136
R4712 VSS.n5708 VSS.t468 9.54089
R4713 VSS.n5709 VSS.t359 9.51568
R4714 VSS.n4923 VSS.t434 9.5154
R4715 VSS.n5707 VSS.t510 9.5085
R4716 VSS.n4946 VSS.t373 9.50824
R4717 VSS.n23 VSS.t461 9.49457
R4718 VSS.n5159 VSS.t426 9.49428
R4719 VSS.n5160 VSS.t449 9.49428
R4720 VSS.n5161 VSS.t474 9.49428
R4721 VSS.n5162 VSS.t458 9.49428
R4722 VSS.n5613 VSS.t498 9.49403
R4723 VSS.n5612 VSS.t506 9.49403
R4724 VSS.n5573 VSS.t441 9.49403
R4725 VSS.n5455 VSS.t423 9.49403
R4726 VSS.n5710 VSS.t429 9.49372
R4727 VSS.n5163 VSS.t384 9.45083
R4728 VSS.n5454 VSS.t508 9.45057
R4729 VSS.n5718 VSS.t405 9.43205
R4730 VSS.n5754 VSS.t472 9.43205
R4731 VSS.n5777 VSS.t439 9.43205
R4732 VSS.n5747 VSS.t451 9.43205
R4733 VSS.n5768 VSS.t349 9.43205
R4734 VSS.n4934 VSS.t453 9.43205
R4735 VSS.n4911 VSS.t367 9.43205
R4736 VSS.n4920 VSS.t407 9.43205
R4737 VSS.n4944 VSS.t485 9.43205
R4738 VSS.n4937 VSS.t398 9.43205
R4739 VSS.n5933 VSS.t503 9.3886
R4740 VSS.n5912 VSS.t419 9.3886
R4741 VSS.n4756 VSS.t395 9.3886
R4742 VSS.n4778 VSS.t390 9.3886
R4743 VSS.n5872 VSS.t415 9.34514
R4744 VSS.n5877 VSS.t412 9.34514
R4745 VSS.n5939 VSS.t370 9.34514
R4746 VSS.n4976 VSS.t431 9.34514
R4747 VSS.n50 VSS.t387 9.34514
R4748 VSS.n4760 VSS.t479 9.34514
R4749 VSS.n7135 VSS.t261 9.24095
R4750 VSS.n971 VSS.n969 9.13939
R4751 VSS.n1544 VSS.n1542 9.13939
R4752 VSS.n649 VSS.n647 9.13939
R4753 VSS.n5554 VSS.n5460 9.13939
R4754 VSS.n5558 VSS.n5554 9.13939
R4755 VSS.n5482 VSS.n5466 9.13939
R4756 VSS.n5484 VSS.n5482 9.13939
R4757 VSS.n5520 VSS.n5503 9.13939
R4758 VSS.n5522 VSS.n5520 9.13939
R4759 VSS.n5595 VSS.n5578 9.13939
R4760 VSS.n5597 VSS.n5595 9.13939
R4761 VSS.n6788 VSS.n6786 9.13939
R4762 VSS.n7591 VSS.n7589 9.13939
R4763 VSS.n6444 VSS.n6442 9.13939
R4764 VSS.n7819 VSS.n5230 9.13939
R4765 VSS.n7819 VSS.n7817 9.13939
R4766 VSS.n7821 VSS.n7820 9.13939
R4767 VSS.n7820 VSS.n5231 9.13939
R4768 VSS.n7794 VSS.n7793 9.02001
R4769 VSS.n0 VSS.t332 8.97995
R4770 VSS.n5233 VSS.t841 8.89703
R4771 VSS.n5237 VSS.n5236 8.78137
R4772 VSS.n5238 VSS.t923 8.5505
R4773 VSS.n5239 VSS.t922 8.5505
R4774 VSS.n5233 VSS.t842 8.5505
R4775 VSS.n1135 VSS.n1134 8.5505
R4776 VSS.n6794 VSS.n6793 8.31252
R4777 VSS.t475 VSS.t459 8.24923
R4778 VSS.n4545 VSS.n4543 8.16717
R4779 VSS.n6751 VSS.n6750 8.16341
R4780 VSS.n7204 VSS.t85 7.92089
R4781 VSS.n1552 VSS.n1550 7.58383
R4782 VSS.n6978 VSS.n6977 7.54047
R4783 VSS.n763 VSS.n762 7.50194
R4784 VSS.n640 VSS.n638 7.48661
R4785 VSS.t939 VSS.t31 7.40369
R4786 VSS.t839 VSS.t32 7.40369
R4787 VSS.n4302 VSS.t173 7.09038
R4788 VSS.n5663 VSS.n5662 7.08994
R4789 VSS.n6129 VSS.t16 7.08994
R4790 VSS.n6981 VSS.n6595 6.8902
R4791 VSS.n6982 VSS.n6594 6.87063
R4792 VSS.n1466 VSS.n1465 6.76077
R4793 VSS.n6977 VSS.t577 6.68867
R4794 VSS.n6610 VSS.t996 6.68867
R4795 VSS.n730 VSS.n729 6.65541
R4796 VSS.n754 VSS.t235 6.65541
R4797 VSS.n607 VSS.n600 6.65541
R4798 VSS.n607 VSS.n601 6.65541
R4799 VSS.n673 VSS.t340 6.65541
R4800 VSS.n673 VSS.t934 6.65541
R4801 VSS.n5533 VSS.t140 6.65541
R4802 VSS.n5508 VSS.n5504 6.65541
R4803 VSS.n5470 VSS.n5467 6.65541
R4804 VSS.n5495 VSS.t55 6.65541
R4805 VSS.n5542 VSS.n5461 6.65541
R4806 VSS.n5569 VSS.t241 6.65541
R4807 VSS.n5608 VSS.t348 6.65541
R4808 VSS.n5583 VSS.n5579 6.65541
R4809 VSS.n6419 VSS.t905 6.65541
R4810 VSS.n6458 VSS.n6437 6.65541
R4811 VSS.n7082 VSS.n7077 6.65541
R4812 VSS.n7182 VSS.t946 6.65541
R4813 VSS.n7835 VSS.n5222 6.65541
R4814 VSS.n7835 VSS.n5223 6.65541
R4815 VSS.n7802 VSS.t307 6.65541
R4816 VSS.n7802 VSS.t546 6.65541
R4817 VSS.n7577 VSS.t160 6.65541
R4818 VSS.n7605 VSS.n5319 6.65541
R4819 VSS.n6774 VSS.t823 6.65541
R4820 VSS.n6803 VSS.n6640 6.65541
R4821 VSS.n1509 VSS.n1502 6.65541
R4822 VSS.n1509 VSS.n1503 6.65541
R4823 VSS.n1566 VSS.t880 6.65541
R4824 VSS.n1566 VSS.t1001 6.65541
R4825 VSS.n4587 VSS.t80 6.65541
R4826 VSS.n4527 VSS.n697 6.65541
R4827 VSS.n1489 VSS.t1005 6.65541
R4828 VSS.n4370 VSS.n1608 6.65541
R4829 VSS.n951 VSS.t276 6.65541
R4830 VSS.n985 VSS.n964 6.65541
R4831 VSS.n5719 VSS.t406 6.63905
R4832 VSS.n4913 VSS.t369 6.63905
R4833 VSS.n5913 VSS.t420 6.63522
R4834 VSS.n5934 VSS.t505 6.63522
R4835 VSS.n4757 VSS.t397 6.63522
R4836 VSS.n4779 VSS.t392 6.63522
R4837 VSS.n5940 VSS.t372 6.63331
R4838 VSS.n4761 VSS.t481 6.63331
R4839 VSS.n6599 VSS.t560 6.62607
R4840 VSS.n6607 VSS.t557 6.62607
R4841 VSS.n6600 VSS.n6596 6.6202
R4842 VSS.n6608 VSS.n6604 6.6202
R4843 VSS.n4977 VSS.t433 6.5299
R4844 VSS.n5873 VSS.t416 6.5165
R4845 VSS.n5878 VSS.t414 6.50525
R4846 VSS.n51 VSS.t389 6.50525
R4847 VSS.n6953 VSS.n6951 6.45211
R4848 VSS.n7537 VSS.t121 6.45211
R4849 VSS.n5930 VSS.t739 6.4265
R4850 VSS.n5874 VSS.t983 6.4265
R4851 VSS.n5869 VSS.t805 6.4265
R4852 VSS.n5767 VSS.t440 6.4265
R4853 VSS.n5449 VSS.n5444 6.4265
R4854 VSS.n5740 VSS.t452 6.4265
R4855 VSS.n5749 VSS.t473 6.4265
R4856 VSS.n5451 VSS.n5443 6.4265
R4857 VSS.n5742 VSS.n5741 6.4265
R4858 VSS.n5769 VSS.t351 6.4265
R4859 VSS.n6602 VSS.n6601 6.4265
R4860 VSS.n6609 VSS.n6603 6.4265
R4861 VSS.n4927 VSS.t801 6.4265
R4862 VSS.n4929 VSS.t864 6.4265
R4863 VSS.n4906 VSS.t796 6.4265
R4864 VSS.n4921 VSS.t454 6.4265
R4865 VSS.n4912 VSS.t408 6.4265
R4866 VSS.n4924 VSS.t486 6.4265
R4867 VSS.n4938 VSS.t400 6.4265
R4868 VSS.n4745 VSS.n4744 6.4265
R4869 VSS.n4975 VSS.n4974 6.4265
R4870 VSS.n47 VSS.n46 6.4265
R4871 VSS.n7302 VSS.n7301 6.33064
R4872 VSS.n1753 VSS.t464 6.19941
R4873 VSS.n5156 VSS.t899 6.17387
R4874 VSS.n4512 VSS.n4511 5.91574
R4875 VSS.n1261 VSS.n1260 5.84933
R4876 VSS.n7142 VSS.n7141 5.81586
R4877 VSS.n219 VSS.n216 5.80511
R4878 VSS.n4128 VSS.n4127 5.76287
R4879 VSS.n355 VSS.n354 5.60395
R4880 VSS.n5235 VSS.n5234 5.4005
R4881 VSS.n5235 VSS.t925 5.4005
R4882 VSS.n7890 VSS.n7889 5.4005
R4883 VSS.n7890 VSS.t331 5.4005
R4884 VSS.n4287 VSS.n4285 5.38343
R4885 VSS.n1733 VSS.n1731 5.38343
R4886 VSS.n167 VSS.n166 5.26318
R4887 VSS.n5265 VSS.n5264 5.24323
R4888 VSS.n758 VSS.n757 5.2005
R4889 VSS.n760 VSS.n759 5.2005
R4890 VSS.n6415 VSS.n6412 5.2005
R4891 VSS.n6414 VSS.n6413 5.2005
R4892 VSS.n6410 VSS.n6394 5.2005
R4893 VSS.n6409 VSS.n6408 5.2005
R4894 VSS.n6408 VSS.n6407 5.2005
R4895 VSS.n6406 VSS.n6405 5.2005
R4896 VSS.n6405 VSS.n6404 5.2005
R4897 VSS.n6486 VSS.n6485 5.2005
R4898 VSS.n6484 VSS.n6483 5.2005
R4899 VSS.n6432 VSS.n6431 5.2005
R4900 VSS.n6434 VSS.n6433 5.2005
R4901 VSS VSS.n7299 5.2005
R4902 VSS.n7842 VSS.n7841 5.2005
R4903 VSS.n5348 VSS.n5347 5.2005
R4904 VSS.n5350 VSS.n5349 5.2005
R4905 VSS.n6944 VSS.n6943 5.2005
R4906 VSS.n6950 VSS.n6949 5.2005
R4907 VSS.n6951 VSS.n6950 5.2005
R4908 VSS.n7243 VSS.n7242 5.2005
R4909 VSS.n7235 VSS.n7234 5.2005
R4910 VSS.n7232 VSS.n7229 5.2005
R4911 VSS.n7231 VSS.n7230 5.2005
R4912 VSS.n7245 VSS.n7244 5.2005
R4913 VSS.n7178 VSS.n7096 5.2005
R4914 VSS.n7177 VSS.n7097 5.2005
R4915 VSS.n7175 VSS.n7120 5.2005
R4916 VSS.n7174 VSS.n7173 5.2005
R4917 VSS.n7173 VSS.n7172 5.2005
R4918 VSS.n7171 VSS.n7170 5.2005
R4919 VSS.n7170 VSS.n7169 5.2005
R4920 VSS.n7616 VSS.n7615 5.2005
R4921 VSS.n7615 VSS.n7614 5.2005
R4922 VSS.n7613 VSS.n7612 5.2005
R4923 VSS.n7612 VSS.n7611 5.2005
R4924 VSS.n7610 VSS.n5307 5.2005
R4925 VSS.n7608 VSS.n5315 5.2005
R4926 VSS.n7607 VSS.n5316 5.2005
R4927 VSS.n6682 VSS.n6681 5.2005
R4928 VSS.n6684 VSS.n6683 5.2005
R4929 VSS.n6742 VSS.n6741 5.2005
R4930 VSS.n6738 VSS.n6737 5.2005
R4931 VSS.n6740 VSS.n6739 5.2005
R4932 VSS.n6630 VSS.n6629 5.2005
R4933 VSS.n6629 VSS.n6628 5.2005
R4934 VSS.n6633 VSS.n6632 5.2005
R4935 VSS.n6632 VSS.n6631 5.2005
R4936 VSS.n6635 VSS.n6634 5.2005
R4937 VSS.n6806 VSS.n6636 5.2005
R4938 VSS.n6805 VSS.n6637 5.2005
R4939 VSS.n183 VSS.n182 5.2005
R4940 VSS.n182 VSS.n181 5.2005
R4941 VSS.n186 VSS.n185 5.2005
R4942 VSS.n185 VSS.n184 5.2005
R4943 VSS.n190 VSS.n188 5.2005
R4944 VSS.n190 VSS.n189 5.2005
R4945 VSS.n175 VSS.n174 5.2005
R4946 VSS.n280 VSS.n279 5.2005
R4947 VSS.n640 VSS.n630 5.2005
R4948 VSS.n640 VSS.n639 5.2005
R4949 VSS.n139 VSS.n138 5.2005
R4950 VSS.n86 VSS.n85 5.2005
R4951 VSS.n85 VSS.n84 5.2005
R4952 VSS.n89 VSS.n88 5.2005
R4953 VSS.n88 VSS.n87 5.2005
R4954 VSS.n157 VSS.n156 5.2005
R4955 VSS.n4545 VSS.n4544 5.2005
R4956 VSS.n4567 VSS.n4566 5.2005
R4957 VSS.n4580 VSS.n4579 5.2005
R4958 VSS.n4607 VSS.n4606 5.2005
R4959 VSS.n4606 VSS.n4605 5.2005
R4960 VSS.n4604 VSS.n4603 5.2005
R4961 VSS.n4603 VSS.n4602 5.2005
R4962 VSS.n4523 VSS.n4522 5.2005
R4963 VSS.n4287 VSS.n4286 5.2005
R4964 VSS.n4289 VSS.n4288 5.2005
R4965 VSS.n4292 VSS.n4291 5.2005
R4966 VSS.n4294 VSS.n4293 5.2005
R4967 VSS.n4296 VSS.n4295 5.2005
R4968 VSS.n4298 VSS.n4297 5.2005
R4969 VSS.n4300 VSS.n4299 5.2005
R4970 VSS.n4303 VSS.n4302 5.2005
R4971 VSS.n4305 VSS.n4304 5.2005
R4972 VSS.n4306 VSS 5.2005
R4973 VSS.n4308 VSS.n4307 5.2005
R4974 VSS.n4311 VSS.n4310 5.2005
R4975 VSS.n4313 VSS.n4312 5.2005
R4976 VSS.n4316 VSS.n4315 5.2005
R4977 VSS.n4318 VSS.n4317 5.2005
R4978 VSS.n4321 VSS.n4320 5.2005
R4979 VSS.n4335 VSS.n4334 5.2005
R4980 VSS.n4337 VSS.n4336 5.2005
R4981 VSS.n4339 VSS.n4338 5.2005
R4982 VSS.n1733 VSS.n1732 5.2005
R4983 VSS.n1735 VSS.n1734 5.2005
R4984 VSS.n1749 VSS.n1748 5.2005
R4985 VSS.n1751 VSS.n1750 5.2005
R4986 VSS.n1755 VSS.n1754 5.2005
R4987 VSS.n1755 VSS.n1753 5.2005
R4988 VSS.n1688 VSS.n1687 5.2005
R4989 VSS.n1691 VSS.n1690 5.2005
R4990 VSS.n1727 VSS.n1726 5.2005
R4991 VSS.n1725 VSS 5.2005
R4992 VSS.n1724 VSS.n1693 5.2005
R4993 VSS.n1716 VSS.n1694 5.2005
R4994 VSS.n1715 VSS.n1695 5.2005
R4995 VSS.n1632 VSS.n1631 5.2005
R4996 VSS.n1713 VSS.n1712 5.2005
R4997 VSS.n1623 VSS.n1622 5.2005
R4998 VSS.n1626 VSS.n1625 5.2005
R4999 VSS.n1630 VSS.n1629 5.2005
R5000 VSS.n1630 VSS.n1628 5.2005
R5001 VSS.n4411 VSS.n4410 5.2005
R5002 VSS.n4405 VSS.n4404 5.2005
R5003 VSS.n4404 VSS.n4403 5.2005
R5004 VSS.n4387 VSS.n4386 5.2005
R5005 VSS.n1600 VSS.n1599 5.2005
R5006 VSS.n1550 VSS.n1549 5.2005
R5007 VSS.n1479 VSS.n1478 5.2005
R5008 VSS.n4511 VSS.n4510 5.2005
R5009 VSS.n4509 VSS.n723 5.2005
R5010 VSS.n1481 VSS.n1480 5.2005
R5011 VSS.n720 VSS.n719 5.2005
R5012 VSS.n4518 VSS.n4517 5.2005
R5013 VSS.n4521 VSS.n4520 5.2005
R5014 VSS.n722 VSS.n721 5.2005
R5015 VSS.n766 VSS.n765 5.2005
R5016 VSS.n770 VSS.n769 5.2005
R5017 VSS.n4592 VSS.n4591 5.2005
R5018 VSS.n4594 VSS.n4593 5.2005
R5019 VSS.n4596 VSS.n4595 5.2005
R5020 VSS.n5241 VSS.n5240 5.2005
R5021 VSS.n5258 VSS.n5257 5.2005
R5022 VSS.n5261 VSS.n5260 5.2005
R5023 VSS.n5263 VSS.n5262 5.2005
R5024 VSS.n947 VSS.n944 5.2005
R5025 VSS.n946 VSS.n945 5.2005
R5026 VSS.n942 VSS.n926 5.2005
R5027 VSS.n941 VSS.n940 5.2005
R5028 VSS.n940 VSS.n939 5.2005
R5029 VSS.n938 VSS.n937 5.2005
R5030 VSS.n937 VSS.n936 5.2005
R5031 VSS.n995 VSS.n994 5.2005
R5032 VSS.n994 VSS.n993 5.2005
R5033 VSS.n998 VSS.n997 5.2005
R5034 VSS.n997 VSS.n996 5.2005
R5035 VSS.n1004 VSS.n1003 5.2005
R5036 VSS.n1002 VSS.n1001 5.2005
R5037 VSS.n1000 VSS.n999 5.2005
R5038 VSS.n1138 VSS.n1137 5.2005
R5039 VSS.n21 VSS.n20 5.2005
R5040 VSS.n7888 VSS.n7887 5.2005
R5041 VSS.n7893 VSS.n7892 5.2005
R5042 VSS.n1 VSS.n0 5.2005
R5043 VSS VSS.n2 5.2005
R5044 VSS.n7909 VSS.n11 5.2005
R5045 VSS.n13 VSS.n12 5.2005
R5046 VSS.n4894 VSS.t970 5.1234
R5047 VSS.n6173 VSS.n6172 5.12337
R5048 VSS.n4893 VSS.t863 5.12337
R5049 VSS.n4775 VSS.n4773 5.12334
R5050 VSS.n5929 VSS.t723 5.12332
R5051 VSS.n5447 VSS.n5445 5.12328
R5052 VSS.n5895 VSS.t954 5.12118
R5053 VSS.n4748 VSS.n4747 5.12105
R5054 VSS.n4256 VSS.n4253 5.11535
R5055 VSS.n1658 VSS.n1655 5.11535
R5056 VSS.n7144 VSS.t826 5.10208
R5057 VSS.n7147 VSS.t262 5.10194
R5058 VSS.n7143 VSS.t39 5.08021
R5059 VSS.n7092 VSS.t824 4.95074
R5060 VSS.n4477 VSS.n1477 4.88533
R5061 VSS.n7226 VSS.n7225 4.88533
R5062 VSS.n83 VSS.n80 4.88449
R5063 VSS.n6492 VSS.n6488 4.88319
R5064 VSS.n992 VSS.n989 4.88319
R5065 VSS.n180 VSS.n177 4.88277
R5066 VSS.n4601 VSS.n4598 4.88215
R5067 VSS.n6747 VSS.n6746 4.88215
R5068 VSS.n6947 VSS.n6946 4.88215
R5069 VSS.n4566 VSS.t82 4.6889
R5070 VSS.n7147 VSS.n7146 4.66114
R5071 VSS.n2354 VSS.n2331 4.50764
R5072 VSS.n2468 VSS.n2467 4.50764
R5073 VSS.n3026 VSS.n3025 4.50622
R5074 VSS.n2944 VSS.n2943 4.50622
R5075 VSS.n2875 VSS.n2874 4.50622
R5076 VSS.n2725 VSS.n2724 4.50565
R5077 VSS.n2238 VSS.n2236 4.50554
R5078 VSS.n2729 VSS.n2728 4.50495
R5079 VSS.n2810 VSS.n2809 4.50484
R5080 VSS.n2660 VSS.n2659 4.5026
R5081 VSS.n2660 VSS.n2656 4.50224
R5082 VSS.n3027 VSS.n3026 4.50095
R5083 VSS.n2946 VSS.n2238 4.50095
R5084 VSS.n2945 VSS.n2944 4.50095
R5085 VSS.n2877 VSS.n2331 4.50095
R5086 VSS.n2876 VSS.n2875 4.50095
R5087 VSS.n2812 VSS.n2468 4.50095
R5088 VSS.n2726 VSS.n2725 4.50089
R5089 VSS.n2811 VSS.n2810 4.50089
R5090 VSS.n2728 VSS.n2727 4.50089
R5091 VSS.n2146 VSS.n2141 4.5005
R5092 VSS.n2156 VSS.n2149 4.5005
R5093 VSS.n3008 VSS.n3007 4.5005
R5094 VSS.n2157 VSS.n2150 4.5005
R5095 VSS.n2951 VSS.n2950 4.5005
R5096 VSS.n2953 VSS.n2952 4.5005
R5097 VSS.n2206 VSS.n2205 4.5005
R5098 VSS.n2982 VSS.n2981 4.5005
R5099 VSS.n2994 VSS.n2993 4.5005
R5100 VSS.n3023 VSS.n3022 4.5005
R5101 VSS.n2969 VSS.n2968 4.5005
R5102 VSS.n2224 VSS.n2215 4.5005
R5103 VSS.n2225 VSS.n2222 4.5005
R5104 VSS.n2967 VSS.n2966 4.5005
R5105 VSS.n2204 VSS.n2203 4.5005
R5106 VSS.n2173 VSS.n2162 4.5005
R5107 VSS.n3006 VSS.n3005 4.5005
R5108 VSS.n2996 VSS.n2995 4.5005
R5109 VSS.n2998 VSS.n2997 4.5005
R5110 VSS.n2181 VSS.n2180 4.5005
R5111 VSS.n2145 VSS.n2142 4.5005
R5112 VSS.n2159 VSS.n2152 4.5005
R5113 VSS.n3012 VSS.n3011 4.5005
R5114 VSS.n3021 VSS.n3020 4.5005
R5115 VSS.n2176 VSS.n2172 4.5005
R5116 VSS.n2980 VSS.n2979 4.5005
R5117 VSS.n2965 VSS.n2964 4.5005
R5118 VSS.n2240 VSS.n2223 4.5005
R5119 VSS.n2971 VSS.n2970 4.5005
R5120 VSS.n2221 VSS.n2217 4.5005
R5121 VSS.n2237 VSS.n2235 4.5005
R5122 VSS.n2955 VSS.n2954 4.5005
R5123 VSS.n2986 VSS.n2985 4.5005
R5124 VSS.n2171 VSS.n2164 4.5005
R5125 VSS.n2163 VSS.n2161 4.5005
R5126 VSS.n2201 VSS.n2199 4.5005
R5127 VSS.n2207 VSS.n2202 4.5005
R5128 VSS.n3014 VSS.n3013 4.5005
R5129 VSS.n2941 VSS.n2940 4.5005
R5130 VSS.n2332 VSS.n2329 4.5005
R5131 VSS.n2287 VSS.n2286 4.5005
R5132 VSS.n2339 VSS.n2335 4.5005
R5133 VSS.n2284 VSS.n2259 4.5005
R5134 VSS.n2290 VSS.n2271 4.5005
R5135 VSS.n2253 VSS.n2248 4.5005
R5136 VSS.n2347 VSS.n2346 4.5005
R5137 VSS.n2345 VSS.n2328 4.5005
R5138 VSS.n2289 VSS.n2270 4.5005
R5139 VSS.n2341 VSS.n2340 4.5005
R5140 VSS.n2350 VSS.n2349 4.5005
R5141 VSS.n2334 VSS.n2316 4.5005
R5142 VSS.n2927 VSS.n2256 4.5005
R5143 VSS.n2315 VSS.n2282 4.5005
R5144 VSS.n2929 VSS.n2928 4.5005
R5145 VSS.n2931 VSS.n2930 4.5005
R5146 VSS.n2285 VSS.n2267 4.5005
R5147 VSS.n2898 VSS.n2897 4.5005
R5148 VSS.n2909 VSS.n2908 4.5005
R5149 VSS.n2266 VSS.n2261 4.5005
R5150 VSS.n2918 VSS.n2917 4.5005
R5151 VSS.n2896 VSS.n2895 4.5005
R5152 VSS.n2348 VSS.n2325 4.5005
R5153 VSS.n2916 VSS.n2915 4.5005
R5154 VSS.n2260 VSS.n2255 4.5005
R5155 VSS.n2337 VSS.n2336 4.5005
R5156 VSS.n2277 VSS.n2273 4.5005
R5157 VSS.n2298 VSS.n2295 4.5005
R5158 VSS.n2881 VSS.n2880 4.5005
R5159 VSS.n2252 VSS.n2249 4.5005
R5160 VSS.n2296 VSS.n2281 4.5005
R5161 VSS.n2884 VSS.n2883 4.5005
R5162 VSS.n2882 VSS.n2327 4.5005
R5163 VSS.n2338 VSS.n2321 4.5005
R5164 VSS.n2939 VSS.n2938 4.5005
R5165 VSS.n2369 VSS.n2364 4.5005
R5166 VSS.n2405 VSS.n2372 4.5005
R5167 VSS.n2453 VSS.n2438 4.5005
R5168 VSS.n2402 VSS.n2398 4.5005
R5169 VSS.n2409 VSS.n2408 4.5005
R5170 VSS.n2839 VSS.n2838 4.5005
R5171 VSS.n2456 VSS.n2455 4.5005
R5172 VSS.n2461 VSS.n2458 4.5005
R5173 VSS.n2417 VSS.n2416 4.5005
R5174 VSS.n2401 VSS.n2400 4.5005
R5175 VSS.n2872 VSS.n2871 4.5005
R5176 VSS.n2383 VSS.n2381 4.5005
R5177 VSS.n2463 VSS.n2462 4.5005
R5178 VSS.n2406 VSS.n2373 4.5005
R5179 VSS.n2852 VSS.n2851 4.5005
R5180 VSS.n2452 VSS.n2437 4.5005
R5181 VSS.n2450 VSS.n2449 4.5005
R5182 VSS.n2850 VSS.n2849 4.5005
R5183 VSS.n2387 VSS.n2385 4.5005
R5184 VSS.n2840 VSS.n2397 4.5005
R5185 VSS.n2368 VSS.n2365 4.5005
R5186 VSS.n2460 VSS.n2447 4.5005
R5187 VSS.n2828 VSS.n2827 4.5005
R5188 VSS.n2436 VSS.n2420 4.5005
R5189 VSS.n2854 VSS.n2853 4.5005
R5190 VSS.n2861 VSS.n2860 4.5005
R5191 VSS.n2459 VSS.n2445 4.5005
R5192 VSS.n2870 VSS.n2869 4.5005
R5193 VSS.n2396 VSS.n2386 4.5005
R5194 VSS.n2817 VSS.n2816 4.5005
R5195 VSS.n2830 VSS.n2829 4.5005
R5196 VSS.n2842 VSS.n2841 4.5005
R5197 VSS.n2407 VSS.n2375 4.5005
R5198 VSS.n2391 VSS.n2382 4.5005
R5199 VSS.n2454 VSS.n2440 4.5005
R5200 VSS.n2863 VSS.n2862 4.5005
R5201 VSS.n2480 VSS.n2473 4.5005
R5202 VSS.n2795 VSS.n2794 4.5005
R5203 VSS.n2745 VSS.n2744 4.5005
R5204 VSS.n2781 VSS.n2780 4.5005
R5205 VSS.n2783 VSS.n2782 4.5005
R5206 VSS.n2495 VSS.n2484 4.5005
R5207 VSS.n2770 VSS.n2769 4.5005
R5208 VSS.n2526 VSS.n2524 4.5005
R5209 VSS.n2732 VSS.n2731 4.5005
R5210 VSS.n2502 VSS.n2500 4.5005
R5211 VSS.n2807 VSS.n2806 4.5005
R5212 VSS.n2793 VSS.n2482 4.5005
R5213 VSS.n2497 VSS.n2496 4.5005
R5214 VSS.n2755 VSS.n2754 4.5005
R5215 VSS.n2743 VSS.n2742 4.5005
R5216 VSS.n2768 VSS.n2515 4.5005
R5217 VSS.n2560 VSS.n2559 4.5005
R5218 VSS.n2547 VSS.n2546 4.5005
R5219 VSS.n2516 VSS.n2514 4.5005
R5220 VSS.n2757 VSS.n2756 4.5005
R5221 VSS.n2805 VSS.n2804 4.5005
R5222 VSS.n2759 VSS.n2758 4.5005
R5223 VSS.n2558 VSS.n2555 4.5005
R5224 VSS.n2508 VSS.n2501 4.5005
R5225 VSS.n2476 VSS.n2474 4.5005
R5226 VSS.n2499 VSS.n2493 4.5005
R5227 VSS.n2491 VSS.n2487 4.5005
R5228 VSS.n2753 VSS.n2752 4.5005
R5229 VSS.n2565 VSS.n2562 4.5005
R5230 VSS.n2544 VSS.n2529 4.5005
R5231 VSS.n2527 VSS.n2525 4.5005
R5232 VSS.n2741 VSS.n2740 4.5005
R5233 VSS.n2734 VSS.n2733 4.5005
R5234 VSS.n2548 VSS.n2545 4.5005
R5235 VSS.n2494 VSS.n2492 4.5005
R5236 VSS.n2779 VSS.n2778 4.5005
R5237 VSS.n2486 VSS.n2479 4.5005
R5238 VSS.n2797 VSS.n2796 4.5005
R5239 VSS.n2692 VSS.n2691 4.5005
R5240 VSS.n2682 VSS.n2681 4.5005
R5241 VSS.n2591 VSS.n2590 4.5005
R5242 VSS.n2722 VSS.n2721 4.5005
R5243 VSS.n2600 VSS.n2593 4.5005
R5244 VSS.n2649 VSS.n2605 4.5005
R5245 VSS.n2695 VSS.n2694 4.5005
R5246 VSS.n2659 VSS.n2658 4.5005
R5247 VSS.n2619 VSS.n2617 4.5005
R5248 VSS.n2616 VSS.n2614 4.5005
R5249 VSS.n2680 VSS.n2679 4.5005
R5250 VSS.n2654 VSS.n2653 4.5005
R5251 VSS.n2720 VSS.n2577 4.5005
R5252 VSS.n2647 VSS.n2645 4.5005
R5253 VSS.n2644 VSS.n2621 4.5005
R5254 VSS.n2606 VSS.n2604 4.5005
R5255 VSS.n2587 VSS.n2585 4.5005
R5256 VSS.n2580 VSS.n2578 4.5005
R5257 VSS.n2678 VSS.n2677 4.5005
R5258 VSS.n2662 VSS.n2661 4.5005
R5259 VSS.n2598 VSS.n2594 4.5005
R5260 VSS.n2657 VSS.n2655 4.5005
R5261 VSS.n2638 VSS.n2618 4.5005
R5262 VSS.n2719 VSS.n2718 4.5005
R5263 VSS.n2611 VSS.n2607 4.5005
R5264 VSS.n2684 VSS.n2683 4.5005
R5265 VSS.n2697 VSS.n2696 4.5005
R5266 VSS.n2634 VSS.n2615 4.5005
R5267 VSS.n2609 VSS.n2608 4.5005
R5268 VSS.n2637 VSS.n2636 4.5005
R5269 VSS.n2714 VSS.n2713 4.5005
R5270 VSS.n2583 VSS.n2582 4.5005
R5271 VSS.n2717 VSS.n2716 4.5005
R5272 VSS.n2635 VSS.n2613 4.5005
R5273 VSS.n2699 VSS.n2698 4.5005
R5274 VSS.n2641 VSS.n2620 4.5005
R5275 VSS.n2687 VSS.n2686 4.5005
R5276 VSS.n2700 VSS.n2595 4.5005
R5277 VSS.n2640 VSS.n2639 4.5005
R5278 VSS.n2664 VSS.n2663 4.5005
R5279 VSS.n2676 VSS.n2675 4.5005
R5280 VSS.n2735 VSS.n2563 4.5005
R5281 VSS.n2739 VSS.n2738 4.5005
R5282 VSS.n2552 VSS.n2543 4.5005
R5283 VSS.n2511 VSS.n2503 4.5005
R5284 VSS.n2530 VSS.n2528 4.5005
R5285 VSS.n2787 VSS.n2786 4.5005
R5286 VSS.n2760 VSS.n2542 4.5005
R5287 VSS.n2513 VSS.n2512 4.5005
R5288 VSS.n2488 VSS.n2478 4.5005
R5289 VSS.n2801 VSS.n2475 4.5005
R5290 VSS.n2507 VSS.n2506 4.5005
R5291 VSS.n2553 VSS.n2549 4.5005
R5292 VSS.n2762 VSS.n2761 4.5005
R5293 VSS.n2774 VSS.n2773 4.5005
R5294 VSS.n2737 VSS.n2736 4.5005
R5295 VSS.n2788 VSS.n2489 4.5005
R5296 VSS.n2510 VSS.n2509 4.5005
R5297 VSS.n2561 VSS.n2554 4.5005
R5298 VSS.n2799 VSS.n2798 4.5005
R5299 VSS.n2803 VSS.n2802 4.5005
R5300 VSS.n2868 VSS.n2867 4.5005
R5301 VSS.n2389 VSS.n2380 4.5005
R5302 VSS.n2376 VSS.n2374 4.5005
R5303 VSS.n2866 VSS.n2366 4.5005
R5304 VSS.n2394 VSS.n2393 4.5005
R5305 VSS.n2859 VSS.n2858 4.5005
R5306 VSS.n2826 VSS.n2825 4.5005
R5307 VSS.n2441 VSS.n2439 4.5005
R5308 VSS.n2819 VSS.n2818 4.5005
R5309 VSS.n2821 VSS.n2820 4.5005
R5310 VSS.n2832 VSS.n2831 4.5005
R5311 VSS.n2845 VSS.n2388 4.5005
R5312 VSS.n2392 VSS.n2390 4.5005
R5313 VSS.n2435 VSS.n2434 4.5005
R5314 VSS.n2844 VSS.n2843 4.5005
R5315 VSS.n2371 VSS.n2367 4.5005
R5316 VSS.n2418 VSS.n2395 4.5005
R5317 VSS.n2448 VSS.n2446 4.5005
R5318 VSS.n2935 VSS.n2250 4.5005
R5319 VSS.n2264 VSS.n2262 4.5005
R5320 VSS.n2319 VSS.n2317 4.5005
R5321 VSS.n2311 VSS.n2297 4.5005
R5322 VSS.n2275 VSS.n2272 4.5005
R5323 VSS.n2359 VSS.n2330 4.5005
R5324 VSS.n2932 VSS.n2251 4.5005
R5325 VSS.n2922 VSS.n2263 4.5005
R5326 VSS.n2910 VSS.n2276 4.5005
R5327 VSS.n2892 VSS.n2318 4.5005
R5328 VSS.n2914 VSS.n2913 4.5005
R5329 VSS.n2900 VSS.n2899 4.5005
R5330 VSS.n2886 VSS.n2885 4.5005
R5331 VSS.n2356 VSS.n2326 4.5005
R5332 VSS.n2894 VSS.n2893 4.5005
R5333 VSS.n2274 VSS.n2269 4.5005
R5334 VSS.n2314 VSS.n2313 4.5005
R5335 VSS.n2937 VSS.n2936 4.5005
R5336 VSS.n2921 VSS.n2920 4.5005
R5337 VSS.n2358 VSS.n2357 4.5005
R5338 VSS.n2210 VSS.n2200 4.5005
R5339 VSS.n2220 VSS.n2219 4.5005
R5340 VSS.n2988 VSS.n2987 4.5005
R5341 VSS.n2974 VSS.n2973 4.5005
R5342 VSS.n3017 VSS.n2143 4.5005
R5343 VSS.n2148 VSS.n2144 4.5005
R5344 VSS.n2999 VSS.n2169 4.5005
R5345 VSS.n2185 VSS.n2179 4.5005
R5346 VSS.n2166 VSS.n2165 4.5005
R5347 VSS.n2153 VSS.n2151 4.5005
R5348 VSS.n2178 VSS.n2170 4.5005
R5349 VSS.n2978 VSS.n2977 4.5005
R5350 VSS.n2241 VSS.n2239 4.5005
R5351 VSS.n2211 VSS.n2208 4.5005
R5352 VSS.n2243 VSS.n2242 4.5005
R5353 VSS.n2972 VSS.n2198 4.5005
R5354 VSS.n2957 VSS.n2956 4.5005
R5355 VSS.n3019 VSS.n3018 4.5005
R5356 VSS.n3001 VSS.n3000 4.5005
R5357 VSS.n2168 VSS.n2167 4.5005
R5358 VSS.n6403 VSS.n6402 4.5005
R5359 VSS.n6402 VSS.n6401 4.5005
R5360 VSS.n6493 VSS.n6492 4.5005
R5361 VSS.n6494 VSS.n6493 4.5005
R5362 VSS.n7840 VSS.n7839 4.5005
R5363 VSS.n6941 VSS.n6940 4.5005
R5364 VSS.n7247 VSS.n7246 4.5005
R5365 VSS.n7168 VSS.n7167 4.5005
R5366 VSS.n7167 VSS.n7166 4.5005
R5367 VSS.n7619 VSS.n7618 4.5005
R5368 VSS.n7618 VSS.n7617 4.5005
R5369 VSS.n6748 VSS.n6747 4.5005
R5370 VSS.n6749 VSS.n6748 4.5005
R5371 VSS.n6627 VSS.n6626 4.5005
R5372 VSS.n6626 VSS.n6625 4.5005
R5373 VSS.n193 VSS.n192 4.5005
R5374 VSS.n192 VSS.n191 4.5005
R5375 VSS.n282 VSS.n281 4.5005
R5376 VSS.n180 VSS.n179 4.5005
R5377 VSS.n179 VSS.n178 4.5005
R5378 VSS.n643 VSS.n636 4.5005
R5379 VSS.n643 VSS.n642 4.5005
R5380 VSS.n83 VSS.n82 4.5005
R5381 VSS.n82 VSS.n81 4.5005
R5382 VSS.n154 VSS.n153 4.5005
R5383 VSS.n153 VSS.n152 4.5005
R5384 VSS.n222 VSS.n221 4.5005
R5385 VSS.n221 VSS.n220 4.5005
R5386 VSS.n4538 VSS.n4537 4.5005
R5387 VSS.n4578 VSS.n4577 4.5005
R5388 VSS.n4601 VSS.n4600 4.5005
R5389 VSS.n4600 VSS.n4599 4.5005
R5390 VSS.n1603 VSS.n1602 4.5005
R5391 VSS.n4400 VSS.n4397 4.5005
R5392 VSS.n4400 VSS.n4399 4.5005
R5393 VSS.n4390 VSS.n4389 4.5005
R5394 VSS.n1500 VSS.n1499 4.5005
R5395 VSS.n4477 VSS.n4476 4.5005
R5396 VSS.n4476 VSS.n4475 4.5005
R5397 VSS.n4514 VSS.n4513 4.5005
R5398 VSS.n4513 VSS.n4512 4.5005
R5399 VSS.n772 VSS.n771 4.5005
R5400 VSS.n935 VSS.n934 4.5005
R5401 VSS.n934 VSS.n933 4.5005
R5402 VSS.n992 VSS.n991 4.5005
R5403 VSS.n991 VSS.n990 4.5005
R5404 VSS.n7893 VSS.t330 4.49023
R5405 VSS.n5025 VSS.t978 4.44646
R5406 VSS.t391 VSS.t396 4.44646
R5407 VSS.n1690 VSS.t304 4.42829
R5408 VSS.n4281 VSS.n4249 4.42582
R5409 VSS.n1682 VSS.n1653 4.42582
R5410 VSS.n1614 VSS.t1 4.411
R5411 VSS.n4201 VSS.t63 4.411
R5412 VSS.n4526 VSS.n4525 4.25879
R5413 VSS.n725 VSS.n724 4.25822
R5414 VSS.n6789 VSS.t41 4.15651
R5415 VSS.t480 VSS.t388 4.12487
R5416 VSS.t388 VSS.t391 4.12487
R5417 VSS.n7816 VSS.t161 4.12487
R5418 VSS.n6974 VSS.t576 4.11964
R5419 VSS.n7300 VSS.n6589 4.11115
R5420 VSS.n7301 VSS.n6587 4.09159
R5421 VSS.n626 VSS.t114 4.04279
R5422 VSS.n651 VSS.t269 4.04279
R5423 VSS.n1541 VSS.t143 4.04279
R5424 VSS.n1557 VSS.t2 4.04279
R5425 VSS.n7101 VSS.t945 3.9607
R5426 VSS.n717 VSS.n716 3.95365
R5427 VSS.n6623 VSS.n6622 3.95365
R5428 VSS.n5306 VSS.n5305 3.95365
R5429 VSS.n777 VSS.n776 3.95358
R5430 VSS.n7124 VSS.n7123 3.95358
R5431 VSS.n6397 VSS.n6396 3.95196
R5432 VSS.n929 VSS.n928 3.95196
R5433 VSS.n4172 VSS.n4171 3.93274
R5434 VSS.n1707 VSS.n1706 3.82995
R5435 VSS.n4328 VSS.n4327 3.82995
R5436 VSS.n4207 VSS.n4206 3.82991
R5437 VSS.n1700 VSS.n1699 3.82991
R5438 VSS.n1613 VSS.n1612 3.82991
R5439 VSS.n4200 VSS.n4199 3.82991
R5440 VSS.n4265 VSS.n4264 3.826
R5441 VSS.n4268 VSS.n4267 3.826
R5442 VSS.n4271 VSS.n4270 3.826
R5443 VSS.n4207 VSS.n4204 3.826
R5444 VSS.n4329 VSS.n4323 3.826
R5445 VSS.n1667 VSS.n1666 3.826
R5446 VSS.n1670 VSS.n1669 3.826
R5447 VSS.n1673 VSS.n1672 3.826
R5448 VSS.n1700 VSS.n1697 3.826
R5449 VSS.n1618 VSS.n1617 3.826
R5450 VSS.n4259 VSS.n4258 3.82596
R5451 VSS.n4262 VSS.n4261 3.82596
R5452 VSS.n1661 VSS.n1660 3.82596
R5453 VSS.n1664 VSS.n1663 3.82596
R5454 VSS.n1708 VSS.n1702 3.82596
R5455 VSS.n1707 VSS.n1704 3.82596
R5456 VSS.n4328 VSS.n4325 3.82596
R5457 VSS.n4210 VSS.n4209 3.82596
R5458 VSS.n4256 VSS.n4255 3.82592
R5459 VSS.n4276 VSS.n4275 3.82592
R5460 VSS.n1719 VSS.n1718 3.82592
R5461 VSS.n1658 VSS.n1657 3.82592
R5462 VSS.n1613 VSS.n1610 3.82592
R5463 VSS.n4200 VSS.n4197 3.82592
R5464 VSS.n4277 VSS.n4273 3.78196
R5465 VSS.n1676 VSS.n1675 3.78196
R5466 VSS.n4588 VSS.t64 3.75122
R5467 VSS.n1615 VSS.t896 3.7355
R5468 VSS.n4202 VSS.t287 3.7355
R5469 VSS.n5237 VSS.n5235 3.68267
R5470 VSS.n7198 VSS.n7197 3.63068
R5471 VSS.n6983 VSS.n6593 3.60687
R5472 VSS.n4662 VSS.n4661 3.59971
R5473 VSS.n4499 VSS.n4498 3.59911
R5474 VSS.n6984 VSS.n6591 3.5873
R5475 VSS.n7891 VSS.n7890 3.48846
R5476 VSS.n4029 VSS.t286 3.45416
R5477 VSS.n1872 VSS.t284 3.45416
R5478 VSS.n1925 VSS.t596 3.41655
R5479 VSS.n2622 VSS.t671 3.41655
R5480 VSS.n2531 VSS.t601 3.41655
R5481 VSS.n2421 VSS.t628 3.41655
R5482 VSS.n2299 VSS.t694 3.41655
R5483 VSS.n2187 VSS.t625 3.41655
R5484 VSS.n2126 VSS.t650 3.41655
R5485 VSS.n1971 VSS.t648 3.41655
R5486 VSS.n1947 VSS.t613 3.41655
R5487 VSS.n1936 VSS.t598 3.41655
R5488 VSS.n5502 VSS.t539 3.41078
R5489 VSS.n5465 VSS.t106 3.41078
R5490 VSS.n5577 VSS.t578 3.41078
R5491 VSS.n5459 VSS.t222 3.41078
R5492 VSS.n5557 VSS.n5555 3.41078
R5493 VSS.n6976 VSS.n6612 3.40289
R5494 VSS.n6714 VSS.n6713 3.40289
R5495 VSS.n1466 VSS.t911 3.38064
R5496 VSS.n4483 VSS.t14 3.38064
R5497 VSS.n728 VSS.n727 3.37941
R5498 VSS.n645 VSS.n632 3.37941
R5499 VSS.n645 VSS.n634 3.37941
R5500 VSS.n5501 VSS.n5500 3.37941
R5501 VSS.n5464 VSS.n5463 3.37941
R5502 VSS.n5458 VSS.n5457 3.37941
R5503 VSS.n5576 VSS.n5575 3.37941
R5504 VSS.n6445 VSS.n6439 3.37941
R5505 VSS.n7095 VSS.n7076 3.37941
R5506 VSS.n5228 VSS.n5225 3.37941
R5507 VSS.n5228 VSS.n5227 3.37941
R5508 VSS.n5346 VSS.n5345 3.37941
R5509 VSS.n6665 VSS.n6664 3.37941
R5510 VSS.n1498 VSS.n1495 3.37941
R5511 VSS.n1498 VSS.n1497 3.37941
R5512 VSS.n4541 VSS.n4540 3.37941
R5513 VSS.n4402 VSS.n4375 3.37941
R5514 VSS.n972 VSS.n966 3.37941
R5515 VSS.n7732 VSS.n7731 3.3685
R5516 VSS.n5368 VSS.n5366 3.3685
R5517 VSS.n6342 VSS.n6340 3.3685
R5518 VSS.n4505 VSS.n4504 3.3685
R5519 VSS.n12 VSS.t924 3.36779
R5520 VSS.n5262 VSS.t840 3.36779
R5521 VSS.n6441 VSS.t563 3.36489
R5522 VSS.n6599 VSS.n6598 3.3442
R5523 VSS.n6607 VSS.n6606 3.3442
R5524 VSS.n23 VSS.t462 3.333
R5525 VSS.n5710 VSS.t430 3.33271
R5526 VSS.n4936 VSS.t502 3.33057
R5527 VSS.n5708 VSS.t469 3.33036
R5528 VSS.n5613 VSS.t500 3.32608
R5529 VSS.n5612 VSS.t507 3.32608
R5530 VSS.n5573 VSS.t443 3.32608
R5531 VSS.n5455 VSS.t425 3.32608
R5532 VSS.n5159 VSS.t428 3.32582
R5533 VSS.n5160 VSS.t450 3.32582
R5534 VSS.n5161 VSS.t476 3.32582
R5535 VSS.n5162 VSS.t460 3.32582
R5536 VSS.n5454 VSS.t509 3.32512
R5537 VSS.n5163 VSS.t386 3.32486
R5538 VSS.n22 VSS.t448 3.31238
R5539 VSS.n5720 VSS.t418 3.31209
R5540 VSS.n4946 VSS.t375 3.31186
R5541 VSS.n5707 VSS.t512 3.3116
R5542 VSS.n4923 VSS.t436 3.31143
R5543 VSS.n5709 VSS.t361 3.31114
R5544 VSS.n727 VSS.t233 3.2765
R5545 VSS.n727 VSS.n726 3.2765
R5546 VSS.n634 VSS.t272 3.2765
R5547 VSS.n634 VSS.n633 3.2765
R5548 VSS.n632 VSS.t115 3.2765
R5549 VSS.n632 VSS.n631 3.2765
R5550 VSS.n5403 VSS.t785 3.2765
R5551 VSS.n5403 VSS.n5402 3.2765
R5552 VSS.n5405 VSS.t969 3.2765
R5553 VSS.n5405 VSS.n5404 3.2765
R5554 VSS.n5415 VSS.t865 3.2765
R5555 VSS.n5415 VSS.n5414 3.2765
R5556 VSS.n5407 VSS.t755 3.2765
R5557 VSS.n5407 VSS.n5406 3.2765
R5558 VSS.n5409 VSS.t971 3.2765
R5559 VSS.n5409 VSS.n5408 3.2765
R5560 VSS.n5822 VSS.t951 3.2765
R5561 VSS.n5822 VSS.n5821 3.2765
R5562 VSS.n5820 VSS.t817 3.2765
R5563 VSS.n5820 VSS.n5819 3.2765
R5564 VSS.n5818 VSS.t871 3.2765
R5565 VSS.n5818 VSS.n5817 3.2765
R5566 VSS.n5500 VSS.t540 3.2765
R5567 VSS.n5500 VSS.n5499 3.2765
R5568 VSS.n5463 VSS.t107 3.2765
R5569 VSS.n5463 VSS.n5462 3.2765
R5570 VSS.n5457 VSS.t223 3.2765
R5571 VSS.n5457 VSS.n5456 3.2765
R5572 VSS.n5575 VSS.t579 3.2765
R5573 VSS.n5575 VSS.n5574 3.2765
R5574 VSS.n5824 VSS.t816 3.2765
R5575 VSS.n5824 VSS.n5823 3.2765
R5576 VSS.n5826 VSS.t870 3.2765
R5577 VSS.n5826 VSS.n5825 3.2765
R5578 VSS.n5425 VSS.t964 3.2765
R5579 VSS.n5425 VSS.n5424 3.2765
R5580 VSS.n5423 VSS.t860 3.2765
R5581 VSS.n5423 VSS.n5422 3.2765
R5582 VSS.n5421 VSS.t733 3.2765
R5583 VSS.n5421 VSS.n5420 3.2765
R5584 VSS.n5427 VSS.t782 3.2765
R5585 VSS.n5427 VSS.n5426 3.2765
R5586 VSS.n5429 VSS.t818 3.2765
R5587 VSS.n5429 VSS.n5428 3.2765
R5588 VSS.n6598 VSS.t559 3.2765
R5589 VSS.n6598 VSS.n6597 3.2765
R5590 VSS.n6591 VSS.t994 3.2765
R5591 VSS.n6591 VSS.n6590 3.2765
R5592 VSS.n6587 VSS.t835 3.2765
R5593 VSS.n6587 VSS.n6586 3.2765
R5594 VSS.n6589 VSS.t535 3.2765
R5595 VSS.n6589 VSS.n6588 3.2765
R5596 VSS.n6593 VSS.t573 3.2765
R5597 VSS.n6593 VSS.n6592 3.2765
R5598 VSS.n6606 VSS.t938 3.2765
R5599 VSS.n6606 VSS.n6605 3.2765
R5600 VSS.n6439 VSS.t988 3.2765
R5601 VSS.n6439 VSS.n6438 3.2765
R5602 VSS.n7076 VSS.t825 3.2765
R5603 VSS.n7076 VSS.n7075 3.2765
R5604 VSS.n6612 VSS.t338 3.2765
R5605 VSS.n6612 VSS.n6611 3.2765
R5606 VSS.n6713 VSS.t75 3.2765
R5607 VSS.n6713 VSS.n6712 3.2765
R5608 VSS.n5005 VSS.t857 3.2765
R5609 VSS.n5005 VSS.n5004 3.2765
R5610 VSS.n5008 VSS.t955 3.2765
R5611 VSS.n5008 VSS.n5007 3.2765
R5612 VSS.n5011 VSS.t735 3.2765
R5613 VSS.n5011 VSS.n5010 3.2765
R5614 VSS.n4955 VSS.t852 3.2765
R5615 VSS.n4955 VSS.n4954 3.2765
R5616 VSS.n4958 VSS.t784 3.2765
R5617 VSS.n4958 VSS.n4957 3.2765
R5618 VSS.n4952 VSS.t960 3.2765
R5619 VSS.n4952 VSS.n4951 3.2765
R5620 VSS.n4888 VSS.t984 3.2765
R5621 VSS.n4888 VSS.n4887 3.2765
R5622 VSS.n4886 VSS.t820 3.2765
R5623 VSS.n4886 VSS.n4885 3.2765
R5624 VSS.n4870 VSS.t791 3.2765
R5625 VSS.n4870 VSS.n4869 3.2765
R5626 VSS.n4961 VSS.t963 3.2765
R5627 VSS.n4961 VSS.n4960 3.2765
R5628 VSS.n4965 VSS.t749 3.2765
R5629 VSS.n4965 VSS.n4964 3.2765
R5630 VSS.n4968 VSS.t794 3.2765
R5631 VSS.n4968 VSS.n4967 3.2765
R5632 VSS.n4971 VSS.t968 3.2765
R5633 VSS.n4971 VSS.n4970 3.2765
R5634 VSS.n4874 VSS.t756 3.2765
R5635 VSS.n4874 VSS.n4873 3.2765
R5636 VSS.n5001 VSS.t728 3.2765
R5637 VSS.n5001 VSS.n5000 3.2765
R5638 VSS.n5227 VSS.t228 3.2765
R5639 VSS.n5227 VSS.n5226 3.2765
R5640 VSS.n5225 VSS.t308 3.2765
R5641 VSS.n5225 VSS.n5224 3.2765
R5642 VSS.n5345 VSS.t761 3.2765
R5643 VSS.n5345 VSS.n5344 3.2765
R5644 VSS.n6664 VSS.t42 3.2765
R5645 VSS.n6664 VSS.n6663 3.2765
R5646 VSS.n1497 VSS.t144 3.2765
R5647 VSS.n1497 VSS.n1496 3.2765
R5648 VSS.n1495 VSS.t878 3.2765
R5649 VSS.n1495 VSS.n1494 3.2765
R5650 VSS.n4540 VSS.t30 3.2765
R5651 VSS.n4540 VSS.n4539 3.2765
R5652 VSS.n4375 VSS.t1003 3.2765
R5653 VSS.n4375 VSS.n4374 3.2765
R5654 VSS.n966 VSS.t274 3.2765
R5655 VSS.n966 VSS.n965 3.2765
R5656 VSS.n5372 VSS.n5370 3.17523
R5657 VSS.n5387 VSS.n5386 3.17523
R5658 VSS.n7737 VSS.n7736 3.17468
R5659 VSS.n4279 VSS.n4252 3.16517
R5660 VSS.n1680 VSS.n1679 3.16517
R5661 VSS.n4219 VSS.n4218 3.1505
R5662 VSS.n4221 VSS.n4220 3.1505
R5663 VSS.n4223 VSS.n4222 3.1505
R5664 VSS.n4225 VSS.n4224 3.1505
R5665 VSS.n4227 VSS.n4226 3.1505
R5666 VSS.n4229 VSS.n4228 3.1505
R5667 VSS.n4231 VSS.n4230 3.1505
R5668 VSS.n4233 VSS.n4232 3.1505
R5669 VSS.n4284 VSS.n4234 3.1505
R5670 VSS.n4283 VSS.n4235 3.1505
R5671 VSS.n4282 VSS.n4236 3.1505
R5672 VSS.n4280 VSS.n4250 3.1505
R5673 VSS.n4216 VSS.n4215 3.1505
R5674 VSS.n1738 VSS.n1737 3.1505
R5675 VSS.n1740 VSS.n1739 3.1505
R5676 VSS.n1746 VSS.n1741 3.1505
R5677 VSS.n1745 VSS.n1742 3.1505
R5678 VSS.n1744 VSS.n1743 3.1505
R5679 VSS.n1634 VSS.n1633 3.1505
R5680 VSS.n1636 VSS.n1635 3.1505
R5681 VSS.n1638 VSS.n1637 3.1505
R5682 VSS.n1686 VSS.n1685 3.1505
R5683 VSS.n1684 VSS.n1639 3.1505
R5684 VSS.n1683 VSS.n1640 3.1505
R5685 VSS.n1681 VSS.n1654 3.1505
R5686 VSS.n1722 VSS.n1721 3.1505
R5687 VSS.n1711 VSS.n1710 3.1505
R5688 VSS.n1621 VSS.n1620 3.1505
R5689 VSS.n5832 VSS.n5818 3.1505
R5690 VSS.n5831 VSS.n5820 3.1505
R5691 VSS.n5828 VSS.n5824 3.1505
R5692 VSS.n5436 VSS.n5421 3.1505
R5693 VSS.n5435 VSS.n5423 3.1505
R5694 VSS.n5432 VSS.n5427 3.1505
R5695 VSS.n5412 VSS.n5407 3.1505
R5696 VSS.n5417 VSS.n5405 3.1505
R5697 VSS.n5418 VSS.n5403 3.1505
R5698 VSS.n4972 VSS.n4971 3.1505
R5699 VSS.n4969 VSS.n4968 3.1505
R5700 VSS.n4962 VSS.n4961 3.1505
R5701 VSS.n5002 VSS.n5001 3.1505
R5702 VSS.n4889 VSS.n4888 3.1505
R5703 VSS.n4959 VSS.n4958 3.1505
R5704 VSS.n4956 VSS.n4955 3.1505
R5705 VSS.n5012 VSS.n5011 3.1505
R5706 VSS.n5009 VSS.n5008 3.1505
R5707 VSS.n4332 VSS.n4331 3.1505
R5708 VSS.n4213 VSS.n4212 3.1505
R5709 VSS.n5368 VSS.n5367 3.11623
R5710 VSS.n7248 VSS.t766 3.08765
R5711 VSS.n7846 VSS.n7845 3.07743
R5712 VSS.n4513 VSS.n722 2.9883
R5713 VSS.n4476 VSS.n1481 2.9883
R5714 VSS.n6748 VSS.n6740 2.9883
R5715 VSS.n7246 VSS.n7245 2.9883
R5716 VSS.n6493 VSS.n6486 2.9883
R5717 VSS.n6942 VSS.n6941 2.9883
R5718 VSS.n5372 VSS.n5371 2.91648
R5719 VSS.n5359 VSS.n5358 2.91633
R5720 VSS.n6361 VSS.n6358 2.86264
R5721 VSS.n811 VSS.n808 2.86264
R5722 VSS.n7142 VSS.n7140 2.85093
R5723 VSS.n5094 VSS.n5093 2.83943
R5724 VSS.n5098 VSS.n5097 2.83943
R5725 VSS.n5207 VSS.n5206 2.83943
R5726 VSS.n5220 VSS.n5219 2.83943
R5727 VSS.n7849 VSS.n7848 2.83943
R5728 VSS.n5765 VSS.n5764 2.83943
R5729 VSS.n5762 VSS.n5761 2.83943
R5730 VSS.n5758 VSS.n5757 2.83943
R5731 VSS.n5738 VSS.n5737 2.83943
R5732 VSS.n5734 VSS.n5733 2.83943
R5733 VSS.n5648 VSS.n5647 2.83943
R5734 VSS.n5644 VSS.n5643 2.83943
R5735 VSS.n5641 VSS.n5640 2.83943
R5736 VSS.n5638 VSS.n5637 2.83943
R5737 VSS.n5634 VSS.n5633 2.83943
R5738 VSS.n7862 VSS.n7861 2.83943
R5739 VSS.n7865 VSS.n7864 2.83943
R5740 VSS.n1391 VSS.n1390 2.81354
R5741 VSS.n9 VSS.n5 2.65705
R5742 VSS.n9 VSS.n8 2.65638
R5743 VSS.n5508 VSS.n5507 2.64393
R5744 VSS.n5470 VSS.n5469 2.64393
R5745 VSS.n5827 VSS.n5826 2.6255
R5746 VSS.n5830 VSS.n5822 2.6255
R5747 VSS.n5434 VSS.n5425 2.6255
R5748 VSS.n5416 VSS.n5415 2.6255
R5749 VSS.n4966 VSS.n4965 2.6255
R5750 VSS.n4890 VSS.n4886 2.6255
R5751 VSS.n4953 VSS.n4952 2.6255
R5752 VSS.n5006 VSS.n5005 2.6255
R5753 VSS.n6211 VSS.n5952 2.61042
R5754 VSS.n6195 VSS.n5954 2.61042
R5755 VSS.n6182 VSS.n5956 2.61042
R5756 VSS.n6042 VSS.n6041 2.60873
R5757 VSS.n4453 VSS.n1483 2.60616
R5758 VSS.n4429 VSS.n4423 2.60562
R5759 VSS.n606 VSS.n603 2.60491
R5760 VSS.n672 VSS.n669 2.60491
R5761 VSS.n1508 VSS.n1505 2.60491
R5762 VSS.n1565 VSS.n1564 2.60491
R5763 VSS.n7795 VSS.n7794 2.60464
R5764 VSS.n5397 VSS.n5396 2.60246
R5765 VSS.n5915 VSS.n5914 2.60244
R5766 VSS.n5936 VSS.n5935 2.60244
R5767 VSS.n7435 VSS.n5381 2.6016
R5768 VSS.n35 VSS.n34 2.60148
R5769 VSS.n4780 VSS.n4772 2.60147
R5770 VSS.n1388 VSS.n764 2.6005
R5771 VSS.n764 VSS.n763 2.6005
R5772 VSS.n1404 VSS.n1403 2.6005
R5773 VSS.n1403 VSS.n1402 2.6005
R5774 VSS.n1400 VSS.n1399 2.6005
R5775 VSS.n1399 VSS.n1398 2.6005
R5776 VSS.n1396 VSS.n1395 2.6005
R5777 VSS.n1395 VSS.n1394 2.6005
R5778 VSS.n1393 VSS.n1392 2.6005
R5779 VSS.n1392 VSS.n1391 2.6005
R5780 VSS.n1406 VSS.n1405 2.6005
R5781 VSS.n732 VSS.n731 2.6005
R5782 VSS.n735 VSS.n734 2.6005
R5783 VSS.n737 VSS.n736 2.6005
R5784 VSS.n739 VSS.n738 2.6005
R5785 VSS VSS.n741 2.6005
R5786 VSS.n743 VSS.n742 2.6005
R5787 VSS.n748 VSS.n747 2.6005
R5788 VSS.n751 VSS.n750 2.6005
R5789 VSS.n753 VSS.n752 2.6005
R5790 VSS.n756 VSS.n755 2.6005
R5791 VSS.n1420 VSS.n1419 2.6005
R5792 VSS.n1418 VSS.n1417 2.6005
R5793 VSS.n1416 VSS.n1415 2.6005
R5794 VSS.n1412 VSS.n1411 2.6005
R5795 VSS.n1410 VSS.n1409 2.6005
R5796 VSS.n6579 VSS.n6578 2.6005
R5797 VSS.n6577 VSS.n6576 2.6005
R5798 VSS.n6574 VSS.n6573 2.6005
R5799 VSS.n6569 VSS.n6568 2.6005
R5800 VSS.n6568 VSS.n6567 2.6005
R5801 VSS.n6572 VSS.n6571 2.6005
R5802 VSS.n6571 VSS.n6570 2.6005
R5803 VSS.n6459 VSS.n6436 2.6005
R5804 VSS.n6436 VSS.n6435 2.6005
R5805 VSS.n6457 VSS.n6456 2.6005
R5806 VSS.n6456 VSS.n6455 2.6005
R5807 VSS.n6454 VSS.n6453 2.6005
R5808 VSS.n6453 VSS.n6452 2.6005
R5809 VSS.n6451 VSS.n6450 2.6005
R5810 VSS.n6450 VSS.n6449 2.6005
R5811 VSS.n6448 VSS.n6447 2.6005
R5812 VSS.n6447 VSS.n6446 2.6005
R5813 VSS VSS.n6444 2.6005
R5814 VSS.n6444 VSS.n6443 2.6005
R5815 VSS.n6442 VSS.n6440 2.6005
R5816 VSS.n6442 VSS.n6441 2.6005
R5817 VSS.n6429 VSS.n6428 2.6005
R5818 VSS.n6428 VSS.n6427 2.6005
R5819 VSS.n6426 VSS.n6425 2.6005
R5820 VSS.n6425 VSS.n6424 2.6005
R5821 VSS.n6423 VSS.n6422 2.6005
R5822 VSS.n6422 VSS.n6421 2.6005
R5823 VSS.n6418 VSS.n6417 2.6005
R5824 VSS.n6417 VSS.n6416 2.6005
R5825 VSS.n6476 VSS.n6475 2.6005
R5826 VSS.n6475 VSS.n6474 2.6005
R5827 VSS.n6479 VSS.n6478 2.6005
R5828 VSS.n6478 VSS.n6477 2.6005
R5829 VSS.n6482 VSS.n6481 2.6005
R5830 VSS.n6481 VSS.n6480 2.6005
R5831 VSS.n6497 VSS.n6496 2.6005
R5832 VSS.n6496 VSS.n6495 2.6005
R5833 VSS.n6500 VSS.n6499 2.6005
R5834 VSS.n6499 VSS.n6498 2.6005
R5835 VSS.n6504 VSS.n6503 2.6005
R5836 VSS.n6503 VSS.n6502 2.6005
R5837 VSS.n6508 VSS.n6507 2.6005
R5838 VSS.n6507 VSS.n6506 2.6005
R5839 VSS.n6511 VSS.n6510 2.6005
R5840 VSS.n6510 VSS.n6509 2.6005
R5841 VSS.n6514 VSS.n6513 2.6005
R5842 VSS.n6513 VSS.n6512 2.6005
R5843 VSS.n6518 VSS.n6517 2.6005
R5844 VSS.n6517 VSS.n6516 2.6005
R5845 VSS.n6521 VSS.n6520 2.6005
R5846 VSS.n6520 VSS.n6519 2.6005
R5847 VSS.n6524 VSS.n6523 2.6005
R5848 VSS.n6523 VSS.n6522 2.6005
R5849 VSS.n6527 VSS.n6526 2.6005
R5850 VSS.n6526 VSS.n6525 2.6005
R5851 VSS.n6530 VSS.n6529 2.6005
R5852 VSS.n6529 VSS.n6528 2.6005
R5853 VSS.n6534 VSS.n6533 2.6005
R5854 VSS.n6533 VSS.n6532 2.6005
R5855 VSS.n6537 VSS.n6536 2.6005
R5856 VSS.n6536 VSS.n6535 2.6005
R5857 VSS.n6540 VSS.n6539 2.6005
R5858 VSS.n6539 VSS.n6538 2.6005
R5859 VSS.n6543 VSS.n6542 2.6005
R5860 VSS.n6542 VSS.n6541 2.6005
R5861 VSS.n6546 VSS.n6545 2.6005
R5862 VSS.n6545 VSS.n6544 2.6005
R5863 VSS.n6549 VSS.n6548 2.6005
R5864 VSS.n6548 VSS.n6547 2.6005
R5865 VSS.n6552 VSS.n6551 2.6005
R5866 VSS.n6551 VSS.n6550 2.6005
R5867 VSS.n6556 VSS.n6555 2.6005
R5868 VSS.n6555 VSS.n6554 2.6005
R5869 VSS.n6559 VSS.n6558 2.6005
R5870 VSS.n6558 VSS.n6557 2.6005
R5871 VSS.n6562 VSS.n6561 2.6005
R5872 VSS.n6561 VSS.n6560 2.6005
R5873 VSS.n6566 VSS.n6565 2.6005
R5874 VSS.n6565 VSS.n6564 2.6005
R5875 VSS.n7323 VSS.n7322 2.6005
R5876 VSS.n7322 VSS.n7321 2.6005
R5877 VSS.n7319 VSS.n7318 2.6005
R5878 VSS.n7318 VSS.n7317 2.6005
R5879 VSS.n7316 VSS.n7315 2.6005
R5880 VSS.n7315 VSS.n7314 2.6005
R5881 VSS.n7313 VSS.n7312 2.6005
R5882 VSS.n7312 VSS.n7311 2.6005
R5883 VSS.n7310 VSS.n7309 2.6005
R5884 VSS.n7306 VSS.n7305 2.6005
R5885 VSS.n6464 VSS.n6463 2.6005
R5886 VSS.n6467 VSS.n6466 2.6005
R5887 VSS.n6469 VSS.n6468 2.6005
R5888 VSS.n6473 VSS.n6472 2.6005
R5889 VSS.n7414 VSS.n7413 2.6005
R5890 VSS.n7397 VSS.n7396 2.6005
R5891 VSS.n7396 VSS.n7395 2.6005
R5892 VSS.n7400 VSS.n7399 2.6005
R5893 VSS.n7399 VSS.n7398 2.6005
R5894 VSS.n7403 VSS.n7402 2.6005
R5895 VSS.n7402 VSS.n7401 2.6005
R5896 VSS.n7406 VSS.n7405 2.6005
R5897 VSS.n7405 VSS.n7404 2.6005
R5898 VSS.n7409 VSS.n7408 2.6005
R5899 VSS.n7408 VSS.n7407 2.6005
R5900 VSS.n7412 VSS.n7411 2.6005
R5901 VSS.n7411 VSS.n7410 2.6005
R5902 VSS.n7415 VSS.n7414 2.6005
R5903 VSS.n7363 VSS.n7362 2.6005
R5904 VSS.n7342 VSS.n7341 2.6005
R5905 VSS.n7341 VSS.n7340 2.6005
R5906 VSS.n7345 VSS.n7344 2.6005
R5907 VSS.n7344 VSS.n7343 2.6005
R5908 VSS.n7349 VSS.n7348 2.6005
R5909 VSS.n7348 VSS.n7347 2.6005
R5910 VSS.n7352 VSS.n7351 2.6005
R5911 VSS.n7351 VSS.n7350 2.6005
R5912 VSS.n7356 VSS.n7355 2.6005
R5913 VSS.n7355 VSS.n7354 2.6005
R5914 VSS.n7359 VSS.n7358 2.6005
R5915 VSS.n7358 VSS.n7357 2.6005
R5916 VSS.n7362 VSS.n7361 2.6005
R5917 VSS.n7063 VSS.n6989 2.6005
R5918 VSS.n6989 VSS.n6988 2.6005
R5919 VSS.n7062 VSS.n7061 2.6005
R5920 VSS.n7061 VSS.n7060 2.6005
R5921 VSS.n7059 VSS.n7058 2.6005
R5922 VSS.n7058 VSS.n7057 2.6005
R5923 VSS.n7056 VSS.n7055 2.6005
R5924 VSS.n7055 VSS.n7054 2.6005
R5925 VSS.n7053 VSS.n7052 2.6005
R5926 VSS.n7052 VSS.n7051 2.6005
R5927 VSS.n7050 VSS.n7049 2.6005
R5928 VSS.n7049 VSS.n7048 2.6005
R5929 VSS.n7017 VSS.n7016 2.6005
R5930 VSS.n7016 VSS.n7015 2.6005
R5931 VSS.n7014 VSS.n7013 2.6005
R5932 VSS.n7013 VSS.n7012 2.6005
R5933 VSS.n7011 VSS.n7010 2.6005
R5934 VSS.n7010 VSS.n7009 2.6005
R5935 VSS.n7008 VSS.n7007 2.6005
R5936 VSS.n7007 VSS.n7006 2.6005
R5937 VSS.n7005 VSS.n7004 2.6005
R5938 VSS.n7004 VSS.n7003 2.6005
R5939 VSS.n7002 VSS.n7001 2.6005
R5940 VSS.n7001 VSS.n7000 2.6005
R5941 VSS.n6999 VSS.n6998 2.6005
R5942 VSS.n6998 VSS.n6997 2.6005
R5943 VSS.n7295 VSS.n7294 2.6005
R5944 VSS.n7281 VSS.n7280 2.6005
R5945 VSS.n7280 VSS.n7279 2.6005
R5946 VSS.n7284 VSS.n7283 2.6005
R5947 VSS.n7283 VSS.n7282 2.6005
R5948 VSS.n7287 VSS.n7286 2.6005
R5949 VSS.n7286 VSS.n7285 2.6005
R5950 VSS.n7290 VSS.n7289 2.6005
R5951 VSS.n7289 VSS.n7288 2.6005
R5952 VSS.n7293 VSS.n7292 2.6005
R5953 VSS.n7292 VSS.n7291 2.6005
R5954 VSS.n7296 VSS.n7295 2.6005
R5955 VSS.t908 VSS.t937 2.6005
R5956 VSS.t937 VSS.t939 2.6005
R5957 VSS.t907 VSS.t936 2.6005
R5958 VSS.t936 VSS.t839 2.6005
R5959 VSS.n7339 VSS.n7338 2.6005
R5960 VSS.n7338 VSS.n7337 2.6005
R5961 VSS.n7335 VSS.n7334 2.6005
R5962 VSS.n7334 VSS.n7333 2.6005
R5963 VSS.n7072 VSS.n7071 2.6005
R5964 VSS.n7071 VSS.n7070 2.6005
R5965 VSS.n7069 VSS.n7068 2.6005
R5966 VSS.n7068 VSS.n7067 2.6005
R5967 VSS.n7066 VSS.n7065 2.6005
R5968 VSS.n7065 VSS.n7064 2.6005
R5969 VSS.n7332 VSS.n7331 2.6005
R5970 VSS.n7328 VSS.n7327 2.6005
R5971 VSS.n7326 VSS.n7325 2.6005
R5972 VSS.n6973 VSS 2.6005
R5973 VSS.n6973 VSS.n6972 2.6005
R5974 VSS VSS.n6975 2.6005
R5975 VSS.n6975 VSS.n6974 2.6005
R5976 VSS.n6715 VSS 2.6005
R5977 VSS.n6716 VSS.n6715 2.6005
R5978 VSS VSS.n6711 2.6005
R5979 VSS.n6711 VSS.n6710 2.6005
R5980 VSS.n5068 VSS.n5067 2.6005
R5981 VSS.n5067 VSS.n5066 2.6005
R5982 VSS.n5065 VSS.n5064 2.6005
R5983 VSS.n5064 VSS.n5063 2.6005
R5984 VSS.n5062 VSS.n5061 2.6005
R5985 VSS.n5061 VSS.n5060 2.6005
R5986 VSS.n5166 VSS.n5165 2.6005
R5987 VSS.n5165 VSS.n5164 2.6005
R5988 VSS.n5169 VSS.n5168 2.6005
R5989 VSS.n5168 VSS.n5167 2.6005
R5990 VSS.n5172 VSS.n5171 2.6005
R5991 VSS.n5171 VSS.n5170 2.6005
R5992 VSS.n5175 VSS.n5174 2.6005
R5993 VSS.n5174 VSS.n5173 2.6005
R5994 VSS.n5178 VSS.n5177 2.6005
R5995 VSS.n5177 VSS.n5176 2.6005
R5996 VSS.n5181 VSS.n5180 2.6005
R5997 VSS.n5180 VSS.n5179 2.6005
R5998 VSS.n5184 VSS.n5183 2.6005
R5999 VSS.n5183 VSS.n5182 2.6005
R6000 VSS.n5187 VSS.n5186 2.6005
R6001 VSS.n5186 VSS.n5185 2.6005
R6002 VSS.n5190 VSS.n5189 2.6005
R6003 VSS.n5189 VSS.n5188 2.6005
R6004 VSS.n5193 VSS.n5192 2.6005
R6005 VSS.n5192 VSS.n5191 2.6005
R6006 VSS.n5196 VSS.n5195 2.6005
R6007 VSS.n5195 VSS.n5194 2.6005
R6008 VSS.n4985 VSS.n4984 2.6005
R6009 VSS.n4984 VSS.n4983 2.6005
R6010 VSS.n4988 VSS.n4987 2.6005
R6011 VSS.n4987 VSS.n4986 2.6005
R6012 VSS.n4982 VSS.n4981 2.6005
R6013 VSS.n4981 VSS.n4980 2.6005
R6014 VSS.n4992 VSS.n4991 2.6005
R6015 VSS.n4991 VSS.n4990 2.6005
R6016 VSS.n4995 VSS.n4994 2.6005
R6017 VSS.n4994 VSS.n4993 2.6005
R6018 VSS.n4998 VSS.n4997 2.6005
R6019 VSS.n4997 VSS.n4996 2.6005
R6020 VSS.n5017 VSS.n5016 2.6005
R6021 VSS.n5016 VSS.n5015 2.6005
R6022 VSS.n5021 VSS.n5020 2.6005
R6023 VSS.n5020 VSS.n5019 2.6005
R6024 VSS.n5024 VSS.n5023 2.6005
R6025 VSS.n5023 VSS.n5022 2.6005
R6026 VSS.n5027 VSS.n5026 2.6005
R6027 VSS.n5026 VSS.n5025 2.6005
R6028 VSS.n5031 VSS.n5030 2.6005
R6029 VSS.n5030 VSS.n5029 2.6005
R6030 VSS.n4949 VSS.n4948 2.6005
R6031 VSS.n4948 VSS.n4947 2.6005
R6032 VSS.n5036 VSS.n5035 2.6005
R6033 VSS.n5035 VSS.n5034 2.6005
R6034 VSS.n5040 VSS.n5039 2.6005
R6035 VSS.n5039 VSS.n5038 2.6005
R6036 VSS.n5043 VSS.n5042 2.6005
R6037 VSS.n5042 VSS.n5041 2.6005
R6038 VSS.n45 VSS.n44 2.6005
R6039 VSS.n41 VSS.n40 2.6005
R6040 VSS.n38 VSS.n37 2.6005
R6041 VSS.n4769 VSS.n4768 2.6005
R6042 VSS.n4767 VSS.n4766 2.6005
R6043 VSS.n4763 VSS.n4762 2.6005
R6044 VSS.n32 VSS.n31 2.6005
R6045 VSS.n5047 VSS.n5046 2.6005
R6046 VSS.n5046 VSS.n5045 2.6005
R6047 VSS.n5050 VSS.n5049 2.6005
R6048 VSS.n5049 VSS.n5048 2.6005
R6049 VSS.n5053 VSS.n5052 2.6005
R6050 VSS.n5052 VSS.n5051 2.6005
R6051 VSS.n5056 VSS.n5055 2.6005
R6052 VSS.n5055 VSS.n5054 2.6005
R6053 VSS.n5059 VSS.n5058 2.6005
R6054 VSS.n5058 VSS.n5057 2.6005
R6055 VSS.n5070 VSS.n5069 2.6005
R6056 VSS.n5077 VSS.n5076 2.6005
R6057 VSS.n5080 VSS.n5079 2.6005
R6058 VSS.n5074 VSS.n5073 2.6005
R6059 VSS.n5085 VSS.n5084 2.6005
R6060 VSS.n5088 VSS.n5087 2.6005
R6061 VSS.n5091 VSS.n5090 2.6005
R6062 VSS.n5095 VSS.n5094 2.6005
R6063 VSS.n5099 VSS.n5098 2.6005
R6064 VSS.n5104 VSS.n5103 2.6005
R6065 VSS.n5199 VSS.n5198 2.6005
R6066 VSS.n5198 VSS.n5197 2.6005
R6067 VSS.n5202 VSS.n5201 2.6005
R6068 VSS.n5204 VSS.n5203 2.6005
R6069 VSS.n5208 VSS.n5207 2.6005
R6070 VSS.n5212 VSS.n5211 2.6005
R6071 VSS.n5215 VSS.n5214 2.6005
R6072 VSS.n5218 VSS.n5217 2.6005
R6073 VSS.n5221 VSS.n5220 2.6005
R6074 VSS.n7850 VSS.n7849 2.6005
R6075 VSS.n7854 VSS.n7853 2.6005
R6076 VSS.n7801 VSS.n5232 2.6005
R6077 VSS.n7834 VSS.n7831 2.6005
R6078 VSS.n7830 VSS.n7827 2.6005
R6079 VSS.n7826 VSS.n7823 2.6005
R6080 VSS.n7822 VSS.n5230 2.6005
R6081 VSS.n5230 VSS.n5229 2.6005
R6082 VSS VSS.n7819 2.6005
R6083 VSS.n7819 VSS.n7818 2.6005
R6084 VSS.n7817 VSS.n7815 2.6005
R6085 VSS.n7817 VSS.n7816 2.6005
R6086 VSS.n7814 VSS.n7811 2.6005
R6087 VSS.n7810 VSS.n7808 2.6005
R6088 VSS.n7808 VSS.n7807 2.6005
R6089 VSS.n7806 VSS.n7804 2.6005
R6090 VSS.n7804 VSS.n7803 2.6005
R6091 VSS.n7844 VSS.n7838 2.6005
R6092 VSS.n7838 VSS.n7837 2.6005
R6093 VSS.n7834 VSS.n7833 2.6005
R6094 VSS.n7833 VSS.n7832 2.6005
R6095 VSS.n7830 VSS.n7829 2.6005
R6096 VSS.n7829 VSS.n7828 2.6005
R6097 VSS.n7826 VSS.n7825 2.6005
R6098 VSS.n7825 VSS.n7824 2.6005
R6099 VSS.n7822 VSS.n7821 2.6005
R6100 VSS.n7820 VSS 2.6005
R6101 VSS.n7814 VSS.n7813 2.6005
R6102 VSS.n7813 VSS.n7812 2.6005
R6103 VSS.n7810 VSS.n7809 2.6005
R6104 VSS.n7806 VSS.n7805 2.6005
R6105 VSS.n7801 VSS.n7800 2.6005
R6106 VSS.n7800 VSS.n7799 2.6005
R6107 VSS.n7844 VSS.n7843 2.6005
R6108 VSS.n7632 VSS.n7631 2.6005
R6109 VSS.n7631 VSS.n7630 2.6005
R6110 VSS.n7554 VSS.n7553 2.6005
R6111 VSS.n7553 VSS.n7552 2.6005
R6112 VSS.n6928 VSS.n6927 2.6005
R6113 VSS.n6927 VSS.n6926 2.6005
R6114 VSS.n6931 VSS.n6930 2.6005
R6115 VSS.n6930 VSS.n6929 2.6005
R6116 VSS.n7551 VSS.n7550 2.6005
R6117 VSS.n7550 VSS.n7549 2.6005
R6118 VSS.n7547 VSS.n7546 2.6005
R6119 VSS.n7546 VSS.n7545 2.6005
R6120 VSS.n7543 VSS.n7542 2.6005
R6121 VSS.n7542 VSS.n7541 2.6005
R6122 VSS.n6916 VSS.n6915 2.6005
R6123 VSS.n6919 VSS.n6918 2.6005
R6124 VSS.n6918 VSS.n6917 2.6005
R6125 VSS.n6915 VSS.n6914 2.6005
R6126 VSS.n7740 VSS.n5299 2.6005
R6127 VSS.n5362 VSS.n5361 2.6005
R6128 VSS.n5364 VSS.n5363 2.6005
R6129 VSS.n5303 VSS.n5302 2.6005
R6130 VSS.n7727 VSS.n7726 2.6005
R6131 VSS.n5379 VSS.n5378 2.6005
R6132 VSS.n5376 VSS.n5375 2.6005
R6133 VSS.n5301 VSS.n5300 2.6005
R6134 VSS.n7265 VSS.n7264 2.6005
R6135 VSS.n7267 VSS.n7266 2.6005
R6136 VSS.n7272 VSS.n7271 2.6005
R6137 VSS.n7262 VSS.n7261 2.6005
R6138 VSS.n7257 VSS.n7256 2.6005
R6139 VSS.n7256 VSS.n7255 2.6005
R6140 VSS.n7254 VSS.n7253 2.6005
R6141 VSS.n7253 VSS.n7252 2.6005
R6142 VSS.n7250 VSS.n7249 2.6005
R6143 VSS.n7249 VSS.n7248 2.6005
R6144 VSS.n7241 VSS.n7240 2.6005
R6145 VSS.n7240 VSS.n7239 2.6005
R6146 VSS.n7238 VSS.n7237 2.6005
R6147 VSS.n7237 VSS.n7236 2.6005
R6148 VSS.n7222 VSS.n7221 2.6005
R6149 VSS.n7221 VSS.n7220 2.6005
R6150 VSS.n7219 VSS.n7218 2.6005
R6151 VSS.n7218 VSS.n7217 2.6005
R6152 VSS.n7216 VSS.n7215 2.6005
R6153 VSS.n7215 VSS.n7214 2.6005
R6154 VSS.n7212 VSS.n7211 2.6005
R6155 VSS.n7211 VSS.n7210 2.6005
R6156 VSS.n7260 VSS.n7259 2.6005
R6157 VSS.n7259 VSS.n7258 2.6005
R6158 VSS.n7274 VSS.n7273 2.6005
R6159 VSS.n7278 VSS.n7277 2.6005
R6160 VSS.n7366 VSS.n7365 2.6005
R6161 VSS.n7365 VSS.n7364 2.6005
R6162 VSS.n7369 VSS.n7368 2.6005
R6163 VSS.n7368 VSS.n7367 2.6005
R6164 VSS.n7372 VSS.n7371 2.6005
R6165 VSS.n7371 VSS.n7370 2.6005
R6166 VSS.n7375 VSS.n7374 2.6005
R6167 VSS.n7374 VSS.n7373 2.6005
R6168 VSS.n7380 VSS.n7379 2.6005
R6169 VSS.n7379 VSS.n7378 2.6005
R6170 VSS.n7383 VSS.n7382 2.6005
R6171 VSS.n7382 VSS.n7381 2.6005
R6172 VSS.n7386 VSS.n7385 2.6005
R6173 VSS.n7385 VSS.n7384 2.6005
R6174 VSS.n7389 VSS.n7388 2.6005
R6175 VSS.n7388 VSS.n7387 2.6005
R6176 VSS.n7392 VSS.n7391 2.6005
R6177 VSS.n7391 VSS.n7390 2.6005
R6178 VSS.n7047 VSS.n7046 2.6005
R6179 VSS.n7046 VSS.n7045 2.6005
R6180 VSS.n7044 VSS.n7043 2.6005
R6181 VSS.n7043 VSS.n7042 2.6005
R6182 VSS.n7041 VSS.n7040 2.6005
R6183 VSS.n7040 VSS.n7039 2.6005
R6184 VSS.n7038 VSS.n7037 2.6005
R6185 VSS.n7037 VSS.n7036 2.6005
R6186 VSS.n7035 VSS.n7034 2.6005
R6187 VSS.n7034 VSS.n7033 2.6005
R6188 VSS.n7032 VSS.n7031 2.6005
R6189 VSS.n7031 VSS.n7030 2.6005
R6190 VSS.n7029 VSS.n7028 2.6005
R6191 VSS.n7028 VSS.n7027 2.6005
R6192 VSS.n7026 VSS.n7025 2.6005
R6193 VSS.n7025 VSS.n7024 2.6005
R6194 VSS.n7023 VSS.n7022 2.6005
R6195 VSS.n7022 VSS.n7021 2.6005
R6196 VSS.n7020 VSS.n7019 2.6005
R6197 VSS.n7019 VSS.n7018 2.6005
R6198 VSS.n6580 VSS.n6392 2.6005
R6199 VSS.n6388 VSS.n6387 2.6005
R6200 VSS.n6385 VSS.n6384 2.6005
R6201 VSS.n6381 VSS.n6380 2.6005
R6202 VSS.n6379 VSS.n6378 2.6005
R6203 VSS.n6376 VSS.n6375 2.6005
R6204 VSS.n6375 VSS.n6374 2.6005
R6205 VSS.n6372 VSS.n6371 2.6005
R6206 VSS.n6370 VSS.n6369 2.6005
R6207 VSS.n6368 VSS.n6367 2.6005
R6208 VSS.n6367 VSS.n6366 2.6005
R6209 VSS.n6585 VSS.n6584 2.6005
R6210 VSS.n6584 VSS.n6583 2.6005
R6211 VSS.n7417 VSS.n7416 2.6005
R6212 VSS.n7421 VSS.n7420 2.6005
R6213 VSS.n6363 VSS.n6362 2.6005
R6214 VSS.n6995 VSS.n6994 2.6005
R6215 VSS.n6993 VSS.n6992 2.6005
R6216 VSS.n6349 VSS.n6348 2.6005
R6217 VSS.n6348 VSS.n6347 2.6005
R6218 VSS.n6346 VSS.n6345 2.6005
R6219 VSS.n6345 VSS.n6344 2.6005
R6220 VSS.n6353 VSS.n6352 2.6005
R6221 VSS.n6352 VSS.n6351 2.6005
R6222 VSS.n6356 VSS.n6355 2.6005
R6223 VSS.n6355 VSS.n6354 2.6005
R6224 VSS.n6360 VSS.n6359 2.6005
R6225 VSS.n6358 VSS.n6357 2.6005
R6226 VSS.n6350 VSS.n6343 2.6005
R6227 VSS.n7085 VSS.n7084 2.6005
R6228 VSS.n7084 VSS.n7083 2.6005
R6229 VSS.n7088 VSS.n7087 2.6005
R6230 VSS.n7087 VSS.n7086 2.6005
R6231 VSS.n7091 VSS.n7090 2.6005
R6232 VSS.n7090 VSS.n7089 2.6005
R6233 VSS.n7094 VSS.n7093 2.6005
R6234 VSS.n7093 VSS.n7092 2.6005
R6235 VSS.n7196 VSS 2.6005
R6236 VSS.n7197 VSS.n7196 2.6005
R6237 VSS.n7195 VSS.n7194 2.6005
R6238 VSS.n7194 VSS.n7193 2.6005
R6239 VSS.n7191 VSS.n7190 2.6005
R6240 VSS.n7190 VSS.n7189 2.6005
R6241 VSS.n7188 VSS.n7187 2.6005
R6242 VSS.n7187 VSS.n7186 2.6005
R6243 VSS.n7185 VSS.n7184 2.6005
R6244 VSS.n7184 VSS.n7183 2.6005
R6245 VSS.n7181 VSS.n7180 2.6005
R6246 VSS.n7180 VSS.n7179 2.6005
R6247 VSS.n7081 VSS.n7080 2.6005
R6248 VSS.n7080 VSS.n7079 2.6005
R6249 VSS.n6332 VSS.n6331 2.6005
R6250 VSS.n6334 VSS.n6333 2.6005
R6251 VSS.n6338 VSS.n6337 2.6005
R6252 VSS.n7209 VSS.n7208 2.6005
R6253 VSS.n7208 VSS.n7207 2.6005
R6254 VSS.n7206 VSS.n7205 2.6005
R6255 VSS.n7205 VSS.n7204 2.6005
R6256 VSS.n7203 VSS.n7202 2.6005
R6257 VSS.n7202 VSS.n7201 2.6005
R6258 VSS.n7200 VSS.n7199 2.6005
R6259 VSS.n7199 VSS.n7198 2.6005
R6260 VSS.n7100 VSS.n7099 2.6005
R6261 VSS.n7099 VSS.n7098 2.6005
R6262 VSS.n7103 VSS.n7102 2.6005
R6263 VSS.n7102 VSS.n7101 2.6005
R6264 VSS.n7106 VSS.n7105 2.6005
R6265 VSS.n7105 VSS.n7104 2.6005
R6266 VSS.n7109 VSS.n7108 2.6005
R6267 VSS.n7108 VSS.n7107 2.6005
R6268 VSS.n7112 VSS.n7111 2.6005
R6269 VSS.n7111 VSS.n7110 2.6005
R6270 VSS.n7115 VSS.n7114 2.6005
R6271 VSS.n7114 VSS.n7113 2.6005
R6272 VSS.n7118 VSS.n7117 2.6005
R6273 VSS.n7117 VSS.n7116 2.6005
R6274 VSS.n7131 VSS.n7130 2.6005
R6275 VSS.n7130 VSS.n7129 2.6005
R6276 VSS.n7134 VSS.n7133 2.6005
R6277 VSS.n7133 VSS.n7132 2.6005
R6278 VSS.n7137 VSS.n7136 2.6005
R6279 VSS.n7136 VSS.n7135 2.6005
R6280 VSS.n7161 VSS.n7160 2.6005
R6281 VSS.n7160 VSS.n7159 2.6005
R6282 VSS.n7157 VSS.n7156 2.6005
R6283 VSS.n7156 VSS.n7155 2.6005
R6284 VSS.n7154 VSS.n7153 2.6005
R6285 VSS.n7153 VSS.n7152 2.6005
R6286 VSS.n5888 VSS.n5887 2.6005
R6287 VSS.n6157 VSS.n6156 2.6005
R6288 VSS.n6221 VSS.n6220 2.6005
R6289 VSS.n6220 VSS.n6219 2.6005
R6290 VSS.n6224 VSS.n6223 2.6005
R6291 VSS.n6223 VSS.n6222 2.6005
R6292 VSS.n5918 VSS.n5917 2.6005
R6293 VSS.n5893 VSS.n5892 2.6005
R6294 VSS.n5886 VSS.n5885 2.6005
R6295 VSS.n5882 VSS.n5881 2.6005
R6296 VSS.n5880 VSS.n5879 2.6005
R6297 VSS.n5944 VSS.n5943 2.6005
R6298 VSS.n5724 VSS.n5723 2.6005
R6299 VSS.n5726 VSS.n5725 2.6005
R6300 VSS.n5712 VSS.n5711 2.6005
R6301 VSS.n5729 VSS.n5728 2.6005
R6302 VSS.n5731 VSS.n5730 2.6005
R6303 VSS.n5735 VSS.n5734 2.6005
R6304 VSS.n5739 VSS.n5738 2.6005
R6305 VSS.n5759 VSS.n5758 2.6005
R6306 VSS.n5763 VSS.n5762 2.6005
R6307 VSS.n5766 VSS.n5765 2.6005
R6308 VSS.n5797 VSS.n5796 2.6005
R6309 VSS.n5796 VSS.n5795 2.6005
R6310 VSS.n5800 VSS.n5799 2.6005
R6311 VSS.n5799 VSS.n5798 2.6005
R6312 VSS.n5803 VSS.n5802 2.6005
R6313 VSS.n5802 VSS.n5801 2.6005
R6314 VSS.n5706 VSS.n5705 2.6005
R6315 VSS.n6114 VSS.n6113 2.6005
R6316 VSS.n6111 VSS.n6110 2.6005
R6317 VSS.n5616 VSS.n5615 2.6005
R6318 VSS.n5618 VSS.n5617 2.6005
R6319 VSS.n5620 VSS.n5619 2.6005
R6320 VSS.n5623 VSS.n5622 2.6005
R6321 VSS.n5625 VSS.n5624 2.6005
R6322 VSS.n5628 VSS.n5627 2.6005
R6323 VSS.n5631 VSS.n5630 2.6005
R6324 VSS.n5635 VSS.n5634 2.6005
R6325 VSS.n5639 VSS.n5638 2.6005
R6326 VSS.n5642 VSS.n5641 2.6005
R6327 VSS.n5645 VSS.n5644 2.6005
R6328 VSS.n5649 VSS.n5648 2.6005
R6329 VSS.n5660 VSS.n5659 2.6005
R6330 VSS.n6116 VSS.n6115 2.6005
R6331 VSS.n5661 VSS.n5453 2.6005
R6332 VSS.n5453 VSS.n5452 2.6005
R6333 VSS.n5665 VSS.n5664 2.6005
R6334 VSS.n5664 VSS.n5663 2.6005
R6335 VSS.n5668 VSS.n5667 2.6005
R6336 VSS.n5667 VSS.n5666 2.6005
R6337 VSS.n5671 VSS.n5670 2.6005
R6338 VSS.n5670 VSS.n5669 2.6005
R6339 VSS.n5674 VSS.n5673 2.6005
R6340 VSS.n5673 VSS.n5672 2.6005
R6341 VSS.n5677 VSS.n5676 2.6005
R6342 VSS.n5676 VSS.n5675 2.6005
R6343 VSS.n5680 VSS.n5679 2.6005
R6344 VSS.n5679 VSS.n5678 2.6005
R6345 VSS.n5683 VSS.n5682 2.6005
R6346 VSS.n5682 VSS.n5681 2.6005
R6347 VSS.n5686 VSS.n5685 2.6005
R6348 VSS.n5685 VSS.n5684 2.6005
R6349 VSS.n5689 VSS.n5688 2.6005
R6350 VSS.n5688 VSS.n5687 2.6005
R6351 VSS.n5692 VSS.n5691 2.6005
R6352 VSS.n5691 VSS.n5690 2.6005
R6353 VSS.n5695 VSS.n5694 2.6005
R6354 VSS.n5694 VSS.n5693 2.6005
R6355 VSS.n5698 VSS.n5697 2.6005
R6356 VSS.n5697 VSS.n5696 2.6005
R6357 VSS.n5701 VSS.n5700 2.6005
R6358 VSS.n5700 VSS.n5699 2.6005
R6359 VSS.n5704 VSS.n5703 2.6005
R6360 VSS.n5703 VSS.n5702 2.6005
R6361 VSS.n5394 VSS.n5393 2.6005
R6362 VSS.n5393 VSS.n5392 2.6005
R6363 VSS.n5391 VSS.n5390 2.6005
R6364 VSS.n5390 VSS.n5389 2.6005
R6365 VSS.n5867 VSS.n5866 2.6005
R6366 VSS.n5866 VSS.n5865 2.6005
R6367 VSS.n5863 VSS.n5862 2.6005
R6368 VSS.n5862 VSS.n5861 2.6005
R6369 VSS.n5860 VSS.n5859 2.6005
R6370 VSS.n5859 VSS.n5858 2.6005
R6371 VSS.n5857 VSS.n5856 2.6005
R6372 VSS.n5856 VSS.n5855 2.6005
R6373 VSS.n5853 VSS.n5852 2.6005
R6374 VSS.n5852 VSS.n5851 2.6005
R6375 VSS.n5850 VSS.n5849 2.6005
R6376 VSS.n5849 VSS.n5848 2.6005
R6377 VSS.n5847 VSS.n5846 2.6005
R6378 VSS.n5846 VSS.n5845 2.6005
R6379 VSS.n5844 VSS.n5843 2.6005
R6380 VSS.n5843 VSS.n5842 2.6005
R6381 VSS.n5442 VSS.n5441 2.6005
R6382 VSS.n5441 VSS.n5440 2.6005
R6383 VSS.n5840 VSS.n5839 2.6005
R6384 VSS.n5839 VSS.n5838 2.6005
R6385 VSS.n5836 VSS.n5835 2.6005
R6386 VSS.n5835 VSS.n5834 2.6005
R6387 VSS.n5816 VSS.n5815 2.6005
R6388 VSS.n5815 VSS.n5814 2.6005
R6389 VSS.n5813 VSS.n5812 2.6005
R6390 VSS.n5812 VSS.n5811 2.6005
R6391 VSS.n5809 VSS.n5808 2.6005
R6392 VSS.n5808 VSS.n5807 2.6005
R6393 VSS.n5806 VSS.n5805 2.6005
R6394 VSS.n5805 VSS.n5804 2.6005
R6395 VSS.n5790 VSS.n5789 2.6005
R6396 VSS.n5787 VSS.n5786 2.6005
R6397 VSS.n5793 VSS.n5792 2.6005
R6398 VSS.n6105 VSS.n6104 2.6005
R6399 VSS.n5948 VSS.n5947 2.6005
R6400 VSS.n6218 VSS.n6217 2.6005
R6401 VSS.n6217 VSS.n6216 2.6005
R6402 VSS.n6214 VSS.n6213 2.6005
R6403 VSS.n6213 VSS.n6212 2.6005
R6404 VSS.n5952 VSS.n5951 2.6005
R6405 VSS.n6210 VSS.n6209 2.6005
R6406 VSS.n6209 VSS.n6208 2.6005
R6407 VSS.n6207 VSS.n6206 2.6005
R6408 VSS.n6206 VSS.n6205 2.6005
R6409 VSS.n6204 VSS.n6203 2.6005
R6410 VSS.n6203 VSS.n6202 2.6005
R6411 VSS.n6201 VSS.n6200 2.6005
R6412 VSS.n6200 VSS.n6199 2.6005
R6413 VSS.n6198 VSS.n6197 2.6005
R6414 VSS.n6197 VSS.n6196 2.6005
R6415 VSS.n5954 VSS.n5953 2.6005
R6416 VSS.n6194 VSS.n6193 2.6005
R6417 VSS.n6193 VSS.n6192 2.6005
R6418 VSS.n6191 VSS.n6190 2.6005
R6419 VSS.n6190 VSS.n6189 2.6005
R6420 VSS.n6188 VSS.n6187 2.6005
R6421 VSS.n6187 VSS.n6186 2.6005
R6422 VSS.n6185 VSS.n6184 2.6005
R6423 VSS.n6184 VSS.n6183 2.6005
R6424 VSS.n5956 VSS.n5955 2.6005
R6425 VSS.n6181 VSS.n6180 2.6005
R6426 VSS.n6180 VSS.n6179 2.6005
R6427 VSS.n6178 VSS.n6177 2.6005
R6428 VSS.n6177 VSS.n6176 2.6005
R6429 VSS.n6170 VSS.n6169 2.6005
R6430 VSS.n6169 VSS.n6168 2.6005
R6431 VSS.n6167 VSS.n6166 2.6005
R6432 VSS.n6166 VSS.n6165 2.6005
R6433 VSS.n6164 VSS.n6163 2.6005
R6434 VSS.n6163 VSS.n6162 2.6005
R6435 VSS.n6161 VSS.n6160 2.6005
R6436 VSS.n6160 VSS.n6159 2.6005
R6437 VSS.n6109 VSS.n6108 2.6005
R6438 VSS.n6108 VSS.n6107 2.6005
R6439 VSS.n6122 VSS.n6121 2.6005
R6440 VSS.n6121 VSS.n6120 2.6005
R6441 VSS.n6125 VSS.n6124 2.6005
R6442 VSS.n6124 VSS.n6123 2.6005
R6443 VSS.n6128 VSS.n6127 2.6005
R6444 VSS.n6127 VSS.n6126 2.6005
R6445 VSS.n6131 VSS.n6130 2.6005
R6446 VSS.n6130 VSS.n6129 2.6005
R6447 VSS.n6134 VSS.n6133 2.6005
R6448 VSS.n6133 VSS.n6132 2.6005
R6449 VSS.n6137 VSS.n6136 2.6005
R6450 VSS.n6136 VSS.n6135 2.6005
R6451 VSS.n6140 VSS.n6139 2.6005
R6452 VSS.n6139 VSS.n6138 2.6005
R6453 VSS.n6143 VSS.n6142 2.6005
R6454 VSS.n6142 VSS.n6141 2.6005
R6455 VSS.n6146 VSS.n6145 2.6005
R6456 VSS.n6145 VSS.n6144 2.6005
R6457 VSS.n6149 VSS.n6148 2.6005
R6458 VSS.n6148 VSS.n6147 2.6005
R6459 VSS.n6152 VSS.n6151 2.6005
R6460 VSS.n6151 VSS.n6150 2.6005
R6461 VSS.n6155 VSS.n6154 2.6005
R6462 VSS.n6154 VSS.n6153 2.6005
R6463 VSS.n6119 VSS.n6118 2.6005
R6464 VSS.n6118 VSS.n6117 2.6005
R6465 VSS.n5401 VSS.n5400 2.6005
R6466 VSS.n7725 VSS.n7724 2.6005
R6467 VSS.n7724 VSS.n7723 2.6005
R6468 VSS.n7722 VSS.n7721 2.6005
R6469 VSS.n7721 VSS.n7720 2.6005
R6470 VSS.n7719 VSS.n7718 2.6005
R6471 VSS.n7718 VSS.n7717 2.6005
R6472 VSS.n7716 VSS.n7715 2.6005
R6473 VSS.n7715 VSS.n7714 2.6005
R6474 VSS.n7713 VSS.n7712 2.6005
R6475 VSS.n7712 VSS.n7711 2.6005
R6476 VSS.n7707 VSS.n7706 2.6005
R6477 VSS.n7706 VSS.n7705 2.6005
R6478 VSS.n7704 VSS.n7703 2.6005
R6479 VSS.n7703 VSS.n7702 2.6005
R6480 VSS.n7701 VSS.n7700 2.6005
R6481 VSS.n7700 VSS.n7699 2.6005
R6482 VSS.n7698 VSS.n7697 2.6005
R6483 VSS.n7697 VSS.n7696 2.6005
R6484 VSS.n7695 VSS.n7694 2.6005
R6485 VSS.n7694 VSS.n7693 2.6005
R6486 VSS.n7692 VSS.n7691 2.6005
R6487 VSS.n7691 VSS.n7690 2.6005
R6488 VSS.n7689 VSS.n7688 2.6005
R6489 VSS.n7688 VSS.n7687 2.6005
R6490 VSS.n7686 VSS.n7685 2.6005
R6491 VSS.n7685 VSS.n7684 2.6005
R6492 VSS.n7683 VSS.n7682 2.6005
R6493 VSS.n7682 VSS.n7681 2.6005
R6494 VSS.n7680 VSS.n7679 2.6005
R6495 VSS.n7679 VSS.n7678 2.6005
R6496 VSS.n7677 VSS.n7676 2.6005
R6497 VSS.n7676 VSS.n7675 2.6005
R6498 VSS.n7744 VSS.n7743 2.6005
R6499 VSS.n7743 VSS.n7742 2.6005
R6500 VSS.n7748 VSS.n7747 2.6005
R6501 VSS.n7747 VSS.n7746 2.6005
R6502 VSS.n7751 VSS.n7750 2.6005
R6503 VSS.n7750 VSS.n7749 2.6005
R6504 VSS.n7754 VSS.n7753 2.6005
R6505 VSS.n7753 VSS.n7752 2.6005
R6506 VSS.n7757 VSS.n7756 2.6005
R6507 VSS.n7756 VSS.n7755 2.6005
R6508 VSS.n7760 VSS.n7759 2.6005
R6509 VSS.n7759 VSS.n7758 2.6005
R6510 VSS.n7763 VSS.n7762 2.6005
R6511 VSS.n7762 VSS.n7761 2.6005
R6512 VSS.n7766 VSS.n7765 2.6005
R6513 VSS.n7765 VSS.n7764 2.6005
R6514 VSS.n7769 VSS.n7768 2.6005
R6515 VSS.n7768 VSS.n7767 2.6005
R6516 VSS.n7772 VSS.n7771 2.6005
R6517 VSS.n7771 VSS.n7770 2.6005
R6518 VSS.n7775 VSS.n7774 2.6005
R6519 VSS.n7774 VSS.n7773 2.6005
R6520 VSS.n7778 VSS.n7777 2.6005
R6521 VSS.n7777 VSS.n7776 2.6005
R6522 VSS.n7781 VSS.n7780 2.6005
R6523 VSS.n7780 VSS.n7779 2.6005
R6524 VSS.n7785 VSS.n7784 2.6005
R6525 VSS.n7784 VSS.n7783 2.6005
R6526 VSS.n7788 VSS.n7787 2.6005
R6527 VSS.n7787 VSS.n7786 2.6005
R6528 VSS.n7791 VSS.n7790 2.6005
R6529 VSS.n7790 VSS.n7789 2.6005
R6530 VSS.n7796 VSS.n7795 2.6005
R6531 VSS.n7606 VSS.n5318 2.6005
R6532 VSS.n5318 VSS.n5317 2.6005
R6533 VSS.n7604 VSS.n7603 2.6005
R6534 VSS.n7603 VSS.n7602 2.6005
R6535 VSS.n7601 VSS.n7600 2.6005
R6536 VSS.n7600 VSS.n7599 2.6005
R6537 VSS.n7598 VSS.n7597 2.6005
R6538 VSS.n7597 VSS.n7596 2.6005
R6539 VSS.n7594 VSS.n7593 2.6005
R6540 VSS.n7593 VSS.n7592 2.6005
R6541 VSS VSS.n7591 2.6005
R6542 VSS.n7591 VSS.n7590 2.6005
R6543 VSS.n7589 VSS.n7587 2.6005
R6544 VSS.n7589 VSS.n7588 2.6005
R6545 VSS.n7586 VSS.n7585 2.6005
R6546 VSS.n7585 VSS.n7584 2.6005
R6547 VSS.n7583 VSS.n7582 2.6005
R6548 VSS.n7582 VSS.n7581 2.6005
R6549 VSS.n7580 VSS.n7579 2.6005
R6550 VSS.n7579 VSS.n7578 2.6005
R6551 VSS.n7576 VSS.n7575 2.6005
R6552 VSS.n7575 VSS.n7574 2.6005
R6553 VSS.n6924 VSS.n6923 2.6005
R6554 VSS.n6923 VSS.n6922 2.6005
R6555 VSS.n7558 VSS.n7557 2.6005
R6556 VSS.n7557 VSS.n7556 2.6005
R6557 VSS.n7571 VSS.n7570 2.6005
R6558 VSS.n7570 VSS.n7569 2.6005
R6559 VSS.n7629 VSS.n7628 2.6005
R6560 VSS.n7628 VSS.n7627 2.6005
R6561 VSS.n7625 VSS.n7624 2.6005
R6562 VSS.n7624 VSS.n7623 2.6005
R6563 VSS.n5310 VSS.n5309 2.6005
R6564 VSS.n5309 VSS.n5308 2.6005
R6565 VSS.n5313 VSS.n5312 2.6005
R6566 VSS.n5312 VSS.n5311 2.6005
R6567 VSS.n5322 VSS.n5321 2.6005
R6568 VSS.n5321 VSS.n5320 2.6005
R6569 VSS.n5325 VSS.n5324 2.6005
R6570 VSS.n5324 VSS.n5323 2.6005
R6571 VSS.n5328 VSS.n5327 2.6005
R6572 VSS.n5327 VSS.n5326 2.6005
R6573 VSS.n5333 VSS.n5332 2.6005
R6574 VSS.n5332 VSS.n5331 2.6005
R6575 VSS.n5336 VSS.n5335 2.6005
R6576 VSS.n5335 VSS.n5334 2.6005
R6577 VSS.n5339 VSS.n5338 2.6005
R6578 VSS.n5338 VSS.n5337 2.6005
R6579 VSS.n5342 VSS.n5341 2.6005
R6580 VSS.n5341 VSS.n5340 2.6005
R6581 VSS.n7561 VSS.n7560 2.6005
R6582 VSS.n7560 VSS.n7559 2.6005
R6583 VSS.n7564 VSS.n7563 2.6005
R6584 VSS.n7563 VSS.n7562 2.6005
R6585 VSS.n6618 VSS.n6617 2.6005
R6586 VSS.n6617 VSS.n6616 2.6005
R6587 VSS.n7567 VSS.n7566 2.6005
R6588 VSS.n7566 VSS.n7565 2.6005
R6589 VSS.n6912 VSS.n6911 2.6005
R6590 VSS.n6911 VSS.n6910 2.6005
R6591 VSS.n6909 VSS.n6908 2.6005
R6592 VSS.n6908 VSS.n6907 2.6005
R6593 VSS.n6906 VSS.n6905 2.6005
R6594 VSS.n6905 VSS.n6904 2.6005
R6595 VSS.n6903 VSS.n6902 2.6005
R6596 VSS.n6902 VSS.n6901 2.6005
R6597 VSS.n6900 VSS.n6899 2.6005
R6598 VSS.n6899 VSS.n6898 2.6005
R6599 VSS.n6896 VSS.n6895 2.6005
R6600 VSS.n6895 VSS.n6894 2.6005
R6601 VSS.n6893 VSS.n6892 2.6005
R6602 VSS.n6892 VSS.n6891 2.6005
R6603 VSS.n6890 VSS.n6889 2.6005
R6604 VSS.n6889 VSS.n6888 2.6005
R6605 VSS.n6887 VSS.n6886 2.6005
R6606 VSS.n6886 VSS.n6885 2.6005
R6607 VSS.n6884 VSS.n6883 2.6005
R6608 VSS.n6883 VSS.n6882 2.6005
R6609 VSS.n6881 VSS.n6880 2.6005
R6610 VSS.n6880 VSS.n6879 2.6005
R6611 VSS.n6878 VSS.n6877 2.6005
R6612 VSS.n6877 VSS.n6876 2.6005
R6613 VSS.n6875 VSS.n6874 2.6005
R6614 VSS.n6874 VSS.n6873 2.6005
R6615 VSS.n6849 VSS.n6848 2.6005
R6616 VSS.n6848 VSS.n6847 2.6005
R6617 VSS.n6852 VSS.n6851 2.6005
R6618 VSS.n6851 VSS.n6850 2.6005
R6619 VSS.n6855 VSS.n6854 2.6005
R6620 VSS.n6854 VSS.n6853 2.6005
R6621 VSS.n6840 VSS.n6839 2.6005
R6622 VSS.n6842 VSS.n6841 2.6005
R6623 VSS.n6846 VSS.n6845 2.6005
R6624 VSS.n6828 VSS.n6827 2.6005
R6625 VSS.n6827 VSS.n6826 2.6005
R6626 VSS.n6825 VSS.n6824 2.6005
R6627 VSS.n6824 VSS.n6823 2.6005
R6628 VSS.n6831 VSS.n6830 2.6005
R6629 VSS.n6833 VSS.n6832 2.6005
R6630 VSS.n6837 VSS.n6836 2.6005
R6631 VSS.n6804 VSS.n6639 2.6005
R6632 VSS.n6639 VSS.n6638 2.6005
R6633 VSS.n6802 VSS.n6801 2.6005
R6634 VSS.n6801 VSS.n6800 2.6005
R6635 VSS.n6799 VSS.n6798 2.6005
R6636 VSS.n6798 VSS.n6797 2.6005
R6637 VSS.n6796 VSS.n6795 2.6005
R6638 VSS.n6795 VSS.n6794 2.6005
R6639 VSS.n6791 VSS.n6790 2.6005
R6640 VSS.n6790 VSS.n6789 2.6005
R6641 VSS VSS.n6788 2.6005
R6642 VSS.n6788 VSS.n6787 2.6005
R6643 VSS.n6786 VSS.n6784 2.6005
R6644 VSS.n6786 VSS.n6785 2.6005
R6645 VSS.n6783 VSS.n6782 2.6005
R6646 VSS.n6782 VSS.n6781 2.6005
R6647 VSS.n6780 VSS.n6779 2.6005
R6648 VSS.n6779 VSS.n6778 2.6005
R6649 VSS.n6777 VSS.n6776 2.6005
R6650 VSS.n6776 VSS.n6775 2.6005
R6651 VSS.n6773 VSS.n6772 2.6005
R6652 VSS.n6772 VSS.n6771 2.6005
R6653 VSS.n6821 VSS.n6820 2.6005
R6654 VSS.n6820 VSS.n6819 2.6005
R6655 VSS.n6817 VSS.n6816 2.6005
R6656 VSS.n6816 VSS.n6815 2.6005
R6657 VSS.n6814 VSS.n6813 2.6005
R6658 VSS.n6813 VSS.n6812 2.6005
R6659 VSS.n6811 VSS.n6810 2.6005
R6660 VSS.n6810 VSS.n6809 2.6005
R6661 VSS.n6643 VSS.n6642 2.6005
R6662 VSS.n6642 VSS.n6641 2.6005
R6663 VSS.n6646 VSS.n6645 2.6005
R6664 VSS.n6645 VSS.n6644 2.6005
R6665 VSS.n6649 VSS.n6648 2.6005
R6666 VSS.n6648 VSS.n6647 2.6005
R6667 VSS.n6652 VSS.n6651 2.6005
R6668 VSS.n6651 VSS.n6650 2.6005
R6669 VSS.n6655 VSS.n6654 2.6005
R6670 VSS.n6654 VSS.n6653 2.6005
R6671 VSS.n6658 VSS.n6657 2.6005
R6672 VSS.n6657 VSS.n6656 2.6005
R6673 VSS.n6661 VSS.n6660 2.6005
R6674 VSS.n6660 VSS.n6659 2.6005
R6675 VSS.n6668 VSS.n6667 2.6005
R6676 VSS.n6667 VSS.n6666 2.6005
R6677 VSS.n6671 VSS.n6670 2.6005
R6678 VSS.n6670 VSS.n6669 2.6005
R6679 VSS.n6674 VSS.n6673 2.6005
R6680 VSS.n6673 VSS.n6672 2.6005
R6681 VSS.n6677 VSS.n6676 2.6005
R6682 VSS.n6676 VSS.n6675 2.6005
R6683 VSS.n6680 VSS.n6679 2.6005
R6684 VSS.n6679 VSS.n6678 2.6005
R6685 VSS.n6768 VSS.n6767 2.6005
R6686 VSS.n6767 VSS.n6766 2.6005
R6687 VSS.n6765 VSS.n6764 2.6005
R6688 VSS.n6764 VSS.n6763 2.6005
R6689 VSS.n6762 VSS.n6761 2.6005
R6690 VSS.n6761 VSS.n6760 2.6005
R6691 VSS.n6758 VSS.n6757 2.6005
R6692 VSS.n6757 VSS.n6756 2.6005
R6693 VSS.n6755 VSS.n6754 2.6005
R6694 VSS.n6754 VSS.n6753 2.6005
R6695 VSS.n6752 VSS.n6751 2.6005
R6696 VSS.n6736 VSS.n6735 2.6005
R6697 VSS.n6735 VSS.n6734 2.6005
R6698 VSS.n6732 VSS.n6731 2.6005
R6699 VSS.n6731 VSS.n6730 2.6005
R6700 VSS.n6729 VSS.n6728 2.6005
R6701 VSS.n6728 VSS.n6727 2.6005
R6702 VSS.n6967 VSS.n6966 2.6005
R6703 VSS.n6966 VSS.n6965 2.6005
R6704 VSS.n6969 VSS.n6968 2.6005
R6705 VSS.n6970 VSS.n6969 2.6005
R6706 VSS.n6615 VSS.n6614 2.6005
R6707 VSS.n6614 VSS.n6613 2.6005
R6708 VSS.n6688 VSS.n6687 2.6005
R6709 VSS.n6687 VSS.n6686 2.6005
R6710 VSS.n6691 VSS.n6690 2.6005
R6711 VSS.n6690 VSS.n6689 2.6005
R6712 VSS.n6694 VSS.n6693 2.6005
R6713 VSS.n6693 VSS.n6692 2.6005
R6714 VSS.n6699 VSS.n6698 2.6005
R6715 VSS.n6698 VSS.n6697 2.6005
R6716 VSS.n6703 VSS.n6702 2.6005
R6717 VSS.n6705 VSS.n6704 2.6005
R6718 VSS.n6708 VSS.n6707 2.6005
R6719 VSS.n6721 VSS.n6720 2.6005
R6720 VSS.n6723 VSS.n6722 2.6005
R6721 VSS.n6726 VSS.n6725 2.6005
R6722 VSS.n6964 VSS.n6963 2.6005
R6723 VSS.n6962 VSS.n6961 2.6005
R6724 VSS.n6958 VSS.n6957 2.6005
R6725 VSS.n6957 VSS.n6956 2.6005
R6726 VSS.n6955 VSS.n6954 2.6005
R6727 VSS.n6954 VSS.n6953 2.6005
R6728 VSS.n6935 VSS.n6934 2.6005
R6729 VSS.n6934 VSS.n6933 2.6005
R6730 VSS.n6938 VSS.n6937 2.6005
R6731 VSS.n6937 VSS.n6936 2.6005
R6732 VSS.n5354 VSS.n5353 2.6005
R6733 VSS.n5353 VSS.n5352 2.6005
R6734 VSS.n7539 VSS.n7538 2.6005
R6735 VSS.n7538 VSS.n7537 2.6005
R6736 VSS.n7536 VSS.n7535 2.6005
R6737 VSS.n7535 VSS.n7534 2.6005
R6738 VSS.n7533 VSS.n7532 2.6005
R6739 VSS.n7531 VSS.n7530 2.6005
R6740 VSS.n7490 VSS.n7489 2.6005
R6741 VSS.n7489 VSS.n7488 2.6005
R6742 VSS.n7493 VSS.n7492 2.6005
R6743 VSS.n7492 VSS.n7491 2.6005
R6744 VSS.n7496 VSS.n7495 2.6005
R6745 VSS.n7495 VSS.n7494 2.6005
R6746 VSS.n7499 VSS.n7498 2.6005
R6747 VSS.n7498 VSS.n7497 2.6005
R6748 VSS.n7502 VSS.n7501 2.6005
R6749 VSS.n7501 VSS.n7500 2.6005
R6750 VSS.n7505 VSS.n7504 2.6005
R6751 VSS.n7504 VSS.n7503 2.6005
R6752 VSS.n7508 VSS.n7507 2.6005
R6753 VSS.n7507 VSS.n7506 2.6005
R6754 VSS.n7511 VSS.n7510 2.6005
R6755 VSS.n7510 VSS.n7509 2.6005
R6756 VSS.n7514 VSS.n7513 2.6005
R6757 VSS.n7513 VSS.n7512 2.6005
R6758 VSS.n7517 VSS.n7516 2.6005
R6759 VSS.n7516 VSS.n7515 2.6005
R6760 VSS.n7520 VSS.n7519 2.6005
R6761 VSS.n7519 VSS.n7518 2.6005
R6762 VSS.n7524 VSS.n7523 2.6005
R6763 VSS.n7523 VSS.n7522 2.6005
R6764 VSS.n7527 VSS.n7526 2.6005
R6765 VSS.n7526 VSS.n7525 2.6005
R6766 VSS.n5356 VSS.n5355 2.6005
R6767 VSS.n7438 VSS.n7437 2.6005
R6768 VSS.n7437 VSS.n7436 2.6005
R6769 VSS.n7441 VSS.n7440 2.6005
R6770 VSS.n7440 VSS.n7439 2.6005
R6771 VSS.n7444 VSS.n7443 2.6005
R6772 VSS.n7443 VSS.n7442 2.6005
R6773 VSS.n7447 VSS.n7446 2.6005
R6774 VSS.n7446 VSS.n7445 2.6005
R6775 VSS.n7450 VSS.n7449 2.6005
R6776 VSS.n7449 VSS.n7448 2.6005
R6777 VSS.n7453 VSS.n7452 2.6005
R6778 VSS.n7452 VSS.n7451 2.6005
R6779 VSS.n7456 VSS.n7455 2.6005
R6780 VSS.n7455 VSS.n7454 2.6005
R6781 VSS.n7459 VSS.n7458 2.6005
R6782 VSS.n7458 VSS.n7457 2.6005
R6783 VSS.n7462 VSS.n7461 2.6005
R6784 VSS.n7461 VSS.n7460 2.6005
R6785 VSS.n7465 VSS.n7464 2.6005
R6786 VSS.n7464 VSS.n7463 2.6005
R6787 VSS.n7468 VSS.n7467 2.6005
R6788 VSS.n7467 VSS.n7466 2.6005
R6789 VSS.n7471 VSS.n7470 2.6005
R6790 VSS.n7470 VSS.n7469 2.6005
R6791 VSS.n7475 VSS.n7474 2.6005
R6792 VSS.n7474 VSS.n7473 2.6005
R6793 VSS.n7478 VSS.n7477 2.6005
R6794 VSS.n7480 VSS.n7479 2.6005
R6795 VSS.n7483 VSS.n7482 2.6005
R6796 VSS.n7430 VSS.n7429 2.6005
R6797 VSS.n6327 VSS.n6326 2.6005
R6798 VSS.n6324 VSS.n6323 2.6005
R6799 VSS.n6322 VSS.n6321 2.6005
R6800 VSS.n6319 VSS.n6318 2.6005
R6801 VSS.n6317 VSS.n6316 2.6005
R6802 VSS.n6314 VSS.n6313 2.6005
R6803 VSS.n6312 VSS.n6311 2.6005
R6804 VSS.n6309 VSS.n6308 2.6005
R6805 VSS.n6307 VSS.n6306 2.6005
R6806 VSS.n6304 VSS.n6303 2.6005
R6807 VSS.n7434 VSS.n7433 2.6005
R6808 VSS.n5381 VSS.n5380 2.6005
R6809 VSS.n6301 VSS.n6300 2.6005
R6810 VSS.n6299 VSS.n6298 2.6005
R6811 VSS.n6296 VSS.n6295 2.6005
R6812 VSS.n6294 VSS.n6293 2.6005
R6813 VSS.n6291 VSS.n6290 2.6005
R6814 VSS.n6289 VSS.n6288 2.6005
R6815 VSS.n6286 VSS.n6285 2.6005
R6816 VSS.n6284 VSS.n6283 2.6005
R6817 VSS.n6282 VSS.n6281 2.6005
R6818 VSS.n6281 VSS.n6280 2.6005
R6819 VSS.n6279 VSS.n6278 2.6005
R6820 VSS.n6272 VSS.n6271 2.6005
R6821 VSS.n6270 VSS.n6269 2.6005
R6822 VSS.n6266 VSS.n6265 2.6005
R6823 VSS.n6237 VSS.n6236 2.6005
R6824 VSS.n6239 VSS.n6238 2.6005
R6825 VSS.n6242 VSS.n6241 2.6005
R6826 VSS.n6244 VSS.n6243 2.6005
R6827 VSS.n6247 VSS.n6246 2.6005
R6828 VSS.n6249 VSS.n6248 2.6005
R6829 VSS.n6263 VSS.n6262 2.6005
R6830 VSS.n6253 VSS.n6252 2.6005
R6831 VSS.n6255 VSS.n6254 2.6005
R6832 VSS.n6258 VSS.n6257 2.6005
R6833 VSS.n6260 VSS.n6259 2.6005
R6834 VSS.n5950 VSS.n5949 2.6005
R6835 VSS.n6033 VSS.n6032 2.6005
R6836 VSS.n6035 VSS.n6034 2.6005
R6837 VSS.n6037 VSS.n6036 2.6005
R6838 VSS.n6039 VSS.n6038 2.6005
R6839 VSS.n6234 VSS.n6233 2.6005
R6840 VSS.n6231 VSS.n6230 2.6005
R6841 VSS.n6227 VSS.n6226 2.6005
R6842 VSS.n6226 VSS.n6225 2.6005
R6843 VSS.n6045 VSS.n6044 2.6005
R6844 VSS.n6044 VSS.n6043 2.6005
R6845 VSS.n6049 VSS.n6048 2.6005
R6846 VSS.n6048 VSS.n6047 2.6005
R6847 VSS.n6052 VSS.n6051 2.6005
R6848 VSS.n6051 VSS.n6050 2.6005
R6849 VSS.n6056 VSS.n6055 2.6005
R6850 VSS.n6055 VSS.n6054 2.6005
R6851 VSS.n6059 VSS.n6058 2.6005
R6852 VSS.n6058 VSS.n6057 2.6005
R6853 VSS.n6062 VSS.n6061 2.6005
R6854 VSS.n6061 VSS.n6060 2.6005
R6855 VSS.n6065 VSS.n6064 2.6005
R6856 VSS.n6064 VSS.n6063 2.6005
R6857 VSS.n6068 VSS.n6067 2.6005
R6858 VSS.n6067 VSS.n6066 2.6005
R6859 VSS.n6071 VSS.n6070 2.6005
R6860 VSS.n6070 VSS.n6069 2.6005
R6861 VSS.n6074 VSS.n6073 2.6005
R6862 VSS.n6073 VSS.t724 2.6005
R6863 VSS.n6077 VSS.n6076 2.6005
R6864 VSS.n6076 VSS.n6075 2.6005
R6865 VSS.n6080 VSS.n6079 2.6005
R6866 VSS.n6079 VSS.n6078 2.6005
R6867 VSS.n6083 VSS.n6082 2.6005
R6868 VSS.n6082 VSS.n6081 2.6005
R6869 VSS.n6086 VSS.n6085 2.6005
R6870 VSS.n6085 VSS.n6084 2.6005
R6871 VSS.n6090 VSS.n6089 2.6005
R6872 VSS.n6089 VSS.n6088 2.6005
R6873 VSS.n6093 VSS.n6092 2.6005
R6874 VSS.n6092 VSS.n6091 2.6005
R6875 VSS.n6096 VSS.n6095 2.6005
R6876 VSS.n6095 VSS.n6094 2.6005
R6877 VSS.n6099 VSS.n6098 2.6005
R6878 VSS.n6098 VSS.n6097 2.6005
R6879 VSS.n6102 VSS.n6101 2.6005
R6880 VSS.n6101 VSS.n6100 2.6005
R6881 VSS.n6031 VSS.n6030 2.6005
R6882 VSS.n6030 VSS.n6029 2.6005
R6883 VSS.n6028 VSS.n6027 2.6005
R6884 VSS.n6027 VSS.n6026 2.6005
R6885 VSS.n6025 VSS.n6024 2.6005
R6886 VSS.n6024 VSS.n6023 2.6005
R6887 VSS.n6022 VSS.n6021 2.6005
R6888 VSS.n6021 VSS.n6020 2.6005
R6889 VSS.n6019 VSS.n6018 2.6005
R6890 VSS.n6018 VSS.n6017 2.6005
R6891 VSS.n6016 VSS.n6015 2.6005
R6892 VSS.n6015 VSS.n6014 2.6005
R6893 VSS.n6013 VSS.n6012 2.6005
R6894 VSS.n6012 VSS.n6011 2.6005
R6895 VSS.n6010 VSS.n6009 2.6005
R6896 VSS.n6009 VSS.n6008 2.6005
R6897 VSS.n6007 VSS.n6006 2.6005
R6898 VSS.n6006 VSS.n6005 2.6005
R6899 VSS.n6004 VSS.n6003 2.6005
R6900 VSS.n6003 VSS.n6002 2.6005
R6901 VSS.n6001 VSS.n6000 2.6005
R6902 VSS.n6000 VSS.n5999 2.6005
R6903 VSS.n5998 VSS.n5997 2.6005
R6904 VSS.n5997 VSS.n5996 2.6005
R6905 VSS.n5995 VSS.n5994 2.6005
R6906 VSS.n5994 VSS.n5993 2.6005
R6907 VSS.n5992 VSS.n5991 2.6005
R6908 VSS.n5991 VSS.n5990 2.6005
R6909 VSS.n5989 VSS.n5988 2.6005
R6910 VSS.n5988 VSS.n5987 2.6005
R6911 VSS.n5986 VSS.n5985 2.6005
R6912 VSS.n5985 VSS.n5984 2.6005
R6913 VSS.n5983 VSS.n5982 2.6005
R6914 VSS.n5982 VSS.n5981 2.6005
R6915 VSS.n5980 VSS.n5979 2.6005
R6916 VSS.n5979 VSS.n5978 2.6005
R6917 VSS.n5977 VSS.n5976 2.6005
R6918 VSS.n5976 VSS.n5975 2.6005
R6919 VSS.n5974 VSS.n5973 2.6005
R6920 VSS.n5973 VSS.n5972 2.6005
R6921 VSS.n5971 VSS.n5970 2.6005
R6922 VSS.n5970 VSS.n5969 2.6005
R6923 VSS.n5968 VSS.n5967 2.6005
R6924 VSS.n5967 VSS.n5966 2.6005
R6925 VSS.n5965 VSS.n5964 2.6005
R6926 VSS.n5964 VSS.n5963 2.6005
R6927 VSS.n5958 VSS.n5957 2.6005
R6928 VSS.n327 VSS.n326 2.6005
R6929 VSS.n331 VSS.n330 2.6005
R6930 VSS.n335 VSS.n334 2.6005
R6931 VSS.n334 VSS.n333 2.6005
R6932 VSS.n338 VSS.n337 2.6005
R6933 VSS.n337 VSS.n336 2.6005
R6934 VSS.n341 VSS.n340 2.6005
R6935 VSS.n340 VSS.n339 2.6005
R6936 VSS.n344 VSS.n343 2.6005
R6937 VSS.n343 VSS.n342 2.6005
R6938 VSS.n347 VSS.n346 2.6005
R6939 VSS.n346 VSS.n345 2.6005
R6940 VSS.n350 VSS.n349 2.6005
R6941 VSS.n349 VSS.n348 2.6005
R6942 VSS.n353 VSS.n352 2.6005
R6943 VSS.n352 VSS.n351 2.6005
R6944 VSS.n357 VSS.n356 2.6005
R6945 VSS.n356 VSS.n355 2.6005
R6946 VSS.n360 VSS.n359 2.6005
R6947 VSS.n359 VSS.n358 2.6005
R6948 VSS.n363 VSS.n362 2.6005
R6949 VSS.n362 VSS.n361 2.6005
R6950 VSS.n366 VSS.n365 2.6005
R6951 VSS.n365 VSS.n364 2.6005
R6952 VSS.n369 VSS.n368 2.6005
R6953 VSS.n368 VSS.n367 2.6005
R6954 VSS.n372 VSS.n371 2.6005
R6955 VSS.n371 VSS.n370 2.6005
R6956 VSS.n375 VSS.n374 2.6005
R6957 VSS.n374 VSS.n373 2.6005
R6958 VSS.n378 VSS.n377 2.6005
R6959 VSS.n377 VSS.n376 2.6005
R6960 VSS.n494 VSS.n493 2.6005
R6961 VSS.n493 VSS.n492 2.6005
R6962 VSS.n497 VSS.n496 2.6005
R6963 VSS.n496 VSS.n495 2.6005
R6964 VSS.n428 VSS.n427 2.6005
R6965 VSS.n427 VSS.n426 2.6005
R6966 VSS.n431 VSS.n430 2.6005
R6967 VSS.n430 VSS.n429 2.6005
R6968 VSS.n434 VSS.n433 2.6005
R6969 VSS.n433 VSS.n432 2.6005
R6970 VSS.n437 VSS.n436 2.6005
R6971 VSS.n436 VSS.n435 2.6005
R6972 VSS.n440 VSS.n439 2.6005
R6973 VSS.n439 VSS.n438 2.6005
R6974 VSS.n443 VSS.n442 2.6005
R6975 VSS.n442 VSS.n441 2.6005
R6976 VSS.n446 VSS.n445 2.6005
R6977 VSS.n445 VSS.n444 2.6005
R6978 VSS.n449 VSS.n448 2.6005
R6979 VSS.n448 VSS.n447 2.6005
R6980 VSS.n452 VSS.n451 2.6005
R6981 VSS.n451 VSS.n450 2.6005
R6982 VSS.n455 VSS.n454 2.6005
R6983 VSS.n454 VSS.n453 2.6005
R6984 VSS.n458 VSS.n457 2.6005
R6985 VSS.n457 VSS.n456 2.6005
R6986 VSS.n461 VSS.n460 2.6005
R6987 VSS.n460 VSS.n459 2.6005
R6988 VSS.n464 VSS.n463 2.6005
R6989 VSS.n463 VSS.n462 2.6005
R6990 VSS.n467 VSS.n466 2.6005
R6991 VSS.n466 VSS.n465 2.6005
R6992 VSS.n470 VSS.n469 2.6005
R6993 VSS.n469 VSS.n468 2.6005
R6994 VSS.n473 VSS.n472 2.6005
R6995 VSS.n472 VSS.n471 2.6005
R6996 VSS.n476 VSS.n475 2.6005
R6997 VSS.n475 VSS.n474 2.6005
R6998 VSS.n479 VSS.n478 2.6005
R6999 VSS.n478 VSS.n477 2.6005
R7000 VSS.n482 VSS.n481 2.6005
R7001 VSS.n481 VSS.n480 2.6005
R7002 VSS.n485 VSS.n484 2.6005
R7003 VSS.n484 VSS.n483 2.6005
R7004 VSS.n488 VSS.n487 2.6005
R7005 VSS.n487 VSS.n486 2.6005
R7006 VSS.n491 VSS.n490 2.6005
R7007 VSS.n490 VSS.n489 2.6005
R7008 VSS.n422 VSS.n421 2.6005
R7009 VSS.n425 VSS.n424 2.6005
R7010 VSS.n398 VSS.n397 2.6005
R7011 VSS.n397 VSS.n396 2.6005
R7012 VSS.n401 VSS.n400 2.6005
R7013 VSS.n400 VSS.n399 2.6005
R7014 VSS.n404 VSS.n403 2.6005
R7015 VSS.n403 VSS.n402 2.6005
R7016 VSS.n407 VSS.n406 2.6005
R7017 VSS.n406 VSS.n405 2.6005
R7018 VSS.n410 VSS.n409 2.6005
R7019 VSS.n409 VSS.n408 2.6005
R7020 VSS.n413 VSS.n412 2.6005
R7021 VSS.n412 VSS.n411 2.6005
R7022 VSS.n416 VSS.n415 2.6005
R7023 VSS.n415 VSS.n414 2.6005
R7024 VSS.n420 VSS.n419 2.6005
R7025 VSS.n419 VSS.n418 2.6005
R7026 VSS.n381 VSS.n380 2.6005
R7027 VSS.n383 VSS.n382 2.6005
R7028 VSS.n386 VSS.n385 2.6005
R7029 VSS.n389 VSS.n388 2.6005
R7030 VSS.n393 VSS.n392 2.6005
R7031 VSS.n5611 VSS.n5610 2.6005
R7032 VSS.n5610 VSS.n5609 2.6005
R7033 VSS.n5586 VSS.n5585 2.6005
R7034 VSS.n5585 VSS.n5584 2.6005
R7035 VSS.n5589 VSS.n5588 2.6005
R7036 VSS.n5588 VSS.n5587 2.6005
R7037 VSS.n5592 VSS.n5591 2.6005
R7038 VSS.n5591 VSS.n5590 2.6005
R7039 VSS.n5593 VSS.n5578 2.6005
R7040 VSS.n5578 VSS.n5577 2.6005
R7041 VSS.n5595 VSS 2.6005
R7042 VSS.n5595 VSS.n5594 2.6005
R7043 VSS.n5598 VSS.n5597 2.6005
R7044 VSS.n5597 VSS.n5596 2.6005
R7045 VSS.n5601 VSS.n5600 2.6005
R7046 VSS.n5600 VSS.n5599 2.6005
R7047 VSS.n5604 VSS.n5603 2.6005
R7048 VSS.n5603 VSS.n5602 2.6005
R7049 VSS.n5607 VSS.n5606 2.6005
R7050 VSS.n5606 VSS.n5605 2.6005
R7051 VSS.n5582 VSS.n5581 2.6005
R7052 VSS.n5581 VSS.n5580 2.6005
R7053 VSS.n5536 VSS.n5535 2.6005
R7054 VSS.n5535 VSS.n5534 2.6005
R7055 VSS.n5511 VSS.n5510 2.6005
R7056 VSS.n5510 VSS.n5509 2.6005
R7057 VSS.n5514 VSS.n5513 2.6005
R7058 VSS.n5513 VSS.n5512 2.6005
R7059 VSS.n5517 VSS.n5516 2.6005
R7060 VSS.n5516 VSS.n5515 2.6005
R7061 VSS.n5518 VSS.n5503 2.6005
R7062 VSS.n5503 VSS.n5502 2.6005
R7063 VSS.n5520 VSS 2.6005
R7064 VSS.n5520 VSS.n5519 2.6005
R7065 VSS.n5523 VSS.n5522 2.6005
R7066 VSS.n5522 VSS.n5521 2.6005
R7067 VSS.n5526 VSS.n5525 2.6005
R7068 VSS.n5525 VSS.n5524 2.6005
R7069 VSS.n5529 VSS.n5528 2.6005
R7070 VSS.n5528 VSS.n5527 2.6005
R7071 VSS.n5532 VSS.n5531 2.6005
R7072 VSS.n5531 VSS.n5530 2.6005
R7073 VSS.n5507 VSS.n5506 2.6005
R7074 VSS.n5469 VSS.n5468 2.6005
R7075 VSS.n5473 VSS.n5472 2.6005
R7076 VSS.n5472 VSS.n5471 2.6005
R7077 VSS.n5476 VSS.n5475 2.6005
R7078 VSS.n5475 VSS.n5474 2.6005
R7079 VSS.n5479 VSS.n5478 2.6005
R7080 VSS.n5478 VSS.n5477 2.6005
R7081 VSS.n5480 VSS.n5466 2.6005
R7082 VSS.n5466 VSS.n5465 2.6005
R7083 VSS.n5482 VSS 2.6005
R7084 VSS.n5482 VSS.n5481 2.6005
R7085 VSS.n5485 VSS.n5484 2.6005
R7086 VSS.n5484 VSS.n5483 2.6005
R7087 VSS.n5488 VSS.n5487 2.6005
R7088 VSS.n5487 VSS.n5486 2.6005
R7089 VSS.n5491 VSS.n5490 2.6005
R7090 VSS.n5490 VSS.n5489 2.6005
R7091 VSS.n5494 VSS.n5493 2.6005
R7092 VSS.n5493 VSS.n5492 2.6005
R7093 VSS.n5498 VSS.n5497 2.6005
R7094 VSS.n5497 VSS.n5496 2.6005
R7095 VSS.n5541 VSS.n5540 2.6005
R7096 VSS.n5540 VSS.n5539 2.6005
R7097 VSS.n5545 VSS.n5544 2.6005
R7098 VSS.n5544 VSS.n5543 2.6005
R7099 VSS.n5548 VSS.n5547 2.6005
R7100 VSS.n5547 VSS.n5546 2.6005
R7101 VSS.n5551 VSS.n5550 2.6005
R7102 VSS.n5550 VSS.n5549 2.6005
R7103 VSS.n5552 VSS.n5460 2.6005
R7104 VSS.n5460 VSS.n5459 2.6005
R7105 VSS.n5554 VSS 2.6005
R7106 VSS.n5554 VSS.n5553 2.6005
R7107 VSS.n5559 VSS.n5558 2.6005
R7108 VSS.n5558 VSS.n5557 2.6005
R7109 VSS.n5562 VSS.n5561 2.6005
R7110 VSS.n5561 VSS.n5560 2.6005
R7111 VSS.n5565 VSS.n5564 2.6005
R7112 VSS.n5564 VSS.n5563 2.6005
R7113 VSS.n5568 VSS.n5567 2.6005
R7114 VSS.n5567 VSS.n5566 2.6005
R7115 VSS.n5572 VSS.n5571 2.6005
R7116 VSS.n5571 VSS.n5570 2.6005
R7117 VSS.n518 VSS.n517 2.6005
R7118 VSS.n582 VSS.n581 2.6005
R7119 VSS.n581 VSS.n580 2.6005
R7120 VSS.n585 VSS.n584 2.6005
R7121 VSS.n584 VSS.n583 2.6005
R7122 VSS.n588 VSS.n587 2.6005
R7123 VSS.n587 VSS.n586 2.6005
R7124 VSS.n591 VSS.n590 2.6005
R7125 VSS.n590 VSS.n589 2.6005
R7126 VSS.n594 VSS.n593 2.6005
R7127 VSS.n593 VSS.n592 2.6005
R7128 VSS.n75 VSS.n74 2.6005
R7129 VSS.n74 VSS.n73 2.6005
R7130 VSS.n578 VSS.n577 2.6005
R7131 VSS.n577 VSS.n576 2.6005
R7132 VSS.n566 VSS.n565 2.6005
R7133 VSS.n565 VSS.n564 2.6005
R7134 VSS.n569 VSS.n568 2.6005
R7135 VSS.n568 VSS.n567 2.6005
R7136 VSS.n572 VSS.n571 2.6005
R7137 VSS.n571 VSS.n570 2.6005
R7138 VSS.n575 VSS.n574 2.6005
R7139 VSS.n574 VSS.n573 2.6005
R7140 VSS.n562 VSS.n561 2.6005
R7141 VSS.n561 VSS.n560 2.6005
R7142 VSS.n540 VSS.n539 2.6005
R7143 VSS.n539 VSS.n538 2.6005
R7144 VSS.n537 VSS.n536 2.6005
R7145 VSS.n536 VSS.n535 2.6005
R7146 VSS.n534 VSS.n533 2.6005
R7147 VSS.n533 VSS.n532 2.6005
R7148 VSS.n531 VSS.n530 2.6005
R7149 VSS.n530 VSS.n529 2.6005
R7150 VSS.n320 VSS.n319 2.6005
R7151 VSS.n323 VSS.n322 2.6005
R7152 VSS.n527 VSS.n526 2.6005
R7153 VSS.n526 VSS.n525 2.6005
R7154 VSS.n524 VSS.n523 2.6005
R7155 VSS.n523 VSS.n522 2.6005
R7156 VSS.n521 VSS.n520 2.6005
R7157 VSS.n520 VSS.n519 2.6005
R7158 VSS.n500 VSS.n499 2.6005
R7159 VSS.n502 VSS.n501 2.6005
R7160 VSS.n505 VSS.n504 2.6005
R7161 VSS.n508 VSS.n507 2.6005
R7162 VSS.n512 VSS.n511 2.6005
R7163 VSS.n514 VSS.n513 2.6005
R7164 VSS.n284 VSS.n283 2.6005
R7165 VSS.n672 VSS.n671 2.6005
R7166 VSS.n671 VSS.n670 2.6005
R7167 VSS.n610 VSS.n609 2.6005
R7168 VSS.n609 VSS.n608 2.6005
R7169 VSS.n616 VSS.n615 2.6005
R7170 VSS.n615 VSS.n614 2.6005
R7171 VSS.n622 VSS.n621 2.6005
R7172 VSS.n621 VSS.n620 2.6005
R7173 VSS.n628 VSS.n627 2.6005
R7174 VSS.n627 VSS.n626 2.6005
R7175 VSS.n647 VSS 2.6005
R7176 VSS.n647 VSS.n646 2.6005
R7177 VSS.n650 VSS.n649 2.6005
R7178 VSS.n649 VSS.n648 2.6005
R7179 VSS.n656 VSS.n655 2.6005
R7180 VSS.n655 VSS.n654 2.6005
R7181 VSS.n663 VSS.n662 2.6005
R7182 VSS.n662 VSS.n661 2.6005
R7183 VSS.n679 VSS.n678 2.6005
R7184 VSS.n678 VSS.n677 2.6005
R7185 VSS.n603 VSS.n602 2.6005
R7186 VSS.n660 VSS.n659 2.6005
R7187 VSS.n659 VSS.n658 2.6005
R7188 VSS.n666 VSS.n665 2.6005
R7189 VSS.n665 VSS.n664 2.6005
R7190 VSS.n676 VSS.n675 2.6005
R7191 VSS.n675 VSS.n674 2.6005
R7192 VSS.n669 VSS.n668 2.6005
R7193 VSS.n644 VSS.n641 2.6005
R7194 VSS.n606 VSS.n605 2.6005
R7195 VSS.n605 VSS.n604 2.6005
R7196 VSS.n613 VSS.n612 2.6005
R7197 VSS.n612 VSS.n611 2.6005
R7198 VSS.n619 VSS.n618 2.6005
R7199 VSS.n618 VSS.n617 2.6005
R7200 VSS.n625 VSS.n624 2.6005
R7201 VSS.n624 VSS.n623 2.6005
R7202 VSS.n638 VSS.n637 2.6005
R7203 VSS VSS.n644 2.6005
R7204 VSS.n653 VSS.n652 2.6005
R7205 VSS.n652 VSS.n651 2.6005
R7206 VSS.n218 VSS.n217 2.6005
R7207 VSS.n158 VSS.n155 2.6005
R7208 VSS.n159 VSS.n158 2.6005
R7209 VSS.n4583 VSS.n4582 2.6005
R7210 VSS.n4582 VSS.n4581 2.6005
R7211 VSS.n4569 VSS.n4568 2.6005
R7212 VSS.n4543 VSS 2.6005
R7213 VSS.n4543 VSS.n4542 2.6005
R7214 VSS.n4573 VSS.n4572 2.6005
R7215 VSS.n4572 VSS.n4571 2.6005
R7216 VSS.n4586 VSS.n4585 2.6005
R7217 VSS.n4590 VSS.n4589 2.6005
R7218 VSS.n4589 VSS.n4588 2.6005
R7219 VSS.n4529 VSS.n4528 2.6005
R7220 VSS.n4532 VSS.n4531 2.6005
R7221 VSS.n4534 VSS.n4533 2.6005
R7222 VSS.n4548 VSS.n4547 2.6005
R7223 VSS.n4547 VSS.n4546 2.6005
R7224 VSS.n4658 VSS.n4657 2.6005
R7225 VSS.n713 VSS.n712 2.6005
R7226 VSS.n711 VSS.n710 2.6005
R7227 VSS.n708 VSS.n707 2.6005
R7228 VSS.n706 VSS.n705 2.6005
R7229 VSS.n704 VSS.n703 2.6005
R7230 VSS.n702 VSS.n701 2.6005
R7231 VSS.n700 VSS.n699 2.6005
R7232 VSS.n699 VSS.n698 2.6005
R7233 VSS.n4612 VSS.n4611 2.6005
R7234 VSS.n4611 VSS.n4610 2.6005
R7235 VSS.n4615 VSS.n4614 2.6005
R7236 VSS.n4614 VSS.n4613 2.6005
R7237 VSS.n4618 VSS.n4617 2.6005
R7238 VSS.n4617 VSS.n4616 2.6005
R7239 VSS.n4643 VSS.n4642 2.6005
R7240 VSS.n4642 VSS.n4641 2.6005
R7241 VSS.n4646 VSS.n4645 2.6005
R7242 VSS.n4645 VSS.n4644 2.6005
R7243 VSS.n4649 VSS.n4648 2.6005
R7244 VSS.n4648 VSS.n4647 2.6005
R7245 VSS.n4652 VSS.n4651 2.6005
R7246 VSS.n4651 VSS.n4650 2.6005
R7247 VSS.n4655 VSS.n4654 2.6005
R7248 VSS.n4654 VSS.n4653 2.6005
R7249 VSS.n4657 VSS.n4656 2.6005
R7250 VSS.n98 VSS.n97 2.6005
R7251 VSS.n97 VSS.n96 2.6005
R7252 VSS.n101 VSS.n100 2.6005
R7253 VSS.n100 VSS.n99 2.6005
R7254 VSS.n104 VSS.n103 2.6005
R7255 VSS.n103 VSS.n102 2.6005
R7256 VSS.n107 VSS.n106 2.6005
R7257 VSS.n106 VSS.n105 2.6005
R7258 VSS.n110 VSS.n109 2.6005
R7259 VSS.n109 VSS.n108 2.6005
R7260 VSS.n113 VSS.n112 2.6005
R7261 VSS.n112 VSS.n111 2.6005
R7262 VSS.n116 VSS.n115 2.6005
R7263 VSS.n115 VSS.n114 2.6005
R7264 VSS.n120 VSS.n119 2.6005
R7265 VSS.n119 VSS.n118 2.6005
R7266 VSS.n123 VSS.n122 2.6005
R7267 VSS.n122 VSS.n121 2.6005
R7268 VSS.n126 VSS.n125 2.6005
R7269 VSS.n125 VSS.n124 2.6005
R7270 VSS.n129 VSS.n128 2.6005
R7271 VSS.n128 VSS.n127 2.6005
R7272 VSS.n132 VSS.n131 2.6005
R7273 VSS.n131 VSS.n130 2.6005
R7274 VSS.n135 VSS.n134 2.6005
R7275 VSS.n134 VSS.n133 2.6005
R7276 VSS.n78 VSS.n77 2.6005
R7277 VSS.n77 VSS.n76 2.6005
R7278 VSS.n230 VSS.n229 2.6005
R7279 VSS.n229 VSS.n228 2.6005
R7280 VSS.n233 VSS.n232 2.6005
R7281 VSS.n232 VSS.n231 2.6005
R7282 VSS.n236 VSS.n235 2.6005
R7283 VSS.n235 VSS.n234 2.6005
R7284 VSS.n241 VSS.n240 2.6005
R7285 VSS.n240 VSS.n239 2.6005
R7286 VSS.n244 VSS.n243 2.6005
R7287 VSS.n243 VSS.n242 2.6005
R7288 VSS.n247 VSS.n246 2.6005
R7289 VSS.n246 VSS.n245 2.6005
R7290 VSS.n250 VSS.n249 2.6005
R7291 VSS.n249 VSS.n248 2.6005
R7292 VSS.n253 VSS.n252 2.6005
R7293 VSS.n252 VSS.n251 2.6005
R7294 VSS.n256 VSS.n255 2.6005
R7295 VSS.n255 VSS.n254 2.6005
R7296 VSS.n259 VSS.n258 2.6005
R7297 VSS.n258 VSS.n257 2.6005
R7298 VSS.n262 VSS.n261 2.6005
R7299 VSS.n261 VSS.n260 2.6005
R7300 VSS.n265 VSS.n264 2.6005
R7301 VSS.n264 VSS.n263 2.6005
R7302 VSS.n268 VSS.n267 2.6005
R7303 VSS.n267 VSS.n266 2.6005
R7304 VSS.n272 VSS.n271 2.6005
R7305 VSS.n271 VSS.n270 2.6005
R7306 VSS.n275 VSS.n274 2.6005
R7307 VSS.n274 VSS.n273 2.6005
R7308 VSS.n278 VSS.n277 2.6005
R7309 VSS.n277 VSS.n276 2.6005
R7310 VSS.n287 VSS.n286 2.6005
R7311 VSS.n286 VSS.n285 2.6005
R7312 VSS.n290 VSS.n289 2.6005
R7313 VSS.n289 VSS.n288 2.6005
R7314 VSS.n293 VSS.n292 2.6005
R7315 VSS.n292 VSS.n291 2.6005
R7316 VSS.n296 VSS.n295 2.6005
R7317 VSS.n295 VSS.n294 2.6005
R7318 VSS.n299 VSS.n298 2.6005
R7319 VSS.n298 VSS.n297 2.6005
R7320 VSS.n301 VSS.n300 2.6005
R7321 VSS.n305 VSS.n304 2.6005
R7322 VSS.n307 VSS.n306 2.6005
R7323 VSS.n72 VSS.n71 2.6005
R7324 VSS.n71 VSS.n70 2.6005
R7325 VSS.n65 VSS.n64 2.6005
R7326 VSS.n64 VSS.n63 2.6005
R7327 VSS.n62 VSS.n61 2.6005
R7328 VSS.n61 VSS.n60 2.6005
R7329 VSS.n59 VSS.n58 2.6005
R7330 VSS.n58 VSS.n57 2.6005
R7331 VSS.n56 VSS.n55 2.6005
R7332 VSS.n55 VSS.n54 2.6005
R7333 VSS.n543 VSS.n542 2.6005
R7334 VSS.n542 VSS.n541 2.6005
R7335 VSS.n559 VSS.n558 2.6005
R7336 VSS.n558 VSS.n557 2.6005
R7337 VSS.n555 VSS.n554 2.6005
R7338 VSS.n554 VSS.n553 2.6005
R7339 VSS.n552 VSS.n551 2.6005
R7340 VSS.n551 VSS.n550 2.6005
R7341 VSS.n549 VSS.n548 2.6005
R7342 VSS.n548 VSS.n547 2.6005
R7343 VSS.n546 VSS.n545 2.6005
R7344 VSS.n545 VSS.n544 2.6005
R7345 VSS.n314 VSS.n313 2.6005
R7346 VSS.n311 VSS.n310 2.6005
R7347 VSS.n310 VSS.n309 2.6005
R7348 VSS.n316 VSS.n315 2.6005
R7349 VSS.n4666 VSS.n4665 2.6005
R7350 VSS.n4668 VSS.n4667 2.6005
R7351 VSS.n4671 VSS.n4670 2.6005
R7352 VSS.n4674 VSS.n4673 2.6005
R7353 VSS.n4673 VSS.n4672 2.6005
R7354 VSS.n4686 VSS.n4685 2.6005
R7355 VSS.n4685 VSS.n4684 2.6005
R7356 VSS.n4683 VSS.n4682 2.6005
R7357 VSS.n4682 VSS.n4681 2.6005
R7358 VSS.n4680 VSS.n4679 2.6005
R7359 VSS.n4679 VSS.n4678 2.6005
R7360 VSS.n4677 VSS.n4676 2.6005
R7361 VSS.n4676 VSS.n4675 2.6005
R7362 VSS.n68 VSS.n67 2.6005
R7363 VSS.n67 VSS.n66 2.6005
R7364 VSS.n4689 VSS.n4688 2.6005
R7365 VSS.n4700 VSS.n4699 2.6005
R7366 VSS.n4695 VSS.n4694 2.6005
R7367 VSS.n4722 VSS.n4721 2.6005
R7368 VSS.n4737 VSS.n4736 2.6005
R7369 VSS.n4733 VSS.n4732 2.6005
R7370 VSS.n4731 VSS.n4730 2.6005
R7371 VSS.n4728 VSS.n4727 2.6005
R7372 VSS.n4725 VSS.n4724 2.6005
R7373 VSS.n4718 VSS.n4717 2.6005
R7374 VSS.n4703 VSS.n4702 2.6005
R7375 VSS.n4707 VSS.n4706 2.6005
R7376 VSS.n4709 VSS.n4708 2.6005
R7377 VSS.n4712 VSS.n4711 2.6005
R7378 VSS.n4715 VSS.n4714 2.6005
R7379 VSS.n1265 VSS.n1264 2.6005
R7380 VSS.n1266 VSS.n1265 2.6005
R7381 VSS.n1269 VSS.n1268 2.6005
R7382 VSS.n1268 VSS.n1267 2.6005
R7383 VSS.n1272 VSS.n1271 2.6005
R7384 VSS.n1271 VSS.n1270 2.6005
R7385 VSS.n1275 VSS.n1274 2.6005
R7386 VSS.n1274 VSS.n1273 2.6005
R7387 VSS.n1278 VSS.n1277 2.6005
R7388 VSS.n1277 VSS.n1276 2.6005
R7389 VSS.n1281 VSS.n1280 2.6005
R7390 VSS.n1280 VSS.n1279 2.6005
R7391 VSS.n1284 VSS.n1283 2.6005
R7392 VSS.n1283 VSS.n1282 2.6005
R7393 VSS.n1487 VSS.n1484 2.6005
R7394 VSS.n1461 VSS.n1460 2.6005
R7395 VSS.n1460 VSS.n1459 2.6005
R7396 VSS.n1604 VSS.n1601 2.6005
R7397 VSS.n4391 VSS.n4388 2.6005
R7398 VSS.n4401 VSS.n4398 2.6005
R7399 VSS.n4414 VSS.n4412 2.6005
R7400 VSS.n4369 VSS.n4368 2.6005
R7401 VSS.n4368 VSS.n4367 2.6005
R7402 VSS.n4373 VSS.n4372 2.6005
R7403 VSS.n4372 VSS.n4371 2.6005
R7404 VSS.n4419 VSS.n4418 2.6005
R7405 VSS.n4418 VSS.n4417 2.6005
R7406 VSS.n4415 VSS.n4414 2.6005
R7407 VSS.n4408 VSS.n4407 2.6005
R7408 VSS.n4407 VSS.n4406 2.6005
R7409 VSS VSS.n4401 2.6005
R7410 VSS.n4396 VSS.n4395 2.6005
R7411 VSS.n4395 VSS.n4394 2.6005
R7412 VSS.n4392 VSS.n4391 2.6005
R7413 VSS.n4382 VSS.n4381 2.6005
R7414 VSS.n4381 VSS.n4380 2.6005
R7415 VSS.n1605 VSS.n1604 2.6005
R7416 VSS.n1453 VSS.n1452 2.6005
R7417 VSS.n1449 VSS.n1448 2.6005
R7418 VSS.n1446 VSS.n1445 2.6005
R7419 VSS.n1443 VSS.n1442 2.6005
R7420 VSS.n1440 VSS.n1439 2.6005
R7421 VSS.n1437 VSS.n1436 2.6005
R7422 VSS.n1434 VSS.n1433 2.6005
R7423 VSS.n1431 VSS.n1430 2.6005
R7424 VSS.n1428 VSS.n1427 2.6005
R7425 VSS.n1425 VSS.n1424 2.6005
R7426 VSS.n1422 VSS.n1421 2.6005
R7427 VSS.n1256 VSS.n1255 2.6005
R7428 VSS.n1259 VSS.n1258 2.6005
R7429 VSS.n1258 VSS.n1257 2.6005
R7430 VSS.n1263 VSS.n1262 2.6005
R7431 VSS.n1262 VSS.n1261 2.6005
R7432 VSS.n1455 VSS.n1454 2.6005
R7433 VSS.n4432 VSS.n4431 2.6005
R7434 VSS.n4431 VSS.n4430 2.6005
R7435 VSS.n4435 VSS.n4434 2.6005
R7436 VSS.n4434 VSS.n4433 2.6005
R7437 VSS.n4438 VSS.n4437 2.6005
R7438 VSS.n4437 VSS.n4436 2.6005
R7439 VSS.n4442 VSS.n4441 2.6005
R7440 VSS.n4441 VSS.n4440 2.6005
R7441 VSS.n4446 VSS.n4445 2.6005
R7442 VSS.n4445 VSS.n4444 2.6005
R7443 VSS.n4449 VSS.n4448 2.6005
R7444 VSS.n4448 VSS.n4447 2.6005
R7445 VSS.n4452 VSS.n4451 2.6005
R7446 VSS.n4451 VSS.n4450 2.6005
R7447 VSS.n1483 VSS.n1482 2.6005
R7448 VSS.n4456 VSS.n4455 2.6005
R7449 VSS.n4455 VSS.n4454 2.6005
R7450 VSS.n4428 VSS.n4427 2.6005
R7451 VSS.n4426 VSS.n4425 2.6005
R7452 VSS.n4365 VSS.n4364 2.6005
R7453 VSS.n4363 VSS.n4362 2.6005
R7454 VSS.n1458 VSS.n1457 2.6005
R7455 VSS.n1457 VSS.n1456 2.6005
R7456 VSS.n4149 VSS.n4148 2.6005
R7457 VSS.n4148 VSS.n4147 2.6005
R7458 VSS.n4152 VSS.n4151 2.6005
R7459 VSS.n4151 VSS.n4150 2.6005
R7460 VSS.n4361 VSS.n4360 2.6005
R7461 VSS.n4360 VSS.n4359 2.6005
R7462 VSS.n4354 VSS.n4353 2.6005
R7463 VSS.n4353 VSS.n4352 2.6005
R7464 VSS.n4351 VSS.n4350 2.6005
R7465 VSS.n4350 VSS.n4349 2.6005
R7466 VSS.n4343 VSS.n4342 2.6005
R7467 VSS.n4345 VSS.n4344 2.6005
R7468 VSS.n4195 VSS.n4194 2.6005
R7469 VSS.n4194 VSS.n4193 2.6005
R7470 VSS.n4192 VSS.n4191 2.6005
R7471 VSS.n4191 VSS.n4190 2.6005
R7472 VSS.n4189 VSS.n4188 2.6005
R7473 VSS.n4188 VSS.n4187 2.6005
R7474 VSS.n4186 VSS.n4185 2.6005
R7475 VSS.n4185 VSS.n4184 2.6005
R7476 VSS.n4183 VSS.n4182 2.6005
R7477 VSS.n4182 VSS.n4181 2.6005
R7478 VSS.n4180 VSS.n4179 2.6005
R7479 VSS.n4179 VSS.n4178 2.6005
R7480 VSS.n4177 VSS.n4176 2.6005
R7481 VSS.n4176 VSS.n4175 2.6005
R7482 VSS.n4174 VSS.n4173 2.6005
R7483 VSS.n4173 VSS.n4172 2.6005
R7484 VSS.n4168 VSS.n4167 2.6005
R7485 VSS.n4167 VSS.n4166 2.6005
R7486 VSS.n4165 VSS.n4164 2.6005
R7487 VSS.n4164 VSS.n4163 2.6005
R7488 VSS.n4162 VSS.n4161 2.6005
R7489 VSS.n4161 VSS.n4160 2.6005
R7490 VSS.n4159 VSS.n4158 2.6005
R7491 VSS.n4158 VSS.n4157 2.6005
R7492 VSS.n4133 VSS.n4132 2.6005
R7493 VSS.n4135 VSS.n4134 2.6005
R7494 VSS.n4139 VSS.n4138 2.6005
R7495 VSS.n4138 VSS.n4137 2.6005
R7496 VSS.n4141 VSS.n4140 2.6005
R7497 VSS.n95 VSS.n94 2.6005
R7498 VSS.n4145 VSS.n4144 2.6005
R7499 VSS.n4155 VSS.n4154 2.6005
R7500 VSS.n4154 VSS.n4153 2.6005
R7501 VSS.n1565 VSS.n1561 2.6005
R7502 VSS.n1561 VSS.n1560 2.6005
R7503 VSS.n1512 VSS.n1511 2.6005
R7504 VSS.n1511 VSS.n1510 2.6005
R7505 VSS.n1518 VSS.n1517 2.6005
R7506 VSS.n1517 VSS.n1516 2.6005
R7507 VSS.n1524 VSS.n1523 2.6005
R7508 VSS.n1523 VSS.n1522 2.6005
R7509 VSS.n1542 VSS.n1540 2.6005
R7510 VSS.n1542 VSS.n1541 2.6005
R7511 VSS VSS.n1544 2.6005
R7512 VSS.n1544 VSS.n1543 2.6005
R7513 VSS.n1556 VSS.n1555 2.6005
R7514 VSS.n1555 VSS.n1554 2.6005
R7515 VSS.n1584 VSS.n1583 2.6005
R7516 VSS.n1583 VSS.n1582 2.6005
R7517 VSS.n1578 VSS.n1577 2.6005
R7518 VSS.n1577 VSS.n1576 2.6005
R7519 VSS.n1572 VSS.n1571 2.6005
R7520 VSS.n1571 VSS.n1570 2.6005
R7521 VSS.n1505 VSS.n1504 2.6005
R7522 VSS VSS.n1552 2.6005
R7523 VSS.n1552 VSS.n1551 2.6005
R7524 VSS.n1559 VSS.n1558 2.6005
R7525 VSS.n1558 VSS.n1557 2.6005
R7526 VSS.n1581 VSS.n1580 2.6005
R7527 VSS.n1580 VSS.n1579 2.6005
R7528 VSS.n1575 VSS.n1574 2.6005
R7529 VSS.n1574 VSS.n1573 2.6005
R7530 VSS.n1569 VSS.n1568 2.6005
R7531 VSS.n1568 VSS.n1567 2.6005
R7532 VSS.n1564 VSS.n1563 2.6005
R7533 VSS.n1508 VSS.n1507 2.6005
R7534 VSS.n1507 VSS.n1506 2.6005
R7535 VSS.n1515 VSS.n1514 2.6005
R7536 VSS.n1514 VSS.n1513 2.6005
R7537 VSS.n1521 VSS.n1520 2.6005
R7538 VSS.n1520 VSS.n1519 2.6005
R7539 VSS.n1527 VSS.n1526 2.6005
R7540 VSS.n1526 VSS.n1525 2.6005
R7541 VSS.n1548 VSS.n1546 2.6005
R7542 VSS.n1548 VSS.n1547 2.6005
R7543 VSS.n1464 VSS.n1463 2.6005
R7544 VSS.n1463 VSS.n1462 2.6005
R7545 VSS.n1468 VSS.n1467 2.6005
R7546 VSS.n1467 VSS.n1466 2.6005
R7547 VSS.n1471 VSS.n1470 2.6005
R7548 VSS.n1470 VSS.n1469 2.6005
R7549 VSS.n1475 VSS.n1474 2.6005
R7550 VSS.n1474 VSS.n1473 2.6005
R7551 VSS.n4485 VSS.n4484 2.6005
R7552 VSS.n4484 VSS.n4483 2.6005
R7553 VSS.n4488 VSS.n4487 2.6005
R7554 VSS.n4487 VSS.n4486 2.6005
R7555 VSS.n4506 VSS.n4490 2.6005
R7556 VSS.n4490 VSS.n4489 2.6005
R7557 VSS.n4503 VSS.n4502 2.6005
R7558 VSS.n4459 VSS.n4458 2.6005
R7559 VSS.n4458 VSS.n4457 2.6005
R7560 VSS.n4473 VSS.n4472 2.6005
R7561 VSS.n4474 VSS.n4473 2.6005
R7562 VSS.n4471 VSS.n4470 2.6005
R7563 VSS.n4470 VSS.n4469 2.6005
R7564 VSS.n4468 VSS.n4467 2.6005
R7565 VSS.n4467 VSS.n4466 2.6005
R7566 VSS.n4465 VSS.n4464 2.6005
R7567 VSS.n4464 VSS.n4463 2.6005
R7568 VSS.n4462 VSS.n4461 2.6005
R7569 VSS.n4461 VSS.n4460 2.6005
R7570 VSS.n4500 VSS.n4492 2.6005
R7571 VSS.n4492 VSS.n4491 2.6005
R7572 VSS.n4495 VSS.n4494 2.6005
R7573 VSS.n1288 VSS.n1287 2.6005
R7574 VSS.n1287 VSS.n1286 2.6005
R7575 VSS.n1291 VSS.n1290 2.6005
R7576 VSS.n1290 VSS.n1289 2.6005
R7577 VSS.n1294 VSS.n1293 2.6005
R7578 VSS.n1293 VSS.n1292 2.6005
R7579 VSS.n1297 VSS.n1296 2.6005
R7580 VSS.n1296 VSS.n1295 2.6005
R7581 VSS.n1300 VSS.n1299 2.6005
R7582 VSS.n1299 VSS.n1298 2.6005
R7583 VSS.n1303 VSS.n1302 2.6005
R7584 VSS.n1302 VSS.n1301 2.6005
R7585 VSS.n1306 VSS.n1305 2.6005
R7586 VSS.n1305 VSS.n1304 2.6005
R7587 VSS.n1309 VSS.n1308 2.6005
R7588 VSS.n1308 VSS.n1307 2.6005
R7589 VSS.n1313 VSS.n1312 2.6005
R7590 VSS.n1312 VSS.n1311 2.6005
R7591 VSS.n1316 VSS.n1315 2.6005
R7592 VSS.n1315 VSS.n1314 2.6005
R7593 VSS.n1319 VSS.n1318 2.6005
R7594 VSS.n1318 VSS.n1317 2.6005
R7595 VSS.n1322 VSS.n1321 2.6005
R7596 VSS.n1321 VSS.n1320 2.6005
R7597 VSS.n1325 VSS.n1324 2.6005
R7598 VSS.n1324 VSS.n1323 2.6005
R7599 VSS.n1328 VSS.n1327 2.6005
R7600 VSS.n1327 VSS.n1326 2.6005
R7601 VSS.n1331 VSS.n1330 2.6005
R7602 VSS.n1330 VSS.n1329 2.6005
R7603 VSS.n1334 VSS.n1333 2.6005
R7604 VSS.n1333 VSS.n1332 2.6005
R7605 VSS.n1387 VSS.n1386 2.6005
R7606 VSS.n1384 VSS.n1383 2.6005
R7607 VSS.n1381 VSS.n1380 2.6005
R7608 VSS.n4620 VSS.n4619 2.6005
R7609 VSS.n4623 VSS.n4622 2.6005
R7610 VSS.n4625 VSS.n4624 2.6005
R7611 VSS.n4629 VSS.n4628 2.6005
R7612 VSS.n1370 VSS.n1369 2.6005
R7613 VSS.n1377 VSS.n1376 2.6005
R7614 VSS.n1376 VSS.n1375 2.6005
R7615 VSS.n1373 VSS.n1372 2.6005
R7616 VSS.n1372 VSS.n1371 2.6005
R7617 VSS.n1336 VSS.n1335 2.6005
R7618 VSS.n1335 VSS.t147 2.6005
R7619 VSS.n1339 VSS.n1338 2.6005
R7620 VSS.n1338 VSS.n1337 2.6005
R7621 VSS.n1342 VSS.n1341 2.6005
R7622 VSS.n1344 VSS.n1343 2.6005
R7623 VSS.n1347 VSS.n1346 2.6005
R7624 VSS.n1349 VSS.n1348 2.6005
R7625 VSS.n1352 VSS.n1351 2.6005
R7626 VSS.n1354 VSS.n1353 2.6005
R7627 VSS.n1357 VSS.n1356 2.6005
R7628 VSS.n1359 VSS.n1358 2.6005
R7629 VSS.n1362 VSS.n1361 2.6005
R7630 VSS.n1364 VSS.n1363 2.6005
R7631 VSS.n1365 VSS.n782 2.6005
R7632 VSS.n4632 VSS.n4631 2.6005
R7633 VSS.n4631 VSS.n4630 2.6005
R7634 VSS.n4635 VSS.n4634 2.6005
R7635 VSS.n4634 VSS.n4633 2.6005
R7636 VSS.n4639 VSS.n4638 2.6005
R7637 VSS.n4638 VSS.n4637 2.6005
R7638 VSS.n1368 VSS.n1367 2.6005
R7639 VSS.n30 VSS.n29 2.6005
R7640 VSS.n784 VSS.n783 2.6005
R7641 VSS.n788 VSS.n787 2.6005
R7642 VSS.n4742 VSS.n4741 2.6005
R7643 VSS.n4739 VSS.n4738 2.6005
R7644 VSS.n7857 VSS.n7856 2.6005
R7645 VSS.n7860 VSS.n7859 2.6005
R7646 VSS.n7863 VSS.n7862 2.6005
R7647 VSS.n7866 VSS.n7865 2.6005
R7648 VSS.n7871 VSS.n7870 2.6005
R7649 VSS.n4796 VSS.n4795 2.6005
R7650 VSS.n4793 VSS.n4792 2.6005
R7651 VSS.n4791 VSS.n4790 2.6005
R7652 VSS.n5107 VSS.n5106 2.6005
R7653 VSS.n5111 VSS.n5110 2.6005
R7654 VSS.n5116 VSS.n5115 2.6005
R7655 VSS.n5114 VSS.n5113 2.6005
R7656 VSS.n5121 VSS.n5120 2.6005
R7657 VSS.n4782 VSS.n4781 2.6005
R7658 VSS.n4787 VSS.n4786 2.6005
R7659 VSS.n6857 VSS.n6856 2.6005
R7660 VSS.n6860 VSS.n6859 2.6005
R7661 VSS.n6862 VSS.n6861 2.6005
R7662 VSS.n6872 VSS.n6871 2.6005
R7663 VSS.n6871 VSS.n6870 2.6005
R7664 VSS.n6869 VSS.n6868 2.6005
R7665 VSS.n6868 VSS.n6867 2.6005
R7666 VSS.n6866 VSS.n6865 2.6005
R7667 VSS.n5295 VSS.n5294 2.6005
R7668 VSS.n7636 VSS.n7635 2.6005
R7669 VSS.n7638 VSS.n7637 2.6005
R7670 VSS.n7641 VSS.n7640 2.6005
R7671 VSS.n7643 VSS.n7642 2.6005
R7672 VSS.n7646 VSS.n7645 2.6005
R7673 VSS.n7648 VSS.n7647 2.6005
R7674 VSS.n7651 VSS.n7650 2.6005
R7675 VSS.n7653 VSS.n7652 2.6005
R7676 VSS.n7656 VSS.n7655 2.6005
R7677 VSS.n7658 VSS.n7657 2.6005
R7678 VSS.n7661 VSS.n7660 2.6005
R7679 VSS.n7663 VSS.n7662 2.6005
R7680 VSS.n7674 VSS.n7673 2.6005
R7681 VSS.n7673 VSS.n7672 2.6005
R7682 VSS.n7671 VSS.n7670 2.6005
R7683 VSS.n7670 VSS.n7669 2.6005
R7684 VSS.n7667 VSS.n7666 2.6005
R7685 VSS.n5298 VSS.n5297 2.6005
R7686 VSS.n5297 VSS.n5296 2.6005
R7687 VSS.n5293 VSS.n5292 2.6005
R7688 VSS.n5292 VSS.n5291 2.6005
R7689 VSS.n5290 VSS.n5289 2.6005
R7690 VSS.n5289 VSS.n5288 2.6005
R7691 VSS.n5287 VSS.n5286 2.6005
R7692 VSS.n5286 VSS.n5285 2.6005
R7693 VSS.n5284 VSS.n5283 2.6005
R7694 VSS.n5283 VSS.n5282 2.6005
R7695 VSS.n5280 VSS.n5279 2.6005
R7696 VSS.n5279 VSS.n5278 2.6005
R7697 VSS.n5277 VSS.n5276 2.6005
R7698 VSS.n5276 VSS.n5275 2.6005
R7699 VSS.n5274 VSS.n5273 2.6005
R7700 VSS.n5273 VSS.n5272 2.6005
R7701 VSS.n5271 VSS.n5270 2.6005
R7702 VSS.n5270 VSS.n5269 2.6005
R7703 VSS.n5268 VSS.n5267 2.6005
R7704 VSS.n5267 VSS.n5266 2.6005
R7705 VSS.n5247 VSS.n5246 2.6005
R7706 VSS.n5246 VSS.n5245 2.6005
R7707 VSS.n5250 VSS.n5249 2.6005
R7708 VSS.n5249 VSS.n5248 2.6005
R7709 VSS.n5253 VSS.n5252 2.6005
R7710 VSS.n5252 VSS.n5251 2.6005
R7711 VSS.n5255 VSS.n5254 2.6005
R7712 VSS.n5256 VSS.n5255 2.6005
R7713 VSS.n5244 VSS.n5243 2.6005
R7714 VSS.n5243 VSS.n5242 2.6005
R7715 VSS.n7905 VSS.n7904 2.6005
R7716 VSS.n7904 VSS.n7903 2.6005
R7717 VSS.n7902 VSS.n7901 2.6005
R7718 VSS.n7901 VSS.n7900 2.6005
R7719 VSS.n7899 VSS.n7898 2.6005
R7720 VSS.n7898 VSS.n7897 2.6005
R7721 VSS.n7896 VSS.n7895 2.6005
R7722 VSS.n7895 VSS.n7894 2.6005
R7723 VSS.n19 VSS.n18 2.6005
R7724 VSS.n18 VSS.n17 2.6005
R7725 VSS.n16 VSS.n15 2.6005
R7726 VSS.n15 VSS.n14 2.6005
R7727 VSS.n802 VSS.n801 2.6005
R7728 VSS.n801 VSS.n800 2.6005
R7729 VSS.n1141 VSS.n1140 2.6005
R7730 VSS.n1140 VSS.n1139 2.6005
R7731 VSS.n1144 VSS.n1143 2.6005
R7732 VSS.n1143 VSS.n1142 2.6005
R7733 VSS.n1147 VSS.n1146 2.6005
R7734 VSS.n1146 VSS.n1145 2.6005
R7735 VSS.n1150 VSS.n1149 2.6005
R7736 VSS.n1149 VSS.n1148 2.6005
R7737 VSS.n1153 VSS.n1152 2.6005
R7738 VSS.n1152 VSS.n1151 2.6005
R7739 VSS.n1156 VSS.n1155 2.6005
R7740 VSS.n1155 VSS.n1154 2.6005
R7741 VSS.n1159 VSS.n1158 2.6005
R7742 VSS.n1158 VSS.n1157 2.6005
R7743 VSS.n1162 VSS.n1161 2.6005
R7744 VSS.n1161 VSS.n1160 2.6005
R7745 VSS.n1165 VSS.n1164 2.6005
R7746 VSS.n1164 VSS.n1163 2.6005
R7747 VSS.n1168 VSS.n1167 2.6005
R7748 VSS.n1167 VSS.n1166 2.6005
R7749 VSS.n1171 VSS.n1170 2.6005
R7750 VSS.n1170 VSS.n1169 2.6005
R7751 VSS.n1174 VSS.n1173 2.6005
R7752 VSS.n1173 VSS.n1172 2.6005
R7753 VSS.n1177 VSS.n1176 2.6005
R7754 VSS.n1176 VSS.n1175 2.6005
R7755 VSS.n1180 VSS.n1179 2.6005
R7756 VSS.n1179 VSS.n1178 2.6005
R7757 VSS.n1183 VSS.n1182 2.6005
R7758 VSS.n1182 VSS.n1181 2.6005
R7759 VSS.n1186 VSS.n1185 2.6005
R7760 VSS.n1185 VSS.n1184 2.6005
R7761 VSS.n1189 VSS.n1188 2.6005
R7762 VSS.n1188 VSS.n1187 2.6005
R7763 VSS.n1192 VSS.n1191 2.6005
R7764 VSS.n1191 VSS.n1190 2.6005
R7765 VSS.n1195 VSS.n1194 2.6005
R7766 VSS.n1194 VSS.n1193 2.6005
R7767 VSS.n1198 VSS.n1197 2.6005
R7768 VSS.n1197 VSS.n1196 2.6005
R7769 VSS.n1201 VSS.n1200 2.6005
R7770 VSS.n1200 VSS.n1199 2.6005
R7771 VSS.n1204 VSS.n1203 2.6005
R7772 VSS.n1203 VSS.n1202 2.6005
R7773 VSS.n1207 VSS.n1206 2.6005
R7774 VSS.n1206 VSS.n1205 2.6005
R7775 VSS.n1210 VSS.n1209 2.6005
R7776 VSS.n1209 VSS.n1208 2.6005
R7777 VSS.n1213 VSS.n1212 2.6005
R7778 VSS.n1212 VSS.n1211 2.6005
R7779 VSS.n1216 VSS.n1215 2.6005
R7780 VSS.n1215 VSS.n1214 2.6005
R7781 VSS.n1219 VSS.n1218 2.6005
R7782 VSS.n1218 VSS.n1217 2.6005
R7783 VSS.n1222 VSS.n1221 2.6005
R7784 VSS.n1221 VSS.n1220 2.6005
R7785 VSS.n1225 VSS.n1224 2.6005
R7786 VSS.n1224 VSS.n1223 2.6005
R7787 VSS.n1228 VSS.n1227 2.6005
R7788 VSS.n1227 VSS.n1226 2.6005
R7789 VSS.n1231 VSS.n1230 2.6005
R7790 VSS.n1230 VSS.n1229 2.6005
R7791 VSS.n1234 VSS.n1233 2.6005
R7792 VSS.n1233 VSS.n1232 2.6005
R7793 VSS.n1237 VSS.n1236 2.6005
R7794 VSS.n1236 VSS.n1235 2.6005
R7795 VSS.n1240 VSS.n1239 2.6005
R7796 VSS.n1239 VSS.n1238 2.6005
R7797 VSS.n1243 VSS.n1242 2.6005
R7798 VSS.n1242 VSS.n1241 2.6005
R7799 VSS.n1246 VSS.n1245 2.6005
R7800 VSS.n1245 VSS.n1244 2.6005
R7801 VSS.n1249 VSS.n1248 2.6005
R7802 VSS.n1248 VSS.n1247 2.6005
R7803 VSS.n1253 VSS.n1252 2.6005
R7804 VSS.n790 VSS.n789 2.6005
R7805 VSS.n793 VSS.n792 2.6005
R7806 VSS.n795 VSS.n794 2.6005
R7807 VSS.n799 VSS.n798 2.6005
R7808 VSS.n7873 VSS.n7872 2.6005
R7809 VSS.n7877 VSS.n7876 2.6005
R7810 VSS.n5131 VSS.n5130 2.6005
R7811 VSS.n5130 VSS.n5129 2.6005
R7812 VSS.n5134 VSS.n5133 2.6005
R7813 VSS.n5133 VSS.n5132 2.6005
R7814 VSS.n5137 VSS.n5136 2.6005
R7815 VSS.n5136 VSS.n5135 2.6005
R7816 VSS.n5140 VSS.n5139 2.6005
R7817 VSS.n5139 VSS.n5138 2.6005
R7818 VSS.n5143 VSS.n5142 2.6005
R7819 VSS.n5142 VSS.n5141 2.6005
R7820 VSS.n5146 VSS.n5145 2.6005
R7821 VSS.n5145 VSS.n5144 2.6005
R7822 VSS.n5149 VSS.n5148 2.6005
R7823 VSS.n5148 VSS.n5147 2.6005
R7824 VSS.n5152 VSS.n5151 2.6005
R7825 VSS.n5151 VSS.n5150 2.6005
R7826 VSS.n5155 VSS.n5154 2.6005
R7827 VSS.n5154 VSS.n5153 2.6005
R7828 VSS.n5158 VSS.n5157 2.6005
R7829 VSS.n5157 VSS.n5156 2.6005
R7830 VSS.n7885 VSS.n7884 2.6005
R7831 VSS.n7886 VSS.n7885 2.6005
R7832 VSS.n7883 VSS.n7882 2.6005
R7833 VSS.n7882 VSS.n7881 2.6005
R7834 VSS.n7880 VSS.n7879 2.6005
R7835 VSS.n7879 VSS.n7878 2.6005
R7836 VSS.n5128 VSS.n5127 2.6005
R7837 VSS.n5127 VSS.n5126 2.6005
R7838 VSS.n4805 VSS.n4804 2.6005
R7839 VSS.n4804 VSS.n4803 2.6005
R7840 VSS.n4802 VSS.n4801 2.6005
R7841 VSS.n4801 VSS.n4800 2.6005
R7842 VSS.n4799 VSS.n4798 2.6005
R7843 VSS.n4798 VSS.n4797 2.6005
R7844 VSS.n4808 VSS.n4807 2.6005
R7845 VSS.n4807 VSS.n4806 2.6005
R7846 VSS.n4812 VSS.n4811 2.6005
R7847 VSS.n4811 VSS.n4810 2.6005
R7848 VSS.n4815 VSS.n4814 2.6005
R7849 VSS.n4814 VSS.n4813 2.6005
R7850 VSS.n4818 VSS.n4817 2.6005
R7851 VSS.n4817 VSS.n4816 2.6005
R7852 VSS.n4821 VSS.n4820 2.6005
R7853 VSS.n4820 VSS.n4819 2.6005
R7854 VSS.n4824 VSS.n4823 2.6005
R7855 VSS.n4823 VSS.n4822 2.6005
R7856 VSS.n4827 VSS.n4826 2.6005
R7857 VSS.n4826 VSS.n4825 2.6005
R7858 VSS.n4830 VSS.n4829 2.6005
R7859 VSS.n4829 VSS.n4828 2.6005
R7860 VSS.n4833 VSS.n4832 2.6005
R7861 VSS.n4832 VSS.n4831 2.6005
R7862 VSS.n4836 VSS.n4835 2.6005
R7863 VSS.n4835 VSS.n4834 2.6005
R7864 VSS.n4840 VSS.n4839 2.6005
R7865 VSS.n4839 VSS.n4838 2.6005
R7866 VSS.n4843 VSS.n4842 2.6005
R7867 VSS.n4842 VSS.n4841 2.6005
R7868 VSS.n4846 VSS.n4845 2.6005
R7869 VSS.n4845 VSS.n4844 2.6005
R7870 VSS.n4849 VSS.n4848 2.6005
R7871 VSS.n4848 VSS.n4847 2.6005
R7872 VSS.n4852 VSS.n4851 2.6005
R7873 VSS.n4851 VSS.n4850 2.6005
R7874 VSS.n4855 VSS.n4854 2.6005
R7875 VSS.n4854 VSS.n4853 2.6005
R7876 VSS.n4867 VSS.n4866 2.6005
R7877 VSS.n4866 VSS.n4865 2.6005
R7878 VSS.n4864 VSS.n4863 2.6005
R7879 VSS.n4863 VSS.n4862 2.6005
R7880 VSS.n4861 VSS.n4860 2.6005
R7881 VSS.n4860 VSS.n4859 2.6005
R7882 VSS.n4858 VSS.n4857 2.6005
R7883 VSS.n4857 VSS.n4856 2.6005
R7884 VSS.n5125 VSS.n5124 2.6005
R7885 VSS.n5124 VSS.n5123 2.6005
R7886 VSS.n860 VSS.n859 2.6005
R7887 VSS.n859 VSS.n858 2.6005
R7888 VSS.n924 VSS.n923 2.6005
R7889 VSS.n923 VSS.n922 2.6005
R7890 VSS.n810 VSS.n809 2.6005
R7891 VSS.n808 VSS.n807 2.6005
R7892 VSS.n805 VSS.n804 2.6005
R7893 VSS.n920 VSS.n919 2.6005
R7894 VSS.n919 VSS.n918 2.6005
R7895 VSS.n917 VSS.n916 2.6005
R7896 VSS.n916 VSS.n915 2.6005
R7897 VSS.n914 VSS.n913 2.6005
R7898 VSS.n913 VSS.n912 2.6005
R7899 VSS.n911 VSS.n910 2.6005
R7900 VSS.n910 VSS.n909 2.6005
R7901 VSS.n908 VSS.n907 2.6005
R7902 VSS.n907 VSS.n906 2.6005
R7903 VSS.n905 VSS.n904 2.6005
R7904 VSS.n904 VSS.n903 2.6005
R7905 VSS.n902 VSS.n901 2.6005
R7906 VSS.n901 VSS.n900 2.6005
R7907 VSS.n899 VSS.n898 2.6005
R7908 VSS.n898 VSS.n897 2.6005
R7909 VSS.n896 VSS.n895 2.6005
R7910 VSS.n895 VSS.n894 2.6005
R7911 VSS.n893 VSS.n892 2.6005
R7912 VSS.n892 VSS.n891 2.6005
R7913 VSS.n890 VSS.n889 2.6005
R7914 VSS.n889 VSS.n888 2.6005
R7915 VSS.n887 VSS.n886 2.6005
R7916 VSS.n886 VSS.n885 2.6005
R7917 VSS.n884 VSS.n883 2.6005
R7918 VSS.n883 VSS.n882 2.6005
R7919 VSS.n881 VSS.n880 2.6005
R7920 VSS.n880 VSS.n879 2.6005
R7921 VSS.n878 VSS.n877 2.6005
R7922 VSS.n877 VSS.n876 2.6005
R7923 VSS.n875 VSS.n874 2.6005
R7924 VSS.n874 VSS.n873 2.6005
R7925 VSS.n872 VSS.n871 2.6005
R7926 VSS.n871 VSS.n870 2.6005
R7927 VSS.n869 VSS.n868 2.6005
R7928 VSS.n868 VSS.n867 2.6005
R7929 VSS.n866 VSS.n865 2.6005
R7930 VSS.n865 VSS.n864 2.6005
R7931 VSS.n863 VSS.n862 2.6005
R7932 VSS.n862 VSS.n861 2.6005
R7933 VSS.n839 VSS.n838 2.6005
R7934 VSS.n838 VSS.n837 2.6005
R7935 VSS.n842 VSS.n841 2.6005
R7936 VSS.n841 VSS.n840 2.6005
R7937 VSS.n845 VSS.n844 2.6005
R7938 VSS.n844 VSS.n843 2.6005
R7939 VSS.n848 VSS.n847 2.6005
R7940 VSS.n847 VSS.n846 2.6005
R7941 VSS.n851 VSS.n850 2.6005
R7942 VSS.n850 VSS.n849 2.6005
R7943 VSS.n854 VSS.n853 2.6005
R7944 VSS.n853 VSS.n852 2.6005
R7945 VSS.n857 VSS.n856 2.6005
R7946 VSS.n856 VSS.n855 2.6005
R7947 VSS.n827 VSS.n826 2.6005
R7948 VSS.n829 VSS.n828 2.6005
R7949 VSS.n836 VSS.n835 2.6005
R7950 VSS.n821 VSS.n820 2.6005
R7951 VSS.n824 VSS.n823 2.6005
R7952 VSS.n819 VSS.n818 2.6005
R7953 VSS.n986 VSS.n963 2.6005
R7954 VSS.n963 VSS.n962 2.6005
R7955 VSS.n984 VSS.n983 2.6005
R7956 VSS.n983 VSS.n982 2.6005
R7957 VSS.n981 VSS.n980 2.6005
R7958 VSS.n980 VSS.n979 2.6005
R7959 VSS.n978 VSS.n977 2.6005
R7960 VSS.n977 VSS.n976 2.6005
R7961 VSS.n975 VSS.n974 2.6005
R7962 VSS.n974 VSS.n973 2.6005
R7963 VSS VSS.n971 2.6005
R7964 VSS.n971 VSS.n970 2.6005
R7965 VSS.n969 VSS.n967 2.6005
R7966 VSS.n969 VSS.n968 2.6005
R7967 VSS.n960 VSS.n959 2.6005
R7968 VSS.n959 VSS.n958 2.6005
R7969 VSS.n957 VSS.n956 2.6005
R7970 VSS.n956 VSS.n955 2.6005
R7971 VSS.n954 VSS.n953 2.6005
R7972 VSS.n953 VSS.n952 2.6005
R7973 VSS.n950 VSS.n949 2.6005
R7974 VSS.n949 VSS.n948 2.6005
R7975 VSS.n817 VSS.n816 2.6005
R7976 VSS.n815 VSS.n814 2.6005
R7977 VSS.n1008 VSS.n1007 2.6005
R7978 VSS.n1007 VSS.n1006 2.6005
R7979 VSS.n1011 VSS.n1010 2.6005
R7980 VSS.n1010 VSS.n1009 2.6005
R7981 VSS.n1014 VSS.n1013 2.6005
R7982 VSS.n1013 VSS.n1012 2.6005
R7983 VSS.n1017 VSS.n1016 2.6005
R7984 VSS.n1016 VSS.n1015 2.6005
R7985 VSS.n1021 VSS.n1020 2.6005
R7986 VSS.n1020 VSS.n1019 2.6005
R7987 VSS.n1024 VSS.n1023 2.6005
R7988 VSS.n1023 VSS.n1022 2.6005
R7989 VSS.n1027 VSS.n1026 2.6005
R7990 VSS.n1026 VSS.n1025 2.6005
R7991 VSS.n1031 VSS.n1030 2.6005
R7992 VSS.n1030 VSS.n1029 2.6005
R7993 VSS.n1034 VSS.n1033 2.6005
R7994 VSS.n1033 VSS.n1032 2.6005
R7995 VSS.n1037 VSS.n1036 2.6005
R7996 VSS.n1036 VSS.n1035 2.6005
R7997 VSS.n1040 VSS.n1039 2.6005
R7998 VSS.n1039 VSS.n1038 2.6005
R7999 VSS.n1043 VSS.n1042 2.6005
R8000 VSS.n1042 VSS.n1041 2.6005
R8001 VSS.n1047 VSS.n1046 2.6005
R8002 VSS.n1046 VSS.n1045 2.6005
R8003 VSS.n1050 VSS.n1049 2.6005
R8004 VSS.n1049 VSS.n1048 2.6005
R8005 VSS.n1053 VSS.n1052 2.6005
R8006 VSS.n1052 VSS.n1051 2.6005
R8007 VSS.n1056 VSS.n1055 2.6005
R8008 VSS.n1055 VSS.n1054 2.6005
R8009 VSS.n1059 VSS.n1058 2.6005
R8010 VSS.n1058 VSS.n1057 2.6005
R8011 VSS.n1062 VSS.n1061 2.6005
R8012 VSS.n1061 VSS.n1060 2.6005
R8013 VSS.n1065 VSS.n1064 2.6005
R8014 VSS.n1064 VSS.n1063 2.6005
R8015 VSS.n1069 VSS.n1068 2.6005
R8016 VSS.n1068 VSS.n1067 2.6005
R8017 VSS.n1072 VSS.n1071 2.6005
R8018 VSS.n1071 VSS.n1070 2.6005
R8019 VSS.n1075 VSS.n1074 2.6005
R8020 VSS.n1074 VSS.n1073 2.6005
R8021 VSS.n1079 VSS.n1078 2.6005
R8022 VSS.n1078 VSS.n1077 2.6005
R8023 VSS.n1082 VSS.n1081 2.6005
R8024 VSS.n1081 VSS.n1080 2.6005
R8025 VSS.n1087 VSS.n1086 2.6005
R8026 VSS.n1086 VSS.n1085 2.6005
R8027 VSS.n1126 VSS.n1125 2.6005
R8028 VSS.n1124 VSS.n1123 2.6005
R8029 VSS.n1123 VSS.n1122 2.6005
R8030 VSS.n1121 VSS.n1120 2.6005
R8031 VSS.n1120 VSS.n1119 2.6005
R8032 VSS.n1118 VSS.n1117 2.6005
R8033 VSS.n1117 VSS.n1116 2.6005
R8034 VSS.n1115 VSS.n1114 2.6005
R8035 VSS.n1114 VSS.n1113 2.6005
R8036 VSS.n1112 VSS.n1111 2.6005
R8037 VSS.n1111 VSS.n1110 2.6005
R8038 VSS.n1109 VSS.n1108 2.6005
R8039 VSS.n1108 VSS.n1107 2.6005
R8040 VSS.n1106 VSS.n1105 2.6005
R8041 VSS.n1101 VSS.n1100 2.6005
R8042 VSS.n1099 VSS.n1098 2.6005
R8043 VSS.n1096 VSS.n1095 2.6005
R8044 VSS.n1092 VSS.n1091 2.6005
R8045 VSS.n1090 VSS.n1089 2.6005
R8046 VSS.n1089 VSS.n1088 2.6005
R8047 VSS.n1129 VSS.n1128 2.6005
R8048 VSS.n7 VSS.n6 2.6005
R8049 VSS.n10 VSS.n9 2.6005
R8050 VSS.n4 VSS.n3 2.6005
R8051 VSS.n4444 VSS.n4443 2.59998
R8052 VSS.n1788 VSS.n1787 2.53192
R8053 VSS.n1424 VSS.n1423 2.48961
R8054 VSS.n1427 VSS.n1426 2.48961
R8055 VSS.n1430 VSS.n1429 2.48961
R8056 VSS.n1433 VSS.n1432 2.48961
R8057 VSS.n1436 VSS.n1435 2.48961
R8058 VSS.n1439 VSS.n1438 2.48961
R8059 VSS.n1442 VSS.n1441 2.48961
R8060 VSS.n1445 VSS.n1444 2.48961
R8061 VSS.n1448 VSS.n1447 2.48961
R8062 VSS.n285 VSS.n284 2.41686
R8063 VSS.n1867 VSS.n1775 2.3405
R8064 VSS.n1868 VSS.n1765 2.33208
R8065 VSS.n1788 VSS.n1783 2.33079
R8066 VSS.n2234 VSS.n2233 2.28632
R8067 VSS.n7482 VSS.n7481 2.28399
R8068 VSS.n385 VSS.n384 2.28399
R8069 VSS.n388 VSS.n387 2.28399
R8070 VSS.n504 VSS.n503 2.28399
R8071 VSS.n507 VSS.n506 2.28399
R8072 VSS.n4092 VSS.n4091 2.27928
R8073 VSS.n2873 VSS.n2363 2.2791
R8074 VSS.n2730 VSS.n2571 2.27836
R8075 VSS.n2353 VSS.n2352 2.27834
R8076 VSS.n7150 VSS.n7149 2.27775
R8077 VSS.n3024 VSS.n2140 2.27413
R8078 VSS.n2942 VSS.n2247 2.27187
R8079 VSS.n2808 VSS.n2472 2.26934
R8080 VSS.n3577 VSS.n3576 2.26031
R8081 VSS.n2466 VSS.n2465 2.25712
R8082 VSS.n5905 VSS.n5904 2.25635
R8083 VSS.n2723 VSS.n2576 2.25613
R8084 VSS.n681 VSS.n680 2.25576
R8085 VSS.n3875 VSS.t617 2.25428
R8086 VSS.n3876 VSS.t614 2.25428
R8087 VSS.n3877 VSS.t603 2.25428
R8088 VSS.n3878 VSS.t678 2.25428
R8089 VSS.n3879 VSS.t670 2.25428
R8090 VSS.n3880 VSS.t691 2.25428
R8091 VSS.n3881 VSS.t621 2.25428
R8092 VSS.n3882 VSS.t620 2.25428
R8093 VSS.n3883 VSS.t693 2.25428
R8094 VSS.n3884 VSS.t685 2.25428
R8095 VSS.n3885 VSS.t588 2.25428
R8096 VSS.n3886 VSS.t631 2.25428
R8097 VSS.n1925 VSS.t664 2.25428
R8098 VSS.n1926 VSS.t642 2.25428
R8099 VSS.n1927 VSS.t654 2.25428
R8100 VSS.n1928 VSS.t698 2.25428
R8101 VSS.n1929 VSS.t701 2.25428
R8102 VSS.n1930 VSS.t651 2.25428
R8103 VSS.n1931 VSS.t629 2.25428
R8104 VSS.n1932 VSS.t639 2.25428
R8105 VSS.n1933 VSS.t683 2.25428
R8106 VSS.n1934 VSS.t335 2.25428
R8107 VSS.n1935 VSS.t336 2.25428
R8108 VSS.n2622 VSS.t626 2.25428
R8109 VSS.n2623 VSS.t605 2.25428
R8110 VSS.n2624 VSS.t615 2.25428
R8111 VSS.n2625 VSS.t655 2.25428
R8112 VSS.n2626 VSS.t658 2.25428
R8113 VSS.n2627 VSS.t611 2.25428
R8114 VSS.n2628 VSS.t591 2.25428
R8115 VSS.n2629 VSS.t719 2.25428
R8116 VSS.n2630 VSS.t640 2.25428
R8117 VSS.n2631 VSS.t647 2.25428
R8118 VSS.n2632 VSS.t649 2.25428
R8119 VSS.n2531 VSS.t673 2.25428
R8120 VSS.n2532 VSS.t652 2.25428
R8121 VSS.n2533 VSS.t660 2.25428
R8122 VSS.n2534 VSS.t587 2.25428
R8123 VSS.n2535 VSS.t589 2.25428
R8124 VSS.n2536 VSS.t659 2.25428
R8125 VSS.n2537 VSS.t638 2.25428
R8126 VSS.n2538 VSS.t644 2.25428
R8127 VSS.n2539 VSS.t776 2.25428
R8128 VSS.n2540 VSS.t777 2.25428
R8129 VSS.n2541 VSS.t778 2.25428
R8130 VSS.n2421 VSS.t704 2.25428
R8131 VSS.n2422 VSS.t680 2.25428
R8132 VSS.n2423 VSS.t689 2.25428
R8133 VSS.n2424 VSS.t618 2.25428
R8134 VSS.n2425 VSS.t619 2.25428
R8135 VSS.n2426 VSS.t687 2.25428
R8136 VSS.n2427 VSS.t665 2.25428
R8137 VSS.n2428 VSS.t676 2.25428
R8138 VSS.n2429 VSS.t600 2.25428
R8139 VSS.n2430 VSS.t609 2.25428
R8140 VSS.n2431 VSS.t612 2.25428
R8141 VSS.n2299 VSS.t643 2.25428
R8142 VSS.n2300 VSS.t627 2.25428
R8143 VSS.n2301 VSS.t633 2.25428
R8144 VSS.n2302 VSS.t677 2.25428
R8145 VSS.n2303 VSS.t679 2.25428
R8146 VSS.n2304 VSS.t630 2.25428
R8147 VSS.n2305 VSS.t616 2.25428
R8148 VSS.n2306 VSS.t622 2.25428
R8149 VSS.n2307 VSS.t663 2.25428
R8150 VSS.n2308 VSS.t672 2.25428
R8151 VSS.n2309 VSS.t674 2.25428
R8152 VSS.n2187 VSS.t696 2.25428
R8153 VSS.n2188 VSS.t675 2.25428
R8154 VSS.n2189 VSS.t684 2.25428
R8155 VSS.n2190 VSS.t608 2.25428
R8156 VSS.n2191 VSS.t610 2.25428
R8157 VSS.n2192 VSS.t681 2.25428
R8158 VSS.n2193 VSS.t661 2.25428
R8159 VSS.n2194 VSS.t668 2.25428
R8160 VSS.n2195 VSS.t595 2.25428
R8161 VSS.n2196 VSS.t602 2.25428
R8162 VSS.n2197 VSS.t606 2.25428
R8163 VSS.n2126 VSS.t607 2.25428
R8164 VSS.n2127 VSS.t586 2.25428
R8165 VSS.n2128 VSS.t594 2.25428
R8166 VSS.n2129 VSS.t635 2.25428
R8167 VSS.n2130 VSS.t637 2.25428
R8168 VSS.n2131 VSS.t593 2.25428
R8169 VSS.n2132 VSS.t690 2.25428
R8170 VSS.n2133 VSS.t699 2.25428
R8171 VSS.n2134 VSS.t624 2.25428
R8172 VSS.n2135 VSS.t720 2.25428
R8173 VSS.n2136 VSS.t721 2.25428
R8174 VSS.n1971 VSS.t604 2.25428
R8175 VSS.n1972 VSS.t705 2.25428
R8176 VSS.n1973 VSS.t592 2.25428
R8177 VSS.n1974 VSS.t634 2.25428
R8178 VSS.n1975 VSS.t636 2.25428
R8179 VSS.n1976 VSS.t590 2.25428
R8180 VSS.n1977 VSS.t688 2.25428
R8181 VSS.n1978 VSS.t697 2.25428
R8182 VSS.n1979 VSS.t623 2.25428
R8183 VSS.n1980 VSS.t717 2.25428
R8184 VSS.n1981 VSS.t718 2.25428
R8185 VSS.n1947 VSS.t682 2.25428
R8186 VSS.n1948 VSS.t662 2.25428
R8187 VSS.n1949 VSS.t669 2.25428
R8188 VSS.n1950 VSS.t597 2.25428
R8189 VSS.n1951 VSS.t599 2.25428
R8190 VSS.n1952 VSS.t667 2.25428
R8191 VSS.n1953 VSS.t646 2.25428
R8192 VSS.n1954 VSS.t657 2.25428
R8193 VSS.n1955 VSS.t702 2.25428
R8194 VSS.n1956 VSS.t541 2.25428
R8195 VSS.n1957 VSS.t542 2.25428
R8196 VSS.n1936 VSS.t666 2.25428
R8197 VSS.n1937 VSS.t645 2.25428
R8198 VSS.n1938 VSS.t656 2.25428
R8199 VSS.n1939 VSS.t700 2.25428
R8200 VSS.n1940 VSS.t703 2.25428
R8201 VSS.n1941 VSS.t653 2.25428
R8202 VSS.n1942 VSS.t632 2.25428
R8203 VSS.n1943 VSS.t641 2.25428
R8204 VSS.n1944 VSS.t686 2.25428
R8205 VSS.n1945 VSS.t692 2.25428
R8206 VSS.n1946 VSS.t695 2.25428
R8207 VSS.n4029 VSS.t281 2.25416
R8208 VSS.n3887 VSS.t283 2.25416
R8209 VSS.n3888 VSS.t285 2.25416
R8210 VSS.n1872 VSS.t282 2.25416
R8211 VSS.n4126 VSS.n4125 2.2531
R8212 VSS.n4091 VSS.n4087 2.2531
R8213 VSS.n4101 VSS.n4100 2.2531
R8214 VSS.n1486 VSS.n1485 2.25285
R8215 VSS.n7622 VSS.n7621 2.25285
R8216 VSS.n6620 VSS.n6619 2.25285
R8217 VSS.n2664 VSS.n2656 2.25113
R8218 VSS.n4110 VSS.n4109 2.25077
R8219 VSS.n4119 VSS.n4118 2.25077
R8220 VSS.n1866 VSS.n1865 2.2505
R8221 VSS.n1801 VSS.n1800 2.2505
R8222 VSS.n1793 VSS.n1792 2.2505
R8223 VSS.n1791 VSS.n1790 2.2505
R8224 VSS.n1799 VSS.n1798 2.2505
R8225 VSS.n3566 VSS.n3538 2.2505
R8226 VSS.n3568 VSS.n3567 2.2505
R8227 VSS.n3557 VSS.n3541 2.2505
R8228 VSS.n3555 VSS.n3554 2.2505
R8229 VSS.n3565 VSS.n3539 2.2505
R8230 VSS.n3547 VSS.n3543 2.2505
R8231 VSS.n3550 VSS.n3542 2.2505
R8232 VSS.n3559 VSS.n3540 2.2505
R8233 VSS.n3237 VSS.n3236 2.2505
R8234 VSS.n3385 VSS.n3374 2.2505
R8235 VSS.n3229 VSS.n3228 2.2505
R8236 VSS.n3390 VSS.n3373 2.2505
R8237 VSS.n3382 VSS.n3376 2.2505
R8238 VSS.n3394 VSS.n3371 2.2505
R8239 VSS.n3072 VSS.n3071 2.2505
R8240 VSS.n3097 VSS.n3096 2.2505
R8241 VSS.n3087 VSS.n3086 2.2505
R8242 VSS.n3076 VSS.n3075 2.2505
R8243 VSS.n3095 VSS.n3094 2.2505
R8244 VSS.n2093 VSS.n2092 2.2505
R8245 VSS.n2114 VSS.n2083 2.2505
R8246 VSS.n2103 VSS.n2085 2.2505
R8247 VSS.n2095 VSS.n2094 2.2505
R8248 VSS.n2104 VSS.n2084 2.2505
R8249 VSS.n2100 VSS.n2086 2.2505
R8250 VSS.n2231 VSS.n2213 2.2505
R8251 VSS.n2155 VSS.n2140 2.2505
R8252 VSS.n2233 VSS.n2216 2.2505
R8253 VSS.n2229 VSS.n2182 2.2505
R8254 VSS.n2226 VSS.n2158 2.2505
R8255 VSS.n2984 VSS.n2983 2.2505
R8256 VSS.n2230 VSS.n2183 2.2505
R8257 VSS.n2227 VSS.n2160 2.2505
R8258 VSS.n2232 VSS.n2214 2.2505
R8259 VSS.n2228 VSS.n2174 2.2505
R8260 VSS.n2288 VSS.n2283 2.2505
R8261 VSS.n2926 VSS.n2258 2.2505
R8262 VSS.n2904 VSS.n2294 2.2505
R8263 VSS.n2292 VSS.n2291 2.2505
R8264 VSS.n2906 VSS.n2905 2.2505
R8265 VSS.n2257 VSS.n2247 2.2505
R8266 VSS.n2293 VSS.n2280 2.2505
R8267 VSS.n2352 VSS.n2351 2.2505
R8268 VSS.n2343 VSS.n2342 2.2505
R8269 VSS.n2344 VSS.n2333 2.2505
R8270 VSS.n2413 VSS.n2384 2.2505
R8271 VSS.n2404 VSS.n2363 2.2505
R8272 VSS.n2457 VSS.n2451 2.2505
R8273 VSS.n2410 VSS.n2403 2.2505
R8274 VSS.n2837 VSS.n2414 2.2505
R8275 VSS.n2412 VSS.n2411 2.2505
R8276 VSS.n2836 VSS.n2415 2.2505
R8277 VSS.n2465 VSS.n2464 2.2505
R8278 VSS.n2792 VSS.n2485 2.2505
R8279 VSS.n2483 VSS.n2472 2.2505
R8280 VSS.n2568 VSS.n2567 2.2505
R8281 VSS.n2767 VSS.n2523 2.2505
R8282 VSS.n2522 VSS.n2521 2.2505
R8283 VSS.n2570 VSS.n2569 2.2505
R8284 VSS.n2571 VSS.n2557 2.2505
R8285 VSS.n2517 VSS.n2498 2.2505
R8286 VSS.n2519 VSS.n2518 2.2505
R8287 VSS.n2772 VSS.n2771 2.2505
R8288 VSS.n2651 VSS.n2650 2.2505
R8289 VSS.n2693 VSS.n2602 2.2505
R8290 VSS.n2648 VSS.n2603 2.2505
R8291 VSS.n2671 VSS.n2652 2.2505
R8292 VSS.n2709 VSS.n2708 2.2505
R8293 VSS.n2706 VSS.n2705 2.2505
R8294 VSS.n2589 VSS.n2576 2.2505
R8295 VSS.n2704 VSS.n2703 2.2505
R8296 VSS.n2711 VSS.n2710 2.2505
R8297 VSS.n2712 VSS.n2584 2.2505
R8298 VSS.n2702 VSS.n2701 2.2505
R8299 VSS.n4111 VSS.n4110 2.2505
R8300 VSS.n4127 VSS.n4126 2.2505
R8301 VSS.n4120 VSS.n4119 2.2505
R8302 VSS.n4102 VSS.n4101 2.2505
R8303 VSS.n7127 VSS.n7126 2.2505
R8304 VSS.n151 VSS.n150 2.2505
R8305 VSS.n223 VSS.n215 2.2505
R8306 VSS.n1539 VSS.n1538 2.2505
R8307 VSS.n1586 VSS.n1585 2.2505
R8308 VSS.n93 VSS.n92 2.2505
R8309 VSS.n4563 VSS.n4562 2.2505
R8310 VSS.n4551 VSS.n4550 2.2505
R8311 VSS.n4384 VSS.n4379 2.2505
R8312 VSS.n1597 VSS.n1596 2.2505
R8313 VSS.n3995 VSS.n1879 2.24994
R8314 VSS.n4098 VSS.n4097 2.24924
R8315 VSS.n6400 VSS.n6399 2.24725
R8316 VSS.n932 VSS.n931 2.24725
R8317 VSS.n778 VSS.n777 2.24654
R8318 VSS.n6398 VSS.n6397 2.24654
R8319 VSS.n7164 VSS.n7124 2.24654
R8320 VSS.n7620 VSS.n5306 2.24654
R8321 VSS.n6624 VSS.n6623 2.24654
R8322 VSS.n718 VSS.n717 2.24654
R8323 VSS.n930 VSS.n929 2.24654
R8324 VSS.n4884 VSS.n4872 2.24592
R8325 VSS.n3994 VSS.n3993 2.24495
R8326 VSS.n4881 VSS.n4875 2.24465
R8327 VSS.n4126 VSS.n4123 2.24449
R8328 VSS.n4091 VSS.n4090 2.24449
R8329 VSS.n283 VSS.n282 2.22001
R8330 VSS.n7140 VSS.t145 2.16717
R8331 VSS.n7140 VSS.n7139 2.16717
R8332 VSS.n7149 VSS 2.0871
R8333 VSS.n192 VSS.n190 2.04928
R8334 VSS.n989 VSS.t898 2.02838
R8335 VSS.n716 VSS.t21 2.02838
R8336 VSS.n6622 VSS.t821 2.02838
R8337 VSS.n6488 VSS.t935 2.02838
R8338 VSS.n5305 VSS.t132 2.02838
R8339 VSS.n1477 VSS.t910 2.02837
R8340 VSS.n80 VSS.t149 2.02837
R8341 VSS.n7225 VSS.t94 2.02837
R8342 VSS.t442 VSS.t499 2.02605
R8343 VSS.t424 VSS.t442 2.02605
R8344 VSS.n5842 VSS.t732 2.02605
R8345 VSS.n4598 VSS.n4597 2.0097
R8346 VSS.n6746 VSS.n6745 2.0097
R8347 VSS.n6396 VSS.n6395 2.0097
R8348 VSS.n6946 VSS.n6945 2.0097
R8349 VSS.n928 VSS.n927 2.0097
R8350 VSS.n776 VSS.n775 2.00969
R8351 VSS.n177 VSS.n176 2.00969
R8352 VSS.n7123 VSS.n7122 2.00969
R8353 VSS.n190 VSS.n175 1.96391
R8354 VSS.n7146 VSS.t830 1.9505
R8355 VSS.n7146 VSS.n7145 1.9505
R8356 VSS.n7801 VSS 1.9362
R8357 VSS.t993 VSS.n6986 1.92522
R8358 VSS.t989 VSS.n6987 1.92522
R8359 VSS.t992 VSS.n6985 1.92328
R8360 VSS.t528 VSS.t525 1.92017
R8361 VSS.t558 VSS.t556 1.92017
R8362 VSS.t531 VSS.t940 1.92017
R8363 VSS.n1398 VSS.n1397 1.87586
R8364 VSS.n4610 VSS.n4609 1.87586
R8365 VSS.n4872 VSS.n4870 1.85787
R8366 VSS.n4875 VSS.n4874 1.85787
R8367 VSS.n5430 VSS.n5429 1.85765
R8368 VSS.n5410 VSS.n5409 1.85765
R8369 VSS.n44 VSS.n43 1.83785
R8370 VSS.n4766 VSS.n4765 1.83785
R8371 VSS.n5917 VSS.n5916 1.83785
R8372 VSS.n5885 VSS.n5884 1.83785
R8373 VSS.n4772 VSS.n4771 1.83724
R8374 VSS.n5943 VSS.n5942 1.83724
R8375 VSS.n5947 VSS.n5946 1.83724
R8376 VSS.n5400 VSS.n5399 1.83724
R8377 VSS.n5120 VSS.n5119 1.83724
R8378 VSS.n7876 VSS.n7875 1.83724
R8379 VSS.n4786 VSS.n4785 1.83716
R8380 VSS.n691 VSS.n690 1.82536
R8381 VSS.n776 VSS.t154 1.82525
R8382 VSS.n177 VSS.t81 1.82525
R8383 VSS.n7123 VSS.t947 1.82525
R8384 VSS.n4598 VSS.t257 1.82525
R8385 VSS.n6746 VSS.t890 1.82525
R8386 VSS.n6396 VSS.t902 1.82525
R8387 VSS.n6946 VSS.t120 1.82525
R8388 VSS.n928 VSS.t123 1.82525
R8389 VSS.n1591 VSS.n1590 1.82479
R8390 VSS.n4219 VSS.n4217 1.81655
R8391 VSS.n1738 VSS.n1736 1.81655
R8392 VSS.n1477 VSS.n1476 1.80405
R8393 VSS.n80 VSS.n79 1.80405
R8394 VSS.n7225 VSS.n7224 1.80405
R8395 VSS.n989 VSS.n988 1.80404
R8396 VSS.n716 VSS.n715 1.80404
R8397 VSS.n6622 VSS.n6621 1.80404
R8398 VSS.n6488 VSS.n6487 1.80404
R8399 VSS.n5305 VSS.n5304 1.80404
R8400 VSS.n710 VSS.n709 1.8001
R8401 VSS.n317 VSS.n314 1.8001
R8402 VSS.n4696 VSS.n4689 1.8001
R8403 VSS.n4425 VSS.n4424 1.8001
R8404 VSS.n4346 VSS.n4343 1.8001
R8405 VSS.n4136 VSS.n4133 1.8001
R8406 VSS.n304 VSS.n303 1.79951
R8407 VSS.n4136 VSS.n4135 1.79951
R8408 VSS.n4144 VSS.n4143 1.79951
R8409 VSS.n317 VSS.n316 1.79951
R8410 VSS.n4662 VSS.n4659 1.79951
R8411 VSS.n4696 VSS.n4695 1.79951
R8412 VSS.n4346 VSS.n4345 1.79951
R8413 VSS.n4499 VSS.n4495 1.79951
R8414 VSS.n4622 VSS.n4621 1.79951
R8415 VSS.n4628 VSS.n4627 1.79942
R8416 VSS.n4670 VSS.n4669 1.79942
R8417 VSS.n283 VSS.n280 1.79318
R8418 VSS.n4414 VSS.n4411 1.7505
R8419 VSS.n37 VSS.n36 1.7445
R8420 VSS.n4423 VSS.n4422 1.7096
R8421 VSS.n1131 VSS.n1130 1.7025
R8422 VSS.n6576 VSS.n6575 1.68478
R8423 VSS.n7732 VSS.n7729 1.68478
R8424 VSS.n6382 VSS.n6381 1.68478
R8425 VSS.n6373 VSS.n6372 1.68478
R8426 VSS.n6342 VSS.n6341 1.68478
R8427 VSS.n1095 VSS.n1094 1.68478
R8428 VSS.n1409 VSS.n1408 1.68421
R8429 VSS.n1415 VSS.n1414 1.68421
R8430 VSS.n7277 VSS.n7276 1.68421
R8431 VSS.n7420 VSS.n7419 1.68421
R8432 VSS.n6373 VSS.n6370 1.68421
R8433 VSS.n6382 VSS.n6379 1.68421
R8434 VSS.n6992 VSS.n6991 1.68421
R8435 VSS.n6961 VSS.n6960 1.68421
R8436 VSS.n7530 VSS.n7529 1.68421
R8437 VSS.n4505 VSS.n4503 1.68421
R8438 VSS.n1367 VSS.n1366 1.68421
R8439 VSS.n6859 VSS.n6858 1.68421
R8440 VSS.n823 VSS.n822 1.68421
R8441 VSS.n1131 VSS.n1129 1.68421
R8442 VSS.n4838 VSS.n4837 1.68415
R8443 VSS.n1351 VSS.n1350 1.68411
R8444 VSS.n1356 VSS.n1355 1.68411
R8445 VSS.n1361 VSS.n1360 1.68411
R8446 VSS.n782 VSS.n781 1.68411
R8447 VSS.n6865 VSS.n6864 1.68411
R8448 VSS.n7645 VSS.n7644 1.68411
R8449 VSS.n7650 VSS.n7649 1.68411
R8450 VSS.n7655 VSS.n7654 1.68411
R8451 VSS.n7660 VSS.n7659 1.68411
R8452 VSS.n7666 VSS.n7665 1.68411
R8453 VSS.n734 VSS.n733 1.65879
R8454 VSS.n740 VSS.n739 1.65879
R8455 VSS.n750 VSS.n749 1.65879
R8456 VSS.n741 VSS.n740 1.65822
R8457 VSS.n747 VSS.n746 1.65822
R8458 VSS.n4531 VSS.n4530 1.65811
R8459 VSS.n644 VSS.n640 1.65328
R8460 VSS.n3887 VSS.n3886 1.65243
R8461 VSS.n158 VSS.n157 1.62245
R8462 VSS.n5331 VSS.n5330 1.6134
R8463 VSS.n5084 VSS.n5083 1.60209
R8464 VSS.n5103 VSS.n5102 1.60209
R8465 VSS.n5211 VSS.n5210 1.60209
R8466 VSS.n7853 VSS.n7852 1.60209
R8467 VSS.n5659 VSS.n5658 1.60209
R8468 VSS.n5786 VSS.n5785 1.60209
R8469 VSS.n7870 VSS.n7869 1.60209
R8470 VSS.n5113 VSS.n5112 1.60209
R8471 VSS.n6113 VSS.n6112 1.60199
R8472 VSS.n5723 VSS.n5722 1.60199
R8473 VSS.n5892 VSS.n5891 1.60199
R8474 VSS.n6230 VSS.n6229 1.60199
R8475 VSS.n7856 VSS.n7855 1.60199
R8476 VSS.n5214 VSS.n5213 1.60199
R8477 VSS.n5201 VSS.n5200 1.60199
R8478 VSS.n5106 VSS.n5105 1.60199
R8479 VSS.n5087 VSS.n5086 1.60199
R8480 VSS.n5076 VSS.n5075 1.60199
R8481 VSS.n4795 VSS.n4794 1.60199
R8482 VSS.n4790 VSS.n4789 1.60199
R8483 VSS.n324 VSS.n320 1.59295
R8484 VSS.n324 VSS.n323 1.5924
R8485 VSS.n4706 VSS.n4705 1.5924
R8486 VSS.n4727 VSS.n4726 1.59228
R8487 VSS.n4711 VSS.n4710 1.59228
R8488 VSS.n4741 VSS.n4740 1.59228
R8489 VSS.n792 VSS.n791 1.59228
R8490 VSS.n798 VSS.n797 1.59228
R8491 VSS.n6326 VSS.n6325 1.58814
R8492 VSS.n6321 VSS.n6320 1.58814
R8493 VSS.n6316 VSS.n6315 1.58814
R8494 VSS.n6311 VSS.n6310 1.58814
R8495 VSS.n6306 VSS.n6305 1.58814
R8496 VSS.n6298 VSS.n6297 1.58814
R8497 VSS.n6293 VSS.n6292 1.58814
R8498 VSS.n6288 VSS.n6287 1.58814
R8499 VSS.n517 VSS.n516 1.58814
R8500 VSS.n7737 VSS.n7734 1.58814
R8501 VSS.n5387 VSS.n5382 1.58814
R8502 VSS.n6278 VSS.n6277 1.58814
R8503 VSS.n7433 VSS.n7432 1.58759
R8504 VSS.n424 VSS.n423 1.58759
R8505 VSS.n5359 VSS.n5357 1.58759
R8506 VSS.n330 VSS.n329 1.58747
R8507 VSS.n6269 VSS.n6268 1.58747
R8508 VSS.n6241 VSS.n6240 1.58747
R8509 VSS.n6246 VSS.n6245 1.58747
R8510 VSS.n6262 VSS.n6261 1.58747
R8511 VSS.n6252 VSS.n6251 1.58747
R8512 VSS.n6257 VSS.n6256 1.58747
R8513 VSS.n222 VSS.n219 1.56241
R8514 VSS.n1550 VSS.n1548 1.55606
R8515 VSS.n7711 VSS.n7710 1.50443
R8516 VSS.n1868 VSS.n1867 1.50266
R8517 VSS.n4081 VSS.n4080 1.50144
R8518 VSS.n1773 VSS.n1772 1.5005
R8519 VSS.n4051 VSS.n4050 1.5005
R8520 VSS.n1878 VSS.n1877 1.5005
R8521 VSS.n3988 VSS.n3987 1.5005
R8522 VSS.n3902 VSS.n3901 1.5005
R8523 VSS.n3955 VSS.n3954 1.5005
R8524 VSS.n3919 VSS.n3918 1.5005
R8525 VSS.n3930 VSS.n3929 1.5005
R8526 VSS.n3975 VSS.n3974 1.5005
R8527 VSS.n1763 VSS.n1762 1.5005
R8528 VSS.n196 VSS.n194 1.5005
R8529 VSS.n4085 VSS.n4084 1.49611
R8530 VSS.n1604 VSS.n1600 1.45883
R8531 VSS.n7843 VSS.n7842 1.45883
R8532 VSS.n4892 VSS.n4891 1.4383
R8533 VSS.n6174 VSS.n6171 1.43813
R8534 VSS.n6472 VSS.n6471 1.43195
R8535 VSS.n6463 VSS.n6462 1.43195
R8536 VSS.n7325 VSS.n7324 1.43195
R8537 VSS.n7271 VSS.n7270 1.43195
R8538 VSS.n6337 VSS.n6336 1.43195
R8539 VSS.n6707 VSS.n6706 1.43195
R8540 VSS.n6725 VSS.n6724 1.43195
R8541 VSS.n1255 VSS.n1254 1.43195
R8542 VSS.n806 VSS.n805 1.43195
R8543 VSS.n1098 VSS.n1097 1.43195
R8544 VSS.n826 VSS.n825 1.43182
R8545 VSS.n835 VSS.n834 1.43182
R8546 VSS.n1105 VSS.n1104 1.43182
R8547 VSS.n811 VSS.n810 1.43182
R8548 VSS.n1452 VSS.n1451 1.43182
R8549 VSS.n1341 VSS.n1340 1.43182
R8550 VSS.n1346 VSS.n1345 1.43182
R8551 VSS.n1386 VSS.n1385 1.43182
R8552 VSS.n1380 VSS.n1379 1.43182
R8553 VSS.n6466 VSS.n6465 1.43182
R8554 VSS.n7309 VSS.n7308 1.43182
R8555 VSS.n7331 VSS.n7330 1.43182
R8556 VSS.n6392 VSS.n6391 1.43182
R8557 VSS.n6384 VSS.n6383 1.43182
R8558 VSS.n6364 VSS.n6363 1.43182
R8559 VSS.n6331 VSS.n6330 1.43182
R8560 VSS.n7264 VSS.n7263 1.43182
R8561 VSS.n6830 VSS.n6829 1.43182
R8562 VSS.n6836 VSS.n6835 1.43182
R8563 VSS.n6839 VSS.n6838 1.43182
R8564 VSS.n6845 VSS.n6844 1.43182
R8565 VSS.n6720 VSS.n6719 1.43182
R8566 VSS.n6702 VSS.n6701 1.43182
R8567 VSS.n5361 VSS.n5360 1.43182
R8568 VSS.n7635 VSS.n7634 1.43182
R8569 VSS.n7640 VSS.n7639 1.43182
R8570 VSS.n6361 VSS.n6360 1.43182
R8571 VSS.n7592 VSS.t760 1.42907
R8572 VSS.n4347 VSS.n4341 1.41664
R8573 VSS.n4092 VSS.n1868 1.38752
R8574 VSS.n4582 VSS.n4580 1.36161
R8575 VSS.n787 VSS.n786 1.33389
R8576 VSS.n29 VSS.n28 1.33375
R8577 VSS.n4736 VSS.n4735 1.33375
R8578 VSS.n4730 VSS.n4729 1.33375
R8579 VSS.n4721 VSS.n4720 1.33375
R8580 VSS.n4714 VSS.n4713 1.33375
R8581 VSS.n392 VSS.n391 1.32883
R8582 VSS.n511 VSS.n510 1.32883
R8583 VSS.n5 VSS.n4 1.32883
R8584 VSS.n499 VSS.n498 1.32869
R8585 VSS.n380 VSS.n379 1.32869
R8586 VSS.n8 VSS.n7 1.32869
R8587 VSS.n5378 VSS.n5377 1.32869
R8588 VSS.n7477 VSS.n7476 1.32869
R8589 VSS.n4904 VSS.n4903 1.28711
R8590 VSS.n5928 VSS.n5927 1.27022
R8591 VSS.n4547 VSS.n4538 1.26439
R8592 VSS.n4568 VSS.n4565 1.26439
R8593 VSS.n5626 VSS.n5611 1.22037
R8594 VSS.n3888 VSS.n3887 1.2005
R8595 VSS.n5784 VSS.n5781 1.18179
R8596 VSS.n5784 VSS.n5782 1.18179
R8597 VSS.n5784 VSS.n5783 1.18179
R8598 VSS.n5657 VSS.n5650 1.18179
R8599 VSS.n5657 VSS.n5651 1.18179
R8600 VSS.n5657 VSS.n5652 1.18179
R8601 VSS.n5657 VSS.n5653 1.18179
R8602 VSS.n5657 VSS.n5654 1.18179
R8603 VSS.n5657 VSS.n5655 1.18179
R8604 VSS.n5657 VSS.n5656 1.18179
R8605 VSS.n4391 VSS.n4387 1.16717
R8606 VSS.n1935 VSS.n1934 1.16276
R8607 VSS.n1934 VSS.n1933 1.16276
R8608 VSS.n1933 VSS.n1932 1.16276
R8609 VSS.n1932 VSS.n1931 1.16276
R8610 VSS.n1931 VSS.n1930 1.16276
R8611 VSS.n1930 VSS.n1929 1.16276
R8612 VSS.n1929 VSS.n1928 1.16276
R8613 VSS.n1928 VSS.n1927 1.16276
R8614 VSS.n1927 VSS.n1926 1.16276
R8615 VSS.n1926 VSS.n1925 1.16276
R8616 VSS.n2632 VSS.n2631 1.16276
R8617 VSS.n2631 VSS.n2630 1.16276
R8618 VSS.n2630 VSS.n2629 1.16276
R8619 VSS.n2629 VSS.n2628 1.16276
R8620 VSS.n2628 VSS.n2627 1.16276
R8621 VSS.n2627 VSS.n2626 1.16276
R8622 VSS.n2626 VSS.n2625 1.16276
R8623 VSS.n2625 VSS.n2624 1.16276
R8624 VSS.n2624 VSS.n2623 1.16276
R8625 VSS.n2623 VSS.n2622 1.16276
R8626 VSS.n2541 VSS.n2540 1.16276
R8627 VSS.n2540 VSS.n2539 1.16276
R8628 VSS.n2539 VSS.n2538 1.16276
R8629 VSS.n2538 VSS.n2537 1.16276
R8630 VSS.n2537 VSS.n2536 1.16276
R8631 VSS.n2536 VSS.n2535 1.16276
R8632 VSS.n2535 VSS.n2534 1.16276
R8633 VSS.n2534 VSS.n2533 1.16276
R8634 VSS.n2533 VSS.n2532 1.16276
R8635 VSS.n2532 VSS.n2531 1.16276
R8636 VSS.n2431 VSS.n2430 1.16276
R8637 VSS.n2430 VSS.n2429 1.16276
R8638 VSS.n2429 VSS.n2428 1.16276
R8639 VSS.n2428 VSS.n2427 1.16276
R8640 VSS.n2427 VSS.n2426 1.16276
R8641 VSS.n2426 VSS.n2425 1.16276
R8642 VSS.n2425 VSS.n2424 1.16276
R8643 VSS.n2424 VSS.n2423 1.16276
R8644 VSS.n2423 VSS.n2422 1.16276
R8645 VSS.n2422 VSS.n2421 1.16276
R8646 VSS.n2309 VSS.n2308 1.16276
R8647 VSS.n2308 VSS.n2307 1.16276
R8648 VSS.n2307 VSS.n2306 1.16276
R8649 VSS.n2306 VSS.n2305 1.16276
R8650 VSS.n2305 VSS.n2304 1.16276
R8651 VSS.n2304 VSS.n2303 1.16276
R8652 VSS.n2303 VSS.n2302 1.16276
R8653 VSS.n2302 VSS.n2301 1.16276
R8654 VSS.n2301 VSS.n2300 1.16276
R8655 VSS.n2300 VSS.n2299 1.16276
R8656 VSS.n2197 VSS.n2196 1.16276
R8657 VSS.n2196 VSS.n2195 1.16276
R8658 VSS.n2195 VSS.n2194 1.16276
R8659 VSS.n2194 VSS.n2193 1.16276
R8660 VSS.n2193 VSS.n2192 1.16276
R8661 VSS.n2192 VSS.n2191 1.16276
R8662 VSS.n2191 VSS.n2190 1.16276
R8663 VSS.n2190 VSS.n2189 1.16276
R8664 VSS.n2189 VSS.n2188 1.16276
R8665 VSS.n2188 VSS.n2187 1.16276
R8666 VSS.n2136 VSS.n2135 1.16276
R8667 VSS.n2135 VSS.n2134 1.16276
R8668 VSS.n2134 VSS.n2133 1.16276
R8669 VSS.n2133 VSS.n2132 1.16276
R8670 VSS.n2132 VSS.n2131 1.16276
R8671 VSS.n2131 VSS.n2130 1.16276
R8672 VSS.n2130 VSS.n2129 1.16276
R8673 VSS.n2129 VSS.n2128 1.16276
R8674 VSS.n2128 VSS.n2127 1.16276
R8675 VSS.n2127 VSS.n2126 1.16276
R8676 VSS.n1981 VSS.n1980 1.16276
R8677 VSS.n1980 VSS.n1979 1.16276
R8678 VSS.n1979 VSS.n1978 1.16276
R8679 VSS.n1978 VSS.n1977 1.16276
R8680 VSS.n1977 VSS.n1976 1.16276
R8681 VSS.n1976 VSS.n1975 1.16276
R8682 VSS.n1975 VSS.n1974 1.16276
R8683 VSS.n1974 VSS.n1973 1.16276
R8684 VSS.n1973 VSS.n1972 1.16276
R8685 VSS.n1972 VSS.n1971 1.16276
R8686 VSS.n1957 VSS.n1956 1.16276
R8687 VSS.n1956 VSS.n1955 1.16276
R8688 VSS.n1955 VSS.n1954 1.16276
R8689 VSS.n1954 VSS.n1953 1.16276
R8690 VSS.n1953 VSS.n1952 1.16276
R8691 VSS.n1952 VSS.n1951 1.16276
R8692 VSS.n1951 VSS.n1950 1.16276
R8693 VSS.n1950 VSS.n1949 1.16276
R8694 VSS.n1949 VSS.n1948 1.16276
R8695 VSS.n1948 VSS.n1947 1.16276
R8696 VSS.n1946 VSS.n1945 1.16276
R8697 VSS.n1945 VSS.n1944 1.16276
R8698 VSS.n1944 VSS.n1943 1.16276
R8699 VSS.n1943 VSS.n1942 1.16276
R8700 VSS.n1942 VSS.n1941 1.16276
R8701 VSS.n1941 VSS.n1940 1.16276
R8702 VSS.n1940 VSS.n1939 1.16276
R8703 VSS.n1939 VSS.n1938 1.16276
R8704 VSS.n1938 VSS.n1937 1.16276
R8705 VSS.n1937 VSS.n1936 1.16276
R8706 VSS.n3876 VSS.n3875 1.16276
R8707 VSS.n3877 VSS.n3876 1.16276
R8708 VSS.n3878 VSS.n3877 1.16276
R8709 VSS.n3879 VSS.n3878 1.16276
R8710 VSS.n3880 VSS.n3879 1.16276
R8711 VSS.n3881 VSS.n3880 1.16276
R8712 VSS.n3882 VSS.n3881 1.16276
R8713 VSS.n3883 VSS.n3882 1.16276
R8714 VSS.n3884 VSS.n3883 1.16276
R8715 VSS.n3885 VSS.n3884 1.16276
R8716 VSS.n3886 VSS.n3885 1.16276
R8717 VSS.n5632 VSS.n5572 1.15537
R8718 VSS.n3760 VSS.n3759 1.13934
R8719 VSS.n2669 VSS.n2652 1.12652
R8720 VSS.n147 VSS.n143 1.12642
R8721 VSS.n3952 VSS.n3947 1.1255
R8722 VSS.n3972 VSS.n3971 1.1255
R8723 VSS.n3916 VSS.n3911 1.1255
R8724 VSS.n3939 VSS.n3938 1.1255
R8725 VSS.n3985 VSS.n3981 1.1255
R8726 VSS.n3899 VSS.n3898 1.1255
R8727 VSS.n3700 VSS.n3699 1.1255
R8728 VSS.n2992 VSS.n2174 1.1255
R8729 VSS.n2182 VSS.n2175 1.1255
R8730 VSS.n2960 VSS.n2216 1.1255
R8731 VSS.n2962 VSS.n2213 1.1255
R8732 VSS.n3009 VSS.n2158 1.1255
R8733 VSS.n3004 VSS.n2160 1.1255
R8734 VSS.n2184 VSS.n2183 1.1255
R8735 VSS.n2961 VSS.n2214 1.1255
R8736 VSS.n2155 VSS.n2147 1.1255
R8737 VSS.n2926 VSS.n2925 1.1255
R8738 VSS.n2288 VSS.n2268 1.1255
R8739 VSS.n2344 VSS.n2323 1.1255
R8740 VSS.n2343 VSS.n2322 1.1255
R8741 VSS.n2907 VSS.n2280 1.1255
R8742 VSS.n2257 VSS.n2254 1.1255
R8743 VSS.n2351 VSS.n2324 1.1255
R8744 VSS.n2848 VSS.n2384 1.1255
R8745 VSS.n2457 VSS.n2443 1.1255
R8746 VSS.n2410 VSS.n2378 1.1255
R8747 VSS.n2837 VSS.n2399 1.1255
R8748 VSS.n2836 VSS.n2835 1.1255
R8749 VSS.n2411 VSS.n2379 1.1255
R8750 VSS.n2464 VSS.n2444 1.1255
R8751 VSS.n2404 VSS.n2370 1.1255
R8752 VSS.n2792 VSS.n2791 1.1255
R8753 VSS.n2568 VSS.n2550 1.1255
R8754 VSS.n2519 VSS.n2504 1.1255
R8755 VSS.n2746 VSS.n2557 1.1255
R8756 VSS.n2569 VSS.n2556 1.1255
R8757 VSS.n2521 VSS.n2520 1.1255
R8758 VSS.n2767 VSS.n2766 1.1255
R8759 VSS.n2784 VSS.n2498 1.1255
R8760 VSS.n2483 VSS.n2481 1.1255
R8761 VSS.n2481 VSS.n2477 1.1255
R8762 VSS.n2707 VSS.n2592 1.1255
R8763 VSS.n2668 VSS.n2667 1.1255
R8764 VSS.n2690 VSS.n2603 1.1255
R8765 VSS.n2670 VSS.n2646 1.1255
R8766 VSS.n2672 VSS.n2671 1.1255
R8767 VSS.n2693 VSS.n2601 1.1255
R8768 VSS.n2589 VSS.n2579 1.1255
R8769 VSS.n2650 VSS.n2612 1.1255
R8770 VSS.n2685 VSS.n2612 1.1255
R8771 VSS.n2575 VSS.n2574 1.1255
R8772 VSS.n2673 VSS.n2672 1.1255
R8773 VSS.n2674 VSS.n2673 1.1255
R8774 VSS.n2599 VSS.n2597 1.1255
R8775 VSS.n2601 VSS.n2599 1.1255
R8776 VSS.n2646 VSS.n2643 1.1255
R8777 VSS.n2643 VSS.n2642 1.1255
R8778 VSS.n2689 VSS.n2688 1.1255
R8779 VSS.n2690 VSS.n2689 1.1255
R8780 VSS.n2574 VSS.n2573 1.1255
R8781 VSS.n2715 VSS.n2581 1.1255
R8782 VSS.n2581 VSS.n2579 1.1255
R8783 VSS.n2666 VSS.n2665 1.1255
R8784 VSS.n2667 VSS.n2666 1.1255
R8785 VSS.n2685 VSS.n2610 1.1255
R8786 VSS.n2800 VSS.n2477 1.1255
R8787 VSS.n2566 VSS.n2564 1.1255
R8788 VSS.n2556 VSS.n2551 1.1255
R8789 VSS.n2520 VSS.n2505 1.1255
R8790 VSS.n2765 VSS.n2764 1.1255
R8791 VSS.n2766 VSS.n2765 1.1255
R8792 VSS.n2748 VSS.n2747 1.1255
R8793 VSS.n2747 VSS.n2746 1.1255
R8794 VSS.n2785 VSS.n2490 1.1255
R8795 VSS.n2785 VSS.n2784 1.1255
R8796 VSS.n2777 VSS.n2504 1.1255
R8797 VSS.n2751 VSS.n2550 1.1255
R8798 VSS.n2777 VSS.n2776 1.1255
R8799 VSS.n2751 VSS.n2750 1.1255
R8800 VSS.n2790 VSS.n2789 1.1255
R8801 VSS.n2791 VSS.n2790 1.1255
R8802 VSS.n2470 VSS.n2469 1.1255
R8803 VSS.n2471 VSS.n2470 1.1255
R8804 VSS.n2775 VSS.n2505 1.1255
R8805 VSS.n2749 VSS.n2551 1.1255
R8806 VSS.n2572 VSS.n2564 1.1255
R8807 VSS.n2362 VSS.n2361 1.1255
R8808 VSS.n2856 VSS.n2378 1.1255
R8809 VSS.n2822 VSS.n2444 1.1255
R8810 VSS.n2823 VSS.n2443 1.1255
R8811 VSS.n2815 VSS.n2814 1.1255
R8812 VSS.n2814 VSS.n2813 1.1255
R8813 VSS.n2432 VSS.n2419 1.1255
R8814 VSS.n2419 VSS.n2399 1.1255
R8815 VSS.n2855 VSS.n2379 1.1255
R8816 VSS.n2835 VSS.n2834 1.1255
R8817 VSS.n2864 VSS.n2370 1.1255
R8818 VSS.n2848 VSS.n2847 1.1255
R8819 VSS.n2847 VSS.n2846 1.1255
R8820 VSS.n2824 VSS.n2823 1.1255
R8821 VSS.n2865 VSS.n2864 1.1255
R8822 VSS.n2855 VSS.n2377 1.1255
R8823 VSS.n2834 VSS.n2833 1.1255
R8824 VSS.n2822 VSS.n2442 1.1255
R8825 VSS.n2857 VSS.n2856 1.1255
R8826 VSS.n2361 VSS.n2360 1.1255
R8827 VSS.n2933 VSS.n2254 1.1255
R8828 VSS.n2911 VSS.n2278 1.1255
R8829 VSS.n2888 VSS.n2324 1.1255
R8830 VSS.n2907 VSS.n2279 1.1255
R8831 VSS.n2879 VSS.n2355 1.1255
R8832 VSS.n2890 VSS.n2322 1.1255
R8833 VSS.n2891 VSS.n2890 1.1255
R8834 VSS.n2879 VSS.n2878 1.1255
R8835 VSS.n2889 VSS.n2323 1.1255
R8836 VSS.n2919 VSS.n2268 1.1255
R8837 VSS.n2903 VSS.n2902 1.1255
R8838 VSS.n2246 VSS.n2245 1.1255
R8839 VSS.n2925 VSS.n2924 1.1255
R8840 VSS.n2310 VSS.n2279 1.1255
R8841 VSS.n2924 VSS.n2923 1.1255
R8842 VSS.n2889 VSS.n2320 1.1255
R8843 VSS.n2245 VSS.n2244 1.1255
R8844 VSS.n2919 VSS.n2265 1.1255
R8845 VSS.n2902 VSS.n2901 1.1255
R8846 VSS.n2888 VSS.n2887 1.1255
R8847 VSS.n2912 VSS.n2911 1.1255
R8848 VSS.n2934 VSS.n2933 1.1255
R8849 VSS.n2961 VSS.n2209 1.1255
R8850 VSS.n2186 VSS.n2184 1.1255
R8851 VSS.n3015 VSS.n2147 1.1255
R8852 VSS.n2177 VSS.n2175 1.1255
R8853 VSS.n2949 VSS.n2948 1.1255
R8854 VSS.n2963 VSS.n2212 1.1255
R8855 VSS.n2963 VSS.n2962 1.1255
R8856 VSS.n2948 VSS.n2947 1.1255
R8857 VSS.n2959 VSS.n2958 1.1255
R8858 VSS.n2960 VSS.n2959 1.1255
R8859 VSS.n2138 VSS.n2137 1.1255
R8860 VSS.n2139 VSS.n2138 1.1255
R8861 VSS.n2989 VSS.n2177 1.1255
R8862 VSS.n3010 VSS.n2154 1.1255
R8863 VSS.n3010 VSS.n3009 1.1255
R8864 VSS.n3004 VSS.n3003 1.1255
R8865 VSS.n2992 VSS.n2991 1.1255
R8866 VSS.n2991 VSS.n2990 1.1255
R8867 VSS.n3016 VSS.n3015 1.1255
R8868 VSS.n3003 VSS.n3002 1.1255
R8869 VSS.n2976 VSS.n2186 1.1255
R8870 VSS.n2218 VSS.n2209 1.1255
R8871 VSS.n2023 VSS.n1998 1.1255
R8872 VSS.n2034 VSS.n1997 1.1255
R8873 VSS.n2042 VSS.n1982 1.1255
R8874 VSS.n2076 VSS.n2075 1.1255
R8875 VSS.n2041 VSS.n1988 1.1255
R8876 VSS.n2066 VSS.n2065 1.1255
R8877 VSS.n2022 VSS.n2007 1.1255
R8878 VSS.n2013 VSS.n2012 1.1255
R8879 VSS.n2025 VSS.n2024 1.1255
R8880 VSS.n2056 VSS.n2055 1.1255
R8881 VSS.n2124 VSS.n2123 1.1255
R8882 VSS.n3128 VSS.n3127 1.1255
R8883 VSS.n3159 VSS.n3156 1.1255
R8884 VSS.n3172 VSS.n3167 1.1255
R8885 VSS.n3223 VSS.n3218 1.1255
R8886 VSS.n3182 VSS.n3181 1.1255
R8887 VSS.n3143 VSS.n3142 1.1255
R8888 VSS.n3106 VSS.n3104 1.1255
R8889 VSS.n3125 VSS.n3118 1.1255
R8890 VSS.n3193 VSS.n3189 1.1255
R8891 VSS.n3206 VSS.n3205 1.1255
R8892 VSS.n3126 VSS.n3125 1.1255
R8893 VSS.n3107 VSS.n3106 1.1255
R8894 VSS.n3144 VSS.n3143 1.1255
R8895 VSS.n3183 VSS.n3182 1.1255
R8896 VSS.n3224 VSS.n3223 1.1255
R8897 VSS.n3207 VSS.n3206 1.1255
R8898 VSS.n3173 VSS.n3172 1.1255
R8899 VSS.n3194 VSS.n3193 1.1255
R8900 VSS.n3160 VSS.n3159 1.1255
R8901 VSS.n3129 VSS.n3128 1.1255
R8902 VSS.n1967 VSS.n1963 1.1255
R8903 VSS.n3270 VSS.n3265 1.1255
R8904 VSS.n3308 VSS.n3307 1.1255
R8905 VSS.n3257 VSS.n3252 1.1255
R8906 VSS.n3301 VSS.n3300 1.1255
R8907 VSS.n3341 VSS.n3336 1.1255
R8908 VSS.n3325 VSS.n3320 1.1255
R8909 VSS.n3362 VSS.n3361 1.1255
R8910 VSS.n3285 VSS.n3280 1.1255
R8911 VSS.n3244 VSS.n3242 1.1255
R8912 VSS.n3363 VSS.n3362 1.1255
R8913 VSS.n3326 VSS.n3325 1.1255
R8914 VSS.n3286 VSS.n3285 1.1255
R8915 VSS.n3245 VSS.n3244 1.1255
R8916 VSS.n3352 VSS.n3351 1.1255
R8917 VSS.n3404 VSS.n3403 1.1255
R8918 VSS.n3405 VSS.n3404 1.1255
R8919 VSS.n3342 VSS.n3341 1.1255
R8920 VSS.n3302 VSS.n3301 1.1255
R8921 VSS.n3258 VSS.n3257 1.1255
R8922 VSS.n3353 VSS.n3352 1.1255
R8923 VSS.n3309 VSS.n3308 1.1255
R8924 VSS.n3271 VSS.n3270 1.1255
R8925 VSS.n3423 VSS.n3422 1.1255
R8926 VSS.n3459 VSS.n3458 1.1255
R8927 VSS.n3500 VSS.n3493 1.1255
R8928 VSS.n3529 VSS.n3528 1.1255
R8929 VSS.n3416 VSS.n3412 1.1255
R8930 VSS.n3463 VSS.n3462 1.1255
R8931 VSS.n3518 VSS.n3517 1.1255
R8932 VSS.n3584 VSS.n3583 1.1255
R8933 VSS.n3503 VSS.n3502 1.1255
R8934 VSS.n3479 VSS.n3476 1.1255
R8935 VSS.n3439 VSS.n3438 1.1255
R8936 VSS.n3504 VSS.n3503 1.1255
R8937 VSS.n3480 VSS.n3479 1.1255
R8938 VSS.n3440 VSS.n3439 1.1255
R8939 VSS.n3585 VSS.n3584 1.1255
R8940 VSS.n3519 VSS.n3518 1.1255
R8941 VSS.n3464 VSS.n3463 1.1255
R8942 VSS.n3417 VSS.n3416 1.1255
R8943 VSS.n3530 VSS.n3529 1.1255
R8944 VSS.n3501 VSS.n3500 1.1255
R8945 VSS.n3460 VSS.n3459 1.1255
R8946 VSS.n3424 VSS.n3423 1.1255
R8947 VSS.n1894 VSS.n1891 1.1255
R8948 VSS.n3872 VSS.n3871 1.1255
R8949 VSS.n1907 VSS.n1906 1.1255
R8950 VSS.n3818 VSS.n3817 1.1255
R8951 VSS.n3807 VSS.n3802 1.1255
R8952 VSS.n3836 VSS.n3835 1.1255
R8953 VSS.n1923 VSS.n1922 1.1255
R8954 VSS.n3793 VSS.n3791 1.1255
R8955 VSS.n1886 VSS.n1885 1.1255
R8956 VSS.n1887 VSS.n1886 1.1255
R8957 VSS.n1924 VSS.n1923 1.1255
R8958 VSS.n3837 VSS.n3836 1.1255
R8959 VSS.n3808 VSS.n3807 1.1255
R8960 VSS.n3794 VSS.n3793 1.1255
R8961 VSS.n3819 VSS.n3818 1.1255
R8962 VSS.n1908 VSS.n1907 1.1255
R8963 VSS.n3856 VSS.n3855 1.1255
R8964 VSS.n3855 VSS.n3854 1.1255
R8965 VSS.n3833 VSS.n3828 1.1255
R8966 VSS.n3834 VSS.n3833 1.1255
R8967 VSS.n3873 VSS.n3872 1.1255
R8968 VSS.n1895 VSS.n1894 1.1255
R8969 VSS.n3973 VSS.n3972 1.1255
R8970 VSS.n3940 VSS.n3939 1.1255
R8971 VSS.n3917 VSS.n3916 1.1255
R8972 VSS.n3986 VSS.n3985 1.1255
R8973 VSS.n3900 VSS.n3899 1.1255
R8974 VSS.n3953 VSS.n3952 1.1255
R8975 VSS.n1863 VSS.n1862 1.1255
R8976 VSS.n1531 VSS.n1530 1.1255
R8977 VSS.n215 VSS.n214 1.1255
R8978 VSS.n1587 VSS.n1586 1.1234
R8979 VSS.n1969 VSS.n1968 1.12321
R8980 VSS.n1775 VSS.n1774 1.12277
R8981 VSS.n1765 VSS.n1764 1.12277
R8982 VSS.n6740 VSS.n6738 1.11026
R8983 VSS.n6950 VSS.n6942 1.11026
R8984 VSS.n213 VSS.n212 1.09796
R8985 VSS.n4401 VSS.n4400 1.06994
R8986 VSS.n4391 VSS.n4390 1.06994
R8987 VSS.n517 VSS.n515 1.03151
R8988 VSS.n722 VSS.n720 1.02489
R8989 VSS.n1481 VSS.n1479 1.02489
R8990 VSS.n7245 VSS.n7243 1.02489
R8991 VSS.n6486 VSS.n6484 1.02489
R8992 VSS.t360 VSS.t511 1.01328
R8993 VSS.n5784 VSS.n5780 1.01328
R8994 VSS.t504 VSS.t413 1.01328
R8995 VSS.t413 VSS.t371 1.01328
R8996 VSS.n1365 VSS.n1253 1.0102
R8997 VSS.n7152 VSS.n7151 0.990549
R8998 VSS.n4547 VSS.n4545 0.972722
R8999 VSS.n4568 VSS.n4567 0.972722
R9000 VSS.n5238 VSS.n5237 0.967979
R9001 VSS.n3060 VSS.n2125 0.960694
R9002 VSS.n4546 VSS.t29 0.93818
R9003 VSS.n1402 VSS.n1401 0.93818
R9004 VSS.n1595 VSS.n1594 0.931667
R9005 VSS.n696 VSS.n695 0.929536
R9006 VSS.n686 VSS.n685 0.928071
R9007 VSS.n1534 VSS.n1533 0.925894
R9008 VSS.n4788 VSS.n4743 0.919029
R9009 VSS.n4723 VSS.n53 0.919029
R9010 VSS.n1136 VSS.n1135 0.910283
R9011 VSS.n1627 VSS.n1615 0.907678
R9012 VSS.n3790 VSS.n3789 0.900727
R9013 VSS.n2354 VSS.n2353 0.900647
R9014 VSS.n2467 VSS.n2466 0.900647
R9015 VSS.n1865 VSS.n1864 0.90054
R9016 VSS.n2291 VSS.n2278 0.9005
R9017 VSS.n2904 VSS.n2903 0.9005
R9018 VSS.n3398 VSS.n3397 0.900483
R9019 VSS.n2809 VSS.n2808 0.900483
R9020 VSS.n3241 VSS.n3240 0.900467
R9021 VSS.n3103 VSS.n3102 0.900467
R9022 VSS.n2730 VSS.n2729 0.900467
R9023 VSS.n3578 VSS.n3577 0.900443
R9024 VSS.n2724 VSS.n2723 0.900442
R9025 VSS.n2236 VSS.n2234 0.900387
R9026 VSS.n2011 VSS.n2010 0.900368
R9027 VSS.n3025 VSS.n3024 0.900365
R9028 VSS.n2943 VSS.n2942 0.900365
R9029 VSS.n2874 VSS.n2873 0.900365
R9030 VSS.n2118 VSS.n2117 0.900347
R9031 VSS.n1778 VSS.n1777 0.900305
R9032 VSS.n92 VSS.n91 0.898922
R9033 VSS.n1962 VSS.n1961 0.898321
R9034 VSS.n211 VSS.n205 0.897993
R9035 VSS.n4891 VSS.n4890 0.895873
R9036 VSS.n1867 VSS.n1866 0.891062
R9037 VSS.n4582 VSS.n4578 0.8755
R9038 VSS.n1624 VSS.n1621 0.869196
R9039 VSS.n4340 VSS.n4202 0.869196
R9040 VSS.n4333 VSS.n4332 0.869196
R9041 VSS.n391 VSS.n390 0.849401
R9042 VSS.n510 VSS.n509 0.849401
R9043 VSS.n786 VSS.n785 0.846031
R9044 VSS.n4720 VSS.n4719 0.845835
R9045 VSS.n4735 VSS.n4734 0.845835
R9046 VSS.n689 VSS.n681 0.830589
R9047 VSS.n7427 VSS.n7426 0.829048
R9048 VSS.n4217 VSS.t422 0.826268
R9049 VSS.n1736 VSS.t378 0.826268
R9050 VSS.n3889 VSS.n3888 0.811705
R9051 VSS.n4526 VSS.n4523 0.79929
R9052 VSS.n1714 VSS.n1711 0.793518
R9053 VSS.n4309 VSS.n4216 0.782913
R9054 VSS.n1723 VSS.n1722 0.782913
R9055 VSS.n6600 VSS.n6599 0.781777
R9056 VSS.n6608 VSS.n6607 0.781777
R9057 VSS.n4314 VSS.n4213 0.781543
R9058 VSS.n6471 VSS.n6470 0.780656
R9059 VSS.n7270 VSS.n7269 0.780656
R9060 VSS.n6336 VSS.n6335 0.780656
R9061 VSS.n812 VSS.n806 0.780656
R9062 VSS.n7308 VSS.n7307 0.780455
R9063 VSS.n7330 VSS.n7329 0.780455
R9064 VSS.n6391 VSS.n6390 0.780455
R9065 VSS.n6365 VSS.n6364 0.780455
R9066 VSS.n6365 VSS.n6361 0.780455
R9067 VSS.n6844 VSS.n6843 0.780455
R9068 VSS.n6835 VSS.n6834 0.780455
R9069 VSS.n6701 VSS.n6700 0.780455
R9070 VSS.n6719 VSS.n6718 0.780455
R9071 VSS.n1451 VSS.n1450 0.780455
R9072 VSS.n1379 VSS.n1378 0.780455
R9073 VSS.n812 VSS.n811 0.780455
R9074 VSS.n834 VSS.n833 0.780455
R9075 VSS.n1104 VSS.n1103 0.780455
R9076 VSS.n1604 VSS.n1603 0.778278
R9077 VSS.n7843 VSS.n7840 0.778278
R9078 VSS.n212 VSS.n211 0.768418
R9079 VSS.n4277 VSS.n4276 0.749848
R9080 VSS.n4592 VSS.n4590 0.726531
R9081 VSS.n4278 VSS.n4271 0.722457
R9082 VSS.n1677 VSS.n1673 0.722457
R9083 VSS.n4271 VSS.n4268 0.708761
R9084 VSS.n1673 VSS.n1670 0.708761
R9085 VSS.n4259 VSS.n4256 0.706804
R9086 VSS.n4262 VSS.n4259 0.706804
R9087 VSS.n4265 VSS.n4262 0.706804
R9088 VSS.n4268 VSS.n4265 0.706804
R9089 VSS.n1661 VSS.n1658 0.706804
R9090 VSS.n1664 VSS.n1661 0.706804
R9091 VSS.n1667 VSS.n1664 0.706804
R9092 VSS.n1670 VSS.n1667 0.706804
R9093 VSS.n1708 VSS.n1700 0.706804
R9094 VSS.n1614 VSS.n1613 0.706804
R9095 VSS.n4201 VSS.n4200 0.706804
R9096 VSS.n4329 VSS.n4328 0.706804
R9097 VSS.n4210 VSS.n4207 0.706804
R9098 VSS.n1708 VSS.n1707 0.704848
R9099 VSS.n1137 VSS.n1133 0.692793
R9100 VSS VSS.n7907 0.683795
R9101 VSS.n1548 VSS.n1500 0.681056
R9102 VSS.n4276 VSS.n4216 0.679996
R9103 VSS.n1722 VSS.n1719 0.679996
R9104 VSS.n1711 VSS.n1708 0.679954
R9105 VSS.n4213 VSS.n4210 0.679954
R9106 VSS.n1621 VSS.n1618 0.679913
R9107 VSS.n1615 VSS.n1614 0.679913
R9108 VSS.n4202 VSS.n4201 0.679913
R9109 VSS.n4332 VSS.n4329 0.679913
R9110 VSS.n6985 VSS.t568 0.678722
R9111 VSS.n4139 VSS.n4131 0.675114
R9112 VSS.n6986 VSS.t572 0.673472
R9113 VSS.n6987 VSS.t569 0.673472
R9114 VSS.n5083 VSS.n5082 0.66722
R9115 VSS.n5102 VSS.n5101 0.66722
R9116 VSS.n5210 VSS.n5209 0.66722
R9117 VSS.n7852 VSS.n7851 0.66722
R9118 VSS.n5785 VSS.n5784 0.66722
R9119 VSS.n5658 VSS.n5657 0.66722
R9120 VSS.n7869 VSS.n7868 0.66722
R9121 VSS.n1747 VSS.n1746 0.659848
R9122 VSS.n4301 VSS.n4284 0.654826
R9123 VSS.n1689 VSS.n1686 0.654826
R9124 VSS.n4036 VSS.n4029 0.652915
R9125 VSS.n4394 VSS.t252 0.65037
R9126 VSS.n7143 VSS.n7142 0.644196
R9127 VSS.n4008 VSS.n1872 0.643803
R9128 VSS.n5832 VSS.n5831 0.642239
R9129 VSS.n5436 VSS.n5435 0.642239
R9130 VSS.n5418 VSS.n5417 0.642239
R9131 VSS.n4972 VSS.n4969 0.642239
R9132 VSS.n4959 VSS.n4956 0.642239
R9133 VSS.n5012 VSS.n5009 0.642239
R9134 VSS.n2975 VSS.n2197 0.615498
R9135 VSS.n2312 VSS.n2309 0.614262
R9136 VSS.n4892 VSS.n4868 0.611348
R9137 VSS.n6175 VSS.n6174 0.610998
R9138 VSS.n2433 VSS.n2431 0.609999
R9139 VSS.n3602 VSS.n1935 0.609008
R9140 VSS.n3148 VSS.n1981 0.608439
R9141 VSS.n3875 VSS.n3874 0.606848
R9142 VSS.n2763 VSS.n2541 0.606843
R9143 VSS.n3311 VSS.n1957 0.606489
R9144 VSS.n3481 VSS.n1946 0.605607
R9145 VSS.n3041 VSS.n2136 0.601243
R9146 VSS.n5417 VSS.n5416 0.597879
R9147 VSS.n5009 VSS.n5006 0.597879
R9148 VSS.n5435 VSS.n5434 0.596788
R9149 VSS.n4969 VSS.n4966 0.596788
R9150 VSS.n5831 VSS.n5830 0.595696
R9151 VSS.n4956 VSS.n4953 0.595696
R9152 VSS.n7428 VSS.n7427 0.594669
R9153 VSS.n2633 VSS.n2632 0.593624
R9154 VSS.n5829 VSS.n5828 0.587128
R9155 VSS.n4963 VSS.n4962 0.586903
R9156 VSS.n5433 VSS.n5432 0.586037
R9157 VSS.n5003 VSS.n5002 0.585812
R9158 VSS.n4212 VSS.t322 0.5855
R9159 VSS.n4212 VSS.n4211 0.5855
R9160 VSS.n4255 VSS.t289 0.5855
R9161 VSS.n4255 VSS.n4254 0.5855
R9162 VSS.n4258 VSS.t182 0.5855
R9163 VSS.n4258 VSS.n4257 0.5855
R9164 VSS.n4261 VSS.t215 0.5855
R9165 VSS.n4261 VSS.n4260 0.5855
R9166 VSS.n4264 VSS.t196 0.5855
R9167 VSS.n4264 VSS.n4263 0.5855
R9168 VSS.n4267 VSS.t317 0.5855
R9169 VSS.n4267 VSS.n4266 0.5855
R9170 VSS.n4270 VSS.t174 0.5855
R9171 VSS.n4270 VSS.n4269 0.5855
R9172 VSS.n4273 VSS.t324 0.5855
R9173 VSS.n4273 VSS.n4272 0.5855
R9174 VSS.n4250 VSS.t402 0.5855
R9175 VSS.n4236 VSS.t495 0.5855
R9176 VSS.n4235 VSS.t404 0.5855
R9177 VSS.n4234 VSS.t438 0.5855
R9178 VSS.n4232 VSS.t353 0.5855
R9179 VSS.n4230 VSS.t394 0.5855
R9180 VSS.n4228 VSS.t488 0.5855
R9181 VSS.n4226 VSS.t514 0.5855
R9182 VSS.n4224 VSS.t380 0.5855
R9183 VSS.n4222 VSS.t478 0.5855
R9184 VSS.n4220 VSS.t516 0.5855
R9185 VSS.n4252 VSS.t363 0.5855
R9186 VSS.n4252 VSS.n4251 0.5855
R9187 VSS.n4275 VSS.t186 0.5855
R9188 VSS.n4275 VSS.n4274 0.5855
R9189 VSS.n4215 VSS.t218 0.5855
R9190 VSS.n4215 VSS.n4214 0.5855
R9191 VSS.n4204 VSS.t188 0.5855
R9192 VSS.n4204 VSS.n4203 0.5855
R9193 VSS.n4206 VSS.t219 0.5855
R9194 VSS.n4206 VSS.n4205 0.5855
R9195 VSS.n4323 VSS.t517 0.5855
R9196 VSS.n4323 VSS.n4322 0.5855
R9197 VSS.n4331 VSS.t217 0.5855
R9198 VSS.n4331 VSS.n4330 0.5855
R9199 VSS.n1718 VSS.t521 0.5855
R9200 VSS.n1718 VSS.n1717 0.5855
R9201 VSS.n1721 VSS.t49 0.5855
R9202 VSS.n1721 VSS.n1720 0.5855
R9203 VSS.n1654 VSS.t497 0.5855
R9204 VSS.n1640 VSS.t491 0.5855
R9205 VSS.n1639 VSS.t471 0.5855
R9206 VSS.n1685 VSS.t484 0.5855
R9207 VSS.n1685 VSS.t493 0.5855
R9208 VSS.n1637 VSS.t465 0.5855
R9209 VSS.n1635 VSS.t445 0.5855
R9210 VSS.n1633 VSS.t411 0.5855
R9211 VSS.n1742 VSS.t457 0.5855
R9212 VSS.n1741 VSS.t366 0.5855
R9213 VSS.n1741 VSS.t383 0.5855
R9214 VSS.n1739 VSS.t355 0.5855
R9215 VSS.n1679 VSS.n1678 0.5855
R9216 VSS.n1657 VSS.t771 0.5855
R9217 VSS.n1657 VSS.n1656 0.5855
R9218 VSS.n1660 VSS.t764 0.5855
R9219 VSS.n1660 VSS.n1659 0.5855
R9220 VSS.n1663 VSS.t843 0.5855
R9221 VSS.n1663 VSS.n1662 0.5855
R9222 VSS.n1666 VSS.t102 0.5855
R9223 VSS.n1666 VSS.n1665 0.5855
R9224 VSS.n1669 VSS.t889 0.5855
R9225 VSS.n1669 VSS.n1668 0.5855
R9226 VSS.n1672 VSS.t305 0.5855
R9227 VSS.n1672 VSS.n1671 0.5855
R9228 VSS.n1675 VSS.t47 0.5855
R9229 VSS.n1675 VSS.n1674 0.5855
R9230 VSS.n1697 VSS.t846 0.5855
R9231 VSS.n1697 VSS.n1696 0.5855
R9232 VSS.n1699 VSS.t100 0.5855
R9233 VSS.n1699 VSS.n1698 0.5855
R9234 VSS.n1702 VSS.t13 0.5855
R9235 VSS.n1702 VSS.n1701 0.5855
R9236 VSS.n1710 VSS.t522 0.5855
R9237 VSS.n1710 VSS.n1709 0.5855
R9238 VSS.n1704 VSS.t109 0.5855
R9239 VSS.n1704 VSS.n1703 0.5855
R9240 VSS.n1706 VSS.t768 0.5855
R9241 VSS.n1706 VSS.n1705 0.5855
R9242 VSS.n1617 VSS.t89 0.5855
R9243 VSS.n1617 VSS.n1616 0.5855
R9244 VSS.n1620 VSS.t518 0.5855
R9245 VSS.n1620 VSS.n1619 0.5855
R9246 VSS.n1610 VSS.t11 0.5855
R9247 VSS.n1610 VSS.n1609 0.5855
R9248 VSS.n1612 VSS.t893 0.5855
R9249 VSS.n1612 VSS.n1611 0.5855
R9250 VSS.n4197 VSS.t716 0.5855
R9251 VSS.n4197 VSS.n4196 0.5855
R9252 VSS.n4199 VSS.t315 0.5855
R9253 VSS.n4199 VSS.n4198 0.5855
R9254 VSS.n4325 VSS.t906 0.5855
R9255 VSS.n4325 VSS.n4324 0.5855
R9256 VSS.n4327 VSS.t184 0.5855
R9257 VSS.n4327 VSS.n4326 0.5855
R9258 VSS.n4209 VSS.t170 0.5855
R9259 VSS.n4209 VSS.n4208 0.5855
R9260 VSS.n5413 VSS.n5412 0.584946
R9261 VSS.n644 VSS.n643 0.583833
R9262 VSS.n5432 VSS.n5431 0.574718
R9263 VSS.n5412 VSS.n5411 0.573627
R9264 VSS.n5002 VSS.n4999 0.573197
R9265 VSS.n3701 VSS.n3700 0.563
R9266 VSS.n2707 VSS.n2588 0.563
R9267 VSS.n2588 VSS.n2586 0.563
R9268 VSS.n2596 VSS.n2586 0.563
R9269 VSS.n3737 VSS.n3701 0.563
R9270 VSS.n3738 VSS.n3737 0.563
R9271 VSS.n1139 VSS.n1138 0.561716
R9272 VSS.n7887 VSS.n7886 0.561716
R9273 VSS.n7894 VSS.n7893 0.561716
R9274 VSS.n11 VSS.n10 0.561716
R9275 VSS.n5257 VSS.n5256 0.561716
R9276 VSS.n5266 VSS.n5265 0.561716
R9277 VSS.n5296 VSS.n5295 0.561716
R9278 VSS.n1789 VSS.n1788 0.551597
R9279 VSS.n5828 VSS.n5827 0.550283
R9280 VSS.n4890 VSS.n4889 0.550283
R9281 VSS.n4891 VSS.n4884 0.54076
R9282 VSS.n6938 VSS.n5354 0.525217
R9283 VSS.n5373 VSS.n5369 0.522718
R9284 VSS.n7738 VSS.n7733 0.522718
R9285 VSS.n7736 VSS.n7735 0.508005
R9286 VSS.n7432 VSS.n7431 0.508005
R9287 VSS.n5373 VSS.n5372 0.508005
R9288 VSS.n7738 VSS.n7737 0.508005
R9289 VSS.n7485 VSS.n5359 0.508005
R9290 VSS.n5388 VSS.n5387 0.508005
R9291 VSS.n5386 VSS.n5385 0.508005
R9292 VSS.n6277 VSS.n6276 0.508005
R9293 VSS.n6276 VSS.n6275 0.507764
R9294 VSS.n6276 VSS.n6274 0.507764
R9295 VSS.n6276 VSS.n6273 0.507764
R9296 VSS.n329 VSS.n328 0.507764
R9297 VSS.n325 VSS.n324 0.505601
R9298 VSS.n4705 VSS.n4704 0.505601
R9299 VSS.n797 VSS.n796 0.50536
R9300 VSS.n7486 VSS.n7485 0.502758
R9301 VSS.n769 VSS.n768 0.502377
R9302 VSS.n5899 VSS.n5898 0.502362
R9303 VSS.n4882 VSS.n4881 0.502362
R9304 VSS.n4879 VSS.n4878 0.497425
R9305 VSS.n5902 VSS.n5901 0.497402
R9306 VSS.n4414 VSS.n4413 0.486611
R9307 VSS.n6979 VSS.n6609 0.477891
R9308 VSS.n3407 VSS.n3406 0.473104
R9309 VSS.n746 VSS.n745 0.472687
R9310 VSS.n4525 VSS.n4524 0.472687
R9311 VSS.n2812 VSS.n2811 0.467151
R9312 VSS.n3587 VSS.n3586 0.465504
R9313 VSS.n1408 VSS.n1407 0.459689
R9314 VSS.n5369 VSS.n5368 0.459689
R9315 VSS.n7733 VSS.n7732 0.459689
R9316 VSS.n7731 VSS.n7730 0.459689
R9317 VSS.n7276 VSS.n7275 0.459689
R9318 VSS.n6386 VSS.n6382 0.459689
R9319 VSS.n6377 VSS.n6373 0.459689
R9320 VSS.n7419 VSS.n7418 0.459689
R9321 VSS.n6991 VSS.n6990 0.459689
R9322 VSS.n6350 VSS.n6342 0.459689
R9323 VSS.n6340 VSS.n6339 0.459689
R9324 VSS.n6960 VSS.n6959 0.459689
R9325 VSS.n7529 VSS.n7528 0.459689
R9326 VSS.n4506 VSS.n4505 0.459689
R9327 VSS.n1094 VSS.n1093 0.459689
R9328 VSS.n1132 VSS.n1131 0.459689
R9329 VSS.n781 VSS.n780 0.459446
R9330 VSS.n6864 VSS.n6863 0.459446
R9331 VSS.n7665 VSS.n7664 0.459446
R9332 VSS.n3992 VSS.n3991 0.459227
R9333 VSS.n3061 VSS.n3060 0.458913
R9334 VSS.n6980 VSS.n6602 0.458326
R9335 VSS.n2877 VSS.n2876 0.456584
R9336 VSS.n2946 VSS.n2945 0.451624
R9337 VSS.n2727 VSS.n2726 0.449946
R9338 VSS.n1487 VSS 0.449668
R9339 VSS.n7144 VSS.n7143 0.449473
R9340 VSS.n4422 VSS.n4421 0.447284
R9341 VSS.n3227 VSS.n3226 0.443676
R9342 VSS.n3745 VSS.n3744 0.441768
R9343 VSS.n4938 VSS.n4937 0.435547
R9344 VSS.n5769 VSS.n5768 0.434956
R9345 VSS.n4506 VSS.n4500 0.4313
R9346 VSS.n5397 VSS.n5394 0.426043
R9347 VSS VSS.n1486 0.405813
R9348 VSS.n4497 VSS.n4496 0.402035
R9349 VSS.n303 VSS.n302 0.402035
R9350 VSS.n4498 VSS.n4497 0.402035
R9351 VSS.n4139 VSS.n4136 0.402035
R9352 VSS.n4143 VSS.n4142 0.402035
R9353 VSS.n318 VSS.n317 0.402035
R9354 VSS.n4663 VSS.n4662 0.402035
R9355 VSS.n4661 VSS.n4660 0.402035
R9356 VSS.n4697 VSS.n4696 0.402035
R9357 VSS.n4500 VSS.n4499 0.402035
R9358 VSS.n4347 VSS.n4346 0.402035
R9359 VSS.n4627 VSS.n4626 0.401791
R9360 VSS.n7426 VSS.n7425 0.39444
R9361 VSS.n6119 VSS.n6116 0.393137
R9362 VSS.n7880 VSS.n7877 0.393137
R9363 VSS.n6182 VSS.n6103 0.391771
R9364 VSS.n75 VSS.n72 0.390642
R9365 VSS.n562 VSS.n559 0.390642
R9366 VSS.n325 VSS.n318 0.390642
R9367 VSS.n4700 VSS.n4697 0.390642
R9368 VSS.n5239 VSS.n5238 0.383479
R9369 VSS.n43 VSS.n42 0.383166
R9370 VSS.n4771 VSS.n4770 0.383166
R9371 VSS.n5399 VSS.n5398 0.383166
R9372 VSS.n5119 VSS.n5118 0.383166
R9373 VSS.n7875 VSS.n7874 0.383166
R9374 VSS.n4785 VSS.n4784 0.382921
R9375 VSS.n5117 VSS.n22 0.376519
R9376 VSS.n5096 VSS.n4923 0.376518
R9377 VSS.n5721 VSS.n5720 0.37489
R9378 VSS.n5736 VSS.n5709 0.374889
R9379 VSS.n5810 VSS.n5451 0.372135
R9380 VSS.n4898 VSS.n4897 0.371392
R9381 VSS.n5925 VSS.n5924 0.371022
R9382 VSS.n5922 VSS.n5921 0.370645
R9383 VSS.n4901 VSS.n4900 0.370645
R9384 VSS.n5706 VSS.n5704 0.358977
R9385 VSS.n5070 VSS.n5068 0.358977
R9386 VSS.n5078 VSS.n4946 0.356537
R9387 VSS.n4931 VSS.n4930 0.356409
R9388 VSS.n5788 VSS.n5707 0.354994
R9389 VSS.n4279 VSS.n4278 0.354579
R9390 VSS.n1680 VSS.n1677 0.354579
R9391 VSS.n5259 VSS.n5239 0.350926
R9392 VSS.n5712 VSS.n5710 0.347591
R9393 VSS.n5264 VSS.n5233 0.342028
R9394 VSS.n4929 VSS.n4928 0.341179
R9395 VSS.n5450 VSS.n5449 0.340476
R9396 VSS.n6250 VSS.n5948 0.331895
R9397 VSS.n6235 VSS.n6234 0.331895
R9398 VSS.n7193 VSS.t831 0.330516
R9399 VSS.n4369 VSS.n4366 0.327038
R9400 VSS.n6041 VSS.n6040 0.326081
R9401 VSS.n5760 VSS.n5708 0.321363
R9402 VSS.n5089 VSS.n4936 0.320022
R9403 VSS.n5448 VSS.n5447 0.31827
R9404 VSS.n5109 VSS.n23 0.313628
R9405 VSS VSS.n3027 0.307487
R9406 VSS.n219 VSS.n218 0.302495
R9407 VSS.n6264 VSS.n5890 0.301198
R9408 VSS.n4217 VSS.t467 0.301111
R9409 VSS.n1736 VSS.t358 0.301111
R9410 VSS.n1252 VSS.n1251 0.3005
R9411 VSS.n5636 VSS.n5455 0.292445
R9412 VSS.n5216 VSS.n5162 0.290903
R9413 VSS.n5646 VSS.n5454 0.289506
R9414 VSS.n5629 VSS.n5573 0.288772
R9415 VSS.n5205 VSS.n5163 0.287963
R9416 VSS.n7847 VSS.n5161 0.287229
R9417 VSS.n5614 VSS.n5613 0.285098
R9418 VSS.n5621 VSS.n5612 0.285098
R9419 VSS.n7867 VSS.n5159 0.283556
R9420 VSS.n7858 VSS.n5160 0.283556
R9421 VSS.n4663 VSS 0.281962
R9422 VSS.n4341 VSS.n4340 0.281213
R9423 VSS.n6581 VSS.n6580 0.280325
R9424 VSS.n5868 VSS.n5419 0.2753
R9425 VSS.n4130 VSS.n4129 0.274556
R9426 VSS.n4027 VSS.n4026 0.274296
R9427 VSS.n5438 VSS.n5437 0.2729
R9428 VSS.n5033 VSS.n4959 0.272046
R9429 VSS.n7360 VSS.n7304 0.271584
R9430 VSS.n5833 VSS.n5832 0.27149
R9431 VSS.n7427 VSS.n6329 0.270078
R9432 VSS.n5870 VSS.n5868 0.269479
R9433 VSS.n4979 VSS.n4978 0.269479
R9434 VSS.n4024 VSS.n4023 0.266088
R9435 VSS.n4907 VSS.n4893 0.254764
R9436 VSS.n4131 VSS.n4130 0.253311
R9437 VSS.n7422 VSS.n7421 0.25175
R9438 VSS.n5438 VSS.n5436 0.250935
R9439 VSS.n5419 VSS.n5418 0.250935
R9440 VSS.n4973 VSS.n4972 0.250935
R9441 VSS.n5013 VSS.n5012 0.250935
R9442 VSS.n5792 VSS.n5791 0.2505
R9443 VSS.n5073 VSS.n5072 0.2505
R9444 VSS.n7422 VSS.n6585 0.250143
R9445 VSS.n4906 VSS.n4905 0.24562
R9446 VSS.n5745 VSS.n5742 0.244911
R9447 VSS.n758 VSS 0.243106
R9448 VSS VSS.n6415 0.243106
R9449 VSS VSS.n7178 0.243106
R9450 VSS VSS.n947 0.243106
R9451 VSS.n7607 VSS 0.242302
R9452 VSS.n6805 VSS 0.242302
R9453 VSS.n6975 VSS.n6973 0.241879
R9454 VSS.n5931 VSS.n5930 0.241152
R9455 VSS.n5745 VSS.n5744 0.239887
R9456 VSS.n4754 VSS.n4745 0.235283
R9457 VSS.n6582 VSS.n6377 0.230988
R9458 VSS.n6581 VSS.n6386 0.230988
R9459 VSS.n4640 VSS.n4608 0.224214
R9460 VSS.n1735 VSS.n1733 0.220012
R9461 VSS.n1751 VSS.n1749 0.220012
R9462 VSS VSS.n1724 0.220012
R9463 VSS.n1716 VSS.n1715 0.220012
R9464 VSS.n4289 VSS.n4287 0.220012
R9465 VSS.n4294 VSS.n4292 0.220012
R9466 VSS.n4296 VSS.n4294 0.220012
R9467 VSS.n4298 VSS.n4296 0.220012
R9468 VSS.n4300 VSS.n4298 0.220012
R9469 VSS.n4305 VSS.n4303 0.220012
R9470 VSS VSS.n4305 0.220012
R9471 VSS.n4308 VSS 0.220012
R9472 VSS.n4313 VSS.n4311 0.220012
R9473 VSS.n1691 VSS.n1689 0.216354
R9474 VSS.n4303 VSS.n4301 0.216354
R9475 VSS.n5033 VSS.n5032 0.2141
R9476 VSS.n4907 VSS.n4906 0.21339
R9477 VSS.n5778 VSS.n5767 0.213053
R9478 VSS.n5755 VSS.n5749 0.213053
R9479 VSS.n5748 VSS.n5740 0.213053
R9480 VSS.n7148 VSS.n7147 0.21214
R9481 VSS.n5752 VSS.n5751 0.211098
R9482 VSS.n4978 VSS.n4975 0.207059
R9483 VSS.n7303 VSS.n7302 0.205724
R9484 VSS.n4519 VSS.n714 0.205426
R9485 VSS.n5870 VSS.n5869 0.205144
R9486 VSS.n5538 VSS.n5537 0.205045
R9487 VSS.n1752 VSS.n1751 0.204646
R9488 VSS.n1747 VSS.n1735 0.20172
R9489 VSS.n4290 VSS.n4289 0.20172
R9490 VSS.n4129 VSS.n4128 0.201552
R9491 VSS.n1723 VSS.n1716 0.200988
R9492 VSS.n4311 VSS.n4309 0.200988
R9493 VSS.n4221 VSS.n4219 0.200065
R9494 VSS.n4223 VSS.n4221 0.200065
R9495 VSS.n4225 VSS.n4223 0.200065
R9496 VSS.n4227 VSS.n4225 0.200065
R9497 VSS.n4229 VSS.n4227 0.200065
R9498 VSS.n4231 VSS.n4229 0.200065
R9499 VSS.n4233 VSS.n4231 0.200065
R9500 VSS.n4284 VSS.n4233 0.200065
R9501 VSS.n4284 VSS.n4283 0.200065
R9502 VSS.n4283 VSS.n4282 0.200065
R9503 VSS.n1740 VSS.n1738 0.200065
R9504 VSS.n1746 VSS.n1740 0.200065
R9505 VSS.n1746 VSS.n1745 0.200065
R9506 VSS.n1745 VSS.n1744 0.200065
R9507 VSS.n1636 VSS.n1634 0.200065
R9508 VSS.n1638 VSS.n1636 0.200065
R9509 VSS.n1686 VSS.n1638 0.200065
R9510 VSS.n1686 VSS.n1684 0.200065
R9511 VSS.n1684 VSS.n1683 0.200065
R9512 VSS.n6602 VSS.n6600 0.200065
R9513 VSS.n6609 VSS.n6608 0.200065
R9514 VSS.n4318 VSS.n4316 0.20001
R9515 VSS.n4905 VSS.n4904 0.199702
R9516 VSS.n7148 VSS.n7144 0.198571
R9517 VSS.n137 VSS.n136 0.1985
R9518 VSS.n5541 VSS.n5538 0.196574
R9519 VSS.n5775 VSS.n5774 0.196132
R9520 VSS.n4439 VSS.n4420 0.193921
R9521 VSS.n4453 VSS.n1607 0.193087
R9522 VSS.n6715 VSS.n6711 0.188841
R9523 VSS.n227 VSS.n226 0.188079
R9524 VSS.n860 VSS.n857 0.188
R9525 VSS.n7072 VSS.n7069 0.188
R9526 VSS.n6967 VSS.n6964 0.188
R9527 VSS.n1259 VSS.n1256 0.188
R9528 VSS.n5437 VSS.n5419 0.1865
R9529 VSS.n5014 VSS.n5013 0.1865
R9530 VSS.n4280 VSS.n4279 0.185391
R9531 VSS.n1681 VSS.n1680 0.185391
R9532 VSS.n145 VSS.n144 0.185092
R9533 VSS.n5439 VSS.n5438 0.1805
R9534 VSS.n5032 VSS.n4973 0.1805
R9535 VSS.n4128 VSS.n1755 0.176444
R9536 VSS.n4129 VSS.n1727 0.176444
R9537 VSS.n4130 VSS.n1632 0.176444
R9538 VSS.n4131 VSS.n1630 0.176444
R9539 VSS.n1133 VSS.n1132 0.17565
R9540 VSS.n4314 VSS.n4313 0.174646
R9541 VSS.n5134 VSS.n5131 0.174181
R9542 VSS.n6155 VSS.n6152 0.17414
R9543 VSS.n4776 VSS.n4775 0.174137
R9544 VSS.n5931 VSS.n5929 0.172819
R9545 VSS.n6460 VSS.n6434 0.169688
R9546 VSS.n4509 VSS.n4508 0.169688
R9547 VSS.n1000 VSS.n987 0.169688
R9548 VSS.n4699 VSS.n4698 0.164562
R9549 VSS.n4021 VSS.n4020 0.163308
R9550 VSS.n5451 VSS.n5450 0.163136
R9551 VSS.n4928 VSS.n4927 0.162433
R9552 VSS.n4594 VSS.n4592 0.161214
R9553 VSS.n760 VSS.n758 0.161214
R9554 VSS.n6415 VSS.n6414 0.161214
R9555 VSS.n6434 VSS.n6432 0.161214
R9556 VSS.n7232 VSS.n7231 0.161214
R9557 VSS.n7178 VSS.n7177 0.161214
R9558 VSS.n5350 VSS.n5348 0.161214
R9559 VSS.n7608 VSS.n7607 0.161214
R9560 VSS.n6684 VSS.n6682 0.161214
R9561 VSS.n6806 VSS.n6805 0.161214
R9562 VSS.n4510 VSS.n4509 0.161214
R9563 VSS.n4523 VSS.n4521 0.161214
R9564 VSS.n947 VSS.n946 0.161214
R9565 VSS.n1001 VSS.n1000 0.161214
R9566 VSS.n311 VSS.n307 0.160198
R9567 VSS.n4780 VSS.n4779 0.157329
R9568 VSS.n5936 VSS.n5934 0.15648
R9569 VSS VSS.n4594 0.155589
R9570 VSS.n5915 VSS.n5913 0.155512
R9571 VSS.n4764 VSS.n4761 0.153637
R9572 VSS.n5449 VSS.n5448 0.153513
R9573 VSS.n4908 VSS.n4907 0.152808
R9574 VSS.n1373 VSS.n1370 0.15275
R9575 VSS.n6831 VSS.n6828 0.15275
R9576 VSS.n6574 VSS.n6572 0.15275
R9577 VSS.n7636 VSS.n7633 0.15275
R9578 VSS.n1090 VSS.n1087 0.15275
R9579 VSS.n4930 VSS.n4929 0.152738
R9580 VSS.n5124 VSS.n5122 0.152674
R9581 VSS.n6490 VSS.n6489 0.151571
R9582 VSS.n7234 VSS.n7228 0.151571
R9583 VSS.n7613 VSS.n7610 0.151571
R9584 VSS.n6635 VSS.n6633 0.151571
R9585 VSS.n4480 VSS.n4479 0.151571
R9586 VSS.n4518 VSS.n4516 0.151571
R9587 VSS.n1004 VSS.n998 0.151571
R9588 VSS.n767 VSS.n766 0.150768
R9589 VSS.n6410 VSS.n6409 0.150768
R9590 VSS.n7175 VSS.n7174 0.150768
R9591 VSS.n6949 VSS.n6944 0.150768
R9592 VSS.n6743 VSS.n6742 0.150768
R9593 VSS.n942 VSS.n941 0.150768
R9594 VSS.n5661 VSS.n5660 0.150235
R9595 VSS.n5202 VSS.n5199 0.150235
R9596 VSS.n6122 VSS.n6119 0.148852
R9597 VSS.n6125 VSS.n6122 0.148852
R9598 VSS.n6128 VSS.n6125 0.148852
R9599 VSS.n6131 VSS.n6128 0.148852
R9600 VSS.n6134 VSS.n6131 0.148852
R9601 VSS.n6137 VSS.n6134 0.148852
R9602 VSS.n6140 VSS.n6137 0.148852
R9603 VSS.n6143 VSS.n6140 0.148852
R9604 VSS.n6146 VSS.n6143 0.148852
R9605 VSS.n6149 VSS.n6146 0.148852
R9606 VSS.n5680 VSS.n5677 0.148852
R9607 VSS.n5683 VSS.n5680 0.148852
R9608 VSS.n5686 VSS.n5683 0.148852
R9609 VSS.n5689 VSS.n5686 0.148852
R9610 VSS.n5692 VSS.n5689 0.148852
R9611 VSS.n5695 VSS.n5692 0.148852
R9612 VSS.n5698 VSS.n5695 0.148852
R9613 VSS.n5701 VSS.n5698 0.148852
R9614 VSS.n5704 VSS.n5701 0.148852
R9615 VSS.n5068 VSS.n5065 0.148852
R9616 VSS.n5065 VSS.n5062 0.148852
R9617 VSS.n5169 VSS.n5166 0.148852
R9618 VSS.n5172 VSS.n5169 0.148852
R9619 VSS.n5175 VSS.n5172 0.148852
R9620 VSS.n5178 VSS.n5175 0.148852
R9621 VSS.n5181 VSS.n5178 0.148852
R9622 VSS.n5184 VSS.n5181 0.148852
R9623 VSS.n5140 VSS.n5137 0.148852
R9624 VSS.n5143 VSS.n5140 0.148852
R9625 VSS.n5146 VSS.n5143 0.148852
R9626 VSS.n5149 VSS.n5146 0.148852
R9627 VSS.n5152 VSS.n5149 0.148852
R9628 VSS.n5155 VSS.n5152 0.148852
R9629 VSS.n5158 VSS.n5155 0.148852
R9630 VSS.n7884 VSS.n5158 0.148852
R9631 VSS.n7884 VSS.n7883 0.148852
R9632 VSS.n7883 VSS.n7880 0.148852
R9633 VSS.n4508 VSS.n725 0.148402
R9634 VSS.n6460 VSS.n6459 0.148402
R9635 VSS.n7081 VSS.n7073 0.148402
R9636 VSS.n7576 VSS.n7573 0.148402
R9637 VSS.n6773 VSS.n6770 0.148402
R9638 VSS.n987 VSS.n986 0.148402
R9639 VSS.n5847 VSS.n5844 0.147239
R9640 VSS.n5850 VSS.n5847 0.147239
R9641 VSS.n5816 VSS.n5813 0.147239
R9642 VSS.n5394 VSS.n5391 0.147239
R9643 VSS.n5860 VSS.n5857 0.147239
R9644 VSS.n5863 VSS.n5860 0.147239
R9645 VSS.n5888 VSS.n5886 0.147239
R9646 VSS.n5882 VSS.n5880 0.147239
R9647 VSS.n4769 VSS.n4767 0.147239
R9648 VSS.n5043 VSS.n5040 0.147239
R9649 VSS.n5024 VSS.n5021 0.147239
R9650 VSS.n5027 VSS.n5024 0.147239
R9651 VSS.n4995 VSS.n4992 0.147239
R9652 VSS.n4998 VSS.n4995 0.147239
R9653 VSS.n45 VSS.n41 0.147239
R9654 VSS.n4988 VSS.n4985 0.147239
R9655 VSS.n4796 VSS.n4793 0.147239
R9656 VSS.n4793 VSS.n4791 0.147239
R9657 VSS.n3028 VSS 0.145448
R9658 VSS.n6227 VSS.n6224 0.144304
R9659 VSS.n4802 VSS.n4799 0.144304
R9660 VSS.n7626 VSS.n7622 0.143986
R9661 VSS.n6818 VSS.n6620 0.143986
R9662 VSS.n5936 VSS.n5918 0.142348
R9663 VSS.n4783 VSS.n4782 0.142348
R9664 VSS.n4782 VSS.n4780 0.14137
R9665 VSS.n6152 VSS.n6149 0.139951
R9666 VSS.n5137 VSS.n5134 0.139951
R9667 VSS.n1382 VSS.n779 0.139082
R9668 VSS.n6563 VSS.n6393 0.139082
R9669 VSS.n7163 VSS.n7162 0.139082
R9670 VSS.n1076 VSS.n925 0.139082
R9671 VSS.n4919 VSS.n4918 0.138862
R9672 VSS.n4754 VSS.n4753 0.136472
R9673 VSS.n5910 VSS.n5909 0.136463
R9674 VSS.n7336 VSS.n7332 0.13325
R9675 VSS.n187 VSS.n186 0.132286
R9676 VSS.n681 VSS.n598 0.132194
R9677 VSS.n4249 VSS.n4248 0.132032
R9678 VSS.n1653 VSS.n1652 0.132032
R9679 VSS.n39 VSS.n33 0.131851
R9680 VSS.n6981 VSS.n6980 0.131118
R9681 VSS.n5050 VSS.n5047 0.130588
R9682 VSS.n51 VSS.n50 0.130302
R9683 VSS.n7490 VSS.n7486 0.13025
R9684 VSS.n5809 VSS.n5806 0.130084
R9685 VSS.n5878 VSS.n5877 0.129374
R9686 VSS.n7262 VSS.n7260 0.12841
R9687 VSS.n1458 VSS.n1455 0.12841
R9688 VSS.n7671 VSS.n7667 0.128
R9689 VSS.n6869 VSS.n6866 0.128
R9690 VSS.n1342 VSS.n1339 0.128
R9691 VSS.n4989 VSS.n4988 0.127674
R9692 VSS.n819 VSS.n817 0.12766
R9693 VSS.n6476 VSS.n6473 0.12766
R9694 VSS.n6729 VSS.n6726 0.12766
R9695 VSS.n7531 VSS.n7527 0.12766
R9696 VSS.n7423 VSS.n7422 0.12665
R9697 VSS.n5876 VSS.n5875 0.125349
R9698 VSS.n4560 VSS.n4559 0.12483
R9699 VSS.n7424 VSS.n7423 0.124735
R9700 VSS.n49 VSS.n48 0.124421
R9701 VSS.n5911 VSS.n5910 0.123458
R9702 VSS.n6329 VSS.n6328 0.123275
R9703 VSS.n4799 VSS.n4796 0.122783
R9704 VSS.n5938 VSS.n5937 0.122669
R9705 VSS.n4755 VSS.n4754 0.122609
R9706 VSS.n1594 VSS.n1593 0.1225
R9707 VSS.n5932 VSS.n5931 0.12249
R9708 VSS.n5873 VSS.n5872 0.121959
R9709 VSS.n5913 VSS.n5912 0.121915
R9710 VSS.n5934 VSS.n5933 0.121915
R9711 VSS.n4757 VSS.n4756 0.121915
R9712 VSS.n4779 VSS.n4778 0.121915
R9713 VSS.n4759 VSS.n4758 0.121893
R9714 VSS.n5875 VSS.n5874 0.121804
R9715 VSS.n48 VSS.n47 0.121804
R9716 VSS.n4777 VSS.n4776 0.121641
R9717 VSS.n5401 VSS.n5397 0.120826
R9718 VSS.n5028 VSS.n4949 0.120826
R9719 VSS.n5660 VSS.n5649 0.119969
R9720 VSS.n5645 VSS.n5642 0.119969
R9721 VSS.n5642 VSS.n5639 0.119969
R9722 VSS.n5625 VSS.n5623 0.119969
R9723 VSS.n5620 VSS.n5618 0.119969
R9724 VSS.n5618 VSS.n5616 0.119969
R9725 VSS.n6114 VSS.n6111 0.119969
R9726 VSS.n6116 VSS.n6114 0.119969
R9727 VSS.n5731 VSS.n5729 0.119969
R9728 VSS.n5793 VSS.n5790 0.119969
R9729 VSS.n5726 VSS.n5724 0.119969
R9730 VSS.n5077 VSS.n5074 0.119969
R9731 VSS.n5116 VSS.n5114 0.119969
R9732 VSS.n5114 VSS.n5111 0.119969
R9733 VSS.n5107 VSS.n5104 0.119969
R9734 VSS.n7877 VSS.n7873 0.119969
R9735 VSS.n7873 VSS.n7871 0.119969
R9736 VSS.n7866 VSS.n7863 0.119969
R9737 VSS.n7863 VSS.n7860 0.119969
R9738 VSS.n7857 VSS.n7854 0.119969
R9739 VSS.n7854 VSS.n7850 0.119969
R9740 VSS.n5221 VSS.n5218 0.119969
R9741 VSS.n5215 VSS.n5212 0.119969
R9742 VSS.n5212 VSS.n5208 0.119969
R9743 VSS.n5204 VSS.n5202 0.119969
R9744 VSS.n5841 VSS.n5840 0.119848
R9745 VSS.n38 VSS.n35 0.119848
R9746 VSS.n4554 VSS.n4553 0.119263
R9747 VSS.n695 VSS.n694 0.119263
R9748 VSS.n5128 VSS.n5125 0.119173
R9749 VSS.n6201 VSS.n6198 0.118921
R9750 VSS.n6204 VSS.n6201 0.118921
R9751 VSS.n6207 VSS.n6204 0.118921
R9752 VSS.n6210 VSS.n6207 0.118921
R9753 VSS.n6188 VSS.n6185 0.118921
R9754 VSS.n6191 VSS.n6188 0.118921
R9755 VSS.n6181 VSS.n6178 0.118921
R9756 VSS.n4815 VSS.n4812 0.118921
R9757 VSS.n4818 VSS.n4815 0.118921
R9758 VSS.n4821 VSS.n4818 0.118921
R9759 VSS.n4824 VSS.n4821 0.118921
R9760 VSS.n4827 VSS.n4824 0.118921
R9761 VSS.n4830 VSS.n4827 0.118921
R9762 VSS.n4833 VSS.n4830 0.118921
R9763 VSS.n4836 VSS.n4833 0.118921
R9764 VSS.n4843 VSS.n4840 0.118921
R9765 VSS.n4846 VSS.n4843 0.118921
R9766 VSS.n4849 VSS.n4846 0.118921
R9767 VSS.n4852 VSS.n4849 0.118921
R9768 VSS.n4855 VSS.n4852 0.118921
R9769 VSS.n5877 VSS.n5876 0.118335
R9770 VSS.n50 VSS.n49 0.118335
R9771 VSS.n7425 VSS.n7424 0.118151
R9772 VSS.n5131 VSS.n5128 0.116783
R9773 VSS.n6214 VSS.n6211 0.116553
R9774 VSS.n6224 VSS.n6221 0.115403
R9775 VSS.n6158 VSS.n6157 0.115328
R9776 VSS.n4805 VSS.n4802 0.115214
R9777 VSS.n1420 VSS.n1418 0.113945
R9778 VSS.n1418 VSS.n1416 0.113945
R9779 VSS.n1412 VSS.n1410 0.113945
R9780 VSS.n1410 VSS.n1406 0.113945
R9781 VSS.n1406 VSS.n1404 0.113945
R9782 VSS.n1404 VSS.n1400 0.113945
R9783 VSS.n1400 VSS.n1396 0.113945
R9784 VSS.n1396 VSS.n1393 0.113945
R9785 VSS.n1388 VSS.n1387 0.113945
R9786 VSS.n1387 VSS.n1384 0.113945
R9787 VSS.n6479 VSS.n6476 0.113945
R9788 VSS.n6482 VSS.n6479 0.113945
R9789 VSS.n6497 VSS.n6482 0.113945
R9790 VSS.n6500 VSS.n6497 0.113945
R9791 VSS.n6504 VSS.n6500 0.113945
R9792 VSS.n6511 VSS.n6508 0.113945
R9793 VSS.n6514 VSS.n6511 0.113945
R9794 VSS.n6521 VSS.n6518 0.113945
R9795 VSS.n6524 VSS.n6521 0.113945
R9796 VSS.n6527 VSS.n6524 0.113945
R9797 VSS.n6530 VSS.n6527 0.113945
R9798 VSS.n6537 VSS.n6534 0.113945
R9799 VSS.n6540 VSS.n6537 0.113945
R9800 VSS.n6543 VSS.n6540 0.113945
R9801 VSS.n6546 VSS.n6543 0.113945
R9802 VSS.n6549 VSS.n6546 0.113945
R9803 VSS.n6552 VSS.n6549 0.113945
R9804 VSS.n6559 VSS.n6556 0.113945
R9805 VSS.n6562 VSS.n6559 0.113945
R9806 VSS.n7260 VSS.n7257 0.113945
R9807 VSS.n7257 VSS.n7254 0.113945
R9808 VSS.n7254 VSS.n7250 0.113945
R9809 VSS.n7250 VSS.n7241 0.113945
R9810 VSS.n7241 VSS.n7238 0.113945
R9811 VSS.n7222 VSS.n7219 0.113945
R9812 VSS.n7219 VSS.n7216 0.113945
R9813 VSS.n7212 VSS.n7209 0.113945
R9814 VSS.n7209 VSS.n7206 0.113945
R9815 VSS.n7206 VSS.n7203 0.113945
R9816 VSS.n7203 VSS.n7200 0.113945
R9817 VSS.n7103 VSS.n7100 0.113945
R9818 VSS.n7106 VSS.n7103 0.113945
R9819 VSS.n7109 VSS.n7106 0.113945
R9820 VSS.n7112 VSS.n7109 0.113945
R9821 VSS.n7115 VSS.n7112 0.113945
R9822 VSS.n7118 VSS.n7115 0.113945
R9823 VSS.n7134 VSS.n7131 0.113945
R9824 VSS.n7137 VSS.n7134 0.113945
R9825 VSS.n7157 VSS.n7154 0.113945
R9826 VSS.n7554 VSS.n7551 0.113945
R9827 VSS.n5313 VSS.n5310 0.113945
R9828 VSS.n5325 VSS.n5322 0.113945
R9829 VSS.n5328 VSS.n5325 0.113945
R9830 VSS.n5333 VSS.n5328 0.113945
R9831 VSS.n5336 VSS.n5333 0.113945
R9832 VSS.n5339 VSS.n5336 0.113945
R9833 VSS.n5342 VSS.n5339 0.113945
R9834 VSS.n7564 VSS.n7561 0.113945
R9835 VSS.n6817 VSS.n6814 0.113945
R9836 VSS.n6814 VSS.n6811 0.113945
R9837 VSS.n6646 VSS.n6643 0.113945
R9838 VSS.n6649 VSS.n6646 0.113945
R9839 VSS.n6652 VSS.n6649 0.113945
R9840 VSS.n6655 VSS.n6652 0.113945
R9841 VSS.n6658 VSS.n6655 0.113945
R9842 VSS.n6661 VSS.n6658 0.113945
R9843 VSS.n6671 VSS.n6668 0.113945
R9844 VSS.n6674 VSS.n6671 0.113945
R9845 VSS.n6677 VSS.n6674 0.113945
R9846 VSS.n6680 VSS.n6677 0.113945
R9847 VSS.n6768 VSS.n6765 0.113945
R9848 VSS.n6765 VSS.n6762 0.113945
R9849 VSS.n6758 VSS.n6755 0.113945
R9850 VSS.n6755 VSS.n6752 0.113945
R9851 VSS.n6752 VSS.n6736 0.113945
R9852 VSS.n6736 VSS.n6732 0.113945
R9853 VSS.n6732 VSS.n6729 0.113945
R9854 VSS.n7539 VSS.n7536 0.113945
R9855 VSS.n7536 VSS.n7533 0.113945
R9856 VSS.n7533 VSS.n7531 0.113945
R9857 VSS.n1461 VSS.n1458 0.113945
R9858 VSS.n1464 VSS.n1461 0.113945
R9859 VSS.n1468 VSS.n1464 0.113945
R9860 VSS.n1471 VSS.n1468 0.113945
R9861 VSS.n1475 VSS.n1471 0.113945
R9862 VSS.n4488 VSS.n4485 0.113945
R9863 VSS.n817 VSS.n815 0.113945
R9864 VSS.n1011 VSS.n1008 0.113945
R9865 VSS.n1014 VSS.n1011 0.113945
R9866 VSS.n1017 VSS.n1014 0.113945
R9867 VSS.n1024 VSS.n1021 0.113945
R9868 VSS.n1027 VSS.n1024 0.113945
R9869 VSS.n1034 VSS.n1031 0.113945
R9870 VSS.n1037 VSS.n1034 0.113945
R9871 VSS.n1040 VSS.n1037 0.113945
R9872 VSS.n1043 VSS.n1040 0.113945
R9873 VSS.n1050 VSS.n1047 0.113945
R9874 VSS.n1053 VSS.n1050 0.113945
R9875 VSS.n1056 VSS.n1053 0.113945
R9876 VSS.n1059 VSS.n1056 0.113945
R9877 VSS.n1062 VSS.n1059 0.113945
R9878 VSS.n1065 VSS.n1062 0.113945
R9879 VSS.n1072 VSS.n1069 0.113945
R9880 VSS.n1075 VSS.n1072 0.113945
R9881 VSS.n1381 VSS.n1377 0.113933
R9882 VSS.n6825 VSS.n6821 0.113933
R9883 VSS.n6569 VSS.n6566 0.113933
R9884 VSS.n7632 VSS.n7629 0.113933
R9885 VSS.n1082 VSS.n1079 0.113933
R9886 VSS.n1624 VSS.n1623 0.113915
R9887 VSS.n6157 VSS.n6155 0.113776
R9888 VSS.n5727 VSS.n5726 0.113597
R9889 VSS.n821 VSS.n819 0.113
R9890 VSS.n824 VSS.n821 0.113
R9891 VSS.n827 VSS.n824 0.113
R9892 VSS.n829 VSS.n827 0.113
R9893 VSS.n836 VSS.n829 0.113
R9894 VSS.n839 VSS.n836 0.113
R9895 VSS.n842 VSS.n839 0.113
R9896 VSS.n845 VSS.n842 0.113
R9897 VSS.n848 VSS.n845 0.113
R9898 VSS.n851 VSS.n848 0.113
R9899 VSS.n854 VSS.n851 0.113
R9900 VSS.n857 VSS.n854 0.113
R9901 VSS.n863 VSS.n860 0.113
R9902 VSS.n866 VSS.n863 0.113
R9903 VSS.n869 VSS.n866 0.113
R9904 VSS.n872 VSS.n869 0.113
R9905 VSS.n875 VSS.n872 0.113
R9906 VSS.n878 VSS.n875 0.113
R9907 VSS.n881 VSS.n878 0.113
R9908 VSS.n884 VSS.n881 0.113
R9909 VSS.n887 VSS.n884 0.113
R9910 VSS.n890 VSS.n887 0.113
R9911 VSS.n893 VSS.n890 0.113
R9912 VSS.n896 VSS.n893 0.113
R9913 VSS.n899 VSS.n896 0.113
R9914 VSS.n902 VSS.n899 0.113
R9915 VSS.n905 VSS.n902 0.113
R9916 VSS.n908 VSS.n905 0.113
R9917 VSS.n911 VSS.n908 0.113
R9918 VSS.n914 VSS.n911 0.113
R9919 VSS.n917 VSS.n914 0.113
R9920 VSS.n920 VSS.n917 0.113
R9921 VSS.n1370 VSS.n1368 0.113
R9922 VSS.n1377 VSS.n1373 0.113
R9923 VSS.n6828 VSS.n6825 0.113
R9924 VSS.n6572 VSS.n6569 0.113
R9925 VSS.n6577 VSS.n6574 0.113
R9926 VSS.n6579 VSS.n6577 0.113
R9927 VSS.n6473 VSS.n6469 0.113
R9928 VSS.n6469 VSS.n6467 0.113
R9929 VSS.n6467 VSS.n6464 0.113
R9930 VSS.n7310 VSS.n7306 0.113
R9931 VSS.n7313 VSS.n7310 0.113
R9932 VSS.n7316 VSS.n7313 0.113
R9933 VSS.n7319 VSS.n7316 0.113
R9934 VSS.n7323 VSS.n7319 0.113
R9935 VSS.n7326 VSS.n7323 0.113
R9936 VSS.n7328 VSS.n7326 0.113
R9937 VSS.n7332 VSS.n7328 0.113
R9938 VSS.n7342 VSS.n7339 0.113
R9939 VSS.n7352 VSS.n7349 0.113
R9940 VSS.n7359 VSS.n7356 0.113
R9941 VSS.n7366 VSS.n7363 0.113
R9942 VSS.n7369 VSS.n7366 0.113
R9943 VSS.n7372 VSS.n7369 0.113
R9944 VSS.n7375 VSS.n7372 0.113
R9945 VSS.n7380 VSS.n7375 0.113
R9946 VSS.n7383 VSS.n7380 0.113
R9947 VSS.n7386 VSS.n7383 0.113
R9948 VSS.n7389 VSS.n7386 0.113
R9949 VSS.n7392 VSS.n7389 0.113
R9950 VSS.n7397 VSS.n7392 0.113
R9951 VSS.n7400 VSS.n7397 0.113
R9952 VSS.n7403 VSS.n7400 0.113
R9953 VSS.n7406 VSS.n7403 0.113
R9954 VSS.n7409 VSS.n7406 0.113
R9955 VSS.n7412 VSS.n7409 0.113
R9956 VSS.n7415 VSS.n7412 0.113
R9957 VSS.n7417 VSS.n7415 0.113
R9958 VSS.n7421 VSS.n7417 0.113
R9959 VSS.n6338 VSS.n6334 0.113
R9960 VSS.n6334 VSS.n6332 0.113
R9961 VSS.n6356 VSS.n6353 0.113
R9962 VSS.n6349 VSS.n6346 0.113
R9963 VSS.n7069 VSS.n7066 0.113
R9964 VSS.n7066 VSS.n7063 0.113
R9965 VSS.n7063 VSS.n7062 0.113
R9966 VSS.n7062 VSS.n7059 0.113
R9967 VSS.n7059 VSS.n7056 0.113
R9968 VSS.n7056 VSS.n7053 0.113
R9969 VSS.n7053 VSS.n7050 0.113
R9970 VSS.n7050 VSS.n7047 0.113
R9971 VSS.n7047 VSS.n7044 0.113
R9972 VSS.n7044 VSS.n7041 0.113
R9973 VSS.n7041 VSS.n7038 0.113
R9974 VSS.n7038 VSS.n7035 0.113
R9975 VSS.n7035 VSS.n7032 0.113
R9976 VSS.n7032 VSS.n7029 0.113
R9977 VSS.n7029 VSS.n7026 0.113
R9978 VSS.n7026 VSS.n7023 0.113
R9979 VSS.n7023 VSS.n7020 0.113
R9980 VSS.n7020 VSS.n7017 0.113
R9981 VSS.n7017 VSS.n7014 0.113
R9982 VSS.n7014 VSS.n7011 0.113
R9983 VSS.n7011 VSS.n7008 0.113
R9984 VSS.n7008 VSS.n7005 0.113
R9985 VSS.n7005 VSS.n7002 0.113
R9986 VSS.n7002 VSS.n6999 0.113
R9987 VSS.n6999 VSS.n6995 0.113
R9988 VSS.n6995 VSS.n6993 0.113
R9989 VSS.n7294 VSS.n7072 0.113
R9990 VSS.n7294 VSS.n7293 0.113
R9991 VSS.n7293 VSS.n7290 0.113
R9992 VSS.n7290 VSS.n7287 0.113
R9993 VSS.n7287 VSS.n7284 0.113
R9994 VSS.n7284 VSS.n7281 0.113
R9995 VSS.n7281 VSS.n7278 0.113
R9996 VSS.n7278 VSS.n7274 0.113
R9997 VSS.n7274 VSS.n7272 0.113
R9998 VSS.n7272 VSS.n7267 0.113
R9999 VSS.n7267 VSS.n7265 0.113
R10000 VSS.n7265 VSS.n7262 0.113
R10001 VSS.n6919 VSS.n6916 0.113
R10002 VSS.n5364 VSS.n5362 0.113
R10003 VSS.n7674 VSS.n7671 0.113
R10004 VSS.n7677 VSS.n7674 0.113
R10005 VSS.n7680 VSS.n7677 0.113
R10006 VSS.n7683 VSS.n7680 0.113
R10007 VSS.n7686 VSS.n7683 0.113
R10008 VSS.n7689 VSS.n7686 0.113
R10009 VSS.n7692 VSS.n7689 0.113
R10010 VSS.n7695 VSS.n7692 0.113
R10011 VSS.n7698 VSS.n7695 0.113
R10012 VSS.n7701 VSS.n7698 0.113
R10013 VSS.n7704 VSS.n7701 0.113
R10014 VSS.n7707 VSS.n7704 0.113
R10015 VSS.n7713 VSS.n7707 0.113
R10016 VSS.n7716 VSS.n7713 0.113
R10017 VSS.n7719 VSS.n7716 0.113
R10018 VSS.n7722 VSS.n7719 0.113
R10019 VSS.n7725 VSS.n7722 0.113
R10020 VSS.n7727 VSS.n7725 0.113
R10021 VSS.n7638 VSS.n7636 0.113
R10022 VSS.n7641 VSS.n7638 0.113
R10023 VSS.n7643 VSS.n7641 0.113
R10024 VSS.n7646 VSS.n7643 0.113
R10025 VSS.n7648 VSS.n7646 0.113
R10026 VSS.n7651 VSS.n7648 0.113
R10027 VSS.n7653 VSS.n7651 0.113
R10028 VSS.n7656 VSS.n7653 0.113
R10029 VSS.n7658 VSS.n7656 0.113
R10030 VSS.n7661 VSS.n7658 0.113
R10031 VSS.n7663 VSS.n7661 0.113
R10032 VSS.n7667 VSS.n7663 0.113
R10033 VSS.n7633 VSS.n7632 0.113
R10034 VSS.n6872 VSS.n6869 0.113
R10035 VSS.n6875 VSS.n6872 0.113
R10036 VSS.n6878 VSS.n6875 0.113
R10037 VSS.n6881 VSS.n6878 0.113
R10038 VSS.n6884 VSS.n6881 0.113
R10039 VSS.n6887 VSS.n6884 0.113
R10040 VSS.n6890 VSS.n6887 0.113
R10041 VSS.n6893 VSS.n6890 0.113
R10042 VSS.n6896 VSS.n6893 0.113
R10043 VSS.n6900 VSS.n6896 0.113
R10044 VSS.n6903 VSS.n6900 0.113
R10045 VSS.n6906 VSS.n6903 0.113
R10046 VSS.n6909 VSS.n6906 0.113
R10047 VSS.n6912 VSS.n6909 0.113
R10048 VSS.n6833 VSS.n6831 0.113
R10049 VSS.n6837 VSS.n6833 0.113
R10050 VSS.n6840 VSS.n6837 0.113
R10051 VSS.n6842 VSS.n6840 0.113
R10052 VSS.n6846 VSS.n6842 0.113
R10053 VSS.n6849 VSS.n6846 0.113
R10054 VSS.n6852 VSS.n6849 0.113
R10055 VSS.n6855 VSS.n6852 0.113
R10056 VSS.n6857 VSS.n6855 0.113
R10057 VSS.n6860 VSS.n6857 0.113
R10058 VSS.n6862 VSS.n6860 0.113
R10059 VSS.n6866 VSS.n6862 0.113
R10060 VSS.n6726 VSS.n6723 0.113
R10061 VSS.n6723 VSS.n6721 0.113
R10062 VSS.n6721 VSS.n6708 0.113
R10063 VSS.n6708 VSS.n6705 0.113
R10064 VSS.n6705 VSS.n6703 0.113
R10065 VSS.n6703 VSS.n6699 0.113
R10066 VSS.n6699 VSS.n6694 0.113
R10067 VSS.n6694 VSS.n6691 0.113
R10068 VSS.n6691 VSS.n6688 0.113
R10069 VSS.n6688 VSS.n6615 0.113
R10070 VSS.n6968 VSS.n6615 0.113
R10071 VSS.n6968 VSS.n6967 0.113
R10072 VSS.n6958 VSS.n6955 0.113
R10073 VSS.n6962 VSS.n6958 0.113
R10074 VSS.n6964 VSS.n6962 0.113
R10075 VSS.n7527 VSS.n7524 0.113
R10076 VSS.n7524 VSS.n7520 0.113
R10077 VSS.n7520 VSS.n7517 0.113
R10078 VSS.n7517 VSS.n7514 0.113
R10079 VSS.n7514 VSS.n7511 0.113
R10080 VSS.n7511 VSS.n7508 0.113
R10081 VSS.n7508 VSS.n7505 0.113
R10082 VSS.n7505 VSS.n7502 0.113
R10083 VSS.n7502 VSS.n7499 0.113
R10084 VSS.n7499 VSS.n7496 0.113
R10085 VSS.n7496 VSS.n7493 0.113
R10086 VSS.n7493 VSS.n7490 0.113
R10087 VSS.n514 VSS.n512 0.113
R10088 VSS.n1344 VSS.n1342 0.113
R10089 VSS.n1347 VSS.n1344 0.113
R10090 VSS.n1349 VSS.n1347 0.113
R10091 VSS.n1352 VSS.n1349 0.113
R10092 VSS.n1354 VSS.n1352 0.113
R10093 VSS.n1357 VSS.n1354 0.113
R10094 VSS.n1359 VSS.n1357 0.113
R10095 VSS.n1362 VSS.n1359 0.113
R10096 VSS.n1364 VSS.n1362 0.113
R10097 VSS.n1263 VSS.n1259 0.113
R10098 VSS.n1266 VSS.n1263 0.113
R10099 VSS.n1269 VSS.n1266 0.113
R10100 VSS.n1272 VSS.n1269 0.113
R10101 VSS.n1275 VSS.n1272 0.113
R10102 VSS.n1278 VSS.n1275 0.113
R10103 VSS.n1281 VSS.n1278 0.113
R10104 VSS.n1284 VSS.n1281 0.113
R10105 VSS.n1288 VSS.n1284 0.113
R10106 VSS.n1291 VSS.n1288 0.113
R10107 VSS.n1294 VSS.n1291 0.113
R10108 VSS.n1297 VSS.n1294 0.113
R10109 VSS.n1300 VSS.n1297 0.113
R10110 VSS.n1303 VSS.n1300 0.113
R10111 VSS.n1306 VSS.n1303 0.113
R10112 VSS.n1309 VSS.n1306 0.113
R10113 VSS.n1313 VSS.n1309 0.113
R10114 VSS.n1316 VSS.n1313 0.113
R10115 VSS.n1319 VSS.n1316 0.113
R10116 VSS.n1322 VSS.n1319 0.113
R10117 VSS.n1325 VSS.n1322 0.113
R10118 VSS.n1328 VSS.n1325 0.113
R10119 VSS.n1331 VSS.n1328 0.113
R10120 VSS.n1334 VSS.n1331 0.113
R10121 VSS.n1336 VSS.n1334 0.113
R10122 VSS.n1339 VSS.n1336 0.113
R10123 VSS.n1425 VSS.n1422 0.113
R10124 VSS.n1428 VSS.n1425 0.113
R10125 VSS.n1431 VSS.n1428 0.113
R10126 VSS.n1434 VSS.n1431 0.113
R10127 VSS.n1437 VSS.n1434 0.113
R10128 VSS.n1440 VSS.n1437 0.113
R10129 VSS.n1443 VSS.n1440 0.113
R10130 VSS.n1446 VSS.n1443 0.113
R10131 VSS.n1449 VSS.n1446 0.113
R10132 VSS.n1453 VSS.n1449 0.113
R10133 VSS.n1455 VSS.n1453 0.113
R10134 VSS.n1087 VSS.n1082 0.113
R10135 VSS.n1092 VSS.n1090 0.113
R10136 VSS.n1096 VSS.n1092 0.113
R10137 VSS.n1099 VSS.n1096 0.113
R10138 VSS.n1101 VSS.n1099 0.113
R10139 VSS.n1106 VSS.n1101 0.113
R10140 VSS.n1109 VSS.n1106 0.113
R10141 VSS.n1112 VSS.n1109 0.113
R10142 VSS.n1115 VSS.n1112 0.113
R10143 VSS.n1118 VSS.n1115 0.113
R10144 VSS.n1121 VSS.n1118 0.113
R10145 VSS.n1124 VSS.n1121 0.113
R10146 VSS.n1126 VSS.n1124 0.113
R10147 VSS.n7573 VSS.n7572 0.112646
R10148 VSS.n1249 VSS.n1246 0.112367
R10149 VSS.n4783 VSS.n4757 0.111845
R10150 VSS.n7356 VSS.n7353 0.1115
R10151 VSS.n5940 VSS.n5939 0.111448
R10152 VSS.n4761 VSS.n4760 0.111448
R10153 VSS.n305 VSS.n301 0.111156
R10154 VSS.n307 VSS.n305 0.111156
R10155 VSS.n7304 VSS.n7303 0.111102
R10156 VSS.n301 VSS.n299 0.11043
R10157 VSS.n4459 VSS.n4456 0.110256
R10158 VSS.n4472 VSS.n4459 0.110256
R10159 VSS.n4472 VSS.n4471 0.110256
R10160 VSS.n4471 VSS.n4468 0.110256
R10161 VSS.n4468 VSS.n4465 0.110256
R10162 VSS.n4465 VSS.n4462 0.110256
R10163 VSS.n4155 VSS.n4152 0.110256
R10164 VSS.n4152 VSS.n4149 0.110256
R10165 VSS.n65 VSS.n62 0.110256
R10166 VSS.n62 VSS.n59 0.110256
R10167 VSS.n59 VSS.n56 0.110256
R10168 VSS.n555 VSS.n552 0.110256
R10169 VSS.n552 VSS.n549 0.110256
R10170 VSS.n549 VSS.n546 0.110256
R10171 VSS.n4145 VSS.n4141 0.110256
R10172 VSS.n98 VSS.n95 0.110256
R10173 VSS.n101 VSS.n98 0.110256
R10174 VSS.n104 VSS.n101 0.110256
R10175 VSS.n107 VSS.n104 0.110256
R10176 VSS.n110 VSS.n107 0.110256
R10177 VSS.n113 VSS.n110 0.110256
R10178 VSS.n116 VSS.n113 0.110256
R10179 VSS.n120 VSS.n116 0.110256
R10180 VSS.n123 VSS.n120 0.110256
R10181 VSS.n126 VSS.n123 0.110256
R10182 VSS.n129 VSS.n126 0.110256
R10183 VSS.n132 VSS.n129 0.110256
R10184 VSS.n135 VSS.n78 0.110256
R10185 VSS.n233 VSS.n230 0.110256
R10186 VSS.n236 VSS.n233 0.110256
R10187 VSS.n241 VSS.n236 0.110256
R10188 VSS.n244 VSS.n241 0.110256
R10189 VSS.n247 VSS.n244 0.110256
R10190 VSS.n250 VSS.n247 0.110256
R10191 VSS.n253 VSS.n250 0.110256
R10192 VSS.n256 VSS.n253 0.110256
R10193 VSS.n259 VSS.n256 0.110256
R10194 VSS.n262 VSS.n259 0.110256
R10195 VSS.n265 VSS.n262 0.110256
R10196 VSS.n268 VSS.n265 0.110256
R10197 VSS.n272 VSS.n268 0.110256
R10198 VSS.n275 VSS.n272 0.110256
R10199 VSS.n278 VSS.n275 0.110256
R10200 VSS.n287 VSS.n278 0.110256
R10201 VSS.n290 VSS.n287 0.110256
R10202 VSS.n293 VSS.n290 0.110256
R10203 VSS.n296 VSS.n293 0.110256
R10204 VSS.n299 VSS.n296 0.110256
R10205 VSS.n713 VSS.n711 0.110256
R10206 VSS.n711 VSS.n708 0.110256
R10207 VSS.n708 VSS.n706 0.110256
R10208 VSS.n706 VSS.n704 0.110256
R10209 VSS.n704 VSS.n702 0.110256
R10210 VSS.n702 VSS.n700 0.110256
R10211 VSS.n4615 VSS.n4612 0.110256
R10212 VSS.n4618 VSS.n4615 0.110256
R10213 VSS.n4620 VSS.n4618 0.110256
R10214 VSS.n4623 VSS.n4620 0.110256
R10215 VSS.n4625 VSS.n4623 0.110256
R10216 VSS.n4629 VSS.n4625 0.110256
R10217 VSS.n4632 VSS.n4629 0.110256
R10218 VSS.n4635 VSS.n4632 0.110256
R10219 VSS.n4639 VSS.n4635 0.110256
R10220 VSS.n4646 VSS.n4643 0.110256
R10221 VSS.n4649 VSS.n4646 0.110256
R10222 VSS.n4652 VSS.n4649 0.110256
R10223 VSS.n4655 VSS.n4652 0.110256
R10224 VSS.n4658 VSS.n4655 0.110256
R10225 VSS.n4668 VSS.n4666 0.110256
R10226 VSS.n4671 VSS.n4668 0.110256
R10227 VSS.n4674 VSS.n4671 0.110256
R10228 VSS.n4686 VSS.n4683 0.110256
R10229 VSS.n4683 VSS.n4680 0.110256
R10230 VSS.n4680 VSS.n4677 0.110256
R10231 VSS.n4435 VSS.n4432 0.110256
R10232 VSS.n4438 VSS.n4435 0.110256
R10233 VSS.n4446 VSS.n4442 0.110256
R10234 VSS.n4449 VSS.n4446 0.110256
R10235 VSS.n4452 VSS.n4449 0.110256
R10236 VSS.n4428 VSS.n4426 0.110256
R10237 VSS.n4365 VSS.n4363 0.110256
R10238 VSS.n4363 VSS.n4361 0.110256
R10239 VSS.n4361 VSS.n4354 0.110256
R10240 VSS.n4354 VSS.n4351 0.110256
R10241 VSS.n4195 VSS.n4192 0.110256
R10242 VSS.n4192 VSS.n4189 0.110256
R10243 VSS.n4189 VSS.n4186 0.110256
R10244 VSS.n4186 VSS.n4183 0.110256
R10245 VSS.n4183 VSS.n4180 0.110256
R10246 VSS.n4180 VSS.n4177 0.110256
R10247 VSS.n4177 VSS.n4174 0.110256
R10248 VSS.n4174 VSS.n4168 0.110256
R10249 VSS.n4168 VSS.n4165 0.110256
R10250 VSS.n4165 VSS.n4162 0.110256
R10251 VSS.n4162 VSS.n4159 0.110256
R10252 VSS.n5872 VSS.n5871 0.109357
R10253 VSS.n4977 VSS.n4976 0.109357
R10254 VSS VSS.n7797 0.109087
R10255 VSS.n1627 VSS.n1626 0.108793
R10256 VSS.n7551 VSS.n7548 0.108651
R10257 VSS.n5941 VSS.n5940 0.108345
R10258 VSS.n5912 VSS.n5911 0.10833
R10259 VSS.n5933 VSS.n5932 0.10833
R10260 VSS.n4756 VSS.n4755 0.10833
R10261 VSS.n4778 VSS.n4777 0.10833
R10262 VSS.n6164 VSS.n6161 0.108109
R10263 VSS.n4861 VSS.n4858 0.108109
R10264 VSS.n312 VSS.n311 0.108061
R10265 VSS.n4439 VSS.n4438 0.108061
R10266 VSS.n1416 VSS.n1413 0.107895
R10267 VSS.n6531 VSS.n6530 0.107895
R10268 VSS.n7200 VSS.n7074 0.107895
R10269 VSS.n7561 VSS.n5343 0.107895
R10270 VSS.n6668 VSS.n6662 0.107895
R10271 VSS.n1044 VSS.n1043 0.107895
R10272 VSS.n924 VSS.n921 0.10775
R10273 VSS.n4337 VSS.n4335 0.107643
R10274 VSS.n4339 VSS.n4337 0.107643
R10275 VSS.n5915 VSS.n5893 0.10713
R10276 VSS.n6195 VSS.n6194 0.107079
R10277 VSS.n140 VSS 0.107055
R10278 VSS.n1626 VSS.n1624 0.106598
R10279 VSS.n5631 VSS.n5629 0.106429
R10280 VSS.n7908 VSS 0.10626
R10281 VSS.n4687 VSS.n4686 0.105134
R10282 VSS.n6221 VSS.n6218 0.104711
R10283 VSS.n4808 VSS.n4805 0.104711
R10284 VSS.n5886 VSS.n5883 0.104196
R10285 VSS.n52 VSS.n45 0.104196
R10286 VSS.n5766 VSS.n5763 0.10383
R10287 VSS.n5088 VSS.n5085 0.103507
R10288 VSS.n6932 VSS.n6928 0.10325
R10289 VSS.n5071 VSS.n5070 0.103243
R10290 VSS.n5803 VSS.n5800 0.103217
R10291 VSS.n5056 VSS.n5053 0.103217
R10292 VSS.n4507 VSS.n4488 0.102601
R10293 VSS.n5628 VSS.n5626 0.102447
R10294 VSS.n5794 VSS.n5706 0.102447
R10295 VSS.n7425 VSS.n6350 0.102303
R10296 VSS.n7424 VSS.n6365 0.102303
R10297 VSS.n5800 VSS.n5797 0.102239
R10298 VSS.n5806 VSS.n5803 0.102239
R10299 VSS.n5053 VSS.n5050 0.102239
R10300 VSS.n5059 VSS.n5056 0.102239
R10301 VSS.n4281 VSS.n4280 0.101261
R10302 VSS.n1682 VSS.n1681 0.101261
R10303 VSS.n3996 VSS.n3995 0.100173
R10304 VSS.n5836 VSS.n5833 0.0999444
R10305 VSS.n5868 VSS.n5867 0.0999444
R10306 VSS.n5036 VSS.n5033 0.0999444
R10307 VSS.n5017 VSS.n5014 0.0999444
R10308 VSS.n4982 VSS.n4979 0.0999444
R10309 VSS.n4282 VSS.n4281 0.0993043
R10310 VSS.n1683 VSS.n1682 0.0993043
R10311 VSS.n5096 VSS.n5095 0.0992611
R10312 VSS.n5939 VSS.n5938 0.0990345
R10313 VSS.n4760 VSS.n4759 0.0990345
R10314 VSS.n27 VSS.n24 0.0986818
R10315 VSS.n5739 VSS.n5736 0.0984646
R10316 VSS.n5727 VSS.n5719 0.0978681
R10317 VSS.n5668 VSS.n5665 0.0974231
R10318 VSS.n5674 VSS.n5671 0.0974231
R10319 VSS.n5677 VSS.n5674 0.0974231
R10320 VSS.n5187 VSS.n5184 0.0974231
R10321 VSS.n5190 VSS.n5187 0.0974231
R10322 VSS.n5196 VSS.n5193 0.0974231
R10323 VSS.n6231 VSS.n6228 0.0973478
R10324 VSS.n6377 VSS.n6376 0.09725
R10325 VSS.n1250 VSS.n1249 0.0968905
R10326 VSS.n1127 VSS.n924 0.0965
R10327 VSS.n6913 VSS.n6912 0.0965
R10328 VSS.n5671 VSS.n5668 0.0964341
R10329 VSS.n5193 VSS.n5190 0.0964341
R10330 VSS.n5918 VSS.n5915 0.0963696
R10331 VSS.n4348 VSS.n4195 0.0963537
R10332 VSS.n7128 VSS.n7127 0.0954541
R10333 VSS.n5623 VSS.n5621 0.0952788
R10334 VSS.n7858 VSS.n7857 0.0952788
R10335 VSS.n7540 VSS.n7539 0.0950378
R10336 VSS.n5714 VSS.n5713 0.0945909
R10337 VSS.n7300 VSS 0.0945618
R10338 VSS.n5889 VSS.n5873 0.0945541
R10339 VSS.n4864 VSS.n4861 0.0942929
R10340 VSS.n6167 VSS.n6164 0.0941041
R10341 VSS.n7158 VSS.n7150 0.0941
R10342 VSS.n7138 VSS.n7128 0.0941
R10343 VSS.n4508 VSS.n4507 0.09365
R10344 VSS.n6350 VSS.n6349 0.09275
R10345 VSS.n5871 VSS.n5870 0.0922143
R10346 VSS.n5121 VSS.n5117 0.0920929
R10347 VSS.n5258 VSS.n5241 0.0914091
R10348 VSS.n5263 VSS.n5261 0.0914091
R10349 VSS.n4978 VSS.n4977 0.0913571
R10350 VSS.n1365 VSS.n1364 0.09125
R10351 VSS.n225 VSS.n224 0.0907679
R10352 VSS.n5636 VSS.n5635 0.0905
R10353 VSS.n5883 VSS.n5878 0.0905
R10354 VSS.n52 VSS.n51 0.0905
R10355 VSS.n4788 VSS.n4787 0.0905
R10356 VSS.n5218 VSS.n5216 0.0905
R10357 VSS.n4159 VSS.n4156 0.0905
R10358 VSS.n4462 VSS.n714 0.0897683
R10359 VSS.n4432 VSS.n4429 0.0897683
R10360 VSS.n5797 VSS.n5794 0.0895217
R10361 VSS.n5788 VSS.n5787 0.0889071
R10362 VSS.n5071 VSS.n5059 0.0885435
R10363 VSS.n1692 VSS.n1691 0.0883049
R10364 VSS.n5080 VSS.n5078 0.0881106
R10365 VSS.n6983 VSS.n6982 0.0877209
R10366 VSS.n6377 VSS.n6368 0.0875
R10367 VSS.n6170 VSS.n6167 0.0873421
R10368 VSS.n4867 VSS.n4864 0.0873421
R10369 VSS.n7161 VSS.n7158 0.0867185
R10370 VSS.n1536 VSS.n1535 0.0862944
R10371 VSS.n1533 VSS.n1532 0.0862944
R10372 VSS.n5992 VSS.n5989 0.0854057
R10373 VSS.n5995 VSS.n5992 0.0854057
R10374 VSS.n5998 VSS.n5995 0.0854057
R10375 VSS.n6001 VSS.n5998 0.0854057
R10376 VSS.n6004 VSS.n6001 0.0854057
R10377 VSS.n6007 VSS.n6004 0.0854057
R10378 VSS.n6010 VSS.n6007 0.0854057
R10379 VSS.n6013 VSS.n6010 0.0854057
R10380 VSS.n6016 VSS.n6013 0.0854057
R10381 VSS.n6019 VSS.n6016 0.0854057
R10382 VSS.n6022 VSS.n6019 0.0854057
R10383 VSS.n6025 VSS.n6022 0.0854057
R10384 VSS.n6028 VSS.n6025 0.0854057
R10385 VSS.n6031 VSS.n6028 0.0854057
R10386 VSS.n6102 VSS.n6099 0.0854057
R10387 VSS.n6099 VSS.n6096 0.0854057
R10388 VSS.n6096 VSS.n6093 0.0854057
R10389 VSS.n6093 VSS.n6090 0.0854057
R10390 VSS.n6086 VSS.n6083 0.0854057
R10391 VSS.n6083 VSS.n6080 0.0854057
R10392 VSS.n6080 VSS.n6077 0.0854057
R10393 VSS.n6077 VSS.n6074 0.0854057
R10394 VSS.n6071 VSS.n6068 0.0854057
R10395 VSS.n6068 VSS.n6065 0.0854057
R10396 VSS.n6065 VSS.n6062 0.0854057
R10397 VSS.n6062 VSS.n6059 0.0854057
R10398 VSS.n6059 VSS.n6056 0.0854057
R10399 VSS.n6052 VSS.n6049 0.0854057
R10400 VSS.n6049 VSS.n6045 0.0854057
R10401 VSS.n4351 VSS.n4348 0.085378
R10402 VSS.n4748 VSS.n4746 0.0846795
R10403 VSS.n5944 VSS.n5941 0.0846304
R10404 VSS.n5989 VSS.n5986 0.0843639
R10405 VSS.n5125 VSS.n5121 0.0841283
R10406 VSS.n7871 VSS.n7867 0.0841283
R10407 VSS.n5756 VSS.n5739 0.0838349
R10408 VSS.n5396 VSS.n5395 0.0838333
R10409 VSS.n5760 VSS.n5759 0.0837469
R10410 VSS.n5091 VSS.n5089 0.0832732
R10411 VSS.n6109 VSS.n6105 0.0832014
R10412 VSS.n5986 VSS.n5983 0.0830864
R10413 VSS.n5095 VSS.n5092 0.0830384
R10414 VSS.n7572 VSS.n7571 0.082937
R10415 VSS.n4913 VSS.n4912 0.0828404
R10416 VSS.n4935 VSS.n4924 0.0828404
R10417 VSS.n4733 VSS.n4731 0.0828171
R10418 VSS.n1246 VSS.n1243 0.0828171
R10419 VSS.n1243 VSS.n1240 0.0828171
R10420 VSS.n1240 VSS.n1237 0.0828171
R10421 VSS.n1237 VSS.n1234 0.0828171
R10422 VSS.n1234 VSS.n1231 0.0828171
R10423 VSS.n1231 VSS.n1228 0.0828171
R10424 VSS.n1228 VSS.n1225 0.0828171
R10425 VSS.n1225 VSS.n1222 0.0828171
R10426 VSS.n1222 VSS.n1219 0.0828171
R10427 VSS.n1219 VSS.n1216 0.0828171
R10428 VSS.n1216 VSS.n1213 0.0828171
R10429 VSS.n1213 VSS.n1210 0.0828171
R10430 VSS.n1210 VSS.n1207 0.0828171
R10431 VSS.n1207 VSS.n1204 0.0828171
R10432 VSS.n1204 VSS.n1201 0.0828171
R10433 VSS.n1201 VSS.n1198 0.0828171
R10434 VSS.n1198 VSS.n1195 0.0828171
R10435 VSS.n1195 VSS.n1192 0.0828171
R10436 VSS.n1192 VSS.n1189 0.0828171
R10437 VSS.n1189 VSS.n1186 0.0828171
R10438 VSS.n1186 VSS.n1183 0.0828171
R10439 VSS.n1183 VSS.n1180 0.0828171
R10440 VSS.n1180 VSS.n1177 0.0828171
R10441 VSS.n1177 VSS.n1174 0.0828171
R10442 VSS.n1174 VSS.n1171 0.0828171
R10443 VSS.n1171 VSS.n1168 0.0828171
R10444 VSS.n1168 VSS.n1165 0.0828171
R10445 VSS.n1165 VSS.n1162 0.0828171
R10446 VSS.n1162 VSS.n1159 0.0828171
R10447 VSS.n1159 VSS.n1156 0.0828171
R10448 VSS.n1156 VSS.n1153 0.0828171
R10449 VSS.n1153 VSS.n1150 0.0828171
R10450 VSS.n1150 VSS.n1147 0.0828171
R10451 VSS.n1147 VSS.n1144 0.0828171
R10452 VSS.n1144 VSS.n1141 0.0828171
R10453 VSS.n1141 VSS.n802 0.0828171
R10454 VSS.n19 VSS.n16 0.0828171
R10455 VSS.n7896 VSS.n19 0.0828171
R10456 VSS.n7899 VSS.n7896 0.0828171
R10457 VSS.n7902 VSS.n7899 0.0828171
R10458 VSS.n5379 VSS.n5376 0.0828171
R10459 VSS.n5254 VSS.n5244 0.0828171
R10460 VSS.n5254 VSS.n5253 0.0828171
R10461 VSS.n5253 VSS.n5250 0.0828171
R10462 VSS.n5250 VSS.n5247 0.0828171
R10463 VSS.n5271 VSS.n5268 0.0828171
R10464 VSS.n5274 VSS.n5271 0.0828171
R10465 VSS.n5277 VSS.n5274 0.0828171
R10466 VSS.n5280 VSS.n5277 0.0828171
R10467 VSS.n5284 VSS.n5280 0.0828171
R10468 VSS.n5287 VSS.n5284 0.0828171
R10469 VSS.n5290 VSS.n5287 0.0828171
R10470 VSS.n5293 VSS.n5290 0.0828171
R10471 VSS.n5298 VSS.n5293 0.0828171
R10472 VSS.n7796 VSS.n7791 0.0828171
R10473 VSS.n7791 VSS.n7788 0.0828171
R10474 VSS.n7788 VSS.n7785 0.0828171
R10475 VSS.n7785 VSS.n7781 0.0828171
R10476 VSS.n7781 VSS.n7778 0.0828171
R10477 VSS.n7778 VSS.n7775 0.0828171
R10478 VSS.n7775 VSS.n7772 0.0828171
R10479 VSS.n7772 VSS.n7769 0.0828171
R10480 VSS.n7769 VSS.n7766 0.0828171
R10481 VSS.n7766 VSS.n7763 0.0828171
R10482 VSS.n7763 VSS.n7760 0.0828171
R10483 VSS.n7760 VSS.n7757 0.0828171
R10484 VSS.n7757 VSS.n7754 0.0828171
R10485 VSS.n7754 VSS.n7751 0.0828171
R10486 VSS.n7751 VSS.n7748 0.0828171
R10487 VSS.n7748 VSS.n7744 0.0828171
R10488 VSS.n7744 VSS.n7740 0.0828171
R10489 VSS.n7483 VSS.n7480 0.0828171
R10490 VSS.n7480 VSS.n7478 0.0828171
R10491 VSS.n7478 VSS.n7475 0.0828171
R10492 VSS.n7475 VSS.n7471 0.0828171
R10493 VSS.n7471 VSS.n7468 0.0828171
R10494 VSS.n7468 VSS.n7465 0.0828171
R10495 VSS.n7465 VSS.n7462 0.0828171
R10496 VSS.n7462 VSS.n7459 0.0828171
R10497 VSS.n7459 VSS.n7456 0.0828171
R10498 VSS.n7456 VSS.n7453 0.0828171
R10499 VSS.n7453 VSS.n7450 0.0828171
R10500 VSS.n7450 VSS.n7447 0.0828171
R10501 VSS.n7447 VSS.n7444 0.0828171
R10502 VSS.n7444 VSS.n7441 0.0828171
R10503 VSS.n7441 VSS.n7438 0.0828171
R10504 VSS.n7434 VSS.n7430 0.0828171
R10505 VSS.n6327 VSS.n6324 0.0828171
R10506 VSS.n6324 VSS.n6322 0.0828171
R10507 VSS.n6322 VSS.n6319 0.0828171
R10508 VSS.n6319 VSS.n6317 0.0828171
R10509 VSS.n6317 VSS.n6314 0.0828171
R10510 VSS.n6314 VSS.n6312 0.0828171
R10511 VSS.n6312 VSS.n6309 0.0828171
R10512 VSS.n6309 VSS.n6307 0.0828171
R10513 VSS.n6307 VSS.n6304 0.0828171
R10514 VSS.n6301 VSS.n6299 0.0828171
R10515 VSS.n6299 VSS.n6296 0.0828171
R10516 VSS.n6296 VSS.n6294 0.0828171
R10517 VSS.n6294 VSS.n6291 0.0828171
R10518 VSS.n6291 VSS.n6289 0.0828171
R10519 VSS.n6289 VSS.n6286 0.0828171
R10520 VSS.n6286 VSS.n6284 0.0828171
R10521 VSS.n6284 VSS.n6282 0.0828171
R10522 VSS.n6282 VSS.n6279 0.0828171
R10523 VSS.n6279 VSS.n6272 0.0828171
R10524 VSS.n6272 VSS.n6270 0.0828171
R10525 VSS.n6263 VSS.n6260 0.0828171
R10526 VSS.n6260 VSS.n6258 0.0828171
R10527 VSS.n6258 VSS.n6255 0.0828171
R10528 VSS.n6255 VSS.n6253 0.0828171
R10529 VSS.n6249 VSS.n6247 0.0828171
R10530 VSS.n6247 VSS.n6244 0.0828171
R10531 VSS.n6244 VSS.n6242 0.0828171
R10532 VSS.n6242 VSS.n6239 0.0828171
R10533 VSS.n6239 VSS.n6237 0.0828171
R10534 VSS.n6033 VSS.n5950 0.0828171
R10535 VSS.n6035 VSS.n6033 0.0828171
R10536 VSS.n6037 VSS.n6035 0.0828171
R10537 VSS.n6039 VSS.n6037 0.0828171
R10538 VSS.n594 VSS.n591 0.0828171
R10539 VSS.n591 VSS.n588 0.0828171
R10540 VSS.n588 VSS.n585 0.0828171
R10541 VSS.n585 VSS.n582 0.0828171
R10542 VSS.n578 VSS.n575 0.0828171
R10543 VSS.n575 VSS.n572 0.0828171
R10544 VSS.n572 VSS.n569 0.0828171
R10545 VSS.n569 VSS.n566 0.0828171
R10546 VSS.n540 VSS.n537 0.0828171
R10547 VSS.n537 VSS.n534 0.0828171
R10548 VSS.n534 VSS.n531 0.0828171
R10549 VSS.n527 VSS.n524 0.0828171
R10550 VSS.n524 VSS.n521 0.0828171
R10551 VSS.n518 VSS.n514 0.0828171
R10552 VSS.n512 VSS.n508 0.0828171
R10553 VSS.n508 VSS.n505 0.0828171
R10554 VSS.n505 VSS.n502 0.0828171
R10555 VSS.n502 VSS.n500 0.0828171
R10556 VSS.n500 VSS.n497 0.0828171
R10557 VSS.n497 VSS.n494 0.0828171
R10558 VSS.n494 VSS.n491 0.0828171
R10559 VSS.n491 VSS.n488 0.0828171
R10560 VSS.n488 VSS.n485 0.0828171
R10561 VSS.n485 VSS.n482 0.0828171
R10562 VSS.n482 VSS.n479 0.0828171
R10563 VSS.n479 VSS.n476 0.0828171
R10564 VSS.n476 VSS.n473 0.0828171
R10565 VSS.n473 VSS.n470 0.0828171
R10566 VSS.n470 VSS.n467 0.0828171
R10567 VSS.n467 VSS.n464 0.0828171
R10568 VSS.n464 VSS.n461 0.0828171
R10569 VSS.n461 VSS.n458 0.0828171
R10570 VSS.n458 VSS.n455 0.0828171
R10571 VSS.n455 VSS.n452 0.0828171
R10572 VSS.n452 VSS.n449 0.0828171
R10573 VSS.n449 VSS.n446 0.0828171
R10574 VSS.n446 VSS.n443 0.0828171
R10575 VSS.n443 VSS.n440 0.0828171
R10576 VSS.n440 VSS.n437 0.0828171
R10577 VSS.n437 VSS.n434 0.0828171
R10578 VSS.n434 VSS.n431 0.0828171
R10579 VSS.n431 VSS.n428 0.0828171
R10580 VSS.n428 VSS.n425 0.0828171
R10581 VSS.n425 VSS.n422 0.0828171
R10582 VSS.n422 VSS.n420 0.0828171
R10583 VSS.n420 VSS.n416 0.0828171
R10584 VSS.n416 VSS.n413 0.0828171
R10585 VSS.n413 VSS.n410 0.0828171
R10586 VSS.n410 VSS.n407 0.0828171
R10587 VSS.n407 VSS.n404 0.0828171
R10588 VSS.n404 VSS.n401 0.0828171
R10589 VSS.n401 VSS.n398 0.0828171
R10590 VSS.n398 VSS.n393 0.0828171
R10591 VSS.n393 VSS.n389 0.0828171
R10592 VSS.n389 VSS.n386 0.0828171
R10593 VSS.n386 VSS.n383 0.0828171
R10594 VSS.n383 VSS.n381 0.0828171
R10595 VSS.n381 VSS.n378 0.0828171
R10596 VSS.n378 VSS.n375 0.0828171
R10597 VSS.n375 VSS.n372 0.0828171
R10598 VSS.n372 VSS.n369 0.0828171
R10599 VSS.n369 VSS.n366 0.0828171
R10600 VSS.n366 VSS.n363 0.0828171
R10601 VSS.n363 VSS.n360 0.0828171
R10602 VSS.n360 VSS.n357 0.0828171
R10603 VSS.n357 VSS.n353 0.0828171
R10604 VSS.n353 VSS.n350 0.0828171
R10605 VSS.n350 VSS.n347 0.0828171
R10606 VSS.n347 VSS.n344 0.0828171
R10607 VSS.n344 VSS.n341 0.0828171
R10608 VSS.n341 VSS.n338 0.0828171
R10609 VSS.n338 VSS.n335 0.0828171
R10610 VSS.n335 VSS.n331 0.0828171
R10611 VSS.n331 VSS.n327 0.0828171
R10612 VSS.n5965 VSS.n5958 0.0828171
R10613 VSS.n5968 VSS.n5965 0.0828171
R10614 VSS.n5971 VSS.n5968 0.0828171
R10615 VSS.n5974 VSS.n5971 0.0828171
R10616 VSS.n5977 VSS.n5974 0.0828171
R10617 VSS.n5980 VSS.n5977 0.0828171
R10618 VSS.n5983 VSS.n5980 0.0828171
R10619 VSS.n799 VSS.n795 0.0828171
R10620 VSS.n795 VSS.n793 0.0828171
R10621 VSS.n793 VSS.n790 0.0828171
R10622 VSS.n790 VSS.n788 0.0828171
R10623 VSS.n788 VSS.n784 0.0828171
R10624 VSS.n784 VSS.n30 0.0828171
R10625 VSS.n4742 VSS.n4739 0.0828171
R10626 VSS.n4739 VSS.n4737 0.0828171
R10627 VSS.n4737 VSS.n4733 0.0828171
R10628 VSS.n4731 VSS.n4728 0.0828171
R10629 VSS.n4728 VSS.n4725 0.0828171
R10630 VSS.n4722 VSS.n4718 0.0828171
R10631 VSS.n4715 VSS.n4712 0.0828171
R10632 VSS.n4712 VSS.n4709 0.0828171
R10633 VSS.n4709 VSS.n4707 0.0828171
R10634 VSS.n4707 VSS.n4703 0.0828171
R10635 VSS.n6232 VSS.n6231 0.0826739
R10636 VSS.n5081 VSS.n5080 0.082242
R10637 VSS.n5241 VSS.n13 0.0820721
R10638 VSS.n4149 VSS.n4145 0.0817195
R10639 VSS.n531 VSS.n528 0.0817195
R10640 VSS.n5040 VSS.n5037 0.0816957
R10641 VSS.n168 VSS.n167 0.0816607
R10642 VSS.n5537 VSS.n5536 0.0815383
R10643 VSS.n6993 VSS.n6365 0.0815
R10644 VSS.n6928 VSS.n6925 0.0815
R10645 VSS.n5787 VSS.n5779 0.0814455
R10646 VSS.n7797 VSS.n5298 0.0811707
R10647 VSS.n5732 VSS.n5731 0.0809425
R10648 VSS.n761 VSS.n760 0.0808571
R10649 VSS.n6414 VSS.n6411 0.0808571
R10650 VSS.n7233 VSS.n7232 0.0808571
R10651 VSS.n7177 VSS.n7176 0.0808571
R10652 VSS.n5351 VSS.n5350 0.0808571
R10653 VSS.n7609 VSS.n7608 0.0808571
R10654 VSS.n6685 VSS.n6684 0.0808571
R10655 VSS.n6807 VSS.n6806 0.0808571
R10656 VSS.n4608 VSS.n4596 0.0808571
R10657 VSS.n4521 VSS.n4519 0.0808571
R10658 VSS.n946 VSS.n943 0.0808571
R10659 VSS.n5837 VSS.n5816 0.0807174
R10660 VSS.n6267 VSS.n6266 0.0806219
R10661 VSS.n4716 VSS 0.0803113
R10662 VSS.n4868 VSS.n4867 0.0802368
R10663 VSS.n5104 VSS.n5100 0.080146
R10664 VSS.n204 VSS.n203 0.079766
R10665 VSS.n6175 VSS.n6170 0.0794474
R10666 VSS.n210 VSS.n209 0.0794283
R10667 VSS VSS.n756 0.07925
R10668 VSS.n6418 VSS 0.07925
R10669 VSS.n6515 VSS.n6460 0.07925
R10670 VSS.n7213 VSS.n7073 0.07925
R10671 VSS.n7181 VSS 0.07925
R10672 VSS.n7728 VSS.n7727 0.07925
R10673 VSS VSS.n7606 0.07925
R10674 VSS.n6770 VSS.n6769 0.07925
R10675 VSS VSS.n6804 0.07925
R10676 VSS.n950 VSS 0.07925
R10677 VSS.n1028 VSS.n987 0.07925
R10678 VSS.n4429 VSS.n4428 0.0787927
R10679 VSS.n5646 VSS.n5645 0.0777566
R10680 VSS.n7428 VSS.n6327 0.0773293
R10681 VSS.n4453 VSS.n4452 0.0773293
R10682 VSS.n5749 VSS.n5748 0.0770957
R10683 VSS.n4922 VSS.n4921 0.0770957
R10684 VSS.n6185 VSS.n6182 0.077079
R10685 VSS.n5208 VSS.n5205 0.0769602
R10686 VSS.n6074 VSS.n6072 0.0769151
R10687 VSS.n6108 VSS.n6106 0.076587
R10688 VSS.n4716 VSS.n4715 0.0762317
R10689 VSS VSS.n6461 0.0760357
R10690 VSS VSS.n7233 0.0760357
R10691 VSS VSS.n7609 0.0760357
R10692 VSS.n6807 VSS 0.0760357
R10693 VSS.n4481 VSS 0.0760357
R10694 VSS.n4519 VSS 0.0760357
R10695 VSS.n1005 VSS 0.0760357
R10696 VSS.n714 VSS.n713 0.0758658
R10697 VSS.n5857 VSS.n5854 0.0758261
R10698 VSS.n1413 VSS.n744 0.0755
R10699 VSS.n6531 VSS.n6430 0.0755
R10700 VSS.n7192 VSS.n7074 0.0755
R10701 VSS.n7595 VSS.n5343 0.0755
R10702 VSS.n6792 VSS.n6662 0.0755
R10703 VSS.n4321 VSS.n4319 0.0755
R10704 VSS.n1044 VSS.n961 0.0755
R10705 VSS.n6515 VSS.n6514 0.0753739
R10706 VSS.n7216 VSS.n7213 0.0753739
R10707 VSS.n6769 VSS.n6768 0.0753739
R10708 VSS.n1028 VSS.n1027 0.0753739
R10709 VSS VSS.n761 0.0752321
R10710 VSS.n6411 VSS 0.0752321
R10711 VSS.n7176 VSS 0.0752321
R10712 VSS VSS.n5351 0.0752321
R10713 VSS VSS.n6685 0.0752321
R10714 VSS.n943 VSS 0.0752321
R10715 VSS.n689 VSS.n686 0.0752
R10716 VSS.n5018 VSS.n4998 0.0748478
R10717 VSS.n6042 VSS.n6039 0.0745854
R10718 VSS.n6194 VSS 0.0739211
R10719 VSS.n5889 VSS.n5888 0.0738696
R10720 VSS.n7728 VSS.n5303 0.07325
R10721 VSS VSS.n4836 0.0731316
R10722 VSS.n173 VSS.n172 0.0728214
R10723 VSS.n6386 VSS.n6385 0.0725
R10724 VSS.n7847 VSS.n7846 0.0721814
R10725 VSS VSS.n7148 0.0718949
R10726 VSS.n1384 VSS.n1382 0.0715924
R10727 VSS.n6563 VSS.n6562 0.0715924
R10728 VSS.n1076 VSS.n1075 0.0715924
R10729 VSS.n5108 VSS.n5107 0.071385
R10730 VSS.n5259 VSS.n5258 0.0709545
R10731 VSS.n7626 VSS.n7625 0.0708361
R10732 VSS.n6818 VSS.n6817 0.0708361
R10733 VSS.n5632 VSS.n5631 0.0705885
R10734 VSS.n93 VSS.n89 0.0704107
R10735 VSS.n139 VSS.n137 0.0704107
R10736 VSS.n4608 VSS.n4607 0.0704107
R10737 VSS.n1714 VSS.n1713 0.0700122
R10738 VSS.n4687 VSS.n4674 0.0700122
R10739 VSS.n4366 VSS.n4365 0.0700122
R10740 VSS.n6235 VSS.n5950 0.0696463
R10741 VSS.n6580 VSS.n6579 0.06875
R10742 VSS.n5718 VSS.n5717 0.0687418
R10743 VSS.n4911 VSS.n4910 0.0687418
R10744 VSS.n4507 VSS.n1420 0.0685672
R10745 VSS.n5314 VSS.n5313 0.0685672
R10746 VSS.n6811 VSS.n6808 0.0685672
R10747 VSS.n5374 VSS.n5301 0.0685488
R10748 VSS.n6253 VSS.n6250 0.0685488
R10749 VSS.n6939 VSS.n6935 0.068
R10750 VSS.n1389 VSS.n1388 0.0678109
R10751 VSS.n6556 VSS.n6553 0.0678109
R10752 VSS.n7131 VSS.n7119 0.0678109
R10753 VSS.n1069 VSS.n1066 0.0678109
R10754 VSS.n1127 VSS.n1126 0.0676677
R10755 VSS.n6182 VSS.n6181 0.0676053
R10756 VSS.n5778 VSS.n5769 0.0675213
R10757 VSS.n4945 VSS.n4938 0.0675213
R10758 VSS.n6218 VSS.n6215 0.0673304
R10759 VSS.n4809 VSS.n4808 0.067297
R10760 VSS.n6161 VSS.n6158 0.0670217
R10761 VSS.n4934 VSS.n4933 0.0666326
R10762 VSS.n7571 VSS.n7568 0.0662983
R10763 VSS.n5754 VSS.n5753 0.0661354
R10764 VSS.n6505 VSS.n6461 0.0656429
R10765 VSS.n7233 VSS.n7223 0.0656429
R10766 VSS.n7544 VSS.n5351 0.0656429
R10767 VSS.n6759 VSS.n6685 0.0656429
R10768 VSS.n4482 VSS.n4481 0.0656429
R10769 VSS.n1018 VSS.n1005 0.0656429
R10770 VSS.n4666 VSS.n4664 0.0656219
R10771 VSS.n6103 VSS.n6102 0.0655943
R10772 VSS.n6053 VSS.n6052 0.0655943
R10773 VSS.n4944 VSS.n4943 0.0649262
R10774 VSS.n7547 VSS.n7544 0.0647857
R10775 VSS.n6762 VSS.n6759 0.0647857
R10776 VSS.n5777 VSS.n5776 0.0644344
R10777 VSS.n6365 VSS.n6356 0.06425
R10778 VSS.n6508 VSS.n6505 0.0640294
R10779 VSS.n7223 VSS.n7222 0.0640294
R10780 VSS.n4918 VSS.n4917 0.0640294
R10781 VSS.n4485 VSS.n4482 0.0640294
R10782 VSS.n1021 VSS.n1018 0.0640294
R10783 VSS.n1389 VSS.n761 0.0639286
R10784 VSS.n6553 VSS.n6411 0.0639286
R10785 VSS.n7176 VSS.n7119 0.0639286
R10786 VSS.n7609 VSS.n5314 0.0639286
R10787 VSS.n6808 VSS.n6807 0.0639286
R10788 VSS.n1066 VSS.n943 0.0639286
R10789 VSS.n5755 VSS.n5754 0.0636492
R10790 VSS.n4935 VSS.n4934 0.0636492
R10791 VSS.n7484 VSS.n7483 0.0636098
R10792 VSS.n7435 VSS.n7434 0.0636098
R10793 VSS.n5719 VSS.n5718 0.0633022
R10794 VSS.n4913 VSS.n4911 0.0633022
R10795 VSS.n5778 VSS.n5777 0.062959
R10796 VSS.n4945 VSS.n4944 0.062959
R10797 VSS.n556 VSS.n555 0.0626951
R10798 VSS.n7739 VSS.n5301 0.0625122
R10799 VSS.n5748 VSS.n5747 0.0622838
R10800 VSS.n4922 VSS.n4920 0.0622838
R10801 VSS.n4780 VSS.n4769 0.0621304
R10802 VSS.n7346 VSS.n7342 0.062
R10803 VSS.n5895 VSS.n5894 0.0618391
R10804 VSS.n207 VSS.n206 0.0616009
R10805 VSS.n199 VSS.n198 0.0616009
R10806 VSS.n5108 VSS.n4913 0.0613736
R10807 VSS.n7360 VSS.n7359 0.06125
R10808 VSS.n5100 VSS.n4922 0.0611892
R10809 VSS.n5021 VSS.n5018 0.0611522
R10810 VSS.n4640 VSS.n4639 0.0605
R10811 VSS.n5813 VSS.n5810 0.0603902
R10812 VSS.n5854 VSS.n5850 0.0601739
R10813 VSS.n735 VSS.n732 0.0596608
R10814 VSS.n737 VSS.n735 0.0596608
R10815 VSS.n738 VSS.n737 0.0596608
R10816 VSS.n743 VSS 0.0596608
R10817 VSS.n751 VSS.n748 0.0596608
R10818 VSS.n753 VSS.n751 0.0596608
R10819 VSS.n5514 VSS.n5511 0.0596608
R10820 VSS.n5517 VSS.n5514 0.0596608
R10821 VSS.n5518 VSS.n5517 0.0596608
R10822 VSS VSS.n5518 0.0596608
R10823 VSS.n5526 VSS.n5523 0.0596608
R10824 VSS.n5529 VSS.n5526 0.0596608
R10825 VSS.n5532 VSS.n5529 0.0596608
R10826 VSS.n5476 VSS.n5473 0.0596608
R10827 VSS.n5479 VSS.n5476 0.0596608
R10828 VSS.n5480 VSS.n5479 0.0596608
R10829 VSS VSS.n5480 0.0596608
R10830 VSS.n5488 VSS.n5485 0.0596608
R10831 VSS.n5491 VSS.n5488 0.0596608
R10832 VSS.n5494 VSS.n5491 0.0596608
R10833 VSS.n5548 VSS.n5545 0.0596608
R10834 VSS.n5551 VSS.n5548 0.0596608
R10835 VSS.n5552 VSS.n5551 0.0596608
R10836 VSS VSS.n5552 0.0596608
R10837 VSS.n5562 VSS.n5559 0.0596608
R10838 VSS.n5565 VSS.n5562 0.0596608
R10839 VSS.n5568 VSS.n5565 0.0596608
R10840 VSS.n5589 VSS.n5586 0.0596608
R10841 VSS.n5592 VSS.n5589 0.0596608
R10842 VSS.n5593 VSS.n5592 0.0596608
R10843 VSS VSS.n5593 0.0596608
R10844 VSS.n5601 VSS.n5598 0.0596608
R10845 VSS.n5604 VSS.n5601 0.0596608
R10846 VSS.n5607 VSS.n5604 0.0596608
R10847 VSS.n6457 VSS.n6454 0.0596608
R10848 VSS.n6454 VSS.n6451 0.0596608
R10849 VSS.n6451 VSS.n6448 0.0596608
R10850 VSS VSS.n6440 0.0596608
R10851 VSS.n6429 VSS.n6426 0.0596608
R10852 VSS.n6426 VSS.n6423 0.0596608
R10853 VSS.n7088 VSS.n7085 0.0596608
R10854 VSS.n7091 VSS.n7088 0.0596608
R10855 VSS.n7094 VSS.n7091 0.0596608
R10856 VSS VSS.n7195 0.0596608
R10857 VSS.n7191 VSS.n7188 0.0596608
R10858 VSS.n7188 VSS.n7185 0.0596608
R10859 VSS.n7604 VSS.n7601 0.0596608
R10860 VSS.n7601 VSS.n7598 0.0596608
R10861 VSS.n7594 VSS 0.0596608
R10862 VSS.n7587 VSS.n7586 0.0596608
R10863 VSS.n7586 VSS.n7583 0.0596608
R10864 VSS.n7583 VSS.n7580 0.0596608
R10865 VSS.n6802 VSS.n6799 0.0596608
R10866 VSS.n6799 VSS.n6796 0.0596608
R10867 VSS.n6791 VSS 0.0596608
R10868 VSS.n6784 VSS.n6783 0.0596608
R10869 VSS.n6783 VSS.n6780 0.0596608
R10870 VSS.n6780 VSS.n6777 0.0596608
R10871 VSS.n4532 VSS.n4529 0.0596608
R10872 VSS.n4534 VSS.n4532 0.0596608
R10873 VSS.n984 VSS.n981 0.0596608
R10874 VSS.n981 VSS.n978 0.0596608
R10875 VSS.n978 VSS.n975 0.0596608
R10876 VSS VSS.n967 0.0596608
R10877 VSS.n960 VSS.n957 0.0596608
R10878 VSS.n957 VSS.n954 0.0596608
R10879 VSS.n5044 VSS.n5043 0.0594119
R10880 VSS.n7125 VSS 0.0589992
R10881 VSS.n69 VSS.n65 0.0583049
R10882 VSS.n7486 VSS.n5356 0.05825
R10883 VSS.n4409 VSS.n4408 0.0574719
R10884 VSS.n4791 VSS.n4788 0.0572391
R10885 VSS.n5665 VSS.n5661 0.0568736
R10886 VSS.n5199 VSS.n5196 0.0568736
R10887 VSS.n6045 VSS.n6042 0.0559717
R10888 VSS.n136 VSS.n132 0.055378
R10889 VSS.n136 VSS.n135 0.055378
R10890 VSS.n227 VSS.n78 0.055378
R10891 VSS.n230 VSS.n227 0.055378
R10892 VSS.n4333 VSS.n4321 0.0552959
R10893 VSS.n5840 VSS.n5837 0.0552826
R10894 VSS.n738 VSS.n728 0.0552552
R10895 VSS.n5523 VSS.n5501 0.0552552
R10896 VSS.n5485 VSS.n5464 0.0552552
R10897 VSS.n5559 VSS.n5458 0.0552552
R10898 VSS.n5598 VSS.n5576 0.0552552
R10899 VSS.n6448 VSS.n6445 0.0552552
R10900 VSS.n7095 VSS.n7094 0.0552552
R10901 VSS.n7587 VSS.n5346 0.0552552
R10902 VSS.n6784 VSS.n6665 0.0552552
R10903 VSS.n975 VSS.n972 0.0552552
R10904 VSS VSS.n5031 0.0549444
R10905 VSS.n5442 VSS 0.0543889
R10906 VSS.n5037 VSS.n4949 0.0543043
R10907 VSS.n4397 VSS.n4396 0.0536953
R10908 VSS VSS.n4536 0.0533671
R10909 VSS.n4573 VSS.n4570 0.0533671
R10910 VSS.n4812 VSS.n4809 0.0530777
R10911 VSS.n6215 VSS.n6214 0.0530398
R10912 VSS.n6582 VSS.n6581 0.0528735
R10913 VSS.n7906 VSS.n7902 0.0526341
R10914 VSS.n4335 VSS.n4333 0.0522857
R10915 VSS.n7363 VSS.n7360 0.05225
R10916 VSS.n4408 VSS.n4405 0.0521084
R10917 VSS.n4396 VSS.n4393 0.0521084
R10918 VSS.n5746 VSS.n5745 0.0514211
R10919 VSS.n5538 VSS.n5498 0.0513891
R10920 VSS.n5890 VSS.n5401 0.0513696
R10921 VSS.n4586 VSS.n4584 0.0508497
R10922 VSS.n4743 VSS.n30 0.050439
R10923 VSS.n7423 VSS.n6582 0.0504242
R10924 VSS.n6505 VSS.n6504 0.050416
R10925 VSS.n7238 VSS.n7223 0.050416
R10926 VSS.n4482 VSS.n1475 0.050416
R10927 VSS.n1018 VSS.n1017 0.050416
R10928 VSS.n4643 VSS.n4640 0.0502561
R10929 VSS.n528 VSS.n527 0.0498902
R10930 VSS.n4723 VSS.n4722 0.0498902
R10931 VSS.n5635 VSS.n5632 0.0498805
R10932 VSS.n692 VSS.n691 0.0496753
R10933 VSS.n7544 VSS.n7543 0.0496597
R10934 VSS.n6759 VSS.n6758 0.0496597
R10935 VSS.n7740 VSS.n7739 0.0493415
R10936 VSS.n814 VSS.n813 0.048782
R10937 VSS.n5264 VSS.n5263 0.0486818
R10938 VSS.n6090 VSS.n6087 0.0486132
R10939 VSS.n4419 VSS.n4416 0.0483322
R10940 VSS.n7484 VSS.n5379 0.0482439
R10941 VSS.n4701 VSS.n594 0.0476951
R10942 VSS.n5365 VSS.n5364 0.047
R10943 VSS.n4933 VSS.n4926 0.0468235
R10944 VSS.n1393 VSS.n1389 0.0466345
R10945 VSS.n6553 VSS.n6552 0.0466345
R10946 VSS.n7119 VSS.n7118 0.0466345
R10947 VSS.n1066 VSS.n1065 0.0466345
R10948 VSS.n4840 VSS 0.0462895
R10949 VSS VSS.n5439 0.0460556
R10950 VSS.n5322 VSS.n5314 0.0458782
R10951 VSS.n4664 VSS.n4658 0.0458659
R10952 VSS.n4316 VSS.n4314 0.0458659
R10953 VSS.n4920 VSS.n4919 0.0457432
R10954 VSS VSS.n6191 0.0455
R10955 VSS.n5945 VSS.n5936 0.0455
R10956 VSS.n5032 VSS 0.0455
R10957 VSS.n5747 VSS.n5746 0.0452568
R10958 VSS.n5776 VSS.n5771 0.04425
R10959 VSS.n4943 VSS.n4940 0.04425
R10960 VSS.n756 VSS.n754 0.0439266
R10961 VSS.n5542 VSS.n5541 0.0439266
R10962 VSS.n5583 VSS.n5582 0.0439266
R10963 VSS.n6419 VSS.n6418 0.0439266
R10964 VSS.n7182 VSS.n7181 0.0439266
R10965 VSS.n7606 VSS.n7605 0.0439266
R10966 VSS.n6804 VSS.n6803 0.0439266
R10967 VSS.n4527 VSS.n4526 0.0439266
R10968 VSS.n951 VSS.n950 0.0439266
R10969 VSS.n7629 VSS.n7626 0.0436092
R10970 VSS.n6821 VSS.n6818 0.0436092
R10971 VSS.n5883 VSS.n5882 0.0435435
R10972 VSS.n5205 VSS.n5204 0.0435088
R10973 VSS.n5376 VSS.n5374 0.0433049
R10974 VSS.n7438 VSS.n7435 0.0433049
R10975 VSS.n7339 VSS.n7336 0.04325
R10976 VSS.n1382 VSS.n1381 0.0428529
R10977 VSS.n6566 VSS.n6563 0.0428529
R10978 VSS.n7162 VSS.n7161 0.0428529
R10979 VSS.n1079 VSS.n1076 0.0428529
R10980 VSS.n5649 VSS.n5646 0.0427124
R10981 VSS.n4916 VSS.n4915 0.0426277
R10982 VSS.n1589 VSS.n1492 0.0425561
R10983 VSS.n6264 VSS.n6263 0.0422073
R10984 VSS.n7568 VSS.n7564 0.0413403
R10985 VSS.n6266 VSS.n6264 0.0411098
R10986 VSS.n27 VSS.n26 0.0407128
R10987 VSS.n5100 VSS.n5099 0.040323
R10988 VSS.n1607 VSS.n1606 0.0401503
R10989 VSS.n5735 VSS.n5732 0.0395266
R10990 VSS.n7349 VSS.n7346 0.0395
R10991 VSS.n7906 VSS.n7905 0.0394634
R10992 VSS.n6518 VSS.n6515 0.0390714
R10993 VSS.n7213 VSS.n7212 0.0390714
R10994 VSS.n6769 VSS.n6680 0.0390714
R10995 VSS.n1031 VSS.n1028 0.0390714
R10996 VSS.n6955 VSS.n6939 0.03875
R10997 VSS.n4767 VSS.n4764 0.0386522
R10998 VSS.n4456 VSS.n4453 0.0385488
R10999 VSS.n6350 VSS.n6338 0.038
R11000 VSS.n744 VSS.n743 0.0376329
R11001 VSS.n6440 VSS.n6430 0.0376329
R11002 VSS.n7195 VSS.n7192 0.0376329
R11003 VSS.n7595 VSS.n7594 0.0376329
R11004 VSS.n6792 VSS.n6791 0.0376329
R11005 VSS.n967 VSS.n961 0.0376329
R11006 VSS.n6198 VSS.n6195 0.0376053
R11007 VSS.n6087 VSS.n6086 0.0372925
R11008 VSS.n1786 VSS.n1785 0.0368785
R11009 VSS.n1790 VSS.n1789 0.0368564
R11010 VSS.n582 VSS.n579 0.0367195
R11011 VSS.n5945 VSS.n5944 0.0366957
R11012 VSS.n5616 VSS.n5614 0.0363407
R11013 VSS.n7867 VSS.n7866 0.0363407
R11014 VSS.n7138 VSS.n7137 0.0360462
R11015 VSS.n7162 VSS.n7138 0.0360462
R11016 VSS.n1488 VSS.n1487 0.0357448
R11017 VSS.n4753 VSS.n4752 0.0352779
R11018 VSS.n5909 VSS.n5908 0.0352465
R11019 VSS.n730 VSS.n725 0.0351154
R11020 VSS.n5536 VSS.n5533 0.0351154
R11021 VSS.n5498 VSS.n5495 0.0351154
R11022 VSS.n5572 VSS.n5569 0.0351154
R11023 VSS.n5611 VSS.n5608 0.0351154
R11024 VSS.n6459 VSS.n6458 0.0351154
R11025 VSS.n7082 VSS.n7081 0.0351154
R11026 VSS.n7577 VSS.n7576 0.0351154
R11027 VSS.n6774 VSS.n6773 0.0351154
R11028 VSS.n4574 VSS.n4573 0.0351154
R11029 VSS.n4590 VSS.n4587 0.0351154
R11030 VSS.n4370 VSS.n4369 0.0351154
R11031 VSS.n986 VSS.n985 0.0351154
R11032 VSS.n7846 VSS.n5221 0.0347478
R11033 VSS.n4383 VSS.n4382 0.034486
R11034 VSS.n4098 VSS.n4094 0.0339302
R11035 VSS.n7620 VSS.n7619 0.0334464
R11036 VSS.n6627 VSS.n6624 0.0334464
R11037 VSS.n4514 VSS.n718 0.0334464
R11038 VSS.n566 VSS.n563 0.0334268
R11039 VSS.n4725 VSS.n4723 0.0334268
R11040 VSS.n5111 VSS.n5109 0.0331549
R11041 VSS.n4743 VSS.n4742 0.032878
R11042 VSS.n4535 VSS.n4534 0.0325979
R11043 VSS.n5078 VSS.n5077 0.0323584
R11044 VSS.n3226 VSS.n1970 0.0323182
R11045 VSS.n1866 VSS.n1801 0.0320446
R11046 VSS.n1772 VSS.n1771 0.032
R11047 VSS.n1878 VSS.n1873 0.032
R11048 VSS.n1762 VSS.n1761 0.032
R11049 VSS.n4420 VSS.n4419 0.0319685
R11050 VSS.n7834 VSS.n7830 0.0318333
R11051 VSS.n7830 VSS.n7826 0.0318333
R11052 VSS.n7826 VSS.n7822 0.0318333
R11053 VSS VSS.n7815 0.0318333
R11054 VSS.n7815 VSS.n7814 0.0318333
R11055 VSS.n7814 VSS.n7810 0.0318333
R11056 VSS.n7810 VSS.n7806 0.0318333
R11057 VSS.n4278 VSS.n4277 0.0318043
R11058 VSS.n1677 VSS.n1676 0.0318043
R11059 VSS.n5790 VSS.n5788 0.0315619
R11060 VSS.n1780 VSS.n1779 0.0309839
R11061 VSS.n6977 VSS.n6976 0.0308614
R11062 VSS.n211 VSS.n210 0.0305726
R11063 VSS.n5639 VSS.n5636 0.029969
R11064 VSS.n5216 VSS.n5215 0.029969
R11065 VSS.n7822 VSS.n5228 0.0295
R11066 VSS.n694 VSS.n693 0.0292629
R11067 VSS.n7888 VSS.n21 0.0291624
R11068 VSS.n7892 VSS.n7888 0.0291624
R11069 VSS VSS.n1 0.0291624
R11070 VSS VSS.n7909 0.0291624
R11071 VSS.n1807 VSS.n1806 0.0291175
R11072 VSS.n1715 VSS.n1714 0.0290366
R11073 VSS.n1136 VSS.n21 0.0290191
R11074 VSS.n2602 VSS.n2592 0.0289279
R11075 VSS.n4541 VSS.n595 0.0288217
R11076 VSS.n3699 VSS.n3693 0.028625
R11077 VSS.n772 VSS.n770 0.028625
R11078 VSS.n183 VSS.n180 0.028625
R11079 VSS.n6406 VSS.n6403 0.028625
R11080 VSS.n6492 VSS.n6491 0.028625
R11081 VSS.n7227 VSS.n7226 0.028625
R11082 VSS.n7171 VSS.n7168 0.028625
R11083 VSS.n6948 VSS.n6947 0.028625
R11084 VSS.n7619 VSS.n7616 0.028625
R11085 VSS.n6747 VSS.n6744 0.028625
R11086 VSS.n6630 VSS.n6627 0.028625
R11087 VSS.n86 VSS.n83 0.028625
R11088 VSS.n4604 VSS.n4601 0.028625
R11089 VSS.n4478 VSS.n4477 0.028625
R11090 VSS.n4515 VSS.n4514 0.028625
R11091 VSS.n938 VSS.n935 0.028625
R11092 VSS.n995 VSS.n992 0.028625
R11093 VSS.n1250 VSS.n799 0.0284878
R11094 VSS.n597 VSS.n596 0.0284
R11095 VSS.n5117 VSS.n5116 0.0283761
R11096 VSS.n693 VSS.n692 0.0283351
R11097 VSS.n6714 VSS.n6610 0.0282695
R11098 VSS.n4420 VSS.n4373 0.0281923
R11099 VSS.n6211 VSS.n6210 0.0281316
R11100 VSS.n7158 VSS.n7157 0.0277269
R11101 VSS.n1834 VSS.n1833 0.0276659
R11102 VSS.n5724 VSS.n5721 0.0275796
R11103 VSS.n1796 VSS.n1795 0.0274585
R11104 VSS.n5744 VSS.n5743 0.0273085
R11105 VSS.n26 VSS.n25 0.0273085
R11106 VSS.n7908 VSS.n13 0.0272994
R11107 VSS.n53 VSS.n32 0.026913
R11108 VSS.n4117 VSS.n4116 0.0266
R11109 VSS.n4108 VSS.n4107 0.0266
R11110 VSS.n4097 VSS.n4096 0.0266
R11111 VSS.n4878 VSS.n4877 0.0265939
R11112 VSS.n1586 VSS.n1493 0.0265748
R11113 VSS.n1532 VSS.n1531 0.0265748
R11114 VSS.n2952 VSS.n2951 0.0262358
R11115 VSS.n5904 VSS.n5902 0.0261799
R11116 VSS.n2001 VSS.n2000 0.0261034
R11117 VSS.n209 VSS.n208 0.0260963
R11118 VSS.n5901 VSS.n5900 0.0259717
R11119 VSS.n4880 VSS.n4879 0.0259717
R11120 VSS.n4074 VSS.n4073 0.0258911
R11121 VSS.n4340 VSS.n4339 0.0258571
R11122 VSS.n1530 VSS.n1529 0.0257336
R11123 VSS.n1531 VSS.n1492 0.0257336
R11124 VSS.n1768 VSS.n1767 0.0257
R11125 VSS.n1875 VSS.n1874 0.0257
R11126 VSS.n1758 VSS.n1757 0.0257
R11127 VSS.n616 VSS.n613 0.0256748
R11128 VSS.n622 VSS.n619 0.0256748
R11129 VSS.n628 VSS.n625 0.0256748
R11130 VSS.n656 VSS.n653 0.0256748
R11131 VSS.n663 VSS.n660 0.0256748
R11132 VSS.n1518 VSS.n1515 0.0256748
R11133 VSS.n1524 VSS.n1521 0.0256748
R11134 VSS.n1581 VSS.n1578 0.0256748
R11135 VSS.n1575 VSS.n1572 0.0256748
R11136 VSS.n1817 VSS.n1816 0.0255922
R11137 VSS.n2342 VSS.n2294 0.0254833
R11138 VSS.n1804 VSS.n1803 0.0253848
R11139 VSS.n688 VSS.n687 0.0253571
R11140 VSS.n2235 VSS.n2223 0.0253328
R11141 VSS.n2451 VSS.n2415 0.0253328
R11142 VSS.n208 VSS.n207 0.0252706
R11143 VSS.n205 VSS.n204 0.0252706
R11144 VSS.n6925 VSS.n6919 0.02525
R11145 VSS.n5621 VSS.n5620 0.0251903
R11146 VSS.n7860 VSS.n7858 0.0251903
R11147 VSS.n2231 VSS.n2230 0.0251823
R11148 VSS.n2016 VSS.n2015 0.0251724
R11149 VSS.n732 VSS.n730 0.0250455
R11150 VSS.n5533 VSS.n5532 0.0250455
R11151 VSS.n5495 VSS.n5494 0.0250455
R11152 VSS.n5569 VSS.n5568 0.0250455
R11153 VSS.n5608 VSS.n5607 0.0250455
R11154 VSS.n6458 VSS.n6457 0.0250455
R11155 VSS.n7085 VSS.n7082 0.0250455
R11156 VSS.n7580 VSS.n7577 0.0250455
R11157 VSS.n6777 VSS.n6774 0.0250455
R11158 VSS.n1585 VSS.n1559 0.0250455
R11159 VSS.n4587 VSS.n4586 0.0250455
R11160 VSS.n4373 VSS.n4370 0.0250455
R11161 VSS.n985 VSS.n984 0.0250455
R11162 VSS.n2592 VSS.n2576 0.0249978
R11163 VSS.n1792 VSS 0.0247376
R11164 VSS.n630 VSS.n629 0.0247308
R11165 VSS.n5908 VSS.n5907 0.0247308
R11166 VSS.n7572 VSS.n7554 0.0247017
R11167 VSS.n91 VSS.n90 0.024574
R11168 VSS.n2242 VSS.n2241 0.0244298
R11169 VSS.n1966 VSS.n1965 0.0243636
R11170 VSS.n1846 VSS.n1845 0.0241406
R11171 VSS.n521 VSS.n518 0.0240976
R11172 VSS.n6228 VSS.n6227 0.0239783
R11173 VSS.n1961 VSS.n1960 0.0236818
R11174 VSS.n1963 VSS.n1959 0.0236818
R11175 VSS.n1827 VSS.n1826 0.0235184
R11176 VSS.n7802 VSS.n7801 0.0235
R11177 VSS.n5897 VSS.n5896 0.0234789
R11178 VSS.n3754 VSS.n3753 0.0233924
R11179 VSS.n5047 VSS.n5044 0.0232368
R11180 VSS VSS.n6984 0.0231603
R11181 VSS.n4884 VSS.n4883 0.0230525
R11182 VSS.n5890 VSS.n5889 0.023
R11183 VSS.n3698 VSS.n3697 0.0228692
R11184 VSS.n3101 VSS.n3100 0.0228692
R11185 VSS.n5810 VSS.n5809 0.0227632
R11186 VSS.n748 VSS.n744 0.022528
R11187 VSS.n6430 VSS.n6429 0.022528
R11188 VSS.n7192 VSS.n7191 0.022528
R11189 VSS.n7598 VSS.n7595 0.022528
R11190 VSS.n6796 VSS.n6792 0.022528
R11191 VSS.n961 VSS.n960 0.022528
R11192 VSS.n2652 VSS.n2651 0.0225087
R11193 VSS.n4062 VSS.n4061 0.0221201
R11194 VSS.n4902 VSS.n4901 0.0220702
R11195 VSS.n1858 VSS.n1857 0.0220668
R11196 VSS.n5736 VSS.n5735 0.0220044
R11197 VSS.n159 VSS.n154 0.0217195
R11198 VSS.n170 VSS.n169 0.0213929
R11199 VSS.n5921 VSS.n5920 0.0213264
R11200 VSS.n5924 VSS.n5923 0.0213264
R11201 VSS.n4899 VSS.n4898 0.0213264
R11202 VSS.n4752 VSS.n4751 0.0212692
R11203 VSS.n5099 VSS.n5096 0.021208
R11204 VSS.n5261 VSS.n5259 0.0209545
R11205 VSS.n5717 VSS.n5714 0.0209545
R11206 VSS.n4910 VSS.n27 0.0209545
R11207 VSS.n4883 VSS.n4882 0.0208774
R11208 VSS.n3060 VSS.n3059 0.020815
R11209 VSS.n143 VSS.n141 0.0207174
R11210 VSS.n214 VSS.n165 0.0207174
R11211 VSS.n1545 VSS 0.0206399
R11212 VSS.n2292 VSS.n2283 0.0205167
R11213 VSS.n2413 VSS.n2412 0.0205167
R11214 VSS.n5089 VSS.n5088 0.0204115
R11215 VSS.n2567 VSS.n2523 0.0203837
R11216 VSS.n197 VSS.n196 0.0203165
R11217 VSS.n6103 VSS.n6031 0.0203113
R11218 VSS.n6056 VSS.n6053 0.0203113
R11219 VSS.n2706 VSS.n2593 0.0201507
R11220 VSS.n39 VSS.n38 0.0200652
R11221 VSS.n143 VSS.n142 0.0200652
R11222 VSS.n214 VSS.n213 0.0200652
R11223 VSS.n6174 VSS.n6173 0.0200447
R11224 VSS.n5898 VSS.n5897 0.0200283
R11225 VSS.n4120 VSS.n4111 0.0200225
R11226 VSS.n4555 VSS.n4554 0.0199845
R11227 VSS.n3670 VSS.n3669 0.0198605
R11228 VSS.n4896 VSS.n4895 0.0198388
R11229 VSS.n194 VSS.n173 0.0197857
R11230 VSS.n4893 VSS.n4892 0.0197025
R11231 VSS.n5763 VSS.n5760 0.019615
R11232 VSS.n4904 VSS.n4894 0.0196091
R11233 VSS.n2731 VSS.n2559 0.0195988
R11234 VSS.n147 VSS.n146 0.0195947
R11235 VSS.n5411 VSS.n5410 0.019555
R11236 VSS.n5431 VSS.n5430 0.019555
R11237 VSS.n1724 VSS.n1723 0.0195244
R11238 VSS.n4309 VSS.n4308 0.0195244
R11239 VSS.n2704 VSS.n2594 0.0193646
R11240 VSS.n5447 VSS.n5446 0.0193395
R11241 VSS.n4872 VSS.n4871 0.0191251
R11242 VSS.n5927 VSS.n5926 0.019095
R11243 VSS.n41 VSS.n39 0.019087
R11244 VSS.n3628 VSS.n3627 0.0190756
R11245 VSS.n4552 VSS.n4551 0.0190567
R11246 VSS.n2872 VSS.n2364 0.0190117
R11247 VSS.n188 VSS.n187 0.0189821
R11248 VSS.n3788 VSS.n3787 0.0189448
R11249 VSS.n149 VSS.n148 0.0188673
R11250 VSS.n2733 VSS.n2565 0.018814
R11251 VSS.n1749 VSS.n1747 0.0187927
R11252 VSS.n4292 VSS.n4290 0.0187927
R11253 VSS.n5830 VSS.n5829 0.0186836
R11254 VSS.n5434 VSS.n5433 0.0186836
R11255 VSS.n5416 VSS.n5413 0.0186836
R11256 VSS.n203 VSS.n202 0.0186651
R11257 VSS.n2702 VSS.n2595 0.0185786
R11258 VSS.n4378 VSS.n4377 0.0185
R11259 VSS.n690 VSS.n689 0.0185
R11260 VSS.n4775 VSS.n4774 0.018485
R11261 VSS.n5926 VSS.n5925 0.0184602
R11262 VSS.n1528 VSS.n1527 0.0184371
R11263 VSS.n2082 VSS.n2081 0.0183448
R11264 VSS.n3617 VSS.n3616 0.0182907
R11265 VSS.n2345 VSS.n2332 0.0182592
R11266 VSS.n4562 VSS.n4561 0.0181289
R11267 VSS.n2870 VSS.n2365 0.0181087
R11268 VSS.n4764 VSS.n4763 0.0181087
R11269 VSS.n5929 VSS.n5928 0.0181073
R11270 VSS.n4897 VSS.n4896 0.0180867
R11271 VSS.n2736 VSS.n2735 0.0180291
R11272 VSS.n5626 VSS.n5625 0.0180221
R11273 VSS.n5794 VSS.n5793 0.0180221
R11274 VSS.n201 VSS.n200 0.0178394
R11275 VSS.n4966 VSS.n4963 0.0178182
R11276 VSS.n4953 VSS.n4950 0.0178182
R11277 VSS.n5006 VSS.n5003 0.0178182
R11278 VSS.n2227 VSS.n2226 0.0178077
R11279 VSS.n607 VSS.n606 0.0178077
R11280 VSS.n673 VSS.n672 0.0178077
R11281 VSS.n1509 VSS.n1508 0.0178077
R11282 VSS.n1566 VSS.n1565 0.0178077
R11283 VSS.n921 VSS.n920 0.01775
R11284 VSS.n2403 VSS.n2363 0.0176572
R11285 VSS.n3695 VSS.n3694 0.0176366
R11286 VSS.n1770 VSS.n1769 0.0175923
R11287 VSS.n1760 VSS.n1759 0.0175923
R11288 VSS.n4379 VSS.n4376 0.0175
R11289 VSS.n680 VSS.n666 0.017493
R11290 VSS.n778 VSS.n773 0.0174458
R11291 VSS.n6400 VSS.n6398 0.0174458
R11292 VSS.n7165 VSS.n7164 0.0174458
R11293 VSS.n932 VSS.n930 0.0174458
R11294 VSS.n6403 VSS.n6400 0.0173807
R11295 VSS.n7168 VSS.n7165 0.0173807
R11296 VSS.n773 VSS.n772 0.0173807
R11297 VSS.n935 VSS.n932 0.0173807
R11298 VSS.n2518 VSS.n2517 0.017375
R11299 VSS.n169 VSS.n168 0.017375
R11300 VSS.n172 VSS.n171 0.017375
R11301 VSS.n2882 VSS.n2881 0.0173562
R11302 VSS.n4319 VSS.n4318 0.0173367
R11303 VSS.n5074 VSS.n5071 0.0172257
R11304 VSS.n2868 VSS.n2366 0.0172057
R11305 VSS.n777 VSS.n774 0.0171955
R11306 VSS.n7124 VSS.n7121 0.0171955
R11307 VSS.n53 VSS.n52 0.0171304
R11308 VSS.n161 VSS.n160 0.0170306
R11309 VSS.n2083 VSS.n2082 0.0169483
R11310 VSS.n3226 VSS.n3225 0.0167984
R11311 VSS.n2228 VSS.n2227 0.0167542
R11312 VSS.n1491 VSS.n1490 0.0165
R11313 VSS.n2226 VSS.n2140 0.0164532
R11314 VSS.n2357 VSS.n2330 0.0164532
R11315 VSS.n5109 VSS.n5108 0.0164292
R11316 VSS.n4559 VSS.n4558 0.0162732
R11317 VSS.n754 VSS.n753 0.0162343
R11318 VSS.n5511 VSS.n5508 0.0162343
R11319 VSS.n5473 VSS.n5470 0.0162343
R11320 VSS.n5545 VSS.n5542 0.0162343
R11321 VSS.n5586 VSS.n5583 0.0162343
R11322 VSS.n6423 VSS.n6419 0.0162343
R11323 VSS.n7185 VSS.n7182 0.0162343
R11324 VSS.n7605 VSS.n7604 0.0162343
R11325 VSS.n6803 VSS.n6802 0.0162343
R11326 VSS.n4529 VSS.n4527 0.0162343
R11327 VSS.n954 VSS.n951 0.0162343
R11328 VSS.n2708 VSS.n2591 0.0162205
R11329 VSS.n5844 VSS.n5841 0.0161522
R11330 VSS.n215 VSS.n164 0.0161122
R11331 VSS.n3572 VSS.n3571 0.0160669
R11332 VSS.n563 VSS.n540 0.0158659
R11333 VSS.n5923 VSS.n5922 0.015852
R11334 VSS.n684 VSS.n683 0.0158
R11335 VSS.n7892 VSS.n7891 0.0156911
R11336 VSS.n1553 VSS 0.0156049
R11337 VSS.n2099 VSS.n2098 0.0155517
R11338 VSS.n1596 VSS.n1491 0.0155
R11339 VSS.n2710 VSS.n2587 0.0154345
R11340 VSS.n2334 VSS.n2282 0.0153997
R11341 VSS.n5900 VSS.n5899 0.015398
R11342 VSS.n2453 VSS.n2452 0.0152492
R11343 VSS.n5028 VSS.n5027 0.0151739
R11344 VSS.n5920 VSS.n5919 0.0151082
R11345 VSS.n4900 VSS.n4899 0.0151082
R11346 VSS.n2968 VSS.n2204 0.0150987
R11347 VSS.n3757 VSS.n3756 0.0150203
R11348 VSS.n3562 VSS.n3561 0.0148895
R11349 VSS.n5729 VSS.n5727 0.0148363
R11350 VSS.n5905 VSS.n5895 0.0148234
R11351 VSS.n4749 VSS.n4748 0.0148073
R11352 VSS.n6250 VSS.n6249 0.0147683
R11353 VSS.n4903 VSS.n4902 0.0147345
R11354 VSS.n650 VSS.n599 0.0146608
R11355 VSS.n2713 VSS.n2712 0.0146485
R11356 VSS.n3782 VSS.n3781 0.0146279
R11357 VSS.n1995 VSS.n1994 0.0146207
R11358 VSS.n4881 VSS.n4880 0.014549
R11359 VSS.n2897 VSS.n2896 0.0144967
R11360 VSS.n2116 VSS.n2115 0.0144655
R11361 VSS.n151 VSS.n140 0.0144024
R11362 VSS.n3071 VSS.n3070 0.0143663
R11363 VSS.n2829 VSS.n2828 0.0143462
R11364 VSS.n2970 VSS.n2201 0.0141957
R11365 VSS.n6979 VSS.n6978 0.0141817
R11366 VSS.n223 VSS.n222 0.0141607
R11367 VSS.n193 VSS 0.0141607
R11368 VSS.n1589 VSS.n1588 0.0141607
R11369 VSS.n3689 VSS.n3688 0.0141047
R11370 VSS.n3023 VSS.n2141 0.0140452
R11371 VSS.n5629 VSS.n5628 0.0140398
R11372 VSS.n7850 VSS.n7847 0.0140398
R11373 VSS.n4090 VSS.n4089 0.0140123
R11374 VSS.n4123 VSS.n4122 0.0140123
R11375 VSS.n7891 VSS.n1 0.0139713
R11376 VSS.n1537 VSS.n1536 0.0139579
R11377 VSS.n7836 VSS.n7835 0.0138333
R11378 VSS.n2681 VSS.n2680 0.0137314
R11379 VSS.n2032 VSS.n2031 0.0136897
R11380 VSS.n6237 VSS.n6235 0.0136707
R11381 VSS.n2317 VSS.n2314 0.0135936
R11382 VSS.n2121 VSS.n2120 0.0135345
R11383 VSS.n7835 VSS.n7834 0.0135
R11384 VSS.n4558 VSS.n4557 0.0134897
R11385 VSS.n2439 VSS.n2435 0.0134431
R11386 VSS.n3658 VSS.n3657 0.0133198
R11387 VSS.n2973 VSS.n2972 0.0132926
R11388 VSS.n1970 VSS.n1969 0.0132273
R11389 VSS.n3089 VSS.n3088 0.013189
R11390 VSS.n3021 VSS.n2142 0.0131421
R11391 VSS.n4550 VSS.n4549 0.0130874
R11392 VSS.n2618 VSS.n2615 0.0129454
R11393 VSS.n2079 VSS.n2078 0.0126034
R11394 VSS.n7543 VSS.n7540 0.0126008
R11395 VSS.n4000 VSS.n3999 0.0125737
R11396 VSS.n579 VSS.n578 0.0125732
R11397 VSS.n3730 VSS.n3729 0.0125349
R11398 VSS.n4379 VSS.n4378 0.0125
R11399 VSS.n4564 VSS.n4563 0.012458
R11400 VSS.n164 VSS.n163 0.0124388
R11401 VSS.n5756 VSS.n5755 0.0124337
R11402 VSS.n4932 VSS.n4931 0.0124337
R11403 VSS.n4909 VSS.n4908 0.0123681
R11404 VSS.n5779 VSS.n5778 0.0123033
R11405 VSS.n4942 VSS.n4941 0.0123033
R11406 VSS.n1538 VSS.n1537 0.0122757
R11407 VSS.n3019 VSS.n2143 0.0122391
R11408 VSS.n683 VSS.n682 0.0122
R11409 VSS.n2639 VSS.n2637 0.0121594
R11410 VSS.n6302 VSS.n6301 0.0120244
R11411 VSS.n4918 VSS.n4916 0.0119894
R11412 VSS.n5752 VSS.n5750 0.0119365
R11413 VSS.n5092 VSS.n4935 0.0119365
R11414 VSS.n5716 VSS.n5715 0.0118736
R11415 VSS.n4416 VSS.n4415 0.0118287
R11416 VSS.n5775 VSS.n5772 0.0118115
R11417 VSS.n5081 VSS.n4945 0.0118115
R11418 VSS.n2941 VSS.n2248 0.0117876
R11419 VSS.n137 VSS.n93 0.01175
R11420 VSS.n2756 VSS.n2524 0.0116192
R11421 VSS.n146 VSS.n145 0.0115204
R11422 VSS.n5774 VSS.n5773 0.0113172
R11423 VSS.n4926 VSS.n4925 0.0113172
R11424 VSS.n4385 VSS.n4384 0.0111993
R11425 VSS.n2243 VSS.n2239 0.0111355
R11426 VSS.n224 VSS.n223 0.0109464
R11427 VSS.n770 VSS.n767 0.0109464
R11428 VSS.n186 VSS.n183 0.0109464
R11429 VSS.n6409 VSS.n6406 0.0109464
R11430 VSS.n7174 VSS.n7171 0.0109464
R11431 VSS.n6949 VSS.n6948 0.0109464
R11432 VSS.n6744 VSS.n6743 0.0109464
R11433 VSS.n4607 VSS.n4604 0.0109464
R11434 VSS.n941 VSS.n938 0.0109464
R11435 VSS.n4102 VSS.n4093 0.0109366
R11436 VSS.n2939 VSS.n2249 0.0108846
R11437 VSS.n2758 VSS.n2544 0.0108343
R11438 VSS VSS.n1692 0.0107439
R11439 VSS.n4561 VSS.n4560 0.0107062
R11440 VSS.n4106 VSS.n4105 0.0106256
R11441 VSS.n2807 VSS.n2473 0.0105727
R11442 VSS.n1556 VSS.n1553 0.0105699
R11443 VSS.n4576 VSS.n4575 0.0105699
R11444 VSS.n4382 VSS.n1607 0.0105699
R11445 VSS.n2290 VSS.n2289 0.0104331
R11446 VSS.n2851 VSS.n2850 0.0104331
R11447 VSS.n3236 VSS.n3235 0.0103111
R11448 VSS.n598 VSS.n597 0.0102958
R11449 VSS.n4115 VSS.n4114 0.0102906
R11450 VSS.n6916 VSS.n6913 0.01025
R11451 VSS.n779 VSS.n778 0.0101429
R11452 VSS.n6398 VSS.n6393 0.0101429
R11453 VSS.n6491 VSS.n6490 0.0101429
R11454 VSS.n7228 VSS.n7227 0.0101429
R11455 VSS.n7164 VSS.n7163 0.0101429
R11456 VSS.n7616 VSS.n7613 0.0101429
R11457 VSS.n6633 VSS.n6630 0.0101429
R11458 VSS.n89 VSS.n86 0.0101429
R11459 VSS.n1590 VSS.n1589 0.0101429
R11460 VSS.n4479 VSS.n4478 0.0101429
R11461 VSS.n4516 VSS.n4515 0.0101429
R11462 VSS.n930 VSS.n925 0.0101429
R11463 VSS.n998 VSS.n995 0.0101429
R11464 VSS.n4017 VSS.n4016 0.0100852
R11465 VSS.n2761 VSS.n2760 0.0100494
R11466 VSS.n3759 VSS.n3758 0.0100494
R11467 VSS.n226 VSS.n159 0.0100122
R11468 VSS.n4084 VSS.n4083 0.0100029
R11469 VSS.n2937 VSS.n2250 0.00998161
R11470 VSS.n5779 VSS.n5766 0.00997368
R11471 VSS.n1606 VSS.n1605 0.00994056
R11472 VSS.n1598 VSS.n1597 0.00994056
R11473 VSS.n4045 VSS.n4044 0.00989535
R11474 VSS.n3959 VSS.n3958 0.00982401
R11475 VSS.n2805 VSS.n2474 0.00978779
R11476 VSS.n4553 VSS.n4552 0.00977835
R11477 VSS.n4562 VSS.n4555 0.00977835
R11478 VSS.n3109 VSS.n3108 0.00974419
R11479 VSS.n150 VSS.n149 0.00968367
R11480 VSS.n2283 VSS.n2258 0.0096806
R11481 VSS.n1799 VSS 0.00958911
R11482 VSS.n2917 VSS.n2916 0.0095301
R11483 VSS.n2385 VSS.n2382 0.0095301
R11484 VSS.n2485 VSS.n2472 0.00952616
R11485 VSS.n5085 VSS.n5081 0.0095
R11486 VSS.n3756 VSS.n3755 0.00939535
R11487 VSS.n4575 VSS.n4574 0.00931119
R11488 VSS.n4584 VSS.n4583 0.00931119
R11489 VSS.n3552 VSS.n3551 0.00926454
R11490 VSS.n5771 VSS.n5770 0.00925
R11491 VSS.n4940 VSS.n4939 0.00925
R11492 VSS.n5092 VSS.n5091 0.00902632
R11493 VSS.n2803 VSS.n2475 0.00900291
R11494 VSS.n6072 VSS.n6071 0.00899057
R11495 VSS.n3680 VSS.n3679 0.00887209
R11496 VSS.n7806 VSS.n7802 0.00883333
R11497 VSS.n7128 VSS.n7125 0.00875688
R11498 VSS.n680 VSS.n679 0.00868182
R11499 VSS.n4549 VSS.n4548 0.00868182
R11500 VSS.n4569 VSS.n4564 0.00868182
R11501 VSS.n1489 VSS.n1488 0.00868182
R11502 VSS.n2258 VSS.n2247 0.00862709
R11503 VSS.n2272 VSS.n2269 0.00862709
R11504 VSS.n2414 VSS.n2413 0.00862709
R11505 VSS.n2393 VSS.n2392 0.00862709
R11506 VSS.n4008 VSS.n4007 0.0086106
R11507 VSS.n2782 VSS.n2781 0.00861047
R11508 VSS.n5759 VSS.n5756 0.00855263
R11509 VSS.n3031 VSS.n3030 0.00855063
R11510 VSS.n4156 VSS.n4155 0.00854878
R11511 VSS.n3454 VSS.n3453 0.00847965
R11512 VSS.n3740 VSS.n3739 0.00840698
R11513 VSS.n2701 VSS.n2700 0.00838571
R11514 VSS.n1774 VSS.n1773 0.00836872
R11515 VSS.n1877 VSS.n1876 0.00836872
R11516 VSS.n1764 VSS.n1763 0.00836872
R11517 VSS.n610 VSS.n607 0.00836713
R11518 VSS.n676 VSS.n673 0.00836713
R11519 VSS.n1512 VSS.n1509 0.00836713
R11520 VSS.n1569 VSS.n1566 0.00836713
R11521 VSS.n2517 VSS.n2485 0.00834884
R11522 VSS.n3923 VSS.n3922 0.00833217
R11523 VSS.n4992 VSS.n4989 0.00832609
R11524 VSS.n2737 VSS.n2563 0.0082907
R11525 VSS.n3644 VSS.n3643 0.00808721
R11526 VSS.n3393 VSS.n3392 0.00808721
R11527 VSS.n4393 VSS.n4392 0.00805245
R11528 VSS.n4384 VSS.n4383 0.00805245
R11529 VSS.n4054 VSS.n4053 0.0080419
R11530 VSS.n2230 VSS.n2229 0.00802508
R11531 VSS.n1368 VSS.n1365 0.008
R11532 VSS.n3796 VSS.n3795 0.00797826
R11533 VSS.n1253 VSS.n1250 0.00795562
R11534 VSS.n2110 VSS.n2109 0.00794828
R11535 VSS.n202 VSS.n201 0.00793119
R11536 VSS.n200 VSS.n199 0.00793119
R11537 VSS.n162 VSS.n161 0.00784694
R11538 VSS.n2501 VSS.n2499 0.00782558
R11539 VSS.n154 VSS.n151 0.00781707
R11540 VSS.n4110 VSS.n4104 0.0077905
R11541 VSS.n4068 VSS.n4067 0.0077905
R11542 VSS.n4058 VSS.n4057 0.0077905
R11543 VSS.n171 VSS.n170 0.00773214
R11544 VSS.n3007 VSS.n3006 0.00772408
R11545 VSS.n3447 VSS.n3446 0.00769477
R11546 VSS.n6178 VSS.n6175 0.00760526
R11547 VSS.n2406 VSS.n2405 0.00757358
R11548 VSS.n1592 VSS.n1591 0.00757142
R11549 VSS.n4091 VSS.n4086 0.00753911
R11550 VSS.n4080 VSS.n4079 0.00753911
R11551 VSS.n2867 VSS.n2866 0.00748113
R11552 VSS.n1588 VSS.n1587 0.00743371
R11553 VSS VSS.n4397 0.00742308
R11554 VSS.n4392 VSS.n4385 0.00742308
R11555 VSS.n689 VSS.n688 0.00735714
R11556 VSS.n5864 VSS.n5863 0.00734783
R11557 VSS.n1832 VSS.n1831 0.00734332
R11558 VSS.n1862 VSS.n1861 0.00734332
R11559 VSS.n2359 VSS.n2358 0.0073277
R11560 VSS.n3716 VSS.n3715 0.00730233
R11561 VSS.n4064 VSS.n4063 0.00728771
R11562 VSS.n1968 VSS.n1967 0.00726364
R11563 VSS.n1830 VSS.n1829 0.00713594
R11564 VSS.n1860 VSS.n1859 0.00713594
R11565 VSS.n69 VSS.n68 0.00708537
R11566 VSS.n4718 VSS.n4716 0.00708537
R11567 VSS.n3086 VSS.n3085 0.0070407
R11568 VSS.n2509 VSS.n2507 0.0070407
R11569 VSS.n4126 VSS.n4124 0.00703631
R11570 VSS.n4076 VSS.n4075 0.00703631
R11571 VSS.n4072 VSS.n4071 0.00703631
R11572 VSS.n3953 VSS.n3944 0.00701869
R11573 VSS.n2063 VSS.n2062 0.00701724
R11574 VSS.n5776 VSS.n5775 0.00689344
R11575 VSS.n2107 VSS.n2106 0.00686207
R11576 VSS.n2161 VSS.n2159 0.00682107
R11577 VSS.n4868 VSS.n4855 0.00681579
R11578 VSS.n3929 VSS.n3928 0.00680841
R11579 VSS.n4550 VSS.n4535 0.00679371
R11580 VSS.n4548 VSS.n4536 0.00679371
R11581 VSS.n4563 VSS.n595 0.00679371
R11582 VSS.n4570 VSS.n4569 0.00679371
R11583 VSS.n4119 VSS.n4113 0.00678492
R11584 VSS.n1870 VSS.n1869 0.00678492
R11585 VSS.n3074 VSS.n3073 0.00677907
R11586 VSS.n3523 VSS.n3522 0.00668497
R11587 VSS.n2714 VSS.n2584 0.00667143
R11588 VSS.n2995 VSS.n2173 0.00667057
R11589 VSS.n2862 VSS.n2861 0.00667057
R11590 VSS.n6976 VSS 0.00664458
R11591 VSS.n2113 VSS.n2112 0.00655172
R11592 VSS.n1413 VSS.n1412 0.00655042
R11593 VSS.n6534 VSS.n6531 0.00655042
R11594 VSS.n7100 VSS.n7074 0.00655042
R11595 VSS.n5343 VSS.n5342 0.00655042
R11596 VSS.n6662 VSS.n6661 0.00655042
R11597 VSS.n1047 VSS.n1044 0.00655042
R11598 VSS VSS.n6714 0.00652231
R11599 VSS.n1779 VSS.n1778 0.00651383
R11600 VSS.n1593 VSS.n1592 0.0065
R11601 VSS.n579 VSS.n75 0.0064434
R11602 VSS.n563 VSS.n562 0.0064434
R11603 VSS.n528 VSS.n325 0.0064434
R11604 VSS.n4701 VSS.n4700 0.0064434
R11605 VSS.n4943 VSS.n4942 0.00640164
R11606 VSS.n2157 VSS.n2156 0.00636957
R11607 VSS.n1865 VSS.n1804 0.00630645
R11608 VSS.n1863 VSS.n1828 0.00630645
R11609 VSS.n198 VSS.n197 0.00627982
R11610 VSS.n2523 VSS.n2522 0.00625581
R11611 VSS.n3773 VSS.n3772 0.00625581
R11612 VSS.n2124 VSS.n2080 0.00624138
R11613 VSS.n2076 VSS.n2070 0.00624138
R11614 VSS.n2066 VSS.n2060 0.00624138
R11615 VSS.n2056 VSS.n2048 0.00624138
R11616 VSS.n2034 VSS.n2033 0.00624138
R11617 VSS.n2013 VSS.n2008 0.00624138
R11618 VSS.n6624 VSS.n6620 0.00622751
R11619 VSS.n7622 VSS.n7620 0.00622751
R11620 VSS.n1486 VSS.n718 0.00622751
R11621 VSS.n2974 VSS.n2198 0.00618562
R11622 VSS.n1787 VSS.n1786 0.00617757
R11623 VSS.n3947 VSS.n3946 0.00617757
R11624 VSS.n3970 VSS.n3969 0.00617757
R11625 VSS.n3952 VSS.n3951 0.00617757
R11626 VSS.n3917 VSS.n3907 0.00617757
R11627 VSS.n3484 VSS.n3483 0.00616474
R11628 VSS.n4583 VSS.n4576 0.00616434
R11629 VSS.n766 VSS 0.006125
R11630 VSS.n188 VSS 0.006125
R11631 VSS VSS.n6410 0.006125
R11632 VSS VSS.n7175 0.006125
R11633 VSS.n6944 VSS 0.006125
R11634 VSS.n6742 VSS 0.006125
R11635 VSS.n4596 VSS 0.006125
R11636 VSS VSS.n942 0.006125
R11637 VSS.n2319 VSS.n2313 0.00610386
R11638 VSS.n2077 VSS.n2076 0.00608621
R11639 VSS.n2067 VSS.n2066 0.00608621
R11640 VSS.n2059 VSS.n2058 0.00608621
R11641 VSS.n2057 VSS.n2056 0.00608621
R11642 VSS.n2014 VSS.n2013 0.00608621
R11643 VSS.n3020 VSS.n2138 0.00606856
R11644 VSS.n3015 VSS.n3014 0.00606856
R11645 VSS.n3010 VSS.n2152 0.00606856
R11646 VSS.n3003 VSS.n2164 0.00606856
R11647 VSS.n2199 VSS.n2186 0.00606856
R11648 VSS.n2948 VSS.n2238 0.00606856
R11649 VSS.n2938 VSS.n2245 0.00606856
R11650 VSS.n2919 VSS.n2918 0.00606856
R11651 VSS.n2879 VSS.n2331 0.00606856
R11652 VSS.n2869 VSS.n2361 0.00606856
R11653 VSS.n2864 VSS.n2863 0.00606856
R11654 VSS.n2814 VSS.n2468 0.00606856
R11655 VSS.n3822 VSS.n3821 0.00606522
R11656 VSS.n3699 VSS.n3698 0.00599419
R11657 VSS.n3203 VSS.n3202 0.00599419
R11658 VSS.n7430 VSS.n7428 0.0059878
R11659 VSS.n5753 VSS.n5752 0.00596961
R11660 VSS.n3938 VSS.n3937 0.00596729
R11661 VSS.n3939 VSS.n3935 0.00596729
R11662 VSS.n3901 VSS.n3893 0.00596729
R11663 VSS.n2053 VSS.n2052 0.00593103
R11664 VSS.n3026 VSS.n2138 0.00591806
R11665 VSS.n3015 VSS.n2145 0.00591806
R11666 VSS.n3011 VSS.n3010 0.00591806
R11667 VSS.n2167 VSS.n2166 0.00591806
R11668 VSS.n3003 VSS.n2163 0.00591806
R11669 VSS.n2948 VSS.n2237 0.00591806
R11670 VSS.n2944 VSS.n2245 0.00591806
R11671 VSS.n2933 VSS.n2252 0.00591806
R11672 VSS.n2880 VSS.n2879 0.00591806
R11673 VSS.n2875 VSS.n2361 0.00591806
R11674 VSS.n2864 VSS.n2368 0.00591806
R11675 VSS.n2847 VSS.n2387 0.00591806
R11676 VSS.n2441 VSS.n2434 0.0059088
R11677 VSS.n1842 VSS.n1841 0.0058917
R11678 VSS.n1854 VSS.n1853 0.0058917
R11679 VSS.n4082 VSS.n4081 0.00588013
R11680 VSS.n3078 VSS.n3077 0.00586337
R11681 VSS.n635 VSS.n599 0.00584965
R11682 VSS.n3605 VSS.n3604 0.00584884
R11683 VSS.n7548 VSS.n7547 0.00579412
R11684 VSS.n2117 VSS.n2116 0.00577586
R11685 VSS.n2114 VSS.n2113 0.00577586
R11686 VSS.n2111 VSS.n2110 0.00577586
R11687 VSS.n2108 VSS.n2107 0.00577586
R11688 VSS.n2100 VSS.n2099 0.00577586
R11689 VSS.n2123 VSS.n2122 0.00577586
R11690 VSS.n2075 VSS.n2074 0.00577586
R11691 VSS.n2065 VSS.n2064 0.00577586
R11692 VSS.n2055 VSS.n2054 0.00577586
R11693 VSS.n1997 VSS.n1996 0.00577586
R11694 VSS.n2997 VSS.n2171 0.00576756
R11695 VSS.n2374 VSS.n2371 0.00576756
R11696 VSS.n3018 VSS.n3017 0.00571739
R11697 VSS.n1838 VSS.n1837 0.00568433
R11698 VSS.n1850 VSS.n1849 0.00568433
R11699 VSS.n2115 VSS.n2114 0.00562069
R11700 VSS.n2112 VSS.n2111 0.00562069
R11701 VSS.n2109 VSS.n2108 0.00562069
R11702 VSS.n2010 VSS.n2009 0.00562069
R11703 VSS.n2073 VSS.n2072 0.00562069
R11704 VSS.n3024 VSS.n3023 0.00561706
R11705 VSS.n2156 VSS.n2155 0.00561706
R11706 VSS.n3007 VSS.n2158 0.00561706
R11707 VSS.n2173 VSS.n2160 0.00561706
R11708 VSS.n2204 VSS.n2183 0.00561706
R11709 VSS.n3022 VSS.n2139 0.00561706
R11710 VSS.n2149 VSS.n2147 0.00561706
R11711 VSS.n3009 VSS.n3008 0.00561706
R11712 VSS.n3004 VSS.n2162 0.00561706
R11713 VSS.n2203 VSS.n2184 0.00561706
R11714 VSS.n2294 VSS.n2293 0.00561706
R11715 VSS.n2942 VSS.n2941 0.00561706
R11716 VSS.n2289 VSS.n2288 0.00561706
R11717 VSS.n2904 VSS.n2282 0.00561706
R11718 VSS.n2940 VSS.n2246 0.00561706
R11719 VSS.n2270 VSS.n2268 0.00561706
R11720 VSS.n2873 VSS.n2872 0.00561706
R11721 VSS.n2405 VSS.n2404 0.00561706
R11722 VSS.n2871 VSS.n2362 0.00561706
R11723 VSS.n2372 VSS.n2370 0.00561706
R11724 VSS.n3069 VSS.n3068 0.00560174
R11725 VSS.n3978 VSS.n3977 0.00554673
R11726 VSS.n1539 VSS.n1528 0.00553496
R11727 VSS.n1546 VSS.n1545 0.00553496
R11728 VSS.n1605 VSS.n1598 0.00553496
R11729 VSS.n4036 VSS.n4035 0.00552326
R11730 VSS.n7844 VSS.n7836 0.0055
R11731 VSS.n4933 VSS.n4932 0.00547238
R11732 VSS.n3867 VSS.n3866 0.00547093
R11733 VSS.n2155 VSS.n2141 0.00546656
R11734 VSS.n2158 VSS.n2157 0.00546656
R11735 VSS.n3006 VSS.n2160 0.00546656
R11736 VSS.n2951 VSS.n2234 0.00546656
R11737 VSS.n2147 VSS.n2146 0.00546656
R11738 VSS.n3013 VSS.n3012 0.00546656
R11739 VSS.n3009 VSS.n2150 0.00546656
R11740 VSS.n3005 VSS.n3004 0.00546656
R11741 VSS.n2950 VSS.n2949 0.00546656
R11742 VSS.n2293 VSS.n2292 0.00546656
R11743 VSS.n2257 VSS.n2248 0.00546656
R11744 VSS.n2291 VSS.n2290 0.00546656
R11745 VSS.n2291 VSS.n2280 0.00546656
R11746 VSS.n2905 VSS.n2904 0.00546656
R11747 VSS.n2353 VSS.n2332 0.00546656
R11748 VSS.n2254 VSS.n2253 0.00546656
R11749 VSS.n2355 VSS.n2329 0.00546656
R11750 VSS.n2404 VSS.n2364 0.00546656
R11751 VSS.n2850 VSS.n2384 0.00546656
R11752 VSS.n2370 VSS.n2369 0.00546656
R11753 VSS.n2849 VSS.n2848 0.00546656
R11754 VSS.n1963 VSS.n1962 0.00546429
R11755 VSS.n2640 VSS.n2633 0.00541429
R11756 VSS.n4787 VSS.n4783 0.0053913
R11757 VSS.n3149 VSS.n3148 0.00538372
R11758 VSS.n2585 VSS.n2581 0.00534716
R11759 VSS.n2703 VSS.n2586 0.00534716
R11760 VSS.n3696 VSS.n3695 0.00534012
R11761 VSS.n3732 VSS.n3731 0.00534012
R11762 VSS.n3713 VSS.n3712 0.00534012
R11763 VSS.n3529 VSS.n3525 0.00534012
R11764 VSS.n3439 VSS.n3432 0.00534012
R11765 VSS.n3404 VSS.n3370 0.00534012
R11766 VSS.n3362 VSS.n3358 0.00534012
R11767 VSS.n3325 VSS.n3324 0.00534012
R11768 VSS.n3285 VSS.n3284 0.00534012
R11769 VSS.n3244 VSS.n3243 0.00534012
R11770 VSS.n3223 VSS.n3222 0.00534012
R11771 VSS.n3206 VSS.n3200 0.00534012
R11772 VSS.n3193 VSS.n3192 0.00534012
R11773 VSS.n3159 VSS.n3158 0.00534012
R11774 VSS.n3106 VSS.n3105 0.00534012
R11775 VSS.n2804 VSS.n2470 0.00534012
R11776 VSS.n2785 VSS.n2493 0.00534012
R11777 VSS.n2765 VSS.n2529 0.00534012
R11778 VSS.n2728 VSS.n2564 0.00534012
R11779 VSS.n3793 VSS.n3792 0.00534012
R11780 VSS.n3911 VSS.n3910 0.00533645
R11781 VSS.n3916 VSS.n3915 0.00533645
R11782 VSS.n3983 VSS.n3982 0.00533645
R11783 VSS.n3963 VSS.n3962 0.00533645
R11784 VSS.n194 VSS.n193 0.00532143
R11785 VSS.n6489 VSS 0.00532143
R11786 VSS.n7234 VSS 0.00532143
R11787 VSS.n7610 VSS 0.00532143
R11788 VSS VSS.n6635 0.00532143
R11789 VSS VSS.n139 0.00532143
R11790 VSS VSS.n4480 0.00532143
R11791 VSS VSS.n4518 0.00532143
R11792 VSS VSS.n1004 0.00532143
R11793 VSS.n1965 VSS.n1964 0.00527273
R11794 VSS.n2725 VSS.n2574 0.00521616
R11795 VSS.n2711 VSS.n2586 0.00521616
R11796 VSS.n3610 VSS.n3609 0.0052093
R11797 VSS.n3615 VSS.n3614 0.0052093
R11798 VSS.n3737 VSS.n3618 0.0052093
R11799 VSS.n3714 VSS.n3713 0.0052093
R11800 VSS.n3584 VSS.n3533 0.0052093
R11801 VSS.n3584 VSS.n3537 0.0052093
R11802 VSS.n3439 VSS.n3428 0.0052093
R11803 VSS.n3404 VSS.n3366 0.0052093
R11804 VSS.n3270 VSS.n3269 0.0052093
R11805 VSS.n3223 VSS.n3211 0.0052093
R11806 VSS.n3199 VSS.n3198 0.0052093
R11807 VSS.n3106 VSS.n3063 0.0052093
R11808 VSS.n2810 VSS.n2470 0.0052093
R11809 VSS.n2477 VSS.n2476 0.0052093
R11810 VSS.n2734 VSS.n2564 0.0052093
R11811 VSS.n1907 VSS.n1902 0.0052093
R11812 VSS.n3855 VSS.n3841 0.0052093
R11813 VSS.n3793 VSS.n3747 0.0052093
R11814 VSS.n2908 VSS.n2278 0.00516555
R11815 VSS.n2315 VSS.n2295 0.00516555
R11816 VSS.n2899 VSS.n2898 0.00516555
R11817 VSS.n3898 VSS.n3897 0.00512617
R11818 VSS.n3899 VSS.n3896 0.00512617
R11819 VSS.n3967 VSS.n3966 0.00512617
R11820 VSS.n5906 VSS.n5905 0.00511538
R11821 VSS.n4750 VSS.n4749 0.00511538
R11822 VSS.n215 VSS.n162 0.00509184
R11823 VSS.n3376 VSS.n3375 0.00507849
R11824 VSS.n3764 VSS.n3763 0.00507849
R11825 VSS.n1794 VSS.n1793 0.00506221
R11826 VSS.n1813 VSS.n1812 0.00506221
R11827 VSS.n1823 VSS.n1822 0.00506221
R11828 VSS.n2277 VSS.n2271 0.00501505
R11829 VSS.n2903 VSS.n2281 0.00501505
R11830 VSS.n2915 VSS.n2914 0.00501505
R11831 VSS.n2047 VSS.n2046 0.005
R11832 VSS.n2591 VSS.n2589 0.00495415
R11833 VSS.n2707 VSS.n2706 0.00495415
R11834 VSS.n2590 VSS.n2579 0.00495415
R11835 VSS.n2705 VSS.n2588 0.00495415
R11836 VSS.n3669 VSS.n3668 0.00494767
R11837 VSS.n3690 VSS.n3689 0.00494767
R11838 VSS.n3681 VSS.n3680 0.00494767
R11839 VSS.n3678 VSS.n3677 0.00494767
R11840 VSS.n3626 VSS.n3625 0.00494767
R11841 VSS.n3660 VSS.n3659 0.00494767
R11842 VSS.n3646 VSS.n3645 0.00494767
R11843 VSS.n3641 VSS.n3640 0.00494767
R11844 VSS.n3612 VSS.n3611 0.00494767
R11845 VSS.n3718 VSS.n3717 0.00494767
R11846 VSS.n3577 VSS.n3575 0.00494767
R11847 VSS.n3573 VSS.n3572 0.00494767
R11848 VSS.n3550 VSS.n3549 0.00494767
R11849 VSS.n3583 VSS.n3582 0.00494767
R11850 VSS.n3528 VSS.n3527 0.00494767
R11851 VSS.n3438 VSS.n3437 0.00494767
R11852 VSS.n3397 VSS.n3396 0.00494767
R11853 VSS.n3394 VSS.n3393 0.00494767
R11854 VSS.n3385 VSS.n3384 0.00494767
R11855 VSS.n3230 VSS.n3229 0.00494767
R11856 VSS.n3233 VSS.n3232 0.00494767
R11857 VSS.n3403 VSS.n3402 0.00494767
R11858 VSS.n3361 VSS.n3360 0.00494767
R11859 VSS.n3320 VSS.n3319 0.00494767
R11860 VSS.n3280 VSS.n3279 0.00494767
R11861 VSS.n3265 VSS.n3264 0.00494767
R11862 VSS.n3068 VSS.n3067 0.00494767
R11863 VSS.n3073 VSS.n3072 0.00494767
R11864 VSS.n3077 VSS.n3076 0.00494767
R11865 VSS.n3088 VSS.n3087 0.00494767
R11866 VSS.n3218 VSS.n3217 0.00494767
R11867 VSS.n3205 VSS.n3204 0.00494767
R11868 VSS.n3189 VSS.n3188 0.00494767
R11869 VSS.n3156 VSS.n3155 0.00494767
R11870 VSS.n2808 VSS.n2807 0.00494767
R11871 VSS.n2794 VSS.n2483 0.00494767
R11872 VSS.n2782 VSS.n2498 0.00494767
R11873 VSS.n2767 VSS.n2524 0.00494767
R11874 VSS.n2806 VSS.n2471 0.00494767
R11875 VSS.n2784 VSS.n2783 0.00494767
R11876 VSS.n2766 VSS.n2526 0.00494767
R11877 VSS.n3766 VSS.n3765 0.00494767
R11878 VSS.n3775 VSS.n3774 0.00494767
R11879 VSS VSS.n728 0.00490559
R11880 VSS.n613 VSS.n610 0.00490559
R11881 VSS.n619 VSS.n616 0.00490559
R11882 VSS.n625 VSS.n622 0.00490559
R11883 VSS.n629 VSS.n628 0.00490559
R11884 VSS.n653 VSS.n650 0.00490559
R11885 VSS.n666 VSS.n663 0.00490559
R11886 VSS.n679 VSS.n676 0.00490559
R11887 VSS VSS.n5501 0.00490559
R11888 VSS VSS.n5464 0.00490559
R11889 VSS VSS.n5458 0.00490559
R11890 VSS VSS.n5576 0.00490559
R11891 VSS.n6445 VSS 0.00490559
R11892 VSS VSS.n7095 0.00490559
R11893 VSS VSS.n5346 0.00490559
R11894 VSS VSS.n6665 0.00490559
R11895 VSS.n1515 VSS.n1512 0.00490559
R11896 VSS.n1521 VSS.n1518 0.00490559
R11897 VSS.n1527 VSS.n1524 0.00490559
R11898 VSS.n1559 VSS.n1556 0.00490559
R11899 VSS.n1584 VSS.n1581 0.00490559
R11900 VSS.n1578 VSS.n1575 0.00490559
R11901 VSS.n1572 VSS.n1569 0.00490559
R11902 VSS VSS.n4541 0.00490559
R11903 VSS.n4402 VSS 0.00490559
R11904 VSS.n972 VSS 0.00490559
R11905 VSS.n226 VSS.n225 0.00489024
R11906 VSS.n3000 VSS.n2999 0.00486455
R11907 VSS.n1596 VSS.n1595 0.00486421
R11908 VSS.n1791 VSS.n1781 0.00485484
R11909 VSS.n1798 VSS.n1797 0.00485484
R11910 VSS.n1811 VSS.n1810 0.00485484
R11911 VSS.n1821 VSS.n1820 0.00485484
R11912 VSS.n2708 VSS.n2707 0.00482314
R11913 VSS.n2709 VSS.n2588 0.00482314
R11914 VSS.n3700 VSS.n3670 0.00481686
R11915 VSS.n3679 VSS.n3678 0.00481686
R11916 VSS.n3701 VSS.n3629 0.00481686
R11917 VSS.n3642 VSS.n3641 0.00481686
R11918 VSS.n3574 VSS.n3573 0.00481686
R11919 VSS.n3551 VSS.n3550 0.00481686
R11920 VSS.n3548 VSS.n3547 0.00481686
R11921 VSS.n3438 VSS.n3433 0.00481686
R11922 VSS.n3395 VSS.n3394 0.00481686
R11923 VSS.n3384 VSS.n3383 0.00481686
R11924 VSS.n3383 VSS.n3382 0.00481686
R11925 VSS.n3232 VSS.n3231 0.00481686
R11926 VSS.n3237 VSS.n3234 0.00481686
R11927 VSS.n3067 VSS.n3066 0.00481686
R11928 VSS.n3072 VSS.n3069 0.00481686
R11929 VSS.n3076 VSS.n3074 0.00481686
R11930 VSS.n3102 VSS.n3101 0.00481686
R11931 VSS.n3218 VSS.n3213 0.00481686
R11932 VSS.n3216 VSS.n3215 0.00481686
R11933 VSS.n3104 VSS.n3065 0.00481686
R11934 VSS.n2483 VSS.n2473 0.00481686
R11935 VSS.n2793 VSS.n2792 0.00481686
R11936 VSS.n2731 VSS.n2730 0.00481686
R11937 VSS.n2481 VSS.n2480 0.00481686
R11938 VSS.n2796 VSS.n2481 0.00481686
R11939 VSS.n2732 VSS.n2566 0.00481686
R11940 VSS.n3765 VSS.n3764 0.00481686
R11941 VSS.n3774 VSS.n3773 0.00481686
R11942 VSS.n3789 VSS.n3788 0.00481686
R11943 VSS.n1906 VSS.n1905 0.00481686
R11944 VSS.n3791 VSS.n3749 0.00481686
R11945 VSS.n3807 VSS.n3806 0.00481686
R11946 VSS.n3040 VSS.n3039 0.0048038
R11947 VSS.n3994 VSS.n3992 0.00476036
R11948 VSS.n4022 VSS.n4021 0.00476036
R11949 VSS.n4025 VSS.n4024 0.00476036
R11950 VSS.n2762 VSS.n2542 0.00474419
R11951 VSS.n2926 VSS.n2259 0.00471405
R11952 VSS.n2911 VSS.n2910 0.00471405
R11953 VSS.n2069 VSS.n2068 0.00468966
R11954 VSS.n3546 VSS.n3545 0.00468605
R11955 VSS.n3411 VSS.n3410 0.00468605
R11956 VSS.n3414 VSS.n3413 0.00468605
R11957 VSS.n3381 VSS.n3380 0.00468605
R11958 VSS.n2791 VSS.n2486 0.00468605
R11959 VSS.n3854 VSS.n3853 0.00468605
R11960 VSS.n3861 VSS.n3860 0.00468605
R11961 VSS.n3818 VSS.n3812 0.00468605
R11962 VSS.n2151 VSS.n2148 0.00456355
R11963 VSS.n2288 VSS.n2287 0.00456355
R11964 VSS.n2902 VSS.n2297 0.00456355
R11965 VSS.n1538 VSS.n1534 0.00456316
R11966 VSS.n2936 VSS.n2935 0.00455797
R11967 VSS.n3735 VSS.n3734 0.00455523
R11968 VSS.n4101 VSS.n4098 0.0045168
R11969 VSS.n3059 VSS.n3058 0.00444937
R11970 VSS.n2718 VSS.n2580 0.00443013
R11971 VSS.n3238 VSS.n3237 0.00442442
R11972 VSS.n2798 VSS.n2477 0.00442442
R11973 VSS.n3786 VSS.n3785 0.00442442
R11974 VSS.n3802 VSS.n3801 0.00442442
R11975 VSS.n2651 VSS.n2648 0.00429913
R11976 VSS.n2681 VSS.n2616 0.00429913
R11977 VSS.n3676 VSS.n3675 0.0042936
R11978 VSS.n3634 VSS.n3633 0.0042936
R11979 VSS.n3706 VSS.n3705 0.0042936
R11980 VSS.n3373 VSS.n3372 0.0042936
R11981 VSS.n3392 VSS.n3391 0.0042936
R11982 VSS.n3390 VSS.n3389 0.0042936
R11983 VSS.n3240 VSS.n3239 0.0042936
R11984 VSS.n3191 VSS.n3190 0.0042936
R11985 VSS.n2522 VSS.n2518 0.0042936
R11986 VSS.n2781 VSS.n2500 0.0042936
R11987 VSS.n2521 VSS.n2519 0.0042936
R11988 VSS.n2520 VSS.n2504 0.0042936
R11989 VSS.n2790 VSS.n2488 0.0042936
R11990 VSS.n2777 VSS.n2505 0.0042936
R11991 VSS.n3763 VSS.n3762 0.0042936
R11992 VSS.n3784 VSS.n3783 0.0042936
R11993 VSS.n1904 VSS.n1903 0.0042936
R11994 VSS.n3817 VSS.n3816 0.0042936
R11995 VSS.n3855 VSS.n3847 0.0042936
R11996 VSS.n2802 VSS.n2801 0.00427907
R11997 VSS.n636 VSS.n635 0.00427622
R11998 VSS.n660 VSS.n657 0.00427622
R11999 VSS.n2925 VSS.n2261 0.00426254
R12000 VSS.n4111 VSS.n4102 0.00418349
R12001 VSS.n3667 VSS.n3666 0.00416279
R12002 VSS.n3623 VSS.n3622 0.00416279
R12003 VSS.n3833 VSS.n3832 0.00416279
R12004 VSS.n1689 VSS.n1688 0.00415854
R12005 VSS.n4301 VSS.n4300 0.00415854
R12006 VSS.n4919 VSS.n4914 0.00414865
R12007 VSS.n2285 VSS.n2268 0.00411204
R12008 VSS.n2855 VSS.n2854 0.00411204
R12009 VSS.n3396 VSS.n3395 0.00403198
R12010 VSS.n3318 VSS.n3317 0.00403198
R12011 VSS.n3252 VSS.n3251 0.00403198
R12012 VSS.n3221 VSS.n3220 0.00403198
R12013 VSS.n2792 VSS.n2484 0.00403198
R12014 VSS.n3758 VSS.n3757 0.00403198
R12015 VSS.n3768 VSS.n3767 0.00403198
R12016 VSS.n3770 VSS.n3769 0.00403198
R12017 VSS.n3772 VSS.n3771 0.00403198
R12018 VSS.n2275 VSS.n2274 0.00397826
R12019 VSS.n4557 VSS.n4556 0.00397013
R12020 VSS.n2856 VSS.n2375 0.00396154
R12021 VSS.n5908 VSS.n5906 0.00396154
R12022 VSS.n2683 VSS.n2682 0.00390611
R12023 VSS.n2634 VSS.n2613 0.00390611
R12024 VSS.n3637 VSS.n3636 0.00390116
R12025 VSS.n3631 VSS.n3630 0.00390116
R12026 VSS.n3709 VSS.n3708 0.00390116
R12027 VSS.n3703 VSS.n3702 0.00390116
R12028 VSS.n3349 VSS.n3348 0.00390116
R12029 VSS.n3345 VSS.n3344 0.00390116
R12030 VSS.n2498 VSS.n2497 0.00390116
R12031 VSS.n2780 VSS.n2779 0.00390116
R12032 VSS.n2508 VSS.n2503 0.00390116
R12033 VSS.n2527 VSS.n2513 0.00390116
R12034 VSS.n1883 VSS.n1882 0.00390116
R12035 VSS.n1889 VSS.n1888 0.00390116
R12036 VSS.n2394 VSS.n2390 0.00389623
R12037 VSS.n3997 VSS.n3996 0.00381797
R12038 VSS.n3999 VSS.n3998 0.00381797
R12039 VSS.n4018 VSS.n4017 0.00381797
R12040 VSS.n4020 VSS.n4019 0.00381797
R12041 VSS.n2924 VSS.n2263 0.00381104
R12042 VSS.n2888 VSS.n2325 0.00381104
R12043 VSS.n3697 VSS.n3696 0.00377035
R12044 VSS.n3692 VSS.n3691 0.00377035
R12045 VSS.n3688 VSS.n3687 0.00377035
R12046 VSS.n3686 VSS.n3685 0.00377035
R12047 VSS.n3683 VSS.n3682 0.00377035
R12048 VSS.n3663 VSS.n3662 0.00377035
R12049 VSS.n3653 VSS.n3652 0.00377035
R12050 VSS.n3780 VSS.n3779 0.00377035
R12051 VSS.n3828 VSS.n3827 0.00377035
R12052 VSS.n4551 VSS.n696 0.00373363
R12053 VSS.n5727 VSS.n5712 0.00371429
R12054 VSS.n3442 VSS.n3441 0.00367919
R12055 VSS.n3930 VSS.n3924 0.00367016
R12056 VSS.n3957 VSS.n3956 0.00367016
R12057 VSS.n6302 VSS.n5388 0.00366159
R12058 VSS.n2928 VSS.n2257 0.00366054
R12059 VSS.n2920 VSS.n2919 0.00366054
R12060 VSS.n2890 VSS.n2321 0.00366054
R12061 VSS.n2411 VSS.n2383 0.00366054
R12062 VSS.n2401 VSS.n2384 0.00366054
R12063 VSS.n2381 VSS.n2379 0.00366054
R12064 VSS.n4415 VSS.n4409 0.00364685
R12065 VSS.n4405 VSS.n4402 0.00364685
R12066 VSS.n2722 VSS.n2577 0.0036441
R12067 VSS.n2721 VSS.n2720 0.0036441
R12068 VSS.n3379 VSS.n3378 0.00363953
R12069 VSS.n3257 VSS.n3256 0.00363953
R12070 VSS.n2791 VSS.n2487 0.00363953
R12071 VSS.n3778 VSS.n3777 0.00363953
R12072 VSS.n1920 VSS.n1919 0.00363953
R12073 VSS.n3869 VSS.n3868 0.00363953
R12074 VSS.n3863 VSS.n3862 0.00363953
R12075 VSS.n4348 VSS.n4347 0.00360345
R12076 VSS.n4034 VSS.n4033 0.00356977
R12077 VSS.n3596 VSS.n3595 0.00352326
R12078 VSS.n2927 VSS.n2926 0.00351003
R12079 VSS.n2410 VSS.n2409 0.00351003
R12080 VSS.n2408 VSS.n2378 0.00351003
R12081 VSS.n2834 VSS.n2420 0.00351003
R12082 VSS.n2823 VSS.n2440 0.00351003
R12083 VSS.n3677 VSS.n3676 0.00350872
R12084 VSS.n3725 VSS.n3724 0.00350872
R12085 VSS.n3553 VSS.n3552 0.00350872
R12086 VSS.n2769 VSS.n2768 0.00350872
R12087 VSS.n2784 VSS.n2494 0.00350872
R12088 VSS.n2770 VSS.n2515 0.00350872
R12089 VSS.n1901 VSS.n1900 0.00350872
R12090 VSS.n6580 VSS.n6388 0.0035
R12091 VSS.n6935 VSS.n6932 0.0035
R12092 VSS.n4037 VSS.n4036 0.00347674
R12093 VSS.n72 VSS.n69 0.0034717
R12094 VSS.n559 VSS.n556 0.0034717
R12095 VSS.n318 VSS.n312 0.0034717
R12096 VSS.n4664 VSS.n4663 0.0034717
R12097 VSS.n4697 VSS.n4687 0.0034717
R12098 VSS.n2043 VSS.n2042 0.00344828
R12099 VSS.n2510 VSS.n2506 0.00340698
R12100 VSS.n3656 VSS.n3655 0.00337791
R12101 VSS.n3648 VSS.n3647 0.00337791
R12102 VSS.n3728 VSS.n3727 0.00337791
R12103 VSS.n3720 VSS.n3719 0.00337791
R12104 VSS.n2991 VSS.n2176 0.00335953
R12105 VSS.n2351 VSS.n2350 0.00335953
R12106 VSS.n2349 VSS.n2324 0.00335953
R12107 VSS.n2931 VSS.n2255 0.00335953
R12108 VSS.n6932 VSS.n6931 0.00333019
R12109 VSS.n6925 VSS.n6924 0.00333019
R12110 VSS.n6913 VSS.n6618 0.00333019
R12111 VSS.n6939 VSS.n6938 0.00333019
R12112 VSS.n3902 VSS.n3890 0.0032972
R12113 VSS.n3921 VSS.n3920 0.0032972
R12114 VSS.n4044 VSS.n4043 0.0032907
R12115 VSS.n4038 VSS.n4037 0.0032907
R12116 VSS.n3995 VSS.n3994 0.00324751
R12117 VSS.n4026 VSS.n4025 0.00324751
R12118 VSS.n4023 VSS.n4022 0.00324751
R12119 VSS.n3401 VSS.n3400 0.00324709
R12120 VSS.n3323 VSS.n3322 0.00324709
R12121 VSS.n2790 VSS.n2489 0.00324709
R12122 VSS.n1915 VSS.n1914 0.00324709
R12123 VSS.n1959 VSS.n1958 0.00322727
R12124 VSS.n7336 VSS.n7335 0.00321084
R12125 VSS.n7346 VSS.n7345 0.00321084
R12126 VSS.n2343 VSS.n2341 0.00320903
R12127 VSS.n2930 VSS.n2254 0.00320903
R12128 VSS.n2340 VSS.n2322 0.00320903
R12129 VSS.n2848 VSS.n2386 0.00320903
R12130 VSS.n4028 VSS.n4027 0.00319767
R12131 VSS.n4046 VSS.n4045 0.00319767
R12132 VSS.n4041 VSS.n4040 0.00319767
R12133 VSS.n3018 VSS.n2137 0.00317559
R12134 VSS.n3016 VSS.n2144 0.00317559
R12135 VSS.n2165 VSS.n2154 0.00317559
R12136 VSS.n3002 VSS.n3001 0.00317559
R12137 VSS.n2947 VSS.n2946 0.00317559
R12138 VSS.n4002 VSS.n4001 0.00317281
R12139 VSS.n4006 VSS.n4005 0.00317281
R12140 VSS.n4011 VSS.n4010 0.00317281
R12141 VSS.n4015 VSS.n4014 0.00317281
R12142 VSS.n7845 VSS.n7844 0.00316667
R12143 VSS.n3356 VSS.n3355 0.00315896
R12144 VSS.n685 VSS.n684 0.00313878
R12145 VSS.n2106 VSS.n2105 0.00313793
R12146 VSS.n2104 VSS.n2103 0.00313793
R12147 VSS.n2103 VSS.n2102 0.00313793
R12148 VSS.n2102 VSS.n2101 0.00313793
R12149 VSS.n2098 VSS.n2097 0.00313793
R12150 VSS.n2095 VSS.n2093 0.00313793
R12151 VSS.n2089 VSS.n2088 0.00313793
R12152 VSS.n2042 VSS.n2041 0.00313793
R12153 VSS.n2025 VSS.n2023 0.00313793
R12154 VSS.n2689 VSS.n2607 0.00312009
R12155 VSS.n3456 VSS.n3455 0.00311628
R12156 VSS.n3449 VSS.n3448 0.00311628
R12157 VSS.n3386 VSS.n3385 0.00311628
R12158 VSS.n3231 VSS.n3230 0.00311628
R12159 VSS.n3280 VSS.n3275 0.00311628
R12160 VSS.n2786 VSS.n2785 0.00311628
R12161 VSS.n3027 VSS.n2137 0.0031087
R12162 VSS.n3017 VSS.n3016 0.0031087
R12163 VSS.n2154 VSS.n2153 0.0031087
R12164 VSS.n3002 VSS.n2168 0.0031087
R12165 VSS.n2947 VSS.n2243 0.0031087
R12166 VSS.n4049 VSS.n4048 0.00310465
R12167 VSS.n1864 VSS.n1863 0.00309859
R12168 VSS.n2936 VSS.n2244 0.00307649
R12169 VSS.n2274 VSS.n2265 0.00307649
R12170 VSS.n2878 VSS.n2877 0.00307649
R12171 VSS.n2229 VSS.n2228 0.00305853
R12172 VSS.n2232 VSS.n2231 0.00305853
R12173 VSS.n2995 VSS.n2994 0.00305853
R12174 VSS.n2182 VSS.n2174 0.00305853
R12175 VSS.n2983 VSS.n2182 0.00305853
R12176 VSS.n2983 VSS.n2982 0.00305853
R12177 VSS.n2968 VSS.n2967 0.00305853
R12178 VSS.n2214 VSS.n2213 0.00305853
R12179 VSS.n2225 VSS.n2224 0.00305853
R12180 VSS.n2992 VSS.n2175 0.00305853
R12181 VSS.n2962 VSS.n2961 0.00305853
R12182 VSS.n2991 VSS.n2177 0.00305853
R12183 VSS.n2963 VSS.n2209 0.00305853
R12184 VSS.n2925 VSS.n2260 0.00305853
R12185 VSS.n2415 VSS.n2414 0.00305853
R12186 VSS.n2837 VSS.n2836 0.00305853
R12187 VSS.n2836 VSS.n2416 0.00305853
R12188 VSS.n2452 VSS.n2416 0.00305853
R12189 VSS.n2457 VSS.n2456 0.00305853
R12190 VSS.n2835 VSS.n2399 0.00305853
R12191 VSS.n2835 VSS.n2417 0.00305853
R12192 VSS.n2455 VSS.n2443 0.00305853
R12193 VSS.n2834 VSS.n2419 0.00305853
R12194 VSS.n1881 VSS.n1880 0.00304301
R12195 VSS.n3960 VSS.n3959 0.00301748
R12196 VSS.n3991 VSS.n3990 0.00301748
R12197 VSS.n2867 VSS.n2360 0.00301572
R12198 VSS.n2865 VSS.n2367 0.00301572
R12199 VSS.n2813 VSS.n2812 0.00301572
R12200 VSS.n2945 VSS.n2244 0.00301208
R12201 VSS.n2935 VSS.n2934 0.00301208
R12202 VSS.n2878 VSS.n2359 0.00301208
R12203 VSS.n2697 VSS.n2599 0.00298908
R12204 VSS.n3299 VSS.n3298 0.00298547
R12205 VSS.n3182 VSS.n3176 0.00298547
R12206 VSS.n2571 VSS.n2570 0.00298547
R12207 VSS.n2755 VSS.n2546 0.00298547
R12208 VSS.n2569 VSS.n2557 0.00298547
R12209 VSS.n2743 VSS.n2559 0.00298547
R12210 VSS.n2746 VSS.n2556 0.00298547
R12211 VSS.n2747 VSS.n2551 0.00298547
R12212 VSS.n2105 VSS.n2104 0.00298276
R12213 VSS.n2101 VSS.n2100 0.00298276
R12214 VSS.n2022 VSS.n2021 0.00298276
R12215 VSS.n5717 VSS.n5716 0.00297253
R12216 VSS.n4910 VSS.n4909 0.00297253
R12217 VSS.n2876 VSS.n2360 0.00295283
R12218 VSS.n2866 VSS.n2865 0.00295283
R12219 VSS.n2846 VSS.n2394 0.00295283
R12220 VSS.n3988 VSS.n3976 0.00292424
R12221 VSS.n2355 VSS.n2354 0.00292012
R12222 VSS.n2815 VSS.n2467 0.00292012
R12223 VSS.n2994 VSS.n2174 0.00290803
R12224 VSS.n2982 VSS.n2183 0.00290803
R12225 VSS.n2993 VSS.n2992 0.00290803
R12226 VSS.n2959 VSS.n2217 0.00290803
R12227 VSS.n2465 VSS.n2451 0.00290803
R12228 VSS.n2838 VSS.n2837 0.00290803
R12229 VSS.n2456 VSS.n2453 0.00290803
R12230 VSS.n2464 VSS.n2457 0.00290803
R12231 VSS.n2458 VSS.n2450 0.00290803
R12232 VSS.n2839 VSS.n2399 0.00290803
R12233 VSS.n2444 VSS.n2443 0.00290803
R12234 VSS.n2823 VSS.n2822 0.00290803
R12235 VSS.n2168 VSS.n2165 0.00290803
R12236 VSS.n3673 VSS.n3672 0.0028968
R12237 VSS.n3760 VSS.n3751 0.0028968
R12238 VSS.n4009 VSS.n4008 0.00289631
R12239 VSS.n3674 VSS.n3673 0.00289361
R12240 VSS.n3761 VSS.n3760 0.00289361
R12241 VSS.n196 VSS.n195 0.00287973
R12242 VSS.n3561 VSS.n3560 0.00285465
R12243 VSS.n3479 VSS.n3469 0.00285465
R12244 VSS.n2975 VSS.n2974 0.00284114
R12245 VSS VSS.n5228 0.00283333
R12246 VSS.n2026 VSS.n2025 0.00282759
R12247 VSS.n2802 VSS.n2469 0.00282558
R12248 VSS.n2506 VSS.n2490 0.00282558
R12249 VSS.n2727 VSS.n2572 0.00282558
R12250 VSS.n3224 VSS.n3209 0.00282558
R12251 VSS.n3207 VSS.n3196 0.00282558
R12252 VSS.n3194 VSS.n3186 0.00282558
R12253 VSS.n3160 VSS.n3149 0.00282558
R12254 VSS.n3107 VSS.n3061 0.00282558
R12255 VSS.n3606 VSS.n3605 0.00282558
R12256 VSS.n3594 VSS.n3593 0.00282558
R12257 VSS.n3794 VSS.n3745 0.00281884
R12258 VSS.n3405 VSS.n3365 0.00281214
R12259 VSS.n3363 VSS.n3356 0.00281214
R12260 VSS.n3326 VSS.n3313 0.00281214
R12261 VSS.n3286 VSS.n3273 0.00281214
R12262 VSS.n3245 VSS.n3227 0.00281214
R12263 VSS.n3530 VSS.n3523 0.00281214
R12264 VSS.n3440 VSS.n3427 0.00281214
R12265 VSS.n4752 VSS.n4750 0.00280769
R12266 VSS.n3791 VSS.n3790 0.00278682
R12267 VSS.n2715 VSS.n2714 0.00278571
R12268 VSS.n2701 VSS.n2596 0.00278571
R12269 VSS.n2811 VSS.n2469 0.00276744
R12270 VSS.n2801 VSS.n2800 0.00276744
R12271 VSS.n2572 VSS.n2563 0.00276744
R12272 VSS.n3225 VSS.n3224 0.00276744
R12273 VSS.n3208 VSS.n3207 0.00276744
R12274 VSS.n3195 VSS.n3194 0.00276744
R12275 VSS.n3108 VSS.n3107 0.00276744
R12276 VSS.n3744 VSS.n3743 0.00276744
R12277 VSS.n3743 VSS.n3742 0.00276744
R12278 VSS.n3741 VSS.n3740 0.00276744
R12279 VSS.n3739 VSS.n3738 0.00276744
R12280 VSS.n3595 VSS.n3594 0.00276744
R12281 VSS.n1908 VSS.n1898 0.00276087
R12282 VSS.n3857 VSS.n3856 0.00276087
R12283 VSS.n3795 VSS.n3794 0.00276087
R12284 VSS.n2964 VSS.n2963 0.00275752
R12285 VSS.n2933 VSS.n2932 0.00275752
R12286 VSS.n2847 VSS.n2388 0.00275752
R12287 VSS.n3406 VSS.n3405 0.00275434
R12288 VSS.n3364 VSS.n3363 0.00275434
R12289 VSS.n3272 VSS.n3271 0.00275434
R12290 VSS.n3586 VSS.n3585 0.00275434
R12291 VSS.n3441 VSS.n3440 0.00275434
R12292 VSS.n2726 VSS.n2573 0.00272857
R12293 VSS.n2596 VSS.n2584 0.00272857
R12294 VSS.n2648 VSS.n2602 0.00272707
R12295 VSS.n2694 VSS.n2593 0.00272707
R12296 VSS.n2649 VSS.n2603 0.00272707
R12297 VSS.n2690 VSS.n2605 0.00272707
R12298 VSS.n2666 VSS.n2655 0.00272707
R12299 VSS.n3639 VSS.n3638 0.00272384
R12300 VSS.n3285 VSS.n3274 0.00272384
R12301 VSS.n3085 VSS.n3084 0.00272384
R12302 VSS.n3094 VSS.n3093 0.00272384
R12303 VSS.n3079 VSS.n3078 0.00272384
R12304 VSS.n3081 VSS.n3080 0.00272384
R12305 VSS.n3082 VSS.n3081 0.00272384
R12306 VSS.n3083 VSS.n3082 0.00272384
R12307 VSS.n3090 VSS.n3089 0.00272384
R12308 VSS.n3095 VSS.n3092 0.00272384
R12309 VSS.n3099 VSS.n3098 0.00272384
R12310 VSS VSS.n645 0.0027028
R12311 VSS.n645 VSS 0.0027028
R12312 VSS.n1540 VSS.n1539 0.0027028
R12313 VSS.n1540 VSS.n1501 0.0027028
R12314 VSS.n1546 VSS.n1501 0.0027028
R12315 VSS VSS.n1498 0.0027028
R12316 VSS VSS.n1498 0.0027028
R12317 VSS.n2376 VSS.n2367 0.00270126
R12318 VSS.n6270 VSS.n6267 0.00269512
R12319 VSS.n556 VSS.n543 0.00269512
R12320 VSS.n4442 VSS.n4439 0.00269512
R12321 VSS.n2900 VSS.n2313 0.00269002
R12322 VSS.n2051 VSS.n2050 0.00267241
R12323 VSS.n1988 VSS.n1987 0.00267241
R12324 VSS.n1985 VSS.n1984 0.00267241
R12325 VSS.n1993 VSS.n1992 0.00267241
R12326 VSS.n2005 VSS.n2004 0.00267241
R12327 VSS.n2045 VSS.n2044 0.00267241
R12328 VSS.n2037 VSS.n2036 0.00267241
R12329 VSS.n2030 VSS.n2029 0.00267241
R12330 VSS.n2020 VSS.n2019 0.00267241
R12331 VSS.n4500 VSS.n714 0.00266
R12332 VSS.n3608 VSS.n3607 0.00265116
R12333 VSS.n3597 VSS.n3596 0.00265116
R12334 VSS.n2913 VSS.n2275 0.0026256
R12335 VSS.n2125 VSS.n2124 0.00260962
R12336 VSS.n2996 VSS.n2172 0.00260702
R12337 VSS.n2985 VSS.n2175 0.00260702
R12338 VSS.n2981 VSS.n2181 0.00260702
R12339 VSS.n2969 VSS.n2202 0.00260702
R12340 VSS.n2222 VSS.n2221 0.00260702
R12341 VSS.n2998 VSS.n2170 0.00260702
R12342 VSS.n2979 VSS.n2185 0.00260702
R12343 VSS.n2971 VSS.n2200 0.00260702
R12344 VSS.n2956 VSS.n2955 0.00260702
R12345 VSS.n2924 VSS.n2262 0.00260702
R12346 VSS.n2437 VSS.n2436 0.00260702
R12347 VSS.n2843 VSS.n2396 0.00260702
R12348 VSS.n2419 VSS.n2418 0.00260702
R12349 VSS.n2831 VSS.n2830 0.00260702
R12350 VSS.n2694 VSS.n2693 0.00259607
R12351 VSS.n2647 VSS.n2617 0.00259607
R12352 VSS.n2695 VSS.n2601 0.00259607
R12353 VSS.n2667 VSS.n2646 0.00259607
R12354 VSS.n2673 VSS.n2621 0.00259607
R12355 VSS.n2666 VSS.n2643 0.00259607
R12356 VSS.n3557 VSS.n3556 0.00259302
R12357 VSS.n3388 VSS.n3387 0.00259302
R12358 VSS.n3291 VSS.n3290 0.00259302
R12359 VSS.n3080 VSS.n3079 0.00259302
R12360 VSS.n3087 VSS.n3083 0.00259302
R12361 VSS.n3181 VSS.n3180 0.00259302
R12362 VSS.n3125 VSS.n3124 0.00259302
R12363 VSS.n2754 VSS.n2753 0.00259302
R12364 VSS.n2741 VSS.n2560 0.00259302
R12365 VSS.n2549 VSS.n2548 0.00259302
R12366 VSS.n2739 VSS.n2562 0.00259302
R12367 VSS.n3196 VSS.n3195 0.00259302
R12368 VSS.n3808 VSS.n3797 0.00258696
R12369 VSS.n3271 VSS.n3260 0.00258092
R12370 VSS.n3585 VSS.n3532 0.00258092
R12371 VSS.n2716 VSS.n2583 0.00255714
R12372 VSS.n1967 VSS.n1966 0.00254545
R12373 VSS.n3820 VSS.n3819 0.00252899
R12374 VSS.n3057 VSS.n3056 0.00252532
R12375 VSS.n3054 VSS.n3053 0.00252532
R12376 VSS.n3051 VSS.n3050 0.00252532
R12377 VSS.n3029 VSS.n3028 0.00252532
R12378 VSS.n3309 VSS.n3302 0.00252312
R12379 VSS.n3259 VSS.n3258 0.00252312
R12380 VSS.n3531 VSS.n3530 0.00252312
R12381 VSS.n3426 VSS.n3425 0.00252312
R12382 VSS.n3424 VSS.n3417 0.00252312
R12383 VSS.n3408 VSS.n3407 0.00252312
R12384 VSS.n2090 VSS.n2089 0.00251724
R12385 VSS.n2007 VSS.n2006 0.00251724
R12386 VSS.n3058 VSS.n3057 0.00247468
R12387 VSS.n3055 VSS.n3054 0.00247468
R12388 VSS.n3052 VSS.n3051 0.00247468
R12389 VSS.n3042 VSS.n3041 0.00247468
R12390 VSS.n3030 VSS.n3029 0.00247468
R12391 VSS.n1909 VSS.n1908 0.00247101
R12392 VSS.n3560 VSS.n3559 0.00246221
R12393 VSS.n3472 VSS.n3471 0.00246221
R12394 VSS.n3476 VSS.n3473 0.00246221
R12395 VSS.n3468 VSS.n3467 0.00246221
R12396 VSS.n3369 VSS.n3368 0.00246221
R12397 VSS.n3143 VSS.n3135 0.00246221
R12398 VSS.n2224 VSS.n2216 0.00245652
R12399 VSS.n2980 VSS.n2184 0.00245652
R12400 VSS.n2960 VSS.n2215 0.00245652
R12401 VSS.n2342 VSS.n2333 0.00245652
R12402 VSS.n2928 VSS.n2927 0.00245652
R12403 VSS.n2335 VSS.n2334 0.00245652
R12404 VSS.n2344 VSS.n2343 0.00245652
R12405 VSS.n2350 VSS.n2346 0.00245652
R12406 VSS.n2929 VSS.n2256 0.00245652
R12407 VSS.n2323 VSS.n2322 0.00245652
R12408 VSS.n2890 VSS.n2889 0.00245652
R12409 VSS.n2412 VSS.n2403 0.00245652
R12410 VSS.n2409 VSS.n2406 0.00245652
R12411 VSS.n2411 VSS.n2410 0.00245652
R12412 VSS.n2851 VSS.n2383 0.00245652
R12413 VSS.n2402 VSS.n2401 0.00245652
R12414 VSS.n2379 VSS.n2378 0.00245652
R12415 VSS.n2400 VSS.n2398 0.00245652
R12416 VSS.n2454 VSS.n2438 0.00245652
R12417 VSS.n2460 VSS.n2449 0.00245652
R12418 VSS.n2856 VSS.n2855 0.00245652
R12419 VSS.n2827 VSS.n2826 0.00245652
R12420 VSS.n2447 VSS.n2445 0.00245652
R12421 VSS.n2818 VSS.n2817 0.00245652
R12422 VSS.n3001 VSS.n2169 0.0024398
R12423 VSS VSS.n636 0.00238811
R12424 VSS.n7909 VSS.n7908 0.00236306
R12425 VSS.n2096 VSS.n2095 0.00236207
R12426 VSS.n3858 VSS.n3857 0.00235507
R12427 VSS.n2668 VSS.n2653 0.00233406
R12428 VSS.n2696 VSS.n2600 0.00233406
R12429 VSS.n2667 VSS.n2654 0.00233406
R12430 VSS.n2698 VSS.n2598 0.00233406
R12431 VSS.n3549 VSS.n3548 0.0023314
R12432 VSS.n3459 VSS.n3450 0.0023314
R12433 VSS.n3278 VSS.n3277 0.0023314
R12434 VSS.n3325 VSS.n3315 0.0023314
R12435 VSS.n3179 VSS.n3178 0.0023314
R12436 VSS.n3167 VSS.n3166 0.0023314
R12437 VSS.n3138 VSS.n3137 0.0023314
R12438 VSS.n3116 VSS.n3115 0.0023314
R12439 VSS.n3175 VSS.n3174 0.0023314
R12440 VSS.n3132 VSS.n3131 0.0023314
R12441 VSS.n3123 VSS.n3122 0.0023314
R12442 VSS.n2747 VSS.n2555 0.0023314
R12443 VSS.n3053 VSS.n3052 0.00232278
R12444 VSS.n5369 VSS.n5365 0.00231452
R12445 VSS.n7733 VSS.n7728 0.00231452
R12446 VSS.n2213 VSS.n2205 0.00230602
R12447 VSS.n2962 VSS.n2206 0.00230602
R12448 VSS.n2267 VSS.n2266 0.00230602
R12449 VSS.n2153 VSS.n2144 0.00230602
R12450 VSS.n2912 VSS.n2276 0.00230354
R12451 VSS.n3834 VSS.n3823 0.0022971
R12452 VSS.n2662 VSS.n2656 0.00224426
R12453 VSS.n2800 VSS.n2799 0.00224419
R12454 VSS.n5904 VSS.n5903 0.00224148
R12455 VSS.n2123 VSS.n2118 0.00222181
R12456 VSS.n2041 VSS.n2040 0.0022069
R12457 VSS.n2693 VSS.n2692 0.00220306
R12458 VSS.n2671 VSS.n2647 0.00220306
R12459 VSS.n2644 VSS.n2619 0.00220306
R12460 VSS.n2672 VSS.n2645 0.00220306
R12461 VSS.n2661 VSS.n2660 0.00220306
R12462 VSS.n2677 VSS.n2676 0.00220306
R12463 VSS.n3570 VSS.n3569 0.00220058
R12464 VSS.n3566 VSS.n3565 0.00220058
R12465 VSS.n3563 VSS.n3562 0.00220058
R12466 VSS.n3387 VSS.n3386 0.00220058
R12467 VSS.n3332 VSS.n3331 0.00220058
R12468 VSS.n3293 VSS.n3292 0.00220058
R12469 VSS.n3098 VSS.n3097 0.00220058
R12470 VSS.n3156 VSS.n3153 0.00220058
R12471 VSS.n3118 VSS.n3117 0.00220058
R12472 VSS.n2492 VSS.n2491 0.00220058
R12473 VSS.n2752 VSS.n2751 0.00220058
R12474 VSS.n2389 VSS.n2377 0.00219811
R12475 VSS.n3025 VSS.n2139 0.00219111
R12476 VSS.n2943 VSS.n2246 0.00219111
R12477 VSS.n2874 VSS.n2362 0.00219111
R12478 VSS.n2789 VSS.n2478 0.00218605
R12479 VSS.n2511 VSS.n2510 0.00218605
R12480 VSS.n2776 VSS.n2775 0.00218605
R12481 VSS.n2530 VSS.n2512 0.00218605
R12482 VSS.n3186 VSS.n3185 0.00218605
R12483 VSS.n3592 VSS.n3591 0.00218605
R12484 VSS.n3590 VSS.n3589 0.00218605
R12485 VSS.n3588 VSS.n3587 0.00218605
R12486 VSS.n1895 VSS.n1887 0.00218116
R12487 VSS.n1897 VSS.n1896 0.00218116
R12488 VSS.n3856 VSS.n3840 0.00218116
R12489 VSS.n3355 VSS.n3354 0.0021763
R12490 VSS.n3353 VSS.n3342 0.0021763
R12491 VSS.n5841 VSS.n5442 0.00216667
R12492 VSS.n5837 VSS.n5836 0.00216667
R12493 VSS.n5854 VSS.n5853 0.00216667
R12494 VSS.n5867 VSS.n5864 0.00216667
R12495 VSS.n1777 VSS.n1776 0.0021589
R12496 VSS.n2636 VSS.n2635 0.00215714
R12497 VSS.n2987 VSS.n2177 0.00215552
R12498 VSS.n2464 VSS.n2463 0.00215552
R12499 VSS.n7797 VSS.n7796 0.00214634
R12500 VSS.n2858 VSS.n2857 0.00213522
R12501 VSS.n3838 VSS.n3837 0.00212319
R12502 VSS.n3312 VSS.n3311 0.0021185
R12503 VSS.n2264 VSS.n2251 0.00211031
R12504 VSS.n2887 VSS.n2886 0.00211031
R12505 VSS.n2650 VSS.n2649 0.00207205
R12506 VSS.n3571 VSS.n3570 0.00206977
R12507 VSS.n3568 VSS.n3566 0.00206977
R12508 VSS.n3564 VSS.n3563 0.00206977
R12509 VSS.n3500 VSS.n3499 0.00206977
R12510 VSS.n3092 VSS.n3091 0.00206977
R12511 VSS.n3142 VSS.n3141 0.00206977
R12512 VSS.n3209 VSS.n3208 0.00206977
R12513 VSS.n3859 VSS.n3858 0.00206522
R12514 VSS.n2724 VSS.n2575 0.0020629
R12515 VSS.n3620 VSS.n3619 0.00206165
R12516 VSS.n3583 VSS.n3578 0.00206165
R12517 VSS.n2012 VSS.n2011 0.0020532
R12518 VSS.n2035 VSS.n2034 0.00205172
R12519 VSS.n2669 VSS.n2668 0.00204803
R12520 VSS.n2670 VSS.n2669 0.00204706
R12521 VSS.n2892 VSS.n2891 0.00204589
R12522 VSS.n2949 VSS.n2236 0.00202155
R12523 VSS.n2978 VSS.n2186 0.00200502
R12524 VSS.n2337 VSS.n2316 0.00200502
R12525 VSS.n2348 VSS.n2347 0.00200502
R12526 VSS.n2895 VSS.n2894 0.00200502
R12527 VSS.n2885 VSS.n2884 0.00200502
R12528 VSS.n2466 VSS.n2450 0.00200502
R12529 VSS.n2407 VSS.n2373 0.00200502
R12530 VSS.n2853 VSS.n2852 0.00200502
R12531 VSS.n2860 VSS.n2859 0.00200502
R12532 VSS.n2391 VSS.n2380 0.00200502
R12533 VSS.n7353 VSS.n7352 0.002
R12534 VSS.n2990 VSS.n2178 0.00197157
R12535 VSS.n3050 VSS.n3049 0.00196835
R12536 VSS.n3604 VSS.n3603 0.00195349
R12537 VSS.n1781 VSS.n1780 0.00195161
R12538 VSS.n1793 VSS.n1791 0.00195161
R12539 VSS.n1795 VSS.n1794 0.00195161
R12540 VSS.n1797 VSS.n1796 0.00195161
R12541 VSS.n1803 VSS.n1802 0.00195161
R12542 VSS.n1812 VSS.n1811 0.00195161
R12543 VSS.n1822 VSS.n1821 0.00195161
R12544 VSS.n2833 VSS.n2832 0.00194654
R12545 VSS.n2825 VSS.n2824 0.00194654
R12546 VSS.n3328 VSS.n3327 0.00194509
R12547 VSS.n3726 VSS.n3725 0.00193895
R12548 VSS.n3722 VSS.n3721 0.00193895
R12549 VSS.n3711 VSS.n3710 0.00193895
R12550 VSS.n3555 VSS.n3553 0.00193895
R12551 VSS.n3458 VSS.n3457 0.00193895
R12552 VSS.n3518 VSS.n3510 0.00193895
R12553 VSS.n3172 VSS.n3171 0.00193895
R12554 VSS.n2744 VSS.n2557 0.00193895
R12555 VSS.n2746 VSS.n2745 0.00193895
R12556 VSS.n2923 VSS.n2922 0.00191707
R12557 VSS.n5948 VSS.n5945 0.00189535
R12558 VSS.n6234 VSS.n6232 0.00189535
R12559 VSS.n3242 VSS.n3241 0.00188813
R12560 VSS.n3104 VSS.n3103 0.00188813
R12561 VSS.n2729 VSS.n2566 0.00188813
R12562 VSS.n3258 VSS.n3247 0.00188728
R12563 VSS.n3056 VSS.n3055 0.00186709
R12564 VSS.n3403 VSS.n3398 0.00186205
R12565 VSS.n2809 VSS.n2471 0.00186205
R12566 VSS.n150 VSS.n147 0.00185388
R12567 VSS.n2921 VSS.n2265 0.00185266
R12568 VSS.n4156 VSS.n4139 0.00185193
R12569 VSS.n1132 VSS.n1127 0.00184731
R12570 VSS.n3602 VSS.n3601 0.00183721
R12571 VSS.n1898 VSS.n1897 0.00183333
R12572 VSS.n3246 VSS.n3245 0.00182948
R12573 VSS.n3443 VSS.n3442 0.00182948
R12574 VSS.n4877 VSS.n4876 0.0018278
R12575 VSS.n2688 VSS.n2687 0.00181429
R12576 VSS.n2723 VSS.n2722 0.00181004
R12577 VSS.n2604 VSS.n2601 0.00181004
R12578 VSS.n3558 VSS.n3557 0.00180814
R12579 VSS.n3515 VSS.n3514 0.00180814
R12580 VSS.n3489 VSS.n3488 0.00180814
R12581 VSS.n3509 VSS.n3508 0.00180814
R12582 VSS.n3496 VSS.n3495 0.00180814
R12583 VSS.n3378 VSS.n3377 0.00180814
R12584 VSS.n3334 VSS.n3333 0.00180814
R12585 VSS.n3297 VSS.n3296 0.00180814
R12586 VSS.n3255 VSS.n3254 0.00180814
R12587 VSS.n3159 VSS.n3151 0.00180814
R12588 VSS.n2768 VSS.n2767 0.00180814
R12589 VSS.n2568 VSS.n2546 0.00180814
R12590 VSS.n2550 VSS.n2547 0.00180814
R12591 VSS.n3872 VSS.n3864 0.00180814
R12592 VSS.n2763 VSS.n2762 0.00177907
R12593 VSS.n3184 VSS.n3183 0.00177907
R12594 VSS.n3599 VSS.n3598 0.00177907
R12595 VSS.n3288 VSS.n3287 0.00177168
R12596 VSS.n3464 VSS.n3461 0.00177168
R12597 VSS.n2958 VSS.n2957 0.0017709
R12598 VSS.n3910 VSS.n3909 0.00176168
R12599 VSS.n3986 VSS.n3979 0.00176168
R12600 VSS.n1597 VSS.n1489 0.00175874
R12601 VSS.n2699 VSS.n2597 0.00175714
R12602 VSS.n1801 VSS.n1799 0.00174752
R12603 VSS.n1840 VSS.n1839 0.00174424
R12604 VSS.n1852 VSS.n1851 0.00174424
R12605 VSS.n2789 VSS.n2788 0.00172093
R12606 VSS.n1911 VSS.n1910 0.00171739
R12607 VSS.n3313 VSS.n3312 0.00171387
R12608 VSS.n2459 VSS.n2444 0.00170401
R12609 VSS.n2212 VSS.n2211 0.00170401
R12610 VSS.n2820 VSS.n2819 0.00169497
R12611 VSS.n2589 VSS.n2577 0.00167904
R12612 VSS.n2612 VSS.n2611 0.00167904
R12613 VSS.n3700 VSS.n3692 0.00167733
R12614 VSS.n3565 VSS.n3564 0.00167733
R12615 VSS.n3513 VSS.n3512 0.00167733
R12616 VSS.n3493 VSS.n3492 0.00167733
R12617 VSS.n3491 VSS.n3490 0.00167733
R12618 VSS.n3507 VSS.n3506 0.00167733
R12619 VSS.n3498 VSS.n3497 0.00167733
R12620 VSS.n3755 VSS.n3754 0.00167733
R12621 VSS.n3777 VSS.n3776 0.00167733
R12622 VSS.n3779 VSS.n3778 0.00167733
R12623 VSS.n3781 VSS.n3780 0.00167733
R12624 VSS.n1923 VSS.n1916 0.00167733
R12625 VSS.n2787 VSS.n2490 0.00166279
R12626 VSS.n2922 VSS.n2921 0.00165942
R12627 VSS.n2312 VSS.n2311 0.00165942
R12628 VSS.n3481 VSS.n3480 0.00165607
R12629 VSS.n2665 VSS.n2664 0.00164286
R12630 VSS.n2178 VSS.n2169 0.00163712
R12631 VSS.n2990 VSS.n2989 0.00163712
R12632 VSS.n2977 VSS.n2179 0.00163712
R12633 VSS.n2210 VSS.n2198 0.00163712
R12634 VSS.n2218 VSS.n2212 0.00163712
R12635 VSS.n2957 VSS.n2219 0.00163712
R12636 VSS.n7572 VSS.n7558 0.00163208
R12637 VSS.n7568 VSS.n7567 0.00163208
R12638 VSS.n7540 VSS.n5354 0.00163208
R12639 VSS.n3911 VSS.n3908 0.00163049
R12640 VSS.n3048 VSS.n3047 0.00161392
R12641 VSS.n5037 VSS.n5036 0.00161111
R12642 VSS.n5031 VSS.n5028 0.00161111
R12643 VSS.n5018 VSS.n5017 0.00161111
R12644 VSS.n4989 VSS.n4982 0.00161111
R12645 VSS.n2788 VSS.n2787 0.00160465
R12646 VSS.n2553 VSS.n2552 0.00160465
R12647 VSS.n2749 VSS.n2748 0.00160465
R12648 VSS.n2738 VSS.n2737 0.00160465
R12649 VSS.n3126 VSS.n3111 0.00160465
R12650 VSS.n3874 VSS.n1924 0.00160145
R12651 VSS.n6304 VSS.n6302 0.00159756
R12652 VSS.n4703 VSS.n4701 0.00159756
R12653 VSS.n2675 VSS.n2674 0.00158571
R12654 VSS.n2845 VSS.n2844 0.00156918
R12655 VSS.n2832 VSS.n2434 0.00156918
R12656 VSS.n2463 VSS.n2458 0.00155351
R12657 VSS.n2462 VSS.n2461 0.00155351
R12658 VSS.n2816 VSS.n2815 0.00155351
R12659 VSS.n3896 VSS.n3895 0.0015514
R12660 VSS.n3966 VSS.n3965 0.0015514
R12661 VSS.n3968 VSS.n3967 0.0015514
R12662 VSS.n3974 VSS.n3964 0.0015514
R12663 VSS.n2685 VSS.n2684 0.00154803
R12664 VSS.n3691 VSS.n3690 0.00154651
R12665 VSS.n3687 VSS.n3686 0.00154651
R12666 VSS.n3654 VSS.n3653 0.00154651
R12667 VSS.n3705 VSS.n3704 0.00154651
R12668 VSS.n3575 VSS.n3574 0.00154651
R12669 VSS.n3569 VSS.n3568 0.00154651
R12670 VSS.n3559 VSS.n3558 0.00154651
R12671 VSS.n3517 VSS.n3516 0.00154651
R12672 VSS.n3436 VSS.n3435 0.00154651
R12673 VSS.n3234 VSS.n3233 0.00154651
R12674 VSS.n3341 VSS.n3340 0.00154651
R12675 VSS.n3283 VSS.n3282 0.00154651
R12676 VSS.n2764 VSS.n2763 0.00154651
R12677 VSS.n3145 VSS.n3144 0.00154651
R12678 VSS.n1894 VSS.n1893 0.00154651
R12679 VSS.n3483 VSS.n3482 0.00154046
R12680 VSS.n921 VSS.n812 0.00153687
R12681 VSS.n1808 VSS.n1807 0.00153687
R12682 VSS.n1810 VSS.n1809 0.00153687
R12683 VSS.n1818 VSS.n1817 0.00153687
R12684 VSS.n1820 VSS.n1819 0.00153687
R12685 VSS.n1828 VSS.n1827 0.00153687
R12686 VSS.n2825 VSS.n2441 0.00150629
R12687 VSS.n2824 VSS.n2442 0.00150629
R12688 VSS.n2819 VSS.n2446 0.00150629
R12689 VSS.n1871 VSS.n1870 0.00150559
R12690 VSS.n4078 VSS.n4077 0.00150559
R12691 VSS.n4073 VSS.n4072 0.00150559
R12692 VSS.n4071 VSS.n4070 0.00150559
R12693 VSS.n2748 VSS.n2554 0.00148837
R12694 VSS.n3185 VSS.n3184 0.00148837
R12695 VSS.n3183 VSS.n3173 0.00148837
R12696 VSS.n3162 VSS.n3161 0.00148837
R12697 VSS.n3147 VSS.n3146 0.00148837
R12698 VSS.n3144 VSS.n3129 0.00148837
R12699 VSS.n3111 VSS.n3110 0.00148837
R12700 VSS.n3287 VSS.n3286 0.00148266
R12701 VSS.n3460 VSS.n3443 0.00148266
R12702 VSS.n2700 VSS.n2699 0.00147143
R12703 VSS.n2934 VSS.n2251 0.00146618
R12704 VSS.n3034 VSS.n3033 0.00146203
R12705 VSS.n4118 VSS.n4117 0.00144995
R12706 VSS.n4109 VSS.n4108 0.00144995
R12707 VSS.n4118 VSS.n4115 0.00144995
R12708 VSS.n4109 VSS.n4106 0.00144995
R12709 VSS VSS.n630 0.00144406
R12710 VSS.n2846 VSS.n2845 0.0014434
R12711 VSS.n2433 VSS.n2432 0.0014434
R12712 VSS.n2039 VSS.n2038 0.00143104
R12713 VSS.n2750 VSS.n2553 0.00143023
R12714 VSS.n3247 VSS.n3246 0.00142485
R12715 VSS.n3465 VSS.n3464 0.00142485
R12716 VSS.n2578 VSS.n2575 0.00141703
R12717 VSS.n2608 VSS.n2599 0.00141703
R12718 VSS.n2689 VSS.n2606 0.00141703
R12719 VSS.n3707 VSS.n3706 0.0014157
R12720 VSS.n3556 VSS.n3555 0.0014157
R12721 VSS.n3352 VSS.n3346 0.0014157
R12722 VSS.n2497 VSS.n2484 0.0014157
R12723 VSS.n2496 VSS.n2495 0.0014157
R12724 VSS.n2766 VSS.n2525 0.0014157
R12725 VSS.n2778 VSS.n2777 0.0014157
R12726 VSS.n3771 VSS.n3770 0.0014157
R12727 VSS.n3871 VSS.n3870 0.0014157
R12728 VSS.n1886 VSS.n1881 0.0014157
R12729 VSS.n2675 VSS.n2641 0.00141429
R12730 VSS.n2665 VSS.n2642 0.00141429
R12731 VSS.n3037 VSS.n3036 0.00141139
R12732 VSS.n2986 VSS.n2180 0.00140301
R12733 VSS.n2287 VSS.n2259 0.00140301
R12734 VSS.n2286 VSS.n2284 0.00140301
R12735 VSS.n2923 VSS.n2264 0.00140177
R12736 VSS.n1775 VSS.n1766 0.0014
R12737 VSS.n1773 VSS.n1768 0.0014
R12738 VSS.n1772 VSS.n1770 0.0014
R12739 VSS.n4089 VSS.n4088 0.0014
R12740 VSS.n4083 VSS.n4082 0.0014
R12741 VSS.n4122 VSS.n4121 0.0014
R12742 VSS.n4097 VSS.n4095 0.0014
R12743 VSS.n1879 VSS.n1878 0.0014
R12744 VSS.n1877 VSS.n1875 0.0014
R12745 VSS.n1783 VSS.n1782 0.0014
R12746 VSS.n1762 VSS.n1760 0.0014
R12747 VSS.n1763 VSS.n1758 0.0014
R12748 VSS.n1765 VSS.n1756 0.0014
R12749 VSS.n2432 VSS.n2395 0.0013805
R12750 VSS.n3600 VSS.n3599 0.00137209
R12751 VSS.n3365 VSS.n3364 0.00136705
R12752 VSS.n3501 VSS.n3486 0.00136705
R12753 VSS.n3049 VSS.n3048 0.00136076
R12754 VSS.n3047 VSS.n3046 0.00136076
R12755 VSS.n3044 VSS.n3043 0.00136076
R12756 VSS.n3039 VSS.n3038 0.00136076
R12757 VSS.n3036 VSS.n3035 0.00136076
R12758 VSS.n3033 VSS.n3032 0.00136076
R12759 VSS.n3915 VSS.n3914 0.00134112
R12760 VSS.n3913 VSS.n3912 0.00134112
R12761 VSS.n3984 VSS.n3983 0.00134112
R12762 VSS.n3893 VSS.n3892 0.00134112
R12763 VSS.n3962 VSS.n3961 0.00134112
R12764 VSS.n3964 VSS.n3963 0.00134112
R12765 VSS.n3975 VSS.n3960 0.00133916
R12766 VSS.n3990 VSS.n3989 0.00133916
R12767 VSS.n2893 VSS.n2319 0.00133736
R12768 VSS.n2891 VSS.n2320 0.00133736
R12769 VSS.n2886 VSS.n2326 0.00133736
R12770 VSS.n1835 VSS.n1834 0.00132949
R12771 VSS.n1837 VSS.n1836 0.00132949
R12772 VSS.n1844 VSS.n1843 0.00132949
R12773 VSS.n1847 VSS.n1846 0.00132949
R12774 VSS.n1849 VSS.n1848 0.00132949
R12775 VSS.n1856 VSS.n1855 0.00132949
R12776 VSS.n1859 VSS.n1858 0.00132949
R12777 VSS.n1806 VSS.n1805 0.00132949
R12778 VSS.n1814 VSS.n1813 0.00132949
R12779 VSS.n1816 VSS.n1815 0.00132949
R12780 VSS.n1824 VSS.n1823 0.00132949
R12781 VSS.n1826 VSS.n1825 0.00132949
R12782 VSS.n2858 VSS.n2376 0.00131761
R12783 VSS.n2857 VSS.n2377 0.00131761
R12784 VSS.n2390 VSS.n2389 0.00131761
R12785 VSS.n3603 VSS.n3602 0.00131395
R12786 VSS.n3327 VSS.n3326 0.00130925
R12787 VSS.n3520 VSS.n3519 0.00130925
R12788 VSS.n2988 VSS.n2179 0.00130268
R12789 VSS.n2719 VSS.n2579 0.00128603
R12790 VSS.n2686 VSS.n2685 0.00128603
R12791 VSS.n3666 VSS.n3665 0.00128488
R12792 VSS.n3701 VSS.n3664 0.00128488
R12793 VSS.n3170 VSS.n3169 0.00128488
R12794 VSS.n2769 VSS.n2516 0.00128488
R12795 VSS.n3767 VSS.n3766 0.00128488
R12796 VSS.n3769 VSS.n3768 0.00128488
R12797 VSS.n1922 VSS.n1921 0.00128488
R12798 VSS.n3826 VSS.n3825 0.00128488
R12799 VSS.n3831 VSS.n3830 0.00128488
R12800 VSS.n6158 VSS.n6109 0.00127586
R12801 VSS.n1755 VSS.n1752 0.00127253
R12802 VSS.n1727 VSS.n1692 0.00127253
R12803 VSS.n1714 VSS.n1632 0.00127253
R12804 VSS.n1630 VSS.n1627 0.00127253
R12805 VSS.n4113 VSS.n4112 0.00125419
R12806 VSS.n4051 VSS.n1871 0.00125419
R12807 VSS.n4077 VSS.n4076 0.00125419
R12808 VSS.n4075 VSS.n4074 0.00125419
R12809 VSS.n4066 VSS.n4065 0.00125419
R12810 VSS.n4065 VSS.n4064 0.00125419
R12811 VSS.n4063 VSS.n4062 0.00125419
R12812 VSS.n4061 VSS.n4060 0.00125419
R12813 VSS.n4059 VSS.n4058 0.00125419
R12814 VSS.n4053 VSS.n4052 0.00125419
R12815 VSS.n3873 VSS.n3859 0.00125362
R12816 VSS.n2822 VSS.n2821 0.00125251
R12817 VSS.n3289 VSS.n3288 0.00125145
R12818 VSS.n3521 VSS.n3520 0.00125145
R12819 VSS.n3504 VSS.n3501 0.00125145
R12820 VSS.n3485 VSS.n3484 0.00125145
R12821 VSS.n2989 VSS.n2988 0.00123579
R12822 VSS.n5374 VSS.n5373 0.00122581
R12823 VSS.n7739 VSS.n7738 0.00122581
R12824 VSS.n7485 VSS.n7484 0.00122581
R12825 VSS.n3163 VSS.n3162 0.00119767
R12826 VSS.n1924 VSS.n1911 0.00119565
R12827 VSS.n3522 VSS.n3521 0.00119364
R12828 VSS.n3519 VSS.n3504 0.00119364
R12829 VSS.n3486 VSS.n3485 0.00119364
R12830 VSS.n2977 VSS.n2976 0.0011689
R12831 VSS.n2650 VSS.n2616 0.00115502
R12832 VSS.n2614 VSS.n2612 0.00115502
R12833 VSS.n3668 VSS.n3667 0.00115407
R12834 VSS.n3684 VSS.n3683 0.00115407
R12835 VSS.n3672 VSS.n3671 0.00115407
R12836 VSS.n3661 VSS.n3660 0.00115407
R12837 VSS.n3650 VSS.n3649 0.00115407
R12838 VSS.n3633 VSS.n3632 0.00115407
R12839 VSS.n3476 VSS.n3475 0.00115407
R12840 VSS.n3389 VSS.n3388 0.00115407
R12841 VSS.n3336 VSS.n3335 0.00115407
R12842 VSS.n2521 VSS.n2516 0.00115407
R12843 VSS.n2520 VSS.n2514 0.00115407
R12844 VSS.n2773 VSS.n2505 0.00115407
R12845 VSS.n3762 VSS.n3761 0.00115407
R12846 VSS.n1891 VSS.n1890 0.00115407
R12847 VSS.n3846 VSS.n3845 0.00115407
R12848 VSS.n4050 VSS.n4028 0.00115116
R12849 VSS.n4047 VSS.n4046 0.00115116
R12850 VSS.n4001 VSS.n4000 0.00114516
R12851 VSS.n4007 VSS.n4006 0.00114516
R12852 VSS.n4010 VSS.n4009 0.00114516
R12853 VSS.n4016 VSS.n4015 0.00114516
R12854 VSS.n3173 VSS.n3163 0.00113953
R12855 VSS.n3593 VSS.n3592 0.00113953
R12856 VSS.n3589 VSS.n3588 0.00113953
R12857 VSS.n1896 VSS.n1895 0.00113768
R12858 VSS.n3342 VSS.n3329 0.00113584
R12859 VSS.n3934 VSS.n3933 0.00113084
R12860 VSS.n3907 VSS.n3906 0.00113084
R12861 VSS.n3906 VSS.n3905 0.00113084
R12862 VSS.n3905 VSS.n3904 0.00113084
R12863 VSS.n3979 VSS.n3978 0.00113084
R12864 VSS.n657 VSS.n656 0.00112937
R12865 VSS.n1585 VSS.n1584 0.00112937
R12866 VSS.n2635 VSS.n2610 0.00112857
R12867 VSS.n1833 VSS.n1832 0.00112212
R12868 VSS.n1836 VSS.n1835 0.00112212
R12869 VSS.n1843 VSS.n1842 0.00112212
R12870 VSS.n1845 VSS.n1844 0.00112212
R12871 VSS.n1848 VSS.n1847 0.00112212
R12872 VSS.n1855 VSS.n1854 0.00112212
R12873 VSS.n1857 VSS.n1856 0.00112212
R12874 VSS.n1815 VSS.n1814 0.00112212
R12875 VSS.n1825 VSS.n1824 0.00112212
R12876 VSS.n2092 VSS.n2091 0.00112069
R12877 VSS.n2097 VSS.n2096 0.00112069
R12878 VSS.n2093 VSS.n2090 0.00112069
R12879 VSS.n2088 VSS.n2087 0.00112069
R12880 VSS.n2023 VSS.n2022 0.00112069
R12881 VSS.n3045 VSS.n3044 0.00110759
R12882 VSS.n2233 VSS.n2232 0.00110201
R12883 VSS.n2967 VSS.n2205 0.00110201
R12884 VSS.n2216 VSS.n2214 0.00110201
R12885 VSS.n2952 VSS.n2225 0.00110201
R12886 VSS.n2961 VSS.n2960 0.00110201
R12887 VSS.n2959 VSS.n2209 0.00110201
R12888 VSS.n2296 VSS.n2279 0.00110201
R12889 VSS.n2838 VSS.n2402 0.00110201
R12890 VSS.n2814 VSS.n2448 0.00110201
R12891 VSS.n2799 VSS.n2478 0.0010814
R12892 VSS.n2776 VSS.n2511 0.0010814
R12893 VSS.n3161 VSS.n3160 0.0010814
R12894 VSS.n3591 VSS.n3590 0.0010814
R12895 VSS.n2901 VSS.n2312 0.00107971
R12896 VSS.n3354 VSS.n3353 0.00107803
R12897 VSS.n2688 VSS.n2609 0.00107143
R12898 VSS.n3890 VSS.n3889 0.00105944
R12899 VSS.n3922 VSS.n3921 0.00105944
R12900 VSS.n4043 VSS.n4042 0.00105814
R12901 VSS.n4039 VSS.n4038 0.00105814
R12902 VSS.n3046 VSS.n3045 0.00105696
R12903 VSS.n4004 VSS.n4003 0.00105299
R12904 VSS.n4013 VSS.n4012 0.00105299
R12905 VSS.n2692 VSS.n2603 0.00102402
R12906 VSS.n2680 VSS.n2617 0.00102402
R12907 VSS.n2671 VSS.n2670 0.00102402
R12908 VSS.n2659 VSS.n2653 0.00102402
R12909 VSS.n2691 VSS.n2690 0.00102402
R12910 VSS.n2672 VSS.n2646 0.00102402
R12911 VSS.n2582 VSS.n2574 0.00102402
R12912 VSS.n2673 VSS.n2643 0.00102402
R12913 VSS.n3685 VSS.n3684 0.00102326
R12914 VSS.n3675 VSS.n3674 0.00102326
R12915 VSS.n3635 VSS.n3634 0.00102326
R12916 VSS.n3458 VSS.n3452 0.00102326
R12917 VSS.n3391 VSS.n3390 0.00102326
R12918 VSS.n3239 VSS.n3238 0.00102326
R12919 VSS.n3351 VSS.n3350 0.00102326
R12920 VSS.n3250 VSS.n3249 0.00102326
R12921 VSS.n3339 VSS.n3338 0.00102326
R12922 VSS.n3091 VSS.n3090 0.00102326
R12923 VSS.n3097 VSS.n3095 0.00102326
R12924 VSS.n3100 VSS.n3099 0.00102326
R12925 VSS.n2570 VSS.n2567 0.00102326
R12926 VSS.n2519 VSS.n2500 0.00102326
R12927 VSS.n2756 VSS.n2755 0.00102326
R12928 VSS.n2569 VSS.n2568 0.00102326
R12929 VSS.n2744 VSS.n2743 0.00102326
R12930 VSS.n2504 VSS.n2502 0.00102326
R12931 VSS.n2556 VSS.n2550 0.00102326
R12932 VSS.n2797 VSS.n2479 0.00102326
R12933 VSS.n2765 VSS.n2528 0.00102326
R12934 VSS.n2751 VSS.n2551 0.00102326
R12935 VSS.n3753 VSS.n3752 0.00102326
R12936 VSS.n3751 VSS.n3750 0.00102326
R12937 VSS.n3783 VSS.n3782 0.00102326
R12938 VSS.n3785 VSS.n3784 0.00102326
R12939 VSS.n3787 VSS.n3786 0.00102326
R12940 VSS.n1885 VSS.n1884 0.00102326
R12941 VSS.n3850 VSS.n3849 0.00102326
R12942 VSS.n4093 VSS.n4092 0.00102326
R12943 VSS.n3840 VSS.n3839 0.00102174
R12944 VSS.n3837 VSS.n3834 0.00102174
R12945 VSS.n3823 VSS.n3822 0.00102174
R12946 VSS.n3043 VSS.n3042 0.00100633
R12947 VSS.n2844 VSS.n2395 0.00100314
R12948 VSS.n4101 VSS.n4099 0.00100279
R12949 VSS.n4070 VSS.n4069 0.00100279
R12950 VSS.n4056 VSS.n4055 0.00100279
R12951 VSS.n3919 VSS.n3903 0.0009662
R12952 VSS.n2122 VSS.n2121 0.000965517
R12953 VSS.n2120 VSS.n2119 0.000965517
R12954 VSS.n2074 VSS.n2073 0.000965517
R12955 VSS.n2072 VSS.n2071 0.000965517
R12956 VSS.n2064 VSS.n2063 0.000965517
R12957 VSS.n2062 VSS.n2061 0.000965517
R12958 VSS.n2054 VSS.n2053 0.000965517
R12959 VSS.n2052 VSS.n2051 0.000965517
R12960 VSS.n2050 VSS.n2049 0.000965517
R12961 VSS.n1987 VSS.n1986 0.000965517
R12962 VSS.n1986 VSS.n1985 0.000965517
R12963 VSS.n1984 VSS.n1983 0.000965517
R12964 VSS.n1996 VSS.n1995 0.000965517
R12965 VSS.n1994 VSS.n1993 0.000965517
R12966 VSS.n1992 VSS.n1991 0.000965517
R12967 VSS.n1990 VSS.n1989 0.000965517
R12968 VSS.n2006 VSS.n2005 0.000965517
R12969 VSS.n2004 VSS.n2003 0.000965517
R12970 VSS.n2002 VSS.n2001 0.000965517
R12971 VSS.n2000 VSS.n1999 0.000965517
R12972 VSS.n2080 VSS.n2079 0.000965517
R12973 VSS.n2078 VSS.n2077 0.000965517
R12974 VSS.n2070 VSS.n2069 0.000965517
R12975 VSS.n2068 VSS.n2067 0.000965517
R12976 VSS.n2060 VSS.n2059 0.000965517
R12977 VSS.n2058 VSS.n2057 0.000965517
R12978 VSS.n2048 VSS.n2047 0.000965517
R12979 VSS.n2046 VSS.n2045 0.000965517
R12980 VSS.n2044 VSS.n2043 0.000965517
R12981 VSS.n2040 VSS.n2039 0.000965517
R12982 VSS.n2038 VSS.n2037 0.000965517
R12983 VSS.n2036 VSS.n2035 0.000965517
R12984 VSS.n2033 VSS.n2032 0.000965517
R12985 VSS.n2031 VSS.n2030 0.000965517
R12986 VSS.n2029 VSS.n2028 0.000965517
R12987 VSS.n2027 VSS.n2026 0.000965517
R12988 VSS.n2021 VSS.n2020 0.000965517
R12989 VSS.n2019 VSS.n2018 0.000965517
R12990 VSS.n2017 VSS.n2016 0.000965517
R12991 VSS.n2015 VSS.n2014 0.000965517
R12992 VSS.n3874 VSS.n3873 0.000963768
R12993 VSS.n3273 VSS.n3272 0.000962428
R12994 VSS.n3022 VSS.n3021 0.000951505
R12995 VSS.n2146 VSS.n2142 0.000951505
R12996 VSS.n3013 VSS.n2149 0.000951505
R12997 VSS.n3012 VSS.n2150 0.000951505
R12998 VSS.n3008 VSS.n2159 0.000951505
R12999 VSS.n3005 VSS.n2161 0.000951505
R13000 VSS.n2171 VSS.n2162 0.000951505
R13001 VSS.n2997 VSS.n2996 0.000951505
R13002 VSS.n2993 VSS.n2172 0.000951505
R13003 VSS.n2985 VSS.n2984 0.000951505
R13004 VSS.n2984 VSS.n2181 0.000951505
R13005 VSS.n2981 VSS.n2980 0.000951505
R13006 VSS.n2203 VSS.n2201 0.000951505
R13007 VSS.n2970 VSS.n2969 0.000951505
R13008 VSS.n2966 VSS.n2202 0.000951505
R13009 VSS.n2965 VSS.n2206 0.000951505
R13010 VSS.n2221 VSS.n2215 0.000951505
R13011 VSS.n2954 VSS.n2222 0.000951505
R13012 VSS.n2953 VSS.n2223 0.000951505
R13013 VSS.n2950 VSS.n2235 0.000951505
R13014 VSS.n3020 VSS.n3019 0.000951505
R13015 VSS.n2145 VSS.n2143 0.000951505
R13016 VSS.n3014 VSS.n2148 0.000951505
R13017 VSS.n3011 VSS.n2151 0.000951505
R13018 VSS.n2166 VSS.n2152 0.000951505
R13019 VSS.n2167 VSS.n2163 0.000951505
R13020 VSS.n3000 VSS.n2164 0.000951505
R13021 VSS.n2999 VSS.n2998 0.000951505
R13022 VSS.n2176 VSS.n2170 0.000951505
R13023 VSS.n2987 VSS.n2986 0.000951505
R13024 VSS.n2185 VSS.n2180 0.000951505
R13025 VSS.n2979 VSS.n2978 0.000951505
R13026 VSS.n2973 VSS.n2199 0.000951505
R13027 VSS.n2972 VSS.n2971 0.000951505
R13028 VSS.n2207 VSS.n2200 0.000951505
R13029 VSS.n2964 VSS.n2208 0.000951505
R13030 VSS.n2956 VSS.n2217 0.000951505
R13031 VSS.n2955 VSS.n2220 0.000951505
R13032 VSS.n2241 VSS.n2240 0.000951505
R13033 VSS.n2242 VSS.n2237 0.000951505
R13034 VSS.n2940 VSS.n2939 0.000951505
R13035 VSS.n2253 VSS.n2249 0.000951505
R13036 VSS.n2930 VSS.n2929 0.000951505
R13037 VSS.n2260 VSS.n2256 0.000951505
R13038 VSS.n2284 VSS.n2261 0.000951505
R13039 VSS.n2286 VSS.n2285 0.000951505
R13040 VSS.n2917 VSS.n2270 0.000951505
R13041 VSS.n2916 VSS.n2271 0.000951505
R13042 VSS.n2278 VSS.n2277 0.000951505
R13043 VSS.n2906 VSS.n2281 0.000951505
R13044 VSS.n2903 VSS.n2295 0.000951505
R13045 VSS.n2897 VSS.n2315 0.000951505
R13046 VSS.n2896 VSS.n2316 0.000951505
R13047 VSS.n2349 VSS.n2348 0.000951505
R13048 VSS.n2881 VSS.n2329 0.000951505
R13049 VSS.n2938 VSS.n2937 0.000951505
R13050 VSS.n2252 VSS.n2250 0.000951505
R13051 VSS.n2932 VSS.n2931 0.000951505
R13052 VSS.n2262 VSS.n2255 0.000951505
R13053 VSS.n2266 VSS.n2263 0.000951505
R13054 VSS.n2920 VSS.n2267 0.000951505
R13055 VSS.n2918 VSS.n2269 0.000951505
R13056 VSS.n2915 VSS.n2272 0.000951505
R13057 VSS.n2914 VSS.n2273 0.000951505
R13058 VSS.n2911 VSS.n2273 0.000951505
R13059 VSS.n2910 VSS.n2909 0.000951505
R13060 VSS.n2297 VSS.n2296 0.000951505
R13061 VSS.n2902 VSS.n2298 0.000951505
R13062 VSS.n2899 VSS.n2298 0.000951505
R13063 VSS.n2898 VSS.n2314 0.000951505
R13064 VSS.n2895 VSS.n2317 0.000951505
R13065 VSS.n2885 VSS.n2325 0.000951505
R13066 VSS.n2880 VSS.n2330 0.000951505
R13067 VSS.n2871 VSS.n2870 0.000951505
R13068 VSS.n2369 VSS.n2365 0.000951505
R13069 VSS.n2862 VSS.n2372 0.000951505
R13070 VSS.n2861 VSS.n2373 0.000951505
R13071 VSS.n2408 VSS.n2407 0.000951505
R13072 VSS.n2853 VSS.n2381 0.000951505
R13073 VSS.n2852 VSS.n2382 0.000951505
R13074 VSS.n2849 VSS.n2385 0.000951505
R13075 VSS.n2400 VSS.n2386 0.000951505
R13076 VSS.n2436 VSS.n2417 0.000951505
R13077 VSS.n2829 VSS.n2437 0.000951505
R13078 VSS.n2828 VSS.n2438 0.000951505
R13079 VSS.n2455 VSS.n2454 0.000951505
R13080 VSS.n2462 VSS.n2459 0.000951505
R13081 VSS.n2461 VSS.n2460 0.000951505
R13082 VSS.n2816 VSS.n2449 0.000951505
R13083 VSS.n2869 VSS.n2868 0.000951505
R13084 VSS.n2368 VSS.n2366 0.000951505
R13085 VSS.n2863 VSS.n2371 0.000951505
R13086 VSS.n2860 VSS.n2374 0.000951505
R13087 VSS.n2859 VSS.n2375 0.000951505
R13088 VSS.n2854 VSS.n2380 0.000951505
R13089 VSS.n2392 VSS.n2391 0.000951505
R13090 VSS.n2393 VSS.n2387 0.000951505
R13091 VSS.n2396 VSS.n2388 0.000951505
R13092 VSS.n2843 VSS.n2842 0.000951505
R13093 VSS.n2418 VSS.n2397 0.000951505
R13094 VSS.n2831 VSS.n2420 0.000951505
R13095 VSS.n2830 VSS.n2435 0.000951505
R13096 VSS.n2827 VSS.n2439 0.000951505
R13097 VSS.n2826 VSS.n2440 0.000951505
R13098 VSS.n2821 VSS.n2445 0.000951505
R13099 VSS.n2818 VSS.n2447 0.000951505
R13100 VSS.n2817 VSS.n2448 0.000951505
R13101 VSS.n2311 VSS.n2310 0.000950886
R13102 VSS.n1785 VSS.n1784 0.000920561
R13103 VSS.n3937 VSS.n3936 0.000920561
R13104 VSS.n3946 VSS.n3945 0.000920561
R13105 VSS.n3981 VSS.n3980 0.000920561
R13106 VSS.n3914 VSS.n3913 0.000920561
R13107 VSS.n3933 VSS.n3932 0.000920561
R13108 VSS.n3935 VSS.n3934 0.000920561
R13109 VSS.n3951 VSS.n3950 0.000920561
R13110 VSS.n3950 VSS.n3949 0.000920561
R13111 VSS.n3949 VSS.n3948 0.000920561
R13112 VSS.n3985 VSS.n3984 0.000920561
R13113 VSS.n3892 VSS.n3891 0.000920561
R13114 VSS.n3926 VSS.n3925 0.000920561
R13115 VSS.n3927 VSS.n3926 0.000920561
R13116 VSS.n3928 VSS.n3927 0.000920561
R13117 VSS.n3944 VSS.n3943 0.000920561
R13118 VSS.n3942 VSS.n3941 0.000920561
R13119 VSS.n1809 VSS.n1808 0.000914747
R13120 VSS.n1819 VSS.n1818 0.000914747
R13121 VSS.n7907 VSS.n7906 0.000914747
R13122 VSS.n3311 VSS.n3310 0.000904624
R13123 VSS.n2609 VSS.n2597 0.0009
R13124 VSS.n2721 VSS.n2578 0.000893013
R13125 VSS.n2720 VSS.n2719 0.000893013
R13126 VSS.n2590 VSS.n2587 0.000893013
R13127 VSS.n2710 VSS.n2709 0.000893013
R13128 VSS.n2705 VSS.n2704 0.000893013
R13129 VSS.n2600 VSS.n2594 0.000893013
R13130 VSS.n2696 VSS.n2695 0.000893013
R13131 VSS.n2691 VSS.n2604 0.000893013
R13132 VSS.n2611 VSS.n2605 0.000893013
R13133 VSS.n2683 VSS.n2614 0.000893013
R13134 VSS.n2682 VSS.n2615 0.000893013
R13135 VSS.n2679 VSS.n2618 0.000893013
R13136 VSS.n2678 VSS.n2619 0.000893013
R13137 VSS.n2645 VSS.n2644 0.000893013
R13138 VSS.n2657 VSS.n2654 0.000893013
R13139 VSS.n2661 VSS.n2658 0.000893013
R13140 VSS.n2582 VSS.n2580 0.000893013
R13141 VSS.n2718 VSS.n2717 0.000893013
R13142 VSS.n2717 VSS.n2581 0.000893013
R13143 VSS.n2713 VSS.n2585 0.000893013
R13144 VSS.n2712 VSS.n2711 0.000893013
R13145 VSS.n2703 VSS.n2702 0.000893013
R13146 VSS.n2598 VSS.n2595 0.000893013
R13147 VSS.n2698 VSS.n2697 0.000893013
R13148 VSS.n2608 VSS.n2606 0.000893013
R13149 VSS.n2686 VSS.n2607 0.000893013
R13150 VSS.n2684 VSS.n2613 0.000893013
R13151 VSS.n2637 VSS.n2634 0.000893013
R13152 VSS.n2639 VSS.n2638 0.000893013
R13153 VSS.n2677 VSS.n2620 0.000893013
R13154 VSS.n2676 VSS.n2621 0.000893013
R13155 VSS.n2663 VSS.n2655 0.000893013
R13156 VSS.n3682 VSS.n3681 0.000892442
R13157 VSS.n3621 VSS.n3620 0.000892442
R13158 VSS.n3622 VSS.n3621 0.000892442
R13159 VSS.n3624 VSS.n3623 0.000892442
R13160 VSS.n3627 VSS.n3626 0.000892442
R13161 VSS.n3629 VSS.n3628 0.000892442
R13162 VSS.n3664 VSS.n3663 0.000892442
R13163 VSS.n3662 VSS.n3661 0.000892442
R13164 VSS.n3659 VSS.n3658 0.000892442
R13165 VSS.n3657 VSS.n3656 0.000892442
R13166 VSS.n3655 VSS.n3654 0.000892442
R13167 VSS.n3651 VSS.n3650 0.000892442
R13168 VSS.n3649 VSS.n3648 0.000892442
R13169 VSS.n3647 VSS.n3646 0.000892442
R13170 VSS.n3645 VSS.n3644 0.000892442
R13171 VSS.n3643 VSS.n3642 0.000892442
R13172 VSS.n3640 VSS.n3639 0.000892442
R13173 VSS.n3638 VSS.n3637 0.000892442
R13174 VSS.n3636 VSS.n3635 0.000892442
R13175 VSS.n3632 VSS.n3631 0.000892442
R13176 VSS.n3611 VSS.n3610 0.000892442
R13177 VSS.n3616 VSS.n3615 0.000892442
R13178 VSS.n3618 VSS.n3617 0.000892442
R13179 VSS.n3737 VSS.n3736 0.000892442
R13180 VSS.n3736 VSS.n3735 0.000892442
R13181 VSS.n3734 VSS.n3733 0.000892442
R13182 VSS.n3731 VSS.n3730 0.000892442
R13183 VSS.n3729 VSS.n3728 0.000892442
R13184 VSS.n3727 VSS.n3726 0.000892442
R13185 VSS.n3721 VSS.n3720 0.000892442
R13186 VSS.n3719 VSS.n3718 0.000892442
R13187 VSS.n3717 VSS.n3716 0.000892442
R13188 VSS.n3715 VSS.n3714 0.000892442
R13189 VSS.n3712 VSS.n3711 0.000892442
R13190 VSS.n3710 VSS.n3709 0.000892442
R13191 VSS.n3708 VSS.n3707 0.000892442
R13192 VSS.n3704 VSS.n3703 0.000892442
R13193 VSS.n3582 VSS.n3581 0.000892442
R13194 VSS.n3580 VSS.n3579 0.000892442
R13195 VSS.n3527 VSS.n3526 0.000892442
R13196 VSS.n3512 VSS.n3511 0.000892442
R13197 VSS.n3514 VSS.n3513 0.000892442
R13198 VSS.n3516 VSS.n3515 0.000892442
R13199 VSS.n3492 VSS.n3491 0.000892442
R13200 VSS.n3490 VSS.n3489 0.000892442
R13201 VSS.n3488 VSS.n3487 0.000892442
R13202 VSS.n3471 VSS.n3470 0.000892442
R13203 VSS.n3473 VSS.n3472 0.000892442
R13204 VSS.n3475 VSS.n3474 0.000892442
R13205 VSS.n3452 VSS.n3451 0.000892442
R13206 VSS.n3457 VSS.n3456 0.000892442
R13207 VSS.n3455 VSS.n3454 0.000892442
R13208 VSS.n3437 VSS.n3436 0.000892442
R13209 VSS.n3435 VSS.n3434 0.000892442
R13210 VSS.n3525 VSS.n3524 0.000892442
R13211 VSS.n3506 VSS.n3505 0.000892442
R13212 VSS.n3508 VSS.n3507 0.000892442
R13213 VSS.n3510 VSS.n3509 0.000892442
R13214 VSS.n3499 VSS.n3498 0.000892442
R13215 VSS.n3497 VSS.n3496 0.000892442
R13216 VSS.n3495 VSS.n3494 0.000892442
R13217 VSS.n3467 VSS.n3466 0.000892442
R13218 VSS.n3469 VSS.n3468 0.000892442
R13219 VSS.n3478 VSS.n3477 0.000892442
R13220 VSS.n3445 VSS.n3444 0.000892442
R13221 VSS.n3450 VSS.n3449 0.000892442
R13222 VSS.n3448 VSS.n3447 0.000892442
R13223 VSS.n3432 VSS.n3431 0.000892442
R13224 VSS.n3430 VSS.n3429 0.000892442
R13225 VSS.n3419 VSS.n3418 0.000892442
R13226 VSS.n3415 VSS.n3414 0.000892442
R13227 VSS.n3402 VSS.n3401 0.000892442
R13228 VSS.n3400 VSS.n3399 0.000892442
R13229 VSS.n3360 VSS.n3359 0.000892442
R13230 VSS.n3348 VSS.n3347 0.000892442
R13231 VSS.n3350 VSS.n3349 0.000892442
R13232 VSS.n3335 VSS.n3334 0.000892442
R13233 VSS.n3333 VSS.n3332 0.000892442
R13234 VSS.n3331 VSS.n3330 0.000892442
R13235 VSS.n3319 VSS.n3318 0.000892442
R13236 VSS.n3317 VSS.n3316 0.000892442
R13237 VSS.n3298 VSS.n3297 0.000892442
R13238 VSS.n3279 VSS.n3278 0.000892442
R13239 VSS.n3277 VSS.n3276 0.000892442
R13240 VSS.n3264 VSS.n3263 0.000892442
R13241 VSS.n3262 VSS.n3261 0.000892442
R13242 VSS.n3251 VSS.n3250 0.000892442
R13243 VSS.n3249 VSS.n3248 0.000892442
R13244 VSS.n3370 VSS.n3369 0.000892442
R13245 VSS.n3368 VSS.n3367 0.000892442
R13246 VSS.n3358 VSS.n3357 0.000892442
R13247 VSS.n3344 VSS.n3343 0.000892442
R13248 VSS.n3346 VSS.n3345 0.000892442
R13249 VSS.n3340 VSS.n3339 0.000892442
R13250 VSS.n3338 VSS.n3337 0.000892442
R13251 VSS.n3315 VSS.n3314 0.000892442
R13252 VSS.n3324 VSS.n3323 0.000892442
R13253 VSS.n3322 VSS.n3321 0.000892442
R13254 VSS.n3304 VSS.n3303 0.000892442
R13255 VSS.n3294 VSS.n3293 0.000892442
R13256 VSS.n3292 VSS.n3291 0.000892442
R13257 VSS.n3284 VSS.n3283 0.000892442
R13258 VSS.n3282 VSS.n3281 0.000892442
R13259 VSS.n3256 VSS.n3255 0.000892442
R13260 VSS.n3254 VSS.n3253 0.000892442
R13261 VSS.n3213 VSS.n3212 0.000892442
R13262 VSS.n3217 VSS.n3216 0.000892442
R13263 VSS.n3215 VSS.n3214 0.000892442
R13264 VSS.n3204 VSS.n3203 0.000892442
R13265 VSS.n3202 VSS.n3201 0.000892442
R13266 VSS.n3188 VSS.n3187 0.000892442
R13267 VSS.n3178 VSS.n3177 0.000892442
R13268 VSS.n3180 VSS.n3179 0.000892442
R13269 VSS.n3166 VSS.n3165 0.000892442
R13270 VSS.n3165 VSS.n3164 0.000892442
R13271 VSS.n3153 VSS.n3152 0.000892442
R13272 VSS.n3155 VSS.n3154 0.000892442
R13273 VSS.n3137 VSS.n3136 0.000892442
R13274 VSS.n3139 VSS.n3138 0.000892442
R13275 VSS.n3141 VSS.n3140 0.000892442
R13276 VSS.n3117 VSS.n3116 0.000892442
R13277 VSS.n3115 VSS.n3114 0.000892442
R13278 VSS.n3113 VSS.n3112 0.000892442
R13279 VSS.n3065 VSS.n3064 0.000892442
R13280 VSS.n3211 VSS.n3210 0.000892442
R13281 VSS.n3222 VSS.n3221 0.000892442
R13282 VSS.n3220 VSS.n3219 0.000892442
R13283 VSS.n3200 VSS.n3199 0.000892442
R13284 VSS.n3198 VSS.n3197 0.000892442
R13285 VSS.n3192 VSS.n3191 0.000892442
R13286 VSS.n3176 VSS.n3175 0.000892442
R13287 VSS.n3171 VSS.n3170 0.000892442
R13288 VSS.n3169 VSS.n3168 0.000892442
R13289 VSS.n3151 VSS.n3150 0.000892442
R13290 VSS.n3158 VSS.n3157 0.000892442
R13291 VSS.n3131 VSS.n3130 0.000892442
R13292 VSS.n3133 VSS.n3132 0.000892442
R13293 VSS.n3135 VSS.n3134 0.000892442
R13294 VSS.n3124 VSS.n3123 0.000892442
R13295 VSS.n3122 VSS.n3121 0.000892442
R13296 VSS.n3120 VSS.n3119 0.000892442
R13297 VSS.n3063 VSS.n3062 0.000892442
R13298 VSS.n2806 VSS.n2805 0.000892442
R13299 VSS.n2480 VSS.n2474 0.000892442
R13300 VSS.n2495 VSS.n2487 0.000892442
R13301 VSS.n2496 VSS.n2494 0.000892442
R13302 VSS.n2783 VSS.n2499 0.000892442
R13303 VSS.n2780 VSS.n2501 0.000892442
R13304 VSS.n2779 VSS.n2502 0.000892442
R13305 VSS.n2771 VSS.n2514 0.000892442
R13306 VSS.n2771 VSS.n2770 0.000892442
R13307 VSS.n2525 VSS.n2515 0.000892442
R13308 VSS.n2544 VSS.n2526 0.000892442
R13309 VSS.n2758 VSS.n2757 0.000892442
R13310 VSS.n2754 VSS.n2545 0.000892442
R13311 VSS.n2753 VSS.n2547 0.000892442
R13312 VSS.n2745 VSS.n2558 0.000892442
R13313 VSS.n2742 VSS.n2741 0.000892442
R13314 VSS.n2565 VSS.n2560 0.000892442
R13315 VSS.n2733 VSS.n2732 0.000892442
R13316 VSS.n2804 VSS.n2803 0.000892442
R13317 VSS.n2476 VSS.n2475 0.000892442
R13318 VSS.n2798 VSS.n2797 0.000892442
R13319 VSS.n2488 VSS.n2479 0.000892442
R13320 VSS.n2491 VSS.n2489 0.000892442
R13321 VSS.n2786 VSS.n2492 0.000892442
R13322 VSS.n2507 VSS.n2493 0.000892442
R13323 VSS.n2509 VSS.n2508 0.000892442
R13324 VSS.n2778 VSS.n2503 0.000892442
R13325 VSS.n2773 VSS.n2772 0.000892442
R13326 VSS.n2772 VSS.n2513 0.000892442
R13327 VSS.n2528 VSS.n2527 0.000892442
R13328 VSS.n2761 VSS.n2529 0.000892442
R13329 VSS.n2760 VSS.n2759 0.000892442
R13330 VSS.n2548 VSS.n2543 0.000892442
R13331 VSS.n2752 VSS.n2549 0.000892442
R13332 VSS.n2561 VSS.n2555 0.000892442
R13333 VSS.n2740 VSS.n2739 0.000892442
R13334 VSS.n2736 VSS.n2562 0.000892442
R13335 VSS.n2735 VSS.n2734 0.000892442
R13336 VSS.n1884 VSS.n1883 0.000892442
R13337 VSS.n1890 VSS.n1889 0.000892442
R13338 VSS.n1905 VSS.n1904 0.000892442
R13339 VSS.n1918 VSS.n1917 0.000892442
R13340 VSS.n1919 VSS.n1918 0.000892442
R13341 VSS.n1921 VSS.n1920 0.000892442
R13342 VSS.n3870 VSS.n3869 0.000892442
R13343 VSS.n3868 VSS.n3867 0.000892442
R13344 VSS.n3866 VSS.n3865 0.000892442
R13345 VSS.n3849 VSS.n3848 0.000892442
R13346 VSS.n3827 VSS.n3826 0.000892442
R13347 VSS.n3825 VSS.n3824 0.000892442
R13348 VSS.n3814 VSS.n3813 0.000892442
R13349 VSS.n3816 VSS.n3815 0.000892442
R13350 VSS.n3801 VSS.n3800 0.000892442
R13351 VSS.n3799 VSS.n3798 0.000892442
R13352 VSS.n3749 VSS.n3748 0.000892442
R13353 VSS.n1893 VSS.n1892 0.000892442
R13354 VSS.n1900 VSS.n1899 0.000892442
R13355 VSS.n1902 VSS.n1901 0.000892442
R13356 VSS.n1913 VSS.n1912 0.000892442
R13357 VSS.n1914 VSS.n1913 0.000892442
R13358 VSS.n1916 VSS.n1915 0.000892442
R13359 VSS.n3864 VSS.n3863 0.000892442
R13360 VSS.n3862 VSS.n3861 0.000892442
R13361 VSS.n3847 VSS.n3846 0.000892442
R13362 VSS.n3832 VSS.n3831 0.000892442
R13363 VSS.n3830 VSS.n3829 0.000892442
R13364 VSS.n3810 VSS.n3809 0.000892442
R13365 VSS.n3812 VSS.n3811 0.000892442
R13366 VSS.n3806 VSS.n3805 0.000892442
R13367 VSS.n3804 VSS.n3803 0.000892442
R13368 VSS.n3747 VSS.n3746 0.000892442
R13369 VSS.n2913 VSS.n2912 0.000886473
R13370 VSS.n2901 VSS.n2900 0.000886473
R13371 VSS.n4127 VSS.n4120 0.000868349
R13372 VSS.n2774 VSS.n2512 0.000848837
R13373 VSS.n1910 VSS.n1909 0.000847826
R13374 VSS.n2687 VSS.n2610 0.000842857
R13375 VSS.n2976 VSS.n2975 0.000834448
R13376 VSS.n2310 VSS.n2276 0.000822061
R13377 VSS.n2820 VSS.n2442 0.000814465
R13378 VSS.n2352 VSS.n2333 0.000801003
R13379 VSS.n2341 VSS.n2335 0.000801003
R13380 VSS.n2351 VSS.n2344 0.000801003
R13381 VSS.n2346 VSS.n2345 0.000801003
R13382 VSS.n2908 VSS.n2907 0.000801003
R13383 VSS.n2338 VSS.n2337 0.000801003
R13384 VSS.n2340 VSS.n2339 0.000801003
R13385 VSS.n2324 VSS.n2323 0.000801003
R13386 VSS.n2347 VSS.n2328 0.000801003
R13387 VSS.n2883 VSS.n2882 0.000801003
R13388 VSS.n2909 VSS.n2279 0.000801003
R13389 VSS.n2894 VSS.n2318 0.000801003
R13390 VSS.n2336 VSS.n2321 0.000801003
R13391 VSS.n2889 VSS.n2888 0.000801003
R13392 VSS.n2884 VSS.n2327 0.000801003
R13393 VSS.n2357 VSS.n2356 0.000801003
R13394 VSS.n2841 VSS.n2840 0.000801003
R13395 VSS.n2842 VSS.n2397 0.000801003
R13396 VSS.n2775 VSS.n2774 0.000790698
R13397 VSS.n3302 VSS.n3289 0.000789017
R13398 VSS.n3417 VSS.n3408 0.000789017
R13399 VSS.n4035 VSS.n4034 0.00077907
R13400 VSS.n2211 VSS.n2210 0.000767559
R13401 VSS.n2958 VSS.n2218 0.000767559
R13402 VSS.n2239 VSS.n2219 0.000767559
R13403 VSS.n3625 VSS.n3624 0.000761628
R13404 VSS.n3613 VSS.n3612 0.000761628
R13405 VSS.n3733 VSS.n3732 0.000761628
R13406 VSS.n3724 VSS.n3723 0.000761628
R13407 VSS.n3547 VSS.n3546 0.000761628
R13408 VSS.n3581 VSS.n3580 0.000761628
R13409 VSS.n3422 VSS.n3421 0.000761628
R13410 VSS.n3412 VSS.n3411 0.000761628
R13411 VSS.n3536 VSS.n3535 0.000761628
R13412 VSS.n3479 VSS.n3478 0.000761628
R13413 VSS.n3431 VSS.n3430 0.000761628
R13414 VSS.n3416 VSS.n3415 0.000761628
R13415 VSS.n3382 VSS.n3381 0.000761628
R13416 VSS.n3307 VSS.n3306 0.000761628
R13417 VSS.n3300 VSS.n3299 0.000761628
R13418 VSS.n3263 VSS.n3262 0.000761628
R13419 VSS.n3301 VSS.n3294 0.000761628
R13420 VSS.n3268 VSS.n3267 0.000761628
R13421 VSS.n2794 VSS.n2793 0.000761628
R13422 VSS.n2795 VSS.n2482 0.000761628
R13423 VSS.n3853 VSS.n3852 0.000761628
R13424 VSS.n3851 VSS.n3850 0.000761628
R13425 VSS.n3844 VSS.n3843 0.000761628
R13426 VSS.n2813 VSS.n2446 0.000751572
R13427 VSS.n4086 VSS.n4085 0.000751397
R13428 VSS.n4110 VSS.n4103 0.000751397
R13429 VSS.n4080 VSS.n4051 0.000751397
R13430 VSS.n4079 VSS.n4078 0.000751397
R13431 VSS.n4069 VSS.n4068 0.000751397
R13432 VSS.n4067 VSS.n4066 0.000751397
R13433 VSS.n4060 VSS.n4059 0.000751397
R13434 VSS.n4057 VSS.n4056 0.000751397
R13435 VSS.n4055 VSS.n4054 0.000751397
R13436 VSS.n4507 VSS.n4506 0.00074
R13437 VSS.n2764 VSS.n2530 0.000732558
R13438 VSS.n2552 VSS.n2542 0.000732558
R13439 VSS.n2750 VSS.n2749 0.000732558
R13440 VSS.n2738 VSS.n2554 0.000732558
R13441 VSS.n3146 VSS.n3145 0.000732558
R13442 VSS.n3129 VSS.n3126 0.000732558
R13443 VSS.n3110 VSS.n3109 0.000732558
R13444 VSS.n3821 VSS.n3820 0.000731884
R13445 VSS.n3819 VSS.n3808 0.000731884
R13446 VSS.n3797 VSS.n3796 0.000731884
R13447 VSS.n3329 VSS.n3328 0.000731214
R13448 VSS.n3310 VSS.n3309 0.000731214
R13449 VSS.n3260 VSS.n3259 0.000731214
R13450 VSS.n3532 VSS.n3531 0.000731214
R13451 VSS.n3425 VSS.n3424 0.000731214
R13452 VSS.n2583 VSS.n2573 0.000728571
R13453 VSS.n2641 VSS.n2640 0.000728571
R13454 VSS.n2674 VSS.n2642 0.000728571
R13455 VSS.n6980 VSS.n6979 0.000713777
R13456 VSS.n6982 VSS.n6981 0.000713777
R13457 VSS.n6984 VSS.n6983 0.000713777
R13458 VSS.n7301 VSS.n7300 0.000713777
R13459 VSS.n3971 VSS.n3970 0.00071028
R13460 VSS.n3895 VSS.n3894 0.00071028
R13461 VSS.n3972 VSS.n3968 0.00071028
R13462 VSS.n3901 VSS.n3900 0.00071028
R13463 VSS.n3918 VSS.n3917 0.00071028
R13464 VSS.n3954 VSS.n3940 0.00071028
R13465 VSS.n3954 VSS.n3953 0.00071028
R13466 VSS.n3943 VSS.n3942 0.00071028
R13467 VSS.n3974 VSS.n3973 0.00071028
R13468 VSS.n3987 VSS.n3986 0.00071028
R13469 VSS.n1831 VSS.n1830 0.000707373
R13470 VSS.n1839 VSS.n1838 0.000707373
R13471 VSS.n1841 VSS.n1840 0.000707373
R13472 VSS.n1851 VSS.n1850 0.000707373
R13473 VSS.n1853 VSS.n1852 0.000707373
R13474 VSS.n1862 VSS.n1860 0.000707373
R13475 VSS.n3038 VSS.n3037 0.000702532
R13476 VSS.n3035 VSS.n3034 0.000702532
R13477 VSS.n3032 VSS.n3031 0.000702532
R13478 VSS.n3924 VSS.n3923 0.00068648
R13479 VSS.n3958 VSS.n3957 0.00068648
R13480 VSS.n4032 VSS.n4031 0.000686047
R13481 VSS.n3738 VSS.n3608 0.000674419
R13482 VSS.n3598 VSS.n3597 0.000674419
R13483 VSS.n2716 VSS.n2715 0.000671429
R13484 VSS.n2636 VSS.n2633 0.000671429
R13485 VSS.n1991 VSS.n1990 0.000655172
R13486 VSS.n2003 VSS.n2002 0.000655172
R13487 VSS.n2028 VSS.n2027 0.000655172
R13488 VSS.n2018 VSS.n2017 0.000655172
R13489 VSS.n2966 VSS.n2965 0.000650502
R13490 VSS.n2954 VSS.n2953 0.000650502
R13491 VSS.n2208 VSS.n2207 0.000650502
R13492 VSS.n2240 VSS.n2220 0.000650502
R13493 VSS.n2905 VSS.n2280 0.000650502
R13494 VSS.n2907 VSS.n2906 0.000650502
R13495 VSS.n2339 VSS.n2338 0.000650502
R13496 VSS.n2883 VSS.n2328 0.000650502
R13497 VSS.n2336 VSS.n2318 0.000650502
R13498 VSS.n2356 VSS.n2327 0.000650502
R13499 VSS.n2841 VSS.n2398 0.000650502
R13500 VSS.n2840 VSS.n2839 0.000650502
R13501 VSS.n1137 VSS.n1136 0.000643312
R13502 VSS.n2679 VSS.n2678 0.000631004
R13503 VSS.n2658 VSS.n2657 0.000631004
R13504 VSS.n2638 VSS.n2620 0.000631004
R13505 VSS.n2663 VSS.n2662 0.000631004
R13506 VSS.n3652 VSS.n3651 0.000630814
R13507 VSS.n3614 VSS.n3613 0.000630814
R13508 VSS.n3723 VSS.n3722 0.000630814
R13509 VSS.n3545 VSS.n3544 0.000630814
R13510 VSS.n3422 VSS.n3420 0.000630814
R13511 VSS.n3412 VSS.n3409 0.000630814
R13512 VSS.n3537 VSS.n3536 0.000630814
R13513 VSS.n3535 VSS.n3534 0.000630814
R13514 VSS.n3459 VSS.n3445 0.000630814
R13515 VSS.n3423 VSS.n3419 0.000630814
R13516 VSS.n3380 VSS.n3379 0.000630814
R13517 VSS.n3307 VSS.n3305 0.000630814
R13518 VSS.n3300 VSS.n3295 0.000630814
R13519 VSS.n3308 VSS.n3304 0.000630814
R13520 VSS.n3269 VSS.n3268 0.000630814
R13521 VSS.n3267 VSS.n3266 0.000630814
R13522 VSS.n3140 VSS.n3139 0.000630814
R13523 VSS.n3114 VSS.n3113 0.000630814
R13524 VSS.n3134 VSS.n3133 0.000630814
R13525 VSS.n3121 VSS.n3120 0.000630814
R13526 VSS.n2796 VSS.n2795 0.000630814
R13527 VSS.n2486 VSS.n2482 0.000630814
R13528 VSS.n2757 VSS.n2545 0.000630814
R13529 VSS.n2742 VSS.n2558 0.000630814
R13530 VSS.n2759 VSS.n2543 0.000630814
R13531 VSS.n2740 VSS.n2561 0.000630814
R13532 VSS.n3776 VSS.n3775 0.000630814
R13533 VSS.n3852 VSS.n3851 0.000630814
R13534 VSS.n3815 VSS.n3814 0.000630814
R13535 VSS.n3800 VSS.n3799 0.000630814
R13536 VSS.n3845 VSS.n3844 0.000630814
R13537 VSS.n3843 VSS.n3842 0.000630814
R13538 VSS.n3811 VSS.n3810 0.000630814
R13539 VSS.n3805 VSS.n3804 0.000630814
R13540 VSS.n2893 VSS.n2892 0.000628824
R13541 VSS.n2887 VSS.n2320 0.000628824
R13542 VSS.n2358 VSS.n2326 0.000628824
R13543 VSS.n2833 VSS.n2433 0.000625786
R13544 VSS.n3607 VSS.n3606 0.000616279
R13545 VSS.n3601 VSS.n3600 0.000616279
R13546 VSS.n3839 VSS.n3838 0.000615942
R13547 VSS.n3480 VSS.n3465 0.000615607
R13548 VSS.n3427 VSS.n3426 0.000615607
R13549 VSS.n3903 VSS.n3902 0.00059324
R13550 VSS.n3920 VSS.n3919 0.00059324
R13551 VSS.n3931 VSS.n3930 0.00059324
R13552 VSS.n3955 VSS.n3931 0.00059324
R13553 VSS.n3956 VSS.n3955 0.00059324
R13554 VSS.n3976 VSS.n3975 0.00059324
R13555 VSS.n3989 VSS.n3988 0.00059324
R13556 VSS.n4050 VSS.n4049 0.000593023
R13557 VSS.n4048 VSS.n4047 0.000593023
R13558 VSS.n4042 VSS.n4041 0.000593023
R13559 VSS.n4040 VSS.n4039 0.000593023
R13560 VSS.n4033 VSS.n4032 0.000593023
R13561 VSS.n4031 VSS.n4030 0.000593023
R13562 VSS.n3998 VSS.n3997 0.000592166
R13563 VSS.n4003 VSS.n4002 0.000592166
R13564 VSS.n4005 VSS.n4004 0.000592166
R13565 VSS.n4012 VSS.n4011 0.000592166
R13566 VSS.n4014 VSS.n4013 0.000592166
R13567 VSS.n4019 VSS.n4018 0.000592166
R13568 VSS.n3148 VSS.n3147 0.00055814
R13569 VSS.n3742 VSS.n3741 0.00055814
R13570 VSS.n3482 VSS.n3481 0.000557804
R13571 VSS.n3461 VSS.n3460 0.000557804
R13572 VSS.n3041 VSS.n3040 0.000550633
R13573 PFD_T2_0.INV_mag_1.OUT.n0 PFD_T2_0.INV_mag_1.OUT.t9 29.3524
R13574 PFD_T2_0.INV_mag_1.OUT.n2 PFD_T2_0.INV_mag_1.OUT.t4 23.3605
R13575 PFD_T2_0.INV_mag_1.OUT.n3 PFD_T2_0.INV_mag_1.OUT.n0 16.8716
R13576 PFD_T2_0.INV_mag_1.OUT.n4 PFD_T2_0.INV_mag_1.OUT.t3 12.4111
R13577 PFD_T2_0.INV_mag_1.OUT.n0 PFD_T2_0.INV_mag_1.OUT.t6 9.0525
R13578 PFD_T2_0.INV_mag_1.OUT.n3 PFD_T2_0.INV_mag_1.OUT.t8 9.0525
R13579 PFD_T2_0.INV_mag_1.OUT.t3 PFD_T2_0.INV_mag_1.OUT.n3 9.0525
R13580 PFD_T2_0.INV_mag_1.OUT.n0 PFD_T2_0.INV_mag_1.OUT.t5 9.0525
R13581 PFD_T2_0.INV_mag_1.OUT.n2 PFD_T2_0.INV_mag_1.OUT.t7 8.7605
R13582 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.OUT.n5 6.74425
R13583 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.OUT.n1 5.41686
R13584 PFD_T2_0.INV_mag_1.OUT.n7 PFD_T2_0.INV_mag_1.OUT.t1 3.6405
R13585 PFD_T2_0.INV_mag_1.OUT.n7 PFD_T2_0.INV_mag_1.OUT.n6 3.6405
R13586 PFD_T2_0.INV_mag_1.OUT.n1 PFD_T2_0.INV_mag_1.OUT.n2 9.03264
R13587 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_1.OUT.n7 3.34789
R13588 PFD_T2_0.INV_mag_1.OUT.n1 PFD_T2_0.INV_mag_1.OUT.n4 1.1347
R13589 PFD_T2_0.Buffer_V_2_0.IN.n1 PFD_T2_0.Buffer_V_2_0.IN.t11 13.2135
R13590 PFD_T2_0.Buffer_V_2_0.IN.n2 PFD_T2_0.Buffer_V_2_0.IN.n1 12.5844
R13591 PFD_T2_0.Buffer_V_2_0.IN.n1 PFD_T2_0.Buffer_V_2_0.IN.t13 9.8555
R13592 PFD_T2_0.Buffer_V_2_0.IN.n2 PFD_T2_0.Buffer_V_2_0.IN.t12 9.71737
R13593 PFD_T2_0.Buffer_V_2_0.IN.n16 PFD_T2_0.Buffer_V_2_0.IN.n7 6.60246
R13594 PFD_T2_0.Buffer_V_2_0.IN.n0 PFD_T2_0.Buffer_V_2_0.IN.n18 4.10693
R13595 PFD_T2_0.Buffer_V_2_0.IN.n0 PFD_T2_0.Buffer_V_2_0.IN.n2 3.78915
R13596 PFD_T2_0.Buffer_V_2_0.IN.n11 PFD_T2_0.Buffer_V_2_0.IN.t5 3.6405
R13597 PFD_T2_0.Buffer_V_2_0.IN.n11 PFD_T2_0.Buffer_V_2_0.IN.n10 3.6405
R13598 PFD_T2_0.Buffer_V_2_0.IN.n13 PFD_T2_0.Buffer_V_2_0.IN.t6 3.6405
R13599 PFD_T2_0.Buffer_V_2_0.IN.n13 PFD_T2_0.Buffer_V_2_0.IN.n12 3.6405
R13600 PFD_T2_0.Buffer_V_2_0.IN.n14 PFD_T2_0.Buffer_V_2_0.IN.n11 3.54941
R13601 PFD_T2_0.Buffer_V_2_0.IN.n15 PFD_T2_0.Buffer_V_2_0.IN.n9 3.33833
R13602 PFD_T2_0.Buffer_V_2_0.IN.n17 PFD_T2_0.Buffer_V_2_0.IN.n6 3.33833
R13603 PFD_T2_0.Buffer_V_2_0.IN.n9 PFD_T2_0.Buffer_V_2_0.IN.t2 3.2765
R13604 PFD_T2_0.Buffer_V_2_0.IN.n9 PFD_T2_0.Buffer_V_2_0.IN.n8 3.2765
R13605 PFD_T2_0.Buffer_V_2_0.IN.n4 PFD_T2_0.Buffer_V_2_0.IN.t10 3.2765
R13606 PFD_T2_0.Buffer_V_2_0.IN.n4 PFD_T2_0.Buffer_V_2_0.IN.n3 3.2765
R13607 PFD_T2_0.Buffer_V_2_0.IN.n6 PFD_T2_0.Buffer_V_2_0.IN.t9 3.2765
R13608 PFD_T2_0.Buffer_V_2_0.IN.n6 PFD_T2_0.Buffer_V_2_0.IN.n5 3.2765
R13609 PFD_T2_0.Buffer_V_2_0.IN.n14 PFD_T2_0.Buffer_V_2_0.IN.n13 2.78441
R13610 PFD_T2_0.Buffer_V_2_0.IN.n18 PFD_T2_0.Buffer_V_2_0.IN.n4 1.8538
R13611 PFD_T2_0.Buffer_V_2_0.IN.n18 PFD_T2_0.Buffer_V_2_0.IN.n17 0.78641
R13612 PFD_T2_0.Buffer_V_2_0.IN.n16 PFD_T2_0.Buffer_V_2_0.IN.n15 0.524848
R13613 PFD_T2_0.Buffer_V_2_0.IN.n15 PFD_T2_0.Buffer_V_2_0.IN.n14 0.358543
R13614 PFD_T2_0.Buffer_V_2_0.IN.n17 PFD_T2_0.Buffer_V_2_0.IN.n16 0.274413
R13615 PFD_T2_0.Buffer_V_2_0.IN PFD_T2_0.Buffer_V_2_0.IN.n0 0.264033
R13616 PFD_T2_0.INV_mag_0.IN.n22 PFD_T2_0.INV_mag_0.IN.t2 219.017
R13617 PFD_T2_0.INV_mag_0.IN.n3 PFD_T2_0.INV_mag_0.IN.t28 116.993
R13618 PFD_T2_0.INV_mag_0.IN.n25 PFD_T2_0.INV_mag_0.IN.t23 33.8279
R13619 PFD_T2_0.INV_mag_0.IN.n26 PFD_T2_0.INV_mag_0.IN.n25 30.2144
R13620 PFD_T2_0.INV_mag_0.IN.t20 PFD_T2_0.INV_mag_0.IN.n1 25.0458
R13621 PFD_T2_0.INV_mag_0.IN.n28 PFD_T2_0.INV_mag_0.IN.n27 16.5048
R13622 PFD_T2_0.INV_mag_0.IN.n29 PFD_T2_0.INV_mag_0.IN.n28 16.5048
R13623 PFD_T2_0.INV_mag_0.IN.n1 PFD_T2_0.INV_mag_0.IN.t24 15.3305
R13624 PFD_T2_0.INV_mag_0.IN.n4 PFD_T2_0.INV_mag_0.IN.t25 15.2644
R13625 PFD_T2_0.INV_mag_0.IN.n1 PFD_T2_0.INV_mag_0.IN.n26 12.8616
R13626 PFD_T2_0.INV_mag_0.IN.n4 PFD_T2_0.INV_mag_0.IN.t17 12.7717
R13627 PFD_T2_0.INV_mag_0.IN.n0 PFD_T2_0.INV_mag_0.IN.t20 12.0785
R13628 PFD_T2_0.INV_mag_0.IN.t18 PFD_T2_0.INV_mag_0.IN.n3 11.3197
R13629 PFD_T2_0.INV_mag_0.IN.n22 PFD_T2_0.INV_mag_0.IN.t4 10.8543
R13630 PFD_T2_0.INV_mag_0.IN.n3 PFD_T2_0.INV_mag_0.IN.t29 10.2935
R13631 PFD_T2_0.INV_mag_0.IN.n27 PFD_T2_0.INV_mag_0.IN.t21 9.4175
R13632 PFD_T2_0.INV_mag_0.IN.n28 PFD_T2_0.INV_mag_0.IN.t31 9.4175
R13633 PFD_T2_0.INV_mag_0.IN.t24 PFD_T2_0.INV_mag_0.IN.n29 9.4175
R13634 PFD_T2_0.INV_mag_0.IN.n27 PFD_T2_0.INV_mag_0.IN.t33 9.1985
R13635 PFD_T2_0.INV_mag_0.IN.n28 PFD_T2_0.INV_mag_0.IN.t26 9.1985
R13636 PFD_T2_0.INV_mag_0.IN.n29 PFD_T2_0.INV_mag_0.IN.t19 9.1985
R13637 PFD_T2_0.INV_mag_0.IN.n30 PFD_T2_0.INV_mag_0.IN.n4 8.99637
R13638 PFD_T2_0.INV_mag_0.IN.n1 PFD_T2_0.INV_mag_0.IN.t32 8.05323
R13639 PFD_T2_0.INV_mag_0.IN.n13 PFD_T2_0.INV_mag_0.IN.n12 6.76657
R13640 PFD_T2_0.INV_mag_0.IN.n2 PFD_T2_0.INV_mag_0.IN.n21 6.46389
R13641 PFD_T2_0.INV_mag_0.IN.n18 PFD_T2_0.INV_mag_0.IN.n6 5.77603
R13642 PFD_T2_0.INV_mag_0.IN.n13 PFD_T2_0.INV_mag_0.IN.n10 5.58741
R13643 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.IN.n30 5.21028
R13644 PFD_T2_0.INV_mag_0.IN.n2 PFD_T2_0.INV_mag_0.IN.n22 4.7386
R13645 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.IN.t18 4.69432
R13646 PFD_T2_0.INV_mag_0.IN.n25 PFD_T2_0.INV_mag_0.IN.t30 3.6505
R13647 PFD_T2_0.INV_mag_0.IN.n26 PFD_T2_0.INV_mag_0.IN.t22 3.6505
R13648 PFD_T2_0.INV_mag_0.IN.n20 PFD_T2_0.INV_mag_0.IN.t12 3.6405
R13649 PFD_T2_0.INV_mag_0.IN.n20 PFD_T2_0.INV_mag_0.IN.n19 3.6405
R13650 PFD_T2_0.INV_mag_0.IN.n8 PFD_T2_0.INV_mag_0.IN.t13 3.6405
R13651 PFD_T2_0.INV_mag_0.IN.n8 PFD_T2_0.INV_mag_0.IN.n7 3.6405
R13652 PFD_T2_0.INV_mag_0.IN.n10 PFD_T2_0.INV_mag_0.IN.t11 3.6405
R13653 PFD_T2_0.INV_mag_0.IN.n10 PFD_T2_0.INV_mag_0.IN.n9 3.6405
R13654 PFD_T2_0.INV_mag_0.IN.n15 PFD_T2_0.INV_mag_0.IN.t16 3.6405
R13655 PFD_T2_0.INV_mag_0.IN.n15 PFD_T2_0.INV_mag_0.IN.n14 3.6405
R13656 PFD_T2_0.INV_mag_0.IN.n6 PFD_T2_0.INV_mag_0.IN.t6 3.6405
R13657 PFD_T2_0.INV_mag_0.IN.n6 PFD_T2_0.INV_mag_0.IN.n5 3.6405
R13658 PFD_T2_0.INV_mag_0.IN.n24 PFD_T2_0.INV_mag_0.IN.t5 3.6405
R13659 PFD_T2_0.INV_mag_0.IN.n24 PFD_T2_0.INV_mag_0.IN.n23 3.6405
R13660 PFD_T2_0.INV_mag_0.IN.n12 PFD_T2_0.INV_mag_0.IN.t0 3.2765
R13661 PFD_T2_0.INV_mag_0.IN.n12 PFD_T2_0.INV_mag_0.IN.n11 3.2765
R13662 PFD_T2_0.INV_mag_0.IN.n18 PFD_T2_0.INV_mag_0.IN.n17 3.15378
R13663 PFD_T2_0.INV_mag_0.IN.n2 PFD_T2_0.INV_mag_0.IN.n24 2.94651
R13664 PFD_T2_0.INV_mag_0.IN.n16 PFD_T2_0.INV_mag_0.IN.n15 2.92863
R13665 PFD_T2_0.INV_mag_0.IN.n17 PFD_T2_0.INV_mag_0.IN.n8 2.6005
R13666 PFD_T2_0.INV_mag_0.IN.n0 PFD_T2_0.INV_mag_0.IN.n20 2.6005
R13667 PFD_T2_0.INV_mag_0.IN.n0 PFD_T2_0.INV_mag_0.IN.n18 2.57308
R13668 PFD_T2_0.INV_mag_0.IN.n16 PFD_T2_0.INV_mag_0.IN.n13 2.26925
R13669 PFD_T2_0.INV_mag_0.IN.n17 PFD_T2_0.INV_mag_0.IN.n16 1.00114
R13670 PFD_T2_0.INV_mag_0.IN.n30 PFD_T2_0.INV_mag_0.IN.n0 3.21412
R13671 PFD_T2_0.INV_mag_0.IN.n0 PFD_T2_0.INV_mag_0.IN.n2 2.10654
R13672 a_24437_9224.n1 a_24437_9224.n0 7.21994
R13673 a_24437_9224.n1 a_24437_9224.t0 7.21316
R13674 a_24437_9224.n2 a_24437_9224.t2 3.6405
R13675 a_24437_9224.n3 a_24437_9224.n2 3.6405
R13676 a_24437_9224.n2 a_24437_9224.n1 2.76192
R13677 a_20903_8375.n0 a_20903_8375.t8 29.2961
R13678 a_20903_8375.n1 a_20903_8375.n0 21.9292
R13679 a_20903_8375.n2 a_20903_8375.n1 18.1271
R13680 a_20903_8375.n2 a_20903_8375.t9 11.1695
R13681 a_20903_8375.n0 a_20903_8375.t7 6.1325
R13682 a_20903_8375.n1 a_20903_8375.t6 6.1325
R13683 a_20903_8375.n6 a_20903_8375.n5 4.93252
R13684 a_20903_8375.n6 a_20903_8375.t3 4.70348
R13685 a_20903_8375.n8 a_20903_8375.n2 4.6311
R13686 a_20903_8375.n10 a_20903_8375.n8 2.85093
R13687 a_20903_8375.n4 a_20903_8375.t4 2.16717
R13688 a_20903_8375.n4 a_20903_8375.n3 2.16717
R13689 a_20903_8375.t0 a_20903_8375.n10 2.16717
R13690 a_20903_8375.n10 a_20903_8375.n9 2.16717
R13691 a_20903_8375.n7 a_20903_8375.n6 1.58582
R13692 a_20903_8375.n7 a_20903_8375.n4 1.24371
R13693 a_20903_8375.n8 a_20903_8375.n7 0.971051
R13694 DIV_OUT.n7 DIV_OUT.t3 5.81586
R13695 DIV_OUT.n4 DIV_OUT.n1 5.10148
R13696 DIV_OUT.n11 DIV_OUT.n10 5.10115
R13697 DIV_OUT.n9 DIV_OUT.n8 5.08021
R13698 DIV_OUT.n4 DIV_OUT.n3 4.66166
R13699 DIV_OUT.n7 DIV_OUT.n6 2.85093
R13700 DIV_OUT.n6 DIV_OUT.t4 2.16717
R13701 DIV_OUT.n6 DIV_OUT.n5 2.16717
R13702 DIV_OUT.n3 DIV_OUT.t0 1.9505
R13703 DIV_OUT.n3 DIV_OUT.n2 1.9505
R13704 DIV_OUT.n0 DIV_OUT 1.94122
R13705 DIV_OUT DIV_OUT.n0 1.5484
R13706 DIV_OUT.n0 DIV_OUT 0.838432
R13707 DIV_OUT.n9 DIV_OUT.n7 0.644196
R13708 DIV_OUT.n11 DIV_OUT.n9 0.45084
R13709 DIV_OUT.n12 DIV_OUT.n4 0.309585
R13710 DIV_OUT.n12 DIV_OUT.n11 0.274999
R13711 DIV_OUT DIV_OUT.n12 0.0936034
R13712 PFD_T2_0.FDIV.n4 PFD_T2_0.FDIV.n3 13.9524
R13713 PFD_T2_0.FDIV.n3 PFD_T2_0.FDIV.t17 12.4105
R13714 PFD_T2_0.FDIV.n3 PFD_T2_0.FDIV.t19 11.5345
R13715 PFD_T2_0.FDIV PFD_T2_0.FDIV.n4 8.4325
R13716 PFD_T2_0.FDIV.n4 PFD_T2_0.FDIV.t16 8.1035
R13717 PFD_T2_0.FDIV.n4 PFD_T2_0.FDIV.t18 7.6655
R13718 PFD_T2_0.FDIV.n0 PFD_T2_0.FDIV.t12 6.74332
R13719 PFD_T2_0.FDIV.n1 PFD_T2_0.FDIV.n21 6.74326
R13720 PFD_T2_0.FDIV.n1 PFD_T2_0.FDIV.n22 5.1005
R13721 PFD_T2_0.FDIV.n0 PFD_T2_0.FDIV.t11 5.1005
R13722 PFD_T2_0.FDIV.n19 PFD_T2_0.FDIV.n16 3.57508
R13723 PFD_T2_0.FDIV.n5 PFD_T2_0.FDIV.n8 3.56654
R13724 PFD_T2_0.FDIV.n1 PFD_T2_0.FDIV.t6 3.40075
R13725 PFD_T2_0.FDIV.n0 PFD_T2_0.FDIV.n11 3.40011
R13726 PFD_T2_0.FDIV.n12 PFD_T2_0.FDIV.t3 3.00158
R13727 PFD_T2_0.FDIV.n23 PFD_T2_0.FDIV.n20 3.00032
R13728 PFD_T2_0.FDIV.n14 PFD_T2_0.FDIV 2.51201
R13729 PFD_T2_0.FDIV.n6 PFD_T2_0.FDIV.n10 2.41287
R13730 PFD_T2_0.FDIV.n25 PFD_T2_0.FDIV.n14 2.36206
R13731 PFD_T2_0.FDIV.n14 PFD_T2_0.FDIV.n13 2.30849
R13732 PFD_T2_0.FDIV.n2 PFD_T2_0.FDIV.n6 2.26352
R13733 PFD_T2_0.FDIV.n8 PFD_T2_0.FDIV.t9 2.16717
R13734 PFD_T2_0.FDIV.n8 PFD_T2_0.FDIV.n7 2.16717
R13735 PFD_T2_0.FDIV.n18 PFD_T2_0.FDIV.t1 2.16717
R13736 PFD_T2_0.FDIV.n18 PFD_T2_0.FDIV.n17 2.16717
R13737 PFD_T2_0.FDIV.n16 PFD_T2_0.FDIV.t15 2.16717
R13738 PFD_T2_0.FDIV.n16 PFD_T2_0.FDIV.n15 2.16717
R13739 PFD_T2_0.FDIV.n10 PFD_T2_0.FDIV.t7 2.16717
R13740 PFD_T2_0.FDIV.n10 PFD_T2_0.FDIV.n9 2.16717
R13741 PFD_T2_0.FDIV.n24 PFD_T2_0.FDIV.n23 1.84797
R13742 PFD_T2_0.FDIV.n2 PFD_T2_0.FDIV.n12 1.82978
R13743 PFD_T2_0.FDIV.n19 PFD_T2_0.FDIV.n18 1.25233
R13744 PFD_T2_0.FDIV.n24 PFD_T2_0.FDIV.n19 1.12574
R13745 PFD_T2_0.FDIV PFD_T2_0.FDIV.n25 0.751569
R13746 PFD_T2_0.FDIV.n13 PFD_T2_0.FDIV 0.736653
R13747 PFD_T2_0.FDIV.n23 PFD_T2_0.FDIV.n1 0.558374
R13748 PFD_T2_0.FDIV.n12 PFD_T2_0.FDIV.n0 0.558372
R13749 PFD_T2_0.FDIV.n13 PFD_T2_0.FDIV.n2 0.394824
R13750 PFD_T2_0.FDIV.n25 PFD_T2_0.FDIV.n24 0.33941
R13751 PFD_T2_0.FDIV.n6 PFD_T2_0.FDIV.n5 0.145661
R13752 a_50528_5246.n77 a_50528_5246.t75 40.255
R13753 a_50528_5246.n36 a_50528_5246.t91 37.7641
R13754 a_50528_5246.t98 a_50528_5246.n34 30.4352
R13755 a_50528_5246.t50 a_50528_5246.n52 28.4705
R13756 a_50528_5246.t26 a_50528_5246.n59 28.4705
R13757 a_50528_5246.t58 a_50528_5246.n66 28.4705
R13758 a_50528_5246.t64 a_50528_5246.n73 28.4705
R13759 a_50528_5246.t38 a_50528_5246.n81 28.4705
R13760 a_50528_5246.n85 a_50528_5246.t117 27.3249
R13761 a_50528_5246.n52 a_50528_5246.t82 27.1982
R13762 a_50528_5246.t117 a_50528_5246.n84 25.4384
R13763 a_50528_5246.n84 a_50528_5246.t94 25.4384
R13764 a_50528_5246.n82 a_50528_5246.t60 25.4045
R13765 a_50528_5246.n76 a_50528_5246.t110 25.4045
R13766 a_50528_5246.n76 a_50528_5246.t87 25.4045
R13767 a_50528_5246.n75 a_50528_5246.t37 25.4045
R13768 a_50528_5246.n75 a_50528_5246.t112 25.4045
R13769 a_50528_5246.n67 a_50528_5246.t80 25.4045
R13770 a_50528_5246.n62 a_50528_5246.t102 25.4045
R13771 a_50528_5246.n62 a_50528_5246.t81 25.4045
R13772 a_50528_5246.n61 a_50528_5246.t57 25.4045
R13773 a_50528_5246.n61 a_50528_5246.t35 25.4045
R13774 a_50528_5246.n12 a_50528_5246.t32 25.4045
R13775 a_50528_5246.n12 a_50528_5246.t104 25.4045
R13776 a_50528_5246.n13 a_50528_5246.t77 25.4045
R13777 a_50528_5246.n13 a_50528_5246.t56 25.4045
R13778 a_50528_5246.n14 a_50528_5246.t53 25.4045
R13779 a_50528_5246.n14 a_50528_5246.t34 25.4045
R13780 a_50528_5246.n15 a_50528_5246.t39 25.4045
R13781 a_50528_5246.n15 a_50528_5246.t113 25.4045
R13782 a_50528_5246.n16 a_50528_5246.t111 25.4045
R13783 a_50528_5246.n16 a_50528_5246.t88 25.4045
R13784 a_50528_5246.n17 a_50528_5246.t61 25.4045
R13785 a_50528_5246.n17 a_50528_5246.t40 25.4045
R13786 a_50528_5246.n18 a_50528_5246.t108 25.4045
R13787 a_50528_5246.n18 a_50528_5246.t85 25.4045
R13788 a_50528_5246.n19 a_50528_5246.t83 25.4045
R13789 a_50528_5246.n19 a_50528_5246.t63 25.4045
R13790 a_50528_5246.n20 a_50528_5246.t67 25.4045
R13791 a_50528_5246.n20 a_50528_5246.t44 25.4045
R13792 a_50528_5246.n21 a_50528_5246.t116 25.4045
R13793 a_50528_5246.n21 a_50528_5246.t93 25.4045
R13794 a_50528_5246.n22 a_50528_5246.t66 25.4045
R13795 a_50528_5246.n22 a_50528_5246.t43 25.4045
R13796 a_50528_5246.n23 a_50528_5246.t115 25.4045
R13797 a_50528_5246.n23 a_50528_5246.t92 25.4045
R13798 a_50528_5246.n35 a_50528_5246.t27 25.4045
R13799 a_50528_5246.n35 a_50528_5246.t98 25.4045
R13800 a_50528_5246.n53 a_50528_5246.t71 25.4045
R13801 a_50528_5246.n48 a_50528_5246.t29 25.4045
R13802 a_50528_5246.n46 a_50528_5246.t74 25.4045
R13803 a_50528_5246.n46 a_50528_5246.t54 25.4045
R13804 a_50528_5246.n48 a_50528_5246.t100 25.4045
R13805 a_50528_5246.n50 a_50528_5246.t73 25.4045
R13806 a_50528_5246.n50 a_50528_5246.t51 25.4045
R13807 a_50528_5246.n51 a_50528_5246.t62 25.4045
R13808 a_50528_5246.t82 a_50528_5246.n51 25.4045
R13809 a_50528_5246.n53 a_50528_5246.t50 25.4045
R13810 a_50528_5246.n54 a_50528_5246.t49 25.4045
R13811 a_50528_5246.n54 a_50528_5246.t28 25.4045
R13812 a_50528_5246.n55 a_50528_5246.t96 25.4045
R13813 a_50528_5246.n55 a_50528_5246.t72 25.4045
R13814 a_50528_5246.n60 a_50528_5246.t47 25.4045
R13815 a_50528_5246.n60 a_50528_5246.t26 25.4045
R13816 a_50528_5246.n67 a_50528_5246.t58 25.4045
R13817 a_50528_5246.n68 a_50528_5246.t31 25.4045
R13818 a_50528_5246.n68 a_50528_5246.t103 25.4045
R13819 a_50528_5246.n69 a_50528_5246.t76 25.4045
R13820 a_50528_5246.n69 a_50528_5246.t55 25.4045
R13821 a_50528_5246.n74 a_50528_5246.t86 25.4045
R13822 a_50528_5246.n74 a_50528_5246.t64 25.4045
R13823 a_50528_5246.n82 a_50528_5246.t38 25.4045
R13824 a_50528_5246.n83 a_50528_5246.t107 25.4045
R13825 a_50528_5246.n83 a_50528_5246.t84 25.4045
R13826 a_50528_5246.n58 a_50528_5246.t59 23.6525
R13827 a_50528_5246.n65 a_50528_5246.t41 23.6525
R13828 a_50528_5246.n72 a_50528_5246.t46 23.6525
R13829 a_50528_5246.n80 a_50528_5246.t45 23.6525
R13830 a_50528_5246.n85 a_50528_5246.t109 23.5689
R13831 a_50528_5246.n86 a_50528_5246.t99 23.5065
R13832 a_50528_5246.n87 a_50528_5246.t52 23.5065
R13833 a_50528_5246.n88 a_50528_5246.t101 23.5065
R13834 a_50528_5246.n89 a_50528_5246.t30 23.5065
R13835 a_50528_5246.n90 a_50528_5246.t79 23.5065
R13836 a_50528_5246.n91 a_50528_5246.t69 23.5065
R13837 a_50528_5246.n92 a_50528_5246.t24 23.5065
R13838 a_50528_5246.n37 a_50528_5246.t89 22.4115
R13839 a_50528_5246.n36 a_50528_5246.t42 22.4115
R13840 a_50528_5246.n57 a_50528_5246.t106 20.4405
R13841 a_50528_5246.n56 a_50528_5246.t36 20.4405
R13842 a_50528_5246.n38 a_50528_5246.t97 20.4405
R13843 a_50528_5246.n39 a_50528_5246.t48 20.4405
R13844 a_50528_5246.n40 a_50528_5246.t25 20.4405
R13845 a_50528_5246.n41 a_50528_5246.t70 20.4405
R13846 a_50528_5246.n42 a_50528_5246.t118 20.4405
R13847 a_50528_5246.n43 a_50528_5246.t33 20.4405
R13848 a_50528_5246.n44 a_50528_5246.t78 20.4405
R13849 a_50528_5246.t54 a_50528_5246.n45 20.4405
R13850 a_50528_5246.t100 a_50528_5246.n47 20.4405
R13851 a_50528_5246.t51 a_50528_5246.n49 20.4405
R13852 a_50528_5246.n63 a_50528_5246.t105 20.4405
R13853 a_50528_5246.n64 a_50528_5246.t90 20.4405
R13854 a_50528_5246.n71 a_50528_5246.t65 20.4405
R13855 a_50528_5246.n70 a_50528_5246.t114 20.4405
R13856 a_50528_5246.n78 a_50528_5246.t119 20.4405
R13857 a_50528_5246.n79 a_50528_5246.t68 20.4405
R13858 a_50528_5246.n77 a_50528_5246.t95 20.4405
R13859 a_50528_5246.n58 a_50528_5246.n57 19.2623
R13860 a_50528_5246.n65 a_50528_5246.n64 19.2623
R13861 a_50528_5246.n72 a_50528_5246.n71 19.2623
R13862 a_50528_5246.n80 a_50528_5246.n79 19.2623
R13863 a_50528_5246.n57 a_50528_5246.n56 17.2497
R13864 a_50528_5246.n64 a_50528_5246.n63 17.2497
R13865 a_50528_5246.n71 a_50528_5246.n70 17.2497
R13866 a_50528_5246.n79 a_50528_5246.n78 17.2497
R13867 a_50528_5246.n82 a_50528_5246.n76 15.8172
R13868 a_50528_5246.n76 a_50528_5246.n75 15.8172
R13869 a_50528_5246.n67 a_50528_5246.n62 15.8172
R13870 a_50528_5246.n62 a_50528_5246.n61 15.8172
R13871 a_50528_5246.n14 a_50528_5246.n13 15.8172
R13872 a_50528_5246.n15 a_50528_5246.n14 15.8172
R13873 a_50528_5246.n16 a_50528_5246.n15 15.8172
R13874 a_50528_5246.n17 a_50528_5246.n16 15.8172
R13875 a_50528_5246.n18 a_50528_5246.n17 15.8172
R13876 a_50528_5246.n19 a_50528_5246.n18 15.8172
R13877 a_50528_5246.n20 a_50528_5246.n19 15.8172
R13878 a_50528_5246.n21 a_50528_5246.n20 15.8172
R13879 a_50528_5246.n22 a_50528_5246.n21 15.8172
R13880 a_50528_5246.n23 a_50528_5246.n22 15.8172
R13881 a_50528_5246.n35 a_50528_5246.n23 15.8172
R13882 a_50528_5246.n53 a_50528_5246.n35 15.8172
R13883 a_50528_5246.n54 a_50528_5246.n53 15.8172
R13884 a_50528_5246.n55 a_50528_5246.n54 15.8172
R13885 a_50528_5246.n60 a_50528_5246.n55 15.8172
R13886 a_50528_5246.n61 a_50528_5246.n60 15.8172
R13887 a_50528_5246.n68 a_50528_5246.n67 15.8172
R13888 a_50528_5246.n69 a_50528_5246.n68 15.8172
R13889 a_50528_5246.n74 a_50528_5246.n69 15.8172
R13890 a_50528_5246.n75 a_50528_5246.n74 15.8172
R13891 a_50528_5246.n83 a_50528_5246.n82 15.8172
R13892 a_50528_5246.n84 a_50528_5246.n83 15.8172
R13893 a_50528_5246.n81 a_50528_5246.n77 15.7165
R13894 a_50528_5246.n13 a_50528_5246.n12 15.4944
R13895 a_50528_5246.n37 a_50528_5246.n36 15.3531
R13896 a_50528_5246.n38 a_50528_5246.n37 15.2373
R13897 a_50528_5246.n39 a_50528_5246.n38 14.4179
R13898 a_50528_5246.n40 a_50528_5246.n39 14.4179
R13899 a_50528_5246.n41 a_50528_5246.n40 14.4179
R13900 a_50528_5246.n42 a_50528_5246.n41 14.4179
R13901 a_50528_5246.n43 a_50528_5246.n42 14.4179
R13902 a_50528_5246.n44 a_50528_5246.n43 14.4179
R13903 a_50528_5246.n45 a_50528_5246.n44 14.3002
R13904 a_50528_5246.n48 a_50528_5246.n46 13.3198
R13905 a_50528_5246.n50 a_50528_5246.n48 13.3198
R13906 a_50528_5246.n51 a_50528_5246.n50 13.3198
R13907 a_50528_5246.n87 a_50528_5246.n86 12.7287
R13908 a_50528_5246.n88 a_50528_5246.n87 12.7287
R13909 a_50528_5246.n89 a_50528_5246.n88 12.7287
R13910 a_50528_5246.n90 a_50528_5246.n89 12.7287
R13911 a_50528_5246.n91 a_50528_5246.n90 12.7287
R13912 a_50528_5246.n92 a_50528_5246.n91 12.7287
R13913 a_50528_5246.n86 a_50528_5246.n85 12.6663
R13914 a_50528_5246.n93 a_50528_5246.n92 4.60781
R13915 a_50528_5246.n101 a_50528_5246.n100 3.69699
R13916 a_50528_5246.n59 a_50528_5246.n58 3.54621
R13917 a_50528_5246.n66 a_50528_5246.n65 3.54621
R13918 a_50528_5246.n73 a_50528_5246.n72 3.54621
R13919 a_50528_5246.n81 a_50528_5246.n80 3.54621
R13920 a_50528_5246.n94 a_50528_5246.n9 3.23924
R13921 a_50528_5246.n95 a_50528_5246.n7 3.23924
R13922 a_50528_5246.n96 a_50528_5246.n5 3.23924
R13923 a_50528_5246.n93 a_50528_5246.n11 3.2392
R13924 a_50528_5246.n102 a_50528_5246.n101 3.2392
R13925 a_50528_5246.n97 a_50528_5246.n3 3.23916
R13926 a_50528_5246.n98 a_50528_5246.n1 3.23916
R13927 a_50528_5246.n28 a_50528_5246.n25 2.91928
R13928 a_50528_5246.n34 a_50528_5246.n33 2.58908
R13929 a_50528_5246.n31 a_50528_5246.n30 2.58711
R13930 a_50528_5246.n28 a_50528_5246.n27 2.58292
R13931 a_50528_5246.n11 a_50528_5246.t15 0.6505
R13932 a_50528_5246.n11 a_50528_5246.n10 0.6505
R13933 a_50528_5246.n9 a_50528_5246.t18 0.6505
R13934 a_50528_5246.n9 a_50528_5246.n8 0.6505
R13935 a_50528_5246.n7 a_50528_5246.t13 0.6505
R13936 a_50528_5246.n7 a_50528_5246.n6 0.6505
R13937 a_50528_5246.n5 a_50528_5246.t20 0.6505
R13938 a_50528_5246.n5 a_50528_5246.n4 0.6505
R13939 a_50528_5246.n3 a_50528_5246.t3 0.6505
R13940 a_50528_5246.n3 a_50528_5246.n2 0.6505
R13941 a_50528_5246.n1 a_50528_5246.t12 0.6505
R13942 a_50528_5246.n1 a_50528_5246.n0 0.6505
R13943 a_50528_5246.n100 a_50528_5246.t10 0.6505
R13944 a_50528_5246.n100 a_50528_5246.n99 0.6505
R13945 a_50528_5246.n102 a_50528_5246.t14 0.6505
R13946 a_50528_5246.n103 a_50528_5246.n102 0.6505
R13947 a_50528_5246.n33 a_50528_5246.t21 0.5855
R13948 a_50528_5246.n33 a_50528_5246.n32 0.5855
R13949 a_50528_5246.n25 a_50528_5246.t7 0.5855
R13950 a_50528_5246.n25 a_50528_5246.n24 0.5855
R13951 a_50528_5246.n27 a_50528_5246.t0 0.5855
R13952 a_50528_5246.n27 a_50528_5246.n26 0.5855
R13953 a_50528_5246.n30 a_50528_5246.t16 0.5855
R13954 a_50528_5246.n30 a_50528_5246.n29 0.5855
R13955 a_50528_5246.n98 a_50528_5246.n97 0.466449
R13956 a_50528_5246.n94 a_50528_5246.n93 0.46531
R13957 a_50528_5246.n95 a_50528_5246.n94 0.46531
R13958 a_50528_5246.n96 a_50528_5246.n95 0.46531
R13959 a_50528_5246.n101 a_50528_5246.n98 0.46531
R13960 a_50528_5246.n97 a_50528_5246.n96 0.464171
R13961 a_50528_5246.n31 a_50528_5246.n28 0.341015
R13962 a_50528_5246.n34 a_50528_5246.n31 0.337297
R13963 OUTB.n8 OUTB.n7 3.74358
R13964 OUTB.n10 OUTB.n1 3.24303
R13965 OUTB.n9 OUTB.n3 3.24286
R13966 OUTB.n8 OUTB.n5 3.24211
R13967 OUTB.n84 OUTB.n21 3.23441
R13968 OUTB.n81 OUTB.n27 3.23441
R13969 OUTB.n76 OUTB.n39 3.23441
R13970 OUTB.n69 OUTB.n55 3.23441
R13971 OUTB.n68 OUTB.n59 3.23441
R13972 OUTB.n81 OUTB.n29 3.23391
R13973 OUTB.n83 OUTB.n23 3.23391
R13974 OUTB.n76 OUTB.n41 3.23387
R13975 OUTB.n73 OUTB.n47 3.23387
R13976 OUTB.n75 OUTB.n43 3.23387
R13977 OUTB.n78 OUTB.n35 3.23387
R13978 OUTB.n80 OUTB.n31 3.23387
R13979 OUTB.n69 OUTB.n57 3.23383
R13980 OUTB.n67 OUTB.n61 3.23383
R13981 OUTB.n71 OUTB.n51 3.23383
R13982 OUTB.n82 OUTB.n25 3.23358
R13983 OUTB.n66 OUTB.n65 3.2335
R13984 OUTB.n85 OUTB.n19 3.23343
R13985 OUTB.n87 OUTB.n15 3.23343
R13986 OUTB.n86 OUTB.n17 3.23337
R13987 OUTB.n79 OUTB.n33 3.23316
R13988 OUTB.n77 OUTB.n37 3.23312
R13989 OUTB.n74 OUTB.n45 3.23312
R13990 OUTB.n72 OUTB.n49 3.23312
R13991 OUTB.n70 OUTB.n53 3.23312
R13992 OUTB.n66 OUTB.n63 3.2315
R13993 OUTB.n100 OUTB.n97 2.98385
R13994 OUTB.n113 OUTB.n95 2.87549
R13995 OUTB.n116 OUTB.n115 2.70972
R13996 OUTB.n119 OUTB.n118 2.62238
R13997 OUTB.n122 OUTB.n121 2.62091
R13998 OUTB.n125 OUTB.n124 2.61945
R13999 OUTB.n131 OUTB.n130 2.61636
R14000 OUTB.n137 OUTB.n136 2.61619
R14001 OUTB.n128 OUTB.n127 2.61619
R14002 OUTB.n134 OUTB.n133 2.61554
R14003 OUTB.n13 OUTB.n12 2.6005
R14004 OUTB.n91 OUTB.n90 2.6005
R14005 OUTB.n100 OUTB.n99 2.58236
R14006 OUTB.n106 OUTB.n105 2.58184
R14007 OUTB.n109 OUTB.n108 2.5817
R14008 OUTB.n103 OUTB.n102 2.58166
R14009 OUTB.n112 OUTB.n111 2.58122
R14010 OUTB.n138 OUTB.n137 1.60202
R14011 OUTB.n138 OUTB.n93 1.34978
R14012 OUTB.n139 OUTB.n138 0.888141
R14013 OUTB.n13 OUTB.n10 0.79069
R14014 OUTB.n84 OUTB.n83 0.781777
R14015 OUTB.n81 OUTB.n80 0.781777
R14016 OUTB.n76 OUTB.n75 0.781777
R14017 OUTB.n69 OUTB.n68 0.781777
R14018 OUTB.n67 OUTB.n66 0.781777
R14019 OUTB.n82 OUTB.n81 0.779862
R14020 OUTB.n79 OUTB.n78 0.779862
R14021 OUTB.n77 OUTB.n76 0.779862
R14022 OUTB.n74 OUTB.n73 0.779862
R14023 OUTB.n72 OUTB.n71 0.779862
R14024 OUTB.n70 OUTB.n69 0.779862
R14025 OUTB.n88 OUTB.n87 0.777947
R14026 OUTB.n86 OUTB.n85 0.777947
R14027 OUTB.n139 OUTB.n91 0.655477
R14028 OUTB.n90 OUTB.t49 0.6505
R14029 OUTB.n90 OUTB.n89 0.6505
R14030 OUTB.n12 OUTB.t32 0.6505
R14031 OUTB.n12 OUTB.n11 0.6505
R14032 OUTB.n1 OUTB.t39 0.6505
R14033 OUTB.n1 OUTB.n0 0.6505
R14034 OUTB.n3 OUTB.t77 0.6505
R14035 OUTB.n3 OUTB.n2 0.6505
R14036 OUTB.n5 OUTB.t91 0.6505
R14037 OUTB.n5 OUTB.n4 0.6505
R14038 OUTB.n7 OUTB.t65 0.6505
R14039 OUTB.n7 OUTB.n6 0.6505
R14040 OUTB.n17 OUTB.t71 0.6505
R14041 OUTB.n17 OUTB.n16 0.6505
R14042 OUTB.n21 OUTB.t86 0.6505
R14043 OUTB.n21 OUTB.n20 0.6505
R14044 OUTB.n25 OUTB.t62 0.6505
R14045 OUTB.n25 OUTB.n24 0.6505
R14046 OUTB.n29 OUTB.t72 0.6505
R14047 OUTB.n29 OUTB.n28 0.6505
R14048 OUTB.n27 OUTB.t59 0.6505
R14049 OUTB.n27 OUTB.n26 0.6505
R14050 OUTB.n33 OUTB.t73 0.6505
R14051 OUTB.n33 OUTB.n32 0.6505
R14052 OUTB.n37 OUTB.t48 0.6505
R14053 OUTB.n37 OUTB.n36 0.6505
R14054 OUTB.n41 OUTB.t78 0.6505
R14055 OUTB.n41 OUTB.n40 0.6505
R14056 OUTB.n39 OUTB.t64 0.6505
R14057 OUTB.n39 OUTB.n38 0.6505
R14058 OUTB.n45 OUTB.t34 0.6505
R14059 OUTB.n45 OUTB.n44 0.6505
R14060 OUTB.n49 OUTB.t33 0.6505
R14061 OUTB.n49 OUTB.n48 0.6505
R14062 OUTB.n53 OUTB.t57 0.6505
R14063 OUTB.n53 OUTB.n52 0.6505
R14064 OUTB.n57 OUTB.t83 0.6505
R14065 OUTB.n57 OUTB.n56 0.6505
R14066 OUTB.n55 OUTB.t70 0.6505
R14067 OUTB.n55 OUTB.n54 0.6505
R14068 OUTB.n59 OUTB.t84 0.6505
R14069 OUTB.n59 OUTB.n58 0.6505
R14070 OUTB.n65 OUTB.t74 0.6505
R14071 OUTB.n65 OUTB.n64 0.6505
R14072 OUTB.n63 OUTB.t61 0.6505
R14073 OUTB.n63 OUTB.n62 0.6505
R14074 OUTB.n61 OUTB.t35 0.6505
R14075 OUTB.n61 OUTB.n60 0.6505
R14076 OUTB.n51 OUTB.t69 0.6505
R14077 OUTB.n51 OUTB.n50 0.6505
R14078 OUTB.n47 OUTB.t50 0.6505
R14079 OUTB.n47 OUTB.n46 0.6505
R14080 OUTB.n43 OUTB.t51 0.6505
R14081 OUTB.n43 OUTB.n42 0.6505
R14082 OUTB.n35 OUTB.t63 0.6505
R14083 OUTB.n35 OUTB.n34 0.6505
R14084 OUTB.n31 OUTB.t87 0.6505
R14085 OUTB.n31 OUTB.n30 0.6505
R14086 OUTB.n23 OUTB.t75 0.6505
R14087 OUTB.n23 OUTB.n22 0.6505
R14088 OUTB.n19 OUTB.t36 0.6505
R14089 OUTB.n19 OUTB.n18 0.6505
R14090 OUTB.n15 OUTB.t85 0.6505
R14091 OUTB.n15 OUTB.n14 0.6505
R14092 OUTB.n91 OUTB.n88 0.633955
R14093 OUTB.n88 OUTB.n13 0.631666
R14094 OUTB.n127 OUTB.t27 0.5855
R14095 OUTB.n127 OUTB.n126 0.5855
R14096 OUTB.n133 OUTB.t0 0.5855
R14097 OUTB.n133 OUTB.n132 0.5855
R14098 OUTB.n136 OUTB.t25 0.5855
R14099 OUTB.n136 OUTB.n135 0.5855
R14100 OUTB.n115 OUTB.t30 0.5855
R14101 OUTB.n115 OUTB.n114 0.5855
R14102 OUTB.n118 OUTB.t11 0.5855
R14103 OUTB.n118 OUTB.n117 0.5855
R14104 OUTB.n121 OUTB.t3 0.5855
R14105 OUTB.n121 OUTB.n120 0.5855
R14106 OUTB.n124 OUTB.t4 0.5855
R14107 OUTB.n124 OUTB.n123 0.5855
R14108 OUTB.n130 OUTB.t18 0.5855
R14109 OUTB.n130 OUTB.n129 0.5855
R14110 OUTB.n97 OUTB.t26 0.5855
R14111 OUTB.n97 OUTB.n96 0.5855
R14112 OUTB.n99 OUTB.t6 0.5855
R14113 OUTB.n99 OUTB.n98 0.5855
R14114 OUTB.n102 OUTB.t31 0.5855
R14115 OUTB.n102 OUTB.n101 0.5855
R14116 OUTB.n105 OUTB.t1 0.5855
R14117 OUTB.n105 OUTB.n104 0.5855
R14118 OUTB.n108 OUTB.t12 0.5855
R14119 OUTB.n108 OUTB.n107 0.5855
R14120 OUTB.n111 OUTB.t5 0.5855
R14121 OUTB.n111 OUTB.n110 0.5855
R14122 OUTB.n95 OUTB.t19 0.5855
R14123 OUTB.n95 OUTB.n94 0.5855
R14124 OUTB.n93 OUTB.t13 0.5855
R14125 OUTB.n93 OUTB.n92 0.5855
R14126 OUTB.n116 OUTB.n113 0.510866
R14127 OUTB.n10 OUTB.n9 0.504747
R14128 OUTB.n9 OUTB.n8 0.504747
R14129 OUTB.n106 OUTB.n103 0.403414
R14130 OUTB.n109 OUTB.n106 0.402304
R14131 OUTB.n112 OUTB.n109 0.400958
R14132 OUTB.n103 OUTB.n100 0.400949
R14133 OUTB OUTB.n139 0.354162
R14134 OUTB.n128 OUTB.n125 0.334681
R14135 OUTB.n131 OUTB.n128 0.334473
R14136 OUTB.n122 OUTB.n119 0.334465
R14137 OUTB.n134 OUTB.n131 0.334064
R14138 OUTB.n137 OUTB.n134 0.333663
R14139 OUTB.n125 OUTB.n122 0.333454
R14140 OUTB.n119 OUTB.n116 0.244714
R14141 OUTB.n113 OUTB.n112 0.107492
R14142 OUTB.n87 OUTB.n86 0.00432979
R14143 OUTB.n85 OUTB.n84 0.00241489
R14144 OUTB.n83 OUTB.n82 0.00241489
R14145 OUTB.n80 OUTB.n79 0.00241489
R14146 OUTB.n78 OUTB.n77 0.00241489
R14147 OUTB.n75 OUTB.n74 0.00241489
R14148 OUTB.n73 OUTB.n72 0.00241489
R14149 OUTB.n71 OUTB.n70 0.00241489
R14150 OUTB.n68 OUTB.n67 0.00241489
R14151 ITAIL.n7 ITAIL.t2 10.9054
R14152 ITAIL.n0 ITAIL.t20 10.8613
R14153 ITAIL.n17 ITAIL.t26 10.773
R14154 ITAIL.n13 ITAIL.t24 10.6003
R14155 ITAIL.n0 ITAIL.t10 10.5984
R14156 ITAIL.n17 ITAIL.t0 10.5336
R14157 ITAIL.n7 ITAIL.t16 10.5336
R14158 ITAIL.n1 ITAIL.t18 10.5334
R14159 ITAIL.n35 ITAIL.t19 10.533
R14160 ITAIL.n34 ITAIL.t14 10.5098
R14161 ITAIL.n18 ITAIL.t21 10.4686
R14162 ITAIL.n16 ITAIL.t4 10.0514
R14163 ITAIL.n10 ITAIL.t8 9.72546
R14164 ITAIL.n4 ITAIL.t12 9.65907
R14165 ITAIL.n36 ITAIL.t6 9.29485
R14166 ITAIL.n37 ITAIL.t25 8.47237
R14167 ITAIL.n29 ITAIL.t13 8.17686
R14168 ITAIL.n24 ITAIL.t5 8.07837
R14169 ITAIL.n25 ITAIL.n23 7.98962
R14170 ITAIL.n30 ITAIL.n28 7.84993
R14171 ITAIL.n29 ITAIL.t11 7.79699
R14172 ITAIL.n32 ITAIL.n26 7.73548
R14173 ITAIL.n24 ITAIL.t1 7.72811
R14174 ITAIL.n31 ITAIL.n27 7.58076
R14175 ITAIL.n39 ITAIL 6.54657
R14176 ITAIL ITAIL.n39 2.524
R14177 ITAIL.n32 ITAIL.n31 1.75757
R14178 ITAIL.n20 ITAIL.n16 1.50725
R14179 ITAIL.n11 ITAIL.n10 1.50717
R14180 ITAIL.n6 ITAIL.n5 1.49748
R14181 ITAIL.n39 ITAIL.n38 0.668
R14182 ITAIL.n31 ITAIL.n30 0.661924
R14183 ITAIL.n14 ITAIL.n6 0.490305
R14184 ITAIL.n21 ITAIL.n14 0.446994
R14185 ITAIL.n37 ITAIL.n36 0.413008
R14186 ITAIL.n1 ITAIL.n0 0.390708
R14187 ITAIL.n36 ITAIL.n35 0.375243
R14188 ITAIL.n18 ITAIL.n17 0.365503
R14189 ITAIL.n19 ITAIL.n18 0.357915
R14190 ITAIL.n2 ITAIL.n1 0.357771
R14191 ITAIL.n13 ITAIL.n12 0.356995
R14192 ITAIL.n8 ITAIL.n7 0.341087
R14193 ITAIL.n33 ITAIL.n32 0.31096
R14194 ITAIL.n25 ITAIL.n24 0.301864
R14195 ITAIL.n30 ITAIL.n29 0.285711
R14196 ITAIL.n38 ITAIL.n22 0.278
R14197 ITAIL.n38 ITAIL.n37 0.244031
R14198 ITAIL.n33 ITAIL.n25 0.2255
R14199 ITAIL.n35 ITAIL.n34 0.201238
R14200 ITAIL.n34 ITAIL.n33 0.1493
R14201 ITAIL.n11 ITAIL.n8 0.028981
R14202 ITAIL.n14 ITAIL.n13 0.0236995
R14203 ITAIL.n21 ITAIL.n20 0.017375
R14204 ITAIL.n12 ITAIL.n11 0.0163348
R14205 ITAIL.n20 ITAIL.n19 0.0150187
R14206 ITAIL.n6 ITAIL.n3 0.013491
R14207 ITAIL.n3 ITAIL.n2 0.0117754
R14208 ITAIL.n22 ITAIL.n21 0.003875
R14209 ITAIL.n16 ITAIL.n15 0.00243623
R14210 ITAIL.n10 ITAIL.n9 0.00242648
R14211 ITAIL.n5 ITAIL.n4 0.00155882
R14212 a_32731_10265.n9 a_32731_10265.n8 10.0413
R14213 a_32731_10265.n6 a_32731_10265.t4 8.81226
R14214 a_32731_10265.n9 a_32731_10265.n7 8.80202
R14215 a_32731_10265.n5 a_32731_10265.t6 8.78441
R14216 a_32731_10265.n0 a_32731_10265.t5 8.6005
R14217 a_32731_10265.n1 a_32731_10265.n10 8.15323
R14218 a_32731_10265.n1 a_32731_10265.n11 8.13693
R14219 a_32731_10265.t7 a_32731_10265.n1 8.00806
R14220 a_32731_10265.n2 a_32731_10265.t2 5.72901
R14221 a_32731_10265.n2 a_32731_10265.t11 5.2005
R14222 a_32731_10265.n3 a_32731_10265.t0 5.2005
R14223 a_32731_10265.n4 a_32731_10265.t1 5.2005
R14224 a_32731_10265.n1 a_32731_10265.n0 3.13877
R14225 a_32731_10265.n0 a_32731_10265.n6 2.42442
R14226 a_32731_10265.n0 a_32731_10265.n9 2.34763
R14227 a_32731_10265.n5 a_32731_10265.n4 1.88322
R14228 a_32731_10265.n6 a_32731_10265.n5 1.10344
R14229 a_32731_10265.n3 a_32731_10265.n2 0.529011
R14230 a_32731_10265.n4 a_32731_10265.n3 0.529011
R14231 CP_1_0.VCTRL.n38 CP_1_0.VCTRL.n37 9.07899
R14232 CP_1_0.VCTRL.t15 CP_1_0.VCTRL.n3 8.83029
R14233 CP_1_0.VCTRL.n40 CP_1_0.VCTRL.n39 8.5505
R14234 CP_1_0.VCTRL.n38 CP_1_0.VCTRL.t30 8.5505
R14235 CP_1_0.VCTRL.n41 CP_1_0.VCTRL.t29 8.03277
R14236 CP_1_0.VCTRL.n1 CP_1_0.VCTRL.t26 6.74332
R14237 CP_1_0.VCTRL.n2 CP_1_0.VCTRL.n10 6.74326
R14238 CP_1_0.VCTRL.n30 CP_1_0.VCTRL.t4 5.81586
R14239 CP_1_0.VCTRL.n36 CP_1_0.VCTRL.n35 5.73034
R14240 CP_1_0.VCTRL.n27 CP_1_0.VCTRL.n24 5.10148
R14241 CP_1_0.VCTRL.n34 CP_1_0.VCTRL.n33 5.10115
R14242 CP_1_0.VCTRL.n1 CP_1_0.VCTRL.t23 5.1005
R14243 CP_1_0.VCTRL.n2 CP_1_0.VCTRL.n11 5.1005
R14244 CP_1_0.VCTRL.n32 CP_1_0.VCTRL.n31 5.08021
R14245 CP_1_0.VCTRL.n27 CP_1_0.VCTRL.n26 4.66166
R14246 CP_1_0.VCTRL.n21 CP_1_0.VCTRL.n20 3.5743
R14247 CP_1_0.VCTRL.n8 CP_1_0.VCTRL.n7 3.5743
R14248 CP_1_0.VCTRL.n2 CP_1_0.VCTRL.t22 3.40065
R14249 CP_1_0.VCTRL.n1 CP_1_0.VCTRL.n15 3.40001
R14250 CP_1_0.VCTRL.n16 CP_1_0.VCTRL.t0 3.00159
R14251 CP_1_0.VCTRL.n12 CP_1_0.VCTRL.n9 3.00034
R14252 CP_1_0.VCTRL.n30 CP_1_0.VCTRL.n29 2.85093
R14253 CP_1_0.VCTRL CP_1_0.VCTRL.n42 2.35764
R14254 CP_1_0.VCTRL.n0 CP_1_0.VCTRL 2.34756
R14255 CP_1_0.VCTRL.n0 CP_1_0.VCTRL.n23 2.25694
R14256 CP_1_0.VCTRL.n0 CP_1_0.VCTRL.n14 2.22474
R14257 CP_1_0.VCTRL.n18 CP_1_0.VCTRL.t8 2.16717
R14258 CP_1_0.VCTRL.n18 CP_1_0.VCTRL.n17 2.16717
R14259 CP_1_0.VCTRL.n20 CP_1_0.VCTRL.t9 2.16717
R14260 CP_1_0.VCTRL.n20 CP_1_0.VCTRL.n19 2.16717
R14261 CP_1_0.VCTRL.n5 CP_1_0.VCTRL.t17 2.16717
R14262 CP_1_0.VCTRL.n5 CP_1_0.VCTRL.n4 2.16717
R14263 CP_1_0.VCTRL.n7 CP_1_0.VCTRL.t10 2.16717
R14264 CP_1_0.VCTRL.n7 CP_1_0.VCTRL.n6 2.16717
R14265 CP_1_0.VCTRL.n29 CP_1_0.VCTRL.t5 2.16717
R14266 CP_1_0.VCTRL.n29 CP_1_0.VCTRL.n28 2.16717
R14267 CP_1_0.VCTRL.n42 CP_1_0.VCTRL.n41 2.01704
R14268 CP_1_0.VCTRL.n26 CP_1_0.VCTRL.t32 1.9505
R14269 CP_1_0.VCTRL.n26 CP_1_0.VCTRL.n25 1.9505
R14270 CP_1_0.VCTRL.n22 CP_1_0.VCTRL.n16 1.84725
R14271 CP_1_0.VCTRL.n13 CP_1_0.VCTRL.n12 1.847
R14272 CP_1_0.VCTRL CP_1_0.VCTRL.t11 1.72887
R14273 CP_1_0.VCTRL.n35 CP_1_0.VCTRL 1.70644
R14274 CP_1_0.VCTRL.n42 CP_1_0.VCTRL.n36 1.39379
R14275 CP_1_0.VCTRL.n21 CP_1_0.VCTRL.n18 1.25225
R14276 CP_1_0.VCTRL.n8 CP_1_0.VCTRL.n5 1.25225
R14277 CP_1_0.VCTRL.n13 CP_1_0.VCTRL.n8 1.12594
R14278 CP_1_0.VCTRL.n22 CP_1_0.VCTRL.n21 1.12575
R14279 CP_1_0.VCTRL.n40 CP_1_0.VCTRL.n38 1.1179
R14280 CP_1_0.VCTRL.n35 CP_1_0.VCTRL 1.06348
R14281 CP_1_0.VCTRL.n14 CP_1_0.VCTRL 0.751569
R14282 CP_1_0.VCTRL.n23 CP_1_0.VCTRL 0.736831
R14283 CP_1_0.VCTRL.t11 CP_1_0.VCTRL.t15 0.683746
R14284 CP_1_0.VCTRL.n32 CP_1_0.VCTRL.n30 0.644196
R14285 CP_1_0.VCTRL.n12 CP_1_0.VCTRL.n2 0.559412
R14286 CP_1_0.VCTRL.n16 CP_1_0.VCTRL.n1 0.55941
R14287 CP_1_0.VCTRL.n41 CP_1_0.VCTRL.n40 0.454295
R14288 CP_1_0.VCTRL.n34 CP_1_0.VCTRL.n32 0.45084
R14289 CP_1_0.VCTRL.n23 CP_1_0.VCTRL.n22 0.378694
R14290 CP_1_0.VCTRL CP_1_0.VCTRL.n34 0.368102
R14291 CP_1_0.VCTRL.n36 CP_1_0.VCTRL.n0 0.364361
R14292 CP_1_0.VCTRL.n14 CP_1_0.VCTRL.n13 0.33941
R14293 CP_1_0.VCTRL CP_1_0.VCTRL.n27 0.309585
R14294 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t41 23.6945
R14295 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t51 23.6945
R14296 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n21 18.8035
R14297 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n16 15.8172
R14298 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n24 15.8172
R14299 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n16 15.8172
R14300 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t56 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n19 14.8925
R14301 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t42 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n16 14.8925
R14302 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t49 14.8925
R14303 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n17 12.2457
R14304 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n18 12.2457
R14305 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n18 12.2457
R14306 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t37 11.6285
R14307 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t34 9.07373
R14308 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t55 8.94903
R14309 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t50 8.91906
R14310 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t32 8.91906
R14311 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t54 8.91906
R14312 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t41 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n20 8.9065
R14313 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t57 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n18 8.9065
R14314 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t36 8.9065
R14315 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t51 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n17 8.9065
R14316 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t43 8.88175
R14317 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t48 8.78051
R14318 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t44 8.78051
R14319 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t38 8.76753
R14320 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t58 8.76753
R14321 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t4 8.71893
R14322 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t52 8.71324
R14323 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t46 8.71324
R14324 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t53 8.6145
R14325 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t40 8.6145
R14326 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t45 8.6145
R14327 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t31 8.59715
R14328 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t35 8.50259
R14329 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t47 8.38837
R14330 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t56 8.3225
R14331 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t42 8.3225
R14332 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n23 8.3225
R14333 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t37 8.3225
R14334 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t33 8.30411
R14335 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t39 7.40199
R14336 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t27 6.43598
R14337 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n14 6.42121
R14338 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t28 6.39767
R14339 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t10 6.02888
R14340 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n32 5.82997
R14341 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n45 8.13848
R14342 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n35 5.23266
R14343 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t14 4.93756
R14344 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t22 4.89657
R14345 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n51 4.89332
R14346 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t6 4.76585
R14347 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n29 4.70534
R14348 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n28 4.70317
R14349 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n26 4.60939
R14350 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n6 4.53389
R14351 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n54 4.22351
R14352 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n43 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n42 4.04842
R14353 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t23 4.00791
R14354 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n57 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n56 3.96274
R14355 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n27 3.95313
R14356 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t5 3.94347
R14357 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t26 3.80888
R14358 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n31 3.77407
R14359 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n59 3.75752
R14360 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 3.73676
R14361 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n58 3.65963
R14362 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t57 3.6505
R14363 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t36 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n22 3.6505
R14364 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t19 3.6405
R14365 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n48 3.6405
R14366 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t13 3.6405
R14367 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n46 3.6405
R14368 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t12 3.6405
R14369 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n39 3.6405
R14370 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n34 3.47613
R14371 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n30 3.47611
R14372 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n33 3.35867
R14373 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n36 3.3208
R14374 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t21 3.31772
R14375 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n13 3.31211
R14376 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n25 3.1807
R14377 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 3.15957
R14378 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n12 3.14573
R14379 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n50 2.97396
R14380 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t2 2.86261
R14381 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.t0 2.8626
R14382 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 2.7938
R14383 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n55 2.75901
R14384 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n15 2.62313
R14385 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 2.36584
R14386 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n37 2.35267
R14387 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n44 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n43 2.24883
R14388 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n52 2.24559
R14389 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n2 2.03424
R14390 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n9 1.9805
R14391 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n10 1.86182
R14392 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n53 1.85837
R14393 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n7 1.81023
R14394 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n41 1.78522
R14395 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n49 4.56052
R14396 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n38 3.16799
R14397 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n3 2.93012
R14398 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 2.786
R14399 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n0 2.75194
R14400 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n1 2.75094
R14401 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 2.62258
R14402 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n47 1.77011
R14403 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n44 1.76105
R14404 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n57 1.5089
R14405 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n40 1.495
R14406 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN.n11 1.47485
R14407 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n2 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t12 15.4917
R14408 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t14 15.3942
R14409 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t16 14.904
R14410 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t15 14.7749
R14411 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t21 13.6019
R14412 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t18 13.5312
R14413 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t19 13.4877
R14414 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t20 13.227
R14415 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n6 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t13 13.1835
R14416 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n2 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t17 8.17943
R14417 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n0 4.7425
R14418 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t7 3.6405
R14419 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n24 3.6405
R14420 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n16 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t5 3.6405
R14421 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n16 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n15 3.6405
R14422 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t9 3.6405
R14423 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n14 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n13 3.6405
R14424 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t11 3.6405
R14425 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n23 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n22 3.6405
R14426 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n21 3.50463
R14427 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n28 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n19 3.50463
R14428 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t1 3.2765
R14429 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n20 3.2765
R14430 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n19 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.t0 3.2765
R14431 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n19 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n18 3.2765
R14432 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n17 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n14 3.06224
R14433 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n23 3.06224
R14434 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n17 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n16 2.6005
R14435 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n25 2.6005
R14436 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT 2.28587
R14437 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n12 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n1 2.2505
R14438 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n4 1.5982
R14439 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n10 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n8 1.18336
R14440 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n10 0.961395
R14441 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n11 0.806561
R14442 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n28 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n27 0.798761
R14443 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n0 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT 0.65726
R14444 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n0 0.56461
R14445 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n28 0.539611
R14446 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n2 0.381495
R14447 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n10 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n9 0.37501
R14448 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n4 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n3 0.355126
R14449 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n6 0.31227
R14450 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n6 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n5 0.298874
R14451 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n7 0.233052
R14452 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n28 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n17 0.18637
R14453 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n26 0.18637
R14454 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT.n12 0.185454
R14455 VCTRL2.n124 VCTRL2.n123 10.0043
R14456 VCTRL2.n124 VCTRL2.n61 9.34779
R14457 VCTRL2.n53 VCTRL2.t66 8.213
R14458 VCTRL2.n26 VCTRL2.t30 8.213
R14459 VCTRL2.n112 VCTRL2.t12 8.16955
R14460 VCTRL2.n99 VCTRL2.t36 8.16955
R14461 VCTRL2.n33 VCTRL2.t23 8.16955
R14462 VCTRL2.n18 VCTRL2.t16 8.16955
R14463 VCTRL2.n22 VCTRL2.t24 8.16955
R14464 VCTRL2.n58 VCTRL2.t34 8.16955
R14465 VCTRL2.n88 VCTRL2.t22 8.1261
R14466 VCTRL2.n81 VCTRL2.t26 8.1261
R14467 VCTRL2.n95 VCTRL2.t17 8.1261
R14468 VCTRL2.n117 VCTRL2.t0 8.1261
R14469 VCTRL2.n44 VCTRL2.t11 8.1261
R14470 VCTRL2.n13 VCTRL2.t67 8.1261
R14471 VCTRL2.n75 VCTRL2.t9 8.08264
R14472 VCTRL2.n67 VCTRL2.t72 8.08264
R14473 VCTRL2.n49 VCTRL2.t15 7.51776
R14474 VCTRL2.n24 VCTRL2.t70 7.51776
R14475 VCTRL2.n108 VCTRL2.t13 7.47431
R14476 VCTRL2.n97 VCTRL2.t44 7.47431
R14477 VCTRL2.n56 VCTRL2.t74 7.47431
R14478 VCTRL2.n29 VCTRL2.t60 7.47431
R14479 VCTRL2.n15 VCTRL2.t54 7.47431
R14480 VCTRL2.n51 VCTRL2.t2 7.47431
R14481 VCTRL2.n20 VCTRL2.t61 7.47431
R14482 VCTRL2.n25 VCTRL2.t48 7.47431
R14483 VCTRL2.n85 VCTRL2.t49 7.43086
R14484 VCTRL2.n78 VCTRL2.t59 7.43086
R14485 VCTRL2.n111 VCTRL2.t1 7.43086
R14486 VCTRL2.n92 VCTRL2.t75 7.43086
R14487 VCTRL2.n115 VCTRL2.t19 7.43086
R14488 VCTRL2.n98 VCTRL2.t27 7.43086
R14489 VCTRL2.n30 VCTRL2.t38 7.43086
R14490 VCTRL2.n16 VCTRL2.t32 7.43086
R14491 VCTRL2.n41 VCTRL2.t45 7.43086
R14492 VCTRL2.n5 VCTRL2.t18 7.43086
R14493 VCTRL2.n21 VCTRL2.t39 7.43086
R14494 VCTRL2.n57 VCTRL2.t51 7.43086
R14495 VCTRL2.n87 VCTRL2.t33 7.3874
R14496 VCTRL2.n80 VCTRL2.t40 7.3874
R14497 VCTRL2.n72 VCTRL2.t8 7.3874
R14498 VCTRL2.n65 VCTRL2.t31 7.3874
R14499 VCTRL2.n93 VCTRL2.t57 7.3874
R14500 VCTRL2.n116 VCTRL2.t7 7.3874
R14501 VCTRL2.n42 VCTRL2.t25 7.3874
R14502 VCTRL2.n11 VCTRL2.t3 7.3874
R14503 VCTRL2.n74 VCTRL2.t73 7.34395
R14504 VCTRL2.n66 VCTRL2.t14 7.34395
R14505 VCTRL2.n76 VCTRL2.t62 7.3005
R14506 VCTRL2.n68 VCTRL2.t42 7.3005
R14507 VCTRL2.n96 VCTRL2.t76 7.25705
R14508 VCTRL2.n89 VCTRL2.t79 7.25705
R14509 VCTRL2.n82 VCTRL2.t4 7.25705
R14510 VCTRL2.t9 VCTRL2.n74 7.25705
R14511 VCTRL2.t72 VCTRL2.n66 7.25705
R14512 VCTRL2.n118 VCTRL2.t52 7.25705
R14513 VCTRL2.n45 VCTRL2.t28 7.25705
R14514 VCTRL2.n14 VCTRL2.t6 7.25705
R14515 VCTRL2.n100 VCTRL2.t10 7.2136
R14516 VCTRL2.t22 VCTRL2.n87 7.2136
R14517 VCTRL2.t26 VCTRL2.n80 7.2136
R14518 VCTRL2.t73 VCTRL2.n72 7.2136
R14519 VCTRL2.t14 VCTRL2.n65 7.2136
R14520 VCTRL2.n113 VCTRL2.t69 7.2136
R14521 VCTRL2.t17 VCTRL2.n93 7.2136
R14522 VCTRL2.t0 VCTRL2.n116 7.2136
R14523 VCTRL2.n34 VCTRL2.t41 7.2136
R14524 VCTRL2.n19 VCTRL2.t35 7.2136
R14525 VCTRL2.t11 VCTRL2.n42 7.2136
R14526 VCTRL2.t67 VCTRL2.n11 7.2136
R14527 VCTRL2.n23 VCTRL2.t43 7.2136
R14528 VCTRL2.n59 VCTRL2.t55 7.2136
R14529 VCTRL2.t33 VCTRL2.n85 7.17014
R14530 VCTRL2.t40 VCTRL2.n78 7.17014
R14531 VCTRL2.t12 VCTRL2.n111 7.17014
R14532 VCTRL2.t57 VCTRL2.n92 7.17014
R14533 VCTRL2.t7 VCTRL2.n115 7.17014
R14534 VCTRL2.t36 VCTRL2.n98 7.17014
R14535 VCTRL2.t23 VCTRL2.n30 7.17014
R14536 VCTRL2.t16 VCTRL2.n16 7.17014
R14537 VCTRL2.t25 VCTRL2.n41 7.17014
R14538 VCTRL2.t3 VCTRL2.n5 7.17014
R14539 VCTRL2.n54 VCTRL2.t5 7.17014
R14540 VCTRL2.t24 VCTRL2.n21 7.17014
R14541 VCTRL2.t34 VCTRL2.n57 7.17014
R14542 VCTRL2.n27 VCTRL2.t50 7.17014
R14543 VCTRL2.t1 VCTRL2.n108 7.12669
R14544 VCTRL2.t27 VCTRL2.n97 7.12669
R14545 VCTRL2.t38 VCTRL2.n29 7.12669
R14546 VCTRL2.t32 VCTRL2.n15 7.12669
R14547 VCTRL2.t66 VCTRL2.n51 7.12669
R14548 VCTRL2.t39 VCTRL2.n20 7.12669
R14549 VCTRL2.t51 VCTRL2.n56 7.12669
R14550 VCTRL2.t30 VCTRL2.n25 7.12669
R14551 VCTRL2.t2 VCTRL2.n49 7.08324
R14552 VCTRL2.n54 VCTRL2.t20 7.08324
R14553 VCTRL2.t48 VCTRL2.n24 7.08324
R14554 VCTRL2.n27 VCTRL2.t71 7.08324
R14555 VCTRL2.n113 VCTRL2.t53 7.03979
R14556 VCTRL2.n100 VCTRL2.t78 7.03979
R14557 VCTRL2.n34 VCTRL2.t63 7.03979
R14558 VCTRL2.n19 VCTRL2.t56 7.03979
R14559 VCTRL2.n23 VCTRL2.t64 7.03979
R14560 VCTRL2.n59 VCTRL2.t77 7.03979
R14561 VCTRL2.n96 VCTRL2.t58 6.99633
R14562 VCTRL2.n89 VCTRL2.t65 6.99633
R14563 VCTRL2.n82 VCTRL2.t68 6.99633
R14564 VCTRL2.n118 VCTRL2.t37 6.99633
R14565 VCTRL2.n45 VCTRL2.t47 6.99633
R14566 VCTRL2.n14 VCTRL2.t21 6.99633
R14567 VCTRL2.n76 VCTRL2.t46 6.95288
R14568 VCTRL2.n68 VCTRL2.t29 6.95288
R14569 VCTRL2.t46 VCTRL2.n75 6.51836
R14570 VCTRL2.t29 VCTRL2.n67 6.51836
R14571 VCTRL2.t58 VCTRL2.n95 6.4749
R14572 VCTRL2.t65 VCTRL2.n88 6.4749
R14573 VCTRL2.t68 VCTRL2.n81 6.4749
R14574 VCTRL2.t37 VCTRL2.n117 6.4749
R14575 VCTRL2.t47 VCTRL2.n44 6.4749
R14576 VCTRL2.t21 VCTRL2.n13 6.4749
R14577 VCTRL2.t53 VCTRL2.n112 6.43145
R14578 VCTRL2.t78 VCTRL2.n99 6.43145
R14579 VCTRL2.t63 VCTRL2.n33 6.43145
R14580 VCTRL2.t56 VCTRL2.n18 6.43145
R14581 VCTRL2.t64 VCTRL2.n22 6.43145
R14582 VCTRL2.t77 VCTRL2.n58 6.43145
R14583 VCTRL2.t20 VCTRL2.n53 6.388
R14584 VCTRL2.t71 VCTRL2.n26 6.388
R14585 VCTRL2.n28 VCTRL2.n27 4.03166
R14586 VCTRL2.n101 VCTRL2.n100 4.0306
R14587 VCTRL2.n119 VCTRL2.n118 3.63007
R14588 VCTRL2.n60 VCTRL2.n59 3.62933
R14589 VCTRL2.n11 VCTRL2.n10 3.62499
R14590 VCTRL2.n102 VCTRL2.n89 3.62466
R14591 VCTRL2.n88 VCTRL2.n83 3.62466
R14592 VCTRL2.n108 VCTRL2.n107 3.62466
R14593 VCTRL2.n5 VCTRL2.n4 3.62466
R14594 VCTRL2.n41 VCTRL2.n40 3.62466
R14595 VCTRL2.n28 VCTRL2.n23 3.62466
R14596 VCTRL2.n36 VCTRL2.n19 3.62466
R14597 VCTRL2.n47 VCTRL2.n14 3.62466
R14598 VCTRL2.n85 VCTRL2.n84 3.62466
R14599 VCTRL2.n87 VCTRL2.n86 3.62466
R14600 VCTRL2.n112 VCTRL2.n106 3.62466
R14601 VCTRL2.n114 VCTRL2.n113 3.62466
R14602 VCTRL2.n111 VCTRL2.n110 3.62466
R14603 VCTRL2.n18 VCTRL2.n17 3.62466
R14604 VCTRL2.n44 VCTRL2.n43 3.62466
R14605 VCTRL2.n46 VCTRL2.n45 3.62466
R14606 VCTRL2.n13 VCTRL2.n12 3.62466
R14607 VCTRL2.n101 VCTRL2.n96 3.62462
R14608 VCTRL2.n103 VCTRL2.n82 3.62462
R14609 VCTRL2.n78 VCTRL2.n77 3.62462
R14610 VCTRL2.n80 VCTRL2.n79 3.62462
R14611 VCTRL2.n75 VCTRL2.n70 3.62462
R14612 VCTRL2.n104 VCTRL2.n76 3.62462
R14613 VCTRL2.n72 VCTRL2.n71 3.62462
R14614 VCTRL2.n74 VCTRL2.n73 3.62462
R14615 VCTRL2.n67 VCTRL2.n63 3.62462
R14616 VCTRL2.n105 VCTRL2.n68 3.62462
R14617 VCTRL2.n65 VCTRL2.n64 3.62462
R14618 VCTRL2.n93 VCTRL2.n90 3.62462
R14619 VCTRL2.n92 VCTRL2.n91 3.62462
R14620 VCTRL2.n95 VCTRL2.n94 3.62462
R14621 VCTRL2.n33 VCTRL2.n32 3.62462
R14622 VCTRL2.n35 VCTRL2.n34 3.62462
R14623 VCTRL2.n49 VCTRL2.n48 3.62462
R14624 VCTRL2.n53 VCTRL2.n52 3.62462
R14625 VCTRL2.n55 VCTRL2.n54 3.62462
R14626 VCTRL2.n51 VCTRL2.n50 3.62462
R14627 VCTRL2.n122 VCTRL2.n121 2.2505
R14628 VCTRL2.n3 VCTRL2.n2 2.2505
R14629 VCTRL2.n125 VCTRL2.n124 1.5049
R14630 VCTRL2 VCTRL2.n0 1.16594
R14631 VCTRL2 VCTRL2.n62 1.16341
R14632 VCTRL2.n122 VCTRL2.n119 1.05045
R14633 VCTRL2.n61 VCTRL2.n60 0.984409
R14634 VCTRL2.n120 VCTRL2 0.936261
R14635 VCTRL2.n1 VCTRL2 0.936261
R14636 VCTRL2.n125 VCTRL2 0.61117
R14637 VCTRL2.n119 VCTRL2.n114 0.442081
R14638 VCTRL2.n60 VCTRL2.n55 0.441056
R14639 VCTRL2.n8 VCTRL2.n7 0.404715
R14640 VCTRL2.n36 VCTRL2.n35 0.404715
R14641 VCTRL2.n103 VCTRL2.n102 0.404539
R14642 VCTRL2.n39 VCTRL2.n38 0.404539
R14643 VCTRL2.n46 VCTRL2.n36 0.401155
R14644 VCTRL2.n9 VCTRL2.n8 0.401155
R14645 VCTRL2.n40 VCTRL2.n39 0.401155
R14646 VCTRL2.n104 VCTRL2.n103 0.400353
R14647 VCTRL2.n70 VCTRL2.n69 0.400178
R14648 VCTRL2.n47 VCTRL2.n46 0.398905
R14649 VCTRL2.n10 VCTRL2.n9 0.398484
R14650 VCTRL2.n55 VCTRL2.n47 0.397919
R14651 VCTRL2.n114 VCTRL2.n105 0.397919
R14652 VCTRL2.n105 VCTRL2.n104 0.397753
R14653 VCTRL2.n110 VCTRL2.n109 0.397744
R14654 VCTRL2.n7 VCTRL2.n6 0.389969
R14655 VCTRL2.n102 VCTRL2.n101 0.389723
R14656 VCTRL2.n38 VCTRL2.n37 0.389723
R14657 VCTRL2.n35 VCTRL2.n28 0.389547
R14658 VCTRL2.n32 VCTRL2.n31 0.389547
R14659 VCTRL2 VCTRL2.n125 0.10046
R14660 VCTRL2.n123 VCTRL2.n62 0.0698976
R14661 VCTRL2.n3 VCTRL2.n0 0.0695909
R14662 VCTRL2.n121 VCTRL2 0.0362534
R14663 VCTRL2.n2 VCTRL2 0.0362534
R14664 VCTRL2.n123 VCTRL2.n122 0.0124277
R14665 VCTRL2.n61 VCTRL2.n3 0.00395428
R14666 VCTRL2.n121 VCTRL2.n120 0.00173288
R14667 VCTRL2.n2 VCTRL2.n1 0.00173288
R14668 a_25706_n567.n90 a_25706_n567.n89 9.67588
R14669 a_25706_n567.n42 a_25706_n567.n41 3.74413
R14670 a_25706_n567.n26 a_25706_n567.n25 3.74025
R14671 a_25706_n567.n8 a_25706_n567.n12 3.72928
R14672 a_25706_n567.n9 a_25706_n567.n14 3.71799
R14673 a_25706_n567.n7 a_25706_n567.n6 3.60834
R14674 a_25706_n567.n21 a_25706_n567.t53 3.2765
R14675 a_25706_n567.n21 a_25706_n567.n20 3.2765
R14676 a_25706_n567.n23 a_25706_n567.t46 3.2765
R14677 a_25706_n567.n23 a_25706_n567.n22 3.2765
R14678 a_25706_n567.n70 a_25706_n567.t56 3.2765
R14679 a_25706_n567.n70 a_25706_n567.n69 3.2765
R14680 a_25706_n567.n67 a_25706_n567.t3 3.2765
R14681 a_25706_n567.n67 a_25706_n567.n66 3.2765
R14682 a_25706_n567.n63 a_25706_n567.t58 3.2765
R14683 a_25706_n567.n63 a_25706_n567.n62 3.2765
R14684 a_25706_n567.n60 a_25706_n567.t11 3.2765
R14685 a_25706_n567.n60 a_25706_n567.n59 3.2765
R14686 a_25706_n567.n56 a_25706_n567.t1 3.2765
R14687 a_25706_n567.n56 a_25706_n567.n55 3.2765
R14688 a_25706_n567.n87 a_25706_n567.t9 3.2765
R14689 a_25706_n567.n87 a_25706_n567.n86 3.2765
R14690 a_25706_n567.n84 a_25706_n567.t13 3.2765
R14691 a_25706_n567.n84 a_25706_n567.n83 3.2765
R14692 a_25706_n567.n80 a_25706_n567.t7 3.2765
R14693 a_25706_n567.n80 a_25706_n567.n79 3.2765
R14694 a_25706_n567.n77 a_25706_n567.t8 3.2765
R14695 a_25706_n567.n77 a_25706_n567.n76 3.2765
R14696 a_25706_n567.n73 a_25706_n567.t12 3.2765
R14697 a_25706_n567.n73 a_25706_n567.n72 3.2765
R14698 a_25706_n567.n36 a_25706_n567.t50 3.2765
R14699 a_25706_n567.n36 a_25706_n567.n35 3.2765
R14700 a_25706_n567.n34 a_25706_n567.t19 3.2765
R14701 a_25706_n567.n34 a_25706_n567.n33 3.2765
R14702 a_25706_n567.n30 a_25706_n567.t49 3.2765
R14703 a_25706_n567.n30 a_25706_n567.n29 3.2765
R14704 a_25706_n567.n28 a_25706_n567.t31 3.2765
R14705 a_25706_n567.n28 a_25706_n567.n27 3.2765
R14706 a_25706_n567.n19 a_25706_n567.t28 3.2765
R14707 a_25706_n567.n19 a_25706_n567.n18 3.2765
R14708 a_25706_n567.n12 a_25706_n567.t21 3.2765
R14709 a_25706_n567.n12 a_25706_n567.n11 3.2765
R14710 a_25706_n567.n16 a_25706_n567.t16 3.2765
R14711 a_25706_n567.n16 a_25706_n567.n15 3.2765
R14712 a_25706_n567.n14 a_25706_n567.t48 3.2765
R14713 a_25706_n567.n14 a_25706_n567.n13 3.2765
R14714 a_25706_n567.n4 a_25706_n567.t36 3.2765
R14715 a_25706_n567.n4 a_25706_n567.n3 3.2765
R14716 a_25706_n567.n39 a_25706_n567.t37 3.2765
R14717 a_25706_n567.n39 a_25706_n567.n38 3.2765
R14718 a_25706_n567.n46 a_25706_n567.t42 3.2765
R14719 a_25706_n567.n46 a_25706_n567.n45 3.2765
R14720 a_25706_n567.n44 a_25706_n567.t23 3.2765
R14721 a_25706_n567.n44 a_25706_n567.n43 3.2765
R14722 a_25706_n567.n41 a_25706_n567.t15 3.2765
R14723 a_25706_n567.n41 a_25706_n567.n40 3.2765
R14724 a_25706_n567.n49 a_25706_n567.t30 3.2765
R14725 a_25706_n567.n49 a_25706_n567.n48 3.2765
R14726 a_25706_n567.n2 a_25706_n567.t40 3.2765
R14727 a_25706_n567.n2 a_25706_n567.n1 3.2765
R14728 a_25706_n567.n52 a_25706_n567.t32 3.2765
R14729 a_25706_n567.n52 a_25706_n567.n51 3.2765
R14730 a_25706_n567.n25 a_25706_n567.t24 3.2765
R14731 a_25706_n567.n25 a_25706_n567.n24 3.2765
R14732 a_25706_n567.n94 a_25706_n567.t47 3.2765
R14733 a_25706_n567.n95 a_25706_n567.n94 3.2765
R14734 a_25706_n567.n74 a_25706_n567.n73 3.1505
R14735 a_25706_n567.n78 a_25706_n567.n77 3.1505
R14736 a_25706_n567.n81 a_25706_n567.n80 3.1505
R14737 a_25706_n567.n85 a_25706_n567.n84 3.1505
R14738 a_25706_n567.n88 a_25706_n567.n87 3.1505
R14739 a_25706_n567.n57 a_25706_n567.n56 3.1505
R14740 a_25706_n567.n61 a_25706_n567.n60 3.1505
R14741 a_25706_n567.n64 a_25706_n567.n63 3.1505
R14742 a_25706_n567.n68 a_25706_n567.n67 3.1505
R14743 a_25706_n567.n71 a_25706_n567.n70 3.1505
R14744 a_25706_n567.n47 a_25706_n567.n46 3.1505
R14745 a_25706_n567.n50 a_25706_n567.n49 3.1505
R14746 a_25706_n567.n53 a_25706_n567.n52 3.1505
R14747 a_25706_n567.n5 a_25706_n567.n4 3.1505
R14748 a_25706_n567.n31 a_25706_n567.n30 3.1505
R14749 a_25706_n567.n37 a_25706_n567.n36 3.1505
R14750 a_25706_n567.n92 a_25706_n567.n23 3.1505
R14751 a_25706_n567.n94 a_25706_n567.n93 3.1505
R14752 a_25706_n567.n17 a_25706_n567.n10 2.34866
R14753 a_25706_n567.n8 a_25706_n567.n19 1.8475
R14754 a_25706_n567.n42 a_25706_n567.n44 1.84743
R14755 a_25706_n567.n6 a_25706_n567.n2 1.84743
R14756 a_25706_n567.n26 a_25706_n567.n28 1.8474
R14757 a_25706_n567.n0 a_25706_n567.n39 1.84737
R14758 a_25706_n567.n32 a_25706_n567.n34 1.84737
R14759 a_25706_n567.n7 a_25706_n567.n21 1.84737
R14760 a_25706_n567.n10 a_25706_n567.n16 1.84618
R14761 a_25706_n567.n8 a_25706_n567.n17 1.48093
R14762 a_25706_n567.n54 a_25706_n567.n53 0.899822
R14763 a_25706_n567.n92 a_25706_n567.n91 0.899822
R14764 a_25706_n567.n81 a_25706_n567.n78 0.758798
R14765 a_25706_n567.n64 a_25706_n567.n61 0.758798
R14766 a_25706_n567.n89 a_25706_n567.n71 0.724996
R14767 a_25706_n567.n88 a_25706_n567.n85 0.7205
R14768 a_25706_n567.n71 a_25706_n567.n68 0.7205
R14769 a_25706_n567.n89 a_25706_n567.n88 0.636952
R14770 a_25706_n567.n93 a_25706_n567.n8 0.618999
R14771 a_25706_n567.n50 a_25706_n567.n0 0.607482
R14772 a_25706_n567.n37 a_25706_n567.n32 0.604163
R14773 a_25706_n567.n7 a_25706_n567.n92 0.60198
R14774 a_25706_n567.n93 a_25706_n567.n7 0.601843
R14775 a_25706_n567.n32 a_25706_n567.n31 0.598752
R14776 a_25706_n567.n31 a_25706_n567.n26 0.597003
R14777 a_25706_n567.n0 a_25706_n567.n47 0.595434
R14778 a_25706_n567.n47 a_25706_n567.n42 0.593116
R14779 a_25706_n567.n6 a_25706_n567.n5 0.593116
R14780 a_25706_n567.n75 a_25706_n567.n74 0.555819
R14781 a_25706_n567.n58 a_25706_n567.n57 0.555819
R14782 a_25706_n567.n85 a_25706_n567.n82 0.551989
R14783 a_25706_n567.n68 a_25706_n567.n65 0.551989
R14784 a_25706_n567.n90 a_25706_n567.n54 0.3917
R14785 a_25706_n567.n82 a_25706_n567.n81 0.283904
R14786 a_25706_n567.n65 a_25706_n567.n64 0.283904
R14787 a_25706_n567.n78 a_25706_n567.n75 0.280074
R14788 a_25706_n567.n61 a_25706_n567.n58 0.280074
R14789 a_25706_n567.n91 a_25706_n567.n90 0.2621
R14790 a_25706_n567.n54 a_25706_n567.n50 0.247022
R14791 a_25706_n567.n91 a_25706_n567.n37 0.247022
R14792 a_25706_n567.n10 a_25706_n567.n9 0.0460206
R14793 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n8 15.8172
R14794 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n10 15.8172
R14795 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n9 15.8172
R14796 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t37 14.8925
R14797 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t43 14.8925
R14798 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n16 12.2457
R14799 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n14 12.2457
R14800 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n12 12.2457
R14801 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t58 11.6285
R14802 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t41 9.5787
R14803 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t45 9.55768
R14804 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t56 8.9065
R14805 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t42 8.9065
R14806 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t47 8.9065
R14807 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t35 8.9065
R14808 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n64 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n60 8.86038
R14809 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t33 8.6145
R14810 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t46 8.6145
R14811 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t39 8.6145
R14812 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t54 8.59715
R14813 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t52 8.57144
R14814 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t57 8.57144
R14815 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n54 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t50 8.57144
R14816 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t5 8.54728
R14817 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t38 8.52112
R14818 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t53 8.52112
R14819 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t32 8.52112
R14820 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t48 8.52112
R14821 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n51 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t55 8.51092
R14822 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t34 8.51092
R14823 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t31 8.51092
R14824 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t40 8.35286
R14825 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t49 8.3225
R14826 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t58 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n17 8.3225
R14827 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t36 8.31073
R14828 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t44 8.31073
R14829 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t51 8.31073
R14830 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n22 7.05764
R14831 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t30 6.83153
R14832 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t25 6.78441
R14833 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n35 6.45366
R14834 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n28 6.20932
R14835 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t26 5.87174
R14836 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n76 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t20 5.30249
R14837 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n42 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n41 5.28839
R14838 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t19 4.92134
R14839 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n58 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t13 4.89657
R14840 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n44 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t16 4.89616
R14841 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n36 4.87698
R14842 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n57 4.63042
R14843 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n56 4.63037
R14844 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n45 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n1 4.22693
R14845 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n18 4.223
R14846 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n46 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n42 4.02972
R14847 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n33 4.0288
R14848 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n73 3.96222
R14849 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t42 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n13 3.6505
R14850 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n15 3.6505
R14851 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n62 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t9 3.6405
R14852 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n62 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n61 3.6405
R14853 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n78 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t17 3.6405
R14854 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n78 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n79 3.6405
R14855 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t14 3.6405
R14856 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n37 3.6405
R14857 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t22 3.6405
R14858 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n32 3.6405
R14859 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t10 3.6405
R14860 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n66 3.6405
R14861 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n23 3.47613
R14862 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n19 3.47609
R14863 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n25 3.47601
R14864 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n20 3.39857
R14865 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n45 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n77 3.27464
R14866 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n11 3.1807
R14867 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n75 3.16877
R14868 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n76 2.96981
R14869 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t0 2.8627
R14870 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t4 2.86263
R14871 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.t28 2.8626
R14872 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n68 2.60609
R14873 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n24 2.48343
R14874 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 2.30073
R14875 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n75 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 2.29178
R14876 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n27 2.24606
R14877 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n69 2.24505
R14878 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n67 4.81682
R14879 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n64 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n63 3.77141
R14880 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n44 2.52627
R14881 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n59 1.8072
R14882 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n40 1.76824
R14883 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n63 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n62 1.65829
R14884 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n38 1.65829
R14885 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n51 1.6131
R14886 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n54 1.57488
R14887 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n44 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n43 1.53436
R14888 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n70 1.51602
R14889 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n58 1.49487
R14890 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n34 1.32452
R14891 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n77 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n78 1.25757
R14892 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n39 1.12313
R14893 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n4 1.05601
R14894 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n29 1.01067
R14895 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n49 0.996664
R14896 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n5 0.992966
R14897 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n21 0.983287
R14898 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n26 0.982856
R14899 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n0 0.975705
R14900 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n72 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n71 0.968726
R14901 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n72 0.955885
R14902 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n52 0.953514
R14903 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n3 0.911933
R14904 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n46 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n45 0.856289
R14905 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n47 0.843442
R14906 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n65 0.8015
R14907 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n6 0.741046
R14908 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n31 0.710717
R14909 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n7 0.698938
R14910 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n72 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n48 0.656959
R14911 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n46 0.398395
R14912 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n64 0.3875
R14913 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n54 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n53 0.364199
R14914 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n30 0.362023
R14915 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n2 0.359267
R14916 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n51 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n50 0.323514
R14917 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n55 0.321048
R14918 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n75 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n74 0.271283
R14919 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 0.147028
R14920 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n72 15.8172
R14921 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n73 15.8172
R14922 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n75 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n74 15.8172
R14923 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t50 14.8925
R14924 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t43 14.8925
R14925 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n81 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n80 12.2457
R14926 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n80 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n78 12.2457
R14927 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n78 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n76 12.2457
R14928 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n82 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t37 11.6285
R14929 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t35 9.07401
R14930 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t45 8.94931
R14931 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t32 8.91612
R14932 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t58 8.91612
R14933 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t40 8.91612
R14934 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n76 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t54 8.9065
R14935 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n78 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t47 8.9065
R14936 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n80 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t36 8.9065
R14937 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n81 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t57 8.9065
R14938 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t53 8.88203
R14939 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t42 8.78079
R14940 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t39 8.78079
R14941 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t46 8.76459
R14942 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t44 8.76459
R14943 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n9 8.71932
R14944 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t55 8.71352
R14945 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t51 8.71352
R14946 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n73 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t49 8.6145
R14947 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n72 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t56 8.6145
R14948 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n74 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t38 8.6145
R14949 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n75 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t31 8.59715
R14950 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t0 8.51681
R14951 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t41 8.50287
R14952 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t52 8.38543
R14953 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n76 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t33 8.3225
R14954 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t37 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n81 8.3225
R14955 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t34 8.30117
R14956 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n6 8.23463
R14957 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t48 7.39905
R14958 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n25 6.43594
R14959 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n19 6.42269
R14960 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n27 6.3977
R14961 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n33 6.02773
R14962 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t20 5.83006
R14963 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n66 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n52 5.43818
R14964 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n14 5.23259
R14965 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n64 4.89653
R14966 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n42 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t15 4.89315
R14967 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t27 4.88822
R14968 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n10 4.72831
R14969 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t19 4.70462
R14970 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t22 4.70346
R14971 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n48 4.53146
R14972 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n82 4.22145
R14973 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t5 4.04969
R14974 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n60 4.00854
R14975 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n44 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n43 4.00757
R14976 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t6 4.00481
R14977 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n8 3.90715
R14978 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n70 3.79925
R14979 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n16 3.77445
R14980 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n46 3.76989
R14981 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n24 3.76191
R14982 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t30 3.7183
R14983 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n77 3.6505
R14984 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t36 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n79 3.6505
R14985 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n62 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t11 3.6405
R14986 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n62 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n61 3.6405
R14987 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n57 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t8 3.6405
R14988 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n57 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n56 3.6405
R14989 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t12 3.6405
R14990 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n51 3.6405
R14991 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t21 3.47629
R14992 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t18 3.47627
R14993 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n20 3.3208
R14994 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.t2 3.26228
R14995 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n23 3.25601
R14996 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n82 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n75 3.1807
R14997 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 3.15982
R14998 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n22 3.14573
R14999 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n59 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n58 2.8959
R15000 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n17 2.88663
R15001 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n15 2.86148
R15002 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n13 2.86147
R15003 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n12 2.83772
R15004 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n49 2.75932
R15005 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n66 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n7 2.62155
R15006 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 2.36584
R15007 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n69 2.35159
R15008 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 2.30603
R15009 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n45 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n44 2.2491
R15010 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n54 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n55 2.24586
R15011 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n67 2.03309
R15012 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n71 1.93478
R15013 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n45 1.85135
R15014 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n63 1.79127
R15015 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n54 1.76701
R15016 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n58 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n57 1.65928
R15017 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n53 1.6295
R15018 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n29 1.50938
R15019 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n63 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n65 1.495
R15020 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n28 1.47463
R15021 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n60 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n62 1.25653
R15022 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n66 1.22576
R15023 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n4 1.19023
R15024 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n59 1.1585
R15025 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n42 1.1379
R15026 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n47 1.00671
R15027 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n28 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n5 0.931417
R15028 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n26 0.878898
R15029 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n50 0.836865
R15030 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n38 0.650226
R15031 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n68 0.597881
R15032 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n21 0.488268
R15033 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n32 0.487486
R15034 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n11 0.477758
R15035 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n18 0.472393
R15036 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n0 0.415098
R15037 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n1 0.384677
R15038 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n3 0.384538
R15039 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n40 0.345705
R15040 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n30 0.345705
R15041 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n41 0.34324
R15042 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n36 0.342007
R15043 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n34 0.342007
R15044 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n2 0.33461
R15045 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n37 0.325979
R15046 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n39 0.318582
R15047 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n31 0.312418
R15048 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN.n35 0.312418
R15049 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n23 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t18 23.6945
R15050 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t20 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n24 23.6945
R15051 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n24 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n23 18.8035
R15052 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n19 15.8172
R15053 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n20 15.8172
R15054 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n16 15.8172
R15055 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n19 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t13 14.8925
R15056 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t21 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n21 14.8925
R15057 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t16 14.8925
R15058 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n17 12.2457
R15059 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n17 12.2457
R15060 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n18 12.2457
R15061 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t15 11.6285
R15062 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n18 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t18 8.9065
R15063 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t17 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n22 8.9065
R15064 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t22 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n17 8.9065
R15065 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t20 8.9065
R15066 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n21 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t19 8.6145
R15067 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n19 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t23 8.6145
R15068 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t14 8.6145
R15069 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n16 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t12 8.59715
R15070 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t13 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n18 8.3225
R15071 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t21 8.3225
R15072 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t16 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n17 8.3225
R15073 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t15 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n25 8.3225
R15074 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n26 4.223
R15075 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n23 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t17 3.6505
R15076 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n24 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t22 3.6505
R15077 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t7 3.6405
R15078 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n10 3.6405
R15079 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t9 3.6405
R15080 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n4 3.6405
R15081 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t4 3.6405
R15082 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n6 3.6405
R15083 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n13 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t6 3.6405
R15084 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n13 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n12 3.6405
R15085 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n1 3.50463
R15086 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n3 3.50463
R15087 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t1 3.2765
R15088 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n0 3.2765
R15089 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.t3 3.2765
R15090 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n2 3.2765
R15091 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n16 3.1807
R15092 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n7 3.06224
R15093 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n14 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n11 3.06224
R15094 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n5 2.6005
R15095 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n14 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n13 2.6005
R15096 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n9 0.798761
R15097 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n15 0.562022
R15098 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n8 0.18637
R15099 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT.n14 0.18637
R15100 a_50630_6066.n26 a_50630_6066.n25 72.9524
R15101 a_50630_6066.n20 a_50630_6066.t23 44.8231
R15102 a_50630_6066.n2 a_50630_6066.t18 36.4904
R15103 a_50630_6066.n26 a_50630_6066.t28 23.7985
R15104 a_50630_6066.n2 a_50630_6066.t22 23.6525
R15105 a_50630_6066.n3 a_50630_6066.t11 23.6525
R15106 a_50630_6066.n4 a_50630_6066.t7 23.6525
R15107 a_50630_6066.n5 a_50630_6066.t20 23.6525
R15108 a_50630_6066.n6 a_50630_6066.t8 23.6525
R15109 a_50630_6066.n7 a_50630_6066.t16 23.6525
R15110 a_50630_6066.n8 a_50630_6066.t29 23.6525
R15111 a_50630_6066.n9 a_50630_6066.t26 23.6525
R15112 a_50630_6066.n10 a_50630_6066.t14 23.6525
R15113 a_50630_6066.n11 a_50630_6066.t27 23.6525
R15114 a_50630_6066.n12 a_50630_6066.t15 23.6525
R15115 a_50630_6066.n13 a_50630_6066.t19 23.6525
R15116 a_50630_6066.n14 a_50630_6066.t24 23.6525
R15117 a_50630_6066.n15 a_50630_6066.t13 23.6525
R15118 a_50630_6066.n16 a_50630_6066.t25 23.6525
R15119 a_50630_6066.n21 a_50630_6066.n20 23.3438
R15120 a_50630_6066.n22 a_50630_6066.n21 23.3438
R15121 a_50630_6066.n23 a_50630_6066.n22 23.3438
R15122 a_50630_6066.n24 a_50630_6066.n23 23.3438
R15123 a_50630_6066.n25 a_50630_6066.n24 23.3438
R15124 a_50630_6066.n20 a_50630_6066.t12 20.4405
R15125 a_50630_6066.n21 a_50630_6066.t9 20.4405
R15126 a_50630_6066.n22 a_50630_6066.t21 20.4405
R15127 a_50630_6066.n23 a_50630_6066.t10 20.4405
R15128 a_50630_6066.n24 a_50630_6066.t17 20.4405
R15129 a_50630_6066.n25 a_50630_6066.t6 20.4405
R15130 a_50630_6066.n3 a_50630_6066.n2 12.8384
R15131 a_50630_6066.n4 a_50630_6066.n3 12.8384
R15132 a_50630_6066.n5 a_50630_6066.n4 12.8384
R15133 a_50630_6066.n6 a_50630_6066.n5 12.8384
R15134 a_50630_6066.n7 a_50630_6066.n6 12.8384
R15135 a_50630_6066.n8 a_50630_6066.n7 12.8384
R15136 a_50630_6066.n9 a_50630_6066.n8 12.8384
R15137 a_50630_6066.n10 a_50630_6066.n9 12.8384
R15138 a_50630_6066.n11 a_50630_6066.n10 12.8384
R15139 a_50630_6066.n12 a_50630_6066.n11 12.8384
R15140 a_50630_6066.n13 a_50630_6066.n12 12.8384
R15141 a_50630_6066.n14 a_50630_6066.n13 12.8384
R15142 a_50630_6066.n15 a_50630_6066.n14 12.8384
R15143 a_50630_6066.n16 a_50630_6066.n15 12.8384
R15144 a_50630_6066.n27 a_50630_6066.n26 6.95492
R15145 a_50630_6066.n17 a_50630_6066.n16 4.78319
R15146 a_50630_6066.n28 a_50630_6066.n27 4.13676
R15147 a_50630_6066.n27 a_50630_6066.n19 3.79615
R15148 a_50630_6066.n17 a_50630_6066.n1 3.22711
R15149 a_50630_6066.n30 a_50630_6066.n28 3.22482
R15150 a_50630_6066.n1 a_50630_6066.t2 0.6505
R15151 a_50630_6066.n1 a_50630_6066.n0 0.6505
R15152 a_50630_6066.t0 a_50630_6066.n30 0.6505
R15153 a_50630_6066.n30 a_50630_6066.n29 0.6505
R15154 a_50630_6066.n19 a_50630_6066.t4 0.5855
R15155 a_50630_6066.n19 a_50630_6066.n18 0.5855
R15156 a_50630_6066.n28 a_50630_6066.n17 0.471269
R15157 a_50708_569.n67 a_50708_569.t44 40.255
R15158 a_50708_569.n26 a_50708_569.t58 37.7641
R15159 a_50708_569.t104 a_50708_569.n24 30.4352
R15160 a_50708_569.t50 a_50708_569.n42 28.4705
R15161 a_50708_569.t36 a_50708_569.n49 28.4705
R15162 a_50708_569.t35 a_50708_569.n56 28.4705
R15163 a_50708_569.t39 a_50708_569.n63 28.4705
R15164 a_50708_569.t115 a_50708_569.n71 28.4705
R15165 a_50708_569.n75 a_50708_569.t87 27.3249
R15166 a_50708_569.n42 a_50708_569.t52 27.1982
R15167 a_50708_569.t87 a_50708_569.n74 25.4384
R15168 a_50708_569.n74 a_50708_569.t67 25.4384
R15169 a_50708_569.n72 a_50708_569.t32 25.4045
R15170 a_50708_569.n66 a_50708_569.t79 25.4045
R15171 a_50708_569.n66 a_50708_569.t61 25.4045
R15172 a_50708_569.n65 a_50708_569.t107 25.4045
R15173 a_50708_569.n65 a_50708_569.t86 25.4045
R15174 a_50708_569.n57 a_50708_569.t49 25.4045
R15175 a_50708_569.n52 a_50708_569.t72 25.4045
R15176 a_50708_569.n52 a_50708_569.t53 25.4045
R15177 a_50708_569.n51 a_50708_569.t30 25.4045
R15178 a_50708_569.n51 a_50708_569.t110 25.4045
R15179 a_50708_569.n2 a_50708_569.t101 25.4045
R15180 a_50708_569.n2 a_50708_569.t80 25.4045
R15181 a_50708_569.n3 a_50708_569.t46 25.4045
R15182 a_50708_569.n3 a_50708_569.t33 25.4045
R15183 a_50708_569.n4 a_50708_569.t56 25.4045
R15184 a_50708_569.n4 a_50708_569.t40 25.4045
R15185 a_50708_569.n5 a_50708_569.t109 25.4045
R15186 a_50708_569.n5 a_50708_569.t88 25.4045
R15187 a_50708_569.n6 a_50708_569.t81 25.4045
R15188 a_50708_569.n6 a_50708_569.t62 25.4045
R15189 a_50708_569.n7 a_50708_569.t34 25.4045
R15190 a_50708_569.n7 a_50708_569.t116 25.4045
R15191 a_50708_569.n8 a_50708_569.t76 25.4045
R15192 a_50708_569.n8 a_50708_569.t59 25.4045
R15193 a_50708_569.n9 a_50708_569.t89 25.4045
R15194 a_50708_569.n9 a_50708_569.t68 25.4045
R15195 a_50708_569.n10 a_50708_569.t38 25.4045
R15196 a_50708_569.n10 a_50708_569.t26 25.4045
R15197 a_50708_569.n11 a_50708_569.t117 25.4045
R15198 a_50708_569.n11 a_50708_569.t94 25.4045
R15199 a_50708_569.n12 a_50708_569.t60 25.4045
R15200 a_50708_569.n12 a_50708_569.t43 25.4045
R15201 a_50708_569.n13 a_50708_569.t114 25.4045
R15202 a_50708_569.n13 a_50708_569.t93 25.4045
R15203 a_50708_569.n25 a_50708_569.t27 25.4045
R15204 a_50708_569.n25 a_50708_569.t104 25.4045
R15205 a_50708_569.n43 a_50708_569.t66 25.4045
R15206 a_50708_569.n38 a_50708_569.t97 25.4045
R15207 a_50708_569.n36 a_50708_569.t45 25.4045
R15208 a_50708_569.n36 a_50708_569.t111 25.4045
R15209 a_50708_569.n38 a_50708_569.t28 25.4045
R15210 a_50708_569.n40 a_50708_569.t75 25.4045
R15211 a_50708_569.n40 a_50708_569.t108 25.4045
R15212 a_50708_569.n41 a_50708_569.t119 25.4045
R15213 a_50708_569.t52 a_50708_569.n41 25.4045
R15214 a_50708_569.n43 a_50708_569.t50 25.4045
R15215 a_50708_569.n44 a_50708_569.t25 25.4045
R15216 a_50708_569.n44 a_50708_569.t102 25.4045
R15217 a_50708_569.n45 a_50708_569.t65 25.4045
R15218 a_50708_569.n45 a_50708_569.t47 25.4045
R15219 a_50708_569.n50 a_50708_569.t51 25.4045
R15220 a_50708_569.n50 a_50708_569.t36 25.4045
R15221 a_50708_569.n57 a_50708_569.t35 25.4045
R15222 a_50708_569.n58 a_50708_569.t100 25.4045
R15223 a_50708_569.n58 a_50708_569.t77 25.4045
R15224 a_50708_569.n59 a_50708_569.t82 25.4045
R15225 a_50708_569.n59 a_50708_569.t63 25.4045
R15226 a_50708_569.n64 a_50708_569.t54 25.4045
R15227 a_50708_569.n64 a_50708_569.t39 25.4045
R15228 a_50708_569.n72 a_50708_569.t115 25.4045
R15229 a_50708_569.n73 a_50708_569.t118 25.4045
R15230 a_50708_569.n73 a_50708_569.t95 25.4045
R15231 a_50708_569.n48 a_50708_569.t31 23.6525
R15232 a_50708_569.n55 a_50708_569.t37 23.6525
R15233 a_50708_569.n62 a_50708_569.t42 23.6525
R15234 a_50708_569.n70 a_50708_569.t24 23.6525
R15235 a_50708_569.n75 a_50708_569.t78 23.5689
R15236 a_50708_569.n76 a_50708_569.t106 23.5065
R15237 a_50708_569.n77 a_50708_569.t29 23.5065
R15238 a_50708_569.n78 a_50708_569.t70 23.5065
R15239 a_50708_569.n79 a_50708_569.t99 23.5065
R15240 a_50708_569.n80 a_50708_569.t48 23.5065
R15241 a_50708_569.n81 a_50708_569.t71 23.5065
R15242 a_50708_569.n82 a_50708_569.t92 23.5065
R15243 a_50708_569.n27 a_50708_569.t55 22.4115
R15244 a_50708_569.n26 a_50708_569.t69 22.4115
R15245 a_50708_569.n47 a_50708_569.t74 20.4405
R15246 a_50708_569.n46 a_50708_569.t105 20.4405
R15247 a_50708_569.n28 a_50708_569.t64 20.4405
R15248 a_50708_569.n29 a_50708_569.t73 20.4405
R15249 a_50708_569.n30 a_50708_569.t84 20.4405
R15250 a_50708_569.n31 a_50708_569.t96 20.4405
R15251 a_50708_569.n32 a_50708_569.t83 20.4405
R15252 a_50708_569.n33 a_50708_569.t90 20.4405
R15253 a_50708_569.n34 a_50708_569.t103 20.4405
R15254 a_50708_569.t111 a_50708_569.n35 20.4405
R15255 a_50708_569.t28 a_50708_569.n37 20.4405
R15256 a_50708_569.t108 a_50708_569.n39 20.4405
R15257 a_50708_569.n53 a_50708_569.t113 20.4405
R15258 a_50708_569.n54 a_50708_569.t85 20.4405
R15259 a_50708_569.n61 a_50708_569.t57 20.4405
R15260 a_50708_569.n60 a_50708_569.t112 20.4405
R15261 a_50708_569.n68 a_50708_569.t91 20.4405
R15262 a_50708_569.n69 a_50708_569.t41 20.4405
R15263 a_50708_569.n67 a_50708_569.t98 20.4405
R15264 a_50708_569.n48 a_50708_569.n47 19.2623
R15265 a_50708_569.n55 a_50708_569.n54 19.2623
R15266 a_50708_569.n62 a_50708_569.n61 19.2623
R15267 a_50708_569.n70 a_50708_569.n69 19.2623
R15268 a_50708_569.n47 a_50708_569.n46 17.2497
R15269 a_50708_569.n54 a_50708_569.n53 17.2497
R15270 a_50708_569.n61 a_50708_569.n60 17.2497
R15271 a_50708_569.n69 a_50708_569.n68 17.2497
R15272 a_50708_569.n72 a_50708_569.n66 15.8172
R15273 a_50708_569.n66 a_50708_569.n65 15.8172
R15274 a_50708_569.n57 a_50708_569.n52 15.8172
R15275 a_50708_569.n52 a_50708_569.n51 15.8172
R15276 a_50708_569.n4 a_50708_569.n3 15.8172
R15277 a_50708_569.n5 a_50708_569.n4 15.8172
R15278 a_50708_569.n6 a_50708_569.n5 15.8172
R15279 a_50708_569.n7 a_50708_569.n6 15.8172
R15280 a_50708_569.n8 a_50708_569.n7 15.8172
R15281 a_50708_569.n9 a_50708_569.n8 15.8172
R15282 a_50708_569.n10 a_50708_569.n9 15.8172
R15283 a_50708_569.n11 a_50708_569.n10 15.8172
R15284 a_50708_569.n12 a_50708_569.n11 15.8172
R15285 a_50708_569.n13 a_50708_569.n12 15.8172
R15286 a_50708_569.n25 a_50708_569.n13 15.8172
R15287 a_50708_569.n43 a_50708_569.n25 15.8172
R15288 a_50708_569.n44 a_50708_569.n43 15.8172
R15289 a_50708_569.n45 a_50708_569.n44 15.8172
R15290 a_50708_569.n50 a_50708_569.n45 15.8172
R15291 a_50708_569.n51 a_50708_569.n50 15.8172
R15292 a_50708_569.n58 a_50708_569.n57 15.8172
R15293 a_50708_569.n59 a_50708_569.n58 15.8172
R15294 a_50708_569.n64 a_50708_569.n59 15.8172
R15295 a_50708_569.n65 a_50708_569.n64 15.8172
R15296 a_50708_569.n73 a_50708_569.n72 15.8172
R15297 a_50708_569.n74 a_50708_569.n73 15.8172
R15298 a_50708_569.n71 a_50708_569.n67 15.7165
R15299 a_50708_569.n3 a_50708_569.n2 15.4944
R15300 a_50708_569.n27 a_50708_569.n26 15.3531
R15301 a_50708_569.n28 a_50708_569.n27 15.2373
R15302 a_50708_569.n29 a_50708_569.n28 14.4179
R15303 a_50708_569.n30 a_50708_569.n29 14.4179
R15304 a_50708_569.n31 a_50708_569.n30 14.4179
R15305 a_50708_569.n32 a_50708_569.n31 14.4179
R15306 a_50708_569.n33 a_50708_569.n32 14.4179
R15307 a_50708_569.n34 a_50708_569.n33 14.4179
R15308 a_50708_569.n35 a_50708_569.n34 14.3002
R15309 a_50708_569.n38 a_50708_569.n36 13.3198
R15310 a_50708_569.n40 a_50708_569.n38 13.3198
R15311 a_50708_569.n41 a_50708_569.n40 13.3198
R15312 a_50708_569.n77 a_50708_569.n76 12.7287
R15313 a_50708_569.n78 a_50708_569.n77 12.7287
R15314 a_50708_569.n79 a_50708_569.n78 12.7287
R15315 a_50708_569.n80 a_50708_569.n79 12.7287
R15316 a_50708_569.n81 a_50708_569.n80 12.7287
R15317 a_50708_569.n82 a_50708_569.n81 12.7287
R15318 a_50708_569.n76 a_50708_569.n75 12.6663
R15319 a_50708_569.n83 a_50708_569.n82 4.60781
R15320 a_50708_569.n96 a_50708_569.n95 3.69699
R15321 a_50708_569.n49 a_50708_569.n48 3.54621
R15322 a_50708_569.n56 a_50708_569.n55 3.54621
R15323 a_50708_569.n63 a_50708_569.n62 3.54621
R15324 a_50708_569.n71 a_50708_569.n70 3.54621
R15325 a_50708_569.n100 a_50708_569.n85 3.23924
R15326 a_50708_569.n99 a_50708_569.n87 3.23924
R15327 a_50708_569.n103 a_50708_569.n101 3.23924
R15328 a_50708_569.n83 a_50708_569.n1 3.2392
R15329 a_50708_569.n96 a_50708_569.n93 3.2392
R15330 a_50708_569.n98 a_50708_569.n89 3.23916
R15331 a_50708_569.n97 a_50708_569.n91 3.23916
R15332 a_50708_569.n18 a_50708_569.n15 2.91928
R15333 a_50708_569.n24 a_50708_569.n23 2.58908
R15334 a_50708_569.n21 a_50708_569.n20 2.58711
R15335 a_50708_569.n18 a_50708_569.n17 2.58292
R15336 a_50708_569.n1 a_50708_569.t12 0.6505
R15337 a_50708_569.n1 a_50708_569.n0 0.6505
R15338 a_50708_569.n85 a_50708_569.t16 0.6505
R15339 a_50708_569.n85 a_50708_569.n84 0.6505
R15340 a_50708_569.n87 a_50708_569.t17 0.6505
R15341 a_50708_569.n87 a_50708_569.n86 0.6505
R15342 a_50708_569.n89 a_50708_569.t20 0.6505
R15343 a_50708_569.n89 a_50708_569.n88 0.6505
R15344 a_50708_569.n91 a_50708_569.t21 0.6505
R15345 a_50708_569.n91 a_50708_569.n90 0.6505
R15346 a_50708_569.n93 a_50708_569.t10 0.6505
R15347 a_50708_569.n93 a_50708_569.n92 0.6505
R15348 a_50708_569.n95 a_50708_569.t3 0.6505
R15349 a_50708_569.n95 a_50708_569.n94 0.6505
R15350 a_50708_569.t1 a_50708_569.n103 0.6505
R15351 a_50708_569.n103 a_50708_569.n102 0.6505
R15352 a_50708_569.n23 a_50708_569.t7 0.5855
R15353 a_50708_569.n23 a_50708_569.n22 0.5855
R15354 a_50708_569.n15 a_50708_569.t19 0.5855
R15355 a_50708_569.n15 a_50708_569.n14 0.5855
R15356 a_50708_569.n17 a_50708_569.t5 0.5855
R15357 a_50708_569.n17 a_50708_569.n16 0.5855
R15358 a_50708_569.n20 a_50708_569.t14 0.5855
R15359 a_50708_569.n20 a_50708_569.n19 0.5855
R15360 a_50708_569.n98 a_50708_569.n97 0.466449
R15361 a_50708_569.n101 a_50708_569.n83 0.46531
R15362 a_50708_569.n101 a_50708_569.n100 0.46531
R15363 a_50708_569.n100 a_50708_569.n99 0.46531
R15364 a_50708_569.n97 a_50708_569.n96 0.46531
R15365 a_50708_569.n99 a_50708_569.n98 0.464171
R15366 a_50708_569.n21 a_50708_569.n18 0.341015
R15367 a_50708_569.n24 a_50708_569.n21 0.337297
R15368 OUT.n8 OUT.n7 3.74358
R15369 OUT.n10 OUT.n1 3.24303
R15370 OUT.n9 OUT.n3 3.24286
R15371 OUT.n8 OUT.n5 3.24211
R15372 OUT.n84 OUT.n21 3.23441
R15373 OUT.n81 OUT.n27 3.23441
R15374 OUT.n76 OUT.n39 3.23441
R15375 OUT.n69 OUT.n55 3.23441
R15376 OUT.n68 OUT.n59 3.23441
R15377 OUT.n81 OUT.n29 3.23391
R15378 OUT.n83 OUT.n23 3.23391
R15379 OUT.n76 OUT.n41 3.23387
R15380 OUT.n73 OUT.n47 3.23387
R15381 OUT.n75 OUT.n43 3.23387
R15382 OUT.n78 OUT.n35 3.23387
R15383 OUT.n80 OUT.n31 3.23387
R15384 OUT.n69 OUT.n57 3.23383
R15385 OUT.n67 OUT.n61 3.23383
R15386 OUT.n71 OUT.n51 3.23383
R15387 OUT.n82 OUT.n25 3.23358
R15388 OUT.n66 OUT.n65 3.2335
R15389 OUT.n85 OUT.n19 3.23343
R15390 OUT.n87 OUT.n15 3.23343
R15391 OUT.n86 OUT.n17 3.23337
R15392 OUT.n79 OUT.n33 3.23316
R15393 OUT.n77 OUT.n37 3.23312
R15394 OUT.n74 OUT.n45 3.23312
R15395 OUT.n72 OUT.n49 3.23312
R15396 OUT.n70 OUT.n53 3.23312
R15397 OUT.n66 OUT.n63 3.2315
R15398 OUT.n100 OUT.n97 2.98385
R15399 OUT.n113 OUT.n95 2.87549
R15400 OUT.n116 OUT.n115 2.70972
R15401 OUT.n119 OUT.n118 2.62238
R15402 OUT.n122 OUT.n121 2.62091
R15403 OUT.n125 OUT.n124 2.61945
R15404 OUT.n131 OUT.n130 2.61636
R15405 OUT.n137 OUT.n136 2.61619
R15406 OUT.n128 OUT.n127 2.61619
R15407 OUT.n134 OUT.n133 2.61554
R15408 OUT.n13 OUT.n12 2.6005
R15409 OUT.n91 OUT.n90 2.6005
R15410 OUT.n100 OUT.n99 2.58236
R15411 OUT.n106 OUT.n105 2.58184
R15412 OUT.n109 OUT.n108 2.5817
R15413 OUT.n103 OUT.n102 2.58166
R15414 OUT.n112 OUT.n111 2.58122
R15415 OUT.n138 OUT.n137 1.60202
R15416 OUT.n138 OUT.n93 1.34978
R15417 OUT.n139 OUT.n138 0.888141
R15418 OUT.n13 OUT.n10 0.79069
R15419 OUT.n84 OUT.n83 0.781777
R15420 OUT.n81 OUT.n80 0.781777
R15421 OUT.n76 OUT.n75 0.781777
R15422 OUT.n69 OUT.n68 0.781777
R15423 OUT.n67 OUT.n66 0.781777
R15424 OUT.n82 OUT.n81 0.779862
R15425 OUT.n79 OUT.n78 0.779862
R15426 OUT.n77 OUT.n76 0.779862
R15427 OUT.n74 OUT.n73 0.779862
R15428 OUT.n72 OUT.n71 0.779862
R15429 OUT.n70 OUT.n69 0.779862
R15430 OUT.n88 OUT.n87 0.777947
R15431 OUT.n86 OUT.n85 0.777947
R15432 OUT.n139 OUT.n91 0.655477
R15433 OUT.n90 OUT.t65 0.6505
R15434 OUT.n90 OUT.n89 0.6505
R15435 OUT.n12 OUT.t52 0.6505
R15436 OUT.n12 OUT.n11 0.6505
R15437 OUT.n1 OUT.t58 0.6505
R15438 OUT.n1 OUT.n0 0.6505
R15439 OUT.n3 OUT.t92 0.6505
R15440 OUT.n3 OUT.n2 0.6505
R15441 OUT.n5 OUT.t45 0.6505
R15442 OUT.n5 OUT.n4 0.6505
R15443 OUT.n7 OUT.t62 0.6505
R15444 OUT.n7 OUT.n6 0.6505
R15445 OUT.n17 OUT.t90 0.6505
R15446 OUT.n17 OUT.n16 0.6505
R15447 OUT.n21 OUT.t39 0.6505
R15448 OUT.n21 OUT.n20 0.6505
R15449 OUT.n25 OUT.t54 0.6505
R15450 OUT.n25 OUT.n24 0.6505
R15451 OUT.n29 OUT.t87 0.6505
R15452 OUT.n29 OUT.n28 0.6505
R15453 OUT.n27 OUT.t78 0.6505
R15454 OUT.n27 OUT.n26 0.6505
R15455 OUT.n33 OUT.t91 0.6505
R15456 OUT.n33 OUT.n32 0.6505
R15457 OUT.n37 OUT.t67 0.6505
R15458 OUT.n37 OUT.n36 0.6505
R15459 OUT.n41 OUT.t77 0.6505
R15460 OUT.n41 OUT.n40 0.6505
R15461 OUT.n39 OUT.t66 0.6505
R15462 OUT.n39 OUT.n38 0.6505
R15463 OUT.n45 OUT.t36 0.6505
R15464 OUT.n45 OUT.n44 0.6505
R15465 OUT.n49 OUT.t33 0.6505
R15466 OUT.n49 OUT.n48 0.6505
R15467 OUT.n53 OUT.t50 0.6505
R15468 OUT.n53 OUT.n52 0.6505
R15469 OUT.n57 OUT.t34 0.6505
R15470 OUT.n57 OUT.n56 0.6505
R15471 OUT.n55 OUT.t88 0.6505
R15472 OUT.n55 OUT.n54 0.6505
R15473 OUT.n59 OUT.t38 0.6505
R15474 OUT.n59 OUT.n58 0.6505
R15475 OUT.n65 OUT.t89 0.6505
R15476 OUT.n65 OUT.n64 0.6505
R15477 OUT.n63 OUT.t81 0.6505
R15478 OUT.n63 OUT.n62 0.6505
R15479 OUT.n61 OUT.t51 0.6505
R15480 OUT.n61 OUT.n60 0.6505
R15481 OUT.n51 OUT.t64 0.6505
R15482 OUT.n51 OUT.n50 0.6505
R15483 OUT.n47 OUT.t47 0.6505
R15484 OUT.n47 OUT.n46 0.6505
R15485 OUT.n43 OUT.t48 0.6505
R15486 OUT.n43 OUT.n42 0.6505
R15487 OUT.n35 OUT.t80 0.6505
R15488 OUT.n35 OUT.n34 0.6505
R15489 OUT.n31 OUT.t37 0.6505
R15490 OUT.n31 OUT.n30 0.6505
R15491 OUT.n23 OUT.t68 0.6505
R15492 OUT.n23 OUT.n22 0.6505
R15493 OUT.n19 OUT.t53 0.6505
R15494 OUT.n19 OUT.n18 0.6505
R15495 OUT.n15 OUT.t35 0.6505
R15496 OUT.n15 OUT.n14 0.6505
R15497 OUT.n91 OUT.n88 0.633955
R15498 OUT.n88 OUT.n13 0.631666
R15499 OUT.n127 OUT.t28 0.5855
R15500 OUT.n127 OUT.n126 0.5855
R15501 OUT.n133 OUT.t10 0.5855
R15502 OUT.n133 OUT.n132 0.5855
R15503 OUT.n136 OUT.t31 0.5855
R15504 OUT.n136 OUT.n135 0.5855
R15505 OUT.n115 OUT.t8 0.5855
R15506 OUT.n115 OUT.n114 0.5855
R15507 OUT.n118 OUT.t23 0.5855
R15508 OUT.n118 OUT.n117 0.5855
R15509 OUT.n121 OUT.t16 0.5855
R15510 OUT.n121 OUT.n120 0.5855
R15511 OUT.n124 OUT.t1 0.5855
R15512 OUT.n124 OUT.n123 0.5855
R15513 OUT.n130 OUT.t21 0.5855
R15514 OUT.n130 OUT.n129 0.5855
R15515 OUT.n97 OUT.t18 0.5855
R15516 OUT.n97 OUT.n96 0.5855
R15517 OUT.n99 OUT.t19 0.5855
R15518 OUT.n99 OUT.n98 0.5855
R15519 OUT.n102 OUT.t13 0.5855
R15520 OUT.n102 OUT.n101 0.5855
R15521 OUT.n105 OUT.t14 0.5855
R15522 OUT.n105 OUT.n104 0.5855
R15523 OUT.n108 OUT.t6 0.5855
R15524 OUT.n108 OUT.n107 0.5855
R15525 OUT.n111 OUT.t30 0.5855
R15526 OUT.n111 OUT.n110 0.5855
R15527 OUT.n95 OUT.t0 0.5855
R15528 OUT.n95 OUT.n94 0.5855
R15529 OUT.n93 OUT.t25 0.5855
R15530 OUT.n93 OUT.n92 0.5855
R15531 OUT.n116 OUT.n113 0.510866
R15532 OUT.n10 OUT.n9 0.504747
R15533 OUT.n9 OUT.n8 0.504747
R15534 OUT.n106 OUT.n103 0.403414
R15535 OUT.n109 OUT.n106 0.402304
R15536 OUT.n112 OUT.n109 0.400958
R15537 OUT.n103 OUT.n100 0.400949
R15538 OUT OUT.n139 0.346655
R15539 OUT.n128 OUT.n125 0.334681
R15540 OUT.n131 OUT.n128 0.334473
R15541 OUT.n122 OUT.n119 0.334465
R15542 OUT.n134 OUT.n131 0.334064
R15543 OUT.n137 OUT.n134 0.333663
R15544 OUT.n125 OUT.n122 0.333454
R15545 OUT.n119 OUT.n116 0.244714
R15546 OUT.n113 OUT.n112 0.107492
R15547 OUT.n87 OUT.n86 0.00432979
R15548 OUT.n85 OUT.n84 0.00241489
R15549 OUT.n83 OUT.n82 0.00241489
R15550 OUT.n80 OUT.n79 0.00241489
R15551 OUT.n78 OUT.n77 0.00241489
R15552 OUT.n75 OUT.n74 0.00241489
R15553 OUT.n73 OUT.n72 0.00241489
R15554 OUT.n71 OUT.n70 0.00241489
R15555 OUT.n68 OUT.n67 0.00241489
R15556 S1.n12 S1.t14 45.6363
R15557 S1.n18 S1.t7 29.6446
R15558 S1.t19 S1.n19 29.6446
R15559 S1.n0 S1.t6 24.6117
R15560 S1.n8 S1.t4 23.6945
R15561 S1.t2 S1.n9 23.6945
R15562 S1.n19 S1.n18 22.2047
R15563 S1.t14 S1.t18 22.1925
R15564 S1.n13 S1.n12 20.9314
R15565 S1.n9 S1.n8 18.8035
R15566 S1 S1.t19 18.5175
R15567 S1.n6 S1.n4 15.8172
R15568 S1.n5 S1.n1 15.8172
R15569 S1.n6 S1.n5 15.8172
R15570 S1.n4 S1.t15 14.8925
R15571 S1.t20 S1.n6 14.8925
R15572 S1.n5 S1.t0 14.8925
R15573 S1.n10 S1.n2 12.2457
R15574 S1.n7 S1.n2 12.2457
R15575 S1.n7 S1.n3 12.2457
R15576 S1.n11 S1.t13 11.6285
R15577 S1.n3 S1.t4 8.9065
R15578 S1.t9 S1.n7 8.9065
R15579 S1.t10 S1.n2 8.9065
R15580 S1.n10 S1.t2 8.9065
R15581 S1.n6 S1.t1 8.6145
R15582 S1.n4 S1.t17 8.6145
R15583 S1.n5 S1.t5 8.6145
R15584 S1.n1 S1.t16 8.59715
R15585 S1.t15 S1.n3 8.3225
R15586 S1.n7 S1.t20 8.3225
R15587 S1.t0 S1.n2 8.3225
R15588 S1.t13 S1.n10 8.3225
R15589 S1.n0 S1.t12 6.1325
R15590 S1.n12 S1.t3 6.1325
R15591 S1.n13 S1.t8 6.1325
R15592 S1.n18 S1.t21 6.1325
R15593 S1.n19 S1.t11 6.1325
R15594 S1.n15 S1.n13 4.86736
R15595 S1.n17 S1.n0 4.79907
R15596 S1 S1.n11 4.223
R15597 S1.n8 S1.t9 3.6505
R15598 S1.n9 S1.t10 3.6505
R15599 S1.n11 S1.n1 3.1807
R15600 S1.n15 S1.n14 1.48152
R15601 S1.n14 S1 0.920438
R15602 S1.n14 S1 0.870565
R15603 S1 S1.n17 0.640368
R15604 S1.n16 S1 0.1655
R15605 S1.n16 S1.n15 0.108008
R15606 S1.n17 S1.n16 0.0592755
R15607 A_MUX_1.Tr_Gate_1.CLK.n1 A_MUX_1.Tr_Gate_1.CLK.t12 45.6363
R15608 A_MUX_1.Tr_Gate_1.CLK.n3 A_MUX_1.Tr_Gate_1.CLK.t20 29.6446
R15609 A_MUX_1.Tr_Gate_1.CLK.t15 A_MUX_1.Tr_Gate_1.CLK.n4 29.6446
R15610 A_MUX_1.Tr_Gate_1.CLK.n5 A_MUX_1.Tr_Gate_1.CLK.t16 24.6117
R15611 A_MUX_1.Tr_Gate_1.CLK.n4 A_MUX_1.Tr_Gate_1.CLK.n3 22.2047
R15612 A_MUX_1.Tr_Gate_1.CLK.t12 A_MUX_1.Tr_Gate_1.CLK.t17 22.1925
R15613 A_MUX_1.Tr_Gate_1.CLK.n2 A_MUX_1.Tr_Gate_1.CLK.n1 20.9314
R15614 A_MUX_1.Tr_Gate_1.CLK A_MUX_1.Tr_Gate_1.CLK.t15 18.5245
R15615 A_MUX_1.Tr_Gate_1.CLK.n1 A_MUX_1.Tr_Gate_1.CLK.t19 6.1325
R15616 A_MUX_1.Tr_Gate_1.CLK.n2 A_MUX_1.Tr_Gate_1.CLK.t13 6.1325
R15617 A_MUX_1.Tr_Gate_1.CLK.n3 A_MUX_1.Tr_Gate_1.CLK.t14 6.1325
R15618 A_MUX_1.Tr_Gate_1.CLK.n4 A_MUX_1.Tr_Gate_1.CLK.t21 6.1325
R15619 A_MUX_1.Tr_Gate_1.CLK.n5 A_MUX_1.Tr_Gate_1.CLK.t18 6.1325
R15620 A_MUX_1.Tr_Gate_1.CLK.n0 A_MUX_1.Tr_Gate_1.CLK.n2 5.28481
R15621 A_MUX_1.Tr_Gate_1.CLK.n0 A_MUX_1.Tr_Gate_1.CLK.n5 4.89628
R15622 A_MUX_1.Tr_Gate_1.CLK.n16 A_MUX_1.Tr_Gate_1.CLK.t7 3.6405
R15623 A_MUX_1.Tr_Gate_1.CLK.n16 A_MUX_1.Tr_Gate_1.CLK.n15 3.6405
R15624 A_MUX_1.Tr_Gate_1.CLK.n9 A_MUX_1.Tr_Gate_1.CLK.t5 3.6405
R15625 A_MUX_1.Tr_Gate_1.CLK.n9 A_MUX_1.Tr_Gate_1.CLK.n8 3.6405
R15626 A_MUX_1.Tr_Gate_1.CLK.n11 A_MUX_1.Tr_Gate_1.CLK.t9 3.6405
R15627 A_MUX_1.Tr_Gate_1.CLK.n11 A_MUX_1.Tr_Gate_1.CLK.n10 3.6405
R15628 A_MUX_1.Tr_Gate_1.CLK.n18 A_MUX_1.Tr_Gate_1.CLK.t11 3.6405
R15629 A_MUX_1.Tr_Gate_1.CLK.n18 A_MUX_1.Tr_Gate_1.CLK.n17 3.6405
R15630 A_MUX_1.Tr_Gate_1.CLK.n20 A_MUX_1.Tr_Gate_1.CLK.n14 3.50463
R15631 A_MUX_1.Tr_Gate_1.CLK.n21 A_MUX_1.Tr_Gate_1.CLK.n7 3.50463
R15632 A_MUX_1.Tr_Gate_1.CLK.n14 A_MUX_1.Tr_Gate_1.CLK.t2 3.2765
R15633 A_MUX_1.Tr_Gate_1.CLK.n14 A_MUX_1.Tr_Gate_1.CLK.n13 3.2765
R15634 A_MUX_1.Tr_Gate_1.CLK.n7 A_MUX_1.Tr_Gate_1.CLK.t0 3.2765
R15635 A_MUX_1.Tr_Gate_1.CLK.n7 A_MUX_1.Tr_Gate_1.CLK.n6 3.2765
R15636 A_MUX_1.Tr_Gate_1.CLK.n12 A_MUX_1.Tr_Gate_1.CLK.n11 3.06224
R15637 A_MUX_1.Tr_Gate_1.CLK.n19 A_MUX_1.Tr_Gate_1.CLK.n16 3.06224
R15638 A_MUX_1.Tr_Gate_1.CLK.n12 A_MUX_1.Tr_Gate_1.CLK.n9 2.6005
R15639 A_MUX_1.Tr_Gate_1.CLK.n19 A_MUX_1.Tr_Gate_1.CLK.n18 2.6005
R15640 A_MUX_1.Tr_Gate_1.CLK.n21 A_MUX_1.Tr_Gate_1.CLK.n20 0.798761
R15641 A_MUX_1.Tr_Gate_1.CLK.n0 A_MUX_1.Tr_Gate_1.CLK 0.629601
R15642 A_MUX_1.Tr_Gate_1.CLK A_MUX_1.Tr_Gate_1.CLK.n21 0.562022
R15643 A_MUX_1.Tr_Gate_1.CLK A_MUX_1.Tr_Gate_1.CLK.n0 0.253378
R15644 A_MUX_1.Tr_Gate_1.CLK.n21 A_MUX_1.Tr_Gate_1.CLK.n12 0.18637
R15645 A_MUX_1.Tr_Gate_1.CLK.n20 A_MUX_1.Tr_Gate_1.CLK.n19 0.18637
R15646 a_43528_12082.t0 a_43528_12082.t1 12.9675
R15647 a_43828_11460.t0 a_43828_11460.t1 12.9675
R15648 VCO_DFF_C_0.OUTB.n13 VCO_DFF_C_0.OUTB.t23 37.6513
R15649 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUTB.n13 33.2393
R15650 VCO_DFF_C_0.OUTB.n10 VCO_DFF_C_0.OUTB.t21 32.7094
R15651 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUTB.n12 25.0644
R15652 VCO_DFF_C_0.OUTB.n10 VCO_DFF_C_0.OUTB.t22 23.2875
R15653 VCO_DFF_C_0.OUTB.n11 VCO_DFF_C_0.OUTB.t24 23.2875
R15654 VCO_DFF_C_0.OUTB.n12 VCO_DFF_C_0.OUTB.t20 20.4405
R15655 VCO_DFF_C_0.OUTB.n13 VCO_DFF_C_0.OUTB.t25 20.4405
R15656 VCO_DFF_C_0.OUTB.n11 VCO_DFF_C_0.OUTB.n10 12.5148
R15657 VCO_DFF_C_0.OUTB.n12 VCO_DFF_C_0.OUTB.n11 12.2081
R15658 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUTB.n3 6.65095
R15659 VCO_DFF_C_0.OUTB.n9 VCO_DFF_C_0.OUTB.n6 5.81586
R15660 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUTB.t4 5.10151
R15661 VCO_DFF_C_0.OUTB.n0 VCO_DFF_C_0.OUTB.t5 5.1005
R15662 VCO_DFF_C_0.OUTB.n0 VCO_DFF_C_0.OUTB.t15 5.08021
R15663 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUTB.n5 4.66164
R15664 VCO_DFF_C_0.OUTB.n17 VCO_DFF_C_0.OUTB.t10 3.6405
R15665 VCO_DFF_C_0.OUTB.n17 VCO_DFF_C_0.OUTB.n16 3.6405
R15666 VCO_DFF_C_0.OUTB.n19 VCO_DFF_C_0.OUTB.t0 3.6405
R15667 VCO_DFF_C_0.OUTB.n19 VCO_DFF_C_0.OUTB.n18 3.6405
R15668 VCO_DFF_C_0.OUTB.n23 VCO_DFF_C_0.OUTB.t9 3.6405
R15669 VCO_DFF_C_0.OUTB.n23 VCO_DFF_C_0.OUTB.n22 3.6405
R15670 VCO_DFF_C_0.OUTB.n25 VCO_DFF_C_0.OUTB.t12 3.6405
R15671 VCO_DFF_C_0.OUTB.n25 VCO_DFF_C_0.OUTB.n24 3.6405
R15672 VCO_DFF_C_0.OUTB.n1 VCO_DFF_C_0.OUTB.n15 3.50463
R15673 VCO_DFF_C_0.OUTB.n2 VCO_DFF_C_0.OUTB.n21 3.50463
R15674 VCO_DFF_C_0.OUTB.n15 VCO_DFF_C_0.OUTB.t11 3.2765
R15675 VCO_DFF_C_0.OUTB.n15 VCO_DFF_C_0.OUTB.n14 3.2765
R15676 VCO_DFF_C_0.OUTB.n21 VCO_DFF_C_0.OUTB.t8 3.2765
R15677 VCO_DFF_C_0.OUTB.n21 VCO_DFF_C_0.OUTB.n20 3.2765
R15678 VCO_DFF_C_0.OUTB.n1 VCO_DFF_C_0.OUTB.n19 3.06224
R15679 VCO_DFF_C_0.OUTB.n2 VCO_DFF_C_0.OUTB.n25 3.06224
R15680 VCO_DFF_C_0.OUTB.n9 VCO_DFF_C_0.OUTB.n8 2.85093
R15681 VCO_DFF_C_0.OUTB.n1 VCO_DFF_C_0.OUTB.n17 2.6005
R15682 VCO_DFF_C_0.OUTB.n2 VCO_DFF_C_0.OUTB.n23 2.6005
R15683 VCO_DFF_C_0.OUTB.n8 VCO_DFF_C_0.OUTB.t14 2.16717
R15684 VCO_DFF_C_0.OUTB.n8 VCO_DFF_C_0.OUTB.n7 2.16717
R15685 VCO_DFF_C_0.OUTB.n5 VCO_DFF_C_0.OUTB.t6 1.9505
R15686 VCO_DFF_C_0.OUTB.n5 VCO_DFF_C_0.OUTB.n4 1.9505
R15687 VCO_DFF_C_0.OUTB.n3 VCO_DFF_C_0.OUTB 1.47848
R15688 VCO_DFF_C_0.OUTB.n0 VCO_DFF_C_0.OUTB.n9 1.09092
R15689 VCO_DFF_C_0.OUTB.n1 VCO_DFF_C_0.OUTB.n2 0.98463
R15690 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUTB.n1 0.908615
R15691 VCO_DFF_C_0.OUTB.n3 VCO_DFF_C_0.OUTB 0.883804
R15692 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUTB.n0 0.787647
R15693 a_32467_10269.t8 a_32467_10269.t7 17.9898
R15694 a_32467_10269.t9 a_32467_10269.t8 17.9898
R15695 a_32467_10269.t6 a_32467_10269.t9 17.9898
R15696 a_32467_10269.n0 a_32467_10269.t6 13.0554
R15697 a_32467_10269.n1 a_32467_10269.n3 8.89703
R15698 a_32467_10269.n0 a_32467_10269.n4 8.71168
R15699 a_32467_10269.n7 a_32467_10269.n1 8.60182
R15700 a_32467_10269.n1 a_32467_10269.n6 8.6005
R15701 a_32467_10269.n0 a_32467_10269.n5 8.6005
R15702 a_32467_10269.n1 a_32467_10269.n2 8.5505
R15703 a_32467_10269.n1 a_32467_10269.n0 2.08339
R15704 RES_74k_1.M.t1 RES_74k_1.M.t6 3.92959
R15705 RES_74k_1.M.t1 RES_74k_1.M.n0 3.19141
R15706 RES_74k_1.M.t1 RES_74k_1.M 8.48731
R15707 RES_74k_1.M RES_74k_1.M.t0 6.14618
R15708 RES_74k_1.M.t1 RES_74k_1.M.t7 5.18834
R15709 RES_74k_1.M.t1 RES_74k_1.M.t3 5.18264
R15710 RES_74k_1.M.t1 RES_74k_1.M.t4 3.07204
R15711 RES_74k_1.M.t1 RES_74k_1.M.t5 3.0618
R15712 RES_74k_1.M.t1 RES_74k_1.M.t2 3.0279
R15713 S2.n12 S2.t8 45.6363
R15714 S2.n18 S2.t13 29.6446
R15715 S2.t15 S2.n19 29.6446
R15716 S2.n0 S2.t5 24.6117
R15717 S2.n8 S2.t12 23.6945
R15718 S2.t1 S2.n9 23.6945
R15719 S2.n19 S2.n18 22.2047
R15720 S2.t8 S2.t20 22.1925
R15721 S2.n13 S2.n12 20.9314
R15722 S2.n9 S2.n8 18.8035
R15723 S2 S2.t15 18.5191
R15724 S2.n6 S2.n4 15.8172
R15725 S2.n6 S2.n5 15.8172
R15726 S2.n5 S2.n1 15.8172
R15727 S2.n4 S2.t9 14.8925
R15728 S2.t16 S2.n6 14.8925
R15729 S2.n5 S2.t4 14.8925
R15730 S2.n10 S2.n2 12.2457
R15731 S2.n7 S2.n2 12.2457
R15732 S2.n7 S2.n3 12.2457
R15733 S2.n11 S2.t21 11.6285
R15734 S2.n3 S2.t12 8.9065
R15735 S2.t0 S2.n7 8.9065
R15736 S2.t11 S2.n2 8.9065
R15737 S2.n10 S2.t1 8.9065
R15738 S2.n6 S2.t14 8.6145
R15739 S2.n4 S2.t6 8.6145
R15740 S2.n5 S2.t3 8.6145
R15741 S2.n1 S2.t18 8.59715
R15742 S2.t9 S2.n3 8.3225
R15743 S2.n7 S2.t16 8.3225
R15744 S2.t4 S2.n2 8.3225
R15745 S2.t21 S2.n10 8.3225
R15746 S2.n0 S2.t7 6.1325
R15747 S2.n12 S2.t17 6.1325
R15748 S2.n13 S2.t19 6.1325
R15749 S2.n18 S2.t2 6.1325
R15750 S2.n19 S2.t10 6.1325
R15751 S2.n14 S2 5.70508
R15752 S2.n15 S2.n13 4.8671
R15753 S2.n17 S2.n0 4.79907
R15754 S2 S2.n11 4.223
R15755 S2.n8 S2.t0 3.6505
R15756 S2.n9 S2.t11 3.6505
R15757 S2.n11 S2.n1 3.1807
R15758 S2.n15 S2.n14 1.48741
R15759 S2.n14 S2 0.93932
R15760 S2 S2.n17 0.640368
R15761 S2.n16 S2 0.1655
R15762 S2.n16 S2.n15 0.108287
R15763 S2.n17 S2.n16 0.0592755
R15764 A_MUX_3.Tr_Gate_1.CLK.n17 A_MUX_3.Tr_Gate_1.CLK.t12 45.6363
R15765 A_MUX_3.Tr_Gate_1.CLK.n19 A_MUX_3.Tr_Gate_1.CLK.t15 29.6446
R15766 A_MUX_3.Tr_Gate_1.CLK.t17 A_MUX_3.Tr_Gate_1.CLK.n20 29.6446
R15767 A_MUX_3.Tr_Gate_1.CLK.n21 A_MUX_3.Tr_Gate_1.CLK.t13 24.6117
R15768 A_MUX_3.Tr_Gate_1.CLK.n20 A_MUX_3.Tr_Gate_1.CLK.n19 22.2047
R15769 A_MUX_3.Tr_Gate_1.CLK.t12 A_MUX_3.Tr_Gate_1.CLK.t19 22.1925
R15770 A_MUX_3.Tr_Gate_1.CLK.n18 A_MUX_3.Tr_Gate_1.CLK.n17 20.9314
R15771 A_MUX_3.Tr_Gate_1.CLK A_MUX_3.Tr_Gate_1.CLK.t17 18.524
R15772 A_MUX_3.Tr_Gate_1.CLK.n21 A_MUX_3.Tr_Gate_1.CLK.t16 6.1325
R15773 A_MUX_3.Tr_Gate_1.CLK.n19 A_MUX_3.Tr_Gate_1.CLK.t20 6.1325
R15774 A_MUX_3.Tr_Gate_1.CLK.n20 A_MUX_3.Tr_Gate_1.CLK.t14 6.1325
R15775 A_MUX_3.Tr_Gate_1.CLK.n17 A_MUX_3.Tr_Gate_1.CLK.t18 6.1325
R15776 A_MUX_3.Tr_Gate_1.CLK.n18 A_MUX_3.Tr_Gate_1.CLK.t21 6.1325
R15777 A_MUX_3.Tr_Gate_1.CLK.n0 A_MUX_3.Tr_Gate_1.CLK.n18 5.28289
R15778 A_MUX_3.Tr_Gate_1.CLK.n0 A_MUX_3.Tr_Gate_1.CLK.n21 4.89628
R15779 A_MUX_3.Tr_Gate_1.CLK.n12 A_MUX_3.Tr_Gate_1.CLK.t5 3.6405
R15780 A_MUX_3.Tr_Gate_1.CLK.n12 A_MUX_3.Tr_Gate_1.CLK.n11 3.6405
R15781 A_MUX_3.Tr_Gate_1.CLK.n6 A_MUX_3.Tr_Gate_1.CLK.t4 3.6405
R15782 A_MUX_3.Tr_Gate_1.CLK.n6 A_MUX_3.Tr_Gate_1.CLK.n5 3.6405
R15783 A_MUX_3.Tr_Gate_1.CLK.n8 A_MUX_3.Tr_Gate_1.CLK.t10 3.6405
R15784 A_MUX_3.Tr_Gate_1.CLK.n8 A_MUX_3.Tr_Gate_1.CLK.n7 3.6405
R15785 A_MUX_3.Tr_Gate_1.CLK.n14 A_MUX_3.Tr_Gate_1.CLK.t11 3.6405
R15786 A_MUX_3.Tr_Gate_1.CLK.n14 A_MUX_3.Tr_Gate_1.CLK.n13 3.6405
R15787 A_MUX_3.Tr_Gate_1.CLK.n16 A_MUX_3.Tr_Gate_1.CLK.n2 3.50463
R15788 A_MUX_3.Tr_Gate_1.CLK.n10 A_MUX_3.Tr_Gate_1.CLK.n4 3.50463
R15789 A_MUX_3.Tr_Gate_1.CLK.n2 A_MUX_3.Tr_Gate_1.CLK.t1 3.2765
R15790 A_MUX_3.Tr_Gate_1.CLK.n2 A_MUX_3.Tr_Gate_1.CLK.n1 3.2765
R15791 A_MUX_3.Tr_Gate_1.CLK.n4 A_MUX_3.Tr_Gate_1.CLK.t0 3.2765
R15792 A_MUX_3.Tr_Gate_1.CLK.n4 A_MUX_3.Tr_Gate_1.CLK.n3 3.2765
R15793 A_MUX_3.Tr_Gate_1.CLK.n9 A_MUX_3.Tr_Gate_1.CLK.n8 3.06224
R15794 A_MUX_3.Tr_Gate_1.CLK.n15 A_MUX_3.Tr_Gate_1.CLK.n14 3.06224
R15795 A_MUX_3.Tr_Gate_1.CLK.n9 A_MUX_3.Tr_Gate_1.CLK.n6 2.6005
R15796 A_MUX_3.Tr_Gate_1.CLK.n15 A_MUX_3.Tr_Gate_1.CLK.n12 2.6005
R15797 A_MUX_3.Tr_Gate_1.CLK.n16 A_MUX_3.Tr_Gate_1.CLK.n10 0.798761
R15798 A_MUX_3.Tr_Gate_1.CLK.n0 A_MUX_3.Tr_Gate_1.CLK 0.629597
R15799 A_MUX_3.Tr_Gate_1.CLK A_MUX_3.Tr_Gate_1.CLK.n16 0.562022
R15800 A_MUX_3.Tr_Gate_1.CLK A_MUX_3.Tr_Gate_1.CLK.n0 0.253378
R15801 A_MUX_3.Tr_Gate_1.CLK.n10 A_MUX_3.Tr_Gate_1.CLK.n9 0.18637
R15802 A_MUX_3.Tr_Gate_1.CLK.n16 A_MUX_3.Tr_Gate_1.CLK.n15 0.18637
R15803 a_25557_8739.n0 a_25557_8739.t3 24.1084
R15804 a_25557_8739.n1 a_25557_8739.t5 12.5565
R15805 a_25557_8739.n0 a_25557_8739.t4 8.6145
R15806 a_25557_8739.n2 a_25557_8739.t0 6.71215
R15807 a_25557_8739.n2 a_25557_8739.n1 4.46748
R15808 a_25557_8739.n3 a_25557_8739.t1 3.6405
R15809 a_25557_8739.n4 a_25557_8739.n3 3.6405
R15810 a_25557_8739.n3 a_25557_8739.n2 2.83724
R15811 a_25557_8739.n1 a_25557_8739.n0 1.8985
R15812 a_34443_2598.n69 a_34443_2598.n51 9.67588
R15813 a_34443_2598.n4 a_34443_2598.n89 3.7286
R15814 a_34443_2598.n15 a_34443_2598.n14 3.71799
R15815 a_34443_2598.n2 a_34443_2598.n59 3.71473
R15816 a_34443_2598.n1 a_34443_2598.n75 3.70973
R15817 a_34443_2598.n87 a_34443_2598.t34 3.2765
R15818 a_34443_2598.n87 a_34443_2598.n86 3.2765
R15819 a_34443_2598.n12 a_34443_2598.t17 3.2765
R15820 a_34443_2598.n12 a_34443_2598.n11 3.2765
R15821 a_34443_2598.n9 a_34443_2598.t39 3.2765
R15822 a_34443_2598.n9 a_34443_2598.n8 3.2765
R15823 a_34443_2598.n7 a_34443_2598.t31 3.2765
R15824 a_34443_2598.n7 a_34443_2598.n6 3.2765
R15825 a_34443_2598.n66 a_34443_2598.t19 3.2765
R15826 a_34443_2598.n66 a_34443_2598.n65 3.2765
R15827 a_34443_2598.n53 a_34443_2598.t23 3.2765
R15828 a_34443_2598.n53 a_34443_2598.n52 3.2765
R15829 a_34443_2598.n55 a_34443_2598.t35 3.2765
R15830 a_34443_2598.n55 a_34443_2598.n54 3.2765
R15831 a_34443_2598.n80 a_34443_2598.t49 3.2765
R15832 a_34443_2598.n80 a_34443_2598.n79 3.2765
R15833 a_34443_2598.n71 a_34443_2598.t43 3.2765
R15834 a_34443_2598.n71 a_34443_2598.n70 3.2765
R15835 a_34443_2598.n18 a_34443_2598.t52 3.2765
R15836 a_34443_2598.n18 a_34443_2598.n17 3.2765
R15837 a_34443_2598.n20 a_34443_2598.t9 3.2765
R15838 a_34443_2598.n20 a_34443_2598.n19 3.2765
R15839 a_34443_2598.n26 a_34443_2598.t1 3.2765
R15840 a_34443_2598.n26 a_34443_2598.n25 3.2765
R15841 a_34443_2598.n22 a_34443_2598.t53 3.2765
R15842 a_34443_2598.n22 a_34443_2598.n21 3.2765
R15843 a_34443_2598.n24 a_34443_2598.t57 3.2765
R15844 a_34443_2598.n24 a_34443_2598.n23 3.2765
R15845 a_34443_2598.n39 a_34443_2598.t6 3.2765
R15846 a_34443_2598.n39 a_34443_2598.n38 3.2765
R15847 a_34443_2598.n41 a_34443_2598.t10 3.2765
R15848 a_34443_2598.n41 a_34443_2598.n40 3.2765
R15849 a_34443_2598.n43 a_34443_2598.t0 3.2765
R15850 a_34443_2598.n43 a_34443_2598.n42 3.2765
R15851 a_34443_2598.n35 a_34443_2598.t7 3.2765
R15852 a_34443_2598.n35 a_34443_2598.n34 3.2765
R15853 a_34443_2598.n37 a_34443_2598.t54 3.2765
R15854 a_34443_2598.n37 a_34443_2598.n36 3.2765
R15855 a_34443_2598.n84 a_34443_2598.t12 3.2765
R15856 a_34443_2598.n84 a_34443_2598.n83 3.2765
R15857 a_34443_2598.n73 a_34443_2598.t15 3.2765
R15858 a_34443_2598.n73 a_34443_2598.n72 3.2765
R15859 a_34443_2598.n77 a_34443_2598.t41 3.2765
R15860 a_34443_2598.n77 a_34443_2598.n76 3.2765
R15861 a_34443_2598.n75 a_34443_2598.t47 3.2765
R15862 a_34443_2598.n75 a_34443_2598.n74 3.2765
R15863 a_34443_2598.n57 a_34443_2598.t44 3.2765
R15864 a_34443_2598.n57 a_34443_2598.n56 3.2765
R15865 a_34443_2598.n61 a_34443_2598.t21 3.2765
R15866 a_34443_2598.n61 a_34443_2598.n60 3.2765
R15867 a_34443_2598.n59 a_34443_2598.t33 3.2765
R15868 a_34443_2598.n59 a_34443_2598.n58 3.2765
R15869 a_34443_2598.n14 a_34443_2598.t29 3.2765
R15870 a_34443_2598.n14 a_34443_2598.n13 3.2765
R15871 a_34443_2598.n91 a_34443_2598.t11 3.2765
R15872 a_34443_2598.n91 a_34443_2598.n90 3.2765
R15873 a_34443_2598.n89 a_34443_2598.t22 3.2765
R15874 a_34443_2598.n89 a_34443_2598.n88 3.2765
R15875 a_34443_2598.n93 a_34443_2598.t24 3.2765
R15876 a_34443_2598.n94 a_34443_2598.n93 3.2765
R15877 a_34443_2598.n49 a_34443_2598.n37 3.1505
R15878 a_34443_2598.n50 a_34443_2598.n35 3.1505
R15879 a_34443_2598.n44 a_34443_2598.n43 3.1505
R15880 a_34443_2598.n46 a_34443_2598.n41 3.1505
R15881 a_34443_2598.n47 a_34443_2598.n39 3.1505
R15882 a_34443_2598.n29 a_34443_2598.n24 3.1505
R15883 a_34443_2598.n30 a_34443_2598.n22 3.1505
R15884 a_34443_2598.n27 a_34443_2598.n26 3.1505
R15885 a_34443_2598.n32 a_34443_2598.n20 3.1505
R15886 a_34443_2598.n33 a_34443_2598.n18 3.1505
R15887 a_34443_2598.n85 a_34443_2598.n84 3.1505
R15888 a_34443_2598.n81 a_34443_2598.n71 3.1505
R15889 a_34443_2598.n78 a_34443_2598.n73 3.1505
R15890 a_34443_2598.n62 a_34443_2598.n57 3.1505
R15891 a_34443_2598.n64 a_34443_2598.n53 3.1505
R15892 a_34443_2598.n67 a_34443_2598.n66 3.1505
R15893 a_34443_2598.n10 a_34443_2598.n9 3.1505
R15894 a_34443_2598.n92 a_34443_2598.n87 3.1505
R15895 a_34443_2598.n4 a_34443_2598.n91 1.84747
R15896 a_34443_2598.n2 a_34443_2598.n61 1.84743
R15897 a_34443_2598.n1 a_34443_2598.n77 1.84737
R15898 a_34443_2598.n0 a_34443_2598.n80 1.84737
R15899 a_34443_2598.n63 a_34443_2598.n55 1.84737
R15900 a_34443_2598.n5 a_34443_2598.n7 1.84732
R15901 a_34443_2598.n93 a_34443_2598.n3 1.84728
R15902 a_34443_2598.n16 a_34443_2598.n12 1.84618
R15903 a_34443_2598.n85 a_34443_2598.n82 0.899822
R15904 a_34443_2598.n68 a_34443_2598.n67 0.899822
R15905 a_34443_2598.n47 a_34443_2598.n46 0.758798
R15906 a_34443_2598.n30 a_34443_2598.n29 0.758798
R15907 a_34443_2598.n51 a_34443_2598.n50 0.724996
R15908 a_34443_2598.n50 a_34443_2598.n49 0.7205
R15909 a_34443_2598.n33 a_34443_2598.n32 0.7205
R15910 a_34443_2598.n51 a_34443_2598.n33 0.636952
R15911 a_34443_2598.n16 a_34443_2598.n10 0.622339
R15912 a_34443_2598.n64 a_34443_2598.n63 0.607482
R15913 a_34443_2598.n81 a_34443_2598.n0 0.604163
R15914 a_34443_2598.n3 a_34443_2598.n85 0.602337
R15915 a_34443_2598.n63 a_34443_2598.n62 0.595434
R15916 a_34443_2598.n45 a_34443_2598.n44 0.555819
R15917 a_34443_2598.n28 a_34443_2598.n27 0.555819
R15918 a_34443_2598.n49 a_34443_2598.n48 0.551989
R15919 a_34443_2598.n32 a_34443_2598.n31 0.551989
R15920 a_34443_2598.n69 a_34443_2598.n68 0.378745
R15921 a_34443_2598.n48 a_34443_2598.n47 0.283904
R15922 a_34443_2598.n31 a_34443_2598.n30 0.283904
R15923 a_34443_2598.n46 a_34443_2598.n45 0.280074
R15924 a_34443_2598.n29 a_34443_2598.n28 0.280074
R15925 a_34443_2598.n82 a_34443_2598.n69 0.248582
R15926 a_34443_2598.n82 a_34443_2598.n81 0.247022
R15927 a_34443_2598.n68 a_34443_2598.n64 0.247022
R15928 a_34443_2598.n16 a_34443_2598.n15 0.0460206
R15929 a_34443_2598.n5 a_34443_2598.n3 3.58925
R15930 a_34443_2598.n78 a_34443_2598.n1 0.627536
R15931 a_34443_2598.n62 a_34443_2598.n2 0.622521
R15932 a_34443_2598.n92 a_34443_2598.n4 0.619689
R15933 a_34443_2598.n10 a_34443_2598.n5 0.609769
R15934 a_34443_2598.n3 a_34443_2598.n92 0.602476
R15935 a_34443_2598.n0 a_34443_2598.n78 0.598753
R15936 RES_74k_1.P.n89 RES_74k_1.P.t68 6.77746
R15937 RES_74k_1.P.n161 RES_74k_1.P.t24 6.1905
R15938 RES_74k_1.P.n114 RES_74k_1.P.t23 6.1905
R15939 RES_74k_1.P.n113 RES_74k_1.P.t48 6.1905
R15940 RES_74k_1.P.n112 RES_74k_1.P.t47 6.1905
R15941 RES_74k_1.P.n111 RES_74k_1.P.t74 6.1905
R15942 RES_74k_1.P.n110 RES_74k_1.P.t73 6.1905
R15943 RES_74k_1.P.n109 RES_74k_1.P.t22 6.1905
R15944 RES_74k_1.P.n108 RES_74k_1.P.t21 6.1905
R15945 RES_74k_1.P.n107 RES_74k_1.P.t56 6.1905
R15946 RES_74k_1.P.n106 RES_74k_1.P.t55 6.1905
R15947 RES_74k_1.P.n104 RES_74k_1.P.t44 6.1905
R15948 RES_74k_1.P.n89 RES_74k_1.P.t94 6.1905
R15949 RES_74k_1.P.n90 RES_74k_1.P.t84 6.1905
R15950 RES_74k_1.P.n91 RES_74k_1.P.t70 6.1905
R15951 RES_74k_1.P.n92 RES_74k_1.P.t96 6.1905
R15952 RES_74k_1.P.n93 RES_74k_1.P.t52 6.1905
R15953 RES_74k_1.P.n94 RES_74k_1.P.t12 6.1905
R15954 RES_74k_1.P.n95 RES_74k_1.P.t72 6.1905
R15955 RES_74k_1.P.n96 RES_74k_1.P.t60 6.1905
R15956 RES_74k_1.P.n97 RES_74k_1.P.t8 6.1905
R15957 RES_74k_1.P.n98 RES_74k_1.P.t42 6.1905
R15958 RES_74k_1.P.n99 RES_74k_1.P.t18 6.1905
R15959 RES_74k_1.P.n100 RES_74k_1.P.t92 6.1905
R15960 RES_74k_1.P.n101 RES_74k_1.P.t36 6.1905
R15961 RES_74k_1.P.n102 RES_74k_1.P.t78 6.1905
R15962 RES_74k_1.P.n103 RES_74k_1.P.t38 6.1905
R15963 RES_74k_1.P.n134 RES_74k_1.P.t29 6.1905
R15964 RES_74k_1.P.n135 RES_74k_1.P.t30 6.1905
R15965 RES_74k_1.P.n136 RES_74k_1.P.t5 6.1905
R15966 RES_74k_1.P.n137 RES_74k_1.P.t6 6.1905
R15967 RES_74k_1.P.n138 RES_74k_1.P.t65 6.1905
R15968 RES_74k_1.P.n139 RES_74k_1.P.t66 6.1905
R15969 RES_74k_1.P.n140 RES_74k_1.P.t15 6.1905
R15970 RES_74k_1.P.n141 RES_74k_1.P.t16 6.1905
R15971 RES_74k_1.P.n142 RES_74k_1.P.t39 6.1905
R15972 RES_74k_1.P.n132 RES_74k_1.P.t40 6.1905
R15973 RES_74k_1.P.n131 RES_74k_1.P.t58 6.1905
R15974 RES_74k_1.P.n130 RES_74k_1.P.t62 6.1905
R15975 RES_74k_1.P.n129 RES_74k_1.P.t46 6.1905
R15976 RES_74k_1.P.n128 RES_74k_1.P.t32 6.1905
R15977 RES_74k_1.P.n127 RES_74k_1.P.t80 6.1905
R15978 RES_74k_1.P.n126 RES_74k_1.P.t10 6.1905
R15979 RES_74k_1.P.n125 RES_74k_1.P.t50 6.1905
R15980 RES_74k_1.P.n124 RES_74k_1.P.t64 6.1905
R15981 RES_74k_1.P.n123 RES_74k_1.P.t14 6.1905
R15982 RES_74k_1.P.n122 RES_74k_1.P.t1 6.1905
R15983 RES_74k_1.P.n121 RES_74k_1.P.t76 6.1905
R15984 RES_74k_1.P.n120 RES_74k_1.P.t89 6.1905
R15985 RES_74k_1.P.n119 RES_74k_1.P.t20 6.1905
R15986 RES_74k_1.P.n118 RES_74k_1.P.t82 6.1905
R15987 RES_74k_1.P.n117 RES_74k_1.P.t34 6.1905
R15988 RES_74k_1.P.n116 RES_74k_1.P.t86 6.1905
R15989 RES_74k_1.P.n115 RES_74k_1.P.t3 6.1905
R15990 RES_74k_1.P.n158 RES_74k_1.P.t57 6.1905
R15991 RES_74k_1.P.n133 RES_74k_1.P.t2 6.1905
R15992 RES_74k_1.P.n143 RES_74k_1.P.t85 6.1905
R15993 RES_74k_1.P.n144 RES_74k_1.P.t33 6.1905
R15994 RES_74k_1.P.n145 RES_74k_1.P.t81 6.1905
R15995 RES_74k_1.P.n146 RES_74k_1.P.t19 6.1905
R15996 RES_74k_1.P.n147 RES_74k_1.P.t88 6.1905
R15997 RES_74k_1.P.n148 RES_74k_1.P.t75 6.1905
R15998 RES_74k_1.P.n149 RES_74k_1.P.t0 6.1905
R15999 RES_74k_1.P.n150 RES_74k_1.P.t13 6.1905
R16000 RES_74k_1.P.n151 RES_74k_1.P.t63 6.1905
R16001 RES_74k_1.P.n152 RES_74k_1.P.t49 6.1905
R16002 RES_74k_1.P.n153 RES_74k_1.P.t9 6.1905
R16003 RES_74k_1.P.n154 RES_74k_1.P.t79 6.1905
R16004 RES_74k_1.P.n155 RES_74k_1.P.t31 6.1905
R16005 RES_74k_1.P.n156 RES_74k_1.P.t45 6.1905
R16006 RES_74k_1.P.n157 RES_74k_1.P.t61 6.1905
R16007 RES_74k_1.P.n72 RES_74k_1.P.t67 6.1905
R16008 RES_74k_1.P.n73 RES_74k_1.P.t93 6.1905
R16009 RES_74k_1.P.n74 RES_74k_1.P.t83 6.1905
R16010 RES_74k_1.P.n75 RES_74k_1.P.t69 6.1905
R16011 RES_74k_1.P.n76 RES_74k_1.P.t95 6.1905
R16012 RES_74k_1.P.n77 RES_74k_1.P.t51 6.1905
R16013 RES_74k_1.P.n78 RES_74k_1.P.t11 6.1905
R16014 RES_74k_1.P.n79 RES_74k_1.P.t71 6.1905
R16015 RES_74k_1.P.n80 RES_74k_1.P.t59 6.1905
R16016 RES_74k_1.P.n81 RES_74k_1.P.t7 6.1905
R16017 RES_74k_1.P.n82 RES_74k_1.P.t41 6.1905
R16018 RES_74k_1.P.n83 RES_74k_1.P.t17 6.1905
R16019 RES_74k_1.P.n84 RES_74k_1.P.t91 6.1905
R16020 RES_74k_1.P.n85 RES_74k_1.P.t35 6.1905
R16021 RES_74k_1.P.n86 RES_74k_1.P.t77 6.1905
R16022 RES_74k_1.P.n87 RES_74k_1.P.t37 6.1905
R16023 RES_74k_1.P.n88 RES_74k_1.P.t43 6.1905
R16024 RES_74k_1.P.n286 RES_74k_1.P.t26 5.81586
R16025 RES_74k_1.P.n278 RES_74k_1.P.n277 5.48458
R16026 RES_74k_1.P.n282 RES_74k_1.P.n279 5.10151
R16027 RES_74k_1.P.n289 RES_74k_1.P.n288 5.10119
R16028 RES_74k_1.P.n287 RES_74k_1.P.n283 5.08021
R16029 RES_74k_1.P.n282 RES_74k_1.P.n281 4.66164
R16030 RES_74k_1.P.n239 RES_74k_1.P.n70 4.5266
R16031 RES_74k_1.P.n62 RES_74k_1.P.n183 4.5266
R16032 RES_74k_1.P.n64 RES_74k_1.P.n173 4.5266
R16033 RES_74k_1.P.n248 RES_74k_1.P.n246 4.5266
R16034 RES_74k_1.P.n210 RES_74k_1.P.n208 4.5266
R16035 RES_74k_1.P.n263 RES_74k_1.P.n170 4.5266
R16036 RES_74k_1.P.n237 RES_74k_1.P.n236 4.52639
R16037 RES_74k_1.P.n217 RES_74k_1.P.n63 4.52502
R16038 RES_74k_1.P.n258 RES_74k_1.P.n66 4.52502
R16039 RES_74k_1.P.n245 RES_74k_1.P.n244 4.52502
R16040 RES_74k_1.P.n207 RES_74k_1.P.n206 4.52502
R16041 RES_74k_1.P.n235 RES_74k_1.P.n171 4.52502
R16042 RES_74k_1.P.n236 RES_74k_1.P.n44 4.5032
R16043 RES_74k_1.P.n42 RES_74k_1.P.n63 4.5032
R16044 RES_74k_1.P.n67 RES_74k_1.P.n66 4.5032
R16045 RES_74k_1.P.n244 RES_74k_1.P.n68 4.5032
R16046 RES_74k_1.P.n206 RES_74k_1.P.n42 4.5032
R16047 RES_74k_1.P.n44 RES_74k_1.P.n235 4.5032
R16048 RES_74k_1.P.n204 RES_74k_1.P.n203 4.50309
R16049 RES_74k_1.P.n26 RES_74k_1.P.n55 2.25075
R16050 RES_74k_1.P.n28 RES_74k_1.P.n30 0.375824
R16051 RES_74k_1.P.n2 RES_74k_1.P.n0 0.207027
R16052 RES_74k_1.P.n24 RES_74k_1.P.n20 0.375425
R16053 RES_74k_1.P.n240 RES_74k_1.P.n239 4.5005
R16054 RES_74k_1.P.n269 RES_74k_1.P.n168 4.5005
R16055 RES_74k_1.P.n35 RES_74k_1.P.n51 0.749789
R16056 RES_74k_1.P.n31 RES_74k_1.P.n54 0.00898642
R16057 RES_74k_1.P.n270 RES_74k_1.P.n268 4.5005
R16058 RES_74k_1.P.n31 RES_74k_1.P.n32 0.372209
R16059 RES_74k_1.P.n28 RES_74k_1.P.n271 4.5005
R16060 RES_74k_1.P.n32 RES_74k_1.P.n50 0.0116877
R16061 RES_74k_1.P.n35 RES_74k_1.P.n58 2.2508
R16062 RES_74k_1.P.n267 RES_74k_1.P.n28 4.5005
R16063 RES_74k_1.P.n216 RES_74k_1.P.n183 4.5005
R16064 RES_74k_1.P.n22 RES_74k_1.P.n16 2.25095
R16065 RES_74k_1.P.n21 RES_74k_1.P.n19 2.25095
R16066 RES_74k_1.P.n201 RES_74k_1.P.n200 4.5005
R16067 RES_74k_1.P.n225 RES_74k_1.P.n224 4.5005
R16068 RES_74k_1.P.n20 RES_74k_1.P.n232 4.5005
R16069 RES_74k_1.P.n18 RES_74k_1.P.n20 4.5005
R16070 RES_74k_1.P.n9 RES_74k_1.P.n178 4.5005
R16071 RES_74k_1.P.n180 RES_74k_1.P.n177 4.5005
R16072 RES_74k_1.P.n14 RES_74k_1.P.n39 0.374407
R16073 RES_74k_1.P.n203 RES_74k_1.P.n202 4.5005
R16074 RES_74k_1.P.n37 RES_74k_1.P.n226 4.5005
R16075 RES_74k_1.P.n231 RES_74k_1.P.n230 4.5005
R16076 RES_74k_1.P.n38 RES_74k_1.P.n176 4.5005
R16077 RES_74k_1.P.n19 RES_74k_1.P.n13 0.00735821
R16078 RES_74k_1.P.n257 RES_74k_1.P.n173 4.5005
R16079 RES_74k_1.P.n249 RES_74k_1.P.n248 4.5005
R16080 RES_74k_1.P.n211 RES_74k_1.P.n210 4.5005
R16081 RES_74k_1.P.n8 RES_74k_1.P.n17 0.749855
R16082 RES_74k_1.P.n190 RES_74k_1.P.n187 4.5005
R16083 RES_74k_1.P.n33 RES_74k_1.P.n52 0.749839
R16084 RES_74k_1.P.n194 RES_74k_1.P.n193 4.5005
R16085 RES_74k_1.P.n3 RES_74k_1.P.n0 0.200279
R16086 RES_74k_1.P.n3 RES_74k_1.P.n33 0.0124268
R16087 RES_74k_1.P.n192 RES_74k_1.P.n0 4.5005
R16088 RES_74k_1.P.n0 RES_74k_1.P.n4 4.5005
R16089 RES_74k_1.P.n12 RES_74k_1.P.n10 0.00311493
R16090 RES_74k_1.P.n27 RES_74k_1.P.n26 1.49652
R16091 RES_74k_1.P.n41 RES_74k_1.P.n6 2.2508
R16092 RES_74k_1.P.n49 RES_74k_1.P.n6 2.25095
R16093 RES_74k_1.P.n26 RES_74k_1.P.n48 4.5005
R16094 RES_74k_1.P.n15 RES_74k_1.P.n21 0.0070381
R16095 RES_74k_1.P.n255 RES_74k_1.P.n233 4.5005
R16096 RES_74k_1.P.n242 RES_74k_1.P.n47 0.00851207
R16097 RES_74k_1.P.n44 RES_74k_1.P.n47 0.896327
R16098 RES_74k_1.P.n47 RES_74k_1.P.n70 4.53411
R16099 RES_74k_1.P.n242 RES_74k_1.P.n241 4.5005
R16100 RES_74k_1.P.n255 RES_74k_1.P.n65 0.0123754
R16101 RES_74k_1.P.n255 RES_74k_1.P.n174 4.5005
R16102 RES_74k_1.P.n255 RES_74k_1.P.n254 4.5005
R16103 RES_74k_1.P.n15 RES_74k_1.P.n26 0.450037
R16104 RES_74k_1.P.n43 RES_74k_1.P.n42 0.896327
R16105 RES_74k_1.P.n214 RES_74k_1.P.n184 4.5005
R16106 RES_74k_1.P.n214 RES_74k_1.P.n43 0.00851207
R16107 RES_74k_1.P.n213 RES_74k_1.P.n46 0.00851207
R16108 RES_74k_1.P.n213 RES_74k_1.P.n205 4.5005
R16109 RES_74k_1.P.n42 RES_74k_1.P.n46 0.896327
R16110 RES_74k_1.P.n252 RES_74k_1.P.n251 4.5005
R16111 RES_74k_1.P.n69 RES_74k_1.P.n68 1.49475
R16112 RES_74k_1.P.n252 RES_74k_1.P.n243 4.5005
R16113 RES_74k_1.P.n253 RES_74k_1.P.n252 4.5005
R16114 RES_74k_1.P.n45 RES_74k_1.P.n266 0.00851206
R16115 RES_74k_1.P.n45 RES_74k_1.P.n44 0.896327
R16116 RES_74k_1.P.n266 RES_74k_1.P.n265 4.5005
R16117 RES_74k_1.P.n264 RES_74k_1.P.n263 4.5005
R16118 RES_74k_1.P.n162 RES_74k_1.P.t90 3.49604
R16119 RES_74k_1.P.n286 RES_74k_1.P.n285 2.85093
R16120 RES_74k_1.P.n277 RES_74k_1.P.n162 2.63074
R16121 RES_74k_1.P.n163 RES_74k_1.P.t97 2.38861
R16122 RES_74k_1.P.n25 RES_74k_1.P.t98 2.38861
R16123 RES_74k_1.P.n40 RES_74k_1.P.t101 2.38861
R16124 RES_74k_1.P.n167 RES_74k_1.P.n166 2.37146
R16125 RES_74k_1.P.n53 RES_74k_1.P.n60 1.15033
R16126 RES_74k_1.P.n247 RES_74k_1.P.n172 2.29119
R16127 RES_74k_1.P.n209 RES_74k_1.P.n182 2.29119
R16128 RES_74k_1.P.n262 RES_74k_1.P.n261 2.28464
R16129 RES_74k_1.P.n166 RES_74k_1.P.n164 2.2505
R16130 RES_74k_1.P.n260 RES_74k_1.P.n259 2.2505
R16131 RES_74k_1.P.n229 RES_74k_1.P.n228 2.2505
R16132 RES_74k_1.P.n227 RES_74k_1.P.n175 2.2505
R16133 RES_74k_1.P.n222 RES_74k_1.P.n221 2.2505
R16134 RES_74k_1.P.n39 RES_74k_1.P.n57 1.12595
R16135 RES_74k_1.P.n220 RES_74k_1.P.n181 2.2505
R16136 RES_74k_1.P.n219 RES_74k_1.P.n218 2.2505
R16137 RES_74k_1.P.n197 RES_74k_1.P.n7 2.2505
R16138 RES_74k_1.P.n199 RES_74k_1.P.n198 2.2505
R16139 RES_74k_1.P.n186 RES_74k_1.P.n185 2.2505
R16140 RES_74k_1.P.n196 RES_74k_1.P.n195 2.2505
R16141 RES_74k_1.P.n163 RES_74k_1.P.t102 2.2505
R16142 RES_74k_1.P.n25 RES_74k_1.P.t100 2.2505
R16143 RES_74k_1.P.n40 RES_74k_1.P.t99 2.2505
R16144 RES_74k_1.P.n238 RES_74k_1.P.n165 2.2505
R16145 RES_74k_1.P.n276 RES_74k_1.P.n275 2.2505
R16146 RES_74k_1.P.n274 RES_74k_1.P.n273 2.2505
R16147 RES_74k_1.P RES_74k_1.P.n60 6.01043
R16148 RES_74k_1.P.n67 RES_74k_1.P.n65 1.49475
R16149 RES_74k_1.P.n69 RES_74k_1.P.n246 4.52828
R16150 RES_74k_1.P.n285 RES_74k_1.P.t25 2.16717
R16151 RES_74k_1.P.n285 RES_74k_1.P.n284 2.16717
R16152 RES_74k_1.P.n281 RES_74k_1.P.t54 1.9505
R16153 RES_74k_1.P.n281 RES_74k_1.P.n280 1.9505
R16154 RES_74k_1.P RES_74k_1.P.n278 1.70663
R16155 RES_74k_1.P.n61 RES_74k_1.P.n54 0.457025
R16156 RES_74k_1.P.n240 RES_74k_1.P.n234 1.5005
R16157 RES_74k_1.P.n216 RES_74k_1.P.n215 1.5005
R16158 RES_74k_1.P.n257 RES_74k_1.P.n256 1.5005
R16159 RES_74k_1.P.n250 RES_74k_1.P.n249 1.5005
R16160 RES_74k_1.P.n212 RES_74k_1.P.n211 1.5005
R16161 RES_74k_1.P.n6 RES_74k_1.P.n50 0.449693
R16162 RES_74k_1.P.n12 RES_74k_1.P.n26 0.562674
R16163 RES_74k_1.P.n264 RES_74k_1.P.n169 1.5005
R16164 RES_74k_1.P.n159 RES_74k_1.P.n131 1.2155
R16165 RES_74k_1.P.n105 RES_74k_1.P.n88 1.2155
R16166 RES_74k_1.P.n132 RES_74k_1.P.n142 1.20532
R16167 RES_74k_1.P.n141 RES_74k_1.P.n140 1.20532
R16168 RES_74k_1.P.n139 RES_74k_1.P.n138 1.20532
R16169 RES_74k_1.P.n137 RES_74k_1.P.n136 1.20532
R16170 RES_74k_1.P.n135 RES_74k_1.P.n134 1.20532
R16171 RES_74k_1.P.n107 RES_74k_1.P.n106 1.20532
R16172 RES_74k_1.P.n109 RES_74k_1.P.n108 1.20532
R16173 RES_74k_1.P.n111 RES_74k_1.P.n110 1.20532
R16174 RES_74k_1.P.n113 RES_74k_1.P.n112 1.20532
R16175 RES_74k_1.P.n160 RES_74k_1.P.n114 1.19574
R16176 RES_74k_1.P.n188 RES_74k_1.P.n185 1.15852
R16177 RES_74k_1.P.n36 RES_74k_1.P.n35 0.750079
R16178 RES_74k_1.P.n272 RES_74k_1.P.n167 1.1255
R16179 RES_74k_1.P.n223 RES_74k_1.P.n222 1.1255
R16180 RES_74k_1.P.n229 RES_74k_1.P.n56 1.1255
R16181 RES_74k_1.P.n181 RES_74k_1.P.n179 1.1255
R16182 RES_74k_1.P.n14 RES_74k_1.P.n13 0.00253734
R16183 RES_74k_1.P.n199 RES_74k_1.P.n17 0.00274448
R16184 RES_74k_1.P.n8 RES_74k_1.P.n5 0.00573346
R16185 RES_74k_1.P.n34 RES_74k_1.P.n33 0.750129
R16186 RES_74k_1.P.n191 RES_74k_1.P.n189 1.1255
R16187 RES_74k_1.P.n52 RES_74k_1.P.n186 0.00277662
R16188 RES_74k_1.P.n10 RES_74k_1.P.n11 0.562854
R16189 RES_74k_1.P.n29 RES_74k_1.P.n28 0.45057
R16190 RES_74k_1.P.n0 RES_74k_1.P.n1 0.450717
R16191 RES_74k_1.P.n11 RES_74k_1.P.n179 0.00229276
R16192 RES_74k_1.P.n16 RES_74k_1.P.n13 0.562901
R16193 RES_74k_1.P.n20 RES_74k_1.P.n23 0.450246
R16194 RES_74k_1.P.n49 RES_74k_1.P.n61 0.00977392
R16195 RES_74k_1.P.n61 RES_74k_1.P.n71 0.452583
R16196 RES_74k_1.P.n51 RES_74k_1.P.n276 0.00286644
R16197 RES_74k_1.P.n238 RES_74k_1.P.n237 1.12295
R16198 RES_74k_1.P.n218 RES_74k_1.P.n217 1.12277
R16199 RES_74k_1.P.n259 RES_74k_1.P.n258 1.12277
R16200 RES_74k_1.P.n247 RES_74k_1.P.n245 1.12277
R16201 RES_74k_1.P.n209 RES_74k_1.P.n207 1.12277
R16202 RES_74k_1.P.n262 RES_74k_1.P.n171 1.12277
R16203 RES_74k_1.P.n197 RES_74k_1.P.n182 1.09572
R16204 RES_74k_1.P.n227 RES_74k_1.P.n172 0.963384
R16205 RES_74k_1.P.n278 RES_74k_1.P 0.922754
R16206 RES_74k_1.P.n220 RES_74k_1.P.n219 0.888704
R16207 RES_74k_1.P.n54 RES_74k_1.P.n53 0.374364
R16208 RES_74k_1.P.n277 RES_74k_1.P 0.717341
R16209 RES_74k_1.P.n287 RES_74k_1.P.n286 0.644196
R16210 RES_74k_1.P.n131 RES_74k_1.P.n130 0.587457
R16211 RES_74k_1.P.n130 RES_74k_1.P.n129 0.587457
R16212 RES_74k_1.P.n129 RES_74k_1.P.n128 0.587457
R16213 RES_74k_1.P.n128 RES_74k_1.P.n127 0.587457
R16214 RES_74k_1.P.n127 RES_74k_1.P.n126 0.587457
R16215 RES_74k_1.P.n126 RES_74k_1.P.n125 0.587457
R16216 RES_74k_1.P.n125 RES_74k_1.P.n124 0.587457
R16217 RES_74k_1.P.n124 RES_74k_1.P.n123 0.587457
R16218 RES_74k_1.P.n123 RES_74k_1.P.n122 0.587457
R16219 RES_74k_1.P.n122 RES_74k_1.P.n121 0.587457
R16220 RES_74k_1.P.n121 RES_74k_1.P.n120 0.587457
R16221 RES_74k_1.P.n120 RES_74k_1.P.n119 0.587457
R16222 RES_74k_1.P.n119 RES_74k_1.P.n118 0.587457
R16223 RES_74k_1.P.n118 RES_74k_1.P.n117 0.587457
R16224 RES_74k_1.P.n117 RES_74k_1.P.n116 0.587457
R16225 RES_74k_1.P.n116 RES_74k_1.P.n115 0.587457
R16226 RES_74k_1.P.n158 RES_74k_1.P.n157 0.587457
R16227 RES_74k_1.P.n157 RES_74k_1.P.n156 0.587457
R16228 RES_74k_1.P.n156 RES_74k_1.P.n155 0.587457
R16229 RES_74k_1.P.n155 RES_74k_1.P.n154 0.587457
R16230 RES_74k_1.P.n154 RES_74k_1.P.n153 0.587457
R16231 RES_74k_1.P.n153 RES_74k_1.P.n152 0.587457
R16232 RES_74k_1.P.n152 RES_74k_1.P.n151 0.587457
R16233 RES_74k_1.P.n151 RES_74k_1.P.n150 0.587457
R16234 RES_74k_1.P.n150 RES_74k_1.P.n149 0.587457
R16235 RES_74k_1.P.n149 RES_74k_1.P.n148 0.587457
R16236 RES_74k_1.P.n148 RES_74k_1.P.n147 0.587457
R16237 RES_74k_1.P.n147 RES_74k_1.P.n146 0.587457
R16238 RES_74k_1.P.n146 RES_74k_1.P.n145 0.587457
R16239 RES_74k_1.P.n145 RES_74k_1.P.n144 0.587457
R16240 RES_74k_1.P.n144 RES_74k_1.P.n143 0.587457
R16241 RES_74k_1.P.n143 RES_74k_1.P.n133 0.587457
R16242 RES_74k_1.P.n88 RES_74k_1.P.n87 0.587457
R16243 RES_74k_1.P.n87 RES_74k_1.P.n86 0.587457
R16244 RES_74k_1.P.n86 RES_74k_1.P.n85 0.587457
R16245 RES_74k_1.P.n85 RES_74k_1.P.n84 0.587457
R16246 RES_74k_1.P.n84 RES_74k_1.P.n83 0.587457
R16247 RES_74k_1.P.n83 RES_74k_1.P.n82 0.587457
R16248 RES_74k_1.P.n82 RES_74k_1.P.n81 0.587457
R16249 RES_74k_1.P.n81 RES_74k_1.P.n80 0.587457
R16250 RES_74k_1.P.n80 RES_74k_1.P.n79 0.587457
R16251 RES_74k_1.P.n79 RES_74k_1.P.n78 0.587457
R16252 RES_74k_1.P.n78 RES_74k_1.P.n77 0.587457
R16253 RES_74k_1.P.n77 RES_74k_1.P.n76 0.587457
R16254 RES_74k_1.P.n76 RES_74k_1.P.n75 0.587457
R16255 RES_74k_1.P.n75 RES_74k_1.P.n74 0.587457
R16256 RES_74k_1.P.n74 RES_74k_1.P.n73 0.587457
R16257 RES_74k_1.P.n73 RES_74k_1.P.n72 0.587457
R16258 RES_74k_1.P.n104 RES_74k_1.P.n103 0.587457
R16259 RES_74k_1.P.n103 RES_74k_1.P.n102 0.587457
R16260 RES_74k_1.P.n102 RES_74k_1.P.n101 0.587457
R16261 RES_74k_1.P.n101 RES_74k_1.P.n100 0.587457
R16262 RES_74k_1.P.n100 RES_74k_1.P.n99 0.587457
R16263 RES_74k_1.P.n99 RES_74k_1.P.n98 0.587457
R16264 RES_74k_1.P.n98 RES_74k_1.P.n97 0.587457
R16265 RES_74k_1.P.n97 RES_74k_1.P.n96 0.587457
R16266 RES_74k_1.P.n96 RES_74k_1.P.n95 0.587457
R16267 RES_74k_1.P.n95 RES_74k_1.P.n94 0.587457
R16268 RES_74k_1.P.n94 RES_74k_1.P.n93 0.587457
R16269 RES_74k_1.P.n93 RES_74k_1.P.n92 0.587457
R16270 RES_74k_1.P.n92 RES_74k_1.P.n91 0.587457
R16271 RES_74k_1.P.n91 RES_74k_1.P.n90 0.587457
R16272 RES_74k_1.P.n90 RES_74k_1.P.n89 0.587457
R16273 RES_74k_1.P.n162 RES_74k_1.P.n161 0.54333
R16274 RES_74k_1.P.n289 RES_74k_1.P.n287 0.4508
R16275 RES_74k_1.P.n261 RES_74k_1.P.n260 0.402623
R16276 RES_74k_1.P.n42 RES_74k_1.P.n2 0.353245
R16277 RES_74k_1.P.n290 RES_74k_1.P.n282 0.309543
R16278 RES_74k_1.P.n290 RES_74k_1.P.n289 0.274999
R16279 RES_74k_1.P.n142 RES_74k_1.P.n141 0.274015
R16280 RES_74k_1.P.n140 RES_74k_1.P.n139 0.274015
R16281 RES_74k_1.P.n138 RES_74k_1.P.n137 0.274015
R16282 RES_74k_1.P.n136 RES_74k_1.P.n135 0.274015
R16283 RES_74k_1.P.n108 RES_74k_1.P.n107 0.274015
R16284 RES_74k_1.P.n110 RES_74k_1.P.n109 0.274015
R16285 RES_74k_1.P.n112 RES_74k_1.P.n111 0.274015
R16286 RES_74k_1.P.n114 RES_74k_1.P.n113 0.274015
R16287 RES_74k_1.P.n133 RES_74k_1.P.n132 0.268344
R16288 RES_74k_1.P.n106 RES_74k_1.P.n105 0.264431
R16289 RES_74k_1.P.n160 RES_74k_1.P.n159 0.254848
R16290 RES_74k_1.P.n253 RES_74k_1.P.n44 0.190884
R16291 RES_74k_1.P.n274 RES_74k_1.P.n165 0.143146
R16292 RES_74k_1.P.n26 RES_74k_1.P.n25 0.0995566
R16293 RES_74k_1.P RES_74k_1.P.n290 0.0936034
R16294 RES_74k_1.P.n2 RES_74k_1.P.n40 0.0946742
R16295 RES_74k_1.P.n71 RES_74k_1.P.n163 0.0692209
R16296 RES_74k_1.P.n198 RES_74k_1.P.n196 0.0366935
R16297 RES_74k_1.P.n221 RES_74k_1.P.n57 0.0355442
R16298 RES_74k_1.P.n236 RES_74k_1.P.n234 0.032
R16299 RES_74k_1.P.n215 RES_74k_1.P.n63 0.032
R16300 RES_74k_1.P.n256 RES_74k_1.P.n66 0.032
R16301 RES_74k_1.P.n250 RES_74k_1.P.n244 0.032
R16302 RES_74k_1.P.n212 RES_74k_1.P.n206 0.032
R16303 RES_74k_1.P.n235 RES_74k_1.P.n169 0.032
R16304 RES_74k_1.P.n159 RES_74k_1.P.n158 0.0298478
R16305 RES_74k_1.P.n105 RES_74k_1.P.n104 0.0298478
R16306 RES_74k_1.P.n161 RES_74k_1.P.n160 0.0298478
R16307 RES_74k_1.P.n241 RES_74k_1.P.n70 0.0257
R16308 RES_74k_1.P.n62 RES_74k_1.P.n184 0.0257
R16309 RES_74k_1.P.n64 RES_74k_1.P.n174 0.0257
R16310 RES_74k_1.P.n246 RES_74k_1.P.n243 0.0257
R16311 RES_74k_1.P.n208 RES_74k_1.P.n205 0.0257
R16312 RES_74k_1.P.n265 RES_74k_1.P.n170 0.0257
R16313 RES_74k_1.P.n39 RES_74k_1.P.n37 0.0241947
R16314 RES_74k_1.P.n3 RES_74k_1.P.n8 0.0143144
R16315 RES_74k_1.P.n225 RES_74k_1.P.n22 0.0230022
R16316 RES_74k_1.P.n51 RES_74k_1.P.n270 0.0266526
R16317 RES_74k_1.P.n19 RES_74k_1.P.n18 0.0204137
R16318 RES_74k_1.P.n271 RES_74k_1.P.n35 0.0197576
R16319 RES_74k_1.P.n275 RES_74k_1.P.n274 0.0197233
R16320 RES_74k_1.P.n32 RES_74k_1.P.n49 0.0169518
R16321 RES_74k_1.P.n60 RES_74k_1.P.n59 0.0100942
R16322 RES_74k_1.P.n43 RES_74k_1.P.n62 4.53411
R16323 RES_74k_1.P.n65 RES_74k_1.P.n64 4.52828
R16324 RES_74k_1.P.n228 RES_74k_1.P.n57 0.0331549
R16325 RES_74k_1.P.n252 RES_74k_1.P.n69 0.0123754
R16326 RES_74k_1.P.n46 RES_74k_1.P.n208 4.53411
R16327 RES_74k_1.P.n45 RES_74k_1.P.n170 4.53411
R16328 RES_74k_1.P.n240 RES_74k_1.P.n237 0.00898995
R16329 RES_74k_1.P.n217 RES_74k_1.P.n216 0.00836872
R16330 RES_74k_1.P.n258 RES_74k_1.P.n257 0.00836872
R16331 RES_74k_1.P.n249 RES_74k_1.P.n245 0.00836872
R16332 RES_74k_1.P.n211 RES_74k_1.P.n207 0.00836872
R16333 RES_74k_1.P.n264 RES_74k_1.P.n171 0.00836872
R16334 RES_74k_1.P.n58 RES_74k_1.P.n50 0.0114122
R16335 RES_74k_1.P.n260 RES_74k_1.P.n172 0.00567241
R16336 RES_74k_1.P.n219 RES_74k_1.P.n182 0.00563308
R16337 RES_74k_1.P.n164 RES_74k_1.P.n36 0.0033494
R16338 RES_74k_1.P.n195 RES_74k_1.P.n34 0.00325857
R16339 RES_74k_1.P.n5 RES_74k_1.P.n7 0.748386
R16340 RES_74k_1.P.n10 RES_74k_1.P.n9 0.0044823
R16341 RES_74k_1.P.n189 RES_74k_1.P.n187 0.00437097
R16342 RES_74k_1.P.n191 RES_74k_1.P.n190 0.00437097
R16343 RES_74k_1.P.n23 RES_74k_1.P.n56 0.00422129
R16344 RES_74k_1.P.n200 RES_74k_1.P.n12 0.00744789
R16345 RES_74k_1.P.n230 RES_74k_1.P.n38 0.00428319
R16346 RES_74k_1.P.n229 RES_74k_1.P.n175 0.00428319
R16347 RES_74k_1.P.n228 RES_74k_1.P.n227 0.00428319
R16348 RES_74k_1.P.n166 RES_74k_1.P.n59 0.0041
R16349 RES_74k_1.P.n269 RES_74k_1.P.n167 0.00384061
R16350 RES_74k_1.P.n272 RES_74k_1.P.n168 0.00384061
R16351 RES_74k_1.P.n261 RES_74k_1.P.n165 0.0037767
R16352 RES_74k_1.P.n223 RES_74k_1.P.n180 0.00368584
R16353 RES_74k_1.P.n222 RES_74k_1.P.n177 0.00368584
R16354 RES_74k_1.P.n202 RES_74k_1.P.n179 0.00348673
R16355 RES_74k_1.P.n175 RES_74k_1.P.n23 0.754339
R16356 RES_74k_1.P.n203 RES_74k_1.P.n181 0.00348673
R16357 RES_74k_1.P.n232 RES_74k_1.P.n176 0.00328761
R16358 RES_74k_1.P.n223 RES_74k_1.P.n11 0.00229276
R16359 RES_74k_1.P.n222 RES_74k_1.P.n181 0.0030885
R16360 RES_74k_1.P.n37 RES_74k_1.P.n177 0.0030885
R16361 RES_74k_1.P.n221 RES_74k_1.P.n220 0.0030885
R16362 RES_74k_1.P.n251 RES_74k_1.P.n67 0.00305754
R16363 RES_74k_1.P.n254 RES_74k_1.P.n68 0.00305754
R16364 RES_74k_1.P.n273 RES_74k_1.P.n167 0.00285808
R16365 RES_74k_1.P.n270 RES_74k_1.P.n269 0.00285808
R16366 RES_74k_1.P.n29 RES_74k_1.P.n272 0.0034252
R16367 RES_74k_1.P.n224 RES_74k_1.P.n48 0.00249115
R16368 RES_74k_1.P.n233 RES_74k_1.P.n24 0.291506
R16369 RES_74k_1.P.n226 RES_74k_1.P.n178 0.00229204
R16370 RES_74k_1.P.n231 RES_74k_1.P.n56 0.00229204
R16371 RES_74k_1.P.n204 RES_74k_1.P.n55 4.50289
R16372 RES_74k_1.P.n230 RES_74k_1.P.n229 0.00229204
R16373 RES_74k_1.P.n194 RES_74k_1.P.n187 0.00224194
R16374 RES_74k_1.P.n191 RES_74k_1.P.n1 0.0030813
R16375 RES_74k_1.P.n204 RES_74k_1.P.n201 0.00209292
R16376 RES_74k_1.P.n268 RES_74k_1.P.n267 0.00207205
R16377 RES_74k_1.P.n29 RES_74k_1.P.n273 0.753891
R16378 RES_74k_1.P.n189 RES_74k_1.P.n188 0.00187029
R16379 RES_74k_1.P.n198 RES_74k_1.P.n197 0.00185484
R16380 RES_74k_1.P.n17 RES_74k_1.P.n34 0.0356736
R16381 RES_74k_1.P.n199 RES_74k_1.P.n7 0.00185484
R16382 RES_74k_1.P.n68 RES_74k_1.P.n67 0.00172762
R16383 RES_74k_1.P.n30 RES_74k_1.P.n6 0.024988
R16384 RES_74k_1.P.n196 RES_74k_1.P.n185 0.00166129
R16385 RES_74k_1.P.n52 RES_74k_1.P.n194 0.027118
R16386 RES_74k_1.P.n195 RES_74k_1.P.n186 0.00166129
R16387 RES_74k_1.P.n251 RES_74k_1.P.n233 0.00162532
R16388 RES_74k_1.P.n254 RES_74k_1.P.n253 0.00162532
R16389 RES_74k_1.P.n202 RES_74k_1.P.n201 0.00149557
R16390 RES_74k_1.P.n18 RES_74k_1.P.n176 0.00149557
R16391 RES_74k_1.P.n232 RES_74k_1.P.n231 0.00149557
R16392 RES_74k_1.P.n275 RES_74k_1.P.n59 0.00148301
R16393 RES_74k_1.P.n193 RES_74k_1.P.n4 0.00146774
R16394 RES_74k_1.P.n239 RES_74k_1.P.n238 0.0014
R16395 RES_74k_1.P.n241 RES_74k_1.P.n240 0.0014
R16396 RES_74k_1.P.n242 RES_74k_1.P.n234 0.0014
R16397 RES_74k_1.P.n215 RES_74k_1.P.n214 0.0014
R16398 RES_74k_1.P.n216 RES_74k_1.P.n184 0.0014
R16399 RES_74k_1.P.n218 RES_74k_1.P.n183 0.0014
R16400 RES_74k_1.P.n256 RES_74k_1.P.n255 0.0014
R16401 RES_74k_1.P.n257 RES_74k_1.P.n174 0.0014
R16402 RES_74k_1.P.n259 RES_74k_1.P.n173 0.0014
R16403 RES_74k_1.P.n252 RES_74k_1.P.n250 0.0014
R16404 RES_74k_1.P.n249 RES_74k_1.P.n243 0.0014
R16405 RES_74k_1.P.n248 RES_74k_1.P.n247 0.0014
R16406 RES_74k_1.P.n213 RES_74k_1.P.n212 0.0014
R16407 RES_74k_1.P.n211 RES_74k_1.P.n205 0.0014
R16408 RES_74k_1.P.n210 RES_74k_1.P.n209 0.0014
R16409 RES_74k_1.P.n266 RES_74k_1.P.n169 0.0014
R16410 RES_74k_1.P.n265 RES_74k_1.P.n264 0.0014
R16411 RES_74k_1.P.n263 RES_74k_1.P.n262 0.0014
R16412 RES_74k_1.P.n180 RES_74k_1.P.n178 0.00129646
R16413 RES_74k_1.P.n226 RES_74k_1.P.n225 0.00129646
R16414 RES_74k_1.P.n22 RES_74k_1.P.n14 0.0106918
R16415 RES_74k_1.P.n200 RES_74k_1.P.n55 0.00269222
R16416 RES_74k_1.P.n276 RES_74k_1.P.n164 0.00128603
R16417 RES_74k_1.P.n267 RES_74k_1.P.n168 0.00128603
R16418 RES_74k_1.P.n271 RES_74k_1.P.n268 0.00128603
R16419 RES_74k_1.P.n58 RES_74k_1.P.n41 0.00228596
R16420 RES_74k_1.P.n1 RES_74k_1.P.n188 0.755076
R16421 RES_74k_1.P.n190 RES_74k_1.P.n4 0.00127419
R16422 RES_74k_1.P.n193 RES_74k_1.P.n192 0.00127419
R16423 RES_74k_1.P.n42 RES_74k_1.P.n26 0.273134
R16424 RES_74k_1.P.n30 RES_74k_1.P.n44 0.140772
R16425 RES_74k_1.P.n24 RES_74k_1.P.n26 0.0443926
R16426 RES_74k_1.P.n21 RES_74k_1.P.n20 0.0387411
R16427 RES_74k_1.P.n35 RES_74k_1.P.n31 0.0378189
R16428 RES_74k_1.P.n41 RES_74k_1.P.n28 0.0371921
R16429 RES_74k_1.P.n192 RES_74k_1.P.n33 0.0351768
R16430 RES_74k_1.P.n39 RES_74k_1.P.n38 0.0341549
R16431 RES_74k_1.P.n53 RES_74k_1.P.n36 0.0338509
R16432 RES_74k_1.P.n9 RES_74k_1.P.n48 0.00109734
R16433 RES_74k_1.P.n224 RES_74k_1.P.n27 0.0156248
R16434 RES_74k_1.P.n71 RES_74k_1.P.n6 0.0133785
R16435 RES_74k_1.P.n16 RES_74k_1.P.n15 0.0122767
R16436 RES_74k_1.P.n27 RES_74k_1.P.n16 0.00921204
R16437 RES_74k_1.P.n5 RES_74k_1.P.n0 2.26254
R16438 A_MUX_0.Tr_Gate_1.CLK.n2 A_MUX_0.Tr_Gate_1.CLK.t21 45.6363
R16439 A_MUX_0.Tr_Gate_1.CLK.n4 A_MUX_0.Tr_Gate_1.CLK.t13 29.6446
R16440 A_MUX_0.Tr_Gate_1.CLK.t17 A_MUX_0.Tr_Gate_1.CLK.n5 29.6446
R16441 A_MUX_0.Tr_Gate_1.CLK.n6 A_MUX_0.Tr_Gate_1.CLK.t15 24.6117
R16442 A_MUX_0.Tr_Gate_1.CLK.n5 A_MUX_0.Tr_Gate_1.CLK.n4 22.2047
R16443 A_MUX_0.Tr_Gate_1.CLK.t21 A_MUX_0.Tr_Gate_1.CLK.t16 22.1925
R16444 A_MUX_0.Tr_Gate_1.CLK.n3 A_MUX_0.Tr_Gate_1.CLK.n2 20.9314
R16445 A_MUX_0.Tr_Gate_1.CLK A_MUX_0.Tr_Gate_1.CLK.t17 18.5231
R16446 A_MUX_0.Tr_Gate_1.CLK.n6 A_MUX_0.Tr_Gate_1.CLK.t18 6.1325
R16447 A_MUX_0.Tr_Gate_1.CLK.n4 A_MUX_0.Tr_Gate_1.CLK.t19 6.1325
R16448 A_MUX_0.Tr_Gate_1.CLK.n5 A_MUX_0.Tr_Gate_1.CLK.t14 6.1325
R16449 A_MUX_0.Tr_Gate_1.CLK.n2 A_MUX_0.Tr_Gate_1.CLK.t20 6.1325
R16450 A_MUX_0.Tr_Gate_1.CLK.n3 A_MUX_0.Tr_Gate_1.CLK.t12 6.1325
R16451 A_MUX_0.Tr_Gate_1.CLK A_MUX_0.Tr_Gate_1.CLK.n3 5.28481
R16452 A_MUX_0.Tr_Gate_1.CLK A_MUX_0.Tr_Gate_1.CLK.n6 4.89628
R16453 A_MUX_0.Tr_Gate_1.CLK.n16 A_MUX_0.Tr_Gate_1.CLK.t7 3.6405
R16454 A_MUX_0.Tr_Gate_1.CLK.n16 A_MUX_0.Tr_Gate_1.CLK.n15 3.6405
R16455 A_MUX_0.Tr_Gate_1.CLK.n12 A_MUX_0.Tr_Gate_1.CLK.t5 3.6405
R16456 A_MUX_0.Tr_Gate_1.CLK.n12 A_MUX_0.Tr_Gate_1.CLK.n11 3.6405
R16457 A_MUX_0.Tr_Gate_1.CLK.n10 A_MUX_0.Tr_Gate_1.CLK.t4 3.6405
R16458 A_MUX_0.Tr_Gate_1.CLK.n10 A_MUX_0.Tr_Gate_1.CLK.n9 3.6405
R16459 A_MUX_0.Tr_Gate_1.CLK.n18 A_MUX_0.Tr_Gate_1.CLK.t0 3.6405
R16460 A_MUX_0.Tr_Gate_1.CLK.n18 A_MUX_0.Tr_Gate_1.CLK.n17 3.6405
R16461 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK.n8 3.50463
R16462 A_MUX_0.Tr_Gate_1.CLK.n0 A_MUX_0.Tr_Gate_1.CLK.n14 3.50463
R16463 A_MUX_0.Tr_Gate_1.CLK.n8 A_MUX_0.Tr_Gate_1.CLK.t1 3.2765
R16464 A_MUX_0.Tr_Gate_1.CLK.n8 A_MUX_0.Tr_Gate_1.CLK.n7 3.2765
R16465 A_MUX_0.Tr_Gate_1.CLK.n14 A_MUX_0.Tr_Gate_1.CLK.t6 3.2765
R16466 A_MUX_0.Tr_Gate_1.CLK.n14 A_MUX_0.Tr_Gate_1.CLK.n13 3.2765
R16467 A_MUX_0.Tr_Gate_1.CLK.n0 A_MUX_0.Tr_Gate_1.CLK.n10 3.06224
R16468 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK.n16 3.06224
R16469 A_MUX_0.Tr_Gate_1.CLK.n0 A_MUX_0.Tr_Gate_1.CLK.n12 2.6005
R16470 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK.n18 2.6005
R16471 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK 1.44401
R16472 A_MUX_0.Tr_Gate_1.CLK.n1 A_MUX_0.Tr_Gate_1.CLK.n0 1.1705
R16473 VCO_DFF_C_0.VCTRL.n4 VCO_DFF_C_0.VCTRL.t20 27.5268
R16474 VCO_DFF_C_0.VCTRL.n17 VCO_DFF_C_0.VCTRL.t17 27.5268
R16475 VCO_DFF_C_0.VCTRL.n19 VCO_DFF_C_0.VCTRL.t24 25.3421
R16476 VCO_DFF_C_0.VCTRL.n7 VCO_DFF_C_0.VCTRL.t32 25.3421
R16477 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCTRL.n16 9.02002
R16478 VCO_DFF_C_0.VCTRL.n21 VCO_DFF_C_0.VCTRL.t34 8.86359
R16479 VCO_DFF_C_0.VCTRL.n9 VCO_DFF_C_0.VCTRL.t21 8.86319
R16480 VCO_DFF_C_0.VCTRL.n30 VCO_DFF_C_0.VCTRL 8.38187
R16481 VCO_DFF_C_0.VCTRL.n11 VCO_DFF_C_0.VCTRL.t31 7.92693
R16482 VCO_DFF_C_0.VCTRL.n24 VCO_DFF_C_0.VCTRL.t28 7.92677
R16483 VCO_DFF_C_0.VCTRL.n8 VCO_DFF_C_0.VCTRL.t16 7.79605
R16484 VCO_DFF_C_0.VCTRL.n22 VCO_DFF_C_0.VCTRL.t19 7.79604
R16485 VCO_DFF_C_0.VCTRL.n5 VCO_DFF_C_0.VCTRL.t30 7.57548
R16486 VCO_DFF_C_0.VCTRL.n18 VCO_DFF_C_0.VCTRL.t26 7.54055
R16487 VCO_DFF_C_0.VCTRL.n6 VCO_DFF_C_0.VCTRL.t27 7.49426
R16488 VCO_DFF_C_0.VCTRL.n23 VCO_DFF_C_0.VCTRL.t29 7.49403
R16489 VCO_DFF_C_0.VCTRL.n0 VCO_DFF_C_0.VCTRL.t15 6.74387
R16490 VCO_DFF_C_0.VCTRL.n1 VCO_DFF_C_0.VCTRL.n48 6.74326
R16491 VCO_DFF_C_0.VCTRL.n12 VCO_DFF_C_0.VCTRL.t23 6.73304
R16492 VCO_DFF_C_0.VCTRL.n25 VCO_DFF_C_0.VCTRL.t18 6.73175
R16493 VCO_DFF_C_0.VCTRL.n1 VCO_DFF_C_0.VCTRL.n49 5.1005
R16494 VCO_DFF_C_0.VCTRL.n0 VCO_DFF_C_0.VCTRL.t12 5.1005
R16495 VCO_DFF_C_0.VCTRL.n5 VCO_DFF_C_0.VCTRL.n4 4.72106
R16496 VCO_DFF_C_0.VCTRL.n18 VCO_DFF_C_0.VCTRL.n17 4.72106
R16497 VCO_DFF_C_0.VCTRL.n10 VCO_DFF_C_0.VCTRL.n7 3.90288
R16498 VCO_DFF_C_0.VCTRL.n20 VCO_DFF_C_0.VCTRL.n19 3.90053
R16499 VCO_DFF_C_0.VCTRL.n46 VCO_DFF_C_0.VCTRL.n43 3.57508
R16500 VCO_DFF_C_0.VCTRL.n34 VCO_DFF_C_0.VCTRL.n37 3.56654
R16501 VCO_DFF_C_0.VCTRL.n1 VCO_DFF_C_0.VCTRL.t0 3.40075
R16502 VCO_DFF_C_0.VCTRL.n0 VCO_DFF_C_0.VCTRL.n38 3.40011
R16503 VCO_DFF_C_0.VCTRL.n39 VCO_DFF_C_0.VCTRL.t14 3.00158
R16504 VCO_DFF_C_0.VCTRL.n50 VCO_DFF_C_0.VCTRL.n47 3.00032
R16505 VCO_DFF_C_0.VCTRL.n15 VCO_DFF_C_0.VCTRL 2.50091
R16506 VCO_DFF_C_0.VCTRL.n28 VCO_DFF_C_0.VCTRL 2.46425
R16507 VCO_DFF_C_0.VCTRL.n35 VCO_DFF_C_0.VCTRL.n33 2.41287
R16508 VCO_DFF_C_0.VCTRL.n52 VCO_DFF_C_0.VCTRL.n41 2.36206
R16509 VCO_DFF_C_0.VCTRL.n16 VCO_DFF_C_0.VCTRL 2.32969
R16510 VCO_DFF_C_0.VCTRL.n41 VCO_DFF_C_0.VCTRL.n40 2.30849
R16511 VCO_DFF_C_0.VCTRL.n3 VCO_DFF_C_0.VCTRL.n35 2.26352
R16512 VCO_DFF_C_0.VCTRL.n19 VCO_DFF_C_0.VCTRL.t22 2.17312
R16513 VCO_DFF_C_0.VCTRL.n4 VCO_DFF_C_0.VCTRL.t35 2.17312
R16514 VCO_DFF_C_0.VCTRL.n7 VCO_DFF_C_0.VCTRL.t25 2.17312
R16515 VCO_DFF_C_0.VCTRL.n17 VCO_DFF_C_0.VCTRL.t33 2.17312
R16516 VCO_DFF_C_0.VCTRL.n37 VCO_DFF_C_0.VCTRL.t2 2.16717
R16517 VCO_DFF_C_0.VCTRL.n37 VCO_DFF_C_0.VCTRL.n36 2.16717
R16518 VCO_DFF_C_0.VCTRL.n33 VCO_DFF_C_0.VCTRL.t1 2.16717
R16519 VCO_DFF_C_0.VCTRL.n33 VCO_DFF_C_0.VCTRL.n32 2.16717
R16520 VCO_DFF_C_0.VCTRL.n45 VCO_DFF_C_0.VCTRL.t8 2.16717
R16521 VCO_DFF_C_0.VCTRL.n45 VCO_DFF_C_0.VCTRL.n44 2.16717
R16522 VCO_DFF_C_0.VCTRL.n43 VCO_DFF_C_0.VCTRL.t6 2.16717
R16523 VCO_DFF_C_0.VCTRL.n43 VCO_DFF_C_0.VCTRL.n42 2.16717
R16524 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCTRL.n28 1.89901
R16525 VCO_DFF_C_0.VCTRL.n26 VCO_DFF_C_0.VCTRL.n25 1.896
R16526 VCO_DFF_C_0.VCTRL.n13 VCO_DFF_C_0.VCTRL.n12 1.89145
R16527 VCO_DFF_C_0.VCTRL.n51 VCO_DFF_C_0.VCTRL.n50 1.84797
R16528 VCO_DFF_C_0.VCTRL.n3 VCO_DFF_C_0.VCTRL.n39 1.82978
R16529 VCO_DFF_C_0.VCTRL.n27 VCO_DFF_C_0.VCTRL.n26 1.5395
R16530 VCO_DFF_C_0.VCTRL.n14 VCO_DFF_C_0.VCTRL.n13 1.5395
R16531 VCO_DFF_C_0.VCTRL.n29 VCO_DFF_C_0.VCTRL 1.4706
R16532 VCO_DFF_C_0.VCTRL.n2 VCO_DFF_C_0.VCTRL 0.663665
R16533 VCO_DFF_C_0.VCTRL.n2 VCO_DFF_C_0.VCTRL.n31 1.25555
R16534 VCO_DFF_C_0.VCTRL.n46 VCO_DFF_C_0.VCTRL.n45 1.25233
R16535 VCO_DFF_C_0.VCTRL.n51 VCO_DFF_C_0.VCTRL.n46 1.12574
R16536 VCO_DFF_C_0.VCTRL.n11 VCO_DFF_C_0.VCTRL.n10 1.05913
R16537 VCO_DFF_C_0.VCTRL.n13 VCO_DFF_C_0.VCTRL.n6 0.957464
R16538 VCO_DFF_C_0.VCTRL.n26 VCO_DFF_C_0.VCTRL.n23 0.95722
R16539 VCO_DFF_C_0.VCTRL.n16 VCO_DFF_C_0.VCTRL.n15 0.798473
R16540 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCTRL.n52 0.751569
R16541 VCO_DFF_C_0.VCTRL.n9 VCO_DFF_C_0.VCTRL.n8 0.749817
R16542 VCO_DFF_C_0.VCTRL.n22 VCO_DFF_C_0.VCTRL.n21 0.749568
R16543 VCO_DFF_C_0.VCTRL.n40 VCO_DFF_C_0.VCTRL 0.736653
R16544 VCO_DFF_C_0.VCTRL.n23 VCO_DFF_C_0.VCTRL.n22 0.622921
R16545 VCO_DFF_C_0.VCTRL.n8 VCO_DFF_C_0.VCTRL.n6 0.622675
R16546 VCO_DFF_C_0.VCTRL.n21 VCO_DFF_C_0.VCTRL.n20 0.602194
R16547 VCO_DFF_C_0.VCTRL.n10 VCO_DFF_C_0.VCTRL.n9 0.602194
R16548 VCO_DFF_C_0.VCTRL.n50 VCO_DFF_C_0.VCTRL.n1 0.558374
R16549 VCO_DFF_C_0.VCTRL.n39 VCO_DFF_C_0.VCTRL.n0 0.558372
R16550 VCO_DFF_C_0.VCTRL.n29 VCO_DFF_C_0.VCTRL 0.550625
R16551 VCO_DFF_C_0.VCTRL.n12 VCO_DFF_C_0.VCTRL.n11 0.453053
R16552 VCO_DFF_C_0.VCTRL.n25 VCO_DFF_C_0.VCTRL.n24 0.451515
R16553 VCO_DFF_C_0.VCTRL.n15 VCO_DFF_C_0.VCTRL.n14 0.43025
R16554 VCO_DFF_C_0.VCTRL.n28 VCO_DFF_C_0.VCTRL.n27 0.43025
R16555 VCO_DFF_C_0.VCTRL.n40 VCO_DFF_C_0.VCTRL.n3 0.394824
R16556 VCO_DFF_C_0.VCTRL.n52 VCO_DFF_C_0.VCTRL.n51 0.33941
R16557 VCO_DFF_C_0.VCTRL.n14 VCO_DFF_C_0.VCTRL.n5 0.266
R16558 VCO_DFF_C_0.VCTRL.n27 VCO_DFF_C_0.VCTRL.n18 0.266
R16559 VCO_DFF_C_0.VCTRL.n41 VCO_DFF_C_0.VCTRL.n2 0.25987
R16560 VCO_DFF_C_0.VCTRL.n31 VCO_DFF_C_0.VCTRL.n30 0.23889
R16561 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCTRL.n29 0.195324
R16562 VCO_DFF_C_0.VCTRL.n35 VCO_DFF_C_0.VCTRL.n34 0.145661
R16563 a_22967_8787.n0 a_22967_8787.t14 33.8126
R16564 a_22967_8787.n1 a_22967_8787.n0 30.3299
R16565 a_22967_8787.n2 a_22967_8787.n1 30.3299
R16566 a_22967_8787.n3 a_22967_8787.n2 30.3299
R16567 a_22967_8787.n4 a_22967_8787.n3 30.3299
R16568 a_22967_8787.n5 a_22967_8787.n4 30.3299
R16569 a_22967_8787.n6 a_22967_8787.n5 30.3299
R16570 a_22967_8787.n7 a_22967_8787.n6 30.3299
R16571 a_22967_8787.n8 a_22967_8787.n7 30.3299
R16572 a_22967_8787.n12 a_22967_8787.t7 26.2202
R16573 a_22967_8787.n9 a_22967_8787.t6 12.8368
R16574 a_22967_8787.n9 a_22967_8787.n8 12.0257
R16575 a_22967_8787.n13 a_22967_8787.n12 8.40022
R16576 a_22967_8787.n14 a_22967_8787.n9 5.21471
R16577 a_22967_8787.n12 a_22967_8787.t15 3.6505
R16578 a_22967_8787.n0 a_22967_8787.t4 3.6505
R16579 a_22967_8787.n1 a_22967_8787.t11 3.6505
R16580 a_22967_8787.n2 a_22967_8787.t5 3.6505
R16581 a_22967_8787.n3 a_22967_8787.t12 3.6505
R16582 a_22967_8787.n4 a_22967_8787.t9 3.6505
R16583 a_22967_8787.n5 a_22967_8787.t16 3.6505
R16584 a_22967_8787.n6 a_22967_8787.t10 3.6505
R16585 a_22967_8787.n7 a_22967_8787.t13 3.6505
R16586 a_22967_8787.n8 a_22967_8787.t8 3.6505
R16587 a_22967_8787.n15 a_22967_8787.t0 3.6405
R16588 a_22967_8787.n16 a_22967_8787.n15 3.6405
R16589 a_22967_8787.n14 a_22967_8787.n13 3.38778
R16590 a_22967_8787.n11 a_22967_8787.t3 3.38774
R16591 a_22967_8787.n11 a_22967_8787.n10 2.97656
R16592 a_22967_8787.n13 a_22967_8787.n11 2.47435
R16593 a_22967_8787.n15 a_22967_8787.n14 1.25578
R16594 a_50810_1389.n26 a_50810_1389.n25 72.9524
R16595 a_50810_1389.n20 a_50810_1389.t21 44.8231
R16596 a_50810_1389.n2 a_50810_1389.t13 36.4904
R16597 a_50810_1389.n26 a_50810_1389.t7 23.7985
R16598 a_50810_1389.n2 a_50810_1389.t20 23.6525
R16599 a_50810_1389.n3 a_50810_1389.t8 23.6525
R16600 a_50810_1389.n4 a_50810_1389.t14 23.6525
R16601 a_50810_1389.n5 a_50810_1389.t17 23.6525
R16602 a_50810_1389.n6 a_50810_1389.t28 23.6525
R16603 a_50810_1389.n7 a_50810_1389.t18 23.6525
R16604 a_50810_1389.n8 a_50810_1389.t29 23.6525
R16605 a_50810_1389.n9 a_50810_1389.t26 23.6525
R16606 a_50810_1389.n10 a_50810_1389.t16 23.6525
R16607 a_50810_1389.n11 a_50810_1389.t27 23.6525
R16608 a_50810_1389.n12 a_50810_1389.t11 23.6525
R16609 a_50810_1389.n13 a_50810_1389.t24 23.6525
R16610 a_50810_1389.n14 a_50810_1389.t22 23.6525
R16611 a_50810_1389.n15 a_50810_1389.t10 23.6525
R16612 a_50810_1389.n16 a_50810_1389.t23 23.6525
R16613 a_50810_1389.n21 a_50810_1389.n20 23.3438
R16614 a_50810_1389.n22 a_50810_1389.n21 23.3438
R16615 a_50810_1389.n23 a_50810_1389.n22 23.3438
R16616 a_50810_1389.n24 a_50810_1389.n23 23.3438
R16617 a_50810_1389.n25 a_50810_1389.n24 23.3438
R16618 a_50810_1389.n20 a_50810_1389.t9 20.4405
R16619 a_50810_1389.n21 a_50810_1389.t15 20.4405
R16620 a_50810_1389.n22 a_50810_1389.t19 20.4405
R16621 a_50810_1389.n23 a_50810_1389.t6 20.4405
R16622 a_50810_1389.n24 a_50810_1389.t12 20.4405
R16623 a_50810_1389.n25 a_50810_1389.t25 20.4405
R16624 a_50810_1389.n3 a_50810_1389.n2 12.8384
R16625 a_50810_1389.n4 a_50810_1389.n3 12.8384
R16626 a_50810_1389.n5 a_50810_1389.n4 12.8384
R16627 a_50810_1389.n6 a_50810_1389.n5 12.8384
R16628 a_50810_1389.n7 a_50810_1389.n6 12.8384
R16629 a_50810_1389.n8 a_50810_1389.n7 12.8384
R16630 a_50810_1389.n9 a_50810_1389.n8 12.8384
R16631 a_50810_1389.n10 a_50810_1389.n9 12.8384
R16632 a_50810_1389.n11 a_50810_1389.n10 12.8384
R16633 a_50810_1389.n12 a_50810_1389.n11 12.8384
R16634 a_50810_1389.n13 a_50810_1389.n12 12.8384
R16635 a_50810_1389.n14 a_50810_1389.n13 12.8384
R16636 a_50810_1389.n15 a_50810_1389.n14 12.8384
R16637 a_50810_1389.n16 a_50810_1389.n15 12.8384
R16638 a_50810_1389.n27 a_50810_1389.n26 6.95492
R16639 a_50810_1389.n17 a_50810_1389.n16 4.78319
R16640 a_50810_1389.n28 a_50810_1389.n27 4.13676
R16641 a_50810_1389.n27 a_50810_1389.n19 3.79615
R16642 a_50810_1389.n17 a_50810_1389.n1 3.22711
R16643 a_50810_1389.n29 a_50810_1389.n28 3.22482
R16644 a_50810_1389.n1 a_50810_1389.t2 0.6505
R16645 a_50810_1389.n1 a_50810_1389.n0 0.6505
R16646 a_50810_1389.n29 a_50810_1389.t4 0.6505
R16647 a_50810_1389.n30 a_50810_1389.n29 0.6505
R16648 a_50810_1389.n19 a_50810_1389.t3 0.5855
R16649 a_50810_1389.n19 a_50810_1389.n18 0.5855
R16650 a_50810_1389.n28 a_50810_1389.n17 0.471269
R16651 PFD_T2_0.FIN.n11 PFD_T2_0.FIN.t18 12.4835
R16652 PFD_T2_0.FIN.n13 PFD_T2_0.FIN.t17 11.5345
R16653 PFD_T2_0.FIN.n11 PFD_T2_0.FIN.t16 11.4615
R16654 PFD_T2_0.FIN.n12 PFD_T2_0.FIN.t19 11.4615
R16655 PFD_T2_0.FIN.n12 PFD_T2_0.FIN.n11 10.6935
R16656 PFD_T2_0.FIN.n0 PFD_T2_0.FIN.t9 6.74332
R16657 PFD_T2_0.FIN.n1 PFD_T2_0.FIN.n21 6.74326
R16658 PFD_T2_0.FIN PFD_T2_0.FIN.n13 5.16904
R16659 PFD_T2_0.FIN.n1 PFD_T2_0.FIN.n22 5.1005
R16660 PFD_T2_0.FIN.n0 PFD_T2_0.FIN.t10 5.1005
R16661 PFD_T2_0.FIN.n8 PFD_T2_0.FIN.n7 3.5743
R16662 PFD_T2_0.FIN.n19 PFD_T2_0.FIN.n18 3.5743
R16663 PFD_T2_0.FIN.n1 PFD_T2_0.FIN.t15 3.40065
R16664 PFD_T2_0.FIN.n0 PFD_T2_0.FIN.n2 3.40001
R16665 PFD_T2_0.FIN.n3 PFD_T2_0.FIN.t8 3.00159
R16666 PFD_T2_0.FIN.n23 PFD_T2_0.FIN.n20 3.00034
R16667 PFD_T2_0.FIN PFD_T2_0.FIN.n26 2.60984
R16668 PFD_T2_0.FIN.n26 PFD_T2_0.FIN.n14 2.46176
R16669 PFD_T2_0.FIN.n26 PFD_T2_0.FIN.n25 2.36206
R16670 PFD_T2_0.FIN.n5 PFD_T2_0.FIN.t3 2.16717
R16671 PFD_T2_0.FIN.n5 PFD_T2_0.FIN.n4 2.16717
R16672 PFD_T2_0.FIN.n7 PFD_T2_0.FIN.t0 2.16717
R16673 PFD_T2_0.FIN.n7 PFD_T2_0.FIN.n6 2.16717
R16674 PFD_T2_0.FIN.n16 PFD_T2_0.FIN.t7 2.16717
R16675 PFD_T2_0.FIN.n16 PFD_T2_0.FIN.n15 2.16717
R16676 PFD_T2_0.FIN.n18 PFD_T2_0.FIN.t6 2.16717
R16677 PFD_T2_0.FIN.n18 PFD_T2_0.FIN.n17 2.16717
R16678 PFD_T2_0.FIN.n9 PFD_T2_0.FIN.n3 1.84725
R16679 PFD_T2_0.FIN.n24 PFD_T2_0.FIN.n23 1.847
R16680 PFD_T2_0.FIN.n14 PFD_T2_0.FIN 1.50801
R16681 PFD_T2_0.FIN.n8 PFD_T2_0.FIN.n5 1.25225
R16682 PFD_T2_0.FIN.n19 PFD_T2_0.FIN.n16 1.25225
R16683 PFD_T2_0.FIN.n24 PFD_T2_0.FIN.n19 1.12594
R16684 PFD_T2_0.FIN.n9 PFD_T2_0.FIN.n8 1.12575
R16685 PFD_T2_0.FIN.n13 PFD_T2_0.FIN.n12 0.9495
R16686 PFD_T2_0.FIN.n25 PFD_T2_0.FIN 0.751569
R16687 PFD_T2_0.FIN.n10 PFD_T2_0.FIN 0.737159
R16688 PFD_T2_0.FIN.n23 PFD_T2_0.FIN.n1 0.559412
R16689 PFD_T2_0.FIN.n3 PFD_T2_0.FIN.n0 0.55941
R16690 PFD_T2_0.FIN.n10 PFD_T2_0.FIN.n9 0.377914
R16691 PFD_T2_0.FIN.n25 PFD_T2_0.FIN.n24 0.33941
R16692 PFD_T2_0.FIN.n14 PFD_T2_0.FIN.n10 0.28138
R16693 PRE_SCALAR.n7 PRE_SCALAR.t2 5.81586
R16694 PRE_SCALAR.n4 PRE_SCALAR.n1 5.10151
R16695 PRE_SCALAR.n11 PRE_SCALAR.n10 5.10119
R16696 PRE_SCALAR.n9 PRE_SCALAR.n8 5.08021
R16697 PRE_SCALAR.n4 PRE_SCALAR.n3 4.66164
R16698 PRE_SCALAR.n7 PRE_SCALAR.n6 2.85093
R16699 PRE_SCALAR.n6 PRE_SCALAR.t1 2.16717
R16700 PRE_SCALAR.n6 PRE_SCALAR.n5 2.16717
R16701 PRE_SCALAR.n3 PRE_SCALAR.t4 1.9505
R16702 PRE_SCALAR.n3 PRE_SCALAR.n2 1.9505
R16703 PRE_SCALAR PRE_SCALAR.n0 1.47796
R16704 PRE_SCALAR.n0 PRE_SCALAR 1.47444
R16705 PRE_SCALAR.n0 PRE_SCALAR 0.838578
R16706 PRE_SCALAR.n9 PRE_SCALAR.n7 0.644196
R16707 PRE_SCALAR.n11 PRE_SCALAR.n9 0.4508
R16708 PRE_SCALAR.n12 PRE_SCALAR.n4 0.309543
R16709 PRE_SCALAR.n12 PRE_SCALAR.n11 0.274999
R16710 PRE_SCALAR PRE_SCALAR.n12 0.0936034
R16711 S6.n14 S6.t18 45.6363
R16712 S6.n0 S6.t5 29.6446
R16713 S6.t16 S6.n1 29.6446
R16714 S6.n2 S6.t12 24.6117
R16715 S6.n8 S6.t20 23.6945
R16716 S6.n9 S6.t1 23.6945
R16717 S6.n1 S6.n0 22.2047
R16718 S6.t18 S6.t11 22.1925
R16719 S6.n15 S6.n14 20.9314
R16720 S6.n9 S6.n8 18.8035
R16721 S6 S6.t16 18.5175
R16722 S6.n6 S6.n3 15.8172
R16723 S6.n12 S6.n11 15.8172
R16724 S6.n11 S6.n3 15.8172
R16725 S6.t6 S6.n6 14.8925
R16726 S6.t21 S6.n3 14.8925
R16727 S6.n11 S6.t4 14.8925
R16728 S6.n10 S6.n4 12.2457
R16729 S6.n10 S6.n5 12.2457
R16730 S6.n7 S6.n5 12.2457
R16731 S6.n13 S6.t9 11.6285
R16732 S6.t20 S6.n7 8.9065
R16733 S6.t7 S6.n5 8.9065
R16734 S6.n10 S6.t15 8.9065
R16735 S6.t1 S6.n4 8.9065
R16736 S6.n6 S6.t0 8.6145
R16737 S6.n3 S6.t10 8.6145
R16738 S6.n11 S6.t17 8.6145
R16739 S6.n12 S6.t2 8.59715
R16740 S6.n7 S6.t6 8.3225
R16741 S6.n5 S6.t21 8.3225
R16742 S6.t4 S6.n10 8.3225
R16743 S6.n4 S6.t9 8.3225
R16744 S6.n2 S6.t8 6.1325
R16745 S6.n0 S6.t3 6.1325
R16746 S6.n1 S6.t13 6.1325
R16747 S6.n14 S6.t19 6.1325
R16748 S6.n15 S6.t14 6.1325
R16749 S6.n17 S6.n15 4.86779
R16750 S6.n19 S6.n2 4.79907
R16751 S6 S6.n13 4.223
R16752 S6.n8 S6.t7 3.6505
R16753 S6.t15 S6.n9 3.6505
R16754 S6.n13 S6.n12 3.1807
R16755 S6.n17 S6.n16 1.49668
R16756 S6.n16 S6 0.992377
R16757 S6.n16 S6 0.850469
R16758 S6 S6.n19 0.640368
R16759 S6.n18 S6 0.1655
R16760 S6.n18 S6.n17 0.109537
R16761 S6.n19 S6.n18 0.0592755
R16762 A_MUX_2.Tr_Gate_1.CLK.n1 A_MUX_2.Tr_Gate_1.CLK.t19 45.6363
R16763 A_MUX_2.Tr_Gate_1.CLK.n3 A_MUX_2.Tr_Gate_1.CLK.t17 29.6446
R16764 A_MUX_2.Tr_Gate_1.CLK.t15 A_MUX_2.Tr_Gate_1.CLK.n4 29.6446
R16765 A_MUX_2.Tr_Gate_1.CLK.n5 A_MUX_2.Tr_Gate_1.CLK.t13 24.6117
R16766 A_MUX_2.Tr_Gate_1.CLK.n4 A_MUX_2.Tr_Gate_1.CLK.n3 22.2047
R16767 A_MUX_2.Tr_Gate_1.CLK.t19 A_MUX_2.Tr_Gate_1.CLK.t14 22.1925
R16768 A_MUX_2.Tr_Gate_1.CLK.n2 A_MUX_2.Tr_Gate_1.CLK.n1 20.9314
R16769 A_MUX_2.Tr_Gate_1.CLK A_MUX_2.Tr_Gate_1.CLK.t15 18.5231
R16770 A_MUX_2.Tr_Gate_1.CLK.n5 A_MUX_2.Tr_Gate_1.CLK.t16 6.1325
R16771 A_MUX_2.Tr_Gate_1.CLK.n3 A_MUX_2.Tr_Gate_1.CLK.t20 6.1325
R16772 A_MUX_2.Tr_Gate_1.CLK.n4 A_MUX_2.Tr_Gate_1.CLK.t12 6.1325
R16773 A_MUX_2.Tr_Gate_1.CLK.n1 A_MUX_2.Tr_Gate_1.CLK.t18 6.1325
R16774 A_MUX_2.Tr_Gate_1.CLK.n2 A_MUX_2.Tr_Gate_1.CLK.t21 6.1325
R16775 A_MUX_2.Tr_Gate_1.CLK.n0 A_MUX_2.Tr_Gate_1.CLK.n2 5.28481
R16776 A_MUX_2.Tr_Gate_1.CLK.n0 A_MUX_2.Tr_Gate_1.CLK.n5 4.89628
R16777 A_MUX_2.Tr_Gate_1.CLK.n18 A_MUX_2.Tr_Gate_1.CLK.t10 3.6405
R16778 A_MUX_2.Tr_Gate_1.CLK.n18 A_MUX_2.Tr_Gate_1.CLK.n17 3.6405
R16779 A_MUX_2.Tr_Gate_1.CLK.n9 A_MUX_2.Tr_Gate_1.CLK.t9 3.6405
R16780 A_MUX_2.Tr_Gate_1.CLK.n9 A_MUX_2.Tr_Gate_1.CLK.n8 3.6405
R16781 A_MUX_2.Tr_Gate_1.CLK.n7 A_MUX_2.Tr_Gate_1.CLK.t5 3.6405
R16782 A_MUX_2.Tr_Gate_1.CLK.n7 A_MUX_2.Tr_Gate_1.CLK.n6 3.6405
R16783 A_MUX_2.Tr_Gate_1.CLK.n16 A_MUX_2.Tr_Gate_1.CLK.t6 3.6405
R16784 A_MUX_2.Tr_Gate_1.CLK.n16 A_MUX_2.Tr_Gate_1.CLK.n15 3.6405
R16785 A_MUX_2.Tr_Gate_1.CLK.n20 A_MUX_2.Tr_Gate_1.CLK.n14 3.50463
R16786 A_MUX_2.Tr_Gate_1.CLK.n21 A_MUX_2.Tr_Gate_1.CLK.n12 3.50463
R16787 A_MUX_2.Tr_Gate_1.CLK.n14 A_MUX_2.Tr_Gate_1.CLK.t0 3.2765
R16788 A_MUX_2.Tr_Gate_1.CLK.n14 A_MUX_2.Tr_Gate_1.CLK.n13 3.2765
R16789 A_MUX_2.Tr_Gate_1.CLK.n12 A_MUX_2.Tr_Gate_1.CLK.t3 3.2765
R16790 A_MUX_2.Tr_Gate_1.CLK.n12 A_MUX_2.Tr_Gate_1.CLK.n11 3.2765
R16791 A_MUX_2.Tr_Gate_1.CLK.n10 A_MUX_2.Tr_Gate_1.CLK.n7 3.06224
R16792 A_MUX_2.Tr_Gate_1.CLK.n19 A_MUX_2.Tr_Gate_1.CLK.n16 3.06224
R16793 A_MUX_2.Tr_Gate_1.CLK.n10 A_MUX_2.Tr_Gate_1.CLK.n9 2.6005
R16794 A_MUX_2.Tr_Gate_1.CLK.n19 A_MUX_2.Tr_Gate_1.CLK.n18 2.6005
R16795 A_MUX_2.Tr_Gate_1.CLK.n21 A_MUX_2.Tr_Gate_1.CLK.n20 0.798761
R16796 A_MUX_2.Tr_Gate_1.CLK.n0 A_MUX_2.Tr_Gate_1.CLK 0.629606
R16797 A_MUX_2.Tr_Gate_1.CLK A_MUX_2.Tr_Gate_1.CLK.n21 0.562022
R16798 A_MUX_2.Tr_Gate_1.CLK A_MUX_2.Tr_Gate_1.CLK.n0 0.253378
R16799 A_MUX_2.Tr_Gate_1.CLK.n21 A_MUX_2.Tr_Gate_1.CLK.n10 0.18637
R16800 A_MUX_2.Tr_Gate_1.CLK.n20 A_MUX_2.Tr_Gate_1.CLK.n19 0.18637
R16801 VCO_DFF_C_0.VCO_C_0.OUTB.n20 VCO_DFF_C_0.VCO_C_0.OUTB.t47 45.6363
R16802 VCO_DFF_C_0.VCO_C_0.OUTB.n26 VCO_DFF_C_0.VCO_C_0.OUTB.t35 45.6363
R16803 VCO_DFF_C_0.VCO_C_0.OUTB.n23 VCO_DFF_C_0.VCO_C_0.OUTB.t48 29.6446
R16804 VCO_DFF_C_0.VCO_C_0.OUTB.t51 VCO_DFF_C_0.VCO_C_0.OUTB.n24 29.6446
R16805 VCO_DFF_C_0.VCO_C_0.OUTB.n29 VCO_DFF_C_0.VCO_C_0.OUTB.t43 29.6446
R16806 VCO_DFF_C_0.VCO_C_0.OUTB.t41 VCO_DFF_C_0.VCO_C_0.OUTB.n30 29.6446
R16807 VCO_DFF_C_0.VCO_C_0.OUTB.n19 VCO_DFF_C_0.VCO_C_0.OUTB.t33 24.6117
R16808 VCO_DFF_C_0.VCO_C_0.OUTB.n28 VCO_DFF_C_0.VCO_C_0.OUTB.t32 24.6117
R16809 VCO_DFF_C_0.VCO_C_0.OUTB.n40 VCO_DFF_C_0.VCO_C_0.OUTB.t28 23.6945
R16810 VCO_DFF_C_0.VCO_C_0.OUTB.t16 VCO_DFF_C_0.VCO_C_0.OUTB.n41 23.6945
R16811 VCO_DFF_C_0.VCO_C_0.OUTB.n24 VCO_DFF_C_0.VCO_C_0.OUTB.n23 22.2047
R16812 VCO_DFF_C_0.VCO_C_0.OUTB.n30 VCO_DFF_C_0.VCO_C_0.OUTB.n29 22.2047
R16813 VCO_DFF_C_0.VCO_C_0.OUTB.t47 VCO_DFF_C_0.VCO_C_0.OUTB.t15 22.1925
R16814 VCO_DFF_C_0.VCO_C_0.OUTB.t35 VCO_DFF_C_0.VCO_C_0.OUTB.t46 22.1925
R16815 VCO_DFF_C_0.VCO_C_0.OUTB.n21 VCO_DFF_C_0.VCO_C_0.OUTB.n20 20.9314
R16816 VCO_DFF_C_0.VCO_C_0.OUTB.n27 VCO_DFF_C_0.VCO_C_0.OUTB.n26 20.9314
R16817 VCO_DFF_C_0.VCO_C_0.OUTB.n41 VCO_DFF_C_0.VCO_C_0.OUTB.n40 18.8035
R16818 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.t41 18.5191
R16819 VCO_DFF_C_0.VCO_C_0.OUTB.n25 VCO_DFF_C_0.VCO_C_0.OUTB.t51 17.9055
R16820 VCO_DFF_C_0.VCO_C_0.OUTB.n38 VCO_DFF_C_0.VCO_C_0.OUTB.n36 15.8172
R16821 VCO_DFF_C_0.VCO_C_0.OUTB.n38 VCO_DFF_C_0.VCO_C_0.OUTB.n37 15.8172
R16822 VCO_DFF_C_0.VCO_C_0.OUTB.n37 VCO_DFF_C_0.VCO_C_0.OUTB.n33 15.8172
R16823 VCO_DFF_C_0.VCO_C_0.OUTB.n46 VCO_DFF_C_0.VCO_C_0.OUTB.t14 15.4917
R16824 VCO_DFF_C_0.VCO_C_0.OUTB.n48 VCO_DFF_C_0.VCO_C_0.OUTB.t18 15.3942
R16825 VCO_DFF_C_0.VCO_C_0.OUTB.n49 VCO_DFF_C_0.VCO_C_0.OUTB.t38 14.9265
R16826 VCO_DFF_C_0.VCO_C_0.OUTB.n36 VCO_DFF_C_0.VCO_C_0.OUTB.t52 14.8925
R16827 VCO_DFF_C_0.VCO_C_0.OUTB.t27 VCO_DFF_C_0.VCO_C_0.OUTB.n38 14.8925
R16828 VCO_DFF_C_0.VCO_C_0.OUTB.n37 VCO_DFF_C_0.VCO_C_0.OUTB.t17 14.8925
R16829 VCO_DFF_C_0.VCO_C_0.OUTB.n53 VCO_DFF_C_0.VCO_C_0.OUTB.t31 14.7749
R16830 VCO_DFF_C_0.VCO_C_0.OUTB.n47 VCO_DFF_C_0.VCO_C_0.OUTB.t50 13.6019
R16831 VCO_DFF_C_0.VCO_C_0.OUTB.n53 VCO_DFF_C_0.VCO_C_0.OUTB.t23 13.5312
R16832 VCO_DFF_C_0.VCO_C_0.OUTB.n51 VCO_DFF_C_0.VCO_C_0.OUTB.t42 13.4877
R16833 VCO_DFF_C_0.VCO_C_0.OUTB.n49 VCO_DFF_C_0.VCO_C_0.OUTB.t30 13.227
R16834 VCO_DFF_C_0.VCO_C_0.OUTB.n50 VCO_DFF_C_0.VCO_C_0.OUTB.t26 13.1835
R16835 VCO_DFF_C_0.VCO_C_0.OUTB.n42 VCO_DFF_C_0.VCO_C_0.OUTB.n34 12.2457
R16836 VCO_DFF_C_0.VCO_C_0.OUTB.n39 VCO_DFF_C_0.VCO_C_0.OUTB.n34 12.2457
R16837 VCO_DFF_C_0.VCO_C_0.OUTB.n39 VCO_DFF_C_0.VCO_C_0.OUTB.n35 12.2457
R16838 VCO_DFF_C_0.VCO_C_0.OUTB.n43 VCO_DFF_C_0.VCO_C_0.OUTB.t36 11.6285
R16839 VCO_DFF_C_0.VCO_C_0.OUTB.n45 VCO_DFF_C_0.VCO_C_0.OUTB.n2 9.0064
R16840 VCO_DFF_C_0.VCO_C_0.OUTB.n35 VCO_DFF_C_0.VCO_C_0.OUTB.t28 8.9065
R16841 VCO_DFF_C_0.VCO_C_0.OUTB.t49 VCO_DFF_C_0.VCO_C_0.OUTB.n39 8.9065
R16842 VCO_DFF_C_0.VCO_C_0.OUTB.t37 VCO_DFF_C_0.VCO_C_0.OUTB.n34 8.9065
R16843 VCO_DFF_C_0.VCO_C_0.OUTB.n42 VCO_DFF_C_0.VCO_C_0.OUTB.t16 8.9065
R16844 VCO_DFF_C_0.VCO_C_0.OUTB.n38 VCO_DFF_C_0.VCO_C_0.OUTB.t24 8.6145
R16845 VCO_DFF_C_0.VCO_C_0.OUTB.n36 VCO_DFF_C_0.VCO_C_0.OUTB.t45 8.6145
R16846 VCO_DFF_C_0.VCO_C_0.OUTB.n37 VCO_DFF_C_0.VCO_C_0.OUTB.t13 8.6145
R16847 VCO_DFF_C_0.VCO_C_0.OUTB.n33 VCO_DFF_C_0.VCO_C_0.OUTB.t34 8.59715
R16848 VCO_DFF_C_0.VCO_C_0.OUTB.t52 VCO_DFF_C_0.VCO_C_0.OUTB.n35 8.3225
R16849 VCO_DFF_C_0.VCO_C_0.OUTB.n39 VCO_DFF_C_0.VCO_C_0.OUTB.t27 8.3225
R16850 VCO_DFF_C_0.VCO_C_0.OUTB.t17 VCO_DFF_C_0.VCO_C_0.OUTB.n34 8.3225
R16851 VCO_DFF_C_0.VCO_C_0.OUTB.t36 VCO_DFF_C_0.VCO_C_0.OUTB.n42 8.3225
R16852 VCO_DFF_C_0.VCO_C_0.OUTB.n2 VCO_DFF_C_0.VCO_C_0.OUTB.n25 8.24338
R16853 VCO_DFF_C_0.VCO_C_0.OUTB.n46 VCO_DFF_C_0.VCO_C_0.OUTB.t53 8.1387
R16854 VCO_DFF_C_0.VCO_C_0.OUTB.n23 VCO_DFF_C_0.VCO_C_0.OUTB.t40 6.1325
R16855 VCO_DFF_C_0.VCO_C_0.OUTB.n24 VCO_DFF_C_0.VCO_C_0.OUTB.t44 6.1325
R16856 VCO_DFF_C_0.VCO_C_0.OUTB.n19 VCO_DFF_C_0.VCO_C_0.OUTB.t22 6.1325
R16857 VCO_DFF_C_0.VCO_C_0.OUTB.n20 VCO_DFF_C_0.VCO_C_0.OUTB.t21 6.1325
R16858 VCO_DFF_C_0.VCO_C_0.OUTB.n21 VCO_DFF_C_0.VCO_C_0.OUTB.t12 6.1325
R16859 VCO_DFF_C_0.VCO_C_0.OUTB.n28 VCO_DFF_C_0.VCO_C_0.OUTB.t39 6.1325
R16860 VCO_DFF_C_0.VCO_C_0.OUTB.n29 VCO_DFF_C_0.VCO_C_0.OUTB.t25 6.1325
R16861 VCO_DFF_C_0.VCO_C_0.OUTB.n30 VCO_DFF_C_0.VCO_C_0.OUTB.t19 6.1325
R16862 VCO_DFF_C_0.VCO_C_0.OUTB.n26 VCO_DFF_C_0.VCO_C_0.OUTB.t20 6.1325
R16863 VCO_DFF_C_0.VCO_C_0.OUTB.n27 VCO_DFF_C_0.VCO_C_0.OUTB.t29 6.1325
R16864 VCO_DFF_C_0.VCO_C_0.OUTB.n32 VCO_DFF_C_0.VCO_C_0.OUTB.n27 5.5044
R16865 VCO_DFF_C_0.VCO_C_0.OUTB.n22 VCO_DFF_C_0.VCO_C_0.OUTB.n21 5.38991
R16866 VCO_DFF_C_0.VCO_C_0.OUTB.n22 VCO_DFF_C_0.VCO_C_0.OUTB.n19 4.83094
R16867 VCO_DFF_C_0.VCO_C_0.OUTB.n31 VCO_DFF_C_0.VCO_C_0.OUTB.n28 4.83094
R16868 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n43 4.223
R16869 VCO_DFF_C_0.VCO_C_0.OUTB.n40 VCO_DFF_C_0.VCO_C_0.OUTB.t49 3.6505
R16870 VCO_DFF_C_0.VCO_C_0.OUTB.n41 VCO_DFF_C_0.VCO_C_0.OUTB.t37 3.6505
R16871 VCO_DFF_C_0.VCO_C_0.OUTB.n14 VCO_DFF_C_0.VCO_C_0.OUTB.t8 3.6405
R16872 VCO_DFF_C_0.VCO_C_0.OUTB.n14 VCO_DFF_C_0.VCO_C_0.OUTB.n13 3.6405
R16873 VCO_DFF_C_0.VCO_C_0.OUTB.n8 VCO_DFF_C_0.VCO_C_0.OUTB.t10 3.6405
R16874 VCO_DFF_C_0.VCO_C_0.OUTB.n8 VCO_DFF_C_0.VCO_C_0.OUTB.n7 3.6405
R16875 VCO_DFF_C_0.VCO_C_0.OUTB.n10 VCO_DFF_C_0.VCO_C_0.OUTB.t6 3.6405
R16876 VCO_DFF_C_0.VCO_C_0.OUTB.n10 VCO_DFF_C_0.VCO_C_0.OUTB.n9 3.6405
R16877 VCO_DFF_C_0.VCO_C_0.OUTB.n16 VCO_DFF_C_0.VCO_C_0.OUTB.t5 3.6405
R16878 VCO_DFF_C_0.VCO_C_0.OUTB.n16 VCO_DFF_C_0.VCO_C_0.OUTB.n15 3.6405
R16879 VCO_DFF_C_0.VCO_C_0.OUTB.n18 VCO_DFF_C_0.VCO_C_0.OUTB.n4 3.50463
R16880 VCO_DFF_C_0.VCO_C_0.OUTB.n12 VCO_DFF_C_0.VCO_C_0.OUTB.n6 3.50463
R16881 VCO_DFF_C_0.VCO_C_0.OUTB.n4 VCO_DFF_C_0.VCO_C_0.OUTB.t1 3.2765
R16882 VCO_DFF_C_0.VCO_C_0.OUTB.n4 VCO_DFF_C_0.VCO_C_0.OUTB.n3 3.2765
R16883 VCO_DFF_C_0.VCO_C_0.OUTB.n6 VCO_DFF_C_0.VCO_C_0.OUTB.t3 3.2765
R16884 VCO_DFF_C_0.VCO_C_0.OUTB.n6 VCO_DFF_C_0.VCO_C_0.OUTB.n5 3.2765
R16885 VCO_DFF_C_0.VCO_C_0.OUTB.n43 VCO_DFF_C_0.VCO_C_0.OUTB.n33 3.1807
R16886 VCO_DFF_C_0.VCO_C_0.OUTB.n11 VCO_DFF_C_0.VCO_C_0.OUTB.n10 3.06224
R16887 VCO_DFF_C_0.VCO_C_0.OUTB.n17 VCO_DFF_C_0.VCO_C_0.OUTB.n14 3.06224
R16888 VCO_DFF_C_0.VCO_C_0.OUTB.n2 VCO_DFF_C_0.VCO_C_0.OUTB.n44 2.82705
R16889 VCO_DFF_C_0.VCO_C_0.OUTB.n11 VCO_DFF_C_0.VCO_C_0.OUTB.n8 2.6005
R16890 VCO_DFF_C_0.VCO_C_0.OUTB.n17 VCO_DFF_C_0.VCO_C_0.OUTB.n16 2.6005
R16891 VCO_DFF_C_0.VCO_C_0.OUTB.n2 VCO_DFF_C_0.VCO_C_0.OUTB 2.36547
R16892 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n56 2.30807
R16893 VCO_DFF_C_0.VCO_C_0.OUTB.n0 VCO_DFF_C_0.VCO_C_0.OUTB.n1 1.10603
R16894 VCO_DFF_C_0.VCO_C_0.OUTB.n56 VCO_DFF_C_0.VCO_C_0.OUTB.n55 2.2505
R16895 VCO_DFF_C_0.VCO_C_0.OUTB.n52 VCO_DFF_C_0.VCO_C_0.OUTB.n48 1.5982
R16896 VCO_DFF_C_0.VCO_C_0.OUTB.n54 VCO_DFF_C_0.VCO_C_0.OUTB.n52 1.18336
R16897 VCO_DFF_C_0.VCO_C_0.OUTB.n55 VCO_DFF_C_0.VCO_C_0.OUTB.n54 0.977746
R16898 VCO_DFF_C_0.VCO_C_0.OUTB.n18 VCO_DFF_C_0.VCO_C_0.OUTB.n12 0.798761
R16899 VCO_DFF_C_0.VCO_C_0.OUTB.n45 VCO_DFF_C_0.VCO_C_0.OUTB.n0 0.66931
R16900 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n22 0.658318
R16901 VCO_DFF_C_0.VCO_C_0.OUTB.n31 VCO_DFF_C_0.VCO_C_0.OUTB 0.637045
R16902 VCO_DFF_C_0.VCO_C_0.OUTB.n25 VCO_DFF_C_0.VCO_C_0.OUTB 0.6125
R16903 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n18 0.562022
R16904 VCO_DFF_C_0.VCO_C_0.OUTB.n32 VCO_DFF_C_0.VCO_C_0.OUTB.n31 0.458758
R16905 VCO_DFF_C_0.VCO_C_0.OUTB.n47 VCO_DFF_C_0.VCO_C_0.OUTB.n46 0.381495
R16906 VCO_DFF_C_0.VCO_C_0.OUTB.n54 VCO_DFF_C_0.VCO_C_0.OUTB.n53 0.37501
R16907 VCO_DFF_C_0.VCO_C_0.OUTB.n48 VCO_DFF_C_0.VCO_C_0.OUTB.n47 0.355126
R16908 VCO_DFF_C_0.VCO_C_0.OUTB.n51 VCO_DFF_C_0.VCO_C_0.OUTB.n50 0.31227
R16909 VCO_DFF_C_0.VCO_C_0.OUTB.n50 VCO_DFF_C_0.VCO_C_0.OUTB.n49 0.298874
R16910 VCO_DFF_C_0.VCO_C_0.OUTB.n56 VCO_DFF_C_0.VCO_C_0.OUTB.n0 0.281082
R16911 VCO_DFF_C_0.VCO_C_0.OUTB.n44 VCO_DFF_C_0.VCO_C_0.OUTB.n32 0.238532
R16912 VCO_DFF_C_0.VCO_C_0.OUTB.n52 VCO_DFF_C_0.VCO_C_0.OUTB.n51 0.233052
R16913 VCO_DFF_C_0.VCO_C_0.OUTB.n12 VCO_DFF_C_0.VCO_C_0.OUTB.n11 0.18637
R16914 VCO_DFF_C_0.VCO_C_0.OUTB.n18 VCO_DFF_C_0.VCO_C_0.OUTB.n17 0.18637
R16915 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB.n1 0.203752
R16916 VCO_DFF_C_0.VCO_C_0.OUTB.n55 VCO_DFF_C_0.VCO_C_0.OUTB.n45 0.137564
R16917 VCO_DFF_C_0.VCO_C_0.OUTB.n44 VCO_DFF_C_0.VCO_C_0.OUTB 0.104622
R16918 VCO_DFF_C_0.VCO_C_0.OUTB.n1 VCO_DFF_C_0.VCO_C_0.OUTB 0.147946
R16919 a_18508_8715.n5 a_18508_8715.t9 29.2961
R16920 a_18508_8715.n6 a_18508_8715.n5 21.9292
R16921 a_18508_8715.n7 a_18508_8715.n6 18.1271
R16922 a_18508_8715.n7 a_18508_8715.t7 11.1695
R16923 a_18508_8715.n3 a_18508_8715.t0 10.2143
R16924 a_18508_8715.n5 a_18508_8715.t8 6.1325
R16925 a_18508_8715.n6 a_18508_8715.t6 6.1325
R16926 a_18508_8715.n3 a_18508_8715.n2 4.68517
R16927 a_18508_8715.n8 a_18508_8715.n7 4.6311
R16928 a_18508_8715.n10 a_18508_8715.n8 2.85093
R16929 a_18508_8715.n1 a_18508_8715.t2 2.16717
R16930 a_18508_8715.n1 a_18508_8715.n0 2.16717
R16931 a_18508_8715.t5 a_18508_8715.n10 2.16717
R16932 a_18508_8715.n10 a_18508_8715.n9 2.16717
R16933 a_18508_8715.n4 a_18508_8715.n3 1.58582
R16934 a_18508_8715.n4 a_18508_8715.n1 1.24371
R16935 a_18508_8715.n8 a_18508_8715.n4 0.971051
R16936 VCO_DFF_C_0.OUT.n4 VCO_DFF_C_0.OUT.t10 37.6513
R16937 VCO_DFF_C_0.OUT VCO_DFF_C_0.OUT.n4 33.1884
R16938 VCO_DFF_C_0.OUT.n1 VCO_DFF_C_0.OUT.t28 32.7094
R16939 VCO_DFF_C_0.OUT VCO_DFF_C_0.OUT.n3 25.211
R16940 VCO_DFF_C_0.OUT.n12 VCO_DFF_C_0.OUT.t24 23.6945
R16941 VCO_DFF_C_0.OUT.t31 VCO_DFF_C_0.OUT.n13 23.6945
R16942 VCO_DFF_C_0.OUT.n23 VCO_DFF_C_0.OUT.t17 23.6945
R16943 VCO_DFF_C_0.OUT.t9 VCO_DFF_C_0.OUT.n24 23.6945
R16944 VCO_DFF_C_0.OUT.n1 VCO_DFF_C_0.OUT.t13 23.2875
R16945 VCO_DFF_C_0.OUT.n2 VCO_DFF_C_0.OUT.t12 23.2875
R16946 VCO_DFF_C_0.OUT.n4 VCO_DFF_C_0.OUT.t26 20.4405
R16947 VCO_DFF_C_0.OUT.n3 VCO_DFF_C_0.OUT.t27 20.4405
R16948 VCO_DFF_C_0.OUT.n13 VCO_DFF_C_0.OUT.n12 18.8035
R16949 VCO_DFF_C_0.OUT.n24 VCO_DFF_C_0.OUT.n23 18.8035
R16950 VCO_DFF_C_0.OUT.n10 VCO_DFF_C_0.OUT.n8 15.8172
R16951 VCO_DFF_C_0.OUT.n9 VCO_DFF_C_0.OUT.n5 15.8172
R16952 VCO_DFF_C_0.OUT.n10 VCO_DFF_C_0.OUT.n9 15.8172
R16953 VCO_DFF_C_0.OUT.n21 VCO_DFF_C_0.OUT.n19 15.8172
R16954 VCO_DFF_C_0.OUT.n21 VCO_DFF_C_0.OUT.n20 15.8172
R16955 VCO_DFF_C_0.OUT.n20 VCO_DFF_C_0.OUT.n16 15.8172
R16956 VCO_DFF_C_0.OUT.n8 VCO_DFF_C_0.OUT.t11 14.8925
R16957 VCO_DFF_C_0.OUT.t19 VCO_DFF_C_0.OUT.n10 14.8925
R16958 VCO_DFF_C_0.OUT.n9 VCO_DFF_C_0.OUT.t35 14.8925
R16959 VCO_DFF_C_0.OUT.n19 VCO_DFF_C_0.OUT.t34 14.8925
R16960 VCO_DFF_C_0.OUT.t18 VCO_DFF_C_0.OUT.n21 14.8925
R16961 VCO_DFF_C_0.OUT.n20 VCO_DFF_C_0.OUT.t32 14.8925
R16962 VCO_DFF_C_0.OUT.n2 VCO_DFF_C_0.OUT.n1 12.5148
R16963 VCO_DFF_C_0.OUT.n14 VCO_DFF_C_0.OUT.n6 12.2457
R16964 VCO_DFF_C_0.OUT.n11 VCO_DFF_C_0.OUT.n6 12.2457
R16965 VCO_DFF_C_0.OUT.n11 VCO_DFF_C_0.OUT.n7 12.2457
R16966 VCO_DFF_C_0.OUT.n25 VCO_DFF_C_0.OUT.n17 12.2457
R16967 VCO_DFF_C_0.OUT.n22 VCO_DFF_C_0.OUT.n17 12.2457
R16968 VCO_DFF_C_0.OUT.n22 VCO_DFF_C_0.OUT.n18 12.2457
R16969 VCO_DFF_C_0.OUT.n3 VCO_DFF_C_0.OUT.n2 12.2081
R16970 VCO_DFF_C_0.OUT.n15 VCO_DFF_C_0.OUT.t20 11.6285
R16971 VCO_DFF_C_0.OUT.n26 VCO_DFF_C_0.OUT.t25 11.6285
R16972 VCO_DFF_C_0.OUT.n7 VCO_DFF_C_0.OUT.t24 8.9065
R16973 VCO_DFF_C_0.OUT.t29 VCO_DFF_C_0.OUT.n11 8.9065
R16974 VCO_DFF_C_0.OUT.t15 VCO_DFF_C_0.OUT.n6 8.9065
R16975 VCO_DFF_C_0.OUT.n14 VCO_DFF_C_0.OUT.t31 8.9065
R16976 VCO_DFF_C_0.OUT.n18 VCO_DFF_C_0.OUT.t17 8.9065
R16977 VCO_DFF_C_0.OUT.t33 VCO_DFF_C_0.OUT.n22 8.9065
R16978 VCO_DFF_C_0.OUT.t16 VCO_DFF_C_0.OUT.n17 8.9065
R16979 VCO_DFF_C_0.OUT.n25 VCO_DFF_C_0.OUT.t9 8.9065
R16980 VCO_DFF_C_0.OUT.n10 VCO_DFF_C_0.OUT.t22 8.6145
R16981 VCO_DFF_C_0.OUT.n8 VCO_DFF_C_0.OUT.t14 8.6145
R16982 VCO_DFF_C_0.OUT.n9 VCO_DFF_C_0.OUT.t8 8.6145
R16983 VCO_DFF_C_0.OUT.n21 VCO_DFF_C_0.OUT.t30 8.6145
R16984 VCO_DFF_C_0.OUT.n19 VCO_DFF_C_0.OUT.t21 8.6145
R16985 VCO_DFF_C_0.OUT.n20 VCO_DFF_C_0.OUT.t6 8.6145
R16986 VCO_DFF_C_0.OUT.n5 VCO_DFF_C_0.OUT.t23 8.59715
R16987 VCO_DFF_C_0.OUT.n16 VCO_DFF_C_0.OUT.t7 8.59715
R16988 VCO_DFF_C_0.OUT.t11 VCO_DFF_C_0.OUT.n7 8.3225
R16989 VCO_DFF_C_0.OUT.n11 VCO_DFF_C_0.OUT.t19 8.3225
R16990 VCO_DFF_C_0.OUT.t35 VCO_DFF_C_0.OUT.n6 8.3225
R16991 VCO_DFF_C_0.OUT.t20 VCO_DFF_C_0.OUT.n14 8.3225
R16992 VCO_DFF_C_0.OUT.t34 VCO_DFF_C_0.OUT.n18 8.3225
R16993 VCO_DFF_C_0.OUT.n22 VCO_DFF_C_0.OUT.t18 8.3225
R16994 VCO_DFF_C_0.OUT.t32 VCO_DFF_C_0.OUT.n17 8.3225
R16995 VCO_DFF_C_0.OUT.t25 VCO_DFF_C_0.OUT.n25 8.3225
R16996 VCO_DFF_C_0.OUT.n0 VCO_DFF_C_0.OUT 4.9636
R16997 VCO_DFF_C_0.OUT VCO_DFF_C_0.OUT.n15 4.223
R16998 VCO_DFF_C_0.OUT VCO_DFF_C_0.OUT.n26 4.223
R16999 VCO_DFF_C_0.OUT.n12 VCO_DFF_C_0.OUT.t29 3.6505
R17000 VCO_DFF_C_0.OUT.n13 VCO_DFF_C_0.OUT.t15 3.6505
R17001 VCO_DFF_C_0.OUT.n23 VCO_DFF_C_0.OUT.t33 3.6505
R17002 VCO_DFF_C_0.OUT.n24 VCO_DFF_C_0.OUT.t16 3.6505
R17003 VCO_DFF_C_0.OUT.n15 VCO_DFF_C_0.OUT.n5 3.1807
R17004 VCO_DFF_C_0.OUT.n26 VCO_DFF_C_0.OUT.n16 3.1807
R17005 VCO_DFF_C_0.OUT.n0 VCO_DFF_C_0.OUT 1.38745
R17006 VCO_DFF_C_0.OUT VCO_DFF_C_0.OUT.n0 0.81407
R17007 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t18 5.81586
R17008 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n23 5.10148
R17009 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n21 5.10116
R17010 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n19 5.08021
R17011 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n25 4.66166
R17012 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t11 3.6405
R17013 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n9 3.6405
R17014 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t12 3.6405
R17015 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n2 3.6405
R17016 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t9 3.6405
R17017 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n4 3.6405
R17018 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t15 3.6405
R17019 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n11 3.6405
R17020 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n8 3.50463
R17021 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n1 3.50463
R17022 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t6 3.2765
R17023 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n7 3.2765
R17024 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t4 3.2765
R17025 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n0 3.2765
R17026 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n5 3.06224
R17027 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n12 3.06224
R17028 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n17 2.85093
R17029 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n3 2.6005
R17030 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n10 2.6005
R17031 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n27 2.36593
R17032 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t17 2.16717
R17033 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n16 2.16717
R17034 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.t1 1.9505
R17035 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n24 1.9505
R17036 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n14 0.798761
R17037 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n18 0.644196
R17038 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n15 0.562022
R17039 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n20 0.450839
R17040 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n26 0.358498
R17041 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n22 0.229792
R17042 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n6 0.18637
R17043 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN.n13 0.18637
R17044 a_43828_11254.t0 a_43828_11254.t1 12.9675
R17045 a_43528_10632.t0 a_43528_10632.t1 12.9675
R17046 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t57 23.6945
R17047 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t40 23.6945
R17048 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n30 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n29 18.8035
R17049 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n24 15.8172
R17050 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n24 15.8172
R17051 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n32 15.8172
R17052 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t41 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n27 14.8925
R17053 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t45 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n24 14.8925
R17054 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t49 14.8925
R17055 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n25 12.2457
R17056 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n26 12.2457
R17057 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n28 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n26 12.2457
R17058 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t43 11.6285
R17059 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t51 9.57577
R17060 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t54 9.55796
R17061 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n66 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t10 9.31704
R17062 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n44 8.94165
R17063 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t57 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n28 8.9065
R17064 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t52 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n26 8.9065
R17065 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n31 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t33 8.9065
R17066 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t40 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n25 8.9065
R17067 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n27 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t32 8.6145
R17068 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t37 8.6145
R17069 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n32 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t44 8.6145
R17070 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n33 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t34 8.59715
R17071 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n10 8.59228
R17072 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n37 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t31 8.56851
R17073 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t39 8.56851
R17074 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t38 8.56851
R17075 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t42 8.5214
R17076 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t35 8.5214
R17077 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t56 8.5214
R17078 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t58 8.5214
R17079 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n42 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t47 8.5112
R17080 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t48 8.5112
R17081 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n40 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t36 8.5112
R17082 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t53 8.34992
R17083 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n28 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t41 8.3225
R17084 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t45 8.3225
R17085 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t49 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n31 8.3225
R17086 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t43 8.3225
R17087 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n72 8.65114
R17088 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t50 8.30779
R17089 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t46 8.30779
R17090 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t55 8.30779
R17091 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n64 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n62 7.40037
R17092 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t26 7.05758
R17093 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n21 6.80072
R17094 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n11 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n9 6.73941
R17095 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t18 6.45366
R17096 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t22 6.2092
R17097 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n15 5.83551
R17098 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n45 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t12 4.89657
R17099 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n64 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n63 4.88218
R17100 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n70 4.87529
R17101 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t11 4.6632
R17102 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t4 4.63112
R17103 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n48 5.42442
R17104 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n58 4.54362
R17105 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n34 4.223
R17106 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n61 4.01867
R17107 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n8 3.9838
R17108 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n36 3.96161
R17109 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n65 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n64 3.87403
R17110 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n29 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t52 3.6505
R17111 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t33 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n30 3.6505
R17112 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t3 3.6405
R17113 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n48 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n47 3.6405
R17114 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t17 3.6405
R17115 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n7 3.6405
R17116 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n58 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t8 3.6405
R17117 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n58 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n57 3.6405
R17118 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n60 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t9 3.6405
R17119 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n60 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n59 3.6405
R17120 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t1 3.6405
R17121 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n52 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n51 3.6405
R17122 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t30 3.47629
R17123 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t29 3.47625
R17124 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.t27 3.47617
R17125 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n14 3.39849
R17126 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n34 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n33 3.1807
R17127 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n19 2.86157
R17128 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n13 2.8615
R17129 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n17 2.86147
R17130 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n18 2.48336
R17131 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n20 2.47781
R17132 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 2.35499
R17133 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 2.30073
R17134 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n5 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n54 2.24532
R17135 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n52 4.81789
R17136 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n54 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n53 2.21522
R17137 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n49 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n46 1.7262
R17138 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n43 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n42 1.61187
R17139 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n43 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n39 1.57365
R17140 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n56 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n55 1.51564
R17141 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n35 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 1.51518
R17142 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n46 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n45 1.49463
R17143 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n71 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n12 1.36952
R17144 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n61 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n60 1.25753
R17145 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n2 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n3 1.05601
R17146 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n22 1.01067
R17147 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n41 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n40 0.996664
R17148 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n0 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n4 0.992966
R17149 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n16 0.983287
R17150 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n0 0.975705
R17151 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n56 0.969569
R17152 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n70 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n69 0.955885
R17153 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n38 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n37 0.953514
R17154 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n2 0.907492
R17155 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n66 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n65 0.856289
R17156 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n68 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n67 0.843096
R17157 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n53 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n50 0.8015
R17158 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n11 0.800717
R17159 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n55 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n5 0.741058
R17160 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n56 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n6 0.69855
R17161 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n69 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n68 0.656716
R17162 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n67 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n66 0.398395
R17163 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n50 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n49 0.3875
R17164 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n39 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n38 0.364199
R17165 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n23 0.362368
R17166 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n1 0.359267
R17167 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n42 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n41 0.323514
R17168 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n43 0.319815
R17169 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n36 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n35 0.193979
R17170 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN.n71 0.147028
R17171 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t18 23.6945
R17172 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t22 23.6945
R17173 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n7 18.8035
R17174 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n2 15.8172
R17175 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n11 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n10 15.8172
R17176 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n2 15.8172
R17177 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n5 14.8925
R17178 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n2 14.8925
R17179 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t23 14.8925
R17180 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n3 12.2457
R17181 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n4 12.2457
R17182 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n4 12.2457
R17183 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t19 11.6285
R17184 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n6 8.9065
R17185 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n4 8.9065
R17186 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t17 8.9065
R17187 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n3 8.9065
R17188 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t16 8.6145
R17189 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n2 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t26 8.6145
R17190 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t24 8.6145
R17191 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n11 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t20 8.59715
R17192 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t27 8.3225
R17193 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n4 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t25 8.3225
R17194 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n9 8.3225
R17195 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t19 8.3225
R17196 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t13 6.74566
R17197 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n0 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t4 6.74332
R17198 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n0 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t2 5.1005
R17199 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t12 5.1005
R17200 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n12 4.223
R17201 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t21 3.6505
R17202 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n8 3.6505
R17203 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n16 3.57508
R17204 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n27 3.5743
R17205 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n0 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n13 3.40011
R17206 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n22 3.40001
R17207 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n11 3.1807
R17208 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t11 3.00159
R17209 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t5 3.00158
R17210 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n20 2.58112
R17211 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n29 2.58112
R17212 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t15 2.16717
R17213 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n17 2.16717
R17214 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t8 2.16717
R17215 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n15 2.16717
R17216 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t7 2.16717
R17217 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n24 2.16717
R17218 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.t0 2.16717
R17219 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n26 2.16717
R17220 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n14 1.84821
R17221 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n29 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n23 1.84725
R17222 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n18 1.25233
R17223 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n25 1.25225
R17224 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n29 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n28 1.12575
R17225 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n19 1.12554
R17226 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n21 0.784521
R17227 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.689881
R17228 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n1 0.55941
R17229 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n0 0.558372
R17230 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.25925
R17231 a_22879_10704.n1 a_22879_10704.t2 7.58276
R17232 a_22879_10704.n3 a_22879_10704.n1 7.16556
R17233 a_22879_10704.n1 a_22879_10704.n0 6.4265
R17234 a_22879_10704.n3 a_22879_10704.n2 3.4179
R17235 a_22879_10704.t1 a_22879_10704.n3 2.93981
R17236 UP_OUT.n25 UP_OUT.n24 14.6005
R17237 UP_OUT.n27 UP_OUT.n26 12.8446
R17238 UP_OUT.n1 UP_OUT.t10 6.74332
R17239 UP_OUT.n17 UP_OUT.n16 6.74326
R17240 UP_OUT.n24 UP_OUT.t18 6.51836
R17241 UP_OUT.n24 UP_OUT.t17 6.51836
R17242 UP_OUT.n25 UP_OUT.t20 6.51836
R17243 UP_OUT.n27 UP_OUT.t19 6.388
R17244 UP_OUT.n26 UP_OUT.t16 6.19246
R17245 UP_OUT.n29 UP_OUT 5.62004
R17246 UP_OUT.n19 UP_OUT.n18 5.1005
R17247 UP_OUT.n2 UP_OUT.t11 5.1005
R17248 UP_OUT.n28 UP_OUT.n27 5.01216
R17249 UP_OUT.n14 UP_OUT.n13 3.5743
R17250 UP_OUT.n8 UP_OUT.n7 3.5743
R17251 UP_OUT.n17 UP_OUT.t3 3.40065
R17252 UP_OUT.n1 UP_OUT.n0 3.40001
R17253 UP_OUT.n3 UP_OUT.t9 3.00159
R17254 UP_OUT.n20 UP_OUT.n15 3.00034
R17255 UP_OUT.n23 UP_OUT 2.61054
R17256 UP_OUT.n23 UP_OUT.n22 2.30818
R17257 UP_OUT.n11 UP_OUT.t6 2.16717
R17258 UP_OUT.n11 UP_OUT.n10 2.16717
R17259 UP_OUT.n13 UP_OUT.t5 2.16717
R17260 UP_OUT.n13 UP_OUT.n12 2.16717
R17261 UP_OUT.n5 UP_OUT.t13 2.16717
R17262 UP_OUT.n5 UP_OUT.n4 2.16717
R17263 UP_OUT.n7 UP_OUT.t14 2.16717
R17264 UP_OUT.n7 UP_OUT.n6 2.16717
R17265 UP_OUT.n30 UP_OUT.n23 1.86359
R17266 UP_OUT.n9 UP_OUT.n3 1.84725
R17267 UP_OUT.n21 UP_OUT.n20 1.847
R17268 UP_OUT.n14 UP_OUT.n11 1.25225
R17269 UP_OUT.n8 UP_OUT.n5 1.25225
R17270 UP_OUT.n28 UP_OUT 1.19735
R17271 UP_OUT.n21 UP_OUT.n14 1.12594
R17272 UP_OUT.n9 UP_OUT.n8 1.12575
R17273 UP_OUT UP_OUT.n31 0.751569
R17274 UP_OUT.n22 UP_OUT 0.736693
R17275 UP_OUT.n20 UP_OUT.n19 0.447297
R17276 UP_OUT.n3 UP_OUT.n2 0.446651
R17277 UP_OUT.n30 UP_OUT.n29 0.412666
R17278 UP_OUT.n22 UP_OUT.n21 0.378912
R17279 UP_OUT.n31 UP_OUT.n30 0.353294
R17280 UP_OUT.n31 UP_OUT.n9 0.339608
R17281 UP_OUT.n26 UP_OUT.n25 0.326393
R17282 UP_OUT.n29 UP_OUT.n28 0.151125
R17283 UP_OUT.n2 UP_OUT.n1 0.11326
R17284 UP_OUT.n19 UP_OUT.n17 0.112615
R17285 a_32939_9624.n7 a_32939_9624.n6 10.1602
R17286 a_32939_9624.n1 a_32939_9624.n0 5.4005
R17287 a_32939_9624.n1 a_32939_9624.t0 5.4005
R17288 a_32939_9624.n5 a_32939_9624.n4 5.4005
R17289 a_32939_9624.n5 a_32939_9624.t5 5.4005
R17290 a_32939_9624.n3 a_32939_9624.n2 5.4005
R17291 a_32939_9624.n3 a_32939_9624.t6 5.4005
R17292 a_32939_9624.n11 a_32939_9624.n10 5.4005
R17293 a_32939_9624.t4 a_32939_9624.n11 5.4005
R17294 a_32939_9624.n11 a_32939_9624.n9 3.51269
R17295 a_32939_9624.n8 a_32939_9624.n3 3.31203
R17296 a_32939_9624.n7 a_32939_9624.n5 3.28072
R17297 a_32939_9624.n9 a_32939_9624.n1 3.1505
R17298 a_32939_9624.n8 a_32939_9624.n7 1.46985
R17299 a_32939_9624.n9 a_32939_9624.n8 1.03855
R17300 PFD_T2_0.INV_mag_0.OUT.n4 PFD_T2_0.INV_mag_0.OUT.n3 34.5741
R17301 PFD_T2_0.INV_mag_0.OUT.n3 PFD_T2_0.INV_mag_0.OUT.t8 33.8279
R17302 PFD_T2_0.INV_mag_0.OUT.n0 PFD_T2_0.INV_mag_0.OUT.t3 30.6524
R17303 PFD_T2_0.INV_mag_0.OUT.n1 PFD_T2_0.INV_mag_0.OUT.t4 30.6524
R17304 PFD_T2_0.INV_mag_0.OUT.n0 PFD_T2_0.INV_mag_0.OUT.t7 9.5635
R17305 PFD_T2_0.INV_mag_0.OUT.n1 PFD_T2_0.INV_mag_0.OUT.t5 9.5635
R17306 PFD_T2_0.INV_mag_0.OUT.n5 PFD_T2_0.INV_mag_0.OUT.n4 9.26523
R17307 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.OUT.n6 6.74425
R17308 PFD_T2_0.INV_mag_0.OUT.n4 PFD_T2_0.INV_mag_0.OUT.t9 6.5705
R17309 PFD_T2_0.INV_mag_0.OUT.n2 PFD_T2_0.INV_mag_0.OUT.n0 5.32623
R17310 PFD_T2_0.INV_mag_0.OUT.n2 PFD_T2_0.INV_mag_0.OUT.n1 4.78052
R17311 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.OUT.n5 4.4032
R17312 PFD_T2_0.INV_mag_0.OUT.n3 PFD_T2_0.INV_mag_0.OUT.t6 3.6505
R17313 PFD_T2_0.INV_mag_0.OUT.n8 PFD_T2_0.INV_mag_0.OUT.t1 3.6405
R17314 PFD_T2_0.INV_mag_0.OUT.n8 PFD_T2_0.INV_mag_0.OUT.n7 3.6405
R17315 PFD_T2_0.INV_mag_0.OUT.n5 PFD_T2_0.INV_mag_0.OUT.n2 3.38996
R17316 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.INV_mag_0.OUT.n8 3.35938
R17317 a_22966_11778.n4 a_22966_11778.t11 33.8126
R17318 a_22966_11778.n5 a_22966_11778.n4 30.3299
R17319 a_22966_11778.n6 a_22966_11778.n5 30.3299
R17320 a_22966_11778.n7 a_22966_11778.n6 30.3299
R17321 a_22966_11778.n8 a_22966_11778.n7 30.3299
R17322 a_22966_11778.n9 a_22966_11778.n8 30.3299
R17323 a_22966_11778.n10 a_22966_11778.n9 30.3299
R17324 a_22966_11778.n11 a_22966_11778.n10 30.3299
R17325 a_22966_11778.n12 a_22966_11778.n11 30.3299
R17326 a_22966_11778.n0 a_22966_11778.t14 26.2932
R17327 a_22966_11778.n13 a_22966_11778.t9 12.8368
R17328 a_22966_11778.n13 a_22966_11778.n12 12.0257
R17329 a_22966_11778.n3 a_22966_11778.n0 8.47283
R17330 a_22966_11778.n14 a_22966_11778.n13 5.21535
R17331 a_22966_11778.n0 a_22966_11778.t5 3.6505
R17332 a_22966_11778.n4 a_22966_11778.t4 3.6505
R17333 a_22966_11778.n5 a_22966_11778.t10 3.6505
R17334 a_22966_11778.n6 a_22966_11778.t15 3.6505
R17335 a_22966_11778.n7 a_22966_11778.t6 3.6505
R17336 a_22966_11778.n8 a_22966_11778.t16 3.6505
R17337 a_22966_11778.n9 a_22966_11778.t7 3.6505
R17338 a_22966_11778.n10 a_22966_11778.t12 3.6505
R17339 a_22966_11778.n11 a_22966_11778.t8 3.6505
R17340 a_22966_11778.n12 a_22966_11778.t13 3.6505
R17341 a_22966_11778.n15 a_22966_11778.t2 3.6405
R17342 a_22966_11778.n16 a_22966_11778.n15 3.6405
R17343 a_22966_11778.n14 a_22966_11778.n3 3.5048
R17344 a_22966_11778.n2 a_22966_11778.t0 3.38775
R17345 a_22966_11778.n2 a_22966_11778.n1 2.97655
R17346 a_22966_11778.n3 a_22966_11778.n2 2.47443
R17347 a_22966_11778.n15 a_22966_11778.n14 1.25594
R17348 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t13 14.1829
R17349 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t12 13.9657
R17350 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t20 13.3574
R17351 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t17 13.1401
R17352 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n1 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t14 12.9025
R17353 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t16 12.6187
R17354 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t21 8.77788
R17355 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t19 8.64752
R17356 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n5 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t15 8.56062
R17357 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n4 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t18 8.43026
R17358 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n6 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n5 6.11825
R17359 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n6 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n4 5.88354
R17360 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n11 4.64372
R17361 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t8 3.6405
R17362 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n22 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n21 3.6405
R17363 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t6 3.6405
R17364 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n14 3.6405
R17365 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n17 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t5 3.6405
R17366 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n17 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n16 3.6405
R17367 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n24 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t7 3.6405
R17368 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n24 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n23 3.6405
R17369 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n20 3.50463
R17370 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n13 3.50463
R17371 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t2 3.2765
R17372 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n20 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n19 3.2765
R17373 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n13 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.t1 3.2765
R17374 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n13 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n12 3.2765
R17375 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n18 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n17 3.06224
R17376 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n24 3.06224
R17377 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n18 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n15 2.6005
R17378 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n25 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n22 2.6005
R17379 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT 2.32194
R17380 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n0 2.31638
R17381 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n0 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n10 2.2505
R17382 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n8 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n7 1.58291
R17383 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n3 1.47586
R17384 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n10 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n9 1.33917
R17385 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n9 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n8 1.23958
R17386 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n26 0.798761
R17387 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n27 0.562022
R17388 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n7 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n6 0.448735
R17389 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n3 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n2 0.386992
R17390 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n2 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n1 0.340685
R17391 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n27 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n18 0.18637
R17392 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n26 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n25 0.18637
R17393 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n11 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT.n0 0.130397
R17394 UP1.n14 UP1.n13 6.76498
R17395 UP1.n3 UP1.n2 5.81586
R17396 UP1.n8 UP1.t3 5.10151
R17397 UP1.n5 UP1.t1 5.1005
R17398 UP1.n4 UP1.t7 5.08021
R17399 UP1.n8 UP1.n7 4.66164
R17400 UP1.n12 UP1.t10 3.6405
R17401 UP1.n12 UP1.n11 3.6405
R17402 UP1.n3 UP1.n1 2.85093
R17403 UP1.n14 UP1.n12 2.78441
R17404 UP1.n15 UP1 2.26578
R17405 UP1.n1 UP1.t4 2.16717
R17406 UP1.n1 UP1.n0 2.16717
R17407 UP1.n7 UP1.t0 1.9505
R17408 UP1.n7 UP1.n6 1.9505
R17409 UP1.n10 UP1 1.3114
R17410 UP1.n10 UP1 1.04229
R17411 UP1.n4 UP1.n3 0.644196
R17412 UP1.n5 UP1.n4 0.447229
R17413 UP1 UP1.n14 0.428459
R17414 UP1 UP1.n10 0.375783
R17415 UP1.n9 UP1.n8 0.254356
R17416 UP1.n9 UP1.n5 0.22163
R17417 UP1 UP1.n9 0.127741
R17418 UP1.n15 UP1 0.12599
R17419 UP1 UP1.n15 0.0125
R17420 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t23 45.6363
R17421 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t30 45.6363
R17422 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t15 29.6446
R17423 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n18 29.6446
R17424 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t20 29.6446
R17425 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n20 29.6446
R17426 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t21 24.6117
R17427 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t28 24.6117
R17428 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n17 22.2047
R17429 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n19 22.2047
R17430 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t29 22.1925
R17431 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t30 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t18 22.1925
R17432 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t16 21.8613
R17433 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n26 20.9314
R17434 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n22 20.9314
R17435 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t19 17.8613
R17436 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n28 10.8592
R17437 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n25 8.94379
R17438 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n16 8.87094
R17439 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n26 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t27 6.1325
R17440 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n27 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t25 6.1325
R17441 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n17 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t31 6.1325
R17442 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n18 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t14 6.1325
R17443 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n16 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t13 6.1325
R17444 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n19 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t17 6.1325
R17445 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n20 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t22 6.1325
R17446 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n21 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t12 6.1325
R17447 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n22 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t24 6.1325
R17448 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n23 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t26 6.1325
R17449 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n23 5.38991
R17450 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n27 5.12094
R17451 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n24 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n21 4.83094
R17452 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t7 3.6405
R17453 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n10 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n9 3.6405
R17454 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t9 3.6405
R17455 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n3 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n2 3.6405
R17456 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t5 3.6405
R17457 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n5 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n4 3.6405
R17458 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t11 3.6405
R17459 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n12 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n11 3.6405
R17460 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n8 3.50463
R17461 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n1 3.50463
R17462 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t1 3.2765
R17463 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n8 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n7 3.2765
R17464 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.t2 3.2765
R17465 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n1 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n0 3.2765
R17466 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n5 3.06224
R17467 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n12 3.06224
R17468 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n6 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n3 2.6005
R17469 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n13 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n10 2.6005
R17470 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n28 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 1.07267
R17471 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n14 0.798761
R17472 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n24 0.658318
R17473 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n25 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 0.628846
R17474 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n15 0.562022
R17475 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n15 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n6 0.18637
R17476 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n14 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK.n13 0.18637
R17477 a_44716_n517.n0 a_44716_n517.t6 29.2961
R17478 a_44716_n517.n1 a_44716_n517.n0 21.9292
R17479 a_44716_n517.n2 a_44716_n517.n1 18.1271
R17480 a_44716_n517.n2 a_44716_n517.t7 11.1695
R17481 a_44716_n517.n0 a_44716_n517.t8 6.1325
R17482 a_44716_n517.n1 a_44716_n517.t9 6.1325
R17483 a_44716_n517.n6 a_44716_n517.n5 4.93252
R17484 a_44716_n517.n6 a_44716_n517.t1 4.70348
R17485 a_44716_n517.n8 a_44716_n517.n2 4.6311
R17486 a_44716_n517.n9 a_44716_n517.n8 2.85093
R17487 a_44716_n517.n4 a_44716_n517.t2 2.16717
R17488 a_44716_n517.n4 a_44716_n517.n3 2.16717
R17489 a_44716_n517.n9 a_44716_n517.t3 2.16717
R17490 a_44716_n517.n10 a_44716_n517.n9 2.16717
R17491 a_44716_n517.n7 a_44716_n517.n6 1.58582
R17492 a_44716_n517.n7 a_44716_n517.n4 1.24371
R17493 a_44716_n517.n8 a_44716_n517.n7 0.971051
R17494 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t16 23.6945
R17495 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t22 23.6945
R17496 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n22 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n21 18.8035
R17497 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n16 15.8172
R17498 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n16 15.8172
R17499 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n24 15.8172
R17500 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t18 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n19 14.8925
R17501 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t20 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n16 14.8925
R17502 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t23 14.8925
R17503 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n17 12.2457
R17504 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n18 12.2457
R17505 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n18 12.2457
R17506 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t13 11.6285
R17507 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t16 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n20 8.9065
R17508 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t17 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n18 8.9065
R17509 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n23 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t15 8.9065
R17510 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t22 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n17 8.9065
R17511 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n19 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t19 8.6145
R17512 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n16 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t21 8.6145
R17513 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n24 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t12 8.6145
R17514 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n25 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t14 8.59715
R17515 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n20 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t18 8.3225
R17516 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n18 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t20 8.3225
R17517 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t23 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n23 8.3225
R17518 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n17 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t13 8.3225
R17519 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n26 4.223
R17520 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n21 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t17 3.6505
R17521 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t15 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n22 3.6505
R17522 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t8 3.6405
R17523 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n12 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n11 3.6405
R17524 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t5 3.6405
R17525 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n1 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n0 3.6405
R17526 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t7 3.6405
R17527 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n3 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n2 3.6405
R17528 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t10 3.6405
R17529 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n10 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n9 3.6405
R17530 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n8 3.50463
R17531 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n6 3.50463
R17532 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t2 3.2765
R17533 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n8 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n7 3.2765
R17534 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.t1 3.2765
R17535 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n6 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n5 3.2765
R17536 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n26 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n25 3.1807
R17537 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n1 3.06224
R17538 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n10 3.06224
R17539 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n4 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n3 2.6005
R17540 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n13 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n12 2.6005
R17541 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n14 0.798761
R17542 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n15 0.562022
R17543 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n15 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n4 0.18637
R17544 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n14 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN.n13 0.18637
R17545 VCO_DFF_C_0.VCO_C_0.OUT.n24 VCO_DFF_C_0.VCO_C_0.OUT.t14 14.1829
R17546 VCO_DFF_C_0.VCO_C_0.OUT.n23 VCO_DFF_C_0.VCO_C_0.OUT.t21 13.9657
R17547 VCO_DFF_C_0.VCO_C_0.OUT.n17 VCO_DFF_C_0.VCO_C_0.OUT.t18 13.3574
R17548 VCO_DFF_C_0.VCO_C_0.OUT.n16 VCO_DFF_C_0.VCO_C_0.OUT.t15 13.1401
R17549 VCO_DFF_C_0.VCO_C_0.OUT.n16 VCO_DFF_C_0.VCO_C_0.OUT.t16 12.9025
R17550 VCO_DFF_C_0.VCO_C_0.OUT.n18 VCO_DFF_C_0.VCO_C_0.OUT.t17 12.6187
R17551 VCO_DFF_C_0.VCO_C_0.OUT.n20 VCO_DFF_C_0.VCO_C_0.OUT.t20 8.77788
R17552 VCO_DFF_C_0.VCO_C_0.OUT.n19 VCO_DFF_C_0.VCO_C_0.OUT.t12 8.64752
R17553 VCO_DFF_C_0.VCO_C_0.OUT.n19 VCO_DFF_C_0.VCO_C_0.OUT.t19 8.56062
R17554 VCO_DFF_C_0.VCO_C_0.OUT.n20 VCO_DFF_C_0.VCO_C_0.OUT.t13 8.43026
R17555 VCO_DFF_C_0.VCO_C_0.OUT.n21 VCO_DFF_C_0.VCO_C_0.OUT.n19 6.11825
R17556 VCO_DFF_C_0.VCO_C_0.OUT.n21 VCO_DFF_C_0.VCO_C_0.OUT.n20 5.88354
R17557 VCO_DFF_C_0.VCO_C_0.OUT.n10 VCO_DFF_C_0.VCO_C_0.OUT.t5 3.6405
R17558 VCO_DFF_C_0.VCO_C_0.OUT.n10 VCO_DFF_C_0.VCO_C_0.OUT.n9 3.6405
R17559 VCO_DFF_C_0.VCO_C_0.OUT.n3 VCO_DFF_C_0.VCO_C_0.OUT.t6 3.6405
R17560 VCO_DFF_C_0.VCO_C_0.OUT.n3 VCO_DFF_C_0.VCO_C_0.OUT.n2 3.6405
R17561 VCO_DFF_C_0.VCO_C_0.OUT.n1 VCO_DFF_C_0.VCO_C_0.OUT.t8 3.6405
R17562 VCO_DFF_C_0.VCO_C_0.OUT.n1 VCO_DFF_C_0.VCO_C_0.OUT.n0 3.6405
R17563 VCO_DFF_C_0.VCO_C_0.OUT.n12 VCO_DFF_C_0.VCO_C_0.OUT.t11 3.6405
R17564 VCO_DFF_C_0.VCO_C_0.OUT.n12 VCO_DFF_C_0.VCO_C_0.OUT.n11 3.6405
R17565 VCO_DFF_C_0.VCO_C_0.OUT.n14 VCO_DFF_C_0.VCO_C_0.OUT.n8 3.50463
R17566 VCO_DFF_C_0.VCO_C_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.OUT.n6 3.50463
R17567 VCO_DFF_C_0.VCO_C_0.OUT.n8 VCO_DFF_C_0.VCO_C_0.OUT.t2 3.2765
R17568 VCO_DFF_C_0.VCO_C_0.OUT.n8 VCO_DFF_C_0.VCO_C_0.OUT.n7 3.2765
R17569 VCO_DFF_C_0.VCO_C_0.OUT.n6 VCO_DFF_C_0.VCO_C_0.OUT.t0 3.2765
R17570 VCO_DFF_C_0.VCO_C_0.OUT.n6 VCO_DFF_C_0.VCO_C_0.OUT.n5 3.2765
R17571 VCO_DFF_C_0.VCO_C_0.OUT.n4 VCO_DFF_C_0.VCO_C_0.OUT.n1 3.06224
R17572 VCO_DFF_C_0.VCO_C_0.OUT.n13 VCO_DFF_C_0.VCO_C_0.OUT.n10 3.06224
R17573 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.OUT.n24 2.91964
R17574 VCO_DFF_C_0.VCO_C_0.OUT.n4 VCO_DFF_C_0.VCO_C_0.OUT.n3 2.6005
R17575 VCO_DFF_C_0.VCO_C_0.OUT.n13 VCO_DFF_C_0.VCO_C_0.OUT.n12 2.6005
R17576 VCO_DFF_C_0.VCO_C_0.OUT.n23 VCO_DFF_C_0.VCO_C_0.OUT.n22 1.58291
R17577 VCO_DFF_C_0.VCO_C_0.OUT.n22 VCO_DFF_C_0.VCO_C_0.OUT.n18 1.47586
R17578 VCO_DFF_C_0.VCO_C_0.OUT.n24 VCO_DFF_C_0.VCO_C_0.OUT.n23 1.23958
R17579 VCO_DFF_C_0.VCO_C_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.OUT.n14 0.798761
R17580 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.OUT.n15 0.561439
R17581 VCO_DFF_C_0.VCO_C_0.OUT.n22 VCO_DFF_C_0.VCO_C_0.OUT.n21 0.448735
R17582 VCO_DFF_C_0.VCO_C_0.OUT.n18 VCO_DFF_C_0.VCO_C_0.OUT.n17 0.386992
R17583 VCO_DFF_C_0.VCO_C_0.OUT.n17 VCO_DFF_C_0.VCO_C_0.OUT.n16 0.340685
R17584 VCO_DFF_C_0.VCO_C_0.OUT.n15 VCO_DFF_C_0.VCO_C_0.OUT.n4 0.18637
R17585 VCO_DFF_C_0.VCO_C_0.OUT.n14 VCO_DFF_C_0.VCO_C_0.OUT.n13 0.18637
R17586 a_22880_9797.t1 a_22880_9797.n3 7.58276
R17587 a_22880_9797.n3 a_22880_9797.n1 7.1657
R17588 a_22880_9797.n3 a_22880_9797.n2 6.4265
R17589 a_22880_9797.n1 a_22880_9797.n0 3.41789
R17590 a_22880_9797.n1 a_22880_9797.t2 2.93982
R17591 DN_OUT.t18 DN_OUT.t20 12.5148
R17592 DN_OUT.n3 DN_OUT.t18 10.215
R17593 DN_OUT.n0 DN_OUT.t21 10.1117
R17594 DN_OUT.n1 DN_OUT.t17 9.54068
R17595 DN_OUT.n2 DN_OUT.t16 9.4755
R17596 DN_OUT.n0 DN_OUT.t19 9.4755
R17597 DN_OUT.n6 DN_OUT.t4 6.74332
R17598 DN_OUT.n23 DN_OUT.n22 6.74326
R17599 DN_OUT.n4 DN_OUT 6.06505
R17600 DN_OUT.n7 DN_OUT.t5 5.1005
R17601 DN_OUT.n25 DN_OUT.n24 5.1005
R17602 DN_OUT DN_OUT.n4 4.78785
R17603 DN_OUT.n13 DN_OUT.n12 3.5743
R17604 DN_OUT.n20 DN_OUT.n19 3.5743
R17605 DN_OUT.n23 DN_OUT.t15 3.40065
R17606 DN_OUT.n6 DN_OUT.n5 3.40001
R17607 DN_OUT.n8 DN_OUT.t10 3.00159
R17608 DN_OUT.n26 DN_OUT.n21 3.00034
R17609 DN_OUT DN_OUT.n29 2.57784
R17610 DN_OUT.n29 DN_OUT.n15 2.36206
R17611 DN_OUT.n29 DN_OUT.n28 2.30818
R17612 DN_OUT.n10 DN_OUT.t12 2.16717
R17613 DN_OUT.n10 DN_OUT.n9 2.16717
R17614 DN_OUT.n12 DN_OUT.t0 2.16717
R17615 DN_OUT.n12 DN_OUT.n11 2.16717
R17616 DN_OUT.n17 DN_OUT.t1 2.16717
R17617 DN_OUT.n17 DN_OUT.n16 2.16717
R17618 DN_OUT.n19 DN_OUT.t6 2.16717
R17619 DN_OUT.n19 DN_OUT.n18 2.16717
R17620 DN_OUT.n14 DN_OUT.n8 1.84725
R17621 DN_OUT.n27 DN_OUT.n26 1.847
R17622 DN_OUT.n13 DN_OUT.n10 1.25225
R17623 DN_OUT.n20 DN_OUT.n17 1.25225
R17624 DN_OUT.n27 DN_OUT.n20 1.12594
R17625 DN_OUT.n14 DN_OUT.n13 1.12575
R17626 DN_OUT.n15 DN_OUT 0.751569
R17627 DN_OUT.n28 DN_OUT 0.736693
R17628 DN_OUT.n2 DN_OUT.n1 0.50481
R17629 DN_OUT.n1 DN_OUT.n0 0.501707
R17630 DN_OUT.n4 DN_OUT 0.498
R17631 DN_OUT.n26 DN_OUT.n25 0.447297
R17632 DN_OUT.n8 DN_OUT.n7 0.446651
R17633 DN_OUT.n3 DN_OUT.n2 0.393086
R17634 DN_OUT.n28 DN_OUT.n27 0.378912
R17635 DN_OUT.n15 DN_OUT.n14 0.339608
R17636 DN_OUT DN_OUT.n3 0.200095
R17637 DN_OUT.n7 DN_OUT.n6 0.11326
R17638 DN_OUT.n25 DN_OUT.n23 0.112615
R17639 A_MUX_4.Tr_Gate_1.CLK.n14 A_MUX_4.Tr_Gate_1.CLK.t19 45.6363
R17640 A_MUX_4.Tr_Gate_1.CLK.n16 A_MUX_4.Tr_Gate_1.CLK.t13 29.6446
R17641 A_MUX_4.Tr_Gate_1.CLK.t15 A_MUX_4.Tr_Gate_1.CLK.n17 29.6446
R17642 A_MUX_4.Tr_Gate_1.CLK.n18 A_MUX_4.Tr_Gate_1.CLK.t16 24.6117
R17643 A_MUX_4.Tr_Gate_1.CLK.n17 A_MUX_4.Tr_Gate_1.CLK.n16 22.2047
R17644 A_MUX_4.Tr_Gate_1.CLK.t19 A_MUX_4.Tr_Gate_1.CLK.t14 22.1925
R17645 A_MUX_4.Tr_Gate_1.CLK.n15 A_MUX_4.Tr_Gate_1.CLK.n14 20.9314
R17646 A_MUX_4.Tr_Gate_1.CLK A_MUX_4.Tr_Gate_1.CLK.t15 18.524
R17647 A_MUX_4.Tr_Gate_1.CLK.n18 A_MUX_4.Tr_Gate_1.CLK.t12 6.1325
R17648 A_MUX_4.Tr_Gate_1.CLK.n16 A_MUX_4.Tr_Gate_1.CLK.t20 6.1325
R17649 A_MUX_4.Tr_Gate_1.CLK.n17 A_MUX_4.Tr_Gate_1.CLK.t17 6.1325
R17650 A_MUX_4.Tr_Gate_1.CLK.n14 A_MUX_4.Tr_Gate_1.CLK.t21 6.1325
R17651 A_MUX_4.Tr_Gate_1.CLK.n15 A_MUX_4.Tr_Gate_1.CLK.t18 6.1325
R17652 A_MUX_4.Tr_Gate_1.CLK A_MUX_4.Tr_Gate_1.CLK.n15 5.28289
R17653 A_MUX_4.Tr_Gate_1.CLK A_MUX_4.Tr_Gate_1.CLK.n18 4.89628
R17654 A_MUX_4.Tr_Gate_1.CLK.n11 A_MUX_4.Tr_Gate_1.CLK.t7 3.6405
R17655 A_MUX_4.Tr_Gate_1.CLK.n11 A_MUX_4.Tr_Gate_1.CLK.n10 3.6405
R17656 A_MUX_4.Tr_Gate_1.CLK.n7 A_MUX_4.Tr_Gate_1.CLK.t8 3.6405
R17657 A_MUX_4.Tr_Gate_1.CLK.n7 A_MUX_4.Tr_Gate_1.CLK.n6 3.6405
R17658 A_MUX_4.Tr_Gate_1.CLK.n9 A_MUX_4.Tr_Gate_1.CLK.t4 3.6405
R17659 A_MUX_4.Tr_Gate_1.CLK.n9 A_MUX_4.Tr_Gate_1.CLK.n8 3.6405
R17660 A_MUX_4.Tr_Gate_1.CLK.n13 A_MUX_4.Tr_Gate_1.CLK.t3 3.6405
R17661 A_MUX_4.Tr_Gate_1.CLK.n13 A_MUX_4.Tr_Gate_1.CLK.n12 3.6405
R17662 A_MUX_4.Tr_Gate_1.CLK.n1 A_MUX_4.Tr_Gate_1.CLK.n3 3.50463
R17663 A_MUX_4.Tr_Gate_1.CLK.n0 A_MUX_4.Tr_Gate_1.CLK.n5 3.50463
R17664 A_MUX_4.Tr_Gate_1.CLK.n3 A_MUX_4.Tr_Gate_1.CLK.t2 3.2765
R17665 A_MUX_4.Tr_Gate_1.CLK.n3 A_MUX_4.Tr_Gate_1.CLK.n2 3.2765
R17666 A_MUX_4.Tr_Gate_1.CLK.n5 A_MUX_4.Tr_Gate_1.CLK.t6 3.2765
R17667 A_MUX_4.Tr_Gate_1.CLK.n5 A_MUX_4.Tr_Gate_1.CLK.n4 3.2765
R17668 A_MUX_4.Tr_Gate_1.CLK.n0 A_MUX_4.Tr_Gate_1.CLK.n9 3.06224
R17669 A_MUX_4.Tr_Gate_1.CLK.n1 A_MUX_4.Tr_Gate_1.CLK.n11 3.06224
R17670 A_MUX_4.Tr_Gate_1.CLK.n0 A_MUX_4.Tr_Gate_1.CLK.n7 2.6005
R17671 A_MUX_4.Tr_Gate_1.CLK.n1 A_MUX_4.Tr_Gate_1.CLK.n13 2.6005
R17672 A_MUX_4.Tr_Gate_1.CLK A_MUX_4.Tr_Gate_1.CLK.n1 1.444
R17673 A_MUX_4.Tr_Gate_1.CLK.n1 A_MUX_4.Tr_Gate_1.CLK.n0 1.1705
R17674 a_27423_7180.n5 a_27423_7180.t8 29.3691
R17675 a_27423_7180.n6 a_27423_7180.n5 21.9292
R17676 a_27423_7180.n7 a_27423_7180.n6 18.1271
R17677 a_27423_7180.n7 a_27423_7180.t7 11.2425
R17678 a_27423_7180.n3 a_27423_7180.t0 10.2135
R17679 a_27423_7180.n5 a_27423_7180.t9 6.1325
R17680 a_27423_7180.n6 a_27423_7180.t6 6.1325
R17681 a_27423_7180.n3 a_27423_7180.n2 4.68398
R17682 a_27423_7180.n8 a_27423_7180.n7 4.6302
R17683 a_27423_7180.n9 a_27423_7180.n8 2.85093
R17684 a_27423_7180.n1 a_27423_7180.t4 2.16717
R17685 a_27423_7180.n1 a_27423_7180.n0 2.16717
R17686 a_27423_7180.n9 a_27423_7180.t2 2.16717
R17687 a_27423_7180.n10 a_27423_7180.n9 2.16717
R17688 a_27423_7180.n4 a_27423_7180.n3 1.58582
R17689 a_27423_7180.n4 a_27423_7180.n1 1.24371
R17690 a_27423_7180.n8 a_27423_7180.n4 0.971051
R17691 a_44728_10426.t0 a_44728_10426.t1 12.9675
R17692 a_44428_9804.t0 a_44428_9804.t1 12.9675
R17693 a_27480_10186.n2 a_27480_10186.t7 29.3691
R17694 a_27480_10186.n3 a_27480_10186.n2 21.9292
R17695 a_27480_10186.n4 a_27480_10186.n3 18.1271
R17696 a_27480_10186.n4 a_27480_10186.t9 11.2425
R17697 a_27480_10186.n7 a_27480_10186.t1 10.2135
R17698 a_27480_10186.n2 a_27480_10186.t6 6.1325
R17699 a_27480_10186.n3 a_27480_10186.t8 6.1325
R17700 a_27480_10186.n7 a_27480_10186.n6 4.68398
R17701 a_27480_10186.n5 a_27480_10186.n4 4.6302
R17702 a_27480_10186.n5 a_27480_10186.n1 2.85093
R17703 a_27480_10186.n1 a_27480_10186.t2 2.16717
R17704 a_27480_10186.n1 a_27480_10186.n0 2.16717
R17705 a_27480_10186.n9 a_27480_10186.t3 2.16717
R17706 a_27480_10186.n10 a_27480_10186.n9 2.16717
R17707 a_27480_10186.n8 a_27480_10186.n7 1.58618
R17708 a_27480_10186.n9 a_27480_10186.n8 1.24388
R17709 a_27480_10186.n8 a_27480_10186.n5 0.97169
R17710 S4.n16 S4.t18 45.6363
R17711 S4.n12 S4.t13 29.6446
R17712 S4.t14 S4.n13 29.6446
R17713 S4.n11 S4.t20 24.6117
R17714 S4.n5 S4.t6 23.6945
R17715 S4.n6 S4.t12 23.6945
R17716 S4.n13 S4.n12 22.2047
R17717 S4.t18 S4.t3 22.1925
R17718 S4.n17 S4.n16 20.9314
R17719 S4.n6 S4.n5 18.8035
R17720 S4 S4.t14 18.5175
R17721 S4.n3 S4.n0 15.8172
R17722 S4.n9 S4.n8 15.8172
R17723 S4.n8 S4.n0 15.8172
R17724 S4.t9 S4.n3 14.8925
R17725 S4.t15 S4.n0 14.8925
R17726 S4.n8 S4.t4 14.8925
R17727 S4.n7 S4.n1 12.2457
R17728 S4.n7 S4.n2 12.2457
R17729 S4.n4 S4.n2 12.2457
R17730 S4.n10 S4.t16 11.6285
R17731 S4.t6 S4.n4 8.9065
R17732 S4.t11 S4.n2 8.9065
R17733 S4.n7 S4.t0 8.9065
R17734 S4.t12 S4.n1 8.9065
R17735 S4.n3 S4.t10 8.6145
R17736 S4.n0 S4.t17 8.6145
R17737 S4.n8 S4.t5 8.6145
R17738 S4.n9 S4.t19 8.59715
R17739 S4.n4 S4.t9 8.3225
R17740 S4.n2 S4.t15 8.3225
R17741 S4.t4 S4.n7 8.3225
R17742 S4.n1 S4.t16 8.3225
R17743 S4.n11 S4.t7 6.1325
R17744 S4.n12 S4.t1 6.1325
R17745 S4.n13 S4.t2 6.1325
R17746 S4.n16 S4.t8 6.1325
R17747 S4.n17 S4.t21 6.1325
R17748 S4.n18 S4.n17 4.86779
R17749 S4.n14 S4.n11 4.79907
R17750 S4 S4.n10 4.223
R17751 S4.n5 S4.t11 3.6505
R17752 S4.t0 S4.n6 3.6505
R17753 S4.n10 S4.n9 3.1807
R17754 S4.n19 S4.n18 2.65123
R17755 S4.n14 S4 0.640368
R17756 S4.n15 S4 0.1655
R17757 S4.n18 S4.n15 0.109537
R17758 S4.n19 S4 0.0733182
R17759 S4.n15 S4.n14 0.0592755
R17760 S4 S4.n19 0.0318393
R17761 a_42628_9598.t0 a_42628_9598.t1 12.9675
R17762 a_42928_8976.t0 a_42928_8976.t1 12.9675
R17763 a_44728_12082.t0 a_44728_12082.t1 12.9675
R17764 a_44428_11460.t0 a_44428_11460.t1 12.9675
R17765 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n3 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n2 5.81586
R17766 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t13 5.10148
R17767 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n5 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t14 5.1005
R17768 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n4 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t3 5.08021
R17769 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n7 4.66266
R17770 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t9 3.6405
R17771 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n18 3.6405
R17772 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t16 3.6405
R17773 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n20 3.6405
R17774 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t17 3.6405
R17775 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n11 3.6405
R17776 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n14 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t7 3.6405
R17777 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n14 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n13 3.6405
R17778 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n17 3.50463
R17779 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n10 3.50463
R17780 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t5 3.2765
R17781 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n16 3.2765
R17782 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t8 3.2765
R17783 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n9 3.2765
R17784 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n21 3.06224
R17785 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n14 3.06224
R17786 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n3 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n1 2.85093
R17787 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n19 2.6005
R17788 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n12 2.6005
R17789 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t1 2.16717
R17790 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n0 2.16717
R17791 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.t15 1.9505
R17792 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n6 1.9505
R17793 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n23 0.798761
R17794 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n4 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n3 0.644196
R17795 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n24 0.562022
R17796 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n5 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n4 0.447229
R17797 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n5 0.392597
R17798 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n8 0.308628
R17799 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n22 0.18637
R17800 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT.n15 0.18637
R17801 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t27 23.6945
R17802 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t16 23.6945
R17803 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n17 18.8035
R17804 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n12 15.8172
R17805 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n20 15.8172
R17806 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n12 15.8172
R17807 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n15 14.8925
R17808 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t25 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n12 14.8925
R17809 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t22 14.8925
R17810 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n13 12.2457
R17811 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n14 12.2457
R17812 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n14 12.2457
R17813 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t20 11.6285
R17814 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n16 8.9065
R17815 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n14 8.9065
R17816 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t24 8.9065
R17817 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n13 8.9065
R17818 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t23 8.6145
R17819 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t21 8.6145
R17820 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t19 8.6145
R17821 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t17 8.59715
R17822 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t26 8.3225
R17823 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n14 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t25 8.3225
R17824 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n19 8.3225
R17825 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n13 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t20 8.3225
R17826 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n33 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 6.97731
R17827 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n0 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n29 6.74326
R17828 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n7 6.74326
R17829 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n0 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n30 5.1005
R17830 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n8 5.1005
R17831 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n22 4.21749
R17832 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t18 3.6505
R17833 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n18 3.6505
R17834 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n24 3.57508
R17835 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n5 3.5743
R17836 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n0 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t13 3.40075
R17837 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t6 3.40065
R17838 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n21 3.1807
R17839 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n9 3.00096
R17840 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n28 3.00032
R17841 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n32 2.58093
R17842 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n11 2.58093
R17843 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t4 2.16717
R17844 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n25 2.16717
R17845 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t1 2.16717
R17846 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n23 2.16717
R17847 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n3 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t0 2.16717
R17848 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n3 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n2 2.16717
R17849 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n5 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.t9 2.16717
R17850 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n5 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n4 2.16717
R17851 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n32 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n31 1.84797
R17852 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n11 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n10 1.84666
R17853 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n27 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n26 1.25233
R17854 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n3 1.25225
R17855 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n11 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n6 1.12594
R17856 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n32 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n27 1.12574
R17857 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n33 0.812356
R17858 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n33 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 0.728851
R17859 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n1 0.558764
R17860 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN.n0 0.558374
R17861 a_41879_1284.n2 a_41879_1284.t6 29.3691
R17862 a_41879_1284.n3 a_41879_1284.n2 21.9292
R17863 a_41879_1284.n4 a_41879_1284.n3 18.1271
R17864 a_41879_1284.n4 a_41879_1284.t8 11.2425
R17865 a_41879_1284.n7 a_41879_1284.t0 10.2135
R17866 a_41879_1284.n2 a_41879_1284.t7 6.1325
R17867 a_41879_1284.n3 a_41879_1284.t9 6.1325
R17868 a_41879_1284.n7 a_41879_1284.n6 4.68398
R17869 a_41879_1284.n5 a_41879_1284.n4 4.6302
R17870 a_41879_1284.n5 a_41879_1284.n1 2.85093
R17871 a_41879_1284.n1 a_41879_1284.t2 2.16717
R17872 a_41879_1284.n1 a_41879_1284.n0 2.16717
R17873 a_41879_1284.n9 a_41879_1284.t3 2.16717
R17874 a_41879_1284.n10 a_41879_1284.n9 2.16717
R17875 a_41879_1284.n8 a_41879_1284.n7 1.58618
R17876 a_41879_1284.n9 a_41879_1284.n8 1.24388
R17877 a_41879_1284.n8 a_41879_1284.n5 0.97169
R17878 a_44428_11254.t0 a_44428_11254.t1 12.9675
R17879 a_44728_10632.t0 a_44728_10632.t1 12.9675
R17880 a_23836_10693.t2 a_23836_10693.n5 6.64563
R17881 a_23836_10693.n5 a_23836_10693.t3 6.61433
R17882 a_23836_10693.n4 a_23836_10693.n3 3.36963
R17883 a_23836_10693.n4 a_23836_10693.n1 3.33833
R17884 a_23836_10693.n3 a_23836_10693.t0 3.2765
R17885 a_23836_10693.n3 a_23836_10693.n2 3.2765
R17886 a_23836_10693.n1 a_23836_10693.t4 3.2765
R17887 a_23836_10693.n1 a_23836_10693.n0 3.2765
R17888 a_23836_10693.n5 a_23836_10693.n4 0.781777
R17889 a_45928_10426.t0 a_45928_10426.t1 12.9675
R17890 a_46228_9804.t0 a_46228_9804.t1 12.9675
R17891 a_44428_9598.t0 a_44428_9598.t1 12.9675
R17892 a_44128_8976.t0 a_44128_8976.t1 12.9675
R17893 a_42763_5679.n5 a_42763_5679.t9 29.2961
R17894 a_42763_5679.n6 a_42763_5679.n5 21.9292
R17895 a_42763_5679.n7 a_42763_5679.n6 18.1271
R17896 a_42763_5679.n7 a_42763_5679.t8 11.1695
R17897 a_42763_5679.n3 a_42763_5679.t0 10.2143
R17898 a_42763_5679.n5 a_42763_5679.t7 6.1325
R17899 a_42763_5679.n6 a_42763_5679.t6 6.1325
R17900 a_42763_5679.n3 a_42763_5679.n2 4.68517
R17901 a_42763_5679.n8 a_42763_5679.n7 4.6311
R17902 a_42763_5679.n10 a_42763_5679.n8 2.85093
R17903 a_42763_5679.n1 a_42763_5679.t2 2.16717
R17904 a_42763_5679.n1 a_42763_5679.n0 2.16717
R17905 a_42763_5679.t5 a_42763_5679.n10 2.16717
R17906 a_42763_5679.n10 a_42763_5679.n9 2.16717
R17907 a_42763_5679.n4 a_42763_5679.n3 1.58582
R17908 a_42763_5679.n4 a_42763_5679.n1 1.24371
R17909 a_42763_5679.n8 a_42763_5679.n4 0.971051
R17910 a_45928_8770.t0 a_45928_8770.t1 12.9675
R17911 a_45628_8148.t0 a_45628_8148.t1 12.9675
R17912 a_42628_8770.t0 a_42628_8770.t1 10.2205
R17913 a_42628_8148.t0 a_42628_8148.t1 12.9675
R17914 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t23 23.6945
R17915 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n21 23.6945
R17916 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n20 18.8035
R17917 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n16 15.8172
R17918 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n17 15.8172
R17919 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n13 15.8172
R17920 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t30 14.8925
R17921 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n18 14.8925
R17922 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t20 14.8925
R17923 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n14 12.2457
R17924 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n14 12.2457
R17925 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n15 12.2457
R17926 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t26 11.6285
R17927 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n15 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t23 8.9065
R17928 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n19 8.9065
R17929 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t28 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n14 8.9065
R17930 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n22 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t21 8.9065
R17931 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n18 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t25 8.6145
R17932 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n16 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t24 8.6145
R17933 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n17 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t27 8.6145
R17934 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n13 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t29 8.59715
R17935 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t30 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n15 8.3225
R17936 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n19 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t22 8.3225
R17937 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n14 8.3225
R17938 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n22 8.3225
R17939 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n12 5.24044
R17940 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n4 5.10151
R17941 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n3 5.10119
R17942 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n2 5.08021
R17943 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n7 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n6 4.66164
R17944 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n23 4.223
R17945 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n20 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t31 3.6505
R17946 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n21 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t28 3.6505
R17947 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n37 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t10 3.6405
R17948 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n37 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n36 3.6405
R17949 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n28 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t7 3.6405
R17950 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n28 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n27 3.6405
R17951 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t6 3.6405
R17952 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n26 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n25 3.6405
R17953 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n35 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t9 3.6405
R17954 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n35 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n34 3.6405
R17955 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n39 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n33 3.50463
R17956 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n40 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n31 3.50463
R17957 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t14 3.40711
R17958 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n33 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t4 3.2765
R17959 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n33 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n32 3.2765
R17960 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t2 3.2765
R17961 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n31 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n30 3.2765
R17962 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n23 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n13 3.1807
R17963 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n26 3.06224
R17964 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n38 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n35 3.06224
R17965 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n11 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n1 2.85093
R17966 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n29 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n28 2.6005
R17967 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n38 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n37 2.6005
R17968 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 2.36593
R17969 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t1 2.16717
R17970 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n1 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n0 2.16717
R17971 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n24 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 2.01183
R17972 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.t19 1.9505
R17973 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n6 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n5 1.9505
R17974 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n12 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n11 1.0205
R17975 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n40 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n39 0.798761
R17976 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n11 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n10 0.644196
R17977 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n40 0.562022
R17978 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n10 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n9 0.450799
R17979 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n7 0.358456
R17980 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n24 0.278326
R17981 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n9 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n8 0.229792
R17982 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n40 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n29 0.18637
R17983 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n39 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT.n38 0.18637
R17984 S5.n16 S5.t17 45.6363
R17985 S5.n12 S5.t20 29.6446
R17986 S5.t8 S5.n13 29.6446
R17987 S5.n11 S5.t10 24.6117
R17988 S5.n7 S5.t2 23.6945
R17989 S5.t13 S5.n8 23.6945
R17990 S5.n13 S5.n12 22.2047
R17991 S5.t17 S5.t7 22.1925
R17992 S5.n17 S5.n16 20.9314
R17993 S5.n8 S5.n7 18.8035
R17994 S5 S5.t8 18.5175
R17995 S5.n5 S5.n3 15.8172
R17996 S5.n4 S5.n0 15.8172
R17997 S5.n5 S5.n4 15.8172
R17998 S5.n3 S5.t14 14.8925
R17999 S5.t0 S5.n5 14.8925
R18000 S5.n4 S5.t15 14.8925
R18001 S5.n9 S5.n1 12.2457
R18002 S5.n6 S5.n1 12.2457
R18003 S5.n6 S5.n2 12.2457
R18004 S5.n10 S5.t5 11.6285
R18005 S5.n2 S5.t2 8.9065
R18006 S5.t11 S5.n6 8.9065
R18007 S5.t3 S5.n1 8.9065
R18008 S5.n9 S5.t13 8.9065
R18009 S5.n5 S5.t4 8.6145
R18010 S5.n3 S5.t18 8.6145
R18011 S5.n4 S5.t19 8.6145
R18012 S5.n0 S5.t6 8.59715
R18013 S5.n19 S5 8.37523
R18014 S5.t14 S5.n2 8.3225
R18015 S5.n6 S5.t0 8.3225
R18016 S5.t15 S5.n1 8.3225
R18017 S5.t5 S5.n9 8.3225
R18018 S5.n11 S5.t1 6.1325
R18019 S5.n16 S5.t21 6.1325
R18020 S5.n17 S5.t12 6.1325
R18021 S5.n12 S5.t9 6.1325
R18022 S5.n13 S5.t16 6.1325
R18023 S5.n18 S5.n17 4.86652
R18024 S5.n14 S5.n11 4.79907
R18025 S5 S5.n10 4.223
R18026 S5.n7 S5.t11 3.6505
R18027 S5.n8 S5.t3 3.6505
R18028 S5.n10 S5.n0 3.1807
R18029 S5.n19 S5.n18 1.77452
R18030 S5 S5.n19 0.867837
R18031 S5.n14 S5 0.640368
R18032 S5.n15 S5 0.1655
R18033 S5.n18 S5.n15 0.108908
R18034 S5.n15 S5.n14 0.0592755
R18035 A_MUX_6.Tr_Gate_1.CLK.n1 A_MUX_6.Tr_Gate_1.CLK.t16 45.6363
R18036 A_MUX_6.Tr_Gate_1.CLK.n3 A_MUX_6.Tr_Gate_1.CLK.t18 29.6446
R18037 A_MUX_6.Tr_Gate_1.CLK.t15 A_MUX_6.Tr_Gate_1.CLK.n4 29.6446
R18038 A_MUX_6.Tr_Gate_1.CLK.n5 A_MUX_6.Tr_Gate_1.CLK.t12 24.6117
R18039 A_MUX_6.Tr_Gate_1.CLK.n4 A_MUX_6.Tr_Gate_1.CLK.n3 22.2047
R18040 A_MUX_6.Tr_Gate_1.CLK.t16 A_MUX_6.Tr_Gate_1.CLK.t21 22.1925
R18041 A_MUX_6.Tr_Gate_1.CLK.n2 A_MUX_6.Tr_Gate_1.CLK.n1 20.9314
R18042 A_MUX_6.Tr_Gate_1.CLK A_MUX_6.Tr_Gate_1.CLK.t15 18.5245
R18043 A_MUX_6.Tr_Gate_1.CLK.n1 A_MUX_6.Tr_Gate_1.CLK.t17 6.1325
R18044 A_MUX_6.Tr_Gate_1.CLK.n2 A_MUX_6.Tr_Gate_1.CLK.t13 6.1325
R18045 A_MUX_6.Tr_Gate_1.CLK.n3 A_MUX_6.Tr_Gate_1.CLK.t14 6.1325
R18046 A_MUX_6.Tr_Gate_1.CLK.n4 A_MUX_6.Tr_Gate_1.CLK.t19 6.1325
R18047 A_MUX_6.Tr_Gate_1.CLK.n5 A_MUX_6.Tr_Gate_1.CLK.t20 6.1325
R18048 A_MUX_6.Tr_Gate_1.CLK.n0 A_MUX_6.Tr_Gate_1.CLK.n2 5.28481
R18049 A_MUX_6.Tr_Gate_1.CLK.n0 A_MUX_6.Tr_Gate_1.CLK.n5 4.89628
R18050 A_MUX_6.Tr_Gate_1.CLK.n17 A_MUX_6.Tr_Gate_1.CLK.t10 3.6405
R18051 A_MUX_6.Tr_Gate_1.CLK.n17 A_MUX_6.Tr_Gate_1.CLK.n16 3.6405
R18052 A_MUX_6.Tr_Gate_1.CLK.n11 A_MUX_6.Tr_Gate_1.CLK.t4 3.6405
R18053 A_MUX_6.Tr_Gate_1.CLK.n11 A_MUX_6.Tr_Gate_1.CLK.n10 3.6405
R18054 A_MUX_6.Tr_Gate_1.CLK.n13 A_MUX_6.Tr_Gate_1.CLK.t9 3.6405
R18055 A_MUX_6.Tr_Gate_1.CLK.n13 A_MUX_6.Tr_Gate_1.CLK.n12 3.6405
R18056 A_MUX_6.Tr_Gate_1.CLK.n19 A_MUX_6.Tr_Gate_1.CLK.t5 3.6405
R18057 A_MUX_6.Tr_Gate_1.CLK.n19 A_MUX_6.Tr_Gate_1.CLK.n18 3.6405
R18058 A_MUX_6.Tr_Gate_1.CLK.n21 A_MUX_6.Tr_Gate_1.CLK.n7 3.50463
R18059 A_MUX_6.Tr_Gate_1.CLK.n15 A_MUX_6.Tr_Gate_1.CLK.n9 3.50463
R18060 A_MUX_6.Tr_Gate_1.CLK.n7 A_MUX_6.Tr_Gate_1.CLK.t1 3.2765
R18061 A_MUX_6.Tr_Gate_1.CLK.n7 A_MUX_6.Tr_Gate_1.CLK.n6 3.2765
R18062 A_MUX_6.Tr_Gate_1.CLK.n9 A_MUX_6.Tr_Gate_1.CLK.t0 3.2765
R18063 A_MUX_6.Tr_Gate_1.CLK.n9 A_MUX_6.Tr_Gate_1.CLK.n8 3.2765
R18064 A_MUX_6.Tr_Gate_1.CLK.n14 A_MUX_6.Tr_Gate_1.CLK.n13 3.06224
R18065 A_MUX_6.Tr_Gate_1.CLK.n20 A_MUX_6.Tr_Gate_1.CLK.n17 3.06224
R18066 A_MUX_6.Tr_Gate_1.CLK.n14 A_MUX_6.Tr_Gate_1.CLK.n11 2.6005
R18067 A_MUX_6.Tr_Gate_1.CLK.n20 A_MUX_6.Tr_Gate_1.CLK.n19 2.6005
R18068 A_MUX_6.Tr_Gate_1.CLK.n21 A_MUX_6.Tr_Gate_1.CLK.n15 0.798761
R18069 A_MUX_6.Tr_Gate_1.CLK.n0 A_MUX_6.Tr_Gate_1.CLK 0.629601
R18070 A_MUX_6.Tr_Gate_1.CLK A_MUX_6.Tr_Gate_1.CLK.n21 0.562022
R18071 A_MUX_6.Tr_Gate_1.CLK A_MUX_6.Tr_Gate_1.CLK.n0 0.253378
R18072 A_MUX_6.Tr_Gate_1.CLK.n15 A_MUX_6.Tr_Gate_1.CLK.n14 0.18637
R18073 A_MUX_6.Tr_Gate_1.CLK.n21 A_MUX_6.Tr_Gate_1.CLK.n20 0.18637
R18074 DN1.n14 DN1.n11 6.76498
R18075 DN1.n3 DN1.n2 5.81586
R18076 DN1.n8 DN1.t1 5.10151
R18077 DN1.n5 DN1.t3 5.1005
R18078 DN1.n4 DN1.t6 5.08021
R18079 DN1.n8 DN1.n7 4.66164
R18080 DN1.n13 DN1.t10 3.6405
R18081 DN1.n13 DN1.n12 3.6405
R18082 DN1.n3 DN1.n1 2.85093
R18083 DN1.n14 DN1.n13 2.78441
R18084 DN1.n15 DN1.n10 2.75034
R18085 DN1.n1 DN1.t4 2.16717
R18086 DN1.n1 DN1.n0 2.16717
R18087 DN1.n7 DN1.t2 1.9505
R18088 DN1.n7 DN1.n6 1.9505
R18089 DN1.n10 DN1 1.50193
R18090 DN1.n10 DN1 0.928286
R18091 DN1.n4 DN1.n3 0.644196
R18092 DN1.n5 DN1.n4 0.447229
R18093 DN1 DN1.n14 0.362337
R18094 DN1.n9 DN1.n8 0.254356
R18095 DN1.n9 DN1.n5 0.22163
R18096 DN1 DN1.n9 0.127741
R18097 DN1.n15 DN1 0.109424
R18098 DN1.n16 DN1.n15 0.0302355
R18099 DN1.n16 DN1 0.00368003
R18100 DN1 DN1.n16 0.00103006
R18101 a_39080_11413.n0 a_39080_11413.t7 29.3691
R18102 a_39080_11413.n1 a_39080_11413.n0 21.9292
R18103 a_39080_11413.n2 a_39080_11413.n1 18.1271
R18104 a_39080_11413.n2 a_39080_11413.t8 11.2425
R18105 a_39080_11413.n6 a_39080_11413.n5 10.1038
R18106 a_39080_11413.n0 a_39080_11413.t9 6.1325
R18107 a_39080_11413.n1 a_39080_11413.t6 6.1325
R18108 a_39080_11413.n6 a_39080_11413.t0 4.70149
R18109 a_39080_11413.n8 a_39080_11413.n2 4.6302
R18110 a_39080_11413.n9 a_39080_11413.n8 2.85093
R18111 a_39080_11413.n4 a_39080_11413.t2 2.16717
R18112 a_39080_11413.n4 a_39080_11413.n3 2.16717
R18113 a_39080_11413.n9 a_39080_11413.t3 2.16717
R18114 a_39080_11413.n10 a_39080_11413.n9 2.16717
R18115 a_39080_11413.n7 a_39080_11413.n6 1.58582
R18116 a_39080_11413.n7 a_39080_11413.n4 1.24371
R18117 a_39080_11413.n8 a_39080_11413.n7 0.971051
R18118 a_24436_11277.n2 a_24436_11277.t2 7.21081
R18119 a_24436_11277.n3 a_24436_11277.n2 7.15165
R18120 a_24436_11277.n1 a_24436_11277.t0 3.6405
R18121 a_24436_11277.n1 a_24436_11277.n0 3.6405
R18122 a_24436_11277.n2 a_24436_11277.n1 2.77149
R18123 a_45158_5339.n0 a_45158_5339.t8 29.2961
R18124 a_45158_5339.n1 a_45158_5339.n0 21.9292
R18125 a_45158_5339.n2 a_45158_5339.n1 18.1271
R18126 a_45158_5339.n2 a_45158_5339.t6 11.1695
R18127 a_45158_5339.n0 a_45158_5339.t7 6.1325
R18128 a_45158_5339.n1 a_45158_5339.t9 6.1325
R18129 a_45158_5339.n6 a_45158_5339.n5 4.93252
R18130 a_45158_5339.n6 a_45158_5339.t0 4.70348
R18131 a_45158_5339.n8 a_45158_5339.n2 4.6311
R18132 a_45158_5339.n10 a_45158_5339.n8 2.85093
R18133 a_45158_5339.n4 a_45158_5339.t4 2.16717
R18134 a_45158_5339.n4 a_45158_5339.n3 2.16717
R18135 a_45158_5339.t5 a_45158_5339.n10 2.16717
R18136 a_45158_5339.n10 a_45158_5339.n9 2.16717
R18137 a_45158_5339.n7 a_45158_5339.n6 1.58582
R18138 a_45158_5339.n7 a_45158_5339.n4 1.24371
R18139 a_45158_5339.n8 a_45158_5339.n7 0.971051
R18140 a_45328_12082.t0 a_45328_12082.t1 12.9675
R18141 a_45628_11460.t0 a_45628_11460.t1 12.9675
R18142 F_IN.n6 F_IN.n5 5.81586
R18143 F_IN.n8 F_IN.t4 5.10208
R18144 F_IN.n2 F_IN.t5 5.10195
R18145 F_IN.n7 F_IN.t0 5.08021
R18146 F_IN.n2 F_IN.n1 4.66211
R18147 F_IN.n6 F_IN.n4 2.85093
R18148 F_IN.n4 F_IN.t1 2.16717
R18149 F_IN.n4 F_IN.n3 2.16717
R18150 F_IN.n10 F_IN 2.0861
R18151 F_IN.n1 F_IN.t6 1.9505
R18152 F_IN.n1 F_IN.n0 1.9505
R18153 F_IN F_IN.n10 0.911144
R18154 F_IN.n7 F_IN.n6 0.644196
R18155 F_IN.n10 F_IN 0.643183
R18156 F_IN.n8 F_IN.n7 0.449473
R18157 F_IN.n9 F_IN.n2 0.212726
R18158 F_IN.n9 F_IN.n8 0.198082
R18159 F_IN F_IN.n9 0.0718702
R18160 S3.n16 S3.t7 45.6363
R18161 S3.n12 S3.t14 29.6446
R18162 S3.t17 S3.n13 29.6446
R18163 S3.n11 S3.t13 24.6117
R18164 S3.n7 S3.t0 23.6945
R18165 S3.t9 S3.n8 23.6945
R18166 S3.n13 S3.n12 22.2047
R18167 S3.t7 S3.t18 22.1925
R18168 S3.n17 S3.n16 20.9314
R18169 S3.n8 S3.n7 18.8035
R18170 S3 S3.t17 18.5191
R18171 S3.n5 S3.n3 15.8172
R18172 S3.n5 S3.n4 15.8172
R18173 S3.n4 S3.n0 15.8172
R18174 S3.n3 S3.t11 14.8925
R18175 S3.t8 S3.n5 14.8925
R18176 S3.n4 S3.t2 14.8925
R18177 S3.n9 S3.n1 12.2457
R18178 S3.n6 S3.n1 12.2457
R18179 S3.n6 S3.n2 12.2457
R18180 S3.n10 S3.t21 11.6285
R18181 S3.n2 S3.t0 8.9065
R18182 S3.t20 S3.n6 8.9065
R18183 S3.t12 S3.n1 8.9065
R18184 S3.n9 S3.t9 8.9065
R18185 S3.n5 S3.t6 8.6145
R18186 S3.n3 S3.t10 8.6145
R18187 S3.n4 S3.t1 8.6145
R18188 S3.n0 S3.t19 8.59715
R18189 S3.t11 S3.n2 8.3225
R18190 S3.n6 S3.t8 8.3225
R18191 S3.t2 S3.n1 8.3225
R18192 S3.t21 S3.n9 8.3225
R18193 S3.n19 S3 8.17889
R18194 S3.n11 S3.t15 6.1325
R18195 S3.n16 S3.t4 6.1325
R18196 S3.n17 S3.t5 6.1325
R18197 S3.n12 S3.t3 6.1325
R18198 S3.n13 S3.t16 6.1325
R18199 S3.n18 S3.n17 4.86652
R18200 S3.n14 S3.n11 4.79907
R18201 S3 S3.n10 4.223
R18202 S3.n7 S3.t20 3.6505
R18203 S3.n8 S3.t12 3.6505
R18204 S3.n10 S3.n0 3.1807
R18205 S3.n19 S3.n18 1.7553
R18206 S3 S3.n19 0.866502
R18207 S3.n14 S3 0.640368
R18208 S3.n15 S3 0.1655
R18209 S3.n18 S3.n15 0.108908
R18210 S3.n15 S3.n14 0.0592755
R18211 a_44128_8770.t0 a_44128_8770.t1 12.9675
R18212 a_43828_8148.t0 a_43828_8148.t1 12.9675
R18213 a_20945_11785.n0 a_20945_11785.t7 29.3691
R18214 a_20945_11785.n1 a_20945_11785.n0 21.9292
R18215 a_20945_11785.n2 a_20945_11785.n1 18.1271
R18216 a_20945_11785.n2 a_20945_11785.t8 11.2425
R18217 a_20945_11785.n6 a_20945_11785.n5 10.1038
R18218 a_20945_11785.n0 a_20945_11785.t9 6.1325
R18219 a_20945_11785.n1 a_20945_11785.t6 6.1325
R18220 a_20945_11785.n6 a_20945_11785.t0 4.70149
R18221 a_20945_11785.n8 a_20945_11785.n2 4.6302
R18222 a_20945_11785.n9 a_20945_11785.n8 2.85093
R18223 a_20945_11785.n4 a_20945_11785.t2 2.16717
R18224 a_20945_11785.n4 a_20945_11785.n3 2.16717
R18225 a_20945_11785.n9 a_20945_11785.t3 2.16717
R18226 a_20945_11785.n10 a_20945_11785.n9 2.16717
R18227 a_20945_11785.n7 a_20945_11785.n6 1.58582
R18228 a_20945_11785.n7 a_20945_11785.n4 1.24371
R18229 a_20945_11785.n8 a_20945_11785.n7 0.971051
R18230 a_36685_10901.n3 a_36685_10901.t6 29.3691
R18231 a_36685_10901.n4 a_36685_10901.n3 21.9292
R18232 a_36685_10901.n5 a_36685_10901.n4 18.1271
R18233 a_36685_10901.n5 a_36685_10901.t9 11.2425
R18234 a_36685_10901.n8 a_36685_10901.t0 10.2135
R18235 a_36685_10901.n3 a_36685_10901.t8 6.1325
R18236 a_36685_10901.n4 a_36685_10901.t7 6.1325
R18237 a_36685_10901.n8 a_36685_10901.n7 4.68398
R18238 a_36685_10901.n6 a_36685_10901.n5 4.6302
R18239 a_36685_10901.n6 a_36685_10901.n2 2.85093
R18240 a_36685_10901.n2 a_36685_10901.t4 2.16717
R18241 a_36685_10901.n2 a_36685_10901.n1 2.16717
R18242 a_36685_10901.t5 a_36685_10901.n10 2.16717
R18243 a_36685_10901.n10 a_36685_10901.n0 2.16717
R18244 a_36685_10901.n9 a_36685_10901.n8 1.58618
R18245 a_36685_10901.n10 a_36685_10901.n9 1.24388
R18246 a_36685_10901.n9 a_36685_10901.n6 0.97169
R18247 ITAIL1.n5 ITAIL1.n4 28.0418
R18248 ITAIL1.n3 ITAIL1.n2 14.6005
R18249 ITAIL1.n13 ITAIL1 9.56592
R18250 ITAIL1.n1 ITAIL1.n0 7.61735
R18251 ITAIL1.n1 ITAIL1.t5 7.20135
R18252 ITAIL1.n8 ITAIL1.n7 6.82463
R18253 ITAIL1.n10 ITAIL1.t6 6.77907
R18254 ITAIL1.n5 ITAIL1.t0 6.71389
R18255 ITAIL1.n2 ITAIL1.t8 6.51836
R18256 ITAIL1.n2 ITAIL1.t2 6.51836
R18257 ITAIL1.n3 ITAIL1.t13 6.51836
R18258 ITAIL1.n10 ITAIL1.t11 6.25764
R18259 ITAIL1.n4 ITAIL1.t4 6.25764
R18260 ITAIL1.n6 ITAIL1.t9 6.19246
R18261 ITAIL1.n11 ITAIL1.t7 5.89613
R18262 ITAIL1.n11 ITAIL1.n10 4.23548
R18263 ITAIL1.n8 ITAIL1.n6 4.21461
R18264 ITAIL1 ITAIL1.n13 2.36014
R18265 ITAIL1.n9 ITAIL1.n8 1.42665
R18266 ITAIL1.n12 ITAIL1.n11 1.13763
R18267 ITAIL1.n13 ITAIL1.n12 0.562798
R18268 ITAIL1.n12 ITAIL1.n9 0.474918
R18269 ITAIL1.n4 ITAIL1.n3 0.261214
R18270 ITAIL1.n9 ITAIL1.n1 0.2105
R18271 ITAIL1.n6 ITAIL1.n5 0.130857
R18272 a_45628_11254.t0 a_45628_11254.t1 12.9675
R18273 a_45328_10632.t0 a_45328_10632.t1 12.9675
R18274 a_22880_10947.n1 a_22880_10947.n0 6.53062
R18275 a_22880_10947.n1 a_22880_10947.t0 6.47087
R18276 a_22880_10947.n2 a_22880_10947.t2 3.357
R18277 a_22880_10947.n3 a_22880_10947.n2 3.0145
R18278 a_22880_10947.n2 a_22880_10947.n1 2.46697
R18279 a_29818_7696.n0 a_29818_7696.t9 29.3691
R18280 a_29818_7696.n1 a_29818_7696.n0 21.9292
R18281 a_29818_7696.n2 a_29818_7696.n1 18.1271
R18282 a_29818_7696.n2 a_29818_7696.t7 11.2425
R18283 a_29818_7696.n6 a_29818_7696.n5 10.1038
R18284 a_29818_7696.n0 a_29818_7696.t8 6.1325
R18285 a_29818_7696.n1 a_29818_7696.t6 6.1325
R18286 a_29818_7696.n6 a_29818_7696.t0 4.70149
R18287 a_29818_7696.n8 a_29818_7696.n2 4.6302
R18288 a_29818_7696.n9 a_29818_7696.n8 2.85093
R18289 a_29818_7696.n4 a_29818_7696.t3 2.16717
R18290 a_29818_7696.n4 a_29818_7696.n3 2.16717
R18291 a_29818_7696.n9 a_29818_7696.t4 2.16717
R18292 a_29818_7696.n10 a_29818_7696.n9 2.16717
R18293 a_29818_7696.n7 a_29818_7696.n6 1.58582
R18294 a_29818_7696.n7 a_29818_7696.n4 1.24371
R18295 a_29818_7696.n8 a_29818_7696.n7 0.971051
R18296 DN_INPUT.n15 DN_INPUT.n14 8.92809
R18297 DN_INPUT.n3 DN_INPUT.n0 8.0105
R18298 DN_INPUT.n17 DN_INPUT 7.17525
R18299 DN_INPUT.n6 DN_INPUT.n0 6.8405
R18300 DN_INPUT.n11 DN_INPUT.t4 5.81586
R18301 DN_INPUT.n5 DN_INPUT.n4 5.1005
R18302 DN_INPUT.n8 DN_INPUT.n7 5.1005
R18303 DN_INPUT.n13 DN_INPUT.n12 5.08021
R18304 DN_INPUT.n3 DN_INPUT.n2 4.6305
R18305 DN_INPUT.n11 DN_INPUT.n10 2.85093
R18306 DN_INPUT.n10 DN_INPUT.t7 2.16717
R18307 DN_INPUT.n10 DN_INPUT.n9 2.16717
R18308 DN_INPUT.n23 DN_INPUT 2.0861
R18309 DN_INPUT.n2 DN_INPUT.t3 1.9505
R18310 DN_INPUT.n2 DN_INPUT.n1 1.9505
R18311 DN_INPUT.n15 DN_INPUT.n6 0.818177
R18312 DN_INPUT.n23 DN_INPUT.n22 0.77774
R18313 DN_INPUT.n34 DN_INPUT.n33 0.667293
R18314 DN_INPUT.n13 DN_INPUT.n11 0.644196
R18315 DN_INPUT.n14 DN_INPUT.n13 0.400713
R18316 DN_INPUT.n16 DN_INPUT.n0 0.368
R18317 DN_INPUT.n8 DN_INPUT.n6 0.248625
R18318 DN_INPUT.n6 DN_INPUT.n5 0.237703
R18319 DN_INPUT DN_INPUT.n16 0.06675
R18320 DN_INPUT.n14 DN_INPUT.n8 0.0502872
R18321 DN_INPUT.n5 DN_INPUT.n3 0.0318043
R18322 DN_INPUT.n33 DN_INPUT.n32 0.0297566
R18323 DN_INPUT.n20 DN_INPUT.n19 0.0264322
R18324 DN_INPUT.n37 DN_INPUT.n36 0.016494
R18325 DN_INPUT.n28 DN_INPUT.n27 0.016494
R18326 DN_INPUT DN_INPUT.n39 0.0149608
R18327 DN_INPUT.n36 DN_INPUT.n35 0.0091747
R18328 DN_INPUT.n29 DN_INPUT.n28 0.0091747
R18329 DN_INPUT.n38 DN_INPUT.n37 0.00890361
R18330 DN_INPUT.n27 DN_INPUT.n26 0.00809036
R18331 DN_INPUT.n33 DN_INPUT.n23 0.00697489
R18332 DN_INPUT.n39 DN_INPUT.n38 0.00600723
R18333 DN_INPUT.n21 DN_INPUT.n20 0.00289709
R18334 DN_INPUT.n31 DN_INPUT.n30 0.00266867
R18335 DN_INPUT.n16 DN_INPUT.n15 0.0013148
R18336 DN_INPUT.n35 DN_INPUT.n34 0.00131325
R18337 DN_INPUT.n30 DN_INPUT.n29 0.00131325
R18338 DN_INPUT.n26 DN_INPUT.n25 0.00131325
R18339 DN_INPUT.n25 DN_INPUT.n24 0.00131325
R18340 DN_INPUT.n19 DN_INPUT.n18 0.00115375
R18341 DN_INPUT.n18 DN_INPUT.n17 0.00115375
R18342 DN_INPUT.n32 DN_INPUT.n31 0.00104217
R18343 DN_INPUT.n22 DN_INPUT.n21 0.000935835
R18344 a_22881_9554.n1 a_22881_9554.n0 6.53012
R18345 a_22881_9554.n1 a_22881_9554.t3 6.47102
R18346 a_22881_9554.t1 a_22881_9554.n3 3.35684
R18347 a_22881_9554.n3 a_22881_9554.n2 3.01376
R18348 a_22881_9554.n3 a_22881_9554.n1 2.46742
R18349 a_29875_10702.n0 a_29875_10702.t9 29.3691
R18350 a_29875_10702.n1 a_29875_10702.n0 21.9292
R18351 a_29875_10702.n2 a_29875_10702.n1 18.1271
R18352 a_29875_10702.n2 a_29875_10702.t7 11.2425
R18353 a_29875_10702.n6 a_29875_10702.n5 10.1038
R18354 a_29875_10702.n0 a_29875_10702.t8 6.1325
R18355 a_29875_10702.n1 a_29875_10702.t6 6.1325
R18356 a_29875_10702.n6 a_29875_10702.t0 4.70149
R18357 a_29875_10702.n8 a_29875_10702.n2 4.6302
R18358 a_29875_10702.n9 a_29875_10702.n8 2.85093
R18359 a_29875_10702.n4 a_29875_10702.t4 2.16717
R18360 a_29875_10702.n4 a_29875_10702.n3 2.16717
R18361 a_29875_10702.n9 a_29875_10702.t3 2.16717
R18362 a_29875_10702.n10 a_29875_10702.n9 2.16717
R18363 a_29875_10702.n7 a_29875_10702.n6 1.58582
R18364 a_29875_10702.n7 a_29875_10702.n4 1.24371
R18365 a_29875_10702.n8 a_29875_10702.n7 0.971051
R18366 a_42628_11460.t0 a_42628_11460.t1 12.9675
R18367 a_46528_12082.t0 a_46528_12082.t1 12.9675
R18368 a_46228_11460.t0 a_46228_11460.t1 12.9675
R18369 UP_INPUT.n0 UP_INPUT 6.382
R18370 UP_INPUT.n10 UP_INPUT.t0 5.81586
R18371 UP_INPUT.n6 UP_INPUT.n5 5.1005
R18372 UP_INPUT.n14 UP_INPUT.n7 5.1005
R18373 UP_INPUT.n12 UP_INPUT.n11 5.08021
R18374 UP_INPUT.n4 UP_INPUT.n3 4.6305
R18375 UP_INPUT.n10 UP_INPUT.n9 2.85093
R18376 UP_INPUT.n9 UP_INPUT.t3 2.16717
R18377 UP_INPUT.n9 UP_INPUT.n8 2.16717
R18378 UP_INPUT.n3 UP_INPUT.t6 1.9505
R18379 UP_INPUT.n3 UP_INPUT.n2 1.9505
R18380 UP_INPUT UP_INPUT.n0 1.71977
R18381 UP_INPUT.n0 UP_INPUT 0.852643
R18382 UP_INPUT.n16 UP_INPUT.n15 0.818177
R18383 UP_INPUT.n12 UP_INPUT.n10 0.644196
R18384 UP_INPUT.n13 UP_INPUT.n12 0.400713
R18385 UP_INPUT.n17 UP_INPUT.n1 0.368
R18386 UP_INPUT.n15 UP_INPUT.n14 0.248625
R18387 UP_INPUT.n15 UP_INPUT.n6 0.237703
R18388 UP_INPUT UP_INPUT.n17 0.06675
R18389 UP_INPUT.n14 UP_INPUT.n13 0.0502872
R18390 UP_INPUT.n6 UP_INPUT.n4 0.0318043
R18391 UP_INPUT.n17 UP_INPUT.n16 0.0013148
R18392 a_45328_10426.t0 a_45328_10426.t1 12.9675
R18393 a_45628_9804.t0 a_45628_9804.t1 12.9675
R18394 PFD_T2_0.Buffer_V_2_1.IN.n3 PFD_T2_0.Buffer_V_2_1.IN.t13 13.1405
R18395 PFD_T2_0.Buffer_V_2_1.IN.n4 PFD_T2_0.Buffer_V_2_1.IN.n3 12.4464
R18396 PFD_T2_0.Buffer_V_2_1.IN.n3 PFD_T2_0.Buffer_V_2_1.IN.t12 9.9285
R18397 PFD_T2_0.Buffer_V_2_1.IN.n22 PFD_T2_0.Buffer_V_2_1.IN.t11 9.7095
R18398 PFD_T2_0.Buffer_V_2_1.IN.n19 PFD_T2_0.Buffer_V_2_1.IN.n18 6.60246
R18399 PFD_T2_0.Buffer_V_2_1.IN.n1 PFD_T2_0.Buffer_V_2_1.IN.n5 4.5005
R18400 PFD_T2_0.Buffer_V_2_1.IN.n1 PFD_T2_0.Buffer_V_2_1.IN.n23 4.25602
R18401 PFD_T2_0.Buffer_V_2_1.IN.n1 PFD_T2_0.Buffer_V_2_1.IN.n2 4.22422
R18402 PFD_T2_0.Buffer_V_2_1.IN.n11 PFD_T2_0.Buffer_V_2_1.IN.t3 3.6405
R18403 PFD_T2_0.Buffer_V_2_1.IN.n11 PFD_T2_0.Buffer_V_2_1.IN.n10 3.6405
R18404 PFD_T2_0.Buffer_V_2_1.IN.n13 PFD_T2_0.Buffer_V_2_1.IN.t4 3.6405
R18405 PFD_T2_0.Buffer_V_2_1.IN.n13 PFD_T2_0.Buffer_V_2_1.IN.n12 3.6405
R18406 PFD_T2_0.Buffer_V_2_1.IN.n14 PFD_T2_0.Buffer_V_2_1.IN.n13 3.54941
R18407 PFD_T2_0.Buffer_V_2_1.IN.n17 PFD_T2_0.Buffer_V_2_1.IN.n16 3.33833
R18408 PFD_T2_0.Buffer_V_2_1.IN.n20 PFD_T2_0.Buffer_V_2_1.IN.n9 3.33833
R18409 PFD_T2_0.Buffer_V_2_1.IN.n16 PFD_T2_0.Buffer_V_2_1.IN.t0 3.2765
R18410 PFD_T2_0.Buffer_V_2_1.IN.n16 PFD_T2_0.Buffer_V_2_1.IN.n15 3.2765
R18411 PFD_T2_0.Buffer_V_2_1.IN.n9 PFD_T2_0.Buffer_V_2_1.IN.t8 3.2765
R18412 PFD_T2_0.Buffer_V_2_1.IN.n9 PFD_T2_0.Buffer_V_2_1.IN.n8 3.2765
R18413 PFD_T2_0.Buffer_V_2_1.IN.n0 PFD_T2_0.Buffer_V_2_1.IN.t9 3.2238
R18414 PFD_T2_0.Buffer_V_2_1.IN.n14 PFD_T2_0.Buffer_V_2_1.IN.n11 2.78441
R18415 PFD_T2_0.Buffer_V_2_1.IN.n7 PFD_T2_0.Buffer_V_2_1.IN.n6 1.9535
R18416 PFD_T2_0.Buffer_V_2_1.IN.n2 PFD_T2_0.Buffer_V_2_1.IN.n0 1.82827
R18417 PFD_T2_0.Buffer_V_2_1.IN.n0 PFD_T2_0.Buffer_V_2_1.IN.n7 1.37516
R18418 PFD_T2_0.Buffer_V_2_1.IN.n2 PFD_T2_0.Buffer_V_2_1.IN.n20 0.891537
R18419 PFD_T2_0.Buffer_V_2_1.IN.n23 PFD_T2_0.Buffer_V_2_1.IN.n21 0.729844
R18420 PFD_T2_0.Buffer_V_2_1.IN.n23 PFD_T2_0.Buffer_V_2_1.IN.n22 0.587069
R18421 PFD_T2_0.Buffer_V_2_1.IN.n19 PFD_T2_0.Buffer_V_2_1.IN.n17 0.524848
R18422 PFD_T2_0.Buffer_V_2_1.IN.n5 PFD_T2_0.Buffer_V_2_1.IN.n4 0.5115
R18423 PFD_T2_0.Buffer_V_2_1.IN.n17 PFD_T2_0.Buffer_V_2_1.IN.n14 0.358543
R18424 PFD_T2_0.Buffer_V_2_1.IN.n20 PFD_T2_0.Buffer_V_2_1.IN.n19 0.274413
R18425 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.Buffer_V_2_1.IN.n1 0.271564
R18426 a_43828_9598.t0 a_43828_9598.t1 12.9675
R18427 a_43528_8976.t0 a_43528_8976.t1 12.9675
R18428 VCTRL_IN.n3 VCTRL_IN.n2 5.81586
R18429 VCTRL_IN.n5 VCTRL_IN.t7 5.10208
R18430 VCTRL_IN.n8 VCTRL_IN.t5 5.10194
R18431 VCTRL_IN.n4 VCTRL_IN.t1 5.08021
R18432 VCTRL_IN.n8 VCTRL_IN.n7 4.66114
R18433 VCTRL_IN.n3 VCTRL_IN.n1 2.85093
R18434 VCTRL_IN.n1 VCTRL_IN.t2 2.16717
R18435 VCTRL_IN.n1 VCTRL_IN.n0 2.16717
R18436 VCTRL_IN.n7 VCTRL_IN.t4 1.9505
R18437 VCTRL_IN.n7 VCTRL_IN.n6 1.9505
R18438 VCTRL_IN.n4 VCTRL_IN.n3 0.644196
R18439 VCTRL_IN.n5 VCTRL_IN.n4 0.449473
R18440 VCTRL_IN.n9 VCTRL_IN.n8 0.21214
R18441 VCTRL_IN.n9 VCTRL_IN.n5 0.198571
R18442 VCTRL_IN VCTRL_IN.n9 0.0718949
R18443 a_42628_11254.t0 a_42628_11254.t1 12.9675
R18444 a_42628_10426.t0 a_42628_10426.t1 10.2205
R18445 a_46228_11254.t0 a_46228_11254.t1 12.9675
R18446 a_46528_10632.t0 a_46528_10632.t1 12.9675
R18447 a_23837_9553.n2 a_23837_9553.t3 6.64563
R18448 a_23837_9553.n2 a_23837_9553.t1 6.61433
R18449 a_23837_9553.n3 a_23837_9553.n1 3.36963
R18450 a_23837_9553.n4 a_23837_9553.n3 3.33833
R18451 a_23837_9553.n1 a_23837_9553.t5 3.2765
R18452 a_23837_9553.n1 a_23837_9553.n0 3.2765
R18453 a_23837_9553.n4 a_23837_9553.t0 3.2765
R18454 a_23837_9553.n5 a_23837_9553.n4 3.2765
R18455 a_23837_9553.n3 a_23837_9553.n2 0.781777
R18456 a_45028_9598.t0 a_45028_9598.t1 12.9675
R18457 a_45328_8976.t0 a_45328_8976.t1 12.9675
R18458 a_46528_8770.t0 a_46528_8770.t1 12.9675
R18459 a_43528_8770.t0 a_43528_8770.t1 12.9675
R18460 a_44716_1837.n3 a_44716_1837.t8 29.3691
R18461 a_44716_1837.n4 a_44716_1837.n3 21.9292
R18462 a_44716_1837.n5 a_44716_1837.n4 18.1271
R18463 a_44716_1837.n5 a_44716_1837.t9 11.2425
R18464 a_44716_1837.n8 a_44716_1837.n7 10.1038
R18465 a_44716_1837.n3 a_44716_1837.t6 6.1325
R18466 a_44716_1837.n4 a_44716_1837.t7 6.1325
R18467 a_44716_1837.n8 a_44716_1837.t0 4.70149
R18468 a_44716_1837.n6 a_44716_1837.n5 4.6302
R18469 a_44716_1837.n6 a_44716_1837.n2 2.85093
R18470 a_44716_1837.n2 a_44716_1837.t2 2.16717
R18471 a_44716_1837.n2 a_44716_1837.n1 2.16717
R18472 a_44716_1837.t5 a_44716_1837.n10 2.16717
R18473 a_44716_1837.n10 a_44716_1837.n0 2.16717
R18474 a_44716_1837.n9 a_44716_1837.n8 1.58618
R18475 a_44716_1837.n10 a_44716_1837.n9 1.24388
R18476 a_44716_1837.n9 a_44716_1837.n6 0.97169
R18477 a_43228_11460.t0 a_43228_11460.t1 12.9675
R18478 LF_OFFCHIP.n10 LF_OFFCHIP 8.48631
R18479 LF_OFFCHIP.n6 LF_OFFCHIP.n5 5.81586
R18480 LF_OFFCHIP.n8 LF_OFFCHIP.t7 5.10208
R18481 LF_OFFCHIP.n2 LF_OFFCHIP.t5 5.10195
R18482 LF_OFFCHIP.n7 LF_OFFCHIP.t0 5.08021
R18483 LF_OFFCHIP.n2 LF_OFFCHIP.n1 4.66211
R18484 LF_OFFCHIP.n6 LF_OFFCHIP.n4 2.85093
R18485 LF_OFFCHIP.n4 LF_OFFCHIP.t1 2.16717
R18486 LF_OFFCHIP.n4 LF_OFFCHIP.n3 2.16717
R18487 LF_OFFCHIP.n1 LF_OFFCHIP.t6 1.9505
R18488 LF_OFFCHIP.n1 LF_OFFCHIP.n0 1.9505
R18489 LF_OFFCHIP.n10 LF_OFFCHIP 1.59267
R18490 LF_OFFCHIP LF_OFFCHIP.n10 0.894244
R18491 LF_OFFCHIP.n7 LF_OFFCHIP.n6 0.644196
R18492 LF_OFFCHIP.n8 LF_OFFCHIP.n7 0.449473
R18493 LF_OFFCHIP.n9 LF_OFFCHIP.n2 0.212726
R18494 LF_OFFCHIP.n9 LF_OFFCHIP.n8 0.198082
R18495 LF_OFFCHIP LF_OFFCHIP.n9 0.0718702
R18496 a_41879_n196.n5 a_41879_n196.t8 29.2961
R18497 a_41879_n196.n6 a_41879_n196.n5 21.9292
R18498 a_41879_n196.n7 a_41879_n196.n6 18.1271
R18499 a_41879_n196.n7 a_41879_n196.t6 11.1695
R18500 a_41879_n196.n3 a_41879_n196.t0 10.2143
R18501 a_41879_n196.n5 a_41879_n196.t9 6.1325
R18502 a_41879_n196.n6 a_41879_n196.t7 6.1325
R18503 a_41879_n196.n3 a_41879_n196.n2 4.68517
R18504 a_41879_n196.n8 a_41879_n196.n7 4.6311
R18505 a_41879_n196.n10 a_41879_n196.n8 2.85093
R18506 a_41879_n196.n1 a_41879_n196.t2 2.16717
R18507 a_41879_n196.n1 a_41879_n196.n0 2.16717
R18508 a_41879_n196.t5 a_41879_n196.n10 2.16717
R18509 a_41879_n196.n10 a_41879_n196.n9 2.16717
R18510 a_41879_n196.n4 a_41879_n196.n3 1.58582
R18511 a_41879_n196.n4 a_41879_n196.n1 1.24371
R18512 a_41879_n196.n8 a_41879_n196.n4 0.971051
R18513 a_43228_11254.t0 a_43228_11254.t1 12.9675
R18514 a_44728_8770.t0 a_44728_8770.t1 12.9675
R18515 a_45028_8148.t0 a_45028_8148.t1 12.9675
R18516 a_18550_11273.n5 a_18550_11273.t8 29.3691
R18517 a_18550_11273.n6 a_18550_11273.n5 21.9292
R18518 a_18550_11273.n7 a_18550_11273.n6 18.1271
R18519 a_18550_11273.n7 a_18550_11273.t6 11.2425
R18520 a_18550_11273.n3 a_18550_11273.t1 10.2135
R18521 a_18550_11273.n5 a_18550_11273.t7 6.1325
R18522 a_18550_11273.n6 a_18550_11273.t9 6.1325
R18523 a_18550_11273.n3 a_18550_11273.n2 4.68398
R18524 a_18550_11273.n8 a_18550_11273.n7 4.6302
R18525 a_18550_11273.n9 a_18550_11273.n8 2.85093
R18526 a_18550_11273.n1 a_18550_11273.t3 2.16717
R18527 a_18550_11273.n1 a_18550_11273.n0 2.16717
R18528 a_18550_11273.n9 a_18550_11273.t2 2.16717
R18529 a_18550_11273.n10 a_18550_11273.n9 2.16717
R18530 a_18550_11273.n4 a_18550_11273.n3 1.58582
R18531 a_18550_11273.n4 a_18550_11273.n1 1.24371
R18532 a_18550_11273.n8 a_18550_11273.n4 0.971051
R18533 a_44128_12082.t0 a_44128_12082.t1 12.9675
R18534 a_25556_11637.n0 a_25556_11637.t5 24.1814
R18535 a_25556_11637.n1 a_25556_11637.t4 12.4835
R18536 a_25556_11637.n0 a_25556_11637.t3 8.6875
R18537 a_25556_11637.n2 a_25556_11637.t0 6.71215
R18538 a_25556_11637.n2 a_25556_11637.n1 4.46748
R18539 a_25556_11637.n3 a_25556_11637.t1 3.6405
R18540 a_25556_11637.n4 a_25556_11637.n3 3.6405
R18541 a_25556_11637.n3 a_25556_11637.n2 2.83724
R18542 a_25556_11637.n1 a_25556_11637.n0 1.8985
R18543 a_44128_10632.t0 a_44128_10632.t1 12.9675
R18544 a_46528_10426.t0 a_46528_10426.t1 12.9675
R18545 a_42928_10426.t0 a_42928_10426.t1 12.9675
R18546 a_43228_9804.t0 a_43228_9804.t1 12.9675
R18547 a_44728_8976.t0 a_44728_8976.t1 12.9675
R18548 a_46228_9598.t0 a_46228_9598.t1 12.9675
R18549 a_45928_8976.t0 a_45928_8976.t1 12.9675
R18550 a_45028_11460.t0 a_45028_11460.t1 12.9675
R18551 a_44428_8148.t0 a_44428_8148.t1 12.9675
R18552 a_45028_11254.t0 a_45028_11254.t1 12.9675
R18553 a_45928_12082.t0 a_45928_12082.t1 12.9675
R18554 a_42628_9804.t0 a_42628_9804.t1 12.9675
R18555 a_45928_10632.t0 a_45928_10632.t1 12.9675
R18556 a_44128_10426.t0 a_44128_10426.t1 12.9675
R18557 a_43828_9804.t0 a_43828_9804.t1 12.9675
R18558 a_45628_9598.t0 a_45628_9598.t1 12.9675
R18559 a_42928_12082.t0 a_42928_12082.t1 12.9675
R18560 a_42928_10632.t0 a_42928_10632.t1 12.9675
R18561 a_45328_8770.t0 a_45328_8770.t1 12.9675
R18562 a_46828_9598.t0 a_46828_9598.t1 10.2205
R18563 a_43528_10426.t0 a_43528_10426.t1 12.9675
R18564 a_45028_9804.t0 a_45028_9804.t1 12.9675
R18565 a_46528_8976.t0 a_46528_8976.t1 12.9675
R18566 a_43228_9598.t0 a_43228_9598.t1 12.9675
R18567 a_46228_8148.t0 a_46228_8148.t1 12.9675
R18568 a_46828_11254.t0 a_46828_11254.t1 10.2205
C0 DN_OUT VCTRL2 0.0165f
C1 VCO_DFF_C_0.OUTB A_MUX_0.Tr_Gate_1.CLK 0.00188f
C2 PFD_T2_0.FDIV PFD_T2_0.Buffer_V_2_0.IN 0.00808f
C3 VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT VDD 2.15f
C4 A_MUX_0.Tr_Gate_1.CLK VDD 1.93f
C5 A_MUX_1.Tr_Gate_1.CLK PFD_T2_0.FIN 0.425f
C6 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN m1_30034_1474# 0.00112f
C7 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 1.57f
C8 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.403f
C9 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.0179f
C10 PFD_T2_0.INV_mag_0.IN UP1 3.35e-19
C11 A_MUX_1.Tr_Gate_1.CLK S1 0.404f
C12 PFD_T2_0.Buffer_V_2_0.IN VDD 1.31f
C13 CP_1_0.VCTRL ITAIL 1.83f
C14 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 0.703f
C15 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCTRL2 0.0917f
C16 S5 ITAIL1 0.00468f
C17 ITAIL DN_OUT 0.00678f
C18 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.0107f
C19 PFD_T2_0.INV_mag_0.IN PFD_T2_0.FDIV 3.6e-22
C20 A_MUX_0.Tr_Gate_1.CLK VCO_DFF_C_0.VCTRL 0.422f
C21 DN_OUT S3 1.83f
C22 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.578f
C23 A_MUX_6.Tr_Gate_1.CLK RES_74k_1.P 0.49f
C24 VCO_DFF_C_0.VCO_C_0.OUTB S4 0.0152f
C25 RES_74k_1.M VDD 0.826f
C26 CP_1_0.VCTRL S4 0.0014f
C27 VCO_DFF_C_0.OUTB VCO_DFF_C_0.VCO_C_0.OUTB 0.725f
C28 RES_74k_1.P S5 8.5e-19
C29 CP_1_0.VCTRL VCO_DFF_C_0.OUTB 0.979f
C30 PFD_T2_0.FDIV S6 0.532f
C31 VCO_DFF_C_0.VCO_C_0.OUTB VDD 5.93f
C32 PFD_T2_0.Buffer_V_2_1.IN UP1 0.013f
C33 CP_1_0.VCTRL VDD 3.53f
C34 VDD DN_OUT 5.44f
C35 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_0.OUT 0.218f
C36 A_MUX_1.Tr_Gate_1.CLK A_MUX_2.Tr_Gate_1.CLK 0.00522f
C37 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 10.3f
C38 UP1 DN_INPUT 0.0798f
C39 PFD_T2_0.INV_mag_0.IN VDD 4.74f
C40 A_MUX_3.Tr_Gate_1.CLK UP1 0.491f
C41 PFD_T2_0.INV_mag_0.IN PRE_SCALAR 6.12e-20
C42 PFD_T2_0.INV_mag_0.OUT DN1 7.95e-19
C43 VDD S6 2.87f
C44 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.OUTB 0.0222f
C45 CP_1_0.VCTRL VCO_DFF_C_0.VCTRL 2.03f
C46 VCO_DFF_C_0.VCTRL DN_OUT 0.0605f
C47 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VDD 12.6f
C48 S3 DN_INPUT 1.24f
C49 S2 DN_OUT 0.012f
C50 PFD_T2_0.Buffer_V_2_1.IN VDD 1.18f
C51 PFD_T2_0.FIN PFD_T2_0.INV_mag_0.IN 0.151f
C52 PFD_T2_0.INV_mag_0.IN S2 0.0485f
C53 VDD DN_INPUT 1.13f
C54 S4 VCTRL_IN 0.548f
C55 PRE_SCALAR DN_INPUT 0.00844f
C56 VCO_DFF_C_0.OUTB VCTRL_IN 0.0234f
C57 PFD_T2_0.FIN S6 4.97e-19
C58 PFD_T2_0.INV_mag_1.IN PFD_T2_0.INV_mag_1.OUT 0.224f
C59 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.381f
C60 A_MUX_3.Tr_Gate_1.CLK VDD 1.86f
C61 VCO_DFF_C_0.OUT OUTB 0.0034f
C62 VDD VCTRL_IN 0.112f
C63 UP1 UP_OUT 1.25f
C64 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 1.27f
C65 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 3.46e-19
C66 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 3.19f
C67 PFD_T2_0.FDIV DIV_OUT 1.29f
C68 PFD_T2_0.FIN PFD_T2_0.Buffer_V_2_1.IN 0.00669f
C69 S1 S6 0.00521f
C70 PFD_T2_0.INV_mag_1.OUT DN1 0.0191f
C71 PFD_T2_0.Buffer_V_2_1.IN S2 0.0215f
C72 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCTRL2 0.0273f
C73 DIV_OUT S3 0.0272f
C74 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 0.382f
C75 ITAIL UP_OUT 1.96f
C76 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.39f
C77 UP_OUT S3 0.361f
C78 S2 DN_INPUT 0.984f
C79 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.Buffer_V_2_0.IN 0.187f
C80 VCO_DFF_C_0.VCTRL VCTRL_IN 1.25f
C81 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 10.4f
C82 A_MUX_3.Tr_Gate_1.CLK S2 0.415f
C83 VDD LF_OFFCHIP 0.519f
C84 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUT 1.19f
C85 VCO_DFF_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.0234f
C86 VDD DIV_OUT 0.404f
C87 A_MUX_2.Tr_Gate_1.CLK S6 0.403f
C88 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.4f
C89 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 1.2f
C90 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VDD 2.59f
C91 VDD UP_OUT 3.43f
C92 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 0.00102f
C93 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.00409f
C94 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 5.91e-19
C95 VCO_DFF_C_0.OUTB VCO_DFF_C_0.OUT 0.487f
C96 VDD F_IN 0.112f
C97 VCO_DFF_C_0.OUT VDD 5.58f
C98 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_0.OUT 0.318f
C99 A_MUX_6.Tr_Gate_1.CLK CP_1_0.VCTRL 0.422f
C100 CP_1_0.VCTRL S5 0.504f
C101 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.652f
C102 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VDD 2.16f
C103 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VDD 0.893f
C104 S2 UP_OUT 0.547f
C105 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.Buffer_V_2_0.IN 0.0183f
C106 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.OUT 0.00184f
C107 PFD_T2_0.FIN F_IN 1.25f
C108 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN m1_30034_1474# 0.103f
C109 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCTRL2 0.108f
C110 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.618f
C111 VCO_DFF_C_0.VCO_C_0.OUT VCO_DFF_C_0.VCO_C_0.OUTB 1.64f
C112 PFD_T2_0.INV_mag_0.OUT DN_INPUT 0.228f
C113 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.13f
C114 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT 0.02f
C115 S1 F_IN 0.612f
C116 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 0.674f
C117 A_MUX_3.Tr_Gate_1.CLK PFD_T2_0.INV_mag_0.OUT 5.43e-20
C118 S3 VCTRL2 0.336f
C119 VCO_DFF_C_0.OUTB OUTB 0.0149f
C120 A_MUX_2.Tr_Gate_1.CLK DIV_OUT 0.496f
C121 VDD OUTB 14.7f
C122 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 1.21f
C123 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_1.OUT 0.404f
C124 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 0.488f
C125 VDD VCTRL2 1.21f
C126 VDD UP1 0.648f
C127 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN VDD 0.921f
C128 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.OUT 0.135f
C129 PFD_T2_0.FDIV VDD 2.12f
C130 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VDD 14.9f
C131 VCO_DFF_C_0.VCTRL VCTRL2 0.283f
C132 PFD_T2_0.INV_mag_1.OUT DN_INPUT 0.293f
C133 VCO_DFF_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK 0.493f
C134 PFD_T2_0.INV_mag_1.IN DN1 2.85e-19
C135 VDD ITAIL 6.22f
C136 VDD S3 3.84f
C137 S5 LF_OFFCHIP 5.4f
C138 RES_74k_1.M m1_53133_19897# 0.782f
C139 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VDD 3.8f
C140 A_MUX_3.Tr_Gate_1.CLK PFD_T2_0.INV_mag_1.OUT 0.00126f
C141 VCO_DFF_C_0.OUTB S4 0.0286f
C142 VDD S4 2.92f
C143 UP1 S2 0.0962f
C144 RES_74k_1.P A_MUX_0.Tr_Gate_1.CLK 0.00665f
C145 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 1.21f
C146 VCO_DFF_C_0.OUTB VDD 2.27f
C147 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN m1_33892_1807# 0.00112f
C148 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 1.63f
C149 VDD PRE_SCALAR 0.135f
C150 PFD_T2_0.FIN PFD_T2_0.FDIV 0.284f
C151 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 0.624f
C152 A_MUX_4.Tr_Gate_1.CLK DN1 0.491f
C153 VCO_DFF_C_0.OUT VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.0191f
C154 VCO_DFF_C_0.VCTRL S3 0.608f
C155 S2 S3 0.00929f
C156 PFD_T2_0.FDIV S1 9.35e-19
C157 VCO_DFF_C_0.VCTRL S4 0.523f
C158 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT 1.64f
C159 VCO_DFF_C_0.OUTB VCO_DFF_C_0.VCTRL 0.0294f
C160 PFD_T2_0.INV_mag_1.OUT UP_OUT 0.0705f
C161 CP_1_0.VCTRL ITAIL1 1.65f
C162 VCO_DFF_C_0.VCTRL VDD 13f
C163 PFD_T2_0.FIN VDD 1.93f
C164 DN_OUT ITAIL1 0.00354f
C165 RES_74k_1.P RES_74k_1.M 0.425f
C166 VDD S2 4.28f
C167 PFD_T2_0.FIN PRE_SCALAR 1.31f
C168 PRE_SCALAR S2 0.173f
C169 CP_1_0.VCTRL RES_74k_1.P 2.14f
C170 PFD_T2_0.FDIV A_MUX_2.Tr_Gate_1.CLK 0.43f
C171 PFD_T2_0.INV_mag_1.IN PFD_T2_0.Buffer_V_2_0.IN 0.595f
C172 VDD S1 2.8f
C173 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.00342f
C174 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 3.46e-19
C175 S1 PRE_SCALAR 0.0855f
C176 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUT 0.385f
C177 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 3.61e-20
C178 PFD_T2_0.Buffer_V_2_0.IN DN1 0.0162f
C179 A_MUX_2.Tr_Gate_1.CLK VDD 1.98f
C180 DN_OUT UP_INPUT 1.06f
C181 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCTRL2 0.198f
C182 PFD_T2_0.INV_mag_0.OUT PFD_T2_0.FDIV 0.0689f
C183 PFD_T2_0.FIN S1 0.528f
C184 PFD_T2_0.INV_mag_0.IN PFD_T2_0.INV_mag_1.IN 1.33f
C185 DN_OUT DN1 1.25f
C186 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.IN 7.97e-19
C187 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.765f
C188 A_MUX_4.Tr_Gate_1.CLK DN_OUT 0.424f
C189 RES_74k_1.P VCTRL_IN 4.84e-20
C190 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_2.IN 0.915f
C191 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCTRL2 0.344f
C192 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.915f
C193 PFD_T2_0.FIN A_MUX_2.Tr_Gate_1.CLK 3.91e-19
C194 VCO_DFF_C_0.VCO_C_0.OUT VCTRL2 0.0145f
C195 PFD_T2_0.INV_mag_0.OUT VDD 0.675f
C196 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_1.IN 0.0388f
C197 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.306f
C198 A_MUX_1.Tr_Gate_1.CLK PFD_T2_0.INV_mag_0.IN 7.22e-21
C199 PFD_T2_0.INV_mag_1.IN DN_INPUT 0.124f
C200 PFD_T2_0.INV_mag_1.OUT UP1 0.0288f
C201 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.419f
C202 A_MUX_6.Tr_Gate_1.CLK VDD 2.1f
C203 LF_OFFCHIP ITAIL1 3.17f
C204 VCO_DFF_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT 0.00852f
C205 VDD S5 3.76f
C206 CP_1_0.VCTRL A_MUX_0.Tr_Gate_1.CLK 0.49f
C207 PFD_T2_0.INV_mag_1.IN A_MUX_3.Tr_Gate_1.CLK 6.92e-19
C208 UP_INPUT DN_INPUT 0.86f
C209 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.OUT VDD 2.87f
C210 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VDD 0.795f
C211 UP_OUT ITAIL1 0.0883f
C212 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.OUT 9.22e-19
C213 DN1 DN_INPUT 0.466f
C214 PFD_T2_0.FIN PFD_T2_0.INV_mag_0.OUT 0.0528f
C215 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN S3 1.8e-19
C216 A_MUX_3.Tr_Gate_1.CLK DN1 8.25e-20
C217 VCO_DFF_C_0.OUT OUT 0.0173f
C218 A_MUX_4.Tr_Gate_1.CLK DN_INPUT 0.0194f
C219 A_MUX_3.Tr_Gate_1.CLK A_MUX_4.Tr_Gate_1.CLK 0.00466f
C220 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VDD 12.5f
C221 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.389f
C222 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT 0.00912f
C223 VCO_DFF_C_0.VCO_C_0.OUT VDD 0.723f
C224 PFD_T2_0.INV_mag_1.OUT VDD 0.705f
C225 PFD_T2_0.INV_mag_0.IN PFD_T2_0.Buffer_V_2_0.IN 0.0412f
C226 PFD_T2_0.INV_mag_1.IN UP_OUT 7.85e-19
C227 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN m1_33892_1807# 0.106f
C228 CP_1_0.VCTRL DN_OUT 1.07e-19
C229 UP_OUT UP_INPUT 1.36f
C230 UP_OUT DN1 0.0248f
C231 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 3.31f
C232 VCO_DFF_C_0.VCTRL VCO_DFF_C_0.VCO_C_0.OUT 0.0471f
C233 PFD_T2_0.INV_mag_1.OUT S2 0.0234f
C234 A_MUX_4.Tr_Gate_1.CLK UP_OUT 0.00217f
C235 m1_33892_1807# VDD 0.0434f
C236 PFD_T2_0.Buffer_V_2_0.IN DN_INPUT 0.0128f
C237 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.348f
C238 m1_30034_1474# VDD 0.0163f
C239 DN_OUT DN_INPUT 1.3f
C240 PFD_T2_0.Buffer_V_2_1.IN PFD_T2_0.INV_mag_0.IN 0.428f
C241 VCO_DFF_C_0.VCO_C_0.OUTB VCTRL_IN 0.00272f
C242 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 0.546f
C243 VCO_DFF_C_0.VCTRL m1_33892_1807# 5.46e-20
C244 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 0.00756f
C245 PFD_T2_0.INV_mag_0.IN DN_INPUT 0.0654f
C246 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_0.IN 0.388f
C247 VCO_DFF_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN 1.27f
C248 PFD_T2_0.INV_mag_0.IN A_MUX_3.Tr_Gate_1.CLK 2.18e-19
C249 ITAIL ITAIL1 2.7f
C250 VCO_DFF_C_0.VCTRL m1_30034_1474# 0.0168f
C251 VCO_DFF_C_0.DFF_3_mag_0.INV_2_1.IN VDD 2.74f
C252 A_MUX_6.Tr_Gate_1.CLK S5 0.397f
C253 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 0.0108f
C254 PFD_T2_0.INV_mag_1.IN UP1 2.09e-20
C255 VDD OUT 14.7f
C256 PFD_T2_0.Buffer_V_2_1.IN DN_INPUT 0.0174f
C257 VDD ITAIL1 1.02f
C258 CP_1_0.VCTRL LF_OFFCHIP 1.27f
C259 RES_74k_1.P S4 0.0103f
C260 PFD_T2_0.INV_mag_1.OUT PFD_T2_0.INV_mag_0.OUT 0.479f
C261 RES_74k_1.P VCO_DFF_C_0.OUTB 0.0107f
C262 VCO_DFF_C_0.VCO_C_0.OUTB VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.OUT 0.403f
C263 CP_1_0.VCTRL UP_OUT 0.00287f
C264 PFD_T2_0.INV_mag_1.IN PFD_T2_0.FDIV 0.161f
C265 RES_74k_1.P VDD 22.6f
C266 UP_OUT DN_OUT 2.18f
C267 A_MUX_3.Tr_Gate_1.CLK DN_INPUT 0.0129f
C268 VCO_DFF_C_0.VCO_C_0.INV_2_5.OUT VCO_DFF_C_0.VCO_C_0.INV_2_5.IN 0.391f
C269 PFD_T2_0.INV_mag_0.IN UP_OUT 9.06e-20
C270 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VCTRL2 0.321f
C271 ITAIL UP_INPUT 7.63e-19
C272 VCO_DFF_C_0.OUT VCO_DFF_C_0.VCO_C_0.OUTB 0.00703f
C273 S6 DIV_OUT 0.0112f
C274 VCO_DFF_C_0.VCO_C_0.INV_2_4.IN VCO_DFF_C_0.VCO_C_0.OUTB 0.00204f
C275 PFD_T2_0.INV_mag_1.IN VDD 5.09f
C276 DN1 S3 8.76e-19
C277 RES_74k_1.P VCO_DFF_C_0.VCTRL 0.105f
C278 A_MUX_1.Tr_Gate_1.CLK PFD_T2_0.FDIV 0.00277f
C279 VDD UP_INPUT 0.798f
C280 PRE_SCALAR UP_INPUT 0.0156f
C281 A_MUX_4.Tr_Gate_1.CLK S3 0.404f
C282 VCO_DFF_C_0.VCO_C_0.INV_2_5.IN VCO_DFF_C_0.VCO_C_0.OUT 0.791f
C283 VDD DN1 0.709f
C284 VCO_DFF_C_0.DFF_3_mag_0.Tr_Gate_0.CLK VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT 0.00977f
C285 UP_OUT DN_INPUT 0.101f
C286 VCO_DFF_C_0.VCO_C_0.INV_2_2.IN VCO_DFF_C_0.VCO_C_0.INV_2_3.OUT 7.5e-19
C287 A_MUX_4.Tr_Gate_1.CLK VDD 1.91f
C288 A_MUX_3.Tr_Gate_1.CLK UP_OUT 0.424f
C289 PFD_T2_0.FIN PFD_T2_0.INV_mag_1.IN 0.00687f
C290 A_MUX_1.Tr_Gate_1.CLK VDD 1.86f
C291 VCO_DFF_C_0.VCO_C_0.INV_2_3.IN VCO_DFF_C_0.VCO_C_0.INV_2_4.IN 2.23e-19
C292 VCO_DFF_C_0.DFF_3_mag_0.INV_2_5.OUT VDD 0.958f
C293 VCO_DFF_C_0.VCO_C_0.INV_2_0.OUT VCO_DFF_C_0.VCO_C_0.INV_2_3.IN 0.809f
C294 PFD_T2_0.INV_mag_1.IN S2 0.00145f
C295 A_MUX_1.Tr_Gate_1.CLK PRE_SCALAR 0.502f
C296 VCO_DFF_C_0.VCO_C_0.INV_2_0.IN VDD 14.8f
C297 S2 UP_INPUT 0.934f
C298 VCO_DFF_C_0.VCO_C_0.OUTB VCTRL2 0.00407f
C299 A_MUX_0.Tr_Gate_1.CLK S4 0.403f
.ends

