magic
tech gf180mcuC
magscale 1 10
timestamp 1693477706
<< nwell >>
rect -36 634 390 733
<< psubdiff >>
rect -231 828 589 842
rect -231 826 -101 828
rect -231 776 -218 826
rect -168 778 -101 826
rect -51 778 24 828
rect 74 778 149 828
rect 199 778 274 828
rect 324 778 399 828
rect 449 778 524 828
rect 574 778 589 828
rect -168 776 589 778
rect -231 764 589 776
rect -231 691 -149 764
rect -231 641 -218 691
rect -168 641 -149 691
rect -231 556 -149 641
rect 508 685 589 764
rect 508 635 526 685
rect 576 635 589 685
rect -231 506 -218 556
rect -168 506 -149 556
rect -231 421 -149 506
rect 508 550 589 635
rect 508 500 526 550
rect 576 500 589 550
rect -231 371 -218 421
rect -168 371 -149 421
rect -231 286 -149 371
rect 508 415 589 500
rect 508 365 526 415
rect 576 365 589 415
rect -231 236 -218 286
rect -168 236 -149 286
rect -231 151 -149 236
rect -231 101 -218 151
rect -168 101 -149 151
rect -231 23 -149 101
rect 508 280 589 365
rect 508 230 526 280
rect 576 230 589 280
rect 508 145 589 230
rect 508 95 526 145
rect 576 95 589 145
rect 508 23 589 95
rect -231 10 589 23
rect -231 -40 -214 10
rect -164 -40 -89 10
rect -39 -40 36 10
rect 86 -40 161 10
rect 211 -40 286 10
rect 336 -40 411 10
rect 461 -40 526 10
rect 576 -40 589 10
rect -231 -55 589 -40
<< nsubdiff >>
rect 13 681 330 694
rect 13 635 29 681
rect 75 635 149 681
rect 195 635 269 681
rect 315 635 330 681
rect 13 618 330 635
<< psubdiffcont >>
rect -218 776 -168 826
rect -101 778 -51 828
rect 24 778 74 828
rect 149 778 199 828
rect 274 778 324 828
rect 399 778 449 828
rect 524 778 574 828
rect -218 641 -168 691
rect 526 635 576 685
rect -218 506 -168 556
rect 526 500 576 550
rect -218 371 -168 421
rect 526 365 576 415
rect -218 236 -168 286
rect -218 101 -168 151
rect 526 230 576 280
rect 526 95 576 145
rect -214 -40 -164 10
rect -89 -40 -39 10
rect 36 -40 86 10
rect 161 -40 211 10
rect 286 -40 336 10
rect 411 -40 461 10
rect 526 -40 576 10
<< nsubdiffcont >>
rect 29 635 75 681
rect 149 635 195 681
rect 269 635 315 681
<< polysilicon >>
rect 142 423 212 436
rect 80 408 212 423
rect 80 342 95 408
rect 152 342 212 408
rect 80 329 212 342
rect 142 302 212 329
<< polycontact >>
rect 95 342 152 408
<< metal1 >>
rect -231 828 589 842
rect -231 826 -101 828
rect -231 776 -218 826
rect -168 778 -101 826
rect -51 778 24 828
rect 74 778 149 828
rect 199 778 274 828
rect 324 778 399 828
rect 449 778 524 828
rect 574 778 589 828
rect -168 776 589 778
rect -231 764 589 776
rect -231 691 -149 764
rect -231 641 -218 691
rect -168 641 -149 691
rect -231 556 -149 641
rect 13 681 330 694
rect 13 635 29 681
rect 75 635 149 681
rect 195 635 269 681
rect 315 635 330 681
rect 13 618 330 635
rect 508 685 589 764
rect 508 635 526 685
rect 576 635 589 685
rect -231 506 -218 556
rect -168 506 -149 556
rect -231 421 -149 506
rect 63 492 120 618
rect 508 550 589 635
rect -231 371 -218 421
rect -168 371 -149 421
rect 95 408 163 420
rect -231 286 -149 371
rect -40 342 95 389
rect 152 342 163 408
rect -40 330 163 342
rect -231 236 -218 286
rect -168 236 -149 286
rect 241 244 302 505
rect 508 500 526 550
rect 576 500 589 550
rect 508 415 589 500
rect 508 365 526 415
rect 576 365 589 415
rect 508 280 589 365
rect -231 151 -149 236
rect 508 230 526 280
rect 576 230 589 280
rect -231 101 -218 151
rect -168 101 -149 151
rect -231 23 -149 101
rect 66 23 113 158
rect 508 145 589 230
rect 508 95 526 145
rect 576 95 589 145
rect 508 23 589 95
rect -231 10 589 23
rect -231 -40 -214 10
rect -164 -40 -89 10
rect -39 -40 36 10
rect 86 -40 161 10
rect 211 -40 286 10
rect 336 -40 411 10
rect 461 -40 526 10
rect 576 -40 589 10
rect -231 -55 589 -40
use nmos_3p3_AQSZEK  nmos_3p3_AQSZEK_0
timestamp 1693477706
transform 1 0 177 0 1 188
box -147 -138 147 138
use pmos_3p3_HBGRPK  pmos_3p3_HBGRPK_0
timestamp 1693477706
transform 1 0 177 0 1 515
box -213 -166 213 166
<< labels >>
flabel metal1 112 662 112 662 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal1 -6 353 -6 353 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 273 357 273 357 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 88 84 88 84 0 FreeSans 320 0 0 0 VSS
port 3 nsew
<< end >>
