magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2083 -2083 5677 8020
<< isosubstrate >>
rect -83 -83 3677 6020
<< nwell >>
rect 173 3038 3421 3147
rect 173 2098 1171 3038
<< psubdiff >>
rect 2577 2630 3594 2720
rect 2577 1960 2667 2630
rect 3504 2440 3594 2630
rect 0 1876 2667 1960
rect 90 1870 2667 1876
<< mvpsubdiff >>
rect 247 3267 1295 5667
<< polysilicon >>
rect 335 3089 475 3223
rect 579 3089 719 3223
rect 335 3005 719 3089
rect 823 3089 963 3223
rect 1067 3089 1207 3223
rect 823 3005 1207 3089
rect 1483 2911 1623 3223
rect 1727 2911 1867 3223
rect 1971 2911 2111 3223
rect 2387 3207 2527 3223
rect 2631 3207 2771 3223
rect 2875 3207 3015 3223
rect 3119 3207 3259 3223
rect 2387 3123 3259 3207
rect 823 2144 963 2244
rect 3119 2272 3259 2450
rect 335 1530 1207 1692
rect 335 1514 475 1530
rect 579 1514 719 1530
rect 823 1514 963 1530
rect 1067 1514 1207 1530
rect 1311 1514 1451 1692
rect 1555 1514 1695 1692
rect 1971 1514 2111 1692
rect 2215 1530 2599 1692
rect 2215 1514 2355 1530
rect 2459 1514 2599 1530
rect 2875 1530 3259 1692
rect 2875 1514 3015 1530
rect 3119 1514 3259 1530
<< metal1 >>
rect 79 5858 165 5926
rect 245 3217 321 5667
rect 489 3267 565 5926
rect 733 3217 809 5667
rect 977 3267 1053 5667
rect 1221 3217 1297 5667
rect 245 3141 1297 3217
rect 367 1522 443 3081
rect 489 2713 1053 2789
rect 489 2528 565 2713
rect 1221 2528 1297 3141
rect 1393 3005 1469 5667
rect 1637 3217 1713 5667
rect 1881 3267 1957 5926
rect 2125 3217 2201 5667
rect 2297 3267 2373 5926
rect 1637 3141 2201 3217
rect 1515 2652 1591 3081
rect 489 2288 794 2528
rect 977 2452 1297 2528
rect 1343 2576 1591 2652
rect 79 11 165 79
rect 245 11 321 1470
rect 489 270 565 2288
rect 733 11 809 2220
rect 977 270 1053 2452
rect 1099 1522 1175 2110
rect 1343 1522 1419 2576
rect 1637 2494 1713 2908
rect 1465 2418 1713 2494
rect 1221 11 1297 1470
rect 1465 212 1541 2418
rect 1759 2350 1835 3081
rect 1587 2274 1835 2350
rect 1587 1522 1663 2274
rect 1709 270 1785 2110
rect 1881 2034 1957 3141
rect 2003 1522 2079 3081
rect 2529 2945 2629 5667
rect 2785 3267 2861 5926
rect 2695 3005 2951 3199
rect 3017 3105 3117 5667
rect 3273 3267 3349 5926
rect 3429 5858 3515 5926
rect 3017 3005 3373 3105
rect 2529 2845 3105 2945
rect 2588 2613 2656 2641
rect 2588 1953 2656 1988
rect 2125 1877 2656 1953
rect 1881 212 1957 1470
rect 2125 270 2201 1877
rect 3029 1824 3105 2845
rect 2369 1748 3105 1824
rect 2247 212 2323 1684
rect 2369 270 2445 1748
rect 1465 136 2323 212
rect 2613 11 2689 1470
rect 2773 219 2873 1470
rect 3029 270 3105 1748
rect 3273 219 3373 3005
rect 3445 2641 3583 2709
rect 3515 2617 3583 2641
rect 2773 129 3373 219
rect 3429 11 3515 79
<< metal2 >>
rect 977 2713 1053 3447
rect 1393 3005 2951 3081
rect 3273 2460 3349 3497
rect 3151 2280 3349 2460
rect 1099 2034 1957 2110
rect 2268 1877 3549 1953
use M1_NWELL_CDNS_40661953145230  M1_NWELL_CDNS_40661953145230_0
timestamp 1713338890
transform 1 0 1797 0 1 5892
box -1726 -128 1726 128
use M1_NWELL_CDNS_40661953145231  M1_NWELL_CDNS_40661953145231_0
timestamp 1713338890
transform 1 0 3549 0 1 4529
box -128 -1491 128 1491
use M1_NWELL_CDNS_40661953145236  M1_NWELL_CDNS_40661953145236_0
timestamp 1713338890
transform 1 0 45 0 1 4059
box -128 -1961 128 1961
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_0
timestamp 1713338890
transform 0 -1 405 1 0 1603
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_1
timestamp 1713338890
transform 1 0 846 0 1 2186
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_2
timestamp 1713338890
transform 0 -1 1625 1 0 1603
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_3
timestamp 1713338890
transform 0 -1 1137 1 0 1603
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_4
timestamp 1713338890
transform 0 -1 1381 1 0 1603
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_5
timestamp 1713338890
transform 0 -1 1553 -1 0 3000
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_6
timestamp 1713338890
transform 0 -1 1797 -1 0 3000
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_7
timestamp 1713338890
transform 0 -1 2285 1 0 1603
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_8
timestamp 1713338890
transform 0 -1 2041 1 0 1603
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_9
timestamp 1713338890
transform 0 -1 2041 -1 0 3000
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_10
timestamp 1713338890
transform 0 -1 2945 1 0 1603
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165346  M1_POLY2_CDNS_69033583165346_11
timestamp 1713338890
transform 0 -1 3189 1 0 2361
box -89 -42 89 42
use M1_POLY2_CDNS_69033583165623  M1_POLY2_CDNS_69033583165623_0
timestamp 1713338890
transform 1 0 533 0 -1 3047
box -136 -42 136 42
use M1_POLY2_CDNS_69033583165623  M1_POLY2_CDNS_69033583165623_1
timestamp 1713338890
transform 1 0 1023 0 -1 3047
box -136 -42 136 42
use M1_POLY2_CDNS_69033583165623  M1_POLY2_CDNS_69033583165623_2
timestamp 1713338890
transform -1 0 2823 0 -1 3165
box -136 -42 136 42
use M1_PSUB_CDNS_6903358316545  M1_PSUB_CDNS_6903358316545_0
timestamp 1713338890
transform 1 0 2622 0 1 2297
box -45 -327 45 327
use M1_PSUB_CDNS_69033583165621  M1_PSUB_CDNS_69033583165621_0
timestamp 1713338890
transform 1 0 2434 0 1 1915
box -233 -45 233 45
use M1_PSUB_CDNS_69033583165624  M1_PSUB_CDNS_69033583165624_0
timestamp 1713338890
transform 1 0 45 0 1 938
box -45 -938 45 938
use M1_PSUB_CDNS_69033583165625  M1_PSUB_CDNS_69033583165625_0
timestamp 1713338890
transform 1 0 771 0 1 1915
box -139 -45 139 45
use M1_PSUB_CDNS_69033583165626  M1_PSUB_CDNS_69033583165626_0
timestamp 1713338890
transform 1 0 3549 0 1 1314
box -45 -1314 45 1314
use M1_PSUB_CDNS_69033583165627  M1_PSUB_CDNS_69033583165627_0
timestamp 1713338890
transform 1 0 2763 0 1 2675
box -186 -45 186 45
use M1_PSUB_CDNS_69033583165628  M1_PSUB_CDNS_69033583165628_0
timestamp 1713338890
transform 1 0 1797 0 1 45
box -1643 -45 1643 45
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_0
timestamp 1713338890
transform 1 0 869 0 1 2991
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_1
timestamp 1713338890
transform 1 0 1015 0 1 2803
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_2
timestamp 1713338890
transform 1 0 1431 0 1 3095
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_3
timestamp 1713338890
transform 1 0 1137 0 1 2124
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_4
timestamp 1713338890
transform 1 0 1675 0 1 2991
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_5
timestamp 1713338890
transform 0 -1 1833 1 0 2072
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_6
timestamp 1713338890
transform 1 0 2945 0 1 1612
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_7
timestamp 1713338890
transform 0 -1 2823 1 0 3043
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_8
timestamp 1713338890
transform 1 0 3189 0 1 2370
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_9
timestamp 1713338890
transform 1 0 1015 0 1 3357
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_10
timestamp 1713338890
transform 1 0 3311 0 1 3407
box -38 -90 38 90
use M2_M1_CDNS_69033583165575  M2_M1_CDNS_69033583165575_0
timestamp 1713338890
transform 1 0 2462 0 1 1915
box -194 -38 194 38
use nmos_6p0_CDNS_4066195314514  nmos_6p0_CDNS_4066195314514_0
timestamp 1713338890
transform 1 0 3119 0 1 1988
box -88 -44 228 284
use nmos_6p0_CDNS_4066195314518  nmos_6p0_CDNS_4066195314518_0
timestamp 1713338890
transform -1 0 1207 0 1 270
box -88 -44 472 1244
use nmos_6p0_CDNS_4066195314518  nmos_6p0_CDNS_4066195314518_1
timestamp 1713338890
transform -1 0 2599 0 1 270
box -88 -44 472 1244
use nmos_6p0_CDNS_4066195314519  nmos_6p0_CDNS_4066195314519_0
timestamp 1713338890
transform -1 0 1695 0 1 270
box -88 -44 228 1244
use nmos_6p0_CDNS_4066195314519  nmos_6p0_CDNS_4066195314519_1
timestamp 1713338890
transform -1 0 1451 0 1 270
box -88 -44 228 1244
use nmos_6p0_CDNS_4066195314519  nmos_6p0_CDNS_4066195314519_2
timestamp 1713338890
transform -1 0 2111 0 1 270
box -88 -44 228 1244
use nmos_6p0_CDNS_4066195314520  nmos_6p0_CDNS_4066195314520_0
timestamp 1713338890
transform -1 0 719 0 1 270
box -88 -44 472 1244
use nmos_6p0_CDNS_4066195314520  nmos_6p0_CDNS_4066195314520_1
timestamp 1713338890
transform -1 0 3259 0 -1 1470
box -88 -44 472 1244
use pmos_6p0_CDNS_4066195314515  pmos_6p0_CDNS_4066195314515_0
timestamp 1713338890
transform -1 0 1867 0 1 3267
box -208 -120 348 2520
use pmos_6p0_CDNS_4066195314515  pmos_6p0_CDNS_4066195314515_1
timestamp 1713338890
transform -1 0 2111 0 1 3267
box -208 -120 348 2520
use pmos_6p0_CDNS_4066195314515  pmos_6p0_CDNS_4066195314515_2
timestamp 1713338890
transform -1 0 1623 0 1 3267
box -208 -120 348 2520
use pmos_6p0_CDNS_4066195314516  pmos_6p0_CDNS_4066195314516_0
timestamp 1713338890
transform 1 0 335 0 1 3267
box -208 -120 592 2520
use pmos_6p0_CDNS_4066195314516  pmos_6p0_CDNS_4066195314516_1
timestamp 1713338890
transform 1 0 2875 0 1 3267
box -208 -120 592 2520
use pmos_6p0_CDNS_4066195314516  pmos_6p0_CDNS_4066195314516_2
timestamp 1713338890
transform 1 0 2387 0 1 3267
box -208 -120 592 2520
use pmos_6p0_CDNS_4066195314517  pmos_6p0_CDNS_4066195314517_0
timestamp 1713338890
transform -1 0 963 0 1 2288
box -208 -120 348 360
use pmos_6p0_CDNS_4066195314521  pmos_6p0_CDNS_4066195314521_0
timestamp 1713338890
transform -1 0 1207 0 -1 5667
box -208 -120 512 2520
<< labels >>
rlabel metal1 s 1632 1726 1632 1726 4 EN
port 1 nsew
rlabel metal1 s 3066 5296 3066 5296 4 PDRIVE_X
port 2 nsew
rlabel metal1 s 2580 5278 2580 5278 4 PDRIVE_Y
port 3 nsew
rlabel metal1 s 772 5265 772 5265 4 NDRIVE_Y
port 4 nsew
rlabel metal1 s 345 5891 345 5891 4 DVDD
port 5 nsew
rlabel metal1 s 2042 1726 2042 1726 4 A
port 6 nsew
rlabel metal1 s 284 47 284 47 4 DVSS
port 7 nsew
rlabel metal1 s 1390 1726 1390 1726 4 ENB
port 8 nsew
rlabel metal1 s 1015 5270 1015 5270 4 NDRIVE_X
port 9 nsew
rlabel metal2 s 2947 1602 2947 1602 4 SLB
port 10 nsew
rlabel metal2 s 869 3046 869 3046 4 SL
port 11 nsew
<< end >>
