magic
tech gf180mcuC
magscale 1 10
timestamp 1693543231
<< nwell >>
rect -2162 -230 2162 230
<< pmos >>
rect -1988 -100 -1888 100
rect -1784 -100 -1684 100
rect -1580 -100 -1480 100
rect -1376 -100 -1276 100
rect -1172 -100 -1072 100
rect -968 -100 -868 100
rect -764 -100 -664 100
rect -560 -100 -460 100
rect -356 -100 -256 100
rect -152 -100 -52 100
rect 52 -100 152 100
rect 256 -100 356 100
rect 460 -100 560 100
rect 664 -100 764 100
rect 868 -100 968 100
rect 1072 -100 1172 100
rect 1276 -100 1376 100
rect 1480 -100 1580 100
rect 1684 -100 1784 100
rect 1888 -100 1988 100
<< pdiff >>
rect -2076 87 -1988 100
rect -2076 -87 -2063 87
rect -2017 -87 -1988 87
rect -2076 -100 -1988 -87
rect -1888 87 -1784 100
rect -1888 -87 -1859 87
rect -1813 -87 -1784 87
rect -1888 -100 -1784 -87
rect -1684 87 -1580 100
rect -1684 -87 -1655 87
rect -1609 -87 -1580 87
rect -1684 -100 -1580 -87
rect -1480 87 -1376 100
rect -1480 -87 -1451 87
rect -1405 -87 -1376 87
rect -1480 -100 -1376 -87
rect -1276 87 -1172 100
rect -1276 -87 -1247 87
rect -1201 -87 -1172 87
rect -1276 -100 -1172 -87
rect -1072 87 -968 100
rect -1072 -87 -1043 87
rect -997 -87 -968 87
rect -1072 -100 -968 -87
rect -868 87 -764 100
rect -868 -87 -839 87
rect -793 -87 -764 87
rect -868 -100 -764 -87
rect -664 87 -560 100
rect -664 -87 -635 87
rect -589 -87 -560 87
rect -664 -100 -560 -87
rect -460 87 -356 100
rect -460 -87 -431 87
rect -385 -87 -356 87
rect -460 -100 -356 -87
rect -256 87 -152 100
rect -256 -87 -227 87
rect -181 -87 -152 87
rect -256 -100 -152 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 152 87 256 100
rect 152 -87 181 87
rect 227 -87 256 87
rect 152 -100 256 -87
rect 356 87 460 100
rect 356 -87 385 87
rect 431 -87 460 87
rect 356 -100 460 -87
rect 560 87 664 100
rect 560 -87 589 87
rect 635 -87 664 87
rect 560 -100 664 -87
rect 764 87 868 100
rect 764 -87 793 87
rect 839 -87 868 87
rect 764 -100 868 -87
rect 968 87 1072 100
rect 968 -87 997 87
rect 1043 -87 1072 87
rect 968 -100 1072 -87
rect 1172 87 1276 100
rect 1172 -87 1201 87
rect 1247 -87 1276 87
rect 1172 -100 1276 -87
rect 1376 87 1480 100
rect 1376 -87 1405 87
rect 1451 -87 1480 87
rect 1376 -100 1480 -87
rect 1580 87 1684 100
rect 1580 -87 1609 87
rect 1655 -87 1684 87
rect 1580 -100 1684 -87
rect 1784 87 1888 100
rect 1784 -87 1813 87
rect 1859 -87 1888 87
rect 1784 -100 1888 -87
rect 1988 87 2076 100
rect 1988 -87 2017 87
rect 2063 -87 2076 87
rect 1988 -100 2076 -87
<< pdiffc >>
rect -2063 -87 -2017 87
rect -1859 -87 -1813 87
rect -1655 -87 -1609 87
rect -1451 -87 -1405 87
rect -1247 -87 -1201 87
rect -1043 -87 -997 87
rect -839 -87 -793 87
rect -635 -87 -589 87
rect -431 -87 -385 87
rect -227 -87 -181 87
rect -23 -87 23 87
rect 181 -87 227 87
rect 385 -87 431 87
rect 589 -87 635 87
rect 793 -87 839 87
rect 997 -87 1043 87
rect 1201 -87 1247 87
rect 1405 -87 1451 87
rect 1609 -87 1655 87
rect 1813 -87 1859 87
rect 2017 -87 2063 87
<< polysilicon >>
rect -1988 100 -1888 144
rect -1784 100 -1684 144
rect -1580 100 -1480 144
rect -1376 100 -1276 144
rect -1172 100 -1072 144
rect -968 100 -868 144
rect -764 100 -664 144
rect -560 100 -460 144
rect -356 100 -256 144
rect -152 100 -52 144
rect 52 100 152 144
rect 256 100 356 144
rect 460 100 560 144
rect 664 100 764 144
rect 868 100 968 144
rect 1072 100 1172 144
rect 1276 100 1376 144
rect 1480 100 1580 144
rect 1684 100 1784 144
rect 1888 100 1988 144
rect -1988 -144 -1888 -100
rect -1784 -144 -1684 -100
rect -1580 -144 -1480 -100
rect -1376 -144 -1276 -100
rect -1172 -144 -1072 -100
rect -968 -144 -868 -100
rect -764 -144 -664 -100
rect -560 -144 -460 -100
rect -356 -144 -256 -100
rect -152 -144 -52 -100
rect 52 -144 152 -100
rect 256 -144 356 -100
rect 460 -144 560 -100
rect 664 -144 764 -100
rect 868 -144 968 -100
rect 1072 -144 1172 -100
rect 1276 -144 1376 -100
rect 1480 -144 1580 -100
rect 1684 -144 1784 -100
rect 1888 -144 1988 -100
<< metal1 >>
rect -2063 87 -2017 98
rect -2063 -98 -2017 -87
rect -1859 87 -1813 98
rect -1859 -98 -1813 -87
rect -1655 87 -1609 98
rect -1655 -98 -1609 -87
rect -1451 87 -1405 98
rect -1451 -98 -1405 -87
rect -1247 87 -1201 98
rect -1247 -98 -1201 -87
rect -1043 87 -997 98
rect -1043 -98 -997 -87
rect -839 87 -793 98
rect -839 -98 -793 -87
rect -635 87 -589 98
rect -635 -98 -589 -87
rect -431 87 -385 98
rect -431 -98 -385 -87
rect -227 87 -181 98
rect -227 -98 -181 -87
rect -23 87 23 98
rect -23 -98 23 -87
rect 181 87 227 98
rect 181 -98 227 -87
rect 385 87 431 98
rect 385 -98 431 -87
rect 589 87 635 98
rect 589 -98 635 -87
rect 793 87 839 98
rect 793 -98 839 -87
rect 997 87 1043 98
rect 997 -98 1043 -87
rect 1201 87 1247 98
rect 1201 -98 1247 -87
rect 1405 87 1451 98
rect 1405 -98 1451 -87
rect 1609 87 1655 98
rect 1609 -98 1655 -87
rect 1813 87 1859 98
rect 1813 -98 1859 -87
rect 2017 87 2063 98
rect 2017 -98 2063 -87
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 1 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
