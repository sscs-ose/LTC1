magic
tech gf180mcuC
magscale 1 10
timestamp 1699895628
<< nwell >>
rect -284 -986 284 986
<< nsubdiff >>
rect -260 890 260 962
rect -260 -890 -188 890
rect 188 -890 260 890
rect -260 -962 260 -890
<< polysilicon >>
rect -100 789 100 802
rect -100 743 -87 789
rect 87 743 100 789
rect -100 700 100 743
rect -100 -743 100 -700
rect -100 -789 -87 -743
rect 87 -789 100 -743
rect -100 -802 100 -789
<< polycontact >>
rect -87 743 87 789
rect -87 -789 87 -743
<< ppolyres >>
rect -100 -700 100 700
<< metal1 >>
rect -98 743 -87 789
rect 87 743 98 789
rect -98 -789 -87 -743
rect 87 -789 98 -743
<< properties >>
string FIXED_BBOX -224 -926 224 926
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 7.0 m 1 nx 1 wmin 0.80 lmin 1.00 rho 315 val 2.37k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
