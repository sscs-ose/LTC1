magic
tech gf180mcuC
magscale 1 10
timestamp 1693911244
<< nwell >>
rect -362 -1902 362 1902
<< pmos >>
rect -188 1172 -132 1772
rect -28 1172 28 1772
rect 132 1172 188 1772
rect -188 436 -132 1036
rect -28 436 28 1036
rect 132 436 188 1036
rect -188 -300 -132 300
rect -28 -300 28 300
rect 132 -300 188 300
rect -188 -1036 -132 -436
rect -28 -1036 28 -436
rect 132 -1036 188 -436
rect -188 -1772 -132 -1172
rect -28 -1772 28 -1172
rect 132 -1772 188 -1172
<< pdiff >>
rect -276 1759 -188 1772
rect -276 1185 -263 1759
rect -217 1185 -188 1759
rect -276 1172 -188 1185
rect -132 1759 -28 1772
rect -132 1185 -103 1759
rect -57 1185 -28 1759
rect -132 1172 -28 1185
rect 28 1759 132 1772
rect 28 1185 57 1759
rect 103 1185 132 1759
rect 28 1172 132 1185
rect 188 1759 276 1772
rect 188 1185 217 1759
rect 263 1185 276 1759
rect 188 1172 276 1185
rect -276 1023 -188 1036
rect -276 449 -263 1023
rect -217 449 -188 1023
rect -276 436 -188 449
rect -132 1023 -28 1036
rect -132 449 -103 1023
rect -57 449 -28 1023
rect -132 436 -28 449
rect 28 1023 132 1036
rect 28 449 57 1023
rect 103 449 132 1023
rect 28 436 132 449
rect 188 1023 276 1036
rect 188 449 217 1023
rect 263 449 276 1023
rect 188 436 276 449
rect -276 287 -188 300
rect -276 -287 -263 287
rect -217 -287 -188 287
rect -276 -300 -188 -287
rect -132 287 -28 300
rect -132 -287 -103 287
rect -57 -287 -28 287
rect -132 -300 -28 -287
rect 28 287 132 300
rect 28 -287 57 287
rect 103 -287 132 287
rect 28 -300 132 -287
rect 188 287 276 300
rect 188 -287 217 287
rect 263 -287 276 287
rect 188 -300 276 -287
rect -276 -449 -188 -436
rect -276 -1023 -263 -449
rect -217 -1023 -188 -449
rect -276 -1036 -188 -1023
rect -132 -449 -28 -436
rect -132 -1023 -103 -449
rect -57 -1023 -28 -449
rect -132 -1036 -28 -1023
rect 28 -449 132 -436
rect 28 -1023 57 -449
rect 103 -1023 132 -449
rect 28 -1036 132 -1023
rect 188 -449 276 -436
rect 188 -1023 217 -449
rect 263 -1023 276 -449
rect 188 -1036 276 -1023
rect -276 -1185 -188 -1172
rect -276 -1759 -263 -1185
rect -217 -1759 -188 -1185
rect -276 -1772 -188 -1759
rect -132 -1185 -28 -1172
rect -132 -1759 -103 -1185
rect -57 -1759 -28 -1185
rect -132 -1772 -28 -1759
rect 28 -1185 132 -1172
rect 28 -1759 57 -1185
rect 103 -1759 132 -1185
rect 28 -1772 132 -1759
rect 188 -1185 276 -1172
rect 188 -1759 217 -1185
rect 263 -1759 276 -1185
rect 188 -1772 276 -1759
<< pdiffc >>
rect -263 1185 -217 1759
rect -103 1185 -57 1759
rect 57 1185 103 1759
rect 217 1185 263 1759
rect -263 449 -217 1023
rect -103 449 -57 1023
rect 57 449 103 1023
rect 217 449 263 1023
rect -263 -287 -217 287
rect -103 -287 -57 287
rect 57 -287 103 287
rect 217 -287 263 287
rect -263 -1023 -217 -449
rect -103 -1023 -57 -449
rect 57 -1023 103 -449
rect 217 -1023 263 -449
rect -263 -1759 -217 -1185
rect -103 -1759 -57 -1185
rect 57 -1759 103 -1185
rect 217 -1759 263 -1185
<< polysilicon >>
rect -188 1772 -132 1816
rect -28 1772 28 1816
rect 132 1772 188 1816
rect -188 1128 -132 1172
rect -28 1128 28 1172
rect 132 1128 188 1172
rect -188 1036 -132 1080
rect -28 1036 28 1080
rect 132 1036 188 1080
rect -188 392 -132 436
rect -28 392 28 436
rect 132 392 188 436
rect -188 300 -132 344
rect -28 300 28 344
rect 132 300 188 344
rect -188 -344 -132 -300
rect -28 -344 28 -300
rect 132 -344 188 -300
rect -188 -436 -132 -392
rect -28 -436 28 -392
rect 132 -436 188 -392
rect -188 -1080 -132 -1036
rect -28 -1080 28 -1036
rect 132 -1080 188 -1036
rect -188 -1172 -132 -1128
rect -28 -1172 28 -1128
rect 132 -1172 188 -1128
rect -188 -1816 -132 -1772
rect -28 -1816 28 -1772
rect 132 -1816 188 -1772
<< metal1 >>
rect -263 1759 -217 1770
rect -263 1174 -217 1185
rect -103 1759 -57 1770
rect -103 1174 -57 1185
rect 57 1759 103 1770
rect 57 1174 103 1185
rect 217 1759 263 1770
rect 217 1174 263 1185
rect -263 1023 -217 1034
rect -263 438 -217 449
rect -103 1023 -57 1034
rect -103 438 -57 449
rect 57 1023 103 1034
rect 57 438 103 449
rect 217 1023 263 1034
rect 217 438 263 449
rect -263 287 -217 298
rect -263 -298 -217 -287
rect -103 287 -57 298
rect -103 -298 -57 -287
rect 57 287 103 298
rect 57 -298 103 -287
rect 217 287 263 298
rect 217 -298 263 -287
rect -263 -449 -217 -438
rect -263 -1034 -217 -1023
rect -103 -449 -57 -438
rect -103 -1034 -57 -1023
rect 57 -449 103 -438
rect 57 -1034 103 -1023
rect 217 -449 263 -438
rect 217 -1034 263 -1023
rect -263 -1185 -217 -1174
rect -263 -1770 -217 -1759
rect -103 -1185 -57 -1174
rect -103 -1770 -57 -1759
rect 57 -1185 103 -1174
rect 57 -1770 103 -1759
rect 217 -1185 263 -1174
rect 217 -1770 263 -1759
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 5 nf 3 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
