magic
tech gf180mcuD
magscale 1 10
timestamp 1713971633
<< checkpaint >>
rect -2265 -4148 24479 4078
<< nwell >>
rect 3381 1155 3507 1735
rect 6847 1155 7123 1735
rect 12283 916 13002 1935
rect 3360 -1918 3502 -1338
rect 6860 -1918 6998 -1338
rect 10342 -1918 10688 -1338
rect 13997 -1918 14178 -1372
rect 15694 -1918 15819 -1372
rect 17325 -1918 17473 -1372
<< pwell >>
rect 13720 -1303 14217 -995
rect 15630 -1329 15857 -1038
<< metal1 >>
rect 12842 2016 14766 2062
rect 10286 1826 11156 1970
rect 12023 1896 12075 1897
rect 12023 1843 12075 1844
rect 12201 1893 12253 1894
rect 12201 1840 12253 1841
rect -265 1619 280 1734
rect -265 -1797 -150 1619
rect 2818 1614 7180 1729
rect 10286 1614 10402 1826
rect 12842 1434 12888 2016
rect 14154 1897 14206 1898
rect 13188 1895 13240 1896
rect 13065 1891 13117 1892
rect 14154 1844 14206 1845
rect 14273 1895 14325 1896
rect 13188 1842 13240 1843
rect 14273 1842 14325 1843
rect 13065 1838 13117 1839
rect 12842 1393 12943 1434
rect 3098 224 3160 226
rect 2945 219 3007 221
rect 2945 167 2950 219
rect 3002 167 3007 219
rect 3098 172 3103 224
rect 3155 172 3160 224
rect 3098 171 3160 172
rect 3252 224 3314 226
rect 3252 172 3257 224
rect 3309 172 3314 224
rect 3252 171 3314 172
rect 2945 166 3007 167
rect 2840 -355 2902 -353
rect 2840 -407 2845 -355
rect 2897 -407 2902 -355
rect 2840 -408 2902 -407
rect 3085 -355 3147 -353
rect 3085 -407 3090 -355
rect 3142 -407 3147 -355
rect 3085 -408 3147 -407
rect 3234 -357 3296 -355
rect 3234 -409 3239 -357
rect 3291 -409 3296 -357
rect 3234 -410 3296 -409
rect 6414 -364 6476 -362
rect 6414 -416 6419 -364
rect 6471 -416 6476 -364
rect 6578 -364 6703 302
rect 10305 -42 10426 254
rect 10731 126 10793 128
rect 10731 74 10736 126
rect 10788 74 10793 126
rect 10731 73 10793 74
rect 12505 122 12555 1361
rect 12842 1347 12950 1393
rect 14567 985 14617 1361
rect 14550 973 14627 985
rect 14550 921 14562 973
rect 14614 921 14627 973
rect 14550 909 14627 921
rect 14541 381 14617 395
rect 14541 374 14553 381
rect 14528 329 14553 374
rect 14605 329 14617 381
rect 14528 317 14617 329
rect 12505 72 12860 122
rect 10305 -49 11057 -42
rect 10259 -163 11057 -49
rect 12318 -101 12903 -42
rect 6578 -412 6593 -364
rect 6414 -417 6476 -416
rect 6588 -416 6593 -412
rect 6645 -412 6703 -364
rect 6746 -363 6808 -361
rect 6645 -416 6650 -412
rect 6746 -415 6751 -363
rect 6803 -415 6808 -363
rect 6746 -416 6808 -415
rect 6588 -417 6650 -416
rect 10259 -446 10384 -163
rect 13698 -461 13823 -43
rect 14528 -216 14574 317
rect 14199 -262 14574 -216
rect 14199 -657 14245 -262
rect 14720 -517 14766 2016
rect 22331 1401 22479 1447
rect 17008 983 17102 1002
rect 17008 931 17029 983
rect 17081 931 17102 983
rect 17008 918 17102 931
rect 15041 868 15126 872
rect 14928 787 15126 868
rect 15041 -317 15126 787
rect 15041 -402 15990 -317
rect 14720 -563 15859 -517
rect 14199 -703 15695 -657
rect 2072 -858 2151 -850
rect 13909 -858 14320 -774
rect 15310 -787 15368 -786
rect 15310 -839 15313 -787
rect 15365 -839 15368 -787
rect 15310 -840 15368 -839
rect 15444 -790 15502 -789
rect 15444 -842 15447 -790
rect 15499 -842 15502 -790
rect 15444 -843 15502 -842
rect 2072 -910 2085 -858
rect 2137 -910 2151 -858
rect 2072 -924 2151 -910
rect 15649 -922 15695 -703
rect 15813 -665 15859 -563
rect 15905 -524 15990 -402
rect 15905 -537 17133 -524
rect 15905 -589 16931 -537
rect 16983 -589 17064 -537
rect 17116 -589 17133 -537
rect 15905 -609 17133 -589
rect 15813 -711 17370 -665
rect 16939 -781 16997 -780
rect 16033 -784 16091 -783
rect 15893 -789 15951 -788
rect 15893 -841 15896 -789
rect 15948 -841 15951 -789
rect 16033 -836 16036 -784
rect 16088 -836 16091 -784
rect 16939 -833 16942 -781
rect 16994 -833 16997 -781
rect 16939 -834 16997 -833
rect 17108 -783 17166 -782
rect 17108 -835 17111 -783
rect 17163 -835 17166 -783
rect 17108 -836 17166 -835
rect 16033 -837 16091 -836
rect 15893 -842 15951 -841
rect 14255 -957 14337 -940
rect 14255 -1009 14270 -957
rect 14322 -1009 14337 -957
rect 14255 -1018 14337 -1009
rect 15550 -968 15695 -922
rect 14150 -1375 14221 -1362
rect 15550 -1370 15596 -968
rect 15759 -969 15843 -956
rect 15759 -1021 15776 -969
rect 15828 -1018 16168 -969
rect 15828 -1021 15843 -1018
rect 15759 -1035 15843 -1021
rect 15764 -1370 15823 -1358
rect 14150 -1427 14165 -1375
rect 14217 -1427 14221 -1375
rect 14150 -1440 14221 -1427
rect 15764 -1371 15834 -1370
rect 15764 -1423 15779 -1371
rect 15831 -1423 15834 -1371
rect 17324 -1391 17370 -711
rect 17711 -778 17769 -777
rect 17589 -780 17647 -779
rect 17589 -832 17592 -780
rect 17644 -832 17647 -780
rect 17711 -830 17714 -778
rect 17766 -830 17769 -778
rect 17711 -831 17769 -830
rect 17589 -833 17647 -832
rect 15764 -1424 15834 -1423
rect 15764 -1436 15823 -1424
rect 17204 -1437 17370 -1391
rect 18279 -1422 18647 -1376
rect -265 -1912 187 -1797
rect 3123 -1912 3729 -1797
rect 6581 -1912 7192 -1797
rect 10064 -1892 16443 -1813
rect 17142 -1892 17665 -1813
rect 2071 -1963 2148 -1958
rect 2071 -2015 2083 -1963
rect 2135 -2015 2148 -1963
rect 2071 -2027 2148 -2015
rect 1031 -2076 1107 -2061
rect 2085 -2076 2131 -2027
rect 18601 -2076 18647 -1422
rect 1031 -2122 18647 -2076
rect 1031 -2137 1107 -2122
<< via1 >>
rect 12023 1844 12075 1896
rect 12201 1841 12253 1893
rect 13065 1839 13117 1891
rect 13188 1843 13240 1895
rect 14154 1845 14206 1897
rect 14273 1843 14325 1895
rect 2950 167 3002 219
rect 3103 172 3155 224
rect 3257 172 3309 224
rect 2845 -407 2897 -355
rect 3090 -407 3142 -355
rect 3239 -409 3291 -357
rect 6419 -416 6471 -364
rect 10736 74 10788 126
rect 14562 921 14614 973
rect 14553 329 14605 381
rect 6593 -416 6645 -364
rect 6751 -415 6803 -363
rect 17029 931 17081 983
rect 15313 -839 15365 -787
rect 15447 -842 15499 -790
rect 2085 -910 2137 -858
rect 16931 -589 16983 -537
rect 17064 -589 17116 -537
rect 15896 -841 15948 -789
rect 16036 -836 16088 -784
rect 16942 -833 16994 -781
rect 17111 -835 17163 -783
rect 14270 -1009 14322 -957
rect 15776 -1021 15828 -969
rect 14165 -1427 14217 -1375
rect 15779 -1423 15831 -1371
rect 17592 -832 17644 -780
rect 17714 -830 17766 -778
rect 2083 -2015 2135 -1963
<< metal2 >>
rect 12000 1896 13265 1903
rect 12000 1844 12023 1896
rect 12075 1895 13265 1896
rect 12075 1893 13188 1895
rect 12075 1844 12201 1893
rect 12000 1841 12201 1844
rect 12253 1891 13188 1893
rect 12253 1841 13065 1891
rect 12000 1839 13065 1841
rect 13117 1843 13188 1891
rect 13240 1843 13265 1895
rect 13117 1839 13265 1843
rect 14128 1897 15175 1902
rect 14128 1845 14154 1897
rect 14206 1895 15175 1897
rect 14206 1845 14273 1895
rect 14128 1843 14273 1845
rect 14325 1843 15175 1895
rect 14128 1839 15175 1843
rect 12000 1833 13265 1839
rect 1059 1747 10879 1803
rect 1059 1034 1115 1747
rect 8181 1523 10579 1579
rect 8181 1335 8237 1523
rect 6979 1279 8237 1335
rect 4672 446 5480 502
rect 2918 224 4016 239
rect 2918 219 3103 224
rect 2918 167 2950 219
rect 3002 172 3103 219
rect 3155 172 3257 224
rect 3309 172 4016 224
rect 3002 167 4016 172
rect 2918 161 4016 167
rect 5424 -56 5480 446
rect 6979 -56 7035 1279
rect 10523 946 10579 1523
rect 10823 1348 10879 1747
rect 17008 985 17102 1002
rect 14550 975 14627 985
rect 10523 890 10923 946
rect 12828 897 12967 958
rect 14550 919 14561 975
rect 14617 919 14627 975
rect 14550 909 14627 919
rect 17008 929 17027 985
rect 17083 929 17102 985
rect 17008 918 17102 929
rect 12828 890 12948 897
rect 8259 446 9057 502
rect 5424 -112 7035 -56
rect 9001 -56 9057 446
rect 12828 385 12889 890
rect 14541 385 14617 395
rect 12828 381 14617 385
rect 12828 329 14553 381
rect 14605 329 14617 381
rect 12828 324 14617 329
rect 14541 317 14617 324
rect 10691 126 10880 134
rect 10691 74 10736 126
rect 10788 78 10880 126
rect 10788 74 10805 78
rect 10691 65 10805 74
rect 10691 -56 10747 65
rect 9001 -112 10747 -56
rect 12439 -113 14180 -57
rect 12439 -196 12495 -113
rect 10450 -252 12495 -196
rect 2793 -355 4014 -344
rect 2793 -407 2845 -355
rect 2897 -407 3090 -355
rect 3142 -357 4014 -355
rect 3142 -407 3239 -357
rect 2793 -409 3239 -407
rect 3291 -409 4014 -357
rect 2793 -422 4014 -409
rect 6384 -363 7657 -344
rect 6384 -364 6751 -363
rect 6384 -416 6419 -364
rect 6471 -416 6593 -364
rect 6645 -415 6751 -364
rect 6803 -415 7657 -363
rect 6645 -416 7657 -415
rect 6384 -422 7657 -416
rect 2072 -857 2150 -844
rect 2072 -913 2082 -857
rect 2138 -913 2150 -857
rect 2072 -924 2150 -913
rect 1041 -2061 1097 -1118
rect 2071 -1961 2148 -1951
rect 2071 -2017 2081 -1961
rect 2137 -2017 2148 -1961
rect 2071 -2027 2148 -2017
rect 4536 -2042 4592 -1196
rect 8023 -1915 8079 -1124
rect 10450 -1915 10506 -252
rect 14124 -959 14180 -113
rect 16912 -526 17134 -524
rect 16910 -537 17134 -526
rect 16910 -589 16931 -537
rect 16983 -589 17064 -537
rect 17116 -589 17134 -537
rect 16910 -609 17134 -589
rect 16910 -771 16992 -609
rect 16910 -773 17815 -771
rect 14925 -784 16167 -775
rect 14925 -787 16036 -784
rect 14925 -839 15313 -787
rect 15365 -789 16036 -787
rect 15365 -790 15896 -789
rect 15365 -839 15447 -790
rect 14925 -842 15447 -839
rect 15499 -841 15896 -790
rect 15948 -836 16036 -789
rect 16088 -836 16167 -784
rect 15948 -841 16167 -836
rect 15499 -842 16167 -841
rect 14925 -856 16167 -842
rect 16911 -778 17815 -773
rect 16911 -780 17714 -778
rect 16911 -781 17592 -780
rect 16911 -833 16942 -781
rect 16994 -783 17592 -781
rect 16994 -833 17111 -783
rect 16911 -835 17111 -833
rect 17163 -832 17592 -783
rect 17644 -830 17714 -780
rect 17766 -830 17815 -778
rect 17644 -832 17815 -830
rect 17163 -835 17815 -832
rect 16911 -846 17815 -835
rect 14255 -957 14342 -940
rect 14255 -959 14270 -957
rect 14124 -1009 14270 -959
rect 14322 -1009 14342 -957
rect 14124 -1015 14342 -1009
rect 14255 -1022 14342 -1015
rect 15759 -969 15843 -956
rect 15759 -1025 15772 -969
rect 15828 -1025 15843 -969
rect 15759 -1035 15843 -1025
rect 11674 -1734 11730 -1146
rect 14150 -1367 14221 -1362
rect 14150 -1372 14268 -1367
rect 15711 -1371 15855 -1364
rect 14079 -1375 14270 -1372
rect 14079 -1427 14165 -1375
rect 14217 -1427 14270 -1375
rect 14079 -1428 14270 -1427
rect 15711 -1423 15779 -1371
rect 15831 -1423 15855 -1371
rect 14079 -1432 14268 -1428
rect 15711 -1432 15855 -1423
rect 14079 -1440 14221 -1432
rect 14079 -1734 14135 -1440
rect 11674 -1790 14135 -1734
rect 8023 -1971 10506 -1915
rect 15711 -2042 15767 -1432
rect 1031 -2071 1107 -2061
rect 1031 -2127 1041 -2071
rect 1097 -2127 1107 -2071
rect 4536 -2098 15767 -2042
rect 1031 -2137 1107 -2127
<< via2 >>
rect 14561 973 14617 975
rect 14561 921 14562 973
rect 14562 921 14614 973
rect 14614 921 14617 973
rect 14561 919 14617 921
rect 17027 983 17083 985
rect 17027 931 17029 983
rect 17029 931 17081 983
rect 17081 931 17083 983
rect 17027 929 17083 931
rect 2082 -858 2138 -857
rect 2082 -910 2085 -858
rect 2085 -910 2137 -858
rect 2137 -910 2138 -858
rect 2082 -913 2138 -910
rect 2081 -1963 2137 -1961
rect 2081 -2015 2083 -1963
rect 2083 -2015 2135 -1963
rect 2135 -2015 2137 -1963
rect 2081 -2017 2137 -2015
rect 15772 -1021 15776 -969
rect 15776 -1021 15828 -969
rect 15772 -1025 15828 -1021
rect 1041 -2127 1097 -2071
<< metal3 >>
rect 14549 984 14629 986
rect 17008 985 17102 1002
rect 17008 984 17027 985
rect 14549 975 17027 984
rect 14549 919 14561 975
rect 14617 929 17027 975
rect 17083 984 17102 985
rect 17083 929 17117 984
rect 14617 921 17117 929
rect 14617 919 14629 921
rect 14549 909 14629 919
rect 17008 918 17102 921
rect 2072 -857 2150 -844
rect 2072 -913 2082 -857
rect 2138 -913 2150 -857
rect 2072 -924 2150 -913
rect 2078 -1949 2140 -924
rect 15759 -964 15843 -956
rect 15759 -969 16118 -964
rect 15759 -1025 15772 -969
rect 15828 -1022 16118 -969
rect 15828 -1025 15855 -1022
rect 15759 -1035 15855 -1025
rect 2070 -1961 2148 -1949
rect 2070 -2017 2081 -1961
rect 2137 -2017 2148 -1961
rect 2070 -2028 2148 -2017
rect 1031 -2071 1107 -2061
rect 1031 -2127 1041 -2071
rect 1097 -2090 1107 -2071
rect 15797 -2090 15855 -1035
rect 1097 -2127 15855 -2090
rect 1031 -2137 15855 -2127
rect 1037 -2148 15855 -2137
use 3_inp_AND_magic  3_inp_AND_magic_0
timestamp 1713349043
transform 1 0 12952 0 1 1400
box -184 -1564 1665 536
use 3_inp_AND_magic  3_inp_AND_magic_1
timestamp 1713349043
transform 1 0 10891 0 1 1400
box -184 -1564 1665 536
use AND2_magic  AND2_magic_0
timestamp 1713185578
transform 1 0 15750 0 -1 -1372
box 35 -598 1575 546
use AND2_magic  AND2_magic_1
timestamp 1713185578
transform 1 0 14120 0 -1 -1372
box 35 -598 1575 546
use inverter_magic  inverter_magic_0
timestamp 1713185578
transform 1 0 17458 0 -1 -1338
box 0 -569 1108 580
use neg_DFF_magic  neg_DFF_magic_0
timestamp 1713971633
transform 1 0 16895 0 1 316
box -2075 -823 5510 1762
use xnor_magic  xnor_magic_0
timestamp 1713971188
transform 1 0 8242 0 1 1186
box -1158 -1186 2262 549
use xnor_magic  xnor_magic_1
timestamp 1713971188
transform 1 0 1140 0 -1 -1369
box -1158 -1186 2262 549
use xnor_magic  xnor_magic_2
timestamp 1713971188
transform 1 0 11773 0 -1 -1369
box -1158 -1186 2262 549
use xnor_magic  xnor_magic_3
timestamp 1713971188
transform 1 0 1158 0 1 1186
box -1158 -1186 2262 549
use xnor_magic  xnor_magic_4
timestamp 1713971188
transform 1 0 4653 0 1 1186
box -1158 -1186 2262 549
use xnor_magic  xnor_magic_5
timestamp 1713971188
transform 1 0 4635 0 -1 -1369
box -1158 -1186 2262 549
use xnor_magic  xnor_magic_6
timestamp 1713971188
transform 1 0 8122 0 -1 -1369
box -1158 -1186 2262 549
<< labels >>
flabel metal1 s 10576 1891 10576 1891 0 FreeSans 750 0 0 0 VDD
port 1 nsew
flabel metal1 s 22451 1421 22451 1421 0 FreeSans 750 0 0 0 P3
port 2 nsew
flabel metal1 s 10326 -267 10326 -267 0 FreeSans 750 0 0 0 VSS
port 3 nsew
<< end >>
