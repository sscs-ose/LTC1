magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2128 -2457 2128 2457
<< nwell >>
rect -128 -457 128 457
<< nsubdiff >>
rect -45 352 45 374
rect -45 -352 -23 352
rect 23 -352 45 352
rect -45 -374 45 -352
<< nsubdiffcont >>
rect -23 -352 23 352
<< metal1 >>
rect -34 352 34 363
rect -34 -352 -23 352
rect 23 -352 34 352
rect -34 -363 34 -352
<< end >>
