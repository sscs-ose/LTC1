magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1357 -1019 1357 1019
<< metal1 >>
rect -357 13 357 19
rect -357 -13 -351 13
rect 351 -13 357 13
rect -357 -19 357 -13
<< via1 >>
rect -351 -13 351 13
<< metal2 >>
rect -357 13 357 19
rect -357 -13 -351 13
rect 351 -13 357 13
rect -357 -19 357 -13
<< end >>
