magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2000 -2569 3108 2580
<< nwell >>
rect 0 484 1108 580
rect 400 470 680 484
rect 407 461 680 470
<< psubdiff >>
rect 401 -507 715 -488
rect 401 -553 527 -507
rect 573 -553 715 -507
rect 401 -569 715 -553
<< nsubdiff >>
rect 407 520 680 535
rect 407 474 514 520
rect 560 474 680 520
rect 407 461 680 474
<< psubdiffcont >>
rect 527 -553 573 -507
<< nsubdiffcont >>
rect 514 474 560 520
<< polysilicon >>
rect 174 387 934 425
rect 390 5 501 89
rect 329 -9 501 5
rect 329 -55 349 -9
rect 395 -55 501 -9
rect 329 -59 501 -55
rect 329 -69 411 -59
rect 390 -391 718 -354
<< polycontact >>
rect 349 -55 395 -9
<< metal1 >>
rect 78 520 1043 536
rect 78 474 514 520
rect 560 474 1043 520
rect 78 459 1043 474
rect 99 143 145 459
rect 315 86 361 144
rect 531 143 577 459
rect 963 143 1009 459
rect 747 86 793 143
rect 315 84 793 86
rect 315 38 900 84
rect 329 -9 410 -8
rect 261 -55 349 -9
rect 395 -55 410 -9
rect 329 -59 410 -55
rect 315 -488 361 -105
rect 531 -116 577 38
rect 747 -488 793 -105
rect 100 -507 1065 -488
rect 100 -553 527 -507
rect 573 -553 1065 -507
rect 100 -569 1065 -553
use nmos_3p3_F2UGVV  nmos_3p3_F2UGVV_0
timestamp 1713185578
transform 1 0 554 0 1 -215
box -276 -180 276 180
use pmos_3p3_VH67F7  pmos_3p3_VH67F7_0
timestamp 1713185578
transform 1 0 554 0 1 242
box -554 -242 554 242
<< labels >>
flabel nsubdiffcont 536 497 536 497 0 FreeSans 750 0 0 0 VDD
flabel psubdiffcont 551 -530 551 -530 0 FreeSans 750 0 0 0 VSS
flabel metal1 s 273 -31 273 -31 0 FreeSans 750 0 0 0 VIN
port 1 nsew
flabel metal1 s 862 59 862 59 0 FreeSans 750 0 0 0 VOUT
port 2 nsew
<< end >>
