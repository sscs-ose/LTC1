magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7486 -2128 7486 2128
<< nwell >>
rect -5486 -128 5486 128
<< nsubdiff >>
rect -5403 23 5403 45
rect -5403 -23 -5381 23
rect 5381 -23 5403 23
rect -5403 -45 5403 -23
<< nsubdiffcont >>
rect -5381 -23 5381 23
<< metal1 >>
rect -5392 23 5392 34
rect -5392 -23 -5381 23
rect 5381 -23 5392 23
rect -5392 -34 5392 -23
<< end >>
