magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2285 -2452 5979 4227
<< nwell >>
rect 1154 811 1332 1134
rect 2392 813 2558 1134
<< psubdiff >>
rect -280 1967 3975 1994
rect -280 1921 -146 1967
rect -100 1921 4 1967
rect 50 1921 154 1967
rect 200 1921 304 1967
rect 350 1921 454 1967
rect 500 1921 604 1967
rect 650 1921 754 1967
rect 800 1921 904 1967
rect 950 1921 1054 1967
rect 1100 1921 1204 1967
rect 1250 1921 1354 1967
rect 1400 1921 1504 1967
rect 1550 1921 1654 1967
rect 1700 1921 1804 1967
rect 1850 1921 1954 1967
rect 2000 1921 2104 1967
rect 2150 1921 2254 1967
rect 2300 1921 2404 1967
rect 2450 1921 2554 1967
rect 2600 1921 2704 1967
rect 2750 1921 2854 1967
rect 2900 1921 3004 1967
rect 3050 1921 3154 1967
rect 3200 1921 3304 1967
rect 3350 1921 3454 1967
rect 3500 1921 3604 1967
rect 3650 1921 3754 1967
rect 3800 1921 3975 1967
rect -280 1884 3975 1921
rect -280 1834 -170 1884
rect -280 1788 -248 1834
rect -202 1788 -170 1834
rect -280 1684 -170 1788
rect -280 1638 -248 1684
rect -202 1638 -170 1684
rect -280 1534 -170 1638
rect -280 1488 -248 1534
rect -202 1488 -170 1534
rect -280 1384 -170 1488
rect -280 1338 -248 1384
rect -202 1338 -170 1384
rect -280 1234 -170 1338
rect -280 1188 -248 1234
rect -202 1188 -170 1234
rect -280 1084 -170 1188
rect -280 1038 -248 1084
rect -202 1038 -170 1084
rect -280 934 -170 1038
rect -280 888 -248 934
rect -202 888 -170 934
rect -280 784 -170 888
rect -280 738 -248 784
rect -202 738 -170 784
rect -280 634 -170 738
rect -280 588 -248 634
rect -202 588 -170 634
rect -280 484 -170 588
rect -280 438 -248 484
rect -202 438 -170 484
rect -280 334 -170 438
rect -280 288 -248 334
rect -202 288 -170 334
rect -280 184 -170 288
rect -280 138 -248 184
rect -202 138 -170 184
rect -280 34 -170 138
rect -280 -12 -248 34
rect -202 -12 -170 34
rect -280 -79 -170 -12
rect 3865 1794 3975 1884
rect 3865 1748 3894 1794
rect 3940 1748 3975 1794
rect 3865 1644 3975 1748
rect 3865 1598 3894 1644
rect 3940 1598 3975 1644
rect 3865 1494 3975 1598
rect 3865 1448 3894 1494
rect 3940 1448 3975 1494
rect 3865 1344 3975 1448
rect 3865 1298 3894 1344
rect 3940 1298 3975 1344
rect 3865 1194 3975 1298
rect 3865 1148 3894 1194
rect 3940 1148 3975 1194
rect 3865 1044 3975 1148
rect 3865 998 3894 1044
rect 3940 998 3975 1044
rect 3865 894 3975 998
rect 3865 848 3894 894
rect 3940 848 3975 894
rect 3865 744 3975 848
rect 3865 698 3894 744
rect 3940 698 3975 744
rect 3865 594 3975 698
rect 3865 548 3894 594
rect 3940 548 3975 594
rect 3865 444 3975 548
rect 3865 398 3894 444
rect 3940 398 3975 444
rect 3865 294 3975 398
rect 3865 248 3894 294
rect 3940 248 3975 294
rect 3865 144 3975 248
rect 3865 98 3894 144
rect 3940 98 3975 144
rect 3865 -6 3975 98
rect 3865 -52 3894 -6
rect 3940 -52 3975 -6
rect 3865 -79 3975 -52
rect -280 -112 3975 -79
rect -280 -158 -129 -112
rect -83 -158 21 -112
rect 67 -158 171 -112
rect 217 -158 321 -112
rect 367 -158 471 -112
rect 517 -158 621 -112
rect 667 -158 771 -112
rect 817 -158 921 -112
rect 967 -158 1071 -112
rect 1117 -158 1221 -112
rect 1267 -158 1371 -112
rect 1417 -158 1521 -112
rect 1567 -158 1671 -112
rect 1717 -158 1821 -112
rect 1867 -158 1971 -112
rect 2017 -158 2121 -112
rect 2167 -158 2271 -112
rect 2317 -158 2421 -112
rect 2467 -158 2571 -112
rect 2617 -158 2721 -112
rect 2767 -158 2871 -112
rect 2917 -158 3021 -112
rect 3067 -158 3171 -112
rect 3217 -158 3321 -112
rect 3367 -158 3471 -112
rect 3517 -158 3621 -112
rect 3667 -158 3771 -112
rect 3817 -158 3975 -112
rect -280 -189 3975 -158
<< psubdiffcont >>
rect -146 1921 -100 1967
rect 4 1921 50 1967
rect 154 1921 200 1967
rect 304 1921 350 1967
rect 454 1921 500 1967
rect 604 1921 650 1967
rect 754 1921 800 1967
rect 904 1921 950 1967
rect 1054 1921 1100 1967
rect 1204 1921 1250 1967
rect 1354 1921 1400 1967
rect 1504 1921 1550 1967
rect 1654 1921 1700 1967
rect 1804 1921 1850 1967
rect 1954 1921 2000 1967
rect 2104 1921 2150 1967
rect 2254 1921 2300 1967
rect 2404 1921 2450 1967
rect 2554 1921 2600 1967
rect 2704 1921 2750 1967
rect 2854 1921 2900 1967
rect 3004 1921 3050 1967
rect 3154 1921 3200 1967
rect 3304 1921 3350 1967
rect 3454 1921 3500 1967
rect 3604 1921 3650 1967
rect 3754 1921 3800 1967
rect -248 1788 -202 1834
rect -248 1638 -202 1684
rect -248 1488 -202 1534
rect -248 1338 -202 1384
rect -248 1188 -202 1234
rect -248 1038 -202 1084
rect -248 888 -202 934
rect -248 738 -202 784
rect -248 588 -202 634
rect -248 438 -202 484
rect -248 288 -202 334
rect -248 138 -202 184
rect -248 -12 -202 34
rect 3894 1748 3940 1794
rect 3894 1598 3940 1644
rect 3894 1448 3940 1494
rect 3894 1298 3940 1344
rect 3894 1148 3940 1194
rect 3894 998 3940 1044
rect 3894 848 3940 894
rect 3894 698 3940 744
rect 3894 548 3940 594
rect 3894 398 3940 444
rect 3894 248 3940 294
rect 3894 98 3940 144
rect 3894 -52 3940 -6
rect -129 -158 -83 -112
rect 21 -158 67 -112
rect 171 -158 217 -112
rect 321 -158 367 -112
rect 471 -158 517 -112
rect 621 -158 667 -112
rect 771 -158 817 -112
rect 921 -158 967 -112
rect 1071 -158 1117 -112
rect 1221 -158 1267 -112
rect 1371 -158 1417 -112
rect 1521 -158 1567 -112
rect 1671 -158 1717 -112
rect 1821 -158 1867 -112
rect 1971 -158 2017 -112
rect 2121 -158 2167 -112
rect 2271 -158 2317 -112
rect 2421 -158 2467 -112
rect 2571 -158 2617 -112
rect 2721 -158 2767 -112
rect 2871 -158 2917 -112
rect 3021 -158 3067 -112
rect 3171 -158 3217 -112
rect 3321 -158 3367 -112
rect 3471 -158 3517 -112
rect 3621 -158 3667 -112
rect 3771 -158 3817 -112
<< metal1 >>
rect 1789 2209 1905 2227
rect 1686 2186 1905 2209
rect 1686 2134 1821 2186
rect 1873 2134 1905 2186
rect 1686 2112 1905 2134
rect 1789 2098 1905 2112
rect -285 1967 3979 1999
rect -285 1921 -146 1967
rect -100 1921 4 1967
rect 50 1921 154 1967
rect 200 1921 304 1967
rect 350 1921 454 1967
rect 500 1921 604 1967
rect 650 1921 754 1967
rect 800 1921 904 1967
rect 950 1921 1054 1967
rect 1100 1921 1204 1967
rect 1250 1921 1354 1967
rect 1400 1921 1504 1967
rect 1550 1921 1654 1967
rect 1700 1921 1804 1967
rect 1850 1921 1954 1967
rect 2000 1921 2104 1967
rect 2150 1921 2254 1967
rect 2300 1921 2404 1967
rect 2450 1921 2554 1967
rect 2600 1921 2704 1967
rect 2750 1921 2854 1967
rect 2900 1921 3004 1967
rect 3050 1921 3154 1967
rect 3200 1921 3304 1967
rect 3350 1921 3454 1967
rect 3500 1921 3604 1967
rect 3650 1921 3754 1967
rect 3800 1921 3979 1967
rect -285 1879 3979 1921
rect -285 1834 -165 1879
rect -285 1788 -248 1834
rect -202 1788 -165 1834
rect -285 1684 -165 1788
rect 3859 1794 3979 1879
rect 1076 1708 2587 1786
rect 3859 1748 3894 1794
rect 3940 1748 3979 1794
rect -285 1638 -248 1684
rect -202 1638 -165 1684
rect -285 1534 -165 1638
rect -285 1488 -248 1534
rect -202 1488 -165 1534
rect -285 1384 -165 1488
rect -285 1338 -248 1384
rect -202 1338 -165 1384
rect -285 1234 -165 1338
rect -285 1188 -248 1234
rect -202 1188 -165 1234
rect -285 1084 -165 1188
rect -285 1038 -248 1084
rect -202 1038 -165 1084
rect -285 934 -165 1038
rect -82 1196 28 1217
rect -82 1144 -60 1196
rect -8 1144 28 1196
rect -82 1084 28 1144
rect 1374 1112 1452 1708
rect 1613 1106 1691 1708
rect 1852 1099 1930 1708
rect 2078 1108 2156 1708
rect 3859 1644 3979 1748
rect 3859 1598 3894 1644
rect 3940 1598 3979 1644
rect 3859 1494 3979 1598
rect 3859 1448 3894 1494
rect 3940 1448 3979 1494
rect 3691 1338 3810 1399
rect 3691 1286 3726 1338
rect 3778 1286 3810 1338
rect 3691 1190 3810 1286
rect 3692 1153 3810 1190
rect 3692 1101 3724 1153
rect 3776 1101 3810 1153
rect -82 1044 67 1084
rect 3692 1080 3810 1101
rect 3648 1076 3810 1080
rect 3859 1344 3979 1448
rect 3859 1298 3894 1344
rect 3940 1298 3979 1344
rect 3859 1194 3979 1298
rect 3859 1148 3894 1194
rect 3940 1148 3979 1194
rect -82 1039 120 1044
rect -82 987 -67 1039
rect -15 987 120 1039
rect -82 982 120 987
rect 3648 983 3799 1076
rect 3859 1044 3979 1148
rect 3859 998 3894 1044
rect 3940 998 3979 1044
rect -82 971 67 982
rect -285 888 -248 934
rect -202 888 -165 934
rect -285 784 -165 888
rect -285 738 -248 784
rect -202 738 -165 784
rect -285 634 -165 738
rect -285 588 -248 634
rect -202 588 -165 634
rect 3859 894 3979 998
rect 3859 848 3894 894
rect 3940 848 3979 894
rect 3859 744 3979 848
rect 3859 698 3894 744
rect 3940 698 3979 744
rect -285 484 -165 588
rect -285 438 -248 484
rect -202 438 -165 484
rect -285 334 -165 438
rect -285 288 -248 334
rect -202 288 -165 334
rect -3 529 98 543
rect 235 529 307 609
rect 3859 594 3979 698
rect 3859 548 3894 594
rect 3940 548 3979 594
rect -3 519 307 529
rect 3735 524 3795 533
rect -3 467 21 519
rect 73 467 307 519
rect 3458 521 3804 524
rect -3 457 307 467
rect -3 363 98 457
rect -3 311 21 363
rect 73 311 98 363
rect 235 358 307 457
rect 1134 459 1232 512
rect 2385 488 2551 503
rect 1134 416 1453 459
rect 2336 442 2551 488
rect 3458 469 3621 521
rect 3673 469 3739 521
rect 3791 469 3804 521
rect 3458 466 3804 469
rect 3735 457 3804 466
rect 2385 430 2551 442
rect 1134 364 1158 416
rect 1210 387 1453 416
rect 1210 364 1232 387
rect -3 296 98 311
rect -285 184 -165 288
rect -285 138 -248 184
rect -202 138 -165 184
rect 1134 247 1232 364
rect 3746 365 3804 457
rect 3746 313 3749 365
rect 3801 313 3804 365
rect 3746 297 3804 313
rect 3859 444 3979 548
rect 3859 398 3894 444
rect 3940 398 3979 444
rect 1134 195 1158 247
rect 1210 195 1232 247
rect 1134 174 1232 195
rect 3859 294 3979 398
rect 3859 248 3894 294
rect 3940 248 3979 294
rect -285 34 -165 138
rect 3859 144 3979 248
rect -285 -12 -248 34
rect -202 -12 -165 34
rect -285 -73 -165 -12
rect -285 -74 46 -73
rect 197 -74 304 107
rect 681 -74 786 105
rect 1054 3 2632 91
rect 1657 -74 1747 3
rect 2451 -74 2539 3
rect 2926 -74 3031 107
rect 3859 98 3894 144
rect 3940 98 3979 144
rect 3859 -6 3979 98
rect 3859 -52 3894 -6
rect 3940 -52 3979 -6
rect 3859 -74 3979 -52
rect -285 -112 3979 -74
rect -285 -158 -129 -112
rect -83 -158 21 -112
rect 67 -158 171 -112
rect 217 -158 321 -112
rect 367 -158 471 -112
rect 517 -158 621 -112
rect 667 -158 771 -112
rect 817 -158 921 -112
rect 967 -158 1071 -112
rect 1117 -158 1221 -112
rect 1267 -158 1371 -112
rect 1417 -158 1521 -112
rect 1567 -158 1671 -112
rect 1717 -158 1821 -112
rect 1867 -158 1971 -112
rect 2017 -158 2121 -112
rect 2167 -158 2271 -112
rect 2317 -158 2421 -112
rect 2467 -158 2571 -112
rect 2617 -158 2721 -112
rect 2767 -158 2871 -112
rect 2917 -158 3021 -112
rect 3067 -158 3171 -112
rect 3217 -158 3321 -112
rect 3367 -158 3471 -112
rect 3517 -158 3621 -112
rect 3667 -158 3771 -112
rect 3817 -158 3979 -112
rect -285 -193 3979 -158
rect -17 -324 392 -297
rect -17 -325 156 -324
rect -17 -377 21 -325
rect 73 -376 156 -325
rect 208 -325 392 -324
rect 208 -376 281 -325
rect 73 -377 281 -376
rect 333 -377 392 -325
rect -17 -403 392 -377
rect 794 -302 972 -301
rect 794 -326 1248 -302
rect 794 -378 866 -326
rect 918 -378 1007 -326
rect 1059 -378 1158 -326
rect 1210 -378 1248 -326
rect 794 -410 1248 -378
rect 3327 -367 3845 -327
rect 3327 -368 3568 -367
rect 794 -413 972 -410
rect 3327 -420 3419 -368
rect 3471 -419 3568 -368
rect 3620 -369 3845 -367
rect 3620 -419 3750 -369
rect 3471 -420 3750 -419
rect 3327 -421 3750 -420
rect 3802 -421 3845 -369
rect 3327 -452 3845 -421
<< via1 >>
rect 1821 2134 1873 2186
rect -60 1144 -8 1196
rect 3726 1286 3778 1338
rect 3724 1101 3776 1153
rect -67 987 -15 1039
rect 21 467 73 519
rect 21 311 73 363
rect 3621 469 3673 521
rect 3739 469 3791 521
rect 1158 364 1210 416
rect 3749 313 3801 365
rect 1158 195 1210 247
rect 21 -377 73 -325
rect 156 -376 208 -324
rect 281 -377 333 -325
rect 866 -378 918 -326
rect 1007 -378 1059 -326
rect 1158 -378 1210 -326
rect 3419 -420 3471 -368
rect 3568 -419 3620 -367
rect 3750 -421 3802 -369
<< metal2 >>
rect 1789 2186 1905 2227
rect 1789 2134 1821 2186
rect 1873 2134 1905 2186
rect 1789 2098 1905 2134
rect 1799 1868 1896 2098
rect -73 1771 3799 1868
rect -69 1217 28 1771
rect 3702 1399 3799 1771
rect -82 1196 28 1217
rect -82 1144 -60 1196
rect -8 1144 28 1196
rect 3691 1338 3810 1399
rect 3691 1286 3726 1338
rect 3778 1286 3810 1338
rect 3691 1190 3810 1286
rect -82 1084 28 1144
rect 3692 1153 3810 1190
rect 3692 1101 3724 1153
rect 3776 1101 3810 1153
rect 3692 1099 3810 1101
rect -82 1044 67 1084
rect 3659 1076 3810 1099
rect -82 1039 78 1044
rect -82 987 -67 1039
rect -15 987 78 1039
rect -82 982 78 987
rect -82 971 67 982
rect 3659 969 3809 1076
rect -3 519 98 543
rect -3 467 21 519
rect 73 467 98 519
rect 3613 521 3816 539
rect -3 363 98 467
rect -3 311 21 363
rect 73 311 98 363
rect -3 296 98 311
rect 1134 416 1232 512
rect 3613 469 3621 521
rect 3673 469 3739 521
rect 3791 469 3816 521
rect 3613 455 3816 469
rect 1134 364 1158 416
rect 1210 364 1232 416
rect 3736 384 3816 455
rect 11 -297 83 296
rect 1134 247 1232 364
rect 1134 195 1158 247
rect 1210 195 1232 247
rect 1134 174 1232 195
rect 3731 365 3822 384
rect 3731 313 3749 365
rect 3801 313 3822 365
rect -17 -324 369 -297
rect 1146 -302 1222 174
rect -17 -325 156 -324
rect -17 -377 21 -325
rect 73 -376 156 -325
rect 208 -325 369 -324
rect 208 -376 281 -325
rect 73 -377 281 -376
rect 333 -377 369 -325
rect -17 -403 369 -377
rect 826 -326 1248 -302
rect 826 -378 866 -326
rect 918 -378 1007 -326
rect 1059 -378 1158 -326
rect 1210 -378 1248 -326
rect 3731 -327 3822 313
rect 826 -410 1248 -378
rect 3378 -367 3845 -327
rect 3378 -368 3568 -367
rect 3378 -420 3419 -368
rect 3471 -419 3568 -368
rect 3620 -369 3845 -367
rect 3620 -419 3750 -369
rect 3471 -420 3750 -419
rect 3378 -421 3750 -420
rect 3802 -421 3845 -369
rect 3378 -452 3845 -421
use INV_2  INV_2_0
timestamp 1713185578
transform 1 0 1311 0 1 486
box 21 -485 1081 648
use Tr_Gate  Tr_Gate_0
timestamp 1713185578
transform -1 0 1154 0 1 1233
box -53 -1233 1187 569
use Tr_Gate  Tr_Gate_1
timestamp 1713185578
transform 1 0 2558 0 1 1235
box -53 -1233 1187 569
<< labels >>
flabel metal1 s 811 -359 811 -359 0 FreeSans 1250 0 0 0 SEL
port 1 nsew
flabel metal1 s 3355 -397 3355 -397 0 FreeSans 1250 0 0 0 IN1
port 2 nsew
flabel metal1 s 377 -354 377 -354 0 FreeSans 1250 0 0 0 IN2
port 3 nsew
flabel metal1 s 1705 1747 1705 1747 0 FreeSans 1250 0 0 0 VDD
port 4 nsew
flabel metal1 s 1288 27 1288 27 0 FreeSans 1250 0 0 0 VSS
port 5 nsew
flabel metal1 s 1728 2158 1728 2158 0 FreeSans 1250 0 0 0 OUT
port 6 nsew
<< end >>
