magic
tech gf180mcuC
magscale 1 10
timestamp 1693548584
<< error_p >>
rect -2063 -48 -2017 48
rect -1859 -48 -1813 48
rect -1655 -48 -1609 48
rect -1451 -48 -1405 48
rect -1247 -48 -1201 48
rect -1043 -48 -997 48
rect -839 -48 -793 48
rect -635 -48 -589 48
rect -431 -48 -385 48
rect -227 -48 -181 48
rect -23 -48 23 48
rect 181 -48 227 48
rect 385 -48 431 48
rect 589 -48 635 48
rect 793 -48 839 48
rect 997 -48 1043 48
rect 1201 -48 1247 48
rect 1405 -48 1451 48
rect 1609 -48 1655 48
rect 1813 -48 1859 48
rect 2017 -48 2063 48
<< nwell >>
rect -2162 -180 2162 180
<< pmos >>
rect -1988 -50 -1888 50
rect -1784 -50 -1684 50
rect -1580 -50 -1480 50
rect -1376 -50 -1276 50
rect -1172 -50 -1072 50
rect -968 -50 -868 50
rect -764 -50 -664 50
rect -560 -50 -460 50
rect -356 -50 -256 50
rect -152 -50 -52 50
rect 52 -50 152 50
rect 256 -50 356 50
rect 460 -50 560 50
rect 664 -50 764 50
rect 868 -50 968 50
rect 1072 -50 1172 50
rect 1276 -50 1376 50
rect 1480 -50 1580 50
rect 1684 -50 1784 50
rect 1888 -50 1988 50
<< pdiff >>
rect -2076 37 -1988 50
rect -2076 -37 -2063 37
rect -2017 -37 -1988 37
rect -2076 -50 -1988 -37
rect -1888 37 -1784 50
rect -1888 -37 -1859 37
rect -1813 -37 -1784 37
rect -1888 -50 -1784 -37
rect -1684 37 -1580 50
rect -1684 -37 -1655 37
rect -1609 -37 -1580 37
rect -1684 -50 -1580 -37
rect -1480 37 -1376 50
rect -1480 -37 -1451 37
rect -1405 -37 -1376 37
rect -1480 -50 -1376 -37
rect -1276 37 -1172 50
rect -1276 -37 -1247 37
rect -1201 -37 -1172 37
rect -1276 -50 -1172 -37
rect -1072 37 -968 50
rect -1072 -37 -1043 37
rect -997 -37 -968 37
rect -1072 -50 -968 -37
rect -868 37 -764 50
rect -868 -37 -839 37
rect -793 -37 -764 37
rect -868 -50 -764 -37
rect -664 37 -560 50
rect -664 -37 -635 37
rect -589 -37 -560 37
rect -664 -50 -560 -37
rect -460 37 -356 50
rect -460 -37 -431 37
rect -385 -37 -356 37
rect -460 -50 -356 -37
rect -256 37 -152 50
rect -256 -37 -227 37
rect -181 -37 -152 37
rect -256 -50 -152 -37
rect -52 37 52 50
rect -52 -37 -23 37
rect 23 -37 52 37
rect -52 -50 52 -37
rect 152 37 256 50
rect 152 -37 181 37
rect 227 -37 256 37
rect 152 -50 256 -37
rect 356 37 460 50
rect 356 -37 385 37
rect 431 -37 460 37
rect 356 -50 460 -37
rect 560 37 664 50
rect 560 -37 589 37
rect 635 -37 664 37
rect 560 -50 664 -37
rect 764 37 868 50
rect 764 -37 793 37
rect 839 -37 868 37
rect 764 -50 868 -37
rect 968 37 1072 50
rect 968 -37 997 37
rect 1043 -37 1072 37
rect 968 -50 1072 -37
rect 1172 37 1276 50
rect 1172 -37 1201 37
rect 1247 -37 1276 37
rect 1172 -50 1276 -37
rect 1376 37 1480 50
rect 1376 -37 1405 37
rect 1451 -37 1480 37
rect 1376 -50 1480 -37
rect 1580 37 1684 50
rect 1580 -37 1609 37
rect 1655 -37 1684 37
rect 1580 -50 1684 -37
rect 1784 37 1888 50
rect 1784 -37 1813 37
rect 1859 -37 1888 37
rect 1784 -50 1888 -37
rect 1988 37 2076 50
rect 1988 -37 2017 37
rect 2063 -37 2076 37
rect 1988 -50 2076 -37
<< pdiffc >>
rect -2063 -37 -2017 37
rect -1859 -37 -1813 37
rect -1655 -37 -1609 37
rect -1451 -37 -1405 37
rect -1247 -37 -1201 37
rect -1043 -37 -997 37
rect -839 -37 -793 37
rect -635 -37 -589 37
rect -431 -37 -385 37
rect -227 -37 -181 37
rect -23 -37 23 37
rect 181 -37 227 37
rect 385 -37 431 37
rect 589 -37 635 37
rect 793 -37 839 37
rect 997 -37 1043 37
rect 1201 -37 1247 37
rect 1405 -37 1451 37
rect 1609 -37 1655 37
rect 1813 -37 1859 37
rect 2017 -37 2063 37
<< polysilicon >>
rect -1988 50 -1888 94
rect -1784 50 -1684 94
rect -1580 50 -1480 94
rect -1376 50 -1276 94
rect -1172 50 -1072 94
rect -968 50 -868 94
rect -764 50 -664 94
rect -560 50 -460 94
rect -356 50 -256 94
rect -152 50 -52 94
rect 52 50 152 94
rect 256 50 356 94
rect 460 50 560 94
rect 664 50 764 94
rect 868 50 968 94
rect 1072 50 1172 94
rect 1276 50 1376 94
rect 1480 50 1580 94
rect 1684 50 1784 94
rect 1888 50 1988 94
rect -1988 -94 -1888 -50
rect -1784 -94 -1684 -50
rect -1580 -94 -1480 -50
rect -1376 -94 -1276 -50
rect -1172 -94 -1072 -50
rect -968 -94 -868 -50
rect -764 -94 -664 -50
rect -560 -94 -460 -50
rect -356 -94 -256 -50
rect -152 -94 -52 -50
rect 52 -94 152 -50
rect 256 -94 356 -50
rect 460 -94 560 -50
rect 664 -94 764 -50
rect 868 -94 968 -50
rect 1072 -94 1172 -50
rect 1276 -94 1376 -50
rect 1480 -94 1580 -50
rect 1684 -94 1784 -50
rect 1888 -94 1988 -50
<< metal1 >>
rect -2063 37 -2017 48
rect -2063 -48 -2017 -37
rect -1859 37 -1813 48
rect -1859 -48 -1813 -37
rect -1655 37 -1609 48
rect -1655 -48 -1609 -37
rect -1451 37 -1405 48
rect -1451 -48 -1405 -37
rect -1247 37 -1201 48
rect -1247 -48 -1201 -37
rect -1043 37 -997 48
rect -1043 -48 -997 -37
rect -839 37 -793 48
rect -839 -48 -793 -37
rect -635 37 -589 48
rect -635 -48 -589 -37
rect -431 37 -385 48
rect -431 -48 -385 -37
rect -227 37 -181 48
rect -227 -48 -181 -37
rect -23 37 23 48
rect -23 -48 23 -37
rect 181 37 227 48
rect 181 -48 227 -37
rect 385 37 431 48
rect 385 -48 431 -37
rect 589 37 635 48
rect 589 -48 635 -37
rect 793 37 839 48
rect 793 -48 839 -37
rect 997 37 1043 48
rect 997 -48 1043 -37
rect 1201 37 1247 48
rect 1201 -48 1247 -37
rect 1405 37 1451 48
rect 1405 -48 1451 -37
rect 1609 37 1655 48
rect 1609 -48 1655 -37
rect 1813 37 1859 48
rect 1813 -48 1859 -37
rect 2017 37 2063 48
rect 2017 -48 2063 -37
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.5 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
