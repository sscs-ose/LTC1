magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1461 -1019 1461 1019
<< metal1 >>
rect -461 13 461 19
rect -461 -13 -455 13
rect 455 -13 461 13
rect -461 -19 461 -13
<< via1 >>
rect -455 -13 455 13
<< metal2 >>
rect -461 13 461 19
rect -461 -13 -455 13
rect 455 -13 461 13
rect -461 -19 461 -13
<< end >>
