* NGSPICE file created from filter_res_magic_flat.ext - technology: gf180mcuC

.subckt filter_res_magic_flat R7_R8_R10_C R3_R7 VDD VIN_N VIN_P VOUT_OPAMP_N VOUT_OPAMP_P
+ VOUT_N VOUT_P
X0 a_947_715.t0 a_1507_153.t0 VDD.t18 ppolyf_u r_width=1u r_length=2.3u
X1 VDD.t28 VDD.t29 VDD.t23 ppolyf_u r_width=1u r_length=2.3u
X2 VOUT_OPAMP_N.t0 VOUT_OPAMP_N.t1 VDD.t9 ppolyf_u r_width=1u r_length=2.3u
X3 VDD.t19 VDD.t20 VDD.t2 ppolyf_u r_width=1u r_length=2.3u
X4 VDD.t21 VDD.t22 VDD.t2 ppolyf_u r_width=1u r_length=2.3u
X5 VOUT_N.t1 VOUT_OPAMP_P.t6 cap_mim_2f0_m4m5_noshield c_width=15.2u c_length=16u
X6 a_387_n202.t2 R3_R7.t7 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X7 VDD.t26 VDD.t27 VDD.t23 ppolyf_u r_width=1u r_length=2.3u
X8 a_667_n202.t1 a_387_n1119.t2 VDD.t7 ppolyf_u r_width=1u r_length=2.3u
X9 VDD.t24 VDD.t25 VDD.t23 ppolyf_u r_width=1u r_length=2.3u
X10 a_387_n3450.t0 R3_R7.t1 VDD.t5 ppolyf_u r_width=1u r_length=2.3u
X11 a_387_n202.t1 a_667_153.t1 VDD.t7 ppolyf_u r_width=1u r_length=2.3u
X12 a_667_n1119.t1 a_387_n1681.t1 VDD.t7 ppolyf_u r_width=1u r_length=2.3u
X13 VDD.t15 VDD.t16 VDD.t2 ppolyf_u r_width=1u r_length=2.3u
X14 R7_R8_R10_C.t3 a_387_n1119.t3 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X15 VDD.t30 VDD.t31 VDD.t23 ppolyf_u r_width=1u r_length=2.3u
X16 VIN_N.t0 a_1507_n4012.t1 VDD.t9 ppolyf_u r_width=1u r_length=2.3u
X17 a_387_n4367.t1 a_947_n4929.t0 VDD.t1 ppolyf_u r_width=1u r_length=2.3u
X18 a_387_n202.t3 R3_R7.t6 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X19 VOUT_OPAMP_P.t0 VOUT_OPAMP_P.t1 VDD.t17 ppolyf_u r_width=1u r_length=2.3u
X20 a_387_n2533.t1 a_667_n3095.t1 VDD.t7 ppolyf_u r_width=1u r_length=2.3u
X21 a_667_n4367.t1 a_1227_n4929.t1 VDD.t8 ppolyf_u r_width=1u r_length=2.3u
X22 a_387_n202.t0 a_387_n764.t1 VDD.t5 ppolyf_u r_width=1u r_length=2.3u
X23 VDD.t34 VDD.t35 VDD.t23 ppolyf_u r_width=1u r_length=2.3u
X24 VOUT_OPAMP_N.t2 VOUT_OPAMP_N.t3 VDD.t17 ppolyf_u r_width=1u r_length=2.3u
X25 a_1787_n4367.t0 a_1227_n4929.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X26 VOUT_P.t1 VOUT_OPAMP_N.t4 cap_mim_2f0_m4m5_noshield c_width=15.2u c_length=16u
X27 R7_R8_R10_C.t0 a_667_n4012.t0 VDD.t7 ppolyf_u r_width=1u r_length=2.3u
X28 a_387_n202.t3 R3_R7.t5 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X29 a_667_n1119.t0 a_947_n1681.t0 VDD.t1 ppolyf_u r_width=1u r_length=2.3u
X30 VOUT_N.t2 VOUT_OPAMP_P.t5 cap_mim_2f0_m4m5_noshield c_width=15.2u c_length=16u
X31 a_1227_n1119.t0 a_947_n1681.t1 VDD.t8 ppolyf_u r_width=1u r_length=2.3u
X32 a_2347_n3450.t1 a_2627_n4367.t0 VDD.t17 ppolyf_u r_width=1u r_length=2.3u
X33 a_387_n202.t3 R3_R7.t4 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X34 VOUT_P.t2 VOUT_OPAMP_N.t5 cap_mim_2f0_m4m5_noshield c_width=15.2u c_length=16u
X35 a_2347_715.t0 a_1787_153.t0 VDD.t6 ppolyf_u r_width=1u r_length=2.3u
X36 a_1507_n4367.t1 a_947_n4929.t1 VDD.t18 ppolyf_u r_width=1u r_length=2.3u
X37 a_1507_n4367.t0 a_2067_n4929.t1 VDD.t12 ppolyf_u r_width=1u r_length=2.3u
X38 a_1227_715.t1 a_1787_153.t1 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X39 a_947_n2533.t0 a_667_n3095.t0 VDD.t1 ppolyf_u r_width=1u r_length=2.3u
X40 a_1227_715.t0 a_667_153.t0 VDD.t8 ppolyf_u r_width=1u r_length=2.3u
X41 a_1787_n1119.t1 a_1507_n1681.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X42 a_947_n2533.t1 a_1227_n3095.t1 VDD.t8 ppolyf_u r_width=1u r_length=2.3u
X43 a_387_n202.t3 R3_R7.t3 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X44 VOUT_N.t0 a_387_153.t0 VDD.t5 ppolyf_u r_width=1u r_length=2.3u
X45 a_947_n3450.t0 R7_R8_R10_C.t2 VDD.t1 ppolyf_u r_width=1u r_length=2.3u
X46 a_1787_n1119.t0 a_2067_n1681.t0 VDD.t12 ppolyf_u r_width=1u r_length=2.3u
X47 a_1507_n2533.t0 a_1787_n3095.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X48 a_1227_n3450.t1 a_667_n4012.t1 VDD.t8 ppolyf_u r_width=1u r_length=2.3u
X49 a_1227_n1119.t1 a_1507_n1681.t1 VDD.t18 ppolyf_u r_width=1u r_length=2.3u
X50 a_1787_n4367.t1 a_2347_n4929.t1 VDD.t6 ppolyf_u r_width=1u r_length=2.3u
X51 a_2347_715.t1 a_2067_n202.t1 VDD.t17 ppolyf_u r_width=1u r_length=2.3u
X52 a_2627_153.t0 a_2347_n764.t1 VDD.t17 ppolyf_u r_width=1u r_length=2.3u
X53 a_2067_n2533.t0 a_1787_n3095.t1 VDD.t12 ppolyf_u r_width=1u r_length=2.3u
X54 a_1227_n3450.t0 a_1787_n4012.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X55 a_1507_n2533.t1 a_1227_n3095.t0 VDD.t18 ppolyf_u r_width=1u r_length=2.3u
X56 VDD.t13 VDD.t14 VDD.t2 ppolyf_u r_width=1u r_length=2.3u
X57 a_1507_n202.t1 a_387_n764.t0 VDD.t18 ppolyf_u r_width=1u r_length=2.3u
X58 R7_R8_R10_C.t4 a_387_n1119.t4 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X59 a_947_715.t1 a_387_153.t1 VDD.t1 ppolyf_u r_width=1u r_length=2.3u
X60 a_947_n3450.t1 a_2067_n4012.t1 VDD.t12 ppolyf_u r_width=1u r_length=2.3u
X61 a_387_n4367.t0 VOUT_P.t0 VDD.t5 ppolyf_u r_width=1u r_length=2.3u
X62 a_2067_715.t0 a_1507_153.t1 VDD.t12 ppolyf_u r_width=1u r_length=2.3u
X63 a_1507_n202.t0 VIN_P.t0 VDD.t9 ppolyf_u r_width=1u r_length=2.3u
X64 VOUT_OPAMP_P.t4 a_2067_n1681.t1 VDD.t6 ppolyf_u r_width=1u r_length=2.3u
X65 a_387_n3450.t1 a_1507_n4012.t0 VDD.t18 ppolyf_u r_width=1u r_length=2.3u
X66 VDD.t3 VDD.t4 VDD.t2 ppolyf_u r_width=1u r_length=2.3u
X67 a_2627_n4367.t1 a_2067_n4929.t0 VDD.t9 ppolyf_u r_width=1u r_length=2.3u
X68 a_667_n202.t0 a_1227_n764.t0 VDD.t8 ppolyf_u r_width=1u r_length=2.3u
X69 a_1787_n202.t1 a_1227_n764.t1 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X70 a_2067_n2533.t1 VOUT_OPAMP_N.t6 VDD.t6 ppolyf_u r_width=1u r_length=2.3u
X71 VDD.t32 VDD.t33 VDD.t23 ppolyf_u r_width=1u r_length=2.3u
X72 a_1787_n202.t0 a_2347_n764.t0 VDD.t6 ppolyf_u r_width=1u r_length=2.3u
X73 a_387_n1119.t0 a_387_n1681.t0 VDD.t5 ppolyf_u r_width=1u r_length=2.3u
X74 VDD.t10 VDD.t11 VDD.t2 ppolyf_u r_width=1u r_length=2.3u
X75 a_2347_n3450.t0 a_1787_n4012.t1 VDD.t6 ppolyf_u r_width=1u r_length=2.3u
X76 a_667_n4367.t0 R3_R7.t0 VDD.t7 ppolyf_u r_width=1u r_length=2.3u
X77 a_387_n202.t2 R3_R7.t2 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X78 a_2067_715.t1 a_2627_153.t1 VDD.t9 ppolyf_u r_width=1u r_length=2.3u
X79 a_387_n1119.t1 a_947_n764.t0 VDD.t1 ppolyf_u r_width=1u r_length=2.3u
X80 VOUT_OPAMP_P.t2 VOUT_OPAMP_P.t3 VDD.t9 ppolyf_u r_width=1u r_length=2.3u
X81 a_387_n2533.t0 R7_R8_R10_C.t1 VDD.t5 ppolyf_u r_width=1u r_length=2.3u
X82 a_2067_n202.t0 a_947_n764.t1 VDD.t12 ppolyf_u r_width=1u r_length=2.3u
X83 a_2067_n4012.t0 a_2347_n4929.t0 VDD.t17 ppolyf_u r_width=1u r_length=2.3u
R0 a_947_715.t0 a_947_715.t1 13.5425
R1 a_1507_153.t0 a_1507_153.t1 13.5425
R2 VDD.n459 VDD.t24 6.87803
R3 VDD.n446 VDD.t25 6.87803
R4 VDD.n440 VDD.t34 6.87803
R5 VDD.n433 VDD.t35 6.87803
R6 VDD.n421 VDD.t33 6.87803
R7 VDD.n535 VDD.t30 6.87803
R8 VDD.n509 VDD.t26 6.87803
R9 VDD.n496 VDD.t27 6.87803
R10 VDD.n489 VDD.t28 6.87803
R11 VDD.n476 VDD.t29 6.87803
R12 VDD.n428 VDD.t32 6.87615
R13 VDD.n519 VDD.t31 6.87615
R14 VDD.n278 VDD.t2 6.83492
R15 VDD.n649 VDD.t8 6.83492
R16 VDD.n137 VDD.t11 6.82906
R17 VDD.n150 VDD.t10 6.82906
R18 VDD.n157 VDD.t22 6.82906
R19 VDD.n176 VDD.t21 6.82906
R20 VDD.n189 VDD.t14 6.82906
R21 VDD.n208 VDD.t13 6.82906
R22 VDD.n22 VDD.t4 6.82906
R23 VDD.n29 VDD.t3 6.82906
R24 VDD.n34 VDD.t16 6.82906
R25 VDD.n42 VDD.t15 6.82906
R26 VDD.n49 VDD.t20 6.82906
R27 VDD.n62 VDD.t19 6.82906
R28 VDD.n286 VDD.t17 6.21361
R29 VDD.n641 VDD.t1 6.21361
R30 VDD.n661 VDD.t18 4.66033
R31 VDD.n298 VDD.t9 4.03902
R32 VDD.n629 VDD.t7 4.03902
R33 VDD.n467 VDD.n466 3.1505
R34 VDD.n68 VDD.n67 3.1505
R35 VDD.n463 VDD.n462 3.1505
R36 VDD.n461 VDD.n460 3.1505
R37 VDD.n458 VDD.n457 3.1505
R38 VDD.n456 VDD.n455 3.1505
R39 VDD.n454 VDD.n453 3.1505
R40 VDD.n452 VDD.n451 3.1505
R41 VDD.n450 VDD.n449 3.1505
R42 VDD.n448 VDD.n447 3.1505
R43 VDD.n445 VDD.n444 3.1505
R44 VDD.n443 VDD.n442 3.1505
R45 VDD.n465 VDD.n464 3.1505
R46 VDD.n70 VDD.n69 3.1505
R47 VDD.n127 VDD.n125 3.1505
R48 VDD.n124 VDD.n122 3.1505
R49 VDD.n121 VDD.n119 3.1505
R50 VDD.n118 VDD.n116 3.1505
R51 VDD.n115 VDD.n113 3.1505
R52 VDD.n112 VDD.n110 3.1505
R53 VDD.n109 VDD.n107 3.1505
R54 VDD.n106 VDD.n104 3.1505
R55 VDD.n103 VDD.n101 3.1505
R56 VDD.n100 VDD.n98 3.1505
R57 VDD.n97 VDD.n95 3.1505
R58 VDD.n94 VDD.n92 3.1505
R59 VDD.n91 VDD.n89 3.1505
R60 VDD.n88 VDD.n86 3.1505
R61 VDD.n85 VDD.n83 3.1505
R62 VDD.n82 VDD.n80 3.1505
R63 VDD.n79 VDD.n77 3.1505
R64 VDD.n76 VDD.n74 3.1505
R65 VDD.n73 VDD.n71 3.1505
R66 VDD.n344 VDD.n342 3.1505
R67 VDD.n347 VDD.n345 3.1505
R68 VDD.n350 VDD.n348 3.1505
R69 VDD.n353 VDD.n351 3.1505
R70 VDD.n356 VDD.n354 3.1505
R71 VDD.n359 VDD.n357 3.1505
R72 VDD.n362 VDD.n360 3.1505
R73 VDD.n365 VDD.n363 3.1505
R74 VDD.n368 VDD.n366 3.1505
R75 VDD.n371 VDD.n369 3.1505
R76 VDD.n374 VDD.n372 3.1505
R77 VDD.n377 VDD.n375 3.1505
R78 VDD.n380 VDD.n378 3.1505
R79 VDD.n383 VDD.n381 3.1505
R80 VDD.n386 VDD.n384 3.1505
R81 VDD.n389 VDD.n387 3.1505
R82 VDD.n392 VDD.n390 3.1505
R83 VDD.n395 VDD.n393 3.1505
R84 VDD.n398 VDD.n396 3.1505
R85 VDD.n66 VDD.n65 3.1505
R86 VDD.n64 VDD.n63 3.1505
R87 VDD.n61 VDD.n60 3.1505
R88 VDD.n59 VDD.n58 3.1505
R89 VDD.n57 VDD.n56 3.1505
R90 VDD.n55 VDD.n54 3.1505
R91 VDD.n53 VDD.n52 3.1505
R92 VDD.n51 VDD.n50 3.1505
R93 VDD.n48 VDD.n47 3.1505
R94 VDD.n46 VDD.n45 3.1505
R95 VDD.n44 VDD.n43 3.1505
R96 VDD.n41 VDD.n40 3.1505
R97 VDD.n266 VDD.n265 3.1505
R98 VDD.n270 VDD.n269 3.1505
R99 VDD.n274 VDD.n273 3.1505
R100 VDD.n278 VDD.n277 3.1505
R101 VDD.n282 VDD.n281 3.1505
R102 VDD.n286 VDD.n285 3.1505
R103 VDD.n290 VDD.n289 3.1505
R104 VDD.n294 VDD.n293 3.1505
R105 VDD.n298 VDD.n297 3.1505
R106 VDD.n302 VDD.n301 3.1505
R107 VDD.n306 VDD.n305 3.1505
R108 VDD.n310 VDD.n309 3.1505
R109 VDD.n314 VDD.n313 3.1505
R110 VDD.n318 VDD.n317 3.1505
R111 VDD.n322 VDD.n321 3.1505
R112 VDD.n326 VDD.n325 3.1505
R113 VDD.n330 VDD.n329 3.1505
R114 VDD.n334 VDD.n333 3.1505
R115 VDD.n338 VDD.n337 3.1505
R116 VDD.n665 VDD.n664 3.1505
R117 VDD.n661 VDD.n660 3.1505
R118 VDD.n657 VDD.n656 3.1505
R119 VDD.n653 VDD.n652 3.1505
R120 VDD.n649 VDD.n648 3.1505
R121 VDD.n645 VDD.n644 3.1505
R122 VDD.n641 VDD.n640 3.1505
R123 VDD.n637 VDD.n636 3.1505
R124 VDD.n633 VDD.n632 3.1505
R125 VDD.n629 VDD.n628 3.1505
R126 VDD.n625 VDD.n624 3.1505
R127 VDD.n621 VDD.n620 3.1505
R128 VDD.n617 VDD.n616 3.1505
R129 VDD.n613 VDD.n612 3.1505
R130 VDD.n609 VDD.n608 3.1505
R131 VDD.n605 VDD.n604 3.1505
R132 VDD.n601 VDD.n600 3.1505
R133 VDD.n597 VDD.n596 3.1505
R134 VDD.n593 VDD.n592 3.1505
R135 VDD.n471 VDD.n341 3.1505
R136 VDD.n538 VDD.n537 3.1505
R137 VDD.n534 VDD.n533 3.1505
R138 VDD.n532 VDD.n531 3.1505
R139 VDD.n529 VDD.n528 3.1505
R140 VDD.n527 VDD.n526 3.1505
R141 VDD.n524 VDD.n523 3.1505
R142 VDD.n522 VDD.n521 3.1505
R143 VDD.n518 VDD.n517 3.1505
R144 VDD.n516 VDD.n515 3.1505
R145 VDD.n513 VDD.n512 3.1505
R146 VDD.n511 VDD.n510 3.1505
R147 VDD.n508 VDD.n507 3.1505
R148 VDD.n506 VDD.n505 3.1505
R149 VDD.n504 VDD.n503 3.1505
R150 VDD.n502 VDD.n501 3.1505
R151 VDD.n500 VDD.n499 3.1505
R152 VDD.n498 VDD.n497 3.1505
R153 VDD.n495 VDD.n494 3.1505
R154 VDD.n493 VDD.n492 3.1505
R155 VDD.n491 VDD.n490 3.1505
R156 VDD.n488 VDD.n487 3.1505
R157 VDD.n486 VDD.n485 3.1505
R158 VDD.n484 VDD.n483 3.1505
R159 VDD.n482 VDD.n481 3.1505
R160 VDD.n480 VDD.n479 3.1505
R161 VDD.n478 VDD.n477 3.1505
R162 VDD.n475 VDD.n474 3.1505
R163 VDD.n473 VDD.n472 3.1505
R164 VDD.n540 VDD.n539 3.1505
R165 VDD.n470 VDD.n469 3.1505
R166 VDD.n127 VDD.n126 3.1505
R167 VDD.n124 VDD.n123 3.1505
R168 VDD.n121 VDD.n120 3.1505
R169 VDD.n118 VDD.n117 3.1505
R170 VDD.n115 VDD.n114 3.1505
R171 VDD.n112 VDD.n111 3.1505
R172 VDD.n109 VDD.n108 3.1505
R173 VDD.n106 VDD.n105 3.1505
R174 VDD.n103 VDD.n102 3.1505
R175 VDD.n100 VDD.n99 3.1505
R176 VDD.n97 VDD.n96 3.1505
R177 VDD.n94 VDD.n93 3.1505
R178 VDD.n91 VDD.n90 3.1505
R179 VDD.n88 VDD.n87 3.1505
R180 VDD.n85 VDD.n84 3.1505
R181 VDD.n82 VDD.n81 3.1505
R182 VDD.n79 VDD.n78 3.1505
R183 VDD.n76 VDD.n75 3.1505
R184 VDD.n73 VDD.n72 3.1505
R185 VDD.n344 VDD.n343 3.1505
R186 VDD.n347 VDD.n346 3.1505
R187 VDD.n350 VDD.n349 3.1505
R188 VDD.n353 VDD.n352 3.1505
R189 VDD.n356 VDD.n355 3.1505
R190 VDD.n359 VDD.n358 3.1505
R191 VDD.n362 VDD.n361 3.1505
R192 VDD.n365 VDD.n364 3.1505
R193 VDD.n368 VDD.n367 3.1505
R194 VDD.n371 VDD.n370 3.1505
R195 VDD.n374 VDD.n373 3.1505
R196 VDD.n377 VDD.n376 3.1505
R197 VDD.n380 VDD.n379 3.1505
R198 VDD.n383 VDD.n382 3.1505
R199 VDD.n386 VDD.n385 3.1505
R200 VDD.n389 VDD.n388 3.1505
R201 VDD.n392 VDD.n391 3.1505
R202 VDD.n395 VDD.n394 3.1505
R203 VDD.n398 VDD.n397 3.1505
R204 VDD.n130 VDD.n129 3.1505
R205 VDD.n132 VDD.n131 3.1505
R206 VDD.n134 VDD.n133 3.1505
R207 VDD.n136 VDD.n135 3.1505
R208 VDD.n139 VDD.n138 3.1505
R209 VDD.n141 VDD.n140 3.1505
R210 VDD.n143 VDD.n142 3.1505
R211 VDD.n145 VDD.n144 3.1505
R212 VDD.n147 VDD.n146 3.1505
R213 VDD.n149 VDD.n148 3.1505
R214 VDD.n152 VDD.n151 3.1505
R215 VDD.n154 VDD.n153 3.1505
R216 VDD.n156 VDD.n155 3.1505
R217 VDD.n160 VDD.n159 3.1505
R218 VDD.n163 VDD.n162 3.1505
R219 VDD.n166 VDD.n165 3.1505
R220 VDD.n169 VDD.n168 3.1505
R221 VDD.n172 VDD.n171 3.1505
R222 VDD.n175 VDD.n174 3.1505
R223 VDD.n179 VDD.n178 3.1505
R224 VDD.n182 VDD.n181 3.1505
R225 VDD.n185 VDD.n184 3.1505
R226 VDD.n188 VDD.n187 3.1505
R227 VDD.n192 VDD.n191 3.1505
R228 VDD.n195 VDD.n194 3.1505
R229 VDD.n198 VDD.n197 3.1505
R230 VDD.n201 VDD.n200 3.1505
R231 VDD.n204 VDD.n203 3.1505
R232 VDD.n207 VDD.n206 3.1505
R233 VDD.n211 VDD.n210 3.1505
R234 VDD.n214 VDD.n213 3.1505
R235 VDD.n264 VDD.n263 3.1505
R236 VDD.n268 VDD.n267 3.1505
R237 VDD.n267 VDD.n266 3.1505
R238 VDD.n272 VDD.n271 3.1505
R239 VDD.n271 VDD.n270 3.1505
R240 VDD.n276 VDD.n275 3.1505
R241 VDD.n275 VDD.n274 3.1505
R242 VDD.n280 VDD.n279 3.1505
R243 VDD.n279 VDD.n278 3.1505
R244 VDD.n284 VDD.n283 3.1505
R245 VDD.n283 VDD.n282 3.1505
R246 VDD.n288 VDD.n287 3.1505
R247 VDD.n287 VDD.n286 3.1505
R248 VDD.n292 VDD.n291 3.1505
R249 VDD.n291 VDD.n290 3.1505
R250 VDD.n296 VDD.n295 3.1505
R251 VDD.n295 VDD.n294 3.1505
R252 VDD.n300 VDD.n299 3.1505
R253 VDD.n299 VDD.n298 3.1505
R254 VDD.n304 VDD.n303 3.1505
R255 VDD.n303 VDD.n302 3.1505
R256 VDD.n308 VDD.n307 3.1505
R257 VDD.n307 VDD.n306 3.1505
R258 VDD.n312 VDD.n311 3.1505
R259 VDD.n311 VDD.n310 3.1505
R260 VDD.n316 VDD.n315 3.1505
R261 VDD.n315 VDD.n314 3.1505
R262 VDD.n320 VDD.n319 3.1505
R263 VDD.n319 VDD.n318 3.1505
R264 VDD.n324 VDD.n323 3.1505
R265 VDD.n323 VDD.n322 3.1505
R266 VDD.n328 VDD.n327 3.1505
R267 VDD.n327 VDD.n326 3.1505
R268 VDD.n332 VDD.n331 3.1505
R269 VDD.n331 VDD.n330 3.1505
R270 VDD.n336 VDD.n335 3.1505
R271 VDD.n335 VDD.n334 3.1505
R272 VDD.n340 VDD.n339 3.1505
R273 VDD.n339 VDD.n338 3.1505
R274 VDD.n667 VDD.n666 3.1505
R275 VDD.n666 VDD.n665 3.1505
R276 VDD.n663 VDD.n662 3.1505
R277 VDD.n662 VDD.n661 3.1505
R278 VDD.n659 VDD.n658 3.1505
R279 VDD.n658 VDD.n657 3.1505
R280 VDD.n655 VDD.n654 3.1505
R281 VDD.n654 VDD.n653 3.1505
R282 VDD.n651 VDD.n650 3.1505
R283 VDD.n650 VDD.n649 3.1505
R284 VDD.n647 VDD.n646 3.1505
R285 VDD.n646 VDD.n645 3.1505
R286 VDD.n643 VDD.n642 3.1505
R287 VDD.n642 VDD.n641 3.1505
R288 VDD.n639 VDD.n638 3.1505
R289 VDD.n638 VDD.n637 3.1505
R290 VDD.n635 VDD.n634 3.1505
R291 VDD.n634 VDD.n633 3.1505
R292 VDD.n631 VDD.n630 3.1505
R293 VDD.n630 VDD.n629 3.1505
R294 VDD.n627 VDD.n626 3.1505
R295 VDD.n626 VDD.n625 3.1505
R296 VDD.n623 VDD.n622 3.1505
R297 VDD.n622 VDD.n621 3.1505
R298 VDD.n619 VDD.n618 3.1505
R299 VDD.n618 VDD.n617 3.1505
R300 VDD.n615 VDD.n614 3.1505
R301 VDD.n614 VDD.n613 3.1505
R302 VDD.n611 VDD.n610 3.1505
R303 VDD.n610 VDD.n609 3.1505
R304 VDD.n607 VDD.n606 3.1505
R305 VDD.n606 VDD.n605 3.1505
R306 VDD.n603 VDD.n602 3.1505
R307 VDD.n602 VDD.n601 3.1505
R308 VDD.n599 VDD.n598 3.1505
R309 VDD.n598 VDD.n597 3.1505
R310 VDD.n595 VDD.n594 3.1505
R311 VDD.n594 VDD.n593 3.1505
R312 VDD.n591 VDD.n590 3.1505
R313 VDD.n334 VDD.t0 2.48574
R314 VDD.n213 VDD.n212 2.39402
R315 VDD.n210 VDD.n209 2.39402
R316 VDD.n206 VDD.n205 2.39402
R317 VDD.n203 VDD.n202 2.39402
R318 VDD.n200 VDD.n199 2.39402
R319 VDD.n197 VDD.n196 2.39402
R320 VDD.n194 VDD.n193 2.39402
R321 VDD.n191 VDD.n190 2.39402
R322 VDD.n187 VDD.n186 2.39402
R323 VDD.n184 VDD.n183 2.39402
R324 VDD.n181 VDD.n180 2.39402
R325 VDD.n178 VDD.n177 2.39402
R326 VDD.n174 VDD.n173 2.39402
R327 VDD.n171 VDD.n170 2.39402
R328 VDD.n168 VDD.n167 2.39402
R329 VDD.n165 VDD.n164 2.39402
R330 VDD.n162 VDD.n161 2.39402
R331 VDD.n159 VDD.n158 2.39402
R332 VDD.n585 VDD.n583 2.27972
R333 VDD.n261 VDD.n250 1.95449
R334 VDD.n261 VDD.n251 1.95449
R335 VDD.n261 VDD.n252 1.95449
R336 VDD.n261 VDD.n253 1.95449
R337 VDD.n261 VDD.n254 1.95449
R338 VDD.n261 VDD.n255 1.95449
R339 VDD.n261 VDD.n256 1.95449
R340 VDD.n261 VDD.n257 1.95449
R341 VDD.n261 VDD.n258 1.95449
R342 VDD.n261 VDD.n259 1.95449
R343 VDD.n261 VDD.n260 1.95449
R344 VDD.n310 VDD.t6 1.86443
R345 VDD.n617 VDD.t5 1.86443
R346 VDD.n559 VDD.n557 1.73593
R347 VDD.n562 VDD.n560 1.73593
R348 VDD.n565 VDD.n563 1.73593
R349 VDD.n568 VDD.n566 1.73593
R350 VDD.n571 VDD.n569 1.73593
R351 VDD.n574 VDD.n572 1.73593
R352 VDD.n577 VDD.n575 1.73593
R353 VDD.n580 VDD.n578 1.73593
R354 VDD.n242 VDD.n240 1.73593
R355 VDD.n239 VDD.n237 1.73593
R356 VDD.n236 VDD.n234 1.73593
R357 VDD.n233 VDD.n231 1.73593
R358 VDD.n230 VDD.n228 1.73593
R359 VDD.n227 VDD.n225 1.73593
R360 VDD.n224 VDD.n222 1.73593
R361 VDD.n221 VDD.n219 1.73593
R362 VDD.n242 VDD.n241 1.73541
R363 VDD.n239 VDD.n238 1.73541
R364 VDD.n236 VDD.n235 1.73541
R365 VDD.n233 VDD.n232 1.73541
R366 VDD.n230 VDD.n229 1.73541
R367 VDD.n227 VDD.n226 1.73541
R368 VDD.n224 VDD.n223 1.73541
R369 VDD.n221 VDD.n220 1.73541
R370 VDD.n580 VDD.n579 1.73541
R371 VDD.n577 VDD.n576 1.73541
R372 VDD.n574 VDD.n573 1.73541
R373 VDD.n571 VDD.n570 1.73541
R374 VDD.n568 VDD.n567 1.73541
R375 VDD.n565 VDD.n564 1.73541
R376 VDD.n562 VDD.n561 1.73541
R377 VDD.n559 VDD.n558 1.73541
R378 VDD.n556 VDD.n555 1.73541
R379 VDD.n537 VDD.n536 1.73527
R380 VDD.n531 VDD.n530 1.73527
R381 VDD.n526 VDD.n525 1.73527
R382 VDD.n521 VDD.n520 1.73527
R383 VDD.n515 VDD.n514 1.73527
R384 VDD.n218 VDD.n216 1.44895
R385 VDD.n218 VDD.n217 1.44847
R386 VDD.n590 VDD.n589 1.4483
R387 VDD.n582 VDD.n581 1.41705
R388 VDD.n588 VDD.n586 1.41673
R389 VDD.n261 VDD.n215 1.41673
R390 VDD.n262 VDD.n261 1.3416
R391 VDD.n588 VDD.n585 1.34143
R392 VDD.n588 VDD.n550 1.15696
R393 VDD.n588 VDD.n582 1.15696
R394 VDD.n263 VDD.n262 1.14056
R395 VDD.n585 VDD.n584 1.14036
R396 VDD.n261 VDD.n249 0.914272
R397 VDD.n588 VDD.n587 0.914044
R398 VDD.n261 VDD.n218 0.852583
R399 VDD.n589 VDD.n588 0.852351
R400 VDD.n588 VDD.n551 0.709103
R401 VDD.n588 VDD.n552 0.709103
R402 VDD.n588 VDD.n553 0.709103
R403 VDD.n588 VDD.n554 0.709103
R404 VDD.n588 VDD.n556 0.709103
R405 VDD.n588 VDD.n559 0.709103
R406 VDD.n588 VDD.n562 0.709103
R407 VDD.n588 VDD.n565 0.709103
R408 VDD.n588 VDD.n568 0.709103
R409 VDD.n588 VDD.n571 0.709103
R410 VDD.n588 VDD.n574 0.709103
R411 VDD.n588 VDD.n577 0.709103
R412 VDD.n588 VDD.n580 0.709103
R413 VDD.n261 VDD.n248 0.709103
R414 VDD.n261 VDD.n247 0.709103
R415 VDD.n261 VDD.n246 0.709103
R416 VDD.n261 VDD.n245 0.709103
R417 VDD.n261 VDD.n244 0.709103
R418 VDD.n261 VDD.n243 0.709103
R419 VDD.n261 VDD.n242 0.709103
R420 VDD.n261 VDD.n239 0.709103
R421 VDD.n261 VDD.n236 0.709103
R422 VDD.n261 VDD.n233 0.709103
R423 VDD.n261 VDD.n230 0.709103
R424 VDD.n261 VDD.n227 0.709103
R425 VDD.n261 VDD.n224 0.709103
R426 VDD.n261 VDD.n221 0.709103
R427 VDD.n588 VDD.n549 0.708865
R428 VDD.n588 VDD.n548 0.708865
R429 VDD.n588 VDD.n547 0.708865
R430 VDD.n588 VDD.n546 0.708865
R431 VDD.n588 VDD.n545 0.708865
R432 VDD.n588 VDD.n544 0.708865
R433 VDD.n588 VDD.n543 0.708865
R434 VDD.n588 VDD.n542 0.708865
R435 VDD.n588 VDD.n541 0.708865
R436 VDD.n322 VDD.t12 0.311155
R437 VDD.n605 VDD.t23 0.311155
R438 VDD.n419 VDD.n418 0.122
R439 VDD.n19 VDD.n18 0.120875
R440 VDD.n268 VDD.n264 0.120875
R441 VDD.n214 VDD.n211 0.11075
R442 VDD.n207 VDD.n204 0.11075
R443 VDD.n204 VDD.n201 0.11075
R444 VDD.n201 VDD.n198 0.11075
R445 VDD.n198 VDD.n195 0.11075
R446 VDD.n195 VDD.n192 0.11075
R447 VDD.n188 VDD.n185 0.11075
R448 VDD.n185 VDD.n182 0.11075
R449 VDD.n182 VDD.n179 0.11075
R450 VDD.n175 VDD.n172 0.11075
R451 VDD.n172 VDD.n169 0.11075
R452 VDD.n169 VDD.n166 0.11075
R453 VDD.n166 VDD.n163 0.11075
R454 VDD.n163 VDD.n160 0.11075
R455 VDD.n156 VDD.n154 0.11075
R456 VDD.n154 VDD.n152 0.11075
R457 VDD.n149 VDD.n147 0.11075
R458 VDD.n147 VDD.n145 0.11075
R459 VDD.n145 VDD.n143 0.11075
R460 VDD.n143 VDD.n141 0.11075
R461 VDD.n141 VDD.n139 0.11075
R462 VDD.n136 VDD.n134 0.11075
R463 VDD.n134 VDD.n132 0.11075
R464 VDD.n18 VDD.n17 0.11075
R465 VDD.n17 VDD.n16 0.11075
R466 VDD.n16 VDD.n15 0.11075
R467 VDD.n15 VDD.n14 0.11075
R468 VDD.n14 VDD.n13 0.11075
R469 VDD.n13 VDD.n12 0.11075
R470 VDD.n12 VDD.n11 0.11075
R471 VDD.n11 VDD.n10 0.11075
R472 VDD.n10 VDD.n9 0.11075
R473 VDD.n9 VDD.n8 0.11075
R474 VDD.n8 VDD.n7 0.11075
R475 VDD.n7 VDD.n6 0.11075
R476 VDD.n6 VDD.n5 0.11075
R477 VDD.n5 VDD.n4 0.11075
R478 VDD.n4 VDD.n3 0.11075
R479 VDD.n3 VDD.n2 0.11075
R480 VDD.n2 VDD.n1 0.11075
R481 VDD.n1 VDD.n0 0.11075
R482 VDD.n400 VDD.n399 0.11075
R483 VDD.n401 VDD.n400 0.11075
R484 VDD.n402 VDD.n401 0.11075
R485 VDD.n403 VDD.n402 0.11075
R486 VDD.n404 VDD.n403 0.11075
R487 VDD.n405 VDD.n404 0.11075
R488 VDD.n406 VDD.n405 0.11075
R489 VDD.n407 VDD.n406 0.11075
R490 VDD.n408 VDD.n407 0.11075
R491 VDD.n409 VDD.n408 0.11075
R492 VDD.n410 VDD.n409 0.11075
R493 VDD.n411 VDD.n410 0.11075
R494 VDD.n412 VDD.n411 0.11075
R495 VDD.n413 VDD.n412 0.11075
R496 VDD.n414 VDD.n413 0.11075
R497 VDD.n415 VDD.n414 0.11075
R498 VDD.n416 VDD.n415 0.11075
R499 VDD.n417 VDD.n416 0.11075
R500 VDD.n68 VDD.n66 0.11075
R501 VDD.n66 VDD.n64 0.11075
R502 VDD.n61 VDD.n59 0.11075
R503 VDD.n59 VDD.n57 0.11075
R504 VDD.n57 VDD.n55 0.11075
R505 VDD.n55 VDD.n53 0.11075
R506 VDD.n53 VDD.n51 0.11075
R507 VDD.n48 VDD.n46 0.11075
R508 VDD.n46 VDD.n44 0.11075
R509 VDD.n41 VDD.n39 0.11075
R510 VDD.n39 VDD.n38 0.11075
R511 VDD.n38 VDD.n37 0.11075
R512 VDD.n37 VDD.n36 0.11075
R513 VDD.n36 VDD.n35 0.11075
R514 VDD.n33 VDD.n32 0.11075
R515 VDD.n32 VDD.n31 0.11075
R516 VDD.n31 VDD.n30 0.11075
R517 VDD.n28 VDD.n27 0.11075
R518 VDD.n27 VDD.n26 0.11075
R519 VDD.n26 VDD.n25 0.11075
R520 VDD.n25 VDD.n24 0.11075
R521 VDD.n24 VDD.n23 0.11075
R522 VDD.n21 VDD.n20 0.11075
R523 VDD.n465 VDD.n463 0.11075
R524 VDD.n463 VDD.n461 0.11075
R525 VDD.n458 VDD.n456 0.11075
R526 VDD.n456 VDD.n454 0.11075
R527 VDD.n454 VDD.n452 0.11075
R528 VDD.n452 VDD.n450 0.11075
R529 VDD.n450 VDD.n448 0.11075
R530 VDD.n445 VDD.n443 0.11075
R531 VDD.n443 VDD.n441 0.11075
R532 VDD.n439 VDD.n438 0.11075
R533 VDD.n438 VDD.n437 0.11075
R534 VDD.n437 VDD.n436 0.11075
R535 VDD.n436 VDD.n435 0.11075
R536 VDD.n435 VDD.n434 0.11075
R537 VDD.n432 VDD.n431 0.11075
R538 VDD.n431 VDD.n430 0.11075
R539 VDD.n430 VDD.n429 0.11075
R540 VDD.n427 VDD.n426 0.11075
R541 VDD.n426 VDD.n425 0.11075
R542 VDD.n425 VDD.n424 0.11075
R543 VDD.n424 VDD.n423 0.11075
R544 VDD.n423 VDD.n422 0.11075
R545 VDD.n420 VDD.n419 0.11075
R546 VDD.n540 VDD.n538 0.11075
R547 VDD.n534 VDD.n532 0.11075
R548 VDD.n532 VDD.n529 0.11075
R549 VDD.n529 VDD.n527 0.11075
R550 VDD.n527 VDD.n524 0.11075
R551 VDD.n524 VDD.n522 0.11075
R552 VDD.n518 VDD.n516 0.11075
R553 VDD.n516 VDD.n513 0.11075
R554 VDD.n513 VDD.n511 0.11075
R555 VDD.n508 VDD.n506 0.11075
R556 VDD.n506 VDD.n504 0.11075
R557 VDD.n504 VDD.n502 0.11075
R558 VDD.n502 VDD.n500 0.11075
R559 VDD.n500 VDD.n498 0.11075
R560 VDD.n495 VDD.n493 0.11075
R561 VDD.n493 VDD.n491 0.11075
R562 VDD.n488 VDD.n486 0.11075
R563 VDD.n486 VDD.n484 0.11075
R564 VDD.n484 VDD.n482 0.11075
R565 VDD.n482 VDD.n480 0.11075
R566 VDD.n480 VDD.n478 0.11075
R567 VDD.n475 VDD.n473 0.11075
R568 VDD.n473 VDD.n471 0.11075
R569 VDD.n471 VDD.n470 0.11075
R570 VDD.n272 VDD.n268 0.11075
R571 VDD.n276 VDD.n272 0.11075
R572 VDD.n280 VDD.n276 0.11075
R573 VDD.n284 VDD.n280 0.11075
R574 VDD.n288 VDD.n284 0.11075
R575 VDD.n292 VDD.n288 0.11075
R576 VDD.n296 VDD.n292 0.11075
R577 VDD.n300 VDD.n296 0.11075
R578 VDD.n304 VDD.n300 0.11075
R579 VDD.n308 VDD.n304 0.11075
R580 VDD.n312 VDD.n308 0.11075
R581 VDD.n316 VDD.n312 0.11075
R582 VDD.n320 VDD.n316 0.11075
R583 VDD.n324 VDD.n320 0.11075
R584 VDD.n328 VDD.n324 0.11075
R585 VDD.n332 VDD.n328 0.11075
R586 VDD.n336 VDD.n332 0.11075
R587 VDD.n340 VDD.n336 0.11075
R588 VDD.n667 VDD.n663 0.11075
R589 VDD.n663 VDD.n659 0.11075
R590 VDD.n659 VDD.n655 0.11075
R591 VDD.n655 VDD.n651 0.11075
R592 VDD.n651 VDD.n647 0.11075
R593 VDD.n647 VDD.n643 0.11075
R594 VDD.n643 VDD.n639 0.11075
R595 VDD.n639 VDD.n635 0.11075
R596 VDD.n635 VDD.n631 0.11075
R597 VDD.n631 VDD.n627 0.11075
R598 VDD.n627 VDD.n623 0.11075
R599 VDD.n623 VDD.n619 0.11075
R600 VDD.n619 VDD.n615 0.11075
R601 VDD.n615 VDD.n611 0.11075
R602 VDD.n611 VDD.n607 0.11075
R603 VDD.n607 VDD.n603 0.11075
R604 VDD.n603 VDD.n599 0.11075
R605 VDD.n599 VDD.n595 0.11075
R606 VDD.n595 VDD.n591 0.11075
R607 VDD.n211 VDD.n208 0.10175
R608 VDD.n22 VDD.n21 0.10175
R609 VDD.n421 VDD.n420 0.10175
R610 VDD.n538 VDD.n535 0.10175
R611 VDD.n192 VDD.n189 0.100625
R612 VDD.n29 VDD.n28 0.100625
R613 VDD.n441 VDD.n440 0.09275
R614 VDD.n496 VDD.n495 0.09275
R615 VDD.n428 VDD.n427 0.08825
R616 VDD.n522 VDD.n519 0.08825
R617 VDD.n157 VDD.n156 0.082625
R618 VDD.n44 VDD.n42 0.082625
R619 VDD.n176 VDD.n175 0.07925
R620 VDD.n35 VDD.n34 0.07925
R621 VDD.n264 VDD.n214 0.077
R622 VDD.n20 VDD.n19 0.077
R623 VDD.n468 VDD.n467 0.077
R624 VDD.n591 VDD.n540 0.077
R625 VDD.n446 VDD.n445 0.075875
R626 VDD.n491 VDD.n489 0.075875
R627 VDD.n434 VDD.n433 0.0725
R628 VDD.n509 VDD.n508 0.0725
R629 VDD.n139 VDD.n137 0.071375
R630 VDD.n62 VDD.n61 0.071375
R631 VDD.n459 VDD.n458 0.071375
R632 VDD.n478 VDD.n476 0.071375
R633 VDD.n152 VDD.n150 0.07025
R634 VDD.n49 VDD.n48 0.07025
R635 VDD.n130 VDD.n128 0.068
R636 VDD.n128 VDD.n70 0.068
R637 VDD.n132 VDD.n130 0.06575
R638 VDD.n418 VDD.n417 0.06575
R639 VDD.n70 VDD.n68 0.06575
R640 VDD.n467 VDD.n465 0.06575
R641 VDD VDD.n340 0.062375
R642 VDD VDD.n667 0.048875
R643 VDD.n150 VDD.n149 0.041
R644 VDD.n51 VDD.n49 0.041
R645 VDD.n137 VDD.n136 0.039875
R646 VDD.n64 VDD.n62 0.039875
R647 VDD.n461 VDD.n459 0.039875
R648 VDD.n476 VDD.n475 0.039875
R649 VDD.n433 VDD.n432 0.03875
R650 VDD.n511 VDD.n509 0.03875
R651 VDD.n127 VDD.n124 0.0369463
R652 VDD.n124 VDD.n121 0.0369463
R653 VDD.n121 VDD.n118 0.0369463
R654 VDD.n118 VDD.n115 0.0369463
R655 VDD.n115 VDD.n112 0.0369463
R656 VDD.n112 VDD.n109 0.0369463
R657 VDD.n109 VDD.n106 0.0369463
R658 VDD.n106 VDD.n103 0.0369463
R659 VDD.n103 VDD.n100 0.0369463
R660 VDD.n100 VDD.n97 0.0369463
R661 VDD.n97 VDD.n94 0.0369463
R662 VDD.n94 VDD.n91 0.0369463
R663 VDD.n91 VDD.n88 0.0369463
R664 VDD.n88 VDD.n85 0.0369463
R665 VDD.n85 VDD.n82 0.0369463
R666 VDD.n82 VDD.n79 0.0369463
R667 VDD.n79 VDD.n76 0.0369463
R668 VDD.n76 VDD.n73 0.0369463
R669 VDD.n347 VDD.n344 0.0369463
R670 VDD.n350 VDD.n347 0.0369463
R671 VDD.n353 VDD.n350 0.0369463
R672 VDD.n356 VDD.n353 0.0369463
R673 VDD.n359 VDD.n356 0.0369463
R674 VDD.n362 VDD.n359 0.0369463
R675 VDD.n365 VDD.n362 0.0369463
R676 VDD.n368 VDD.n365 0.0369463
R677 VDD.n371 VDD.n368 0.0369463
R678 VDD.n374 VDD.n371 0.0369463
R679 VDD.n377 VDD.n374 0.0369463
R680 VDD.n380 VDD.n377 0.0369463
R681 VDD.n383 VDD.n380 0.0369463
R682 VDD.n386 VDD.n383 0.0369463
R683 VDD.n389 VDD.n386 0.0369463
R684 VDD.n392 VDD.n389 0.0369463
R685 VDD.n395 VDD.n392 0.0369463
R686 VDD.n398 VDD.n395 0.0369463
R687 VDD.n448 VDD.n446 0.035375
R688 VDD.n489 VDD.n488 0.035375
R689 VDD.n179 VDD.n176 0.032
R690 VDD.n34 VDD.n33 0.032
R691 VDD.n470 VDD.n468 0.032
R692 VDD.n160 VDD.n157 0.028625
R693 VDD.n42 VDD.n41 0.028625
R694 VDD.n429 VDD.n428 0.023
R695 VDD.n519 VDD.n518 0.023
R696 VDD.n440 VDD.n439 0.0185
R697 VDD.n498 VDD.n496 0.0185
R698 VDD.n128 VDD.n127 0.0179793
R699 VDD.n468 VDD.n398 0.011657
R700 VDD.n189 VDD.n188 0.010625
R701 VDD.n30 VDD.n29 0.010625
R702 VDD.n208 VDD.n207 0.0095
R703 VDD.n23 VDD.n22 0.0095
R704 VDD.n422 VDD.n421 0.0095
R705 VDD.n535 VDD.n534 0.0095
R706 VOUT_OPAMP_N.n0 VOUT_OPAMP_N.t6 6.52638
R707 VOUT_OPAMP_N.n2 VOUT_OPAMP_N.t2 6.43144
R708 VOUT_OPAMP_N.n1 VOUT_OPAMP_N.t0 6.43144
R709 VOUT_OPAMP_N.n0 VOUT_OPAMP_N.t1 6.43144
R710 VOUT_OPAMP_N.n3 VOUT_OPAMP_N.t3 3.18932
R711 VOUT_OPAMP_N.n6 VOUT_OPAMP_N.t5 2.73371
R712 VOUT_OPAMP_N.n6 VOUT_OPAMP_N.t4 2.4088
R713 VOUT_OPAMP_N VOUT_OPAMP_N.n10 1.65759
R714 VOUT_OPAMP_N VOUT_OPAMP_N.n3 1.65341
R715 VOUT_OPAMP_N.n5 VOUT_OPAMP_N.n4 1.4964
R716 VOUT_OPAMP_N.n8 VOUT_OPAMP_N.n7 1.49069
R717 VOUT_OPAMP_N.n10 VOUT_OPAMP_N.n9 1.14993
R718 VOUT_OPAMP_N.n10 VOUT_OPAMP_N.n5 1.14978
R719 VOUT_OPAMP_N.n3 VOUT_OPAMP_N.n2 0.302215
R720 VOUT_OPAMP_N.n1 VOUT_OPAMP_N.n0 0.289625
R721 VOUT_OPAMP_N.n2 VOUT_OPAMP_N.n1 0.069461
R722 VOUT_OPAMP_N.n7 VOUT_OPAMP_N.n6 0.0608233
R723 VOUT_OPAMP_N.n9 VOUT_OPAMP_N.n8 0.0164591
R724 VOUT_N VOUT_N.t0 4.20169
R725 VOUT_N VOUT_N.n0 3.47982
R726 VOUT_N.n0 VOUT_N.t1 2.38651
R727 VOUT_N.n0 VOUT_N.t2 2.2505
R728 VOUT_OPAMP_P.n17 VOUT_OPAMP_P.t4 6.55774
R729 VOUT_OPAMP_P.n19 VOUT_OPAMP_P.t1 6.43045
R730 VOUT_OPAMP_P.n18 VOUT_OPAMP_P.t3 6.42009
R731 VOUT_OPAMP_P.n17 VOUT_OPAMP_P.t2 6.4095
R732 VOUT_OPAMP_P.n12 VOUT_OPAMP_P.n11 2.82778
R733 VOUT_OPAMP_P.n2 VOUT_OPAMP_P.t5 2.73276
R734 VOUT_OPAMP_P.n2 VOUT_OPAMP_P.t6 2.40975
R735 VOUT_OPAMP_P.n21 VOUT_OPAMP_P.n20 2.2505
R736 VOUT_OPAMP_P.n11 VOUT_OPAMP_P.t0 2.1905
R737 VOUT_OPAMP_P VOUT_OPAMP_P.n6 1.67937
R738 VOUT_OPAMP_P.n1 VOUT_OPAMP_P.n0 1.4964
R739 VOUT_OPAMP_P.n4 VOUT_OPAMP_P.n3 1.49069
R740 VOUT_OPAMP_P.n6 VOUT_OPAMP_P.n5 1.14993
R741 VOUT_OPAMP_P.n6 VOUT_OPAMP_P.n1 1.14978
R742 VOUT_OPAMP_P VOUT_OPAMP_P.n21 0.878717
R743 VOUT_OPAMP_P.n20 VOUT_OPAMP_P.n19 0.245262
R744 VOUT_OPAMP_P.n18 VOUT_OPAMP_P.n17 0.212047
R745 VOUT_OPAMP_P.n12 VOUT_OPAMP_P.n10 0.141929
R746 VOUT_OPAMP_P.n14 VOUT_OPAMP_P.n13 0.121357
R747 VOUT_OPAMP_P.n19 VOUT_OPAMP_P.n18 0.0830882
R748 VOUT_OPAMP_P.n3 VOUT_OPAMP_P.n2 0.0608233
R749 VOUT_OPAMP_P.n10 VOUT_OPAMP_P.n9 0.051948
R750 VOUT_OPAMP_P.n14 VOUT_OPAMP_P.n12 0.0210714
R751 VOUT_OPAMP_P.n5 VOUT_OPAMP_P.n4 0.0164591
R752 VOUT_OPAMP_P.n21 VOUT_OPAMP_P.n8 0.0108185
R753 VOUT_OPAMP_P.n16 VOUT_OPAMP_P.n15 0.00764286
R754 VOUT_OPAMP_P.n8 VOUT_OPAMP_P.n7 0.00623248
R755 VOUT_OPAMP_P.n15 VOUT_OPAMP_P.n14 0.00240476
R756 VOUT_OPAMP_P.n20 VOUT_OPAMP_P.n16 0.00192857
R757 a_387_n202.t3 a_387_n202.t2 5.9203
R758 a_387_n202.t3 a_387_n202.t1 4.57473
R759 a_387_n202.t0 a_387_n202.t3 3.89251
R760 R3_R7.n3 R3_R7.t4 5.14152
R761 R3_R7.n0 R3_R7.t0 4.72867
R762 R3_R7.n0 R3_R7.t1 3.99183
R763 R3_R7.n5 R3_R7.n4 2.88446
R764 R3_R7.n7 R3_R7.t6 2.27001
R765 R3_R7.n6 R3_R7.t5 2.25756
R766 R3_R7.n5 R3_R7.t7 2.25756
R767 R3_R7.n6 R3_R7.n5 1.44088
R768 R3_R7.n12 R3_R7.n1 1.14829
R769 R3_R7.n11 R3_R7.n10 1.1255
R770 R3_R7.n13 R3_R7.n12 0.608075
R771 R3_R7.n7 R3_R7.n6 0.582009
R772 R3_R7.n9 R3_R7.n8 0.577293
R773 R3_R7.n4 R3_R7.n3 0.352858
R774 R3_R7 R3_R7.n0 0.299466
R775 R3_R7 R3_R7.n13 0.152486
R776 R3_R7.n8 R3_R7.n7 0.0937076
R777 R3_R7.n11 R3_R7.n2 0.0450755
R778 R3_R7.n10 R3_R7.n9 0.0226677
R779 R3_R7.n12 R3_R7.n11 0.0224383
R780 R3_R7.n3 R3_R7.t3 0.00755556
R781 R3_R7.n4 R3_R7.t2 0.00755556
R782 a_667_n202.t0 a_667_n202.t1 13.5425
R783 a_387_n1119.n2 a_387_n1119.t1 7.26507
R784 a_387_n1119.n0 a_387_n1119.t0 3.89298
R785 a_387_n1119.t3 a_387_n1119.t4 3.06722
R786 a_387_n1119.n5 a_387_n1119.t2 2.3
R787 a_387_n1119.t4 a_387_n1119.n1 1.76691
R788 a_387_n1119.n3 a_387_n1119.n5 1.72527
R789 a_387_n1119.t4 a_387_n1119.n7 1.1255
R790 a_387_n1119.n1 a_387_n1119.n0 0.657163
R791 a_387_n1119.n4 a_387_n1119.n2 0.0210063
R792 a_387_n1119.n4 a_387_n1119.n3 0.0118924
R793 a_387_n1119.n4 a_387_n1119.n0 2.47036
R794 a_387_n1119.t4 a_387_n1119.n6 1.73255
R795 a_387_n3450.t0 a_387_n3450.t1 14.32
R796 a_667_153.t0 a_667_153.t1 13.5425
R797 a_667_n1119.t0 a_667_n1119.t1 12.9821
R798 a_387_n1681.t0 a_387_n1681.t1 12.9821
R799 R7_R8_R10_C.n3 R7_R8_R10_C.t2 7.26507
R800 R7_R8_R10_C.n11 R7_R8_R10_C.t1 3.97272
R801 R7_R8_R10_C.n14 R7_R8_R10_C.t3 2.3855
R802 R7_R8_R10_C.n0 R7_R8_R10_C.t0 2.3
R803 R7_R8_R10_C.n14 R7_R8_R10_C.t4 2.2505
R804 R7_R8_R10_C.n9 R7_R8_R10_C.n6 2.2501
R805 R7_R8_R10_C R7_R8_R10_C.n24 2.06348
R806 R7_R8_R10_C.n1 R7_R8_R10_C.n0 1.72411
R807 R7_R8_R10_C.n22 R7_R8_R10_C.n12 1.148
R808 R7_R8_R10_C.n19 R7_R8_R10_C.n18 1.1255
R809 R7_R8_R10_C.n21 R7_R8_R10_C.n20 1.1255
R810 R7_R8_R10_C.n23 R7_R8_R10_C.n22 0.6075
R811 R7_R8_R10_C.n17 R7_R8_R10_C.n16 0.577112
R812 R7_R8_R10_C R7_R8_R10_C.n11 0.299909
R813 R7_R8_R10_C.n11 R7_R8_R10_C.n10 0.155122
R814 R7_R8_R10_C.n15 R7_R8_R10_C.n14 0.0793189
R815 R7_R8_R10_C.n19 R7_R8_R10_C.n13 0.0445
R816 R7_R8_R10_C.n21 R7_R8_R10_C.n19 0.0445
R817 R7_R8_R10_C.n24 R7_R8_R10_C.n23 0.0445
R818 R7_R8_R10_C.n5 R7_R8_R10_C.n4 0.0335186
R819 R7_R8_R10_C.n18 R7_R8_R10_C.n17 0.0223956
R820 R7_R8_R10_C.n22 R7_R8_R10_C.n21 0.0221719
R821 R7_R8_R10_C.n4 R7_R8_R10_C.n3 0.0198671
R822 R7_R8_R10_C.n6 R7_R8_R10_C.n5 0.0126852
R823 R7_R8_R10_C.n2 R7_R8_R10_C.n1 0.00961392
R824 R7_R8_R10_C.n8 R7_R8_R10_C.n7 0.0095
R825 R7_R8_R10_C.n16 R7_R8_R10_C.n15 0.00903333
R826 R7_R8_R10_C.n4 R7_R8_R10_C.n2 0.00391772
R827 R7_R8_R10_C.n9 R7_R8_R10_C.n8 0.00279928
R828 R7_R8_R10_C.n10 R7_R8_R10_C.n9 0.00279928
R829 VIN_N VIN_N.t0 5.04285
R830 a_1507_n4012.t0 a_1507_n4012.t1 14.4367
R831 a_387_n4367.t0 a_387_n4367.t1 13.5444
R832 a_947_n4929.t0 a_947_n4929.t1 13.5425
R833 a_387_n2533.t0 a_387_n2533.t1 12.9821
R834 a_667_n3095.t0 a_667_n3095.t1 12.9821
R835 a_667_n4367.t0 a_667_n4367.t1 13.5425
R836 a_1227_n4929.t0 a_1227_n4929.t1 13.5444
R837 a_387_n764.t0 a_387_n764.t1 14.32
R838 a_1787_n4367.t0 a_1787_n4367.t1 13.5425
R839 VOUT_P VOUT_P.t0 4.25927
R840 VOUT_P VOUT_P.n0 3.4605
R841 VOUT_P.n0 VOUT_P.t1 2.38651
R842 VOUT_P.n0 VOUT_P.t2 2.2505
R843 a_667_n4012.t0 a_667_n4012.t1 13.5425
R844 a_947_n1681.t0 a_947_n1681.t1 12.9821
R845 a_1227_n1119.t0 a_1227_n1119.t1 12.98
R846 a_2347_n3450.t0 a_2347_n3450.t1 13.5425
R847 a_2627_n4367.t0 a_2627_n4367.t1 10.1673
R848 a_2347_715.t0 a_2347_715.t1 13.5444
R849 a_1787_153.t0 a_1787_153.t1 13.5425
R850 a_1507_n4367.t0 a_1507_n4367.t1 13.5425
R851 a_2067_n4929.t0 a_2067_n4929.t1 13.5425
R852 a_1227_715.t0 a_1227_715.t1 13.5444
R853 a_947_n2533.t0 a_947_n2533.t1 12.9821
R854 a_1787_n1119.t0 a_1787_n1119.t1 12.9667
R855 a_1507_n1681.t0 a_1507_n1681.t1 13.0109
R856 a_1227_n3095.t0 a_1227_n3095.t1 12.9821
R857 a_387_153.t0 a_387_153.t1 13.5444
R858 a_947_n3450.t0 a_947_n3450.t1 14.6442
R859 a_2067_n1681.t0 a_2067_n1681.t1 12.9667
R860 a_1507_n2533.t0 a_1507_n2533.t1 12.9821
R861 a_1787_n3095.t0 a_1787_n3095.t1 12.9821
R862 a_1227_n3450.t0 a_1227_n3450.t1 13.5425
R863 a_2347_n4929.t0 a_2347_n4929.t1 13.5444
R864 a_2067_n202.t0 a_2067_n202.t1 8.88555
R865 a_2627_153.t0 a_2627_153.t1 10.1324
R866 a_2347_n764.t0 a_2347_n764.t1 13.5425
R867 a_2067_n2533.t0 a_2067_n2533.t1 12.9821
R868 a_1787_n4012.t0 a_1787_n4012.t1 13.5425
R869 a_1507_n202.t0 a_1507_n202.t1 14.4367
R870 a_2067_n4012.t0 a_2067_n4012.t1 8.92045
R871 a_2067_715.t0 a_2067_715.t1 13.5425
R872 VIN_P VIN_P.t0 5.25526
R873 a_1227_n764.t0 a_1227_n764.t1 13.5425
R874 a_1787_n202.t0 a_1787_n202.t1 13.5425
R875 a_947_n764.t0 a_947_n764.t1 14.6442
C0 R3_R7 VOUT_P 0.551f
C1 VDD VIN_P 0.641f
C2 VOUT_OPAMP_N VOUT_P 3.76f
C3 VDD R3_R7 0.943f
C4 VOUT_N R7_R8_R10_C 0.00657f
C5 VDD VOUT_OPAMP_N 2.04f
C6 VOUT_N VOUT_OPAMP_P 3.76f
C7 VDD VOUT_P 0.457f
C8 VIN_P R7_R8_R10_C 0.00311f
C9 VIN_P VOUT_OPAMP_P 0.0407f
C10 R7_R8_R10_C R3_R7 1.53f
C11 R7_R8_R10_C VOUT_OPAMP_N 6.07e-19
C12 VOUT_OPAMP_P VOUT_OPAMP_N 0.0476f
C13 R3_R7 VIN_N 0.234f
C14 VOUT_OPAMP_N VIN_N 0.0413f
C15 VDD R7_R8_R10_C 1.03f
C16 m3_n2949_2707# R7_R8_R10_C 0.0764f
C17 VDD VOUT_OPAMP_P 2.04f
C18 VDD VIN_N 0.648f
C19 VDD VOUT_N 0.457f
C20 R7_R8_R10_C VIN_N 0.407f
C21 VOUT_OPAMP_N R3_R7 0.351f
C22 VOUT_P VSUBS 7.38f
C23 VIN_N VSUBS 0.364f
C24 R3_R7 VSUBS 11.4f
C25 VOUT_OPAMP_N VSUBS 6.25f
C26 R7_R8_R10_C VSUBS 7.3f
C27 VOUT_OPAMP_P VSUBS 6.15f
C28 VIN_P VSUBS 0.376f
C29 VOUT_N VSUBS 7.38f
C30 VDD VSUBS 81.4f
C31 m3_n2949_2707# VSUBS 0.0548f $ **FLOATING
C32 VOUT_P.t0 VSUBS 0.00201f
C33 VOUT_P.t1 VSUBS 1.03f
C34 VOUT_P.t2 VSUBS 0.976f
C35 VOUT_P.n0 VSUBS 1.74f
C36 R7_R8_R10_C.t1 VSUBS 0.0015f
C37 R7_R8_R10_C.t0 VSUBS 6.22e-19
C38 R7_R8_R10_C.n0 VSUBS 0.00133f
C39 R7_R8_R10_C.n1 VSUBS 2.94e-19
C40 R7_R8_R10_C.n2 VSUBS 4.28e-20
C41 R7_R8_R10_C.t2 VSUBS 0.00191f
C42 R7_R8_R10_C.n3 VSUBS 0.00629f
C43 R7_R8_R10_C.n4 VSUBS 4.95e-19
C44 R7_R8_R10_C.n6 VSUBS 4.53e-19
C45 R7_R8_R10_C.n7 VSUBS 5.72e-19
C46 R7_R8_R10_C.n8 VSUBS 2.76e-19
C47 R7_R8_R10_C.n10 VSUBS 0.00424f
C48 R7_R8_R10_C.n11 VSUBS 0.0135f
C49 R7_R8_R10_C.n12 VSUBS 0.00228f
C50 R7_R8_R10_C.n13 VSUBS 0.00215f
C51 R7_R8_R10_C.t3 VSUBS 1.01f
C52 R7_R8_R10_C.t4 VSUBS 0.959f
C53 R7_R8_R10_C.n14 VSUBS 1.64f
C54 R7_R8_R10_C.n15 VSUBS 0.0575f
C55 R7_R8_R10_C.n16 VSUBS 0.00612f
C56 R7_R8_R10_C.n17 VSUBS 0.00226f
C57 R7_R8_R10_C.n18 VSUBS 0.00244f
C58 R7_R8_R10_C.n19 VSUBS 0.00244f
C59 R7_R8_R10_C.n20 VSUBS 0.00244f
C60 R7_R8_R10_C.n21 VSUBS 0.00244f
C61 R7_R8_R10_C.n22 VSUBS 0.00259f
C62 R7_R8_R10_C.n23 VSUBS 0.00669f
C63 R7_R8_R10_C.n24 VSUBS 0.0361f
C64 a_387_n1119.t4 VSUBS 2.01f
C65 a_387_n1119.t0 VSUBS 0.00839f
C66 a_387_n1119.n0 VSUBS 0.125f
C67 a_387_n1119.n1 VSUBS 0.127f
C68 a_387_n1119.t1 VSUBS 0.0109f
C69 a_387_n1119.n2 VSUBS 0.0359f
C70 a_387_n1119.n3 VSUBS 0.00168f
C71 a_387_n1119.n4 VSUBS 0.00678f
C72 a_387_n1119.t2 VSUBS 0.00355f
C73 a_387_n1119.n5 VSUBS 0.0076f
C74 a_387_n1119.n6 VSUBS 0.0116f
C75 a_387_n1119.n7 VSUBS 0.013f
C76 a_387_n1119.t3 VSUBS 1.43f
C77 R3_R7.t1 VSUBS 0.0109f
C78 R3_R7.t0 VSUBS 0.0204f
C79 R3_R7.n0 VSUBS 0.154f
C80 R3_R7.n1 VSUBS 0.0143f
C81 R3_R7.n2 VSUBS 0.0149f
C82 R3_R7.t6 VSUBS 1.65f
C83 R3_R7.t5 VSUBS 1.65f
C84 R3_R7.t4 VSUBS 2.15f
C85 R3_R7.t3 VSUBS 1.12f
C86 R3_R7.n3 VSUBS 1.1f
C87 R3_R7.t2 VSUBS 1.12f
C88 R3_R7.n4 VSUBS 0.707f
C89 R3_R7.t7 VSUBS 1.65f
C90 R3_R7.n5 VSUBS 1.24f
C91 R3_R7.n6 VSUBS 0.821f
C92 R3_R7.n7 VSUBS 0.546f
C93 R3_R7.n8 VSUBS 0.074f
C94 R3_R7.n9 VSUBS 0.0156f
C95 R3_R7.n10 VSUBS 0.0158f
C96 R3_R7.n11 VSUBS 0.0158f
C97 R3_R7.n12 VSUBS 0.0157f
C98 R3_R7.n13 VSUBS 0.0485f
C99 a_387_n202.t2 VSUBS 3.53f
C100 a_387_n202.t3 VSUBS 10.7f
C101 a_387_n202.t1 VSUBS 0.00327f
C102 a_387_n202.t0 VSUBS 0.00186f
C103 VOUT_OPAMP_P.n0 VSUBS 0.0178f
C104 VOUT_OPAMP_P.n1 VSUBS 0.0184f
C105 VOUT_OPAMP_P.t6 VSUBS 1.88f
C106 VOUT_OPAMP_P.t5 VSUBS 1.95f
C107 VOUT_OPAMP_P.n2 VSUBS 1.05f
C108 VOUT_OPAMP_P.n3 VSUBS 0.0276f
C109 VOUT_OPAMP_P.n5 VSUBS 0.0181f
C110 VOUT_OPAMP_P.n6 VSUBS 0.136f
C111 VOUT_OPAMP_P.n7 VSUBS 0.00374f
C112 VOUT_OPAMP_P.n8 VSUBS -2.49e-19
C113 VOUT_OPAMP_P.n9 VSUBS 3.66e-19
C114 VOUT_OPAMP_P.n10 VSUBS 0.0015f
C115 VOUT_OPAMP_P.t0 VSUBS 0.00476f
C116 VOUT_OPAMP_P.n11 VSUBS 0.0108f
C117 VOUT_OPAMP_P.n12 VSUBS 0.00149f
C118 VOUT_OPAMP_P.n13 VSUBS 0.00189f
C119 VOUT_OPAMP_P.n14 VSUBS 0.00106f
C120 VOUT_OPAMP_P.n15 VSUBS 0.00142f
C121 VOUT_OPAMP_P.n16 VSUBS 0.00195f
C122 VOUT_OPAMP_P.t2 VSUBS 0.0121f
C123 VOUT_OPAMP_P.t4 VSUBS 0.0129f
C124 VOUT_OPAMP_P.n17 VSUBS 0.0894f
C125 VOUT_OPAMP_P.t3 VSUBS 0.0121f
C126 VOUT_OPAMP_P.n18 VSUBS 0.0511f
C127 VOUT_OPAMP_P.t1 VSUBS 0.0121f
C128 VOUT_OPAMP_P.n19 VSUBS 0.0636f
C129 VOUT_OPAMP_P.n20 VSUBS 0.0388f
C130 VOUT_OPAMP_P.n21 VSUBS 0.108f
C131 VOUT_N.t1 VSUBS 1.03f
C132 VOUT_N.t2 VSUBS 0.976f
C133 VOUT_N.n0 VSUBS 1.74f
C134 VOUT_N.t0 VSUBS 0.00196f
C135 VOUT_OPAMP_N.t0 VSUBS 0.0122f
C136 VOUT_OPAMP_N.t6 VSUBS 0.0126f
C137 VOUT_OPAMP_N.t1 VSUBS 0.0122f
C138 VOUT_OPAMP_N.n0 VSUBS 0.0845f
C139 VOUT_OPAMP_N.n1 VSUBS 0.0515f
C140 VOUT_OPAMP_N.t2 VSUBS 0.0122f
C141 VOUT_OPAMP_N.n2 VSUBS 0.0523f
C142 VOUT_OPAMP_N.t3 VSUBS 0.00815f
C143 VOUT_OPAMP_N.n3 VSUBS 0.112f
C144 VOUT_OPAMP_N.n4 VSUBS 0.0178f
C145 VOUT_OPAMP_N.n5 VSUBS 0.0181f
C146 VOUT_OPAMP_N.t4 VSUBS 1.89f
C147 VOUT_OPAMP_N.t5 VSUBS 1.96f
C148 VOUT_OPAMP_N.n6 VSUBS 1.05f
C149 VOUT_OPAMP_N.n7 VSUBS 0.0277f
C150 VOUT_OPAMP_N.n9 VSUBS 0.0185f
C151 VOUT_OPAMP_N.n10 VSUBS 0.135f
C152 VDD.t13 VSUBS 0.00209f
C153 VDD.t14 VSUBS 0.00209f
C154 VDD.t21 VSUBS 0.00209f
C155 VDD.t22 VSUBS 0.00209f
C156 VDD.t10 VSUBS 0.00209f
C157 VDD.t11 VSUBS 0.00209f
C158 VDD.t19 VSUBS 0.00209f
C159 VDD.t20 VSUBS 0.00209f
C160 VDD.t15 VSUBS 0.00209f
C161 VDD.t16 VSUBS 0.00209f
C162 VDD.t3 VSUBS 0.00209f
C163 VDD.t4 VSUBS 0.00209f
C164 VDD.n0 VSUBS 9.88e-19
C165 VDD.n1 VSUBS 9.88e-19
C166 VDD.n2 VSUBS 9.88e-19
C167 VDD.n3 VSUBS 9.88e-19
C168 VDD.n4 VSUBS 9.88e-19
C169 VDD.n5 VSUBS 9.88e-19
C170 VDD.n6 VSUBS 9.88e-19
C171 VDD.n7 VSUBS 9.88e-19
C172 VDD.n8 VSUBS 9.88e-19
C173 VDD.n9 VSUBS 9.88e-19
C174 VDD.n10 VSUBS 9.88e-19
C175 VDD.n11 VSUBS 9.88e-19
C176 VDD.n12 VSUBS 9.88e-19
C177 VDD.n13 VSUBS 9.88e-19
C178 VDD.n14 VSUBS 9.88e-19
C179 VDD.n15 VSUBS 9.88e-19
C180 VDD.n16 VSUBS 9.88e-19
C181 VDD.n17 VSUBS 9.88e-19
C182 VDD.n18 VSUBS 0.00103f
C183 VDD.n19 VSUBS 0.00129f
C184 VDD.n20 VSUBS 8.37e-19
C185 VDD.n21 VSUBS 9.48e-19
C186 VDD.n22 VSUBS 0.00452f
C187 VDD.n23 VSUBS 5.35e-19
C188 VDD.n24 VSUBS 9.88e-19
C189 VDD.n25 VSUBS 9.88e-19
C190 VDD.n26 VSUBS 9.88e-19
C191 VDD.n27 VSUBS 9.88e-19
C192 VDD.n28 VSUBS 9.43e-19
C193 VDD.n29 VSUBS 0.00455f
C194 VDD.n30 VSUBS 5.4e-19
C195 VDD.n31 VSUBS 9.88e-19
C196 VDD.n32 VSUBS 9.88e-19
C197 VDD.n33 VSUBS 6.35e-19
C198 VDD.n34 VSUBS 0.00454f
C199 VDD.n35 VSUBS 8.47e-19
C200 VDD.n36 VSUBS 9.88e-19
C201 VDD.n37 VSUBS 9.88e-19
C202 VDD.n38 VSUBS 9.88e-19
C203 VDD.n39 VSUBS 9.88e-19
C204 VDD.n40 VSUBS 9.88e-19
C205 VDD.n41 VSUBS 6.2e-19
C206 VDD.n42 VSUBS 0.00455f
C207 VDD.n43 VSUBS 9.88e-19
C208 VDD.n44 VSUBS 8.62e-19
C209 VDD.n45 VSUBS 9.88e-19
C210 VDD.n46 VSUBS 9.88e-19
C211 VDD.n47 VSUBS 9.88e-19
C212 VDD.n48 VSUBS 8.07e-19
C213 VDD.n49 VSUBS 0.00455f
C214 VDD.n50 VSUBS 9.88e-19
C215 VDD.n51 VSUBS 6.76e-19
C216 VDD.n52 VSUBS 9.88e-19
C217 VDD.n53 VSUBS 9.88e-19
C218 VDD.n54 VSUBS 9.88e-19
C219 VDD.n55 VSUBS 9.88e-19
C220 VDD.n56 VSUBS 9.88e-19
C221 VDD.n57 VSUBS 9.88e-19
C222 VDD.n58 VSUBS 9.88e-19
C223 VDD.n59 VSUBS 9.88e-19
C224 VDD.n60 VSUBS 9.88e-19
C225 VDD.n61 VSUBS 8.12e-19
C226 VDD.n62 VSUBS 0.00455f
C227 VDD.n63 VSUBS 9.88e-19
C228 VDD.n64 VSUBS 6.71e-19
C229 VDD.n65 VSUBS 9.88e-19
C230 VDD.n66 VSUBS 9.88e-19
C231 VDD.n67 VSUBS 7.87e-19
C232 VDD.n68 VSUBS 7.87e-19
C233 VDD.n69 VSUBS 0.00124f
C234 VDD.n70 VSUBS 9.98e-19
C235 VDD.n71 VSUBS 9.88e-19
C236 VDD.n72 VSUBS 9.88e-19
C237 VDD.n73 VSUBS 0.00299f
C238 VDD.n74 VSUBS 9.88e-19
C239 VDD.n75 VSUBS 9.88e-19
C240 VDD.n76 VSUBS 0.00299f
C241 VDD.n77 VSUBS 9.88e-19
C242 VDD.n78 VSUBS 9.88e-19
C243 VDD.n79 VSUBS 0.00299f
C244 VDD.n80 VSUBS 9.88e-19
C245 VDD.n81 VSUBS 9.88e-19
C246 VDD.n82 VSUBS 0.00299f
C247 VDD.n83 VSUBS 9.88e-19
C248 VDD.n84 VSUBS 9.88e-19
C249 VDD.n85 VSUBS 0.00299f
C250 VDD.n86 VSUBS 9.88e-19
C251 VDD.n87 VSUBS 9.88e-19
C252 VDD.n88 VSUBS 0.00299f
C253 VDD.n89 VSUBS 9.88e-19
C254 VDD.n90 VSUBS 9.88e-19
C255 VDD.n91 VSUBS 0.00299f
C256 VDD.n92 VSUBS 9.88e-19
C257 VDD.n93 VSUBS 9.88e-19
C258 VDD.n94 VSUBS 0.00299f
C259 VDD.n95 VSUBS 9.88e-19
C260 VDD.n96 VSUBS 9.88e-19
C261 VDD.n97 VSUBS 0.00299f
C262 VDD.n98 VSUBS 9.88e-19
C263 VDD.n99 VSUBS 9.88e-19
C264 VDD.n100 VSUBS 0.00299f
C265 VDD.n101 VSUBS 9.88e-19
C266 VDD.n102 VSUBS 9.88e-19
C267 VDD.n103 VSUBS 0.00299f
C268 VDD.n104 VSUBS 9.88e-19
C269 VDD.n105 VSUBS 9.88e-19
C270 VDD.n106 VSUBS 0.00299f
C271 VDD.n107 VSUBS 9.88e-19
C272 VDD.n108 VSUBS 9.88e-19
C273 VDD.n109 VSUBS 0.00299f
C274 VDD.n110 VSUBS 9.88e-19
C275 VDD.n111 VSUBS 9.88e-19
C276 VDD.n112 VSUBS 0.00299f
C277 VDD.n113 VSUBS 9.88e-19
C278 VDD.n114 VSUBS 9.88e-19
C279 VDD.n115 VSUBS 0.00299f
C280 VDD.n116 VSUBS 9.88e-19
C281 VDD.n117 VSUBS 9.88e-19
C282 VDD.n118 VSUBS 0.00299f
C283 VDD.n119 VSUBS 9.88e-19
C284 VDD.n120 VSUBS 9.88e-19
C285 VDD.n121 VSUBS 0.00299f
C286 VDD.n122 VSUBS 9.88e-19
C287 VDD.n123 VSUBS 9.88e-19
C288 VDD.n124 VSUBS 0.00299f
C289 VDD.n125 VSUBS 0.00103f
C290 VDD.n126 VSUBS 0.00103f
C291 VDD.n127 VSUBS 0.00221f
C292 VDD.n128 VSUBS 0.00132f
C293 VDD.n129 VSUBS 0.00124f
C294 VDD.n130 VSUBS 9.98e-19
C295 VDD.n131 VSUBS 7.87e-19
C296 VDD.n132 VSUBS 7.87e-19
C297 VDD.n133 VSUBS 9.88e-19
C298 VDD.n134 VSUBS 9.88e-19
C299 VDD.n135 VSUBS 9.88e-19
C300 VDD.n136 VSUBS 6.71e-19
C301 VDD.n137 VSUBS 0.00455f
C302 VDD.n138 VSUBS 9.88e-19
C303 VDD.n139 VSUBS 8.12e-19
C304 VDD.n140 VSUBS 9.88e-19
C305 VDD.n141 VSUBS 9.88e-19
C306 VDD.n142 VSUBS 9.88e-19
C307 VDD.n143 VSUBS 9.88e-19
C308 VDD.n144 VSUBS 9.88e-19
C309 VDD.n145 VSUBS 9.88e-19
C310 VDD.n146 VSUBS 9.88e-19
C311 VDD.n147 VSUBS 9.88e-19
C312 VDD.n148 VSUBS 9.88e-19
C313 VDD.n149 VSUBS 6.76e-19
C314 VDD.n150 VSUBS 0.00455f
C315 VDD.n151 VSUBS 9.88e-19
C316 VDD.n152 VSUBS 8.07e-19
C317 VDD.n153 VSUBS 9.88e-19
C318 VDD.n154 VSUBS 9.88e-19
C319 VDD.n155 VSUBS 9.88e-19
C320 VDD.n156 VSUBS 8.62e-19
C321 VDD.n157 VSUBS 0.00455f
C322 VDD.n159 VSUBS 9.88e-19
C323 VDD.n160 VSUBS 6.2e-19
C324 VDD.n162 VSUBS 9.88e-19
C325 VDD.n163 VSUBS 9.88e-19
C326 VDD.n165 VSUBS 9.88e-19
C327 VDD.n166 VSUBS 9.88e-19
C328 VDD.n168 VSUBS 9.88e-19
C329 VDD.n169 VSUBS 9.88e-19
C330 VDD.n171 VSUBS 9.88e-19
C331 VDD.n172 VSUBS 9.88e-19
C332 VDD.n174 VSUBS 9.88e-19
C333 VDD.n175 VSUBS 8.47e-19
C334 VDD.n176 VSUBS 0.00454f
C335 VDD.n178 VSUBS 9.88e-19
C336 VDD.n179 VSUBS 6.35e-19
C337 VDD.n181 VSUBS 9.88e-19
C338 VDD.n182 VSUBS 9.88e-19
C339 VDD.n184 VSUBS 9.88e-19
C340 VDD.n185 VSUBS 9.88e-19
C341 VDD.n187 VSUBS 9.88e-19
C342 VDD.n188 VSUBS 5.4e-19
C343 VDD.n189 VSUBS 0.00455f
C344 VDD.n191 VSUBS 9.88e-19
C345 VDD.n192 VSUBS 9.43e-19
C346 VDD.n194 VSUBS 9.88e-19
C347 VDD.n195 VSUBS 9.88e-19
C348 VDD.n197 VSUBS 9.88e-19
C349 VDD.n198 VSUBS 9.88e-19
C350 VDD.n200 VSUBS 9.88e-19
C351 VDD.n201 VSUBS 9.88e-19
C352 VDD.n203 VSUBS 9.88e-19
C353 VDD.n204 VSUBS 9.88e-19
C354 VDD.n206 VSUBS 9.88e-19
C355 VDD.n207 VSUBS 5.35e-19
C356 VDD.n208 VSUBS 0.00452f
C357 VDD.n210 VSUBS 9.88e-19
C358 VDD.n211 VSUBS 9.48e-19
C359 VDD.n213 VSUBS 8.37e-19
C360 VDD.n214 VSUBS 8.37e-19
C361 VDD.n216 VSUBS 8.37e-19
C362 VDD.n217 VSUBS 0.00129f
C363 VDD.n219 VSUBS 9.88e-19
C364 VDD.n220 VSUBS 9.88e-19
C365 VDD.n222 VSUBS 9.88e-19
C366 VDD.n223 VSUBS 9.88e-19
C367 VDD.n225 VSUBS 9.88e-19
C368 VDD.n226 VSUBS 9.88e-19
C369 VDD.n228 VSUBS 9.88e-19
C370 VDD.n229 VSUBS 9.88e-19
C371 VDD.n231 VSUBS 9.88e-19
C372 VDD.n232 VSUBS 9.88e-19
C373 VDD.n234 VSUBS 9.88e-19
C374 VDD.n235 VSUBS 9.88e-19
C375 VDD.n237 VSUBS 9.88e-19
C376 VDD.n238 VSUBS 9.88e-19
C377 VDD.n240 VSUBS 9.88e-19
C378 VDD.n241 VSUBS 9.88e-19
C379 VDD.n261 VSUBS 0.116f
C380 VDD.n263 VSUBS 0.00129f
C381 VDD.n264 VSUBS 0.00129f
C382 VDD.n265 VSUBS 0.00103f
C383 VDD.n266 VSUBS 0.0832f
C384 VDD.n267 VSUBS 0.00103f
C385 VDD.n268 VSUBS 0.00103f
C386 VDD.n269 VSUBS 9.88e-19
C387 VDD.n270 VSUBS 0.0795f
C388 VDD.n271 VSUBS 9.88e-19
C389 VDD.n272 VSUBS 9.88e-19
C390 VDD.n273 VSUBS 9.88e-19
C391 VDD.n274 VSUBS 0.0617f
C392 VDD.n275 VSUBS 9.88e-19
C393 VDD.n276 VSUBS 9.88e-19
C394 VDD.t2 VSUBS 0.0398f
C395 VDD.n277 VSUBS 9.88e-19
C396 VDD.n278 VSUBS 0.0576f
C397 VDD.n279 VSUBS 9.88e-19
C398 VDD.n280 VSUBS 9.88e-19
C399 VDD.n281 VSUBS 9.88e-19
C400 VDD.n282 VSUBS 0.0795f
C401 VDD.n283 VSUBS 9.88e-19
C402 VDD.n284 VSUBS 9.88e-19
C403 VDD.t17 VSUBS 0.0398f
C404 VDD.n285 VSUBS 9.88e-19
C405 VDD.n286 VSUBS 0.056f
C406 VDD.n287 VSUBS 9.88e-19
C407 VDD.n288 VSUBS 9.88e-19
C408 VDD.n289 VSUBS 9.88e-19
C409 VDD.n290 VSUBS 0.0633f
C410 VDD.n291 VSUBS 9.88e-19
C411 VDD.n292 VSUBS 9.88e-19
C412 VDD.n293 VSUBS 9.88e-19
C413 VDD.n294 VSUBS 0.0795f
C414 VDD.n295 VSUBS 9.88e-19
C415 VDD.n296 VSUBS 9.88e-19
C416 VDD.t9 VSUBS 0.0398f
C417 VDD.n297 VSUBS 9.88e-19
C418 VDD.n298 VSUBS 0.0503f
C419 VDD.n299 VSUBS 9.88e-19
C420 VDD.n300 VSUBS 9.88e-19
C421 VDD.n301 VSUBS 9.88e-19
C422 VDD.n302 VSUBS 0.069f
C423 VDD.n303 VSUBS 9.88e-19
C424 VDD.n304 VSUBS 9.88e-19
C425 VDD.n305 VSUBS 9.88e-19
C426 VDD.n306 VSUBS 0.0795f
C427 VDD.n307 VSUBS 9.88e-19
C428 VDD.n308 VSUBS 9.88e-19
C429 VDD.t6 VSUBS 0.0398f
C430 VDD.n309 VSUBS 9.88e-19
C431 VDD.n310 VSUBS 0.0446f
C432 VDD.n311 VSUBS 9.88e-19
C433 VDD.n312 VSUBS 9.88e-19
C434 VDD.n313 VSUBS 9.88e-19
C435 VDD.n314 VSUBS 0.0747f
C436 VDD.n315 VSUBS 9.88e-19
C437 VDD.n316 VSUBS 9.88e-19
C438 VDD.n317 VSUBS 9.88e-19
C439 VDD.n318 VSUBS 0.0787f
C440 VDD.n319 VSUBS 9.88e-19
C441 VDD.n320 VSUBS 9.88e-19
C442 VDD.t12 VSUBS 0.0398f
C443 VDD.n321 VSUBS 9.88e-19
C444 VDD.n322 VSUBS 0.0406f
C445 VDD.n323 VSUBS 9.88e-19
C446 VDD.n324 VSUBS 9.88e-19
C447 VDD.n325 VSUBS 9.88e-19
C448 VDD.n326 VSUBS 0.0795f
C449 VDD.n327 VSUBS 9.88e-19
C450 VDD.n328 VSUBS 9.88e-19
C451 VDD.n329 VSUBS 9.88e-19
C452 VDD.n330 VSUBS 0.073f
C453 VDD.n331 VSUBS 9.88e-19
C454 VDD.n332 VSUBS 9.88e-19
C455 VDD.t0 VSUBS 0.0398f
C456 VDD.n333 VSUBS 9.88e-19
C457 VDD.n334 VSUBS 0.0463f
C458 VDD.n335 VSUBS 9.88e-19
C459 VDD.n336 VSUBS 9.88e-19
C460 VDD.n337 VSUBS 9.88e-19
C461 VDD.n338 VSUBS 0.0795f
C462 VDD.n339 VSUBS 9.88e-19
C463 VDD.n340 VSUBS 7.72e-19
C464 VDD.t30 VSUBS 0.00212f
C465 VDD.t31 VSUBS 0.00212f
C466 VDD.t26 VSUBS 0.00212f
C467 VDD.t27 VSUBS 0.00212f
C468 VDD.t28 VSUBS 0.00212f
C469 VDD.t29 VSUBS 0.00212f
C470 VDD.n341 VSUBS 7.87e-19
C471 VDD.n342 VSUBS 9.88e-19
C472 VDD.n343 VSUBS 9.88e-19
C473 VDD.n344 VSUBS 0.00299f
C474 VDD.n345 VSUBS 9.88e-19
C475 VDD.n346 VSUBS 9.88e-19
C476 VDD.n347 VSUBS 0.00299f
C477 VDD.n348 VSUBS 9.88e-19
C478 VDD.n349 VSUBS 9.88e-19
C479 VDD.n350 VSUBS 0.00299f
C480 VDD.n351 VSUBS 9.88e-19
C481 VDD.n352 VSUBS 9.88e-19
C482 VDD.n353 VSUBS 0.00299f
C483 VDD.n354 VSUBS 9.88e-19
C484 VDD.n355 VSUBS 9.88e-19
C485 VDD.n356 VSUBS 0.00299f
C486 VDD.n357 VSUBS 9.88e-19
C487 VDD.n358 VSUBS 9.88e-19
C488 VDD.n359 VSUBS 0.00299f
C489 VDD.n360 VSUBS 9.88e-19
C490 VDD.n361 VSUBS 9.88e-19
C491 VDD.n362 VSUBS 0.00299f
C492 VDD.n363 VSUBS 9.88e-19
C493 VDD.n364 VSUBS 9.88e-19
C494 VDD.n365 VSUBS 0.00299f
C495 VDD.n366 VSUBS 9.88e-19
C496 VDD.n367 VSUBS 9.88e-19
C497 VDD.n368 VSUBS 0.00299f
C498 VDD.n369 VSUBS 9.88e-19
C499 VDD.n370 VSUBS 9.88e-19
C500 VDD.n371 VSUBS 0.00299f
C501 VDD.n372 VSUBS 9.88e-19
C502 VDD.n373 VSUBS 9.88e-19
C503 VDD.n374 VSUBS 0.00299f
C504 VDD.n375 VSUBS 9.88e-19
C505 VDD.n376 VSUBS 9.88e-19
C506 VDD.n377 VSUBS 0.00299f
C507 VDD.n378 VSUBS 9.88e-19
C508 VDD.n379 VSUBS 9.88e-19
C509 VDD.n380 VSUBS 0.00299f
C510 VDD.n381 VSUBS 9.88e-19
C511 VDD.n382 VSUBS 9.88e-19
C512 VDD.n383 VSUBS 0.00299f
C513 VDD.n384 VSUBS 9.88e-19
C514 VDD.n385 VSUBS 9.88e-19
C515 VDD.n386 VSUBS 0.00299f
C516 VDD.n387 VSUBS 9.88e-19
C517 VDD.n388 VSUBS 9.88e-19
C518 VDD.n389 VSUBS 0.00299f
C519 VDD.n390 VSUBS 9.88e-19
C520 VDD.n391 VSUBS 9.88e-19
C521 VDD.n392 VSUBS 0.00299f
C522 VDD.n393 VSUBS 9.88e-19
C523 VDD.n394 VSUBS 9.88e-19
C524 VDD.n395 VSUBS 0.00299f
C525 VDD.n396 VSUBS 9.88e-19
C526 VDD.n397 VSUBS 9.88e-19
C527 VDD.n398 VSUBS 0.00195f
C528 VDD.t24 VSUBS 0.00212f
C529 VDD.t25 VSUBS 0.00212f
C530 VDD.t34 VSUBS 0.00212f
C531 VDD.t35 VSUBS 0.00212f
C532 VDD.t32 VSUBS 0.00212f
C533 VDD.t33 VSUBS 0.00212f
C534 VDD.n399 VSUBS 9.88e-19
C535 VDD.n400 VSUBS 9.88e-19
C536 VDD.n401 VSUBS 9.88e-19
C537 VDD.n402 VSUBS 9.88e-19
C538 VDD.n403 VSUBS 9.88e-19
C539 VDD.n404 VSUBS 9.88e-19
C540 VDD.n405 VSUBS 9.88e-19
C541 VDD.n406 VSUBS 9.88e-19
C542 VDD.n407 VSUBS 9.88e-19
C543 VDD.n408 VSUBS 9.88e-19
C544 VDD.n409 VSUBS 9.88e-19
C545 VDD.n410 VSUBS 9.88e-19
C546 VDD.n411 VSUBS 9.88e-19
C547 VDD.n412 VSUBS 9.88e-19
C548 VDD.n413 VSUBS 9.88e-19
C549 VDD.n414 VSUBS 9.88e-19
C550 VDD.n415 VSUBS 9.88e-19
C551 VDD.n416 VSUBS 9.88e-19
C552 VDD.n417 VSUBS 7.87e-19
C553 VDD.n418 VSUBS 0.00124f
C554 VDD.n419 VSUBS 0.00104f
C555 VDD.n420 VSUBS 9.48e-19
C556 VDD.n421 VSUBS 0.00482f
C557 VDD.n422 VSUBS 5.35e-19
C558 VDD.n423 VSUBS 9.88e-19
C559 VDD.n424 VSUBS 9.88e-19
C560 VDD.n425 VSUBS 9.88e-19
C561 VDD.n426 VSUBS 9.88e-19
C562 VDD.n427 VSUBS 8.88e-19
C563 VDD.n428 VSUBS 0.00483f
C564 VDD.n429 VSUBS 5.95e-19
C565 VDD.n430 VSUBS 9.88e-19
C566 VDD.n431 VSUBS 9.88e-19
C567 VDD.n432 VSUBS 6.66e-19
C568 VDD.n433 VSUBS 0.00482f
C569 VDD.n434 VSUBS 8.17e-19
C570 VDD.n435 VSUBS 9.88e-19
C571 VDD.n436 VSUBS 9.88e-19
C572 VDD.n437 VSUBS 9.88e-19
C573 VDD.n438 VSUBS 9.88e-19
C574 VDD.n439 VSUBS 5.75e-19
C575 VDD.n440 VSUBS 0.00482f
C576 VDD.n441 VSUBS 9.08e-19
C577 VDD.n442 VSUBS 9.88e-19
C578 VDD.n443 VSUBS 9.88e-19
C579 VDD.n444 VSUBS 9.88e-19
C580 VDD.n445 VSUBS 8.32e-19
C581 VDD.n446 VSUBS 0.00482f
C582 VDD.n447 VSUBS 9.88e-19
C583 VDD.n448 VSUBS 6.51e-19
C584 VDD.n449 VSUBS 9.88e-19
C585 VDD.n450 VSUBS 9.88e-19
C586 VDD.n451 VSUBS 9.88e-19
C587 VDD.n452 VSUBS 9.88e-19
C588 VDD.n453 VSUBS 9.88e-19
C589 VDD.n454 VSUBS 9.88e-19
C590 VDD.n455 VSUBS 9.88e-19
C591 VDD.n456 VSUBS 9.88e-19
C592 VDD.n457 VSUBS 9.88e-19
C593 VDD.n458 VSUBS 8.12e-19
C594 VDD.n459 VSUBS 0.00483f
C595 VDD.n460 VSUBS 9.88e-19
C596 VDD.n461 VSUBS 6.71e-19
C597 VDD.n462 VSUBS 9.88e-19
C598 VDD.n463 VSUBS 9.88e-19
C599 VDD.n464 VSUBS 7.87e-19
C600 VDD.n465 VSUBS 7.87e-19
C601 VDD.n466 VSUBS 0.00119f
C602 VDD.n467 VSUBS 0.00104f
C603 VDD.n468 VSUBS 9.42e-19
C604 VDD.n469 VSUBS 0.00119f
C605 VDD.n470 VSUBS 0.00104f
C606 VDD.n471 VSUBS 9.88e-19
C607 VDD.n472 VSUBS 9.88e-19
C608 VDD.n473 VSUBS 9.88e-19
C609 VDD.n474 VSUBS 9.88e-19
C610 VDD.n475 VSUBS 6.71e-19
C611 VDD.n476 VSUBS 0.00483f
C612 VDD.n477 VSUBS 9.88e-19
C613 VDD.n478 VSUBS 8.12e-19
C614 VDD.n479 VSUBS 9.88e-19
C615 VDD.n480 VSUBS 9.88e-19
C616 VDD.n481 VSUBS 9.88e-19
C617 VDD.n482 VSUBS 9.88e-19
C618 VDD.n483 VSUBS 9.88e-19
C619 VDD.n484 VSUBS 9.88e-19
C620 VDD.n485 VSUBS 9.88e-19
C621 VDD.n486 VSUBS 9.88e-19
C622 VDD.n487 VSUBS 9.88e-19
C623 VDD.n488 VSUBS 6.51e-19
C624 VDD.n489 VSUBS 0.00482f
C625 VDD.n490 VSUBS 9.88e-19
C626 VDD.n491 VSUBS 8.32e-19
C627 VDD.n492 VSUBS 9.88e-19
C628 VDD.n493 VSUBS 9.88e-19
C629 VDD.n494 VSUBS 9.88e-19
C630 VDD.n495 VSUBS 9.08e-19
C631 VDD.n496 VSUBS 0.00482f
C632 VDD.n497 VSUBS 9.88e-19
C633 VDD.n498 VSUBS 5.75e-19
C634 VDD.n499 VSUBS 9.88e-19
C635 VDD.n500 VSUBS 9.88e-19
C636 VDD.n501 VSUBS 9.88e-19
C637 VDD.n502 VSUBS 9.88e-19
C638 VDD.n503 VSUBS 9.88e-19
C639 VDD.n504 VSUBS 9.88e-19
C640 VDD.n505 VSUBS 9.88e-19
C641 VDD.n506 VSUBS 9.88e-19
C642 VDD.n507 VSUBS 9.88e-19
C643 VDD.n508 VSUBS 8.17e-19
C644 VDD.n509 VSUBS 0.00482f
C645 VDD.n510 VSUBS 9.88e-19
C646 VDD.n511 VSUBS 6.66e-19
C647 VDD.n512 VSUBS 9.88e-19
C648 VDD.n513 VSUBS 9.88e-19
C649 VDD.n515 VSUBS 9.88e-19
C650 VDD.n516 VSUBS 9.88e-19
C651 VDD.n517 VSUBS 9.88e-19
C652 VDD.n518 VSUBS 5.95e-19
C653 VDD.n519 VSUBS 0.00483f
C654 VDD.n521 VSUBS 9.88e-19
C655 VDD.n522 VSUBS 8.88e-19
C656 VDD.n523 VSUBS 9.88e-19
C657 VDD.n524 VSUBS 9.88e-19
C658 VDD.n526 VSUBS 9.88e-19
C659 VDD.n527 VSUBS 9.88e-19
C660 VDD.n528 VSUBS 9.88e-19
C661 VDD.n529 VSUBS 9.88e-19
C662 VDD.n531 VSUBS 9.88e-19
C663 VDD.n532 VSUBS 9.88e-19
C664 VDD.n533 VSUBS 9.88e-19
C665 VDD.n534 VSUBS 5.35e-19
C666 VDD.n535 VSUBS 0.00482f
C667 VDD.n537 VSUBS 9.88e-19
C668 VDD.n538 VSUBS 9.48e-19
C669 VDD.n539 VSUBS 8.37e-19
C670 VDD.n540 VSUBS 8.37e-19
C671 VDD.n555 VSUBS 9.88e-19
C672 VDD.n557 VSUBS 9.88e-19
C673 VDD.n558 VSUBS 9.88e-19
C674 VDD.n560 VSUBS 9.88e-19
C675 VDD.n561 VSUBS 9.88e-19
C676 VDD.n563 VSUBS 9.88e-19
C677 VDD.n564 VSUBS 9.88e-19
C678 VDD.n566 VSUBS 9.88e-19
C679 VDD.n567 VSUBS 9.88e-19
C680 VDD.n569 VSUBS 9.88e-19
C681 VDD.n570 VSUBS 9.88e-19
C682 VDD.n572 VSUBS 9.88e-19
C683 VDD.n573 VSUBS 9.88e-19
C684 VDD.n575 VSUBS 9.88e-19
C685 VDD.n576 VSUBS 9.88e-19
C686 VDD.n578 VSUBS 9.88e-19
C687 VDD.n579 VSUBS 9.88e-19
C688 VDD.n581 VSUBS 9.88e-19
C689 VDD.n583 VSUBS 8.37e-19
C690 VDD.n584 VSUBS 0.00124f
C691 VDD.n588 VSUBS 0.113f
C692 VDD.n590 VSUBS 0.00124f
C693 VDD.n591 VSUBS 0.00124f
C694 VDD.n592 VSUBS 9.88e-19
C695 VDD.n593 VSUBS 0.0795f
C696 VDD.n594 VSUBS 9.88e-19
C697 VDD.n595 VSUBS 9.88e-19
C698 VDD.n596 VSUBS 9.88e-19
C699 VDD.n597 VSUBS 0.0795f
C700 VDD.n598 VSUBS 9.88e-19
C701 VDD.n599 VSUBS 9.88e-19
C702 VDD.n600 VSUBS 9.88e-19
C703 VDD.n601 VSUBS 0.0795f
C704 VDD.n602 VSUBS 9.88e-19
C705 VDD.n603 VSUBS 9.88e-19
C706 VDD.t23 VSUBS 0.0398f
C707 VDD.n604 VSUBS 9.88e-19
C708 VDD.n605 VSUBS 0.0406f
C709 VDD.n606 VSUBS 9.88e-19
C710 VDD.n607 VSUBS 9.88e-19
C711 VDD.n608 VSUBS 9.88e-19
C712 VDD.n609 VSUBS 0.0787f
C713 VDD.n610 VSUBS 9.88e-19
C714 VDD.n611 VSUBS 9.88e-19
C715 VDD.n612 VSUBS 9.88e-19
C716 VDD.n613 VSUBS 0.0747f
C717 VDD.n614 VSUBS 9.88e-19
C718 VDD.n615 VSUBS 9.88e-19
C719 VDD.t5 VSUBS 0.0398f
C720 VDD.n616 VSUBS 9.88e-19
C721 VDD.n617 VSUBS 0.0446f
C722 VDD.n618 VSUBS 9.88e-19
C723 VDD.n619 VSUBS 9.88e-19
C724 VDD.n620 VSUBS 9.88e-19
C725 VDD.n621 VSUBS 0.0795f
C726 VDD.n622 VSUBS 9.88e-19
C727 VDD.n623 VSUBS 9.88e-19
C728 VDD.n624 VSUBS 9.88e-19
C729 VDD.n625 VSUBS 0.069f
C730 VDD.n626 VSUBS 9.88e-19
C731 VDD.n627 VSUBS 9.88e-19
C732 VDD.t7 VSUBS 0.0398f
C733 VDD.n628 VSUBS 9.88e-19
C734 VDD.n629 VSUBS 0.0503f
C735 VDD.n630 VSUBS 9.88e-19
C736 VDD.n631 VSUBS 9.88e-19
C737 VDD.n632 VSUBS 9.88e-19
C738 VDD.n633 VSUBS 0.0795f
C739 VDD.n634 VSUBS 9.88e-19
C740 VDD.n635 VSUBS 9.88e-19
C741 VDD.n636 VSUBS 9.88e-19
C742 VDD.n637 VSUBS 0.0633f
C743 VDD.n638 VSUBS 9.88e-19
C744 VDD.n639 VSUBS 9.88e-19
C745 VDD.t1 VSUBS 0.0398f
C746 VDD.n640 VSUBS 9.88e-19
C747 VDD.n641 VSUBS 0.056f
C748 VDD.n642 VSUBS 9.88e-19
C749 VDD.n643 VSUBS 9.88e-19
C750 VDD.n644 VSUBS 9.88e-19
C751 VDD.n645 VSUBS 0.0795f
C752 VDD.n646 VSUBS 9.88e-19
C753 VDD.n647 VSUBS 9.88e-19
C754 VDD.t8 VSUBS 0.0398f
C755 VDD.n648 VSUBS 9.88e-19
C756 VDD.n649 VSUBS 0.0576f
C757 VDD.n650 VSUBS 9.88e-19
C758 VDD.n651 VSUBS 9.88e-19
C759 VDD.n652 VSUBS 9.88e-19
C760 VDD.n653 VSUBS 0.0617f
C761 VDD.n654 VSUBS 9.88e-19
C762 VDD.n655 VSUBS 9.88e-19
C763 VDD.n656 VSUBS 9.88e-19
C764 VDD.n657 VSUBS 0.0795f
C765 VDD.n658 VSUBS 9.88e-19
C766 VDD.n659 VSUBS 9.88e-19
C767 VDD.t18 VSUBS 0.0398f
C768 VDD.n660 VSUBS 9.88e-19
C769 VDD.n661 VSUBS 0.0519f
C770 VDD.n662 VSUBS 9.88e-19
C771 VDD.n663 VSUBS 9.88e-19
C772 VDD.n664 VSUBS 9.88e-19
C773 VDD.n665 VSUBS 0.0674f
C774 VDD.n666 VSUBS 9.88e-19
C775 VDD.n667 VSUBS 7.11e-19
.ends

