* NGSPICE file created from NOR_Layout_flat.ext - technology: gf180mcuC

.subckt NOR_Layout_flat A B OUT VDD VSS
X0 VDD A.t0 a_86_440.t2 VDD.t4 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 OUT A.t1 VSS.t4 VSS.t3 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 OUT B.t1 a_86_440.t1 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 VSS B.t2 OUT.t2 VSS.t0 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
R0 A.n0 A.t2 32.1987
R1 A.n1 A.t0 31.1559
R2 A.n1 A.n0 19.8148
R3 A.n0 A.t1 15.513
R4 A A.n1 4.11202
R5 a_86_440.n2 a_86_440.t2 5.61007
R6 a_86_440.n3 a_86_440.n2 5.61007
R7 a_86_440.n2 a_86_440.n1 2.6005
R8 a_86_440.n1 a_86_440.t1 1.8205
R9 a_86_440.n1 a_86_440.n0 1.8205
R10 VDD.n6 VDD.t1 135.364
R11 VDD.n2 VDD.t0 75.6093
R12 VDD.n12 VDD.t4 75.608
R13 VDD.t1 VDD.n5 23.6892
R14 VDD.n14 VDD.t2 23.6892
R15 VDD.n7 VDD.n4 8.2255
R16 VDD.n15 VDD.n7 8.2255
R17 VDD VDD.n7 6.3005
R18 VDD VDD.n7 6.3005
R19 VDD.n1 VDD.n0 3.1505
R20 VDD.n4 VDD.n3 3.1505
R21 VDD.n5 VDD.n4 3.1505
R22 VDD.n7 VDD.n6 3.1505
R23 VDD.n16 VDD.n15 3.1505
R24 VDD.n15 VDD.n14 3.1505
R25 VDD.n11 VDD.n10 3.1505
R26 VDD.n13 VDD.n9 3.06224
R27 VDD.n2 VDD.n1 1.87215
R28 VDD.n12 VDD.n11 1.87197
R29 VDD.n9 VDD.t3 1.8205
R30 VDD.n9 VDD.n8 1.8205
R31 VDD.n3 VDD.n2 0.641733
R32 VDD.n13 VDD.n12 0.588896
R33 VDD VDD.n3 0.0760357
R34 VDD VDD.n16 0.0760357
R35 VDD.n16 VDD.n13 0.0535357
R36 B.n0 B.t2 26.3326
R37 B.n1 B.t0 21.3791
R38 B.n0 B.t1 21.3791
R39 B.n1 B.n0 20.8576
R40 B B.n1 17.6592
R41 OUT.n4 OUT.n3 3.64746
R42 OUT.n3 OUT.t2 3.2765
R43 OUT.n3 OUT.n2 3.2765
R44 OUT.n4 OUT.n1 3.15224
R45 OUT.n1 OUT.t1 1.8205
R46 OUT.n1 OUT.n0 1.8205
R47 OUT OUT.n4 0.155065
R48 VSS.n3 VSS.t0 254.148
R49 VSS.n8 VSS.t3 254.148
R50 VSS.n2 VSS.n0 6.67264
R51 VSS.n7 VSS.t4 6.67264
R52 VSS.n7 VSS.n6 2.6005
R53 VSS.n5 VSS.n4 2.6005
R54 VSS.n4 VSS.n3 2.6005
R55 VSS.n10 VSS.n9 2.6005
R56 VSS.n9 VSS.n8 2.6005
R57 VSS.n2 VSS.n1 2.6005
R58 VSS.n5 VSS.n2 0.0760357
R59 VSS.n10 VSS.n7 0.0760357
R60 VSS VSS.n5 0.0422857
R61 VSS VSS.n10 0.03425
C0 OUT VDD 0.0163f
C1 VDD A 0.223f
C2 B OUT 0.0855f
C3 B A 0.0431f
C4 OUT A 0.0214f
C5 B VDD 0.276f
.ends

