magic
tech gf180mcuC
magscale 1 10
timestamp 1699872198
<< metal1 >>
rect 31218 15420 31505 15718
rect 31608 15433 33394 15717
rect 32632 14847 34298 15131
rect 1805 14328 2238 14334
rect 1805 14321 3090 14328
rect 1802 14265 1812 14321
rect 1868 14265 1922 14321
rect 1978 14265 2032 14321
rect 2088 14265 2142 14321
rect 2198 14265 3090 14321
rect 1805 14211 3090 14265
rect 5741 14220 5901 14474
rect 6013 14230 6173 14490
rect 15658 14393 17304 14728
rect 1805 14155 1812 14211
rect 1868 14155 1922 14211
rect 1978 14155 2032 14211
rect 2088 14155 2142 14211
rect 2198 14168 3090 14211
rect 2198 14155 2238 14168
rect 1805 14101 2238 14155
rect 1805 14045 1812 14101
rect 1868 14045 1922 14101
rect 1978 14045 2032 14101
rect 2088 14045 2142 14101
rect 2198 14045 2238 14101
rect 1805 14031 2238 14045
rect 2338 13819 2630 13979
rect 37919 13913 39343 14244
rect -720 13122 2569 13200
rect -721 13046 2892 13122
rect -721 12962 2902 13046
rect -720 12801 2902 12962
rect -3602 10407 -3416 10415
rect -3604 10351 -3594 10407
rect -3538 10351 -3484 10407
rect -3428 10369 -3416 10407
rect -720 10369 -288 12801
rect 67186 12776 67702 13060
rect 11649 10953 11809 11220
rect -3428 10351 -288 10369
rect -3602 10297 -288 10351
rect -3602 10241 -3594 10297
rect -3538 10241 -3484 10297
rect -3428 10241 -288 10297
rect -3602 10187 -288 10241
rect -3602 10131 -3594 10187
rect -3538 10131 -3484 10187
rect -3428 10131 -288 10187
rect -3602 10077 -288 10131
rect -3602 10021 -3594 10077
rect -3538 10021 -3484 10077
rect -3428 10021 -288 10077
rect -3602 9967 -288 10021
rect -3602 9911 -3594 9967
rect -3538 9911 -3484 9967
rect -3428 9931 -288 9967
rect -3428 9911 -3416 9931
rect -3602 9896 -3416 9911
rect -3882 9079 575 9529
rect 0 7545 160 7585
rect 8443 6251 8740 6411
rect 14854 5553 15150 5713
rect 2343 5152 2640 5312
rect 3057 5200 3217 5470
rect 5312 5303 5620 5463
rect 11150 5286 11700 5446
rect 6554 4101 6714 4390
rect 3087 1958 3253 2004
rect 11473 1846 11780 2006
rect 8837 1502 9293 1548
rect 12186 971 12480 1131
rect 21903 500 22472 784
rect 15828 0 16342 284
<< via1 >>
rect 1812 14265 1868 14321
rect 1922 14265 1978 14321
rect 2032 14265 2088 14321
rect 2142 14265 2198 14321
rect 1812 14155 1868 14211
rect 1922 14155 1978 14211
rect 2032 14155 2088 14211
rect 2142 14155 2198 14211
rect 1812 14045 1868 14101
rect 1922 14045 1978 14101
rect 2032 14045 2088 14101
rect 2142 14045 2198 14101
rect -3594 10351 -3538 10407
rect -3484 10351 -3428 10407
rect -3594 10241 -3538 10297
rect -3484 10241 -3428 10297
rect -3594 10131 -3538 10187
rect -3484 10131 -3428 10187
rect -3594 10021 -3538 10077
rect -3484 10021 -3428 10077
rect -3594 9911 -3538 9967
rect -3484 9911 -3428 9967
<< metal2 >>
rect 31218 15706 31505 15718
rect 31218 15650 31226 15706
rect 31282 15650 31336 15706
rect 31392 15650 31446 15706
rect 31502 15650 31505 15706
rect 31218 15596 31505 15650
rect 31218 15540 31226 15596
rect 31282 15540 31336 15596
rect 31392 15540 31446 15596
rect 31502 15540 31505 15596
rect 31218 15486 31505 15540
rect 31218 15430 31226 15486
rect 31282 15430 31336 15486
rect 31392 15430 31446 15486
rect 31502 15430 31505 15486
rect 31218 15420 31505 15430
rect 826 14773 1083 14774
rect -7190 14772 1260 14773
rect -7190 14742 1700 14772
rect -7190 14686 1233 14742
rect 1289 14686 1343 14742
rect 1399 14686 1453 14742
rect 1509 14686 1563 14742
rect 1619 14686 1700 14742
rect -7190 14632 1700 14686
rect -7190 14576 1233 14632
rect 1289 14576 1343 14632
rect 1399 14576 1453 14632
rect 1509 14576 1563 14632
rect 1619 14576 1700 14632
rect -7190 14490 1700 14576
rect -7190 12588 -6907 14490
rect 976 14489 1700 14490
rect 1224 14488 1700 14489
rect 1803 14325 2238 14334
rect -3119 14321 2238 14325
rect -3119 14265 1812 14321
rect 1868 14265 1922 14321
rect 1978 14265 2032 14321
rect 2088 14265 2142 14321
rect 2198 14265 2238 14321
rect -3119 14211 2238 14265
rect -3119 14206 1812 14211
rect -3120 14155 1812 14206
rect 1868 14155 1922 14211
rect 1978 14155 2032 14211
rect 2088 14155 2142 14211
rect 2198 14155 2238 14211
rect -3120 14101 2238 14155
rect -3120 14049 1812 14101
rect -3594 10415 -3538 10417
rect -3602 10407 -3416 10415
rect -3602 10351 -3594 10407
rect -3538 10351 -3484 10407
rect -3428 10351 -3416 10407
rect -3602 10297 -3416 10351
rect -3602 10241 -3594 10297
rect -3538 10241 -3484 10297
rect -3428 10241 -3416 10297
rect -3602 10187 -3416 10241
rect -3602 10131 -3594 10187
rect -3538 10131 -3484 10187
rect -3428 10131 -3416 10187
rect -3602 10077 -3416 10131
rect -3602 10021 -3594 10077
rect -3538 10021 -3484 10077
rect -3428 10021 -3416 10077
rect -3602 9967 -3416 10021
rect -3602 9911 -3594 9967
rect -3538 9911 -3484 9967
rect -3428 9911 -3416 9967
rect -3602 9896 -3416 9911
rect -16674 8972 -7712 9200
rect -8066 8577 -7634 8749
rect -3119 6955 -2860 14049
rect 1805 14045 1812 14049
rect 1868 14045 1922 14101
rect 1978 14045 2032 14101
rect 2088 14045 2142 14101
rect 2198 14045 2238 14101
rect 1805 14031 2238 14045
rect 527 13794 1084 13795
rect -1867 13763 1084 13794
rect -1867 13707 554 13763
rect 610 13707 664 13763
rect 720 13707 774 13763
rect 830 13707 884 13763
rect 940 13707 994 13763
rect 1050 13707 1084 13763
rect -1867 13653 1084 13707
rect -1869 13597 554 13653
rect 610 13597 664 13653
rect 720 13597 774 13653
rect 830 13597 884 13653
rect 940 13597 994 13653
rect 1050 13597 1084 13653
rect -1869 13496 1084 13597
rect -4565 6798 -2860 6955
rect -3659 6703 -2860 6798
rect -8166 6243 -7794 6415
rect -16479 5777 -7620 6020
rect -7575 5362 -7205 5532
rect -1867 2259 -1568 13496
rect 11381 11470 11541 12170
rect -8069 1978 -1434 2259
<< via2 >>
rect 31226 15650 31282 15706
rect 31336 15650 31392 15706
rect 31446 15650 31502 15706
rect 31226 15540 31282 15596
rect 31336 15540 31392 15596
rect 31446 15540 31502 15596
rect 31226 15430 31282 15486
rect 31336 15430 31392 15486
rect 31446 15430 31502 15486
rect 1233 14686 1289 14742
rect 1343 14686 1399 14742
rect 1453 14686 1509 14742
rect 1563 14686 1619 14742
rect 1233 14576 1289 14632
rect 1343 14576 1399 14632
rect 1453 14576 1509 14632
rect 1563 14576 1619 14632
rect 554 13707 610 13763
rect 664 13707 720 13763
rect 774 13707 830 13763
rect 884 13707 940 13763
rect 994 13707 1050 13763
rect 554 13597 610 13653
rect 664 13597 720 13653
rect 774 13597 830 13653
rect 884 13597 940 13653
rect 994 13597 1050 13653
<< metal3 >>
rect 374 15706 31505 15718
rect 374 15650 31226 15706
rect 31282 15650 31336 15706
rect 31392 15650 31446 15706
rect 31502 15650 31505 15706
rect 374 15596 31505 15650
rect 374 15540 31226 15596
rect 31282 15540 31336 15596
rect 31392 15540 31446 15596
rect 31502 15540 31505 15596
rect 374 15491 31505 15540
rect 374 15486 31509 15491
rect 374 15430 31226 15486
rect 31282 15430 31336 15486
rect 31392 15430 31446 15486
rect 31502 15430 31509 15486
rect 374 15207 31509 15430
rect 374 13795 957 15207
rect 1233 14772 9208 14935
rect 1224 14742 9208 14772
rect 1223 14686 1233 14742
rect 1289 14686 1343 14742
rect 1399 14686 1453 14742
rect 1509 14686 1563 14742
rect 1619 14686 9208 14742
rect 1224 14632 9208 14686
rect 1224 14576 1233 14632
rect 1289 14576 1343 14632
rect 1399 14576 1453 14632
rect 1509 14576 1563 14632
rect 1619 14576 9208 14632
rect 1224 14488 9208 14576
rect 374 13763 1084 13795
rect 374 13707 554 13763
rect 610 13707 664 13763
rect 720 13707 774 13763
rect 830 13707 884 13763
rect 940 13707 994 13763
rect 1050 13707 1084 13763
rect 374 13653 1084 13707
rect 374 13597 554 13653
rect 610 13597 664 13653
rect 720 13597 774 13653
rect 830 13597 884 13653
rect 940 13597 994 13653
rect 1050 13597 1084 13653
rect 374 13509 1084 13597
rect 527 13497 1084 13509
rect 8788 13105 9208 14488
rect 8788 12886 18923 13105
rect 8788 12602 20892 12886
rect -3303 5884 9735 6044
rect -3303 5277 -3143 5884
rect -16666 5117 -3143 5277
rect 17588 4192 18122 4476
rect 30954 3657 31976 4149
rect 17578 1984 18112 2268
rect 32404 1645 33506 2137
rect 9670 717 10450 877
<< metal5 >>
rect -8154 7874 -7942 8396
use filter_res_magic  filter_res_magic_0
timestamp 1699205295
transform 1 0 -7493 0 1 9552
box -8879 -9282 6514 5616
use Folded_Diff_Op_Amp_Layout  Folded_Diff_Op_Amp_Layout_0
timestamp 1699707096
transform 1 0 486 0 1 9157
box -486 -9157 67202 6560
<< labels >>
flabel metal1 33652 15036 33652 15036 0 FreeSans 1600 0 0 0 VOUT_N
port 5 nsew
flabel metal1 32948 15654 32948 15654 0 FreeSans 1600 0 0 0 VOUT_P
port 6 nsew
flabel metal1 38509 14010 38509 14010 0 FreeSans 1600 0 0 0 VDD
port 7 nsew
flabel metal1 16460 14550 16460 14550 0 FreeSans 1600 0 0 0 VSS
port 9 nsew
flabel metal1 -1080 10090 -1080 10090 0 FreeSans 1600 0 0 0 VOUT_OPAMP_P
port 11 nsew
flabel metal2 -3040 7540 -3040 7540 0 FreeSans 1600 0 0 0 VOUT_OPAMP_N
port 12 nsew
flabel metal2 -16437 5875 -16437 5875 0 FreeSans 1600 0 0 0 VIN_N1
port 1 nsew
flabel metal3 -16560 5220 -16560 5220 0 FreeSans 1600 0 0 0 VCM1
port 13 nsew
flabel metal2 -16600 9060 -16600 9060 0 FreeSans 1600 0 0 0 VIN_P1
port 14 nsew
flabel metal2 -7400 5460 -7400 5460 0 FreeSans 1600 0 0 0 R3_R7_1
port 15 nsew
flabel metal2 -7980 6330 -7980 6330 0 FreeSans 1600 0 0 0 R7_R8_R10_C1
port 16 nsew
flabel metal1 3160 1980 3160 1980 0 FreeSans 1600 0 0 0 IB21
port 17 nsew
flabel metal1 2440 5270 2440 5270 0 FreeSans 1600 0 0 0 IBIAS11
port 18 nsew
flabel metal1 3130 5380 3130 5380 0 FreeSans 1600 0 0 0 VBM1
port 19 nsew
flabel metal1 5490 5430 5490 5430 0 FreeSans 1600 0 0 0 VBIASN1
port 20 nsew
flabel metal1 8940 1510 8940 1510 0 FreeSans 1600 0 0 0 IB31
port 21 nsew
flabel metal3 9880 760 9880 760 0 FreeSans 1600 0 0 0 IBS1
port 22 nsew
flabel metal1 12290 1080 12290 1080 0 FreeSans 1600 0 0 0 VB21
port 23 nsew
flabel metal1 11560 1940 11560 1940 0 FreeSans 1600 0 0 0 VB31
port 24 nsew
flabel metal1 8540 6320 8540 6320 0 FreeSans 1600 0 0 0 VB41
port 25 nsew
flabel metal1 6620 4310 6620 4310 0 FreeSans 1600 0 0 0 VCD1
port 26 nsew
flabel metal1 5800 14420 5800 14420 0 FreeSans 1600 0 0 0 IND1
port 27 nsew
flabel metal1 6130 14390 6130 14390 0 FreeSans 1600 0 0 0 IPD1
port 28 nsew
flabel metal2 11480 12040 11480 12040 0 FreeSans 1600 0 0 0 OUT2_1
port 29 nsew
flabel metal1 11710 11070 11710 11070 0 FreeSans 1600 0 0 0 OUT1_1
port 30 nsew
flabel metal1 16030 180 16030 180 0 FreeSans 1600 0 0 0 IBIAS3_1
port 32 nsew
flabel metal3 17890 4430 17890 4430 0 FreeSans 1600 0 0 0 IB4_1
port 33 nsew
flabel metal1 22190 700 22190 700 0 FreeSans 1600 0 0 0 IBIAS4_1
port 34 nsew
flabel metal3 17870 2220 17870 2220 0 FreeSans 1600 0 0 0 IVS_1
port 35 nsew
flabel metal1 67400 13010 67400 13010 0 FreeSans 1600 0 0 0 IBIAS2_1
port 36 nsew
flabel metal1 14950 5670 14950 5670 0 FreeSans 1600 0 0 0 VB1_1
port 37 nsew
flabel metal1 2400 13930 2400 13930 0 FreeSans 1600 0 0 0 BD_1
port 38 nsew
flabel metal2 -7820 8650 -7820 8650 0 FreeSans 1600 0 0 0 R_1
port 39 nsew
flabel metal5 -8120 8070 -8120 8070 0 FreeSans 1600 0 0 0 R11_1
port 40 nsew
flabel metal3 32800 1940 32800 1940 0 FreeSans 1600 0 0 0 OPAMP_C_1
port 41 nsew
flabel metal3 31560 3900 31560 3900 0 FreeSans 1600 0 0 0 OPAMP_C1_1
port 42 nsew
flabel metal1 11360 5390 11360 5390 0 FreeSans 1600 0 0 0 VOUT_1_1
port 43 nsew
<< end >>
