magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2233 -2045 2233 2045
<< psubdiff >>
rect -233 23 233 45
rect -233 -23 -211 23
rect 211 -23 233 23
rect -233 -45 233 -23
<< psubdiffcont >>
rect -211 -23 211 23
<< metal1 >>
rect -222 23 222 34
rect -222 -23 -211 23
rect 211 -23 222 23
rect -222 -34 222 -23
<< end >>
