magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2044 -2000 3584 10000
<< metal1 >>
rect -44 0 200 8000
rect 340 0 1584 8000
<< metal2 >>
rect -44 0 200 8000
rect 340 0 1584 8000
use M2_M1_CDNS_69033583165692  M2_M1_CDNS_69033583165692_0
timestamp 1713338890
transform 1 0 78 0 1 3994
box -90 -3944 90 3944
use M2_M1_CDNS_69033583165693  M2_M1_CDNS_69033583165693_0
timestamp 1713338890
transform 1 0 962 0 1 3994
box -596 -3944 596 3944
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_0
timestamp 1713338890
transform 1 0 78 0 1 5502
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165605  M3_M2_CDNS_69033583165605_1
timestamp 1713338890
transform 1 0 78 0 1 2315
box -109 -1458 109 1458
use M3_M2_CDNS_69033583165657  M3_M2_CDNS_69033583165657_0
timestamp 1713338890
transform 1 0 78 0 1 309
box -109 -251 109 251
use M3_M2_CDNS_69033583165685  M3_M2_CDNS_69033583165685_0
timestamp 1713338890
transform 1 0 78 0 1 7603
box -109 -322 109 322
<< end >>
