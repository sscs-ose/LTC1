* NGSPICE file created from pga_res_magice_parallel_flat.ext - technology: gf180mcuC

.subckt pex_pga_res_magice_parallel A B C D E F G H VDD
X0 a_7877_692.t1 a_7597_390.t1 VDD.t12 ppolyf_u r_width=1u r_length=1u
X1 a_2277_692.t0 a_2277_390.t0 VDD.t30 ppolyf_u r_width=1u r_length=1u
X2 a_1437_n1796.t1 a_2837_n794.t1 VDD.t37 ppolyf_u r_width=1u r_length=1u
X3 C.t0 a_1997_1042.t0 VDD.t0 ppolyf_u r_width=1u r_length=1u
X4 G.t8 G.t9 VDD.t36 ppolyf_u r_width=1u r_length=1u
X5 a_3957_1344.t0 a_3957_1042.t1 VDD.t26 ppolyf_u r_width=1u r_length=1u
X6 a_7317_692.t0 a_5917_1694.t0 VDD.t21 ppolyf_u r_width=1u r_length=1u
X7 a_1437_n1796.t0 E.t3 VDD.t36 ppolyf_u r_width=1u r_length=1u
X8 a_4517_n794.t0 a_4237_n2098.t0 VDD.t20 ppolyf_u r_width=1u r_length=1u
X9 a_5917_1344.t0 a_5917_1042.t0 VDD.t8 ppolyf_u r_width=1u r_length=1u
X10 a_3957_n1796.t1 a_2557_n2098.t0 VDD.t26 ppolyf_u r_width=1u r_length=1u
X11 a_6757_692.t1 a_6757_390.t1 VDD.t39 ppolyf_u r_width=1u r_length=1u
X12 a_7597_n1144.t0 a_6477_n2098.t0 VDD.t4 ppolyf_u r_width=1u r_length=1u
X13 E.t7 a_1157_390.t3 VDD.t5 ppolyf_u r_width=1u r_length=1u
X14 a_8437_n1446.t0 a_6197_n2098.t1 VDD.t2 ppolyf_u r_width=1u r_length=1u
X15 a_4237_n1144.t1 a_4517_n1446.t1 VDD.t32 ppolyf_u r_width=1u r_length=1u
X16 G.t1 G.t2 VDD.t0 ppolyf_u r_width=1u r_length=1u
X17 a_1157_n492.t0 a_1157_n492.t1 VDD.t36 ppolyf_u r_width=1u r_length=1u
X18 a_3957_n492.t0 a_3957_n794.t0 VDD.t26 ppolyf_u r_width=1u r_length=1u
X19 a_8157_n1446.t1 a_8717_n2098.t0 VDD.t11 ppolyf_u r_width=1u r_length=1u
X20 a_5637_n492.t1 a_5917_n794.t0 VDD.t8 ppolyf_u r_width=1u r_length=1u
X21 a_1717_1694.t0 a_1717_692.t0 VDD.t34 ppolyf_u r_width=1u r_length=1u
X22 a_4517_1344.t0 a_4237_1042.t1 VDD.t32 ppolyf_u r_width=1u r_length=1u
X23 a_5357_692.t0 a_5637_390.t0 VDD.t1 ppolyf_u r_width=1u r_length=1u
X24 a_1157_n1446.t0 a_1997_n2098.t2 VDD.t0 ppolyf_u r_width=1u r_length=1u
X25 a_1717_n794.t0 a_1717_n1796.t0 VDD.t34 ppolyf_u r_width=1u r_length=1u
X26 C.t1 a_1717_n1144.t0 VDD.t34 ppolyf_u r_width=1u r_length=1u
X27 a_3677_n1446.t1 a_4237_n2098.t1 VDD.t31 ppolyf_u r_width=1u r_length=1u
X28 a_4517_n492.t1 a_4517_n794.t1 VDD.t32 ppolyf_u r_width=1u r_length=1u
X29 a_1157_1344.t1 A.t1 VDD.t5 ppolyf_u r_width=1u r_length=1u
X30 a_3677_1344.t0 a_3677_1042.t0 VDD.t27 ppolyf_u r_width=1u r_length=1u
X31 a_4517_692.t1 a_4517_390.t1 VDD.t32 ppolyf_u r_width=1u r_length=1u
X32 a_6757_n1796.t1 a_5917_n1446.t1 VDD.t39 ppolyf_u r_width=1u r_length=1u
X33 a_1997_1996.t0 a_1997_1996.t1 VDD.t7 ppolyf_u r_width=1u r_length=1u
X34 a_5637_1344.t0 a_5357_1042.t1 VDD.t1 ppolyf_u r_width=1u r_length=1u
X35 a_6757_n794.t0 a_6757_n1796.t0 VDD.t21 ppolyf_u r_width=1u r_length=1u
X36 a_3957_692.t0 a_3957_390.t0 VDD.t26 ppolyf_u r_width=1u r_length=1u
X37 a_1717_1996.t0 a_1717_1694.t1 VDD.t33 ppolyf_u r_width=1u r_length=1u
X38 B.t1 a_8997_n1796.t1 VDD.t35 ppolyf_u r_width=1u r_length=1u
X39 a_1157_n492.t2 E.t6 VDD.t5 ppolyf_u r_width=1u r_length=1u
X40 a_3677_n492.t0 a_3397_n794.t0 VDD.t27 ppolyf_u r_width=1u r_length=1u
X41 a_2277_n1796.t1 G.t3 VDD.t30 ppolyf_u r_width=1u r_length=1u
X42 a_3117_n492.t1 a_2837_n794.t0 VDD.t7 ppolyf_u r_width=1u r_length=1u
X43 a_2277_1344.t1 a_1997_1042.t1 VDD.t30 ppolyf_u r_width=1u r_length=1u
X44 a_5637_n492.t0 a_5357_n794.t0 VDD.t1 ppolyf_u r_width=1u r_length=1u
X45 a_3957_1694.t1 a_3957_692.t1 VDD.t38 ppolyf_u r_width=1u r_length=1u
X46 a_3957_n1446.t1 a_1717_n2098.t1 VDD.t38 ppolyf_u r_width=1u r_length=1u
X47 a_2277_1344.t0 a_4237_1042.t0 VDD.t31 ppolyf_u r_width=1u r_length=1u
X48 a_2837_692.t1 a_1437_1694.t1 VDD.t37 ppolyf_u r_width=1u r_length=1u
X49 a_1717_n1796.t1 a_1717_n2098.t0 VDD.t33 ppolyf_u r_width=1u r_length=1u
X50 a_6757_1344.t1 a_6477_1042.t1 VDD.t39 ppolyf_u r_width=1u r_length=1u
X51 a_5357_n1144.t1 a_4517_n1796.t1 VDD.t6 ppolyf_u r_width=1u r_length=1u
X52 a_2837_1996.t0 a_1157_390.t0 VDD.t37 ppolyf_u r_width=1u r_length=1u
X53 a_6197_n1446.t1 a_7037_n2098.t0 VDD.t18 ppolyf_u r_width=1u r_length=1u
X54 a_6757_1344.t0 a_8717_1042.t1 VDD.t11 ppolyf_u r_width=1u r_length=1u
X55 a_7597_n1144.t1 a_7877_n1446.t1 VDD.t12 ppolyf_u r_width=1u r_length=1u
X56 a_2277_n492.t0 a_2277_n794.t1 VDD.t30 ppolyf_u r_width=1u r_length=1u
X57 a_8157_n492.t1 a_9557_n2098.t1 VDD.t19 ppolyf_u r_width=1u r_length=1u
X58 a_4797_n492.t1 a_3957_n1144.t1 VDD.t38 ppolyf_u r_width=1u r_length=1u
X59 a_1717_692.t1 G.t11 VDD.t33 ppolyf_u r_width=1u r_length=1u
X60 a_2277_n492.t1 a_3677_n1144.t1 VDD.t31 ppolyf_u r_width=1u r_length=1u
X61 a_1997_1996.t2 a_1997_1996.t3 VDD.t29 ppolyf_u r_width=1u r_length=1u
X62 a_6757_n492.t1 a_6757_n794.t1 VDD.t39 ppolyf_u r_width=1u r_length=1u
X63 a_1997_1996.t4 a_1157_1344.t0 VDD.t0 ppolyf_u r_width=1u r_length=1u
X64 a_4517_1694.t0 a_5357_1042.t0 VDD.t6 ppolyf_u r_width=1u r_length=1u
X65 a_7877_1344.t0 a_7597_1042.t0 VDD.t12 ppolyf_u r_width=1u r_length=1u
X66 a_8437_1042.t0 F.t0 VDD.t2 ppolyf_u r_width=1u r_length=1u
X67 a_6757_n492.t0 a_8157_n1144.t1 VDD.t11 ppolyf_u r_width=1u r_length=1u
X68 E.t2 a_1437_1694.t0 VDD.t36 ppolyf_u r_width=1u r_length=1u
X69 VDD.t16 VDD.t17 VDD.t13 ppolyf_u r_width=1u r_length=1u
X70 a_2557_1996.t0 a_3957_1694.t0 VDD.t26 ppolyf_u r_width=1u r_length=1u
X71 a_6757_1694.t0 a_6757_692.t0 VDD.t21 ppolyf_u r_width=1u r_length=1u
X72 a_8997_1694.t1 B.t3 VDD.t35 ppolyf_u r_width=1u r_length=1u
X73 a_1997_n2098.t4 a_1997_n2098.t5 VDD.t29 ppolyf_u r_width=1u r_length=1u
X74 a_3677_n492.t1 a_5077_n2098.t0 VDD.t20 ppolyf_u r_width=1u r_length=1u
X75 a_5637_1996.t0 a_5917_1694.t1 VDD.t8 ppolyf_u r_width=1u r_length=1u
X76 a_3117_n492.t0 a_3397_n794.t1 VDD.t29 ppolyf_u r_width=1u r_length=1u
X77 VDD.t40 VDD.t41 VDD.t22 ppolyf_u r_width=1u r_length=1u
X78 a_7597_n1796.t1 a_7317_n2098.t0 VDD.t4 ppolyf_u r_width=1u r_length=1u
X79 a_2277_n794.t0 a_2277_n1796.t0 VDD.t37 ppolyf_u r_width=1u r_length=1u
X80 a_4517_n1796.t0 a_1997_n2098.t3 VDD.t32 ppolyf_u r_width=1u r_length=1u
X81 a_7597_n492.t1 a_7877_n794.t1 VDD.t12 ppolyf_u r_width=1u r_length=1u
X82 a_5077_n492.t1 a_5357_n794.t1 VDD.t6 ppolyf_u r_width=1u r_length=1u
X83 VDD.t44 VDD.t45 VDD.t13 ppolyf_u r_width=1u r_length=1u
X84 a_7877_692.t0 a_8157_390.t0 VDD.t25 ppolyf_u r_width=1u r_length=1u
X85 VDD.t50 VDD.t51 VDD.t13 ppolyf_u r_width=1u r_length=1u
X86 a_8157_n1144.t0 a_8157_n1446.t0 VDD.t25 ppolyf_u r_width=1u r_length=1u
X87 a_4517_1344.t1 a_6477_1042.t0 VDD.t3 ppolyf_u r_width=1u r_length=1u
X88 a_9557_n492.t1 F.t2 VDD.t35 ppolyf_u r_width=1u r_length=1u
X89 a_5917_n1796.t0 a_7317_n794.t1 VDD.t21 ppolyf_u r_width=1u r_length=1u
X90 B.t0 a_8717_1042.t0 VDD.t10 ppolyf_u r_width=1u r_length=1u
X91 a_7317_692.t1 a_7597_390.t0 VDD.t4 ppolyf_u r_width=1u r_length=1u
X92 a_2557_1996.t1 a_1717_1344.t1 VDD.t34 ppolyf_u r_width=1u r_length=1u
X93 a_8437_1344.t1 a_8437_1042.t1 VDD.t28 ppolyf_u r_width=1u r_length=1u
X94 VDD.t42 VDD.t43 VDD.t22 ppolyf_u r_width=1u r_length=1u
X95 a_1997_1996.t5 a_4517_1694.t1 VDD.t32 ppolyf_u r_width=1u r_length=1u
X96 a_6197_1042.t1 a_3957_390.t1 VDD.t18 ppolyf_u r_width=1u r_length=1u
X97 a_4517_n492.t0 a_5917_n1144.t0 VDD.t3 ppolyf_u r_width=1u r_length=1u
X98 a_1717_n1446.t0 a_2557_n2098.t1 VDD.t34 ppolyf_u r_width=1u r_length=1u
X99 H.t1 a_8997_n794.t0 VDD.t10 ppolyf_u r_width=1u r_length=1u
X100 a_4237_1996.t0 a_4517_692.t0 VDD.t20 ppolyf_u r_width=1u r_length=1u
X101 a_5917_1042.t1 a_4517_390.t0 VDD.t3 ppolyf_u r_width=1u r_length=1u
X102 a_6197_n1144.t0 a_6197_n1446.t0 VDD.t9 ppolyf_u r_width=1u r_length=1u
X103 D.t3 a_8437_n794.t1 VDD.t28 ppolyf_u r_width=1u r_length=1u
X104 a_6477_1996.t0 a_7597_1042.t1 VDD.t4 ppolyf_u r_width=1u r_length=1u
X105 E.t0 E.t1 VDD.t5 ppolyf_u r_width=1u r_length=1u
X106 a_6197_1694.t1 a_6197_692.t1 VDD.t18 ppolyf_u r_width=1u r_length=1u
X107 a_1997_n2098.t0 a_1997_n2098.t1 VDD.t7 ppolyf_u r_width=1u r_length=1u
X108 a_3397_1996.t1 a_3677_1694.t0 VDD.t27 ppolyf_u r_width=1u r_length=1u
X109 a_8717_1996.t1 a_8997_692.t0 VDD.t19 ppolyf_u r_width=1u r_length=1u
X110 a_2837_1996.t1 a_3117_1694.t1 VDD.t7 ppolyf_u r_width=1u r_length=1u
X111 a_5357_n1144.t0 a_5637_n1446.t1 VDD.t1 ppolyf_u r_width=1u r_length=1u
X112 a_5637_1996.t1 a_5357_1694.t1 VDD.t1 ppolyf_u r_width=1u r_length=1u
X113 a_5917_n794.t1 a_7317_n2098.t1 VDD.t21 ppolyf_u r_width=1u r_length=1u
X114 a_5077_n492.t0 a_3677_n1796.t0 VDD.t20 ppolyf_u r_width=1u r_length=1u
X115 a_5357_692.t1 a_5077_390.t0 VDD.t6 ppolyf_u r_width=1u r_length=1u
X116 D.t2 a_9557_n2098.t0 VDD.t35 ppolyf_u r_width=1u r_length=1u
X117 VDD.t23 VDD.t24 VDD.t22 ppolyf_u r_width=1u r_length=1u
X118 a_7597_n492.t0 a_7317_n794.t0 VDD.t4 ppolyf_u r_width=1u r_length=1u
X119 VDD.t14 VDD.t15 VDD.t13 ppolyf_u r_width=1u r_length=1u
X120 a_3957_n492.t1 a_6197_n1144.t1 VDD.t18 ppolyf_u r_width=1u r_length=1u
X121 a_6197_1344.t1 a_6197_1042.t0 VDD.t9 ppolyf_u r_width=1u r_length=1u
X122 a_9557_n492.t0 a_8157_n1796.t1 VDD.t19 ppolyf_u r_width=1u r_length=1u
X123 a_3957_1042.t0 a_4797_390.t0 VDD.t38 ppolyf_u r_width=1u r_length=1u
X124 G.t0 a_2277_1694.t0 VDD.t30 ppolyf_u r_width=1u r_length=1u
X125 a_1717_1996.t1 a_3957_1344.t1 VDD.t38 ppolyf_u r_width=1u r_length=1u
X126 a_8157_1344.t1 a_8157_1042.t0 VDD.t25 ppolyf_u r_width=1u r_length=1u
X127 A.t0 a_1157_n1446.t1 VDD.t5 ppolyf_u r_width=1u r_length=1u
X128 a_4237_1996.t1 a_3677_1344.t1 VDD.t31 ppolyf_u r_width=1u r_length=1u
X129 a_5917_1344.t1 a_6757_1694.t1 VDD.t39 ppolyf_u r_width=1u r_length=1u
X130 F.t3 a_9557_390.t1 VDD.t35 ppolyf_u r_width=1u r_length=1u
X131 a_3677_n1144.t0 a_3677_n1446.t0 VDD.t27 ppolyf_u r_width=1u r_length=1u
X132 a_3677_1042.t1 a_2277_390.t1 VDD.t31 ppolyf_u r_width=1u r_length=1u
X133 a_5357_n1796.t1 a_5077_n2098.t1 VDD.t6 ppolyf_u r_width=1u r_length=1u
X134 a_8717_1996.t0 a_8157_1344.t0 VDD.t11 ppolyf_u r_width=1u r_length=1u
X135 a_4797_n492.t0 a_6197_n794.t1 VDD.t9 ppolyf_u r_width=1u r_length=1u
X136 a_7597_n1796.t0 a_7877_n2098.t0 VDD.t12 ppolyf_u r_width=1u r_length=1u
X137 a_3397_692.t1 a_3677_390.t0 VDD.t27 ppolyf_u r_width=1u r_length=1u
X138 a_8157_n492.t0 a_7877_n794.t0 VDD.t25 ppolyf_u r_width=1u r_length=1u
X139 a_8437_n1144.t1 a_8437_n1446.t1 VDD.t28 ppolyf_u r_width=1u r_length=1u
X140 a_3397_1996.t0 a_3117_1694.t0 VDD.t29 ppolyf_u r_width=1u r_length=1u
X141 a_8437_1694.t1 a_8437_692.t1 VDD.t2 ppolyf_u r_width=1u r_length=1u
X142 a_8157_1042.t1 a_6757_390.t0 VDD.t11 ppolyf_u r_width=1u r_length=1u
X143 a_5077_1996.t0 a_5357_1694.t0 VDD.t6 ppolyf_u r_width=1u r_length=1u
X144 a_2837_692.t0 a_3117_390.t1 VDD.t7 ppolyf_u r_width=1u r_length=1u
X145 VDD.t52 VDD.t53 VDD.t13 ppolyf_u r_width=1u r_length=1u
X146 a_7877_1996.t0 a_7597_1694.t1 VDD.t12 ppolyf_u r_width=1u r_length=1u
X147 a_7317_1996.t1 a_5917_692.t1 VDD.t21 ppolyf_u r_width=1u r_length=1u
X148 a_3117_n1796.t1 a_3397_n2098.t1 VDD.t29 ppolyf_u r_width=1u r_length=1u
X149 a_9557_1996.t0 D.t1 VDD.t35 ppolyf_u r_width=1u r_length=1u
X150 a_1717_1042.t1 C.t2 VDD.t34 ppolyf_u r_width=1u r_length=1u
X151 VDD.t46 VDD.t47 VDD.t22 ppolyf_u r_width=1u r_length=1u
X152 F.t1 a_8437_n1144.t0 VDD.t2 ppolyf_u r_width=1u r_length=1u
X153 G.t4 G.t5 VDD.t0 ppolyf_u r_width=1u r_length=1u
X154 a_1157_n492.t3 a_2837_n2098.t1 VDD.t37 ppolyf_u r_width=1u r_length=1u
X155 a_6477_n1144.t0 a_4517_n1446.t0 VDD.t3 ppolyf_u r_width=1u r_length=1u
X156 a_8157_n1796.t0 a_7877_n2098.t1 VDD.t25 ppolyf_u r_width=1u r_length=1u
X157 a_6477_1996.t1 a_5637_1344.t1 VDD.t3 ppolyf_u r_width=1u r_length=1u
X158 a_8717_n1144.t1 B.t2 VDD.t10 ppolyf_u r_width=1u r_length=1u
X159 a_7877_1344.t1 a_8997_1694.t0 VDD.t10 ppolyf_u r_width=1u r_length=1u
X160 a_1157_390.t1 a_1157_390.t2 VDD.t36 ppolyf_u r_width=1u r_length=1u
X161 a_5917_n1144.t1 a_5917_n1446.t0 VDD.t8 ppolyf_u r_width=1u r_length=1u
X162 a_7037_1996.t1 a_8437_1694.t0 VDD.t28 ppolyf_u r_width=1u r_length=1u
X163 a_5917_692.t0 a_5637_390.t1 VDD.t8 ppolyf_u r_width=1u r_length=1u
X164 a_5077_1996.t1 a_3677_390.t1 VDD.t20 ppolyf_u r_width=1u r_length=1u
X165 a_6197_n1796.t0 a_6197_n2098.t0 VDD.t9 ppolyf_u r_width=1u r_length=1u
X166 G.t6 G.t7 VDD.t36 ppolyf_u r_width=1u r_length=1u
X167 a_7317_1996.t0 a_7597_1694.t0 VDD.t4 ppolyf_u r_width=1u r_length=1u
X168 a_3117_n1796.t0 a_2837_n2098.t0 VDD.t7 ppolyf_u r_width=1u r_length=1u
X169 a_7037_1996.t0 a_6197_1344.t0 VDD.t18 ppolyf_u r_width=1u r_length=1u
X170 a_3957_n1144.t0 a_3957_n1446.t0 VDD.t26 ppolyf_u r_width=1u r_length=1u
X171 a_9557_1996.t1 a_8157_390.t1 VDD.t19 ppolyf_u r_width=1u r_length=1u
X172 a_5357_n1796.t0 a_5637_n2098.t0 VDD.t1 ppolyf_u r_width=1u r_length=1u
X173 a_8437_n794.t0 a_8437_n1796.t0 VDD.t2 ppolyf_u r_width=1u r_length=1u
X174 VDD.t48 VDD.t49 VDD.t22 ppolyf_u r_width=1u r_length=1u
X175 VDD.t56 VDD.t57 VDD.t13 ppolyf_u r_width=1u r_length=1u
X176 a_8717_n1144.t0 a_6757_n1446.t0 VDD.t11 ppolyf_u r_width=1u r_length=1u
X177 a_6197_1996.t1 a_6197_1694.t0 VDD.t9 ppolyf_u r_width=1u r_length=1u
X178 a_7877_1996.t1 a_8157_1694.t1 VDD.t25 ppolyf_u r_width=1u r_length=1u
X179 E.t4 E.t5 VDD.t5 ppolyf_u r_width=1u r_length=1u
X180 a_6197_692.t0 a_4797_390.t1 VDD.t9 ppolyf_u r_width=1u r_length=1u
X181 a_1997_n1144.t1 C.t3 VDD.t0 ppolyf_u r_width=1u r_length=1u
X182 a_3677_n1796.t1 a_3397_n2098.t0 VDD.t27 ppolyf_u r_width=1u r_length=1u
X183 a_4237_n1144.t0 a_2277_n1446.t0 VDD.t31 ppolyf_u r_width=1u r_length=1u
X184 a_6477_n1144.t1 a_6757_n1446.t1 VDD.t39 ppolyf_u r_width=1u r_length=1u
X185 VDD.t54 VDD.t55 VDD.t22 ppolyf_u r_width=1u r_length=1u
X186 a_8437_n1796.t1 a_7037_n2098.t1 VDD.t28 ppolyf_u r_width=1u r_length=1u
X187 a_6197_1996.t0 a_8437_1344.t0 VDD.t2 ppolyf_u r_width=1u r_length=1u
X188 a_3677_1694.t1 a_5077_390.t1 VDD.t20 ppolyf_u r_width=1u r_length=1u
X189 a_1717_1344.t0 a_1717_1042.t0 VDD.t33 ppolyf_u r_width=1u r_length=1u
X190 a_8157_1694.t0 a_9557_390.t0 VDD.t19 ppolyf_u r_width=1u r_length=1u
X191 a_1997_n1144.t0 a_2277_n1446.t1 VDD.t30 ppolyf_u r_width=1u r_length=1u
X192 a_3957_n794.t1 a_3957_n1796.t0 VDD.t38 ppolyf_u r_width=1u r_length=1u
X193 a_8997_692.t1 H.t0 VDD.t10 ppolyf_u r_width=1u r_length=1u
X194 G.t10 a_1717_n794.t1 VDD.t33 ppolyf_u r_width=1u r_length=1u
X195 a_5637_n1446.t0 a_6477_n2098.t1 VDD.t3 ppolyf_u r_width=1u r_length=1u
X196 a_3397_692.t0 a_3117_390.t0 VDD.t29 ppolyf_u r_width=1u r_length=1u
X197 a_1717_n1144.t1 a_1717_n1446.t1 VDD.t33 ppolyf_u r_width=1u r_length=1u
X198 a_8997_n1796.t0 a_7877_n1446.t0 VDD.t10 ppolyf_u r_width=1u r_length=1u
X199 a_2277_1694.t1 a_2277_692.t1 VDD.t37 ppolyf_u r_width=1u r_length=1u
X200 a_6197_n794.t0 a_6197_n1796.t1 VDD.t18 ppolyf_u r_width=1u r_length=1u
X201 a_8437_692.t0 D.t0 VDD.t28 ppolyf_u r_width=1u r_length=1u
X202 a_5917_n1796.t1 a_5637_n2098.t1 VDD.t8 ppolyf_u r_width=1u r_length=1u
X203 a_8997_n794.t1 a_8717_n2098.t1 VDD.t19 ppolyf_u r_width=1u r_length=1u
R0 a_7877_692.t0 a_7877_692.t1 13.3663
R1 a_7597_390.t0 a_7597_390.t1 13.3663
R2 VDD.n353 VDD.t35 9.01689
R3 VDD.n273 VDD.t12 9.01689
R4 VDD.n140 VDD.t8 9.01689
R5 VDD.n990 VDD.t26 9.01689
R6 VDD.n852 VDD.t0 9.01689
R7 VDD.n345 VDD.t19 8.19722
R8 VDD.n261 VDD.t4 8.19722
R9 VDD.n126 VDD.t1 8.19722
R10 VDD.n978 VDD.t27 8.19722
R11 VDD.n838 VDD.t33 8.19722
R12 VDD.n736 VDD.t44 7.09079
R13 VDD.n82 VDD.t51 7.09079
R14 VDD.n536 VDD.t43 7.0013
R15 VDD.n451 VDD.t54 7.0013
R16 VDD.n507 VDD.t49 7.00054
R17 VDD.n405 VDD.t46 7.00054
R18 VDD.n514 VDD.t48 7.00019
R19 VDD.n418 VDD.t47 7.00019
R20 VDD.n521 VDD.t24 6.99979
R21 VDD.n428 VDD.t40 6.99979
R22 VDD.n529 VDD.t23 6.99941
R23 VDD.n441 VDD.t41 6.99941
R24 VDD.n543 VDD.t42 6.99677
R25 VDD.n458 VDD.t55 6.99677
R26 VDD.n729 VDD.t45 6.99412
R27 VDD.n86 VDD.t50 6.99412
R28 VDD.n753 VDD.t16 6.92009
R29 VDD.n73 VDD.t15 6.92009
R30 VDD.n745 VDD.t17 6.91844
R31 VDD.n77 VDD.t14 6.91844
R32 VDD.n50 VDD.t56 6.84254
R33 VDD.n1 VDD.t53 6.84254
R34 VDD.n50 VDD.t57 6.4095
R35 VDD.n1 VDD.t52 6.4095
R36 VDD.n364 VDD.t22 6.14804
R37 VDD.n285 VDD.t25 6.14804
R38 VDD.n163 VDD.t9 6.14804
R39 VDD.n1013 VDD.t31 6.14804
R40 VDD.n872 VDD.t30 6.14804
R41 VDD.n333 VDD.t2 5.32837
R42 VDD.n243 VDD.t21 5.32837
R43 VDD.n105 VDD.t6 5.32837
R44 VDD.n956 VDD.t29 5.32837
R45 VDD.n818 VDD.t36 5.32837
R46 VDD.n297 VDD.t28 3.27919
R47 VDD.n184 VDD.t3 3.27919
R48 VDD.n1034 VDD.t32 3.27919
R49 VDD.n890 VDD.t34 3.27919
R50 VDD.n401 VDD.n400 3.1505
R51 VDD.n464 VDD.n463 3.1505
R52 VDD.n462 VDD.n461 3.1505
R53 VDD.n460 VDD.n459 3.1505
R54 VDD.n457 VDD.n456 3.1505
R55 VDD.n455 VDD.n454 3.1505
R56 VDD.n453 VDD.n452 3.1505
R57 VDD.n450 VDD.n449 3.1505
R58 VDD.n447 VDD.n446 3.1505
R59 VDD.n444 VDD.n443 3.1505
R60 VDD.n440 VDD.n439 3.1505
R61 VDD.n437 VDD.n436 3.1505
R62 VDD.n434 VDD.n433 3.1505
R63 VDD.n431 VDD.n430 3.1505
R64 VDD.n427 VDD.n426 3.1505
R65 VDD.n424 VDD.n423 3.1505
R66 VDD.n421 VDD.n420 3.1505
R67 VDD.n417 VDD.n416 3.1505
R68 VDD.n414 VDD.n413 3.1505
R69 VDD.n411 VDD.n410 3.1505
R70 VDD.n408 VDD.n407 3.1505
R71 VDD.n404 VDD.n403 3.1505
R72 VDD.n549 VDD.n548 3.1505
R73 VDD.n547 VDD.n546 3.1505
R74 VDD.n545 VDD.n544 3.1505
R75 VDD.n542 VDD.n541 3.1505
R76 VDD.n540 VDD.n539 3.1505
R77 VDD.n538 VDD.n537 3.1505
R78 VDD.n535 VDD.n534 3.1505
R79 VDD.n533 VDD.n532 3.1505
R80 VDD.n531 VDD.n530 3.1505
R81 VDD.n529 VDD.n528 3.1505
R82 VDD.n527 VDD.n526 3.1505
R83 VDD.n525 VDD.n524 3.1505
R84 VDD.n523 VDD.n522 3.1505
R85 VDD.n520 VDD.n519 3.1505
R86 VDD.n518 VDD.n517 3.1505
R87 VDD.n516 VDD.n515 3.1505
R88 VDD.n513 VDD.n512 3.1505
R89 VDD.n511 VDD.n510 3.1505
R90 VDD.n503 VDD.n502 3.1505
R91 VDD.n501 VDD.n500 3.1505
R92 VDD.n499 VDD.n498 3.1505
R93 VDD.n497 VDD.n496 3.1505
R94 VDD.n361 VDD.n360 3.1505
R95 VDD.n357 VDD.n356 3.1505
R96 VDD.n353 VDD.n352 3.1505
R97 VDD.n349 VDD.n348 3.1505
R98 VDD.n345 VDD.n344 3.1505
R99 VDD.n341 VDD.n340 3.1505
R100 VDD.n337 VDD.n336 3.1505
R101 VDD.n333 VDD.n332 3.1505
R102 VDD.n329 VDD.n328 3.1505
R103 VDD.n325 VDD.n324 3.1505
R104 VDD.n321 VDD.n320 3.1505
R105 VDD.n317 VDD.n316 3.1505
R106 VDD.n313 VDD.n312 3.1505
R107 VDD.n309 VDD.n308 3.1505
R108 VDD.n305 VDD.n304 3.1505
R109 VDD.n301 VDD.n300 3.1505
R110 VDD.n297 VDD.n296 3.1505
R111 VDD.n293 VDD.n292 3.1505
R112 VDD.n289 VDD.n288 3.1505
R113 VDD.n285 VDD.n284 3.1505
R114 VDD.n281 VDD.n280 3.1505
R115 VDD.n277 VDD.n276 3.1505
R116 VDD.n273 VDD.n270 3.1505
R117 VDD.n267 VDD.n264 3.1505
R118 VDD.n261 VDD.n258 3.1505
R119 VDD.n255 VDD.n252 3.1505
R120 VDD.n249 VDD.n246 3.1505
R121 VDD.n243 VDD.n240 3.1505
R122 VDD.n237 VDD.n234 3.1505
R123 VDD.n231 VDD.n228 3.1505
R124 VDD.n225 VDD.n222 3.1505
R125 VDD.n219 VDD.n216 3.1505
R126 VDD.n213 VDD.n210 3.1505
R127 VDD.n204 VDD.n203 3.1505
R128 VDD.n207 VDD.n204 3.1505
R129 VDD.n196 VDD.n193 3.1505
R130 VDD.n190 VDD.n187 3.1505
R131 VDD.n181 VDD.n180 3.1505
R132 VDD.n184 VDD.n181 3.1505
R133 VDD.n175 VDD.n172 3.1505
R134 VDD.n169 VDD.n166 3.1505
R135 VDD.n160 VDD.n159 3.1505
R136 VDD.n163 VDD.n160 3.1505
R137 VDD.n151 VDD.n150 3.1505
R138 VDD.n154 VDD.n151 3.1505
R139 VDD.n144 VDD.n143 3.1505
R140 VDD.n147 VDD.n144 3.1505
R141 VDD.n137 VDD.n136 3.1505
R142 VDD.n140 VDD.n137 3.1505
R143 VDD.n130 VDD.n129 3.1505
R144 VDD.n133 VDD.n130 3.1505
R145 VDD.n126 VDD.n123 3.1505
R146 VDD.n117 VDD.n116 3.1505
R147 VDD.n120 VDD.n117 3.1505
R148 VDD.n109 VDD.n108 3.1505
R149 VDD.n112 VDD.n109 3.1505
R150 VDD.n102 VDD.n101 3.1505
R151 VDD.n105 VDD.n102 3.1505
R152 VDD.n95 VDD.n94 3.1505
R153 VDD.n98 VDD.n95 3.1505
R154 VDD.n1077 VDD.n1076 3.1505
R155 VDD.n1076 VDD.n1075 3.1505
R156 VDD.n1079 VDD.n1078 3.1505
R157 VDD.n1082 VDD.n1079 3.1505
R158 VDD.n1066 VDD.n1065 3.1505
R159 VDD.n1069 VDD.n1066 3.1505
R160 VDD.n1059 VDD.n1058 3.1505
R161 VDD.n1062 VDD.n1059 3.1505
R162 VDD.n1052 VDD.n1051 3.1505
R163 VDD.n1055 VDD.n1052 3.1505
R164 VDD.n1046 VDD.n1043 3.1505
R165 VDD.n1040 VDD.n1037 3.1505
R166 VDD.n1031 VDD.n1030 3.1505
R167 VDD.n1034 VDD.n1031 3.1505
R168 VDD.n1026 VDD.n1023 3.1505
R169 VDD.n1017 VDD.n1016 3.1505
R170 VDD.n1020 VDD.n1017 3.1505
R171 VDD.n1010 VDD.n1009 3.1505
R172 VDD.n1013 VDD.n1010 3.1505
R173 VDD.n1003 VDD.n1002 3.1505
R174 VDD.n1006 VDD.n1003 3.1505
R175 VDD.n996 VDD.n993 3.1505
R176 VDD.n990 VDD.n987 3.1505
R177 VDD.n984 VDD.n981 3.1505
R178 VDD.n975 VDD.n974 3.1505
R179 VDD.n978 VDD.n975 3.1505
R180 VDD.n968 VDD.n965 3.1505
R181 VDD.n962 VDD.n959 3.1505
R182 VDD.n956 VDD.n953 3.1505
R183 VDD.n947 VDD.n946 3.1505
R184 VDD.n950 VDD.n947 3.1505
R185 VDD.n932 VDD.n929 3.1505
R186 VDD.n926 VDD.n923 3.1505
R187 VDD.n920 VDD.n917 3.1505
R188 VDD.n914 VDD.n911 3.1505
R189 VDD.n908 VDD.n905 3.1505
R190 VDD.n902 VDD.n899 3.1505
R191 VDD.n896 VDD.n893 3.1505
R192 VDD.n890 VDD.n887 3.1505
R193 VDD.n884 VDD.n881 3.1505
R194 VDD.n878 VDD.n875 3.1505
R195 VDD.n872 VDD.n869 3.1505
R196 VDD.n863 VDD.n862 3.1505
R197 VDD.n866 VDD.n863 3.1505
R198 VDD.n858 VDD.n855 3.1505
R199 VDD.n849 VDD.n848 3.1505
R200 VDD.n852 VDD.n849 3.1505
R201 VDD.n842 VDD.n841 3.1505
R202 VDD.n845 VDD.n842 3.1505
R203 VDD.n835 VDD.n834 3.1505
R204 VDD.n838 VDD.n835 3.1505
R205 VDD.n828 VDD.n827 3.1505
R206 VDD.n831 VDD.n828 3.1505
R207 VDD.n824 VDD.n821 3.1505
R208 VDD.n818 VDD.n815 3.1505
R209 VDD.n812 VDD.n809 3.1505
R210 VDD.n806 VDD.n805 3.1505
R211 VDD.n802 VDD.n801 3.1505
R212 VDD.n798 VDD.n797 3.1505
R213 VDD.n794 VDD.n793 3.1505
R214 VDD.n789 VDD.n788 3.1505
R215 VDD.n785 VDD.n784 3.1505
R216 VDD.n781 VDD.n780 3.1505
R217 VDD.n777 VDD.n776 3.1505
R218 VDD.n373 VDD.n93 3.1505
R219 VDD.n93 VDD.n92 3.1505
R220 VDD.n779 VDD.n778 3.1505
R221 VDD.n778 VDD.n777 3.1505
R222 VDD.n783 VDD.n782 3.1505
R223 VDD.n782 VDD.n781 3.1505
R224 VDD.n787 VDD.n786 3.1505
R225 VDD.n786 VDD.n785 3.1505
R226 VDD.n791 VDD.n790 3.1505
R227 VDD.n790 VDD.n789 3.1505
R228 VDD.n796 VDD.n795 3.1505
R229 VDD.n795 VDD.n794 3.1505
R230 VDD.n800 VDD.n799 3.1505
R231 VDD.n799 VDD.n798 3.1505
R232 VDD.n804 VDD.n803 3.1505
R233 VDD.n803 VDD.n802 3.1505
R234 VDD.n808 VDD.n807 3.1505
R235 VDD.n807 VDD.n806 3.1505
R236 VDD.n814 VDD.n813 3.1505
R237 VDD.n813 VDD.n812 3.1505
R238 VDD.n820 VDD.n819 3.1505
R239 VDD.n819 VDD.n818 3.1505
R240 VDD.n826 VDD.n825 3.1505
R241 VDD.n825 VDD.n824 3.1505
R242 VDD.n833 VDD.n832 3.1505
R243 VDD.n832 VDD.n831 3.1505
R244 VDD.n840 VDD.n839 3.1505
R245 VDD.n839 VDD.n838 3.1505
R246 VDD.n847 VDD.n846 3.1505
R247 VDD.n846 VDD.n845 3.1505
R248 VDD.n854 VDD.n853 3.1505
R249 VDD.n853 VDD.n852 3.1505
R250 VDD.n860 VDD.n859 3.1505
R251 VDD.n859 VDD.n858 3.1505
R252 VDD.n868 VDD.n867 3.1505
R253 VDD.n867 VDD.n866 3.1505
R254 VDD.n874 VDD.n873 3.1505
R255 VDD.n873 VDD.n872 3.1505
R256 VDD.n880 VDD.n879 3.1505
R257 VDD.n879 VDD.n878 3.1505
R258 VDD.n886 VDD.n885 3.1505
R259 VDD.n885 VDD.n884 3.1505
R260 VDD.n892 VDD.n891 3.1505
R261 VDD.n891 VDD.n890 3.1505
R262 VDD.n898 VDD.n897 3.1505
R263 VDD.n897 VDD.n896 3.1505
R264 VDD.n904 VDD.n903 3.1505
R265 VDD.n903 VDD.n902 3.1505
R266 VDD.n910 VDD.n909 3.1505
R267 VDD.n909 VDD.n908 3.1505
R268 VDD.n916 VDD.n915 3.1505
R269 VDD.n915 VDD.n914 3.1505
R270 VDD.n922 VDD.n921 3.1505
R271 VDD.n921 VDD.n920 3.1505
R272 VDD.n928 VDD.n927 3.1505
R273 VDD.n927 VDD.n926 3.1505
R274 VDD.n934 VDD.n933 3.1505
R275 VDD.n933 VDD.n932 3.1505
R276 VDD.n952 VDD.n951 3.1505
R277 VDD.n951 VDD.n950 3.1505
R278 VDD.n958 VDD.n957 3.1505
R279 VDD.n957 VDD.n956 3.1505
R280 VDD.n964 VDD.n963 3.1505
R281 VDD.n963 VDD.n962 3.1505
R282 VDD.n970 VDD.n969 3.1505
R283 VDD.n969 VDD.n968 3.1505
R284 VDD.n980 VDD.n979 3.1505
R285 VDD.n979 VDD.n978 3.1505
R286 VDD.n986 VDD.n985 3.1505
R287 VDD.n985 VDD.n984 3.1505
R288 VDD.n992 VDD.n991 3.1505
R289 VDD.n991 VDD.n990 3.1505
R290 VDD.n998 VDD.n997 3.1505
R291 VDD.n997 VDD.n996 3.1505
R292 VDD.n1008 VDD.n1007 3.1505
R293 VDD.n1007 VDD.n1006 3.1505
R294 VDD.n1015 VDD.n1014 3.1505
R295 VDD.n1014 VDD.n1013 3.1505
R296 VDD.n1022 VDD.n1021 3.1505
R297 VDD.n1021 VDD.n1020 3.1505
R298 VDD.n1028 VDD.n1027 3.1505
R299 VDD.n1027 VDD.n1026 3.1505
R300 VDD.n1036 VDD.n1035 3.1505
R301 VDD.n1035 VDD.n1034 3.1505
R302 VDD.n1042 VDD.n1041 3.1505
R303 VDD.n1041 VDD.n1040 3.1505
R304 VDD.n1048 VDD.n1047 3.1505
R305 VDD.n1047 VDD.n1046 3.1505
R306 VDD.n1057 VDD.n1056 3.1505
R307 VDD.n1056 VDD.n1055 3.1505
R308 VDD.n1064 VDD.n1063 3.1505
R309 VDD.n1063 VDD.n1062 3.1505
R310 VDD.n1071 VDD.n1070 3.1505
R311 VDD.n1070 VDD.n1069 3.1505
R312 VDD.n1084 VDD.n1083 3.1505
R313 VDD.n1083 VDD.n1082 3.1505
R314 VDD.n1074 VDD.n0 3.1505
R315 VDD.n1075 VDD.n1074 3.1505
R316 VDD.n100 VDD.n99 3.1505
R317 VDD.n99 VDD.n98 3.1505
R318 VDD.n107 VDD.n106 3.1505
R319 VDD.n106 VDD.n105 3.1505
R320 VDD.n114 VDD.n113 3.1505
R321 VDD.n113 VDD.n112 3.1505
R322 VDD.n122 VDD.n121 3.1505
R323 VDD.n121 VDD.n120 3.1505
R324 VDD.n128 VDD.n127 3.1505
R325 VDD.n127 VDD.n126 3.1505
R326 VDD.n135 VDD.n134 3.1505
R327 VDD.n134 VDD.n133 3.1505
R328 VDD.n142 VDD.n141 3.1505
R329 VDD.n141 VDD.n140 3.1505
R330 VDD.n149 VDD.n148 3.1505
R331 VDD.n148 VDD.n147 3.1505
R332 VDD.n156 VDD.n155 3.1505
R333 VDD.n155 VDD.n154 3.1505
R334 VDD.n165 VDD.n164 3.1505
R335 VDD.n164 VDD.n163 3.1505
R336 VDD.n171 VDD.n170 3.1505
R337 VDD.n170 VDD.n169 3.1505
R338 VDD.n177 VDD.n176 3.1505
R339 VDD.n176 VDD.n175 3.1505
R340 VDD.n186 VDD.n185 3.1505
R341 VDD.n185 VDD.n184 3.1505
R342 VDD.n192 VDD.n191 3.1505
R343 VDD.n191 VDD.n190 3.1505
R344 VDD.n198 VDD.n197 3.1505
R345 VDD.n197 VDD.n196 3.1505
R346 VDD.n209 VDD.n208 3.1505
R347 VDD.n208 VDD.n207 3.1505
R348 VDD.n215 VDD.n214 3.1505
R349 VDD.n214 VDD.n213 3.1505
R350 VDD.n221 VDD.n220 3.1505
R351 VDD.n220 VDD.n219 3.1505
R352 VDD.n227 VDD.n226 3.1505
R353 VDD.n226 VDD.n225 3.1505
R354 VDD.n233 VDD.n232 3.1505
R355 VDD.n232 VDD.n231 3.1505
R356 VDD.n239 VDD.n238 3.1505
R357 VDD.n238 VDD.n237 3.1505
R358 VDD.n245 VDD.n244 3.1505
R359 VDD.n244 VDD.n243 3.1505
R360 VDD.n251 VDD.n250 3.1505
R361 VDD.n250 VDD.n249 3.1505
R362 VDD.n257 VDD.n256 3.1505
R363 VDD.n256 VDD.n255 3.1505
R364 VDD.n263 VDD.n262 3.1505
R365 VDD.n262 VDD.n261 3.1505
R366 VDD.n269 VDD.n268 3.1505
R367 VDD.n268 VDD.n267 3.1505
R368 VDD.n275 VDD.n274 3.1505
R369 VDD.n274 VDD.n273 3.1505
R370 VDD.n279 VDD.n278 3.1505
R371 VDD.n278 VDD.n277 3.1505
R372 VDD.n283 VDD.n282 3.1505
R373 VDD.n282 VDD.n281 3.1505
R374 VDD.n287 VDD.n286 3.1505
R375 VDD.n286 VDD.n285 3.1505
R376 VDD.n291 VDD.n290 3.1505
R377 VDD.n290 VDD.n289 3.1505
R378 VDD.n295 VDD.n294 3.1505
R379 VDD.n294 VDD.n293 3.1505
R380 VDD.n299 VDD.n298 3.1505
R381 VDD.n298 VDD.n297 3.1505
R382 VDD.n303 VDD.n302 3.1505
R383 VDD.n302 VDD.n301 3.1505
R384 VDD.n307 VDD.n306 3.1505
R385 VDD.n306 VDD.n305 3.1505
R386 VDD.n311 VDD.n310 3.1505
R387 VDD.n310 VDD.n309 3.1505
R388 VDD.n315 VDD.n314 3.1505
R389 VDD.n314 VDD.n313 3.1505
R390 VDD.n319 VDD.n318 3.1505
R391 VDD.n318 VDD.n317 3.1505
R392 VDD.n323 VDD.n322 3.1505
R393 VDD.n322 VDD.n321 3.1505
R394 VDD.n327 VDD.n326 3.1505
R395 VDD.n326 VDD.n325 3.1505
R396 VDD.n331 VDD.n330 3.1505
R397 VDD.n330 VDD.n329 3.1505
R398 VDD.n335 VDD.n334 3.1505
R399 VDD.n334 VDD.n333 3.1505
R400 VDD.n339 VDD.n338 3.1505
R401 VDD.n338 VDD.n337 3.1505
R402 VDD.n343 VDD.n342 3.1505
R403 VDD.n342 VDD.n341 3.1505
R404 VDD.n347 VDD.n346 3.1505
R405 VDD.n346 VDD.n345 3.1505
R406 VDD.n351 VDD.n350 3.1505
R407 VDD.n350 VDD.n349 3.1505
R408 VDD.n355 VDD.n354 3.1505
R409 VDD.n354 VDD.n353 3.1505
R410 VDD.n359 VDD.n358 3.1505
R411 VDD.n358 VDD.n357 3.1505
R412 VDD.n363 VDD.n362 3.1505
R413 VDD.n362 VDD.n361 3.1505
R414 VDD.n366 VDD.n365 3.1505
R415 VDD.n365 VDD.n364 3.1505
R416 VDD.n369 VDD.n368 3.1505
R417 VDD.n368 VDD.n367 3.1505
R418 VDD.n372 VDD.n371 3.1505
R419 VDD.n371 VDD.n370 3.1505
R420 VDD.n399 VDD.n398 3.1505
R421 VDD.n49 VDD.n48 3.1505
R422 VDD.n772 VDD.n771 3.1505
R423 VDD.n769 VDD.n768 3.1505
R424 VDD.n767 VDD.n766 3.1505
R425 VDD.n764 VDD.n763 3.1505
R426 VDD.n762 VDD.n761 3.1505
R427 VDD.n759 VDD.n758 3.1505
R428 VDD.n757 VDD.n756 3.1505
R429 VDD.n755 VDD.n754 3.1505
R430 VDD.n752 VDD.n751 3.1505
R431 VDD.n750 VDD.n749 3.1505
R432 VDD.n747 VDD.n746 3.1505
R433 VDD.n744 VDD.n743 3.1505
R434 VDD.n742 VDD.n741 3.1505
R435 VDD.n740 VDD.n739 3.1505
R436 VDD.n738 VDD.n737 3.1505
R437 VDD.n735 VDD.n734 3.1505
R438 VDD.n733 VDD.n732 3.1505
R439 VDD.n731 VDD.n730 3.1505
R440 VDD.n728 VDD.n727 3.1505
R441 VDD.n726 VDD.n725 3.1505
R442 VDD.n774 VDD.n773 3.1505
R443 VDD.n91 VDD.n90 3.1505
R444 VDD.n46 VDD.n5 3.1505
R445 VDD.n466 VDD.n465 3.1505
R446 VDD.n551 VDD.n550 3.1505
R447 VDD.n555 VDD.n553 3.1505
R448 VDD.n558 VDD.n556 3.1505
R449 VDD.n561 VDD.n559 3.1505
R450 VDD.n564 VDD.n562 3.1505
R451 VDD.n567 VDD.n565 3.1505
R452 VDD.n570 VDD.n568 3.1505
R453 VDD.n573 VDD.n571 3.1505
R454 VDD.n576 VDD.n574 3.1505
R455 VDD.n579 VDD.n577 3.1505
R456 VDD.n582 VDD.n580 3.1505
R457 VDD.n585 VDD.n583 3.1505
R458 VDD.n588 VDD.n586 3.1505
R459 VDD.n591 VDD.n589 3.1505
R460 VDD.n594 VDD.n592 3.1505
R461 VDD.n597 VDD.n595 3.1505
R462 VDD.n600 VDD.n598 3.1505
R463 VDD.n603 VDD.n601 3.1505
R464 VDD.n606 VDD.n604 3.1505
R465 VDD.n609 VDD.n607 3.1505
R466 VDD.n612 VDD.n610 3.1505
R467 VDD.n615 VDD.n613 3.1505
R468 VDD.n618 VDD.n616 3.1505
R469 VDD.n621 VDD.n619 3.1505
R470 VDD.n624 VDD.n622 3.1505
R471 VDD.n627 VDD.n625 3.1505
R472 VDD.n630 VDD.n628 3.1505
R473 VDD.n273 VDD.n272 3.1505
R474 VDD.n267 VDD.n266 3.1505
R475 VDD.n261 VDD.n260 3.1505
R476 VDD.n255 VDD.n254 3.1505
R477 VDD.n249 VDD.n248 3.1505
R478 VDD.n243 VDD.n242 3.1505
R479 VDD.n237 VDD.n236 3.1505
R480 VDD.n231 VDD.n230 3.1505
R481 VDD.n225 VDD.n224 3.1505
R482 VDD.n219 VDD.n218 3.1505
R483 VDD.n213 VDD.n212 3.1505
R484 VDD.n207 VDD.n206 3.1505
R485 VDD.n196 VDD.n195 3.1505
R486 VDD.n190 VDD.n189 3.1505
R487 VDD.n184 VDD.n183 3.1505
R488 VDD.n175 VDD.n174 3.1505
R489 VDD.n169 VDD.n168 3.1505
R490 VDD.n163 VDD.n162 3.1505
R491 VDD.n154 VDD.n153 3.1505
R492 VDD.n147 VDD.n146 3.1505
R493 VDD.n140 VDD.n139 3.1505
R494 VDD.n133 VDD.n132 3.1505
R495 VDD.n126 VDD.n125 3.1505
R496 VDD.n120 VDD.n119 3.1505
R497 VDD.n112 VDD.n111 3.1505
R498 VDD.n105 VDD.n104 3.1505
R499 VDD.n98 VDD.n97 3.1505
R500 VDD.n1075 VDD.n1073 3.1505
R501 VDD.n1082 VDD.n1081 3.1505
R502 VDD.n1069 VDD.n1068 3.1505
R503 VDD.n1062 VDD.n1061 3.1505
R504 VDD.n1055 VDD.n1054 3.1505
R505 VDD.n1046 VDD.n1045 3.1505
R506 VDD.n1040 VDD.n1039 3.1505
R507 VDD.n1034 VDD.n1033 3.1505
R508 VDD.n1026 VDD.n1025 3.1505
R509 VDD.n1020 VDD.n1019 3.1505
R510 VDD.n1013 VDD.n1012 3.1505
R511 VDD.n1006 VDD.n1005 3.1505
R512 VDD.n996 VDD.n995 3.1505
R513 VDD.n990 VDD.n989 3.1505
R514 VDD.n984 VDD.n983 3.1505
R515 VDD.n978 VDD.n977 3.1505
R516 VDD.n968 VDD.n967 3.1505
R517 VDD.n962 VDD.n961 3.1505
R518 VDD.n956 VDD.n955 3.1505
R519 VDD.n950 VDD.n949 3.1505
R520 VDD.n932 VDD.n931 3.1505
R521 VDD.n926 VDD.n925 3.1505
R522 VDD.n920 VDD.n919 3.1505
R523 VDD.n914 VDD.n913 3.1505
R524 VDD.n908 VDD.n907 3.1505
R525 VDD.n902 VDD.n901 3.1505
R526 VDD.n896 VDD.n895 3.1505
R527 VDD.n890 VDD.n889 3.1505
R528 VDD.n884 VDD.n883 3.1505
R529 VDD.n878 VDD.n877 3.1505
R530 VDD.n872 VDD.n871 3.1505
R531 VDD.n866 VDD.n865 3.1505
R532 VDD.n858 VDD.n857 3.1505
R533 VDD.n852 VDD.n851 3.1505
R534 VDD.n845 VDD.n844 3.1505
R535 VDD.n838 VDD.n837 3.1505
R536 VDD.n831 VDD.n830 3.1505
R537 VDD.n824 VDD.n823 3.1505
R538 VDD.n818 VDD.n817 3.1505
R539 VDD.n812 VDD.n811 3.1505
R540 VDD.n700 VDD.n698 3.1505
R541 VDD.n703 VDD.n701 3.1505
R542 VDD.n706 VDD.n704 3.1505
R543 VDD.n709 VDD.n707 3.1505
R544 VDD.n712 VDD.n710 3.1505
R545 VDD.n715 VDD.n713 3.1505
R546 VDD.n718 VDD.n716 3.1505
R547 VDD.n721 VDD.n719 3.1505
R548 VDD.n555 VDD.n554 3.1505
R549 VDD.n558 VDD.n557 3.1505
R550 VDD.n561 VDD.n560 3.1505
R551 VDD.n564 VDD.n563 3.1505
R552 VDD.n567 VDD.n566 3.1505
R553 VDD.n570 VDD.n569 3.1505
R554 VDD.n573 VDD.n572 3.1505
R555 VDD.n576 VDD.n575 3.1505
R556 VDD.n579 VDD.n578 3.1505
R557 VDD.n582 VDD.n581 3.1505
R558 VDD.n585 VDD.n584 3.1505
R559 VDD.n588 VDD.n587 3.1505
R560 VDD.n591 VDD.n590 3.1505
R561 VDD.n594 VDD.n593 3.1505
R562 VDD.n597 VDD.n596 3.1505
R563 VDD.n600 VDD.n599 3.1505
R564 VDD.n603 VDD.n602 3.1505
R565 VDD.n606 VDD.n605 3.1505
R566 VDD.n609 VDD.n608 3.1505
R567 VDD.n612 VDD.n611 3.1505
R568 VDD.n615 VDD.n614 3.1505
R569 VDD.n618 VDD.n617 3.1505
R570 VDD.n621 VDD.n620 3.1505
R571 VDD.n624 VDD.n623 3.1505
R572 VDD.n627 VDD.n626 3.1505
R573 VDD.n630 VDD.n629 3.1505
R574 VDD.n273 VDD.n271 3.1505
R575 VDD.n267 VDD.n265 3.1505
R576 VDD.n261 VDD.n259 3.1505
R577 VDD.n255 VDD.n253 3.1505
R578 VDD.n249 VDD.n247 3.1505
R579 VDD.n243 VDD.n241 3.1505
R580 VDD.n237 VDD.n235 3.1505
R581 VDD.n231 VDD.n229 3.1505
R582 VDD.n225 VDD.n223 3.1505
R583 VDD.n219 VDD.n217 3.1505
R584 VDD.n213 VDD.n211 3.1505
R585 VDD.n207 VDD.n205 3.1505
R586 VDD.n196 VDD.n194 3.1505
R587 VDD.n190 VDD.n188 3.1505
R588 VDD.n184 VDD.n182 3.1505
R589 VDD.n175 VDD.n173 3.1505
R590 VDD.n169 VDD.n167 3.1505
R591 VDD.n163 VDD.n161 3.1505
R592 VDD.n154 VDD.n152 3.1505
R593 VDD.n147 VDD.n145 3.1505
R594 VDD.n140 VDD.n138 3.1505
R595 VDD.n133 VDD.n131 3.1505
R596 VDD.n126 VDD.n124 3.1505
R597 VDD.n120 VDD.n118 3.1505
R598 VDD.n112 VDD.n110 3.1505
R599 VDD.n105 VDD.n103 3.1505
R600 VDD.n98 VDD.n96 3.1505
R601 VDD.n1075 VDD.n1072 3.1505
R602 VDD.n1082 VDD.n1080 3.1505
R603 VDD.n1069 VDD.n1067 3.1505
R604 VDD.n1062 VDD.n1060 3.1505
R605 VDD.n1055 VDD.n1053 3.1505
R606 VDD.n1046 VDD.n1044 3.1505
R607 VDD.n1040 VDD.n1038 3.1505
R608 VDD.n1034 VDD.n1032 3.1505
R609 VDD.n1026 VDD.n1024 3.1505
R610 VDD.n1020 VDD.n1018 3.1505
R611 VDD.n1013 VDD.n1011 3.1505
R612 VDD.n1006 VDD.n1004 3.1505
R613 VDD.n996 VDD.n994 3.1505
R614 VDD.n990 VDD.n988 3.1505
R615 VDD.n984 VDD.n982 3.1505
R616 VDD.n978 VDD.n976 3.1505
R617 VDD.n968 VDD.n966 3.1505
R618 VDD.n962 VDD.n960 3.1505
R619 VDD.n956 VDD.n954 3.1505
R620 VDD.n950 VDD.n948 3.1505
R621 VDD.n932 VDD.n930 3.1505
R622 VDD.n926 VDD.n924 3.1505
R623 VDD.n920 VDD.n918 3.1505
R624 VDD.n914 VDD.n912 3.1505
R625 VDD.n908 VDD.n906 3.1505
R626 VDD.n902 VDD.n900 3.1505
R627 VDD.n896 VDD.n894 3.1505
R628 VDD.n890 VDD.n888 3.1505
R629 VDD.n884 VDD.n882 3.1505
R630 VDD.n878 VDD.n876 3.1505
R631 VDD.n872 VDD.n870 3.1505
R632 VDD.n866 VDD.n864 3.1505
R633 VDD.n858 VDD.n856 3.1505
R634 VDD.n852 VDD.n850 3.1505
R635 VDD.n845 VDD.n843 3.1505
R636 VDD.n838 VDD.n836 3.1505
R637 VDD.n831 VDD.n829 3.1505
R638 VDD.n824 VDD.n822 3.1505
R639 VDD.n818 VDD.n816 3.1505
R640 VDD.n812 VDD.n810 3.1505
R641 VDD.n700 VDD.n699 3.1505
R642 VDD.n703 VDD.n702 3.1505
R643 VDD.n706 VDD.n705 3.1505
R644 VDD.n709 VDD.n708 3.1505
R645 VDD.n712 VDD.n711 3.1505
R646 VDD.n715 VDD.n714 3.1505
R647 VDD.n718 VDD.n717 3.1505
R648 VDD.n721 VDD.n720 3.1505
R649 VDD.n321 VDD.t10 2.45952
R650 VDD.n225 VDD.t18 2.45952
R651 VDD.n1082 VDD.t20 2.45952
R652 VDD.n926 VDD.t7 2.45952
R653 VDD.n802 VDD.t5 2.45952
R654 VDD.n407 VDD.n406 2.39402
R655 VDD.n410 VDD.n409 2.39402
R656 VDD.n413 VDD.n412 2.39402
R657 VDD.n416 VDD.n415 2.39402
R658 VDD.n420 VDD.n419 2.39402
R659 VDD.n423 VDD.n422 2.39402
R660 VDD.n426 VDD.n425 2.39402
R661 VDD.n430 VDD.n429 2.39402
R662 VDD.n433 VDD.n432 2.39402
R663 VDD.n436 VDD.n435 2.39402
R664 VDD.n439 VDD.n438 2.39402
R665 VDD.n443 VDD.n442 2.39402
R666 VDD.n446 VDD.n445 2.39402
R667 VDD.n449 VDD.n448 2.39402
R668 VDD.n396 VDD.n392 1.95449
R669 VDD.n396 VDD.n393 1.95449
R670 VDD.n396 VDD.n394 1.95449
R671 VDD.n396 VDD.n395 1.95449
R672 VDD.n379 VDD.n377 1.73593
R673 VDD.n4 VDD.n2 1.73593
R674 VDD.n381 VDD.n380 1.73541
R675 VDD.n379 VDD.n378 1.73541
R676 VDD.n4 VDD.n3 1.73541
R677 VDD.n35 VDD.n33 1.73527
R678 VDD.n32 VDD.n30 1.73527
R679 VDD.n29 VDD.n27 1.73527
R680 VDD.n26 VDD.n24 1.73527
R681 VDD.n23 VDD.n21 1.73527
R682 VDD.n20 VDD.n18 1.73527
R683 VDD.n17 VDD.n15 1.73527
R684 VDD.n14 VDD.n12 1.73527
R685 VDD.n11 VDD.n9 1.73527
R686 VDD.n8 VDD.n6 1.73527
R687 VDD.n771 VDD.n770 1.73527
R688 VDD.n766 VDD.n765 1.73527
R689 VDD.n761 VDD.n760 1.73527
R690 VDD.n32 VDD.n31 1.73527
R691 VDD.n29 VDD.n28 1.73527
R692 VDD.n26 VDD.n25 1.73527
R693 VDD.n23 VDD.n22 1.73527
R694 VDD.n20 VDD.n19 1.73527
R695 VDD.n17 VDD.n16 1.73527
R696 VDD.n14 VDD.n13 1.73527
R697 VDD.n11 VDD.n10 1.73527
R698 VDD.n8 VDD.n7 1.73527
R699 VDD.n35 VDD.n34 1.73527
R700 VDD.n403 VDD.n402 1.41722
R701 VDD.n376 VDD.n374 1.377
R702 VDD.n48 VDD.n47 1.377
R703 VDD.n376 VDD.n375 1.37653
R704 VDD.n398 VDD.n397 1.37653
R705 VDD.n38 VDD.n36 1.32491
R706 VDD.n38 VDD.n37 1.32491
R707 VDD.n396 VDD.n391 1.15696
R708 VDD.n396 VDD.n390 0.914272
R709 VDD.n46 VDD.n38 0.914044
R710 VDD.n396 VDD.n376 0.888554
R711 VDD.n397 VDD.n396 0.888554
R712 VDD.n47 VDD.n46 0.888554
R713 VDD.n396 VDD.n389 0.709103
R714 VDD.n396 VDD.n388 0.709103
R715 VDD.n396 VDD.n387 0.709103
R716 VDD.n396 VDD.n386 0.709103
R717 VDD.n396 VDD.n385 0.709103
R718 VDD.n396 VDD.n384 0.709103
R719 VDD.n396 VDD.n383 0.709103
R720 VDD.n396 VDD.n382 0.709103
R721 VDD.n396 VDD.n381 0.709103
R722 VDD.n396 VDD.n379 0.709103
R723 VDD.n46 VDD.n4 0.709102
R724 VDD.n46 VDD.n45 0.708865
R725 VDD.n46 VDD.n44 0.708865
R726 VDD.n46 VDD.n43 0.708865
R727 VDD.n46 VDD.n42 0.708865
R728 VDD.n46 VDD.n41 0.708865
R729 VDD.n46 VDD.n40 0.708865
R730 VDD.n46 VDD.n39 0.708865
R731 VDD.n46 VDD.n35 0.708865
R732 VDD.n46 VDD.n32 0.708865
R733 VDD.n46 VDD.n29 0.708865
R734 VDD.n46 VDD.n26 0.708865
R735 VDD.n46 VDD.n23 0.708865
R736 VDD.n46 VDD.n20 0.708865
R737 VDD.n46 VDD.n17 0.708865
R738 VDD.n46 VDD.n14 0.708865
R739 VDD.n46 VDD.n11 0.708865
R740 VDD.n46 VDD.n8 0.708865
R741 VDD.n309 VDD.t11 0.410336
R742 VDD.n207 VDD.t39 0.410336
R743 VDD.n1055 VDD.t38 0.410336
R744 VDD.n908 VDD.t37 0.410336
R745 VDD.n789 VDD.t13 0.410336
R746 VDD.n58 VDD.n50 0.329196
R747 VDD.n792 VDD.n1 0.329196
R748 VDD.n64 VDD.n63 0.220012
R749 VDD.n774 VDD.n772 0.215622
R750 VDD.n772 VDD.n769 0.215622
R751 VDD.n769 VDD.n767 0.215622
R752 VDD.n767 VDD.n764 0.215622
R753 VDD.n764 VDD.n762 0.215622
R754 VDD.n762 VDD.n759 0.215622
R755 VDD.n759 VDD.n757 0.215622
R756 VDD.n757 VDD.n755 0.215622
R757 VDD.n752 VDD.n750 0.215622
R758 VDD.n744 VDD.n742 0.215622
R759 VDD.n742 VDD.n740 0.215622
R760 VDD.n740 VDD.n738 0.215622
R761 VDD.n735 VDD.n733 0.215622
R762 VDD.n733 VDD.n731 0.215622
R763 VDD.n728 VDD.n726 0.215622
R764 VDD.n726 VDD.n724 0.215622
R765 VDD.n724 VDD.n723 0.215622
R766 VDD.n91 VDD.n89 0.215622
R767 VDD.n89 VDD.n88 0.215622
R768 VDD.n88 VDD.n87 0.215622
R769 VDD.n85 VDD.n84 0.215622
R770 VDD.n84 VDD.n83 0.215622
R771 VDD.n81 VDD.n80 0.215622
R772 VDD.n80 VDD.n79 0.215622
R773 VDD.n79 VDD.n78 0.215622
R774 VDD.n76 VDD.n75 0.215622
R775 VDD.n75 VDD.n74 0.215622
R776 VDD.n72 VDD.n71 0.215622
R777 VDD.n71 VDD.n70 0.215622
R778 VDD.n70 VDD.n69 0.215622
R779 VDD.n69 VDD.n68 0.215622
R780 VDD.n68 VDD.n67 0.215622
R781 VDD.n67 VDD.n66 0.215622
R782 VDD.n66 VDD.n65 0.215622
R783 VDD.n65 VDD.n64 0.215622
R784 VDD.n723 VDD.n722 0.211232
R785 VDD.n722 VDD.n91 0.211232
R786 VDD.n750 VDD.n748 0.191476
R787 VDD.n747 VDD.n745 0.187085
R788 VDD.n77 VDD.n76 0.187085
R789 VDD.n83 VDD.n82 0.165134
R790 VDD.n736 VDD.n735 0.162939
R791 VDD.n504 VDD.n503 0.14675
R792 VDD.n399 VDD.n373 0.14675
R793 VDD.n775 VDD.n774 0.136598
R794 VDD.n731 VDD.n729 0.134402
R795 VDD.n86 VDD.n85 0.132207
R796 VDD.n755 VDD.n753 0.130012
R797 VDD.n73 VDD.n72 0.130012
R798 VDD.n552 VDD.n466 0.12875
R799 VDD.n552 VDD.n551 0.12875
R800 VDD.n503 VDD.n501 0.11075
R801 VDD.n501 VDD.n499 0.11075
R802 VDD.n499 VDD.n497 0.11075
R803 VDD.n497 VDD.n495 0.11075
R804 VDD.n495 VDD.n494 0.11075
R805 VDD.n494 VDD.n493 0.11075
R806 VDD.n493 VDD.n492 0.11075
R807 VDD.n492 VDD.n491 0.11075
R808 VDD.n491 VDD.n490 0.11075
R809 VDD.n490 VDD.n489 0.11075
R810 VDD.n489 VDD.n488 0.11075
R811 VDD.n488 VDD.n487 0.11075
R812 VDD.n487 VDD.n486 0.11075
R813 VDD.n486 VDD.n485 0.11075
R814 VDD.n485 VDD.n484 0.11075
R815 VDD.n484 VDD.n483 0.11075
R816 VDD.n483 VDD.n482 0.11075
R817 VDD.n482 VDD.n481 0.11075
R818 VDD.n481 VDD.n480 0.11075
R819 VDD.n480 VDD.n479 0.11075
R820 VDD.n479 VDD.n478 0.11075
R821 VDD.n478 VDD.n477 0.11075
R822 VDD.n477 VDD.n476 0.11075
R823 VDD.n476 VDD.n475 0.11075
R824 VDD.n475 VDD.n474 0.11075
R825 VDD.n474 VDD.n473 0.11075
R826 VDD.n473 VDD.n472 0.11075
R827 VDD.n472 VDD.n471 0.11075
R828 VDD.n471 VDD.n470 0.11075
R829 VDD.n470 VDD.n469 0.11075
R830 VDD.n469 VDD.n468 0.11075
R831 VDD.n468 VDD.n467 0.11075
R832 VDD.n200 VDD.n199 0.11075
R833 VDD.n201 VDD.n200 0.11075
R834 VDD.n202 VDD.n201 0.11075
R835 VDD.n203 VDD.n202 0.11075
R836 VDD.n179 VDD.n178 0.11075
R837 VDD.n180 VDD.n179 0.11075
R838 VDD.n158 VDD.n157 0.11075
R839 VDD.n159 VDD.n158 0.11075
R840 VDD.n116 VDD.n115 0.11075
R841 VDD.n1051 VDD.n1050 0.11075
R842 VDD.n1050 VDD.n1049 0.11075
R843 VDD.n1030 VDD.n1029 0.11075
R844 VDD.n1002 VDD.n1001 0.11075
R845 VDD.n1001 VDD.n1000 0.11075
R846 VDD.n1000 VDD.n999 0.11075
R847 VDD.n974 VDD.n973 0.11075
R848 VDD.n973 VDD.n972 0.11075
R849 VDD.n972 VDD.n971 0.11075
R850 VDD.n946 VDD.n945 0.11075
R851 VDD.n945 VDD.n944 0.11075
R852 VDD.n944 VDD.n943 0.11075
R853 VDD.n943 VDD.n942 0.11075
R854 VDD.n942 VDD.n941 0.11075
R855 VDD.n941 VDD.n940 0.11075
R856 VDD.n940 VDD.n939 0.11075
R857 VDD.n939 VDD.n938 0.11075
R858 VDD.n938 VDD.n937 0.11075
R859 VDD.n937 VDD.n936 0.11075
R860 VDD.n936 VDD.n935 0.11075
R861 VDD.n862 VDD.n861 0.11075
R862 VDD.n52 VDD.n51 0.11075
R863 VDD.n53 VDD.n52 0.11075
R864 VDD.n54 VDD.n53 0.11075
R865 VDD.n55 VDD.n54 0.11075
R866 VDD.n56 VDD.n55 0.11075
R867 VDD.n57 VDD.n56 0.11075
R868 VDD.n60 VDD.n59 0.11075
R869 VDD.n61 VDD.n60 0.11075
R870 VDD.n62 VDD.n61 0.11075
R871 VDD.n549 VDD.n547 0.11075
R872 VDD.n547 VDD.n545 0.11075
R873 VDD.n542 VDD.n540 0.11075
R874 VDD.n540 VDD.n538 0.11075
R875 VDD.n535 VDD.n533 0.11075
R876 VDD.n533 VDD.n531 0.11075
R877 VDD.n531 VDD.n529 0.11075
R878 VDD.n529 VDD.n527 0.11075
R879 VDD.n527 VDD.n525 0.11075
R880 VDD.n525 VDD.n523 0.11075
R881 VDD.n520 VDD.n518 0.11075
R882 VDD.n518 VDD.n516 0.11075
R883 VDD.n513 VDD.n511 0.11075
R884 VDD.n511 VDD.n509 0.11075
R885 VDD.n509 VDD.n508 0.11075
R886 VDD.n506 VDD.n505 0.11075
R887 VDD.n404 VDD.n401 0.11075
R888 VDD.n411 VDD.n408 0.11075
R889 VDD.n414 VDD.n411 0.11075
R890 VDD.n417 VDD.n414 0.11075
R891 VDD.n424 VDD.n421 0.11075
R892 VDD.n427 VDD.n424 0.11075
R893 VDD.n434 VDD.n431 0.11075
R894 VDD.n437 VDD.n434 0.11075
R895 VDD.n440 VDD.n437 0.11075
R896 VDD.n447 VDD.n444 0.11075
R897 VDD.n450 VDD.n447 0.11075
R898 VDD.n455 VDD.n453 0.11075
R899 VDD.n457 VDD.n455 0.11075
R900 VDD.n462 VDD.n460 0.11075
R901 VDD.n464 VDD.n462 0.11075
R902 VDD.n373 VDD.n372 0.11075
R903 VDD.n372 VDD.n369 0.11075
R904 VDD.n369 VDD.n366 0.11075
R905 VDD.n366 VDD.n363 0.11075
R906 VDD.n363 VDD.n359 0.11075
R907 VDD.n359 VDD.n355 0.11075
R908 VDD.n355 VDD.n351 0.11075
R909 VDD.n351 VDD.n347 0.11075
R910 VDD.n347 VDD.n343 0.11075
R911 VDD.n343 VDD.n339 0.11075
R912 VDD.n339 VDD.n335 0.11075
R913 VDD.n335 VDD.n331 0.11075
R914 VDD.n331 VDD.n327 0.11075
R915 VDD.n327 VDD.n323 0.11075
R916 VDD.n323 VDD.n319 0.11075
R917 VDD.n319 VDD.n315 0.11075
R918 VDD.n315 VDD.n311 0.11075
R919 VDD.n311 VDD.n307 0.11075
R920 VDD.n307 VDD.n303 0.11075
R921 VDD.n303 VDD.n299 0.11075
R922 VDD.n299 VDD.n295 0.11075
R923 VDD.n295 VDD.n291 0.11075
R924 VDD.n291 VDD.n287 0.11075
R925 VDD.n287 VDD.n283 0.11075
R926 VDD.n283 VDD.n279 0.11075
R927 VDD.n279 VDD.n275 0.11075
R928 VDD.n275 VDD.n269 0.11075
R929 VDD.n269 VDD.n263 0.11075
R930 VDD.n263 VDD.n257 0.11075
R931 VDD.n257 VDD.n251 0.11075
R932 VDD.n251 VDD.n245 0.11075
R933 VDD.n245 VDD.n239 0.11075
R934 VDD.n239 VDD.n233 0.11075
R935 VDD.n233 VDD.n227 0.11075
R936 VDD.n227 VDD.n221 0.11075
R937 VDD.n221 VDD.n215 0.11075
R938 VDD.n215 VDD.n209 0.11075
R939 VDD.n209 VDD.n198 0.11075
R940 VDD.n198 VDD.n192 0.11075
R941 VDD.n192 VDD.n186 0.11075
R942 VDD.n186 VDD.n177 0.11075
R943 VDD.n177 VDD.n171 0.11075
R944 VDD.n171 VDD.n165 0.11075
R945 VDD.n165 VDD.n156 0.11075
R946 VDD.n156 VDD.n149 0.11075
R947 VDD.n149 VDD.n142 0.11075
R948 VDD.n142 VDD.n135 0.11075
R949 VDD.n135 VDD.n128 0.11075
R950 VDD.n128 VDD.n122 0.11075
R951 VDD.n122 VDD.n114 0.11075
R952 VDD.n114 VDD.n107 0.11075
R953 VDD.n107 VDD.n100 0.11075
R954 VDD.n100 VDD.n0 0.11075
R955 VDD.n1084 VDD.n1071 0.11075
R956 VDD.n1071 VDD.n1064 0.11075
R957 VDD.n1064 VDD.n1057 0.11075
R958 VDD.n1057 VDD.n1048 0.11075
R959 VDD.n1048 VDD.n1042 0.11075
R960 VDD.n1042 VDD.n1036 0.11075
R961 VDD.n1036 VDD.n1028 0.11075
R962 VDD.n1028 VDD.n1022 0.11075
R963 VDD.n1022 VDD.n1015 0.11075
R964 VDD.n1015 VDD.n1008 0.11075
R965 VDD.n1008 VDD.n998 0.11075
R966 VDD.n998 VDD.n992 0.11075
R967 VDD.n992 VDD.n986 0.11075
R968 VDD.n986 VDD.n980 0.11075
R969 VDD.n980 VDD.n970 0.11075
R970 VDD.n970 VDD.n964 0.11075
R971 VDD.n964 VDD.n958 0.11075
R972 VDD.n958 VDD.n952 0.11075
R973 VDD.n952 VDD.n934 0.11075
R974 VDD.n934 VDD.n928 0.11075
R975 VDD.n928 VDD.n922 0.11075
R976 VDD.n922 VDD.n916 0.11075
R977 VDD.n916 VDD.n910 0.11075
R978 VDD.n910 VDD.n904 0.11075
R979 VDD.n904 VDD.n898 0.11075
R980 VDD.n898 VDD.n892 0.11075
R981 VDD.n892 VDD.n886 0.11075
R982 VDD.n886 VDD.n880 0.11075
R983 VDD.n880 VDD.n874 0.11075
R984 VDD.n874 VDD.n868 0.11075
R985 VDD.n868 VDD.n860 0.11075
R986 VDD.n860 VDD.n854 0.11075
R987 VDD.n854 VDD.n847 0.11075
R988 VDD.n847 VDD.n840 0.11075
R989 VDD.n840 VDD.n833 0.11075
R990 VDD.n833 VDD.n826 0.11075
R991 VDD.n826 VDD.n820 0.11075
R992 VDD.n820 VDD.n814 0.11075
R993 VDD.n814 VDD.n808 0.11075
R994 VDD.n808 VDD.n804 0.11075
R995 VDD.n804 VDD.n800 0.11075
R996 VDD.n800 VDD.n796 0.11075
R997 VDD.n791 VDD.n787 0.11075
R998 VDD.n787 VDD.n783 0.11075
R999 VDD.n783 VDD.n779 0.11075
R1000 VDD.n444 VDD.n441 0.109625
R1001 VDD.n405 VDD.n404 0.104
R1002 VDD.n507 VDD.n506 0.102875
R1003 VDD.n58 VDD.n57 0.0995
R1004 VDD.n796 VDD.n792 0.0995
R1005 VDD.n779 VDD.n775 0.089375
R1006 VDD.n753 VDD.n752 0.0861098
R1007 VDD.n74 VDD.n73 0.0861098
R1008 VDD.n87 VDD.n86 0.0839146
R1009 VDD.n538 VDD.n536 0.08375
R1010 VDD.n516 VDD.n514 0.082625
R1011 VDD.n453 VDD.n451 0.082625
R1012 VDD.n729 VDD.n728 0.0817195
R1013 VDD.n421 VDD.n418 0.0815
R1014 VDD.n505 VDD.n504 0.07025
R1015 VDD.n401 VDD.n399 0.07025
R1016 VDD.n63 VDD.n62 0.0701402
R1017 VDD.n458 VDD.n457 0.069125
R1018 VDD.n543 VDD.n542 0.068
R1019 VDD.n551 VDD.n549 0.06575
R1020 VDD.n466 VDD.n464 0.06575
R1021 VDD.n428 VDD.n427 0.062375
R1022 VDD.n521 VDD.n520 0.06125
R1023 VDD VDD.n1077 0.05675
R1024 VDD VDD.n0 0.05675
R1025 VDD.n1078 VDD 0.0545
R1026 VDD VDD.n1084 0.0545
R1027 VDD.n738 VDD.n736 0.0531829
R1028 VDD.n82 VDD.n81 0.0509878
R1029 VDD.n523 VDD.n521 0.05
R1030 VDD.n431 VDD.n428 0.048875
R1031 VDD.n545 VDD.n543 0.04325
R1032 VDD.n460 VDD.n458 0.042125
R1033 VDD.n558 VDD.n555 0.0329265
R1034 VDD.n561 VDD.n558 0.0329265
R1035 VDD.n564 VDD.n561 0.0329265
R1036 VDD.n567 VDD.n564 0.0329265
R1037 VDD.n570 VDD.n567 0.0329265
R1038 VDD.n573 VDD.n570 0.0329265
R1039 VDD.n576 VDD.n573 0.0329265
R1040 VDD.n579 VDD.n576 0.0329265
R1041 VDD.n582 VDD.n579 0.0329265
R1042 VDD.n585 VDD.n582 0.0329265
R1043 VDD.n588 VDD.n585 0.0329265
R1044 VDD.n591 VDD.n588 0.0329265
R1045 VDD.n594 VDD.n591 0.0329265
R1046 VDD.n597 VDD.n594 0.0329265
R1047 VDD.n600 VDD.n597 0.0329265
R1048 VDD.n603 VDD.n600 0.0329265
R1049 VDD.n606 VDD.n603 0.0329265
R1050 VDD.n609 VDD.n606 0.0329265
R1051 VDD.n612 VDD.n609 0.0329265
R1052 VDD.n615 VDD.n612 0.0329265
R1053 VDD.n618 VDD.n615 0.0329265
R1054 VDD.n621 VDD.n618 0.0329265
R1055 VDD.n624 VDD.n621 0.0329265
R1056 VDD.n627 VDD.n624 0.0329265
R1057 VDD.n630 VDD.n627 0.0329265
R1058 VDD.n631 VDD.n630 0.0329265
R1059 VDD.n632 VDD.n631 0.0329265
R1060 VDD.n633 VDD.n632 0.0329265
R1061 VDD.n634 VDD.n633 0.0329265
R1062 VDD.n635 VDD.n634 0.0329265
R1063 VDD.n636 VDD.n635 0.0329265
R1064 VDD.n637 VDD.n636 0.0329265
R1065 VDD.n638 VDD.n637 0.0329265
R1066 VDD.n639 VDD.n638 0.0329265
R1067 VDD.n640 VDD.n639 0.0329265
R1068 VDD.n641 VDD.n640 0.0329265
R1069 VDD.n642 VDD.n641 0.0329265
R1070 VDD.n643 VDD.n642 0.0329265
R1071 VDD.n644 VDD.n643 0.0329265
R1072 VDD.n645 VDD.n644 0.0329265
R1073 VDD.n646 VDD.n645 0.0329265
R1074 VDD.n647 VDD.n646 0.0329265
R1075 VDD.n648 VDD.n647 0.0329265
R1076 VDD.n649 VDD.n648 0.0329265
R1077 VDD.n650 VDD.n649 0.0329265
R1078 VDD.n651 VDD.n650 0.0329265
R1079 VDD.n652 VDD.n651 0.0329265
R1080 VDD.n653 VDD.n652 0.0329265
R1081 VDD.n654 VDD.n653 0.0329265
R1082 VDD.n655 VDD.n654 0.0329265
R1083 VDD.n656 VDD.n655 0.0329265
R1084 VDD.n657 VDD.n656 0.0329265
R1085 VDD.n658 VDD.n657 0.0329265
R1086 VDD.n659 VDD.n658 0.0329265
R1087 VDD.n660 VDD.n659 0.0329265
R1088 VDD.n661 VDD.n660 0.0329265
R1089 VDD.n662 VDD.n661 0.0329265
R1090 VDD.n663 VDD.n662 0.0329265
R1091 VDD.n664 VDD.n663 0.0329265
R1092 VDD.n665 VDD.n664 0.0329265
R1093 VDD.n666 VDD.n665 0.0329265
R1094 VDD.n667 VDD.n666 0.0329265
R1095 VDD.n669 VDD.n668 0.0329265
R1096 VDD.n670 VDD.n669 0.0329265
R1097 VDD.n671 VDD.n670 0.0329265
R1098 VDD.n672 VDD.n671 0.0329265
R1099 VDD.n673 VDD.n672 0.0329265
R1100 VDD.n674 VDD.n673 0.0329265
R1101 VDD.n675 VDD.n674 0.0329265
R1102 VDD.n676 VDD.n675 0.0329265
R1103 VDD.n677 VDD.n676 0.0329265
R1104 VDD.n678 VDD.n677 0.0329265
R1105 VDD.n679 VDD.n678 0.0329265
R1106 VDD.n680 VDD.n679 0.0329265
R1107 VDD.n681 VDD.n680 0.0329265
R1108 VDD.n682 VDD.n681 0.0329265
R1109 VDD.n683 VDD.n682 0.0329265
R1110 VDD.n684 VDD.n683 0.0329265
R1111 VDD.n685 VDD.n684 0.0329265
R1112 VDD.n686 VDD.n685 0.0329265
R1113 VDD.n687 VDD.n686 0.0329265
R1114 VDD.n688 VDD.n687 0.0329265
R1115 VDD.n689 VDD.n688 0.0329265
R1116 VDD.n690 VDD.n689 0.0329265
R1117 VDD.n691 VDD.n690 0.0329265
R1118 VDD.n692 VDD.n691 0.0329265
R1119 VDD.n693 VDD.n692 0.0329265
R1120 VDD.n694 VDD.n693 0.0329265
R1121 VDD.n695 VDD.n694 0.0329265
R1122 VDD.n696 VDD.n695 0.0329265
R1123 VDD.n697 VDD.n696 0.0329265
R1124 VDD.n700 VDD.n697 0.0329265
R1125 VDD.n703 VDD.n700 0.0329265
R1126 VDD.n706 VDD.n703 0.0329265
R1127 VDD.n709 VDD.n706 0.0329265
R1128 VDD.n712 VDD.n709 0.0329265
R1129 VDD.n715 VDD.n712 0.0329265
R1130 VDD.n718 VDD.n715 0.0329265
R1131 VDD.n721 VDD.n718 0.0329265
R1132 VDD.n418 VDD.n417 0.02975
R1133 VDD.n745 VDD.n744 0.0290366
R1134 VDD.n78 VDD.n77 0.0290366
R1135 VDD.n514 VDD.n513 0.028625
R1136 VDD.n451 VDD.n450 0.028625
R1137 VDD.n536 VDD.n535 0.0275
R1138 VDD.n748 VDD.n747 0.0246463
R1139 VDD.n668 VDD 0.023
R1140 VDD.n775 VDD.n49 0.021875
R1141 VDD.n722 VDD.n721 0.0196912
R1142 VDD.n59 VDD.n58 0.01175
R1143 VDD.n792 VDD.n791 0.01175
R1144 VDD VDD.n667 0.0104265
R1145 VDD.n508 VDD.n507 0.008375
R1146 VDD.n408 VDD.n405 0.00725
R1147 VDD.n555 VDD.n552 0.00579412
R1148 VDD.n441 VDD.n440 0.001625
R1149 a_2277_692.t0 a_2277_692.t1 9.02698
R1150 a_2277_390.t0 a_2277_390.t1 16.5556
R1151 a_1437_n1796.t0 a_1437_n1796.t1 12.7444
R1152 a_2837_n794.t0 a_2837_n794.t1 13.3663
R1153 C.n0 C.t2 14.2685
R1154 C.n2 C.t1 14.2681
R1155 C.n0 C.t0 10.016
R1156 C.n2 C.t3 10.0155
R1157 C.n3 C 4.01446
R1158 C C.n1 2.05447
R1159 C.n1 C.n0 0.501554
R1160 C.n3 C.n2 0.501256
R1161 C.n1 C 0.00595455
R1162 C C.n3 0.00595455
R1163 a_1997_1042.t0 a_1997_1042.t1 13.3663
R1164 G.n2 G.t3 8.07794
R1165 G.n10 G.t0 8.04282
R1166 G.n17 G.t11 6.5735
R1167 G.n8 G.t10 6.5725
R1168 G.n11 G.t9 5.27447
R1169 G.n3 G.t6 5.27433
R1170 G.n2 G.t7 5.07258
R1171 G.n10 G.t8 5.07252
R1172 G G.n17 3.34772
R1173 G G.n8 3.34772
R1174 G.n16 G.t5 3.25137
R1175 G.n0 G.t2 3.22368
R1176 G.n7 G.t1 3.2166
R1177 G.n13 G.t4 3.18852
R1178 G.n12 G.n9 2.35569
R1179 G.n14 G.n12 2.27388
R1180 G.n5 G.n4 2.27388
R1181 G.n14 G.n13 1.56636
R1182 G.n13 G.n9 1.56434
R1183 G.n1 G.n0 1.56406
R1184 G.n16 G.n15 1.08603
R1185 G.n7 G.n6 1.08567
R1186 G.n12 G.n11 0.835821
R1187 G.n4 G.n3 0.835821
R1188 G.n8 G.n7 0.457759
R1189 G.n17 G.n16 0.45775
R1190 G.n3 G.n2 0.197719
R1191 G.n11 G.n10 0.197719
R1192 G.n15 G.n9 0.0647857
R1193 G.n15 G.n14 0.0647857
R1194 G.n6 G.n1 0.0647857
R1195 G.n6 G.n5 0.0647857
R1196 a_3957_1344.t0 a_3957_1344.t1 15.1072
R1197 a_3957_1042.t0 a_3957_1042.t1 15.1112
R1198 a_7317_692.t0 a_7317_692.t1 13.3663
R1199 a_5917_1694.t0 a_5917_1694.t1 12.7437
R1200 E.n5 E.t7 7.96203
R1201 E.n2 E.t6 7.96203
R1202 E.n3 E.t2 6.95733
R1203 E.n0 E.t3 6.95733
R1204 E.n4 E.t1 6.42124
R1205 E.n1 E.t4 6.42124
R1206 E.n3 E.t0 6.4095
R1207 E.n0 E.t5 6.4095
R1208 E.n2 E.n1 2.56058
R1209 E.n5 E.n4 2.55977
R1210 E E.n5 0.838955
R1211 E E.n2 0.838955
R1212 E.n4 E.n3 0.381128
R1213 E.n1 E.n0 0.381128
R1214 a_4517_n794.t0 a_4517_n794.t1 11.2748
R1215 a_4237_n2098.t0 a_4237_n2098.t1 12.2092
R1216 a_5917_1344.t0 a_5917_1344.t1 12.1738
R1217 a_5917_1042.t0 a_5917_1042.t1 11.2391
R1218 a_3957_n1796.t0 a_3957_n1796.t1 13.318
R1219 a_2557_n2098.t0 a_2557_n2098.t1 15.6157
R1220 a_6757_692.t0 a_6757_692.t1 9.02706
R1221 a_6757_390.t0 a_6757_390.t1 16.5556
R1222 a_7597_n1144.t0 a_7597_n1144.t1 13.3663
R1223 a_6477_n2098.t0 a_6477_n2098.t1 14.7079
R1224 a_1157_390.n1 a_1157_390.t0 8.50661
R1225 a_1157_390.n0 a_1157_390.t3 6.84437
R1226 a_1157_390.t1 a_1157_390.n1 5.39199
R1227 a_1157_390.n0 a_1157_390.t2 3.14625
R1228 a_1157_390.n1 a_1157_390.n0 2.04585
R1229 a_8437_n1446.t0 a_8437_n1446.t1 15.1072
R1230 a_6197_n2098.t0 a_6197_n2098.t1 18.2801
R1231 a_4237_n1144.t0 a_4237_n1144.t1 13.3663
R1232 a_4517_n1446.t0 a_4517_n1446.t1 16.7065
R1233 a_1157_n492.n0 a_1157_n492.t3 8.4719
R1234 a_1157_n492.n1 a_1157_n492.t2 6.84402
R1235 a_1157_n492.n0 a_1157_n492.t1 5.39309
R1236 a_1157_n492.t0 a_1157_n492.n1 3.11188
R1237 a_1157_n492.n1 a_1157_n492.n0 2.04473
R1238 a_3957_n492.t0 a_3957_n492.t1 18.9537
R1239 a_3957_n794.t0 a_3957_n794.t1 14.6446
R1240 a_8157_n1446.t0 a_8157_n1446.t1 8.9401
R1241 a_8717_n2098.t0 a_8717_n2098.t1 12.2097
R1242 a_5637_n492.t0 a_5637_n492.t1 13.3663
R1243 a_5917_n794.t0 a_5917_n794.t1 13.8639
R1244 a_1717_1694.t0 a_1717_1694.t1 15.1072
R1245 a_1717_692.t0 a_1717_692.t1 15.1112
R1246 a_4517_1344.t0 a_4517_1344.t1 16.7065
R1247 a_4237_1042.t0 a_4237_1042.t1 13.3663
R1248 a_5357_692.t0 a_5357_692.t1 13.5463
R1249 a_5637_390.t0 a_5637_390.t1 13.3663
R1250 a_1157_n1446.t0 a_1157_n1446.t1 15.278
R1251 a_1997_n2098.n1 a_1997_n2098.t2 10.5961
R1252 a_1997_n2098.n2 a_1997_n2098.t3 10.5913
R1253 a_1997_n2098.n1 a_1997_n2098.t1 4.11102
R1254 a_1997_n2098.n2 a_1997_n2098.t5 4.11058
R1255 a_1997_n2098.t0 a_1997_n2098.n0 3.25271
R1256 a_1997_n2098.n0 a_1997_n2098.t4 3.25063
R1257 a_1997_n2098.n0 a_1997_n2098.n1 2.26965
R1258 a_1997_n2098.n0 a_1997_n2098.n2 2.25979
R1259 a_1717_n794.t0 a_1717_n794.t1 15.1112
R1260 a_1717_n1796.t0 a_1717_n1796.t1 15.1072
R1261 a_1717_n1144.t0 a_1717_n1144.t1 14.6445
R1262 a_3677_n1446.t0 a_3677_n1446.t1 8.9401
R1263 a_4517_n492.t0 a_4517_n492.t1 16.5391
R1264 a_1157_1344.t0 a_1157_1344.t1 15.3135
R1265 A A.t1 9.04183
R1266 A A.t0 9.04183
R1267 a_3677_1344.t0 a_3677_1344.t1 8.90503
R1268 a_3677_1042.t0 a_3677_1042.t1 9.02687
R1269 a_4517_692.t0 a_4517_692.t1 11.2396
R1270 a_4517_390.t0 a_4517_390.t1 16.5391
R1271 a_6757_n1796.t0 a_6757_n1796.t1 8.94028
R1272 a_5917_n1446.t0 a_5917_n1446.t1 12.2093
R1273 a_1997_1996.n2 a_1997_1996.t4 10.5962
R1274 a_1997_1996.n1 a_1997_1996.t5 10.5913
R1275 a_1997_1996.t0 a_1997_1996.n2 4.07589
R1276 a_1997_1996.n1 a_1997_1996.t2 4.07553
R1277 a_1997_1996.n0 a_1997_1996.t1 3.2869
R1278 a_1997_1996.n0 a_1997_1996.t3 3.2859
R1279 a_1997_1996.n2 a_1997_1996.n0 2.26982
R1280 a_1997_1996.n0 a_1997_1996.n1 2.25987
R1281 a_5637_1344.t0 a_5637_1344.t1 15.3126
R1282 a_5357_1042.t0 a_5357_1042.t1 13.5463
R1283 a_6757_n794.t0 a_6757_n794.t1 8.99186
R1284 a_3957_692.t0 a_3957_692.t1 14.6794
R1285 a_3957_390.t0 a_3957_390.t1 18.9537
R1286 a_1717_1996.t0 a_1717_1996.t1 18.2801
R1287 B.n1 B.t2 7.9449
R1288 B.n0 B.t0 7.9449
R1289 B.n1 B.t1 6.789
R1290 B.n0 B.t3 6.789
R1291 B B.n2 4.26687
R1292 B.n2 B.n1 2.25045
R1293 B.n3 B.n0 2.25045
R1294 B.n3 B 1.49544
R1295 B.n2 B 0.1892
R1296 B B.n3 0.1892
R1297 a_8997_n1796.t0 a_8997_n1796.t1 15.2785
R1298 a_3677_n492.t0 a_3677_n492.t1 12.746
R1299 a_3397_n794.t0 a_3397_n794.t1 13.3663
R1300 a_2277_n1796.t0 a_2277_n1796.t1 8.94028
R1301 a_3117_n492.t0 a_3117_n492.t1 13.3663
R1302 a_2277_1344.t0 a_2277_1344.t1 16.6921
R1303 a_5357_n794.t0 a_5357_n794.t1 13.5463
R1304 a_3957_1694.t0 a_3957_1694.t1 13.3172
R1305 a_3957_n1446.t0 a_3957_n1446.t1 15.1072
R1306 a_1717_n2098.t0 a_1717_n2098.t1 18.2801
R1307 a_2837_692.t0 a_2837_692.t1 13.3663
R1308 a_1437_1694.t0 a_1437_1694.t1 12.7436
R1309 a_6757_1344.t0 a_6757_1344.t1 16.6921
R1310 a_6477_1042.t0 a_6477_1042.t1 13.3663
R1311 a_5357_n1144.t0 a_5357_n1144.t1 13.5463
R1312 a_4517_n1796.t0 a_4517_n1796.t1 15.2785
R1313 a_2837_1996.t0 a_2837_1996.t1 13.3663
R1314 a_6197_n1446.t0 a_6197_n1446.t1 13.317
R1315 a_7037_n2098.t0 a_7037_n2098.t1 15.6157
R1316 a_8717_1042.t0 a_8717_1042.t1 13.3663
R1317 a_7877_n1446.t0 a_7877_n1446.t1 14.7052
R1318 a_2277_n492.t0 a_2277_n492.t1 16.5556
R1319 a_2277_n794.t0 a_2277_n794.t1 8.99186
R1320 a_8157_n492.t0 a_8157_n492.t1 12.746
R1321 a_9557_n2098.t0 a_9557_n2098.t1 13.3663
R1322 a_4797_n492.t0 a_4797_n492.t1 15.3136
R1323 a_3957_n1144.t0 a_3957_n1144.t1 15.1112
R1324 a_3677_n1144.t0 a_3677_n1144.t1 8.99184
R1325 a_6757_n492.t0 a_6757_n492.t1 16.5556
R1326 a_4517_1694.t0 a_4517_1694.t1 15.3118
R1327 a_7877_1344.t0 a_7877_1344.t1 14.6723
R1328 a_7597_1042.t0 a_7597_1042.t1 13.3663
R1329 a_8437_1042.t0 a_8437_1042.t1 15.1112
R1330 F.n0 F.t1 8.86329
R1331 F.n1 F.t0 8.86329
R1332 F.n0 F.t2 8.403
R1333 F.n1 F.t3 8.402
R1334 F F.n0 0.727136
R1335 F F.n1 0.727136
R1336 a_8157_n1144.t0 a_8157_n1144.t1 8.99184
R1337 a_2557_1996.t0 a_2557_1996.t1 15.6157
R1338 a_6757_1694.t0 a_6757_1694.t1 8.90405
R1339 a_8997_1694.t0 a_8997_1694.t1 15.3132
R1340 a_5077_n2098.t0 a_5077_n2098.t1 13.3663
R1341 a_5637_1996.t0 a_5637_1996.t1 13.3663
R1342 a_7597_n1796.t0 a_7597_n1796.t1 13.3663
R1343 a_7317_n2098.t0 a_7317_n2098.t1 13.3663
R1344 a_7597_n492.t0 a_7597_n492.t1 13.3663
R1345 a_7877_n794.t0 a_7877_n794.t1 13.3663
R1346 a_5077_n492.t0 a_5077_n492.t1 13.3663
R1347 a_8157_390.t0 a_8157_390.t1 12.746
R1348 a_9557_n492.t0 a_9557_n492.t1 13.3663
R1349 a_5917_n1796.t0 a_5917_n1796.t1 12.7436
R1350 a_7317_n794.t0 a_7317_n794.t1 13.3663
R1351 a_1717_1344.t0 a_1717_1344.t1 13.3171
R1352 a_8437_1344.t0 a_8437_1344.t1 15.1072
R1353 a_6197_1042.t0 a_6197_1042.t1 14.6793
R1354 a_5917_n1144.t0 a_5917_n1144.t1 11.2743
R1355 a_1717_n1446.t0 a_1717_n1446.t1 13.3151
R1356 H H.t0 10.2549
R1357 H H.t1 10.2549
R1358 a_8997_n794.t0 a_8997_n794.t1 11.2747
R1359 a_4237_1996.t0 a_4237_1996.t1 12.1742
R1360 a_6197_n1144.t0 a_6197_n1144.t1 14.6447
R1361 D.n0 D.t1 11.6419
R1362 D.n1 D.t2 11.6419
R1363 D.n1 D.t3 11.1324
R1364 D.n0 D.t0 11.1319
R1365 D D.n1 0.355623
R1366 D D.n0 0.355326
R1367 a_8437_n794.t0 a_8437_n794.t1 14.6447
R1368 a_6477_1996.t0 a_6477_1996.t1 14.6732
R1369 a_6197_1694.t0 a_6197_1694.t1 15.1072
R1370 a_6197_692.t0 a_6197_692.t1 15.1112
R1371 a_3397_1996.t0 a_3397_1996.t1 13.3663
R1372 a_3677_1694.t0 a_3677_1694.t1 13.8988
R1373 a_8717_1996.t0 a_8717_1996.t1 12.1749
R1374 a_8997_692.t0 a_8997_692.t1 11.2396
R1375 a_3117_1694.t0 a_3117_1694.t1 13.3663
R1376 a_5637_n1446.t0 a_5637_n1446.t1 15.278
R1377 a_5357_1694.t0 a_5357_1694.t1 13.5463
R1378 a_3677_n1796.t0 a_3677_n1796.t1 13.8645
R1379 a_5077_390.t0 a_5077_390.t1 13.3663
R1380 a_6197_1344.t0 a_6197_1344.t1 13.3162
R1381 a_8157_n1796.t0 a_8157_n1796.t1 13.865
R1382 a_4797_390.t0 a_4797_390.t1 15.3136
R1383 a_2277_1694.t0 a_2277_1694.t1 8.90503
R1384 a_8157_1344.t0 a_8157_1344.t1 8.90515
R1385 a_8157_1042.t0 a_8157_1042.t1 9.02687
R1386 a_9557_390.t0 a_9557_390.t1 13.3663
R1387 a_5357_n1796.t0 a_5357_n1796.t1 13.5463
R1388 a_6197_n794.t0 a_6197_n794.t1 15.1112
R1389 a_7877_n2098.t0 a_7877_n2098.t1 13.3663
R1390 a_3397_692.t0 a_3397_692.t1 13.3663
R1391 a_3677_390.t0 a_3677_390.t1 12.746
R1392 a_8437_n1144.t0 a_8437_n1144.t1 15.1112
R1393 a_8437_1694.t0 a_8437_1694.t1 13.3172
R1394 a_8437_692.t0 a_8437_692.t1 14.6794
R1395 a_5077_1996.t0 a_5077_1996.t1 13.3663
R1396 a_3117_390.t0 a_3117_390.t1 13.3663
R1397 a_7877_1996.t0 a_7877_1996.t1 13.3663
R1398 a_7597_1694.t0 a_7597_1694.t1 13.3663
R1399 a_7317_1996.t0 a_7317_1996.t1 13.3663
R1400 a_5917_692.t0 a_5917_692.t1 13.8981
R1401 a_3117_n1796.t0 a_3117_n1796.t1 13.3663
R1402 a_3397_n2098.t0 a_3397_n2098.t1 13.3663
R1403 a_9557_1996.t0 a_9557_1996.t1 13.3663
R1404 a_1717_1042.t0 a_1717_1042.t1 14.6793
R1405 a_2837_n2098.t0 a_2837_n2098.t1 13.3663
R1406 a_6477_n1144.t0 a_6477_n1144.t1 13.3663
R1407 a_8717_n1144.t0 a_8717_n1144.t1 13.3663
R1408 a_7037_1996.t0 a_7037_1996.t1 15.6157
R1409 a_6197_n1796.t0 a_6197_n1796.t1 15.1072
R1410 a_5637_n2098.t0 a_5637_n2098.t1 13.3663
R1411 a_8437_n1796.t0 a_8437_n1796.t1 13.318
R1412 a_6757_n1446.t0 a_6757_n1446.t1 16.6921
R1413 a_6197_1996.t0 a_6197_1996.t1 18.2801
R1414 a_8157_1694.t0 a_8157_1694.t1 13.8986
R1415 a_1997_n1144.t0 a_1997_n1144.t1 13.3663
R1416 a_2277_n1446.t0 a_2277_n1446.t1 16.6921
C0 E C 0.727f
C1 G A 0.181f
C2 F H 1.59f
C3 E G 1.12f
C4 VDD C 4.48f
C5 VDD G 4.52f
C6 E A 2.94f
C7 F B 0.215f
C8 VDD F 1.92f
C9 B H 0.0563f
C10 VDD H 2.55f
C11 F D 3.26f
C12 D H 0.201f
C13 VDD A 1.77f
C14 G C 1.78f
C15 VDD E 3.24f
C16 VDD B 4f
C17 D B 2.2f
C18 A C 2.87f
C19 VDD D 3.41f
C20 F VSUBS 1.68f
C21 H VSUBS 2.62f
C22 B VSUBS 2.45f
C23 C VSUBS 2.42f
C24 A VSUBS 5.44f
C25 D VSUBS 2.99f
C26 G VSUBS 2.25f
C27 E VSUBS 3.17f
C28 VDD VSUBS 0.154p
C29 D.t0 VSUBS 0.536f
C30 D.t1 VSUBS 0.574f
C31 D.n0 VSUBS 2.43f
C32 D.t2 VSUBS 0.574f
C33 D.t3 VSUBS 0.536f
C34 D.n1 VSUBS 2.43f
C35 H.t0 VSUBS 0.264f
C36 H.t1 VSUBS 0.264f
C37 F.t2 VSUBS 0.141f
C38 F.t1 VSUBS 0.173f
C39 F.n0 VSUBS 0.822f
C40 F.t3 VSUBS 0.141f
C41 F.t0 VSUBS 0.173f
C42 F.n1 VSUBS 0.822f
C43 B.t0 VSUBS 0.228f
C44 B.t3 VSUBS 0.189f
C45 B.n0 VSUBS 1.06f
C46 B.t2 VSUBS 0.228f
C47 B.t1 VSUBS 0.189f
C48 B.n1 VSUBS 1.06f
C49 B.n2 VSUBS 1.22f
C50 B.n3 VSUBS 0.604f
C51 a_1997_1996.n0 VSUBS 0.352f
C52 a_1997_1996.t4 VSUBS 0.161f
C53 a_1997_1996.t1 VSUBS 0.0425f
C54 a_1997_1996.t5 VSUBS 0.161f
C55 a_1997_1996.t2 VSUBS 0.0629f
C56 a_1997_1996.n1 VSUBS 0.613f
C57 a_1997_1996.t3 VSUBS 0.0425f
C58 a_1997_1996.n2 VSUBS 0.603f
C59 a_1997_1996.t0 VSUBS 0.0629f
C60 A.t0 VSUBS 0.433f
C61 A.t1 VSUBS 0.433f
C62 a_1997_n2098.n0 VSUBS 0.353f
C63 a_1997_n2098.t2 VSUBS 0.161f
C64 a_1997_n2098.t1 VSUBS 0.0628f
C65 a_1997_n2098.n1 VSUBS 0.603f
C66 a_1997_n2098.t3 VSUBS 0.161f
C67 a_1997_n2098.t5 VSUBS 0.0628f
C68 a_1997_n2098.n2 VSUBS 0.613f
C69 a_1997_n2098.t4 VSUBS 0.0423f
C70 a_1997_n2098.t0 VSUBS 0.0423f
C71 E.t4 VSUBS 0.122f
C72 E.t3 VSUBS 0.132f
C73 E.t5 VSUBS 0.121f
C74 E.n0 VSUBS 0.332f
C75 E.n1 VSUBS 0.463f
C76 E.t6 VSUBS 0.166f
C77 E.n2 VSUBS 0.817f
C78 E.t7 VSUBS 0.166f
C79 E.t1 VSUBS 0.122f
C80 E.t2 VSUBS 0.132f
C81 E.t0 VSUBS 0.121f
C82 E.n3 VSUBS 0.332f
C83 E.n4 VSUBS 0.463f
C84 E.n5 VSUBS 0.817f
C85 G.t1 VSUBS 0.0334f
C86 G.t2 VSUBS 0.0321f
C87 G.n0 VSUBS 0.079f
C88 G.n1 VSUBS 0.0203f
C89 G.t3 VSUBS 0.189f
C90 G.t7 VSUBS 0.0737f
C91 G.n2 VSUBS 0.49f
C92 G.t6 VSUBS 0.0727f
C93 G.n3 VSUBS 0.236f
C94 G.n4 VSUBS 0.134f
C95 G.n5 VSUBS 0.0179f
C96 G.n6 VSUBS 0.114f
C97 G.n7 VSUBS 0.128f
C98 G.t10 VSUBS 0.0488f
C99 G.n8 VSUBS 0.237f
C100 G.t5 VSUBS 0.0335f
C101 G.n9 VSUBS 0.0203f
C102 G.t0 VSUBS 0.189f
C103 G.t8 VSUBS 0.0737f
C104 G.n10 VSUBS 0.489f
C105 G.t9 VSUBS 0.0727f
C106 G.n11 VSUBS 0.236f
C107 G.n12 VSUBS 0.134f
C108 G.t4 VSUBS 0.032f
C109 G.n13 VSUBS 0.0791f
C110 G.n14 VSUBS 0.0179f
C111 G.n15 VSUBS 0.114f
C112 G.n16 VSUBS 0.128f
C113 G.t11 VSUBS 0.0488f
C114 G.n17 VSUBS 0.237f
C115 C.t2 VSUBS 0.64f
C116 C.t0 VSUBS 0.274f
C117 C.n0 VSUBS 1.83f
C118 C.n1 VSUBS 0.279f
C119 C.t3 VSUBS 0.274f
C120 C.t1 VSUBS 0.639f
C121 C.n2 VSUBS 1.83f
C122 C.n3 VSUBS 0.601f
C123 VDD.n0 VSUBS 0.00262f
C124 VDD.t52 VSUBS 0.00673f
C125 VDD.t53 VSUBS 0.00708f
C126 VDD.n1 VSUBS 0.0138f
C127 VDD.n2 VSUBS 0.00283f
C128 VDD.n3 VSUBS 0.00347f
C129 VDD.n5 VSUBS 0.00425f
C130 VDD.n6 VSUBS 0.00347f
C131 VDD.n7 VSUBS 0.00347f
C132 VDD.n9 VSUBS 0.00347f
C133 VDD.n10 VSUBS 0.00347f
C134 VDD.n12 VSUBS 0.00347f
C135 VDD.n13 VSUBS 0.00347f
C136 VDD.n15 VSUBS 0.00347f
C137 VDD.n16 VSUBS 0.00347f
C138 VDD.n18 VSUBS 0.00347f
C139 VDD.n19 VSUBS 0.00347f
C140 VDD.n21 VSUBS 0.00347f
C141 VDD.n22 VSUBS 0.00347f
C142 VDD.n24 VSUBS 0.00347f
C143 VDD.n25 VSUBS 0.00347f
C144 VDD.n27 VSUBS 0.00347f
C145 VDD.n28 VSUBS 0.00347f
C146 VDD.n30 VSUBS 0.00347f
C147 VDD.n31 VSUBS 0.00347f
C148 VDD.n33 VSUBS 0.00347f
C149 VDD.n34 VSUBS 0.00276f
C150 VDD.n36 VSUBS 0.00418f
C151 VDD.n37 VSUBS 0.00276f
C152 VDD.n46 VSUBS 0.3f
C153 VDD.n48 VSUBS 0.00425f
C154 VDD.n49 VSUBS 0.0111f
C155 VDD.t16 VSUBS 0.00739f
C156 VDD.t17 VSUBS 0.00739f
C157 VDD.t44 VSUBS 0.0075f
C158 VDD.t45 VSUBS 0.00743f
C159 VDD.t50 VSUBS 0.00743f
C160 VDD.t51 VSUBS 0.0075f
C161 VDD.t14 VSUBS 0.00739f
C162 VDD.t15 VSUBS 0.00739f
C163 VDD.t56 VSUBS 0.00708f
C164 VDD.t57 VSUBS 0.00673f
C165 VDD.n50 VSUBS 0.0138f
C166 VDD.n51 VSUBS 0.00347f
C167 VDD.n52 VSUBS 0.00347f
C168 VDD.n53 VSUBS 0.00347f
C169 VDD.n54 VSUBS 0.00347f
C170 VDD.n55 VSUBS 0.00347f
C171 VDD.n56 VSUBS 0.00347f
C172 VDD.n57 VSUBS 0.00329f
C173 VDD.n58 VSUBS 0.00558f
C174 VDD.n59 VSUBS 0.00191f
C175 VDD.n60 VSUBS 0.00347f
C176 VDD.n61 VSUBS 0.00347f
C177 VDD.n62 VSUBS 0.00287f
C178 VDD.n63 VSUBS 0.00259f
C179 VDD.n64 VSUBS 0.0018f
C180 VDD.n65 VSUBS 0.00178f
C181 VDD.n66 VSUBS 0.00178f
C182 VDD.n67 VSUBS 0.00178f
C183 VDD.n68 VSUBS 0.00178f
C184 VDD.n69 VSUBS 0.00178f
C185 VDD.n70 VSUBS 0.00178f
C186 VDD.n71 VSUBS 0.00178f
C187 VDD.n72 VSUBS 0.00142f
C188 VDD.n73 VSUBS 0.0145f
C189 VDD.n74 VSUBS 0.00124f
C190 VDD.n75 VSUBS -0.0192f
C191 VDD.n76 VSUBS -0.0177f
C192 VDD.n77 VSUBS 0.0145f
C193 VDD.n78 VSUBS 0.00101f
C194 VDD.n79 VSUBS 0.00178f
C195 VDD.n80 VSUBS 0.00178f
C196 VDD.n81 VSUBS 0.0011f
C197 VDD.n82 VSUBS 0.0117f
C198 VDD.n83 VSUBS 0.00157f
C199 VDD.n84 VSUBS 0.00178f
C200 VDD.n85 VSUBS 0.00143f
C201 VDD.n86 VSUBS 0.0131f
C202 VDD.n87 VSUBS 0.00123f
C203 VDD.n88 VSUBS 0.00178f
C204 VDD.n89 VSUBS 0.00178f
C205 VDD.n90 VSUBS 0.00418f
C206 VDD.n91 VSUBS 0.00176f
C207 VDD.t55 VSUBS 0.00743f
C208 VDD.t54 VSUBS 0.00743f
C209 VDD.t41 VSUBS 0.00743f
C210 VDD.t40 VSUBS 0.00743f
C211 VDD.t47 VSUBS 0.00743f
C212 VDD.t46 VSUBS 0.00743f
C213 VDD.n92 VSUBS 0.246f
C214 VDD.n93 VSUBS 0.00404f
C215 VDD.n94 VSUBS 0.00347f
C216 VDD.n95 VSUBS 0.00347f
C217 VDD.n96 VSUBS 0.00347f
C218 VDD.n97 VSUBS 0.00347f
C219 VDD.n98 VSUBS 0.184f
C220 VDD.n99 VSUBS 0.00347f
C221 VDD.n100 VSUBS 0.00347f
C222 VDD.t6 VSUBS 0.106f
C223 VDD.n101 VSUBS 0.00347f
C224 VDD.n102 VSUBS 0.00347f
C225 VDD.n103 VSUBS 0.00347f
C226 VDD.n104 VSUBS 0.00347f
C227 VDD.n105 VSUBS 0.134f
C228 VDD.n106 VSUBS 0.00347f
C229 VDD.n107 VSUBS 0.00347f
C230 VDD.n108 VSUBS 0.00347f
C231 VDD.n109 VSUBS 0.00347f
C232 VDD.n110 VSUBS 0.00347f
C233 VDD.n111 VSUBS 0.00347f
C234 VDD.n112 VSUBS 0.212f
C235 VDD.n113 VSUBS 0.00347f
C236 VDD.n114 VSUBS 0.00347f
C237 VDD.n115 VSUBS 0.00347f
C238 VDD.n116 VSUBS 0.00347f
C239 VDD.n117 VSUBS 0.00347f
C240 VDD.n118 VSUBS 0.00347f
C241 VDD.n119 VSUBS 0.00347f
C242 VDD.n120 VSUBS 0.168f
C243 VDD.n121 VSUBS 0.00347f
C244 VDD.n122 VSUBS 0.00347f
C245 VDD.t1 VSUBS 0.106f
C246 VDD.n123 VSUBS 0.00347f
C247 VDD.n124 VSUBS 0.00347f
C248 VDD.n125 VSUBS 0.00347f
C249 VDD.n126 VSUBS 0.149f
C250 VDD.n127 VSUBS 0.00347f
C251 VDD.n128 VSUBS 0.00347f
C252 VDD.n129 VSUBS 0.00347f
C253 VDD.n130 VSUBS 0.00347f
C254 VDD.n131 VSUBS 0.00347f
C255 VDD.n132 VSUBS 0.00347f
C256 VDD.n133 VSUBS 0.212f
C257 VDD.n134 VSUBS 0.00347f
C258 VDD.n135 VSUBS 0.00347f
C259 VDD.t8 VSUBS 0.106f
C260 VDD.n136 VSUBS 0.00347f
C261 VDD.n137 VSUBS 0.00347f
C262 VDD.n138 VSUBS 0.00347f
C263 VDD.n139 VSUBS 0.00347f
C264 VDD.n140 VSUBS 0.153f
C265 VDD.n141 VSUBS 0.00347f
C266 VDD.n142 VSUBS 0.00347f
C267 VDD.n143 VSUBS 0.00347f
C268 VDD.n144 VSUBS 0.00347f
C269 VDD.n145 VSUBS 0.00347f
C270 VDD.n146 VSUBS 0.00347f
C271 VDD.n147 VSUBS 0.164f
C272 VDD.n148 VSUBS 0.00347f
C273 VDD.n149 VSUBS 0.00347f
C274 VDD.n150 VSUBS 0.00347f
C275 VDD.n151 VSUBS 0.00347f
C276 VDD.n152 VSUBS 0.00347f
C277 VDD.n153 VSUBS 0.00347f
C278 VDD.n154 VSUBS 0.212f
C279 VDD.n155 VSUBS 0.00347f
C280 VDD.n156 VSUBS 0.00347f
C281 VDD.t9 VSUBS 0.106f
C282 VDD.n157 VSUBS 0.00347f
C283 VDD.n158 VSUBS 0.00347f
C284 VDD.n159 VSUBS 0.00347f
C285 VDD.n160 VSUBS 0.00347f
C286 VDD.n161 VSUBS 0.00347f
C287 VDD.n162 VSUBS 0.00347f
C288 VDD.n163 VSUBS 0.138f
C289 VDD.n164 VSUBS 0.00347f
C290 VDD.n165 VSUBS 0.00347f
C291 VDD.n166 VSUBS 0.00347f
C292 VDD.n167 VSUBS 0.00347f
C293 VDD.n168 VSUBS 0.00347f
C294 VDD.n169 VSUBS 0.179f
C295 VDD.n170 VSUBS 0.00347f
C296 VDD.n171 VSUBS 0.00347f
C297 VDD.n172 VSUBS 0.00347f
C298 VDD.n173 VSUBS 0.00347f
C299 VDD.n174 VSUBS 0.00347f
C300 VDD.n175 VSUBS 0.212f
C301 VDD.n176 VSUBS 0.00347f
C302 VDD.n177 VSUBS 0.00347f
C303 VDD.t3 VSUBS 0.106f
C304 VDD.n178 VSUBS 0.00347f
C305 VDD.n179 VSUBS 0.00347f
C306 VDD.n180 VSUBS 0.00347f
C307 VDD.n181 VSUBS 0.00347f
C308 VDD.n182 VSUBS 0.00347f
C309 VDD.n183 VSUBS 0.00347f
C310 VDD.n184 VSUBS 0.123f
C311 VDD.n185 VSUBS 0.00347f
C312 VDD.n186 VSUBS 0.00347f
C313 VDD.n187 VSUBS 0.00347f
C314 VDD.n188 VSUBS 0.00347f
C315 VDD.n189 VSUBS 0.00347f
C316 VDD.n190 VSUBS 0.194f
C317 VDD.n191 VSUBS 0.00347f
C318 VDD.n192 VSUBS 0.00347f
C319 VDD.n193 VSUBS 0.00347f
C320 VDD.n194 VSUBS 0.00347f
C321 VDD.n195 VSUBS 0.00347f
C322 VDD.n196 VSUBS 0.212f
C323 VDD.n197 VSUBS 0.00347f
C324 VDD.n198 VSUBS 0.00347f
C325 VDD.t39 VSUBS 0.106f
C326 VDD.n199 VSUBS 0.00347f
C327 VDD.n200 VSUBS 0.00347f
C328 VDD.n201 VSUBS 0.00347f
C329 VDD.n202 VSUBS 0.00347f
C330 VDD.n203 VSUBS 0.00347f
C331 VDD.n204 VSUBS 0.00347f
C332 VDD.n205 VSUBS 0.00347f
C333 VDD.n206 VSUBS 0.00347f
C334 VDD.n207 VSUBS 0.108f
C335 VDD.n208 VSUBS 0.00347f
C336 VDD.n209 VSUBS 0.00347f
C337 VDD.n210 VSUBS 0.00347f
C338 VDD.n211 VSUBS 0.00347f
C339 VDD.n212 VSUBS 0.00347f
C340 VDD.n213 VSUBS 0.21f
C341 VDD.n214 VSUBS 0.00347f
C342 VDD.n215 VSUBS 0.00347f
C343 VDD.n216 VSUBS 0.00347f
C344 VDD.n217 VSUBS 0.00347f
C345 VDD.n218 VSUBS 0.00347f
C346 VDD.n219 VSUBS 0.199f
C347 VDD.n220 VSUBS 0.00347f
C348 VDD.n221 VSUBS 0.00347f
C349 VDD.t18 VSUBS 0.106f
C350 VDD.n222 VSUBS 0.00347f
C351 VDD.n223 VSUBS 0.00347f
C352 VDD.n224 VSUBS 0.00347f
C353 VDD.n225 VSUBS 0.119f
C354 VDD.n226 VSUBS 0.00347f
C355 VDD.n227 VSUBS 0.00347f
C356 VDD.n228 VSUBS 0.00347f
C357 VDD.n229 VSUBS 0.00347f
C358 VDD.n230 VSUBS 0.00347f
C359 VDD.n231 VSUBS 0.212f
C360 VDD.n232 VSUBS 0.00347f
C361 VDD.n233 VSUBS 0.00347f
C362 VDD.n234 VSUBS 0.00347f
C363 VDD.n235 VSUBS 0.00347f
C364 VDD.n236 VSUBS 0.00347f
C365 VDD.n237 VSUBS 0.184f
C366 VDD.n238 VSUBS 0.00347f
C367 VDD.n239 VSUBS 0.00347f
C368 VDD.t21 VSUBS 0.106f
C369 VDD.n240 VSUBS 0.00347f
C370 VDD.n241 VSUBS 0.00347f
C371 VDD.n242 VSUBS 0.00347f
C372 VDD.n243 VSUBS 0.134f
C373 VDD.n244 VSUBS 0.00347f
C374 VDD.n245 VSUBS 0.00347f
C375 VDD.n246 VSUBS 0.00347f
C376 VDD.n247 VSUBS 0.00347f
C377 VDD.n248 VSUBS 0.00347f
C378 VDD.n249 VSUBS 0.212f
C379 VDD.n250 VSUBS 0.00347f
C380 VDD.n251 VSUBS 0.00347f
C381 VDD.n252 VSUBS 0.00347f
C382 VDD.n253 VSUBS 0.00347f
C383 VDD.n254 VSUBS 0.00347f
C384 VDD.n255 VSUBS 0.168f
C385 VDD.n256 VSUBS 0.00347f
C386 VDD.n257 VSUBS 0.00347f
C387 VDD.t4 VSUBS 0.106f
C388 VDD.n258 VSUBS 0.00347f
C389 VDD.n259 VSUBS 0.00347f
C390 VDD.n260 VSUBS 0.00347f
C391 VDD.n261 VSUBS 0.149f
C392 VDD.n262 VSUBS 0.00347f
C393 VDD.n263 VSUBS 0.00347f
C394 VDD.n264 VSUBS 0.00347f
C395 VDD.n265 VSUBS 0.00347f
C396 VDD.n266 VSUBS 0.00347f
C397 VDD.n267 VSUBS 0.212f
C398 VDD.n268 VSUBS 0.00347f
C399 VDD.n269 VSUBS 0.00347f
C400 VDD.t12 VSUBS 0.106f
C401 VDD.n270 VSUBS 0.00347f
C402 VDD.n271 VSUBS 0.00347f
C403 VDD.n272 VSUBS 0.00347f
C404 VDD.n273 VSUBS 0.153f
C405 VDD.n274 VSUBS 0.00347f
C406 VDD.n275 VSUBS 0.00347f
C407 VDD.n276 VSUBS 0.00347f
C408 VDD.n277 VSUBS 0.164f
C409 VDD.n278 VSUBS 0.00347f
C410 VDD.n279 VSUBS 0.00347f
C411 VDD.n280 VSUBS 0.00347f
C412 VDD.n281 VSUBS 0.212f
C413 VDD.n282 VSUBS 0.00347f
C414 VDD.n283 VSUBS 0.00347f
C415 VDD.t25 VSUBS 0.106f
C416 VDD.n284 VSUBS 0.00347f
C417 VDD.n285 VSUBS 0.138f
C418 VDD.n286 VSUBS 0.00347f
C419 VDD.n287 VSUBS 0.00347f
C420 VDD.n288 VSUBS 0.00347f
C421 VDD.n289 VSUBS 0.179f
C422 VDD.n290 VSUBS 0.00347f
C423 VDD.n291 VSUBS 0.00347f
C424 VDD.n292 VSUBS 0.00347f
C425 VDD.n293 VSUBS 0.212f
C426 VDD.n294 VSUBS 0.00347f
C427 VDD.n295 VSUBS 0.00347f
C428 VDD.t28 VSUBS 0.106f
C429 VDD.n296 VSUBS 0.00347f
C430 VDD.n297 VSUBS 0.123f
C431 VDD.n298 VSUBS 0.00347f
C432 VDD.n299 VSUBS 0.00347f
C433 VDD.n300 VSUBS 0.00347f
C434 VDD.n301 VSUBS 0.194f
C435 VDD.n302 VSUBS 0.00347f
C436 VDD.n303 VSUBS 0.00347f
C437 VDD.n304 VSUBS 0.00347f
C438 VDD.n305 VSUBS 0.212f
C439 VDD.n306 VSUBS 0.00347f
C440 VDD.n307 VSUBS 0.00347f
C441 VDD.t11 VSUBS 0.106f
C442 VDD.n308 VSUBS 0.00347f
C443 VDD.n309 VSUBS 0.108f
C444 VDD.n310 VSUBS 0.00347f
C445 VDD.n311 VSUBS 0.00347f
C446 VDD.n312 VSUBS 0.00347f
C447 VDD.n313 VSUBS 0.21f
C448 VDD.n314 VSUBS 0.00347f
C449 VDD.n315 VSUBS 0.00347f
C450 VDD.n316 VSUBS 0.00347f
C451 VDD.n317 VSUBS 0.199f
C452 VDD.n318 VSUBS 0.00347f
C453 VDD.n319 VSUBS 0.00347f
C454 VDD.t10 VSUBS 0.106f
C455 VDD.n320 VSUBS 0.00347f
C456 VDD.n321 VSUBS 0.119f
C457 VDD.n322 VSUBS 0.00347f
C458 VDD.n323 VSUBS 0.00347f
C459 VDD.n324 VSUBS 0.00347f
C460 VDD.n325 VSUBS 0.212f
C461 VDD.n326 VSUBS 0.00347f
C462 VDD.n327 VSUBS 0.00347f
C463 VDD.n328 VSUBS 0.00347f
C464 VDD.n329 VSUBS 0.184f
C465 VDD.n330 VSUBS 0.00347f
C466 VDD.n331 VSUBS 0.00347f
C467 VDD.t2 VSUBS 0.106f
C468 VDD.n332 VSUBS 0.00347f
C469 VDD.n333 VSUBS 0.134f
C470 VDD.n334 VSUBS 0.00347f
C471 VDD.n335 VSUBS 0.00347f
C472 VDD.n336 VSUBS 0.00347f
C473 VDD.n337 VSUBS 0.212f
C474 VDD.n338 VSUBS 0.00347f
C475 VDD.n339 VSUBS 0.00347f
C476 VDD.n340 VSUBS 0.00347f
C477 VDD.n341 VSUBS 0.168f
C478 VDD.n342 VSUBS 0.00347f
C479 VDD.n343 VSUBS 0.00347f
C480 VDD.t19 VSUBS 0.106f
C481 VDD.n344 VSUBS 0.00347f
C482 VDD.n345 VSUBS 0.149f
C483 VDD.n346 VSUBS 0.00347f
C484 VDD.n347 VSUBS 0.00347f
C485 VDD.n348 VSUBS 0.00347f
C486 VDD.n349 VSUBS 0.212f
C487 VDD.n350 VSUBS 0.00347f
C488 VDD.n351 VSUBS 0.00347f
C489 VDD.t35 VSUBS 0.106f
C490 VDD.n352 VSUBS 0.00347f
C491 VDD.n353 VSUBS 0.153f
C492 VDD.n354 VSUBS 0.00347f
C493 VDD.n355 VSUBS 0.00347f
C494 VDD.n356 VSUBS 0.00347f
C495 VDD.n357 VSUBS 0.164f
C496 VDD.n358 VSUBS 0.00347f
C497 VDD.n359 VSUBS 0.00347f
C498 VDD.n360 VSUBS 0.00347f
C499 VDD.n361 VSUBS 0.212f
C500 VDD.n362 VSUBS 0.00347f
C501 VDD.n363 VSUBS 0.00347f
C502 VDD.t22 VSUBS 0.106f
C503 VDD.n364 VSUBS 0.138f
C504 VDD.n365 VSUBS 0.00347f
C505 VDD.n366 VSUBS 0.00347f
C506 VDD.n367 VSUBS 0.179f
C507 VDD.n368 VSUBS 0.00347f
C508 VDD.n369 VSUBS 0.00347f
C509 VDD.n370 VSUBS 0.212f
C510 VDD.n371 VSUBS 0.00347f
C511 VDD.n372 VSUBS 0.00347f
C512 VDD.n373 VSUBS 0.00404f
C513 VDD.n374 VSUBS 0.00482f
C514 VDD.n375 VSUBS 0.00283f
C515 VDD.n377 VSUBS 0.00347f
C516 VDD.n378 VSUBS 0.00347f
C517 VDD.n380 VSUBS 0.00347f
C518 VDD.n396 VSUBS 0.335f
C519 VDD.n398 VSUBS 0.00482f
C520 VDD.n399 VSUBS 0.00482f
C521 VDD.n400 VSUBS 0.00283f
C522 VDD.n401 VSUBS 0.00283f
C523 VDD.n403 VSUBS 0.00347f
C524 VDD.n404 VSUBS 0.00336f
C525 VDD.n405 VSUBS 0.0139f
C526 VDD.n407 VSUBS 0.00347f
C527 VDD.n408 VSUBS 0.00184f
C528 VDD.n410 VSUBS 0.00347f
C529 VDD.n411 VSUBS 0.00347f
C530 VDD.n413 VSUBS 0.00347f
C531 VDD.n414 VSUBS 0.00347f
C532 VDD.n416 VSUBS 0.00347f
C533 VDD.n417 VSUBS 0.0022f
C534 VDD.n418 VSUBS 0.0139f
C535 VDD.n420 VSUBS 0.00347f
C536 VDD.n421 VSUBS 0.00301f
C537 VDD.n423 VSUBS 0.00347f
C538 VDD.n424 VSUBS 0.00347f
C539 VDD.n426 VSUBS 0.00347f
C540 VDD.n427 VSUBS 0.00271f
C541 VDD.n428 VSUBS 0.0139f
C542 VDD.n430 VSUBS 0.00347f
C543 VDD.n431 VSUBS 0.0025f
C544 VDD.n433 VSUBS 0.00347f
C545 VDD.n434 VSUBS 0.00347f
C546 VDD.n436 VSUBS 0.00347f
C547 VDD.n437 VSUBS 0.00347f
C548 VDD.n439 VSUBS 0.00347f
C549 VDD.n440 VSUBS 0.00175f
C550 VDD.n441 VSUBS 0.0139f
C551 VDD.n443 VSUBS 0.00347f
C552 VDD.n444 VSUBS 0.00345f
C553 VDD.n446 VSUBS 0.00347f
C554 VDD.n447 VSUBS 0.00347f
C555 VDD.n449 VSUBS 0.00347f
C556 VDD.n450 VSUBS 0.00218f
C557 VDD.n451 VSUBS 0.0138f
C558 VDD.n452 VSUBS 0.00347f
C559 VDD.n453 VSUBS 0.00303f
C560 VDD.n454 VSUBS 0.00347f
C561 VDD.n455 VSUBS 0.00347f
C562 VDD.n456 VSUBS 0.00347f
C563 VDD.n457 VSUBS 0.00282f
C564 VDD.n458 VSUBS 0.0139f
C565 VDD.n459 VSUBS 0.00347f
C566 VDD.n460 VSUBS 0.00239f
C567 VDD.n461 VSUBS 0.00347f
C568 VDD.n462 VSUBS 0.00347f
C569 VDD.n463 VSUBS 0.00276f
C570 VDD.n464 VSUBS 0.00276f
C571 VDD.n465 VSUBS 0.00475f
C572 VDD.n466 VSUBS 0.00446f
C573 VDD.t42 VSUBS 0.00743f
C574 VDD.t43 VSUBS 0.00743f
C575 VDD.t23 VSUBS 0.00743f
C576 VDD.t24 VSUBS 0.00743f
C577 VDD.t48 VSUBS 0.00743f
C578 VDD.t49 VSUBS 0.00743f
C579 VDD.n467 VSUBS 0.00347f
C580 VDD.n468 VSUBS 0.00347f
C581 VDD.n469 VSUBS 0.00347f
C582 VDD.n470 VSUBS 0.00347f
C583 VDD.n471 VSUBS 0.00347f
C584 VDD.n472 VSUBS 0.00347f
C585 VDD.n473 VSUBS 0.00347f
C586 VDD.n474 VSUBS 0.00347f
C587 VDD.n475 VSUBS 0.00347f
C588 VDD.n476 VSUBS 0.00347f
C589 VDD.n477 VSUBS 0.00347f
C590 VDD.n478 VSUBS 0.00347f
C591 VDD.n479 VSUBS 0.00347f
C592 VDD.n480 VSUBS 0.00347f
C593 VDD.n481 VSUBS 0.00347f
C594 VDD.n482 VSUBS 0.00347f
C595 VDD.n483 VSUBS 0.00347f
C596 VDD.n484 VSUBS 0.00347f
C597 VDD.n485 VSUBS 0.00347f
C598 VDD.n486 VSUBS 0.00347f
C599 VDD.n487 VSUBS 0.00347f
C600 VDD.n488 VSUBS 0.00347f
C601 VDD.n489 VSUBS 0.00347f
C602 VDD.n490 VSUBS 0.00347f
C603 VDD.n491 VSUBS 0.00347f
C604 VDD.n492 VSUBS 0.00347f
C605 VDD.n493 VSUBS 0.00347f
C606 VDD.n494 VSUBS 0.00347f
C607 VDD.n495 VSUBS 0.00347f
C608 VDD.n496 VSUBS 0.00347f
C609 VDD.n497 VSUBS 0.00347f
C610 VDD.n498 VSUBS 0.00347f
C611 VDD.n499 VSUBS 0.00347f
C612 VDD.n500 VSUBS 0.00347f
C613 VDD.n501 VSUBS 0.00347f
C614 VDD.n502 VSUBS 0.00404f
C615 VDD.n503 VSUBS 0.00404f
C616 VDD.n504 VSUBS 0.00482f
C617 VDD.n505 VSUBS 0.00283f
C618 VDD.n506 VSUBS 0.00335f
C619 VDD.n507 VSUBS 0.0139f
C620 VDD.n508 VSUBS 0.00186f
C621 VDD.n509 VSUBS 0.00347f
C622 VDD.n510 VSUBS 0.00347f
C623 VDD.n511 VSUBS 0.00347f
C624 VDD.n512 VSUBS 0.00347f
C625 VDD.n513 VSUBS 0.00218f
C626 VDD.n514 VSUBS 0.0139f
C627 VDD.n515 VSUBS 0.00347f
C628 VDD.n516 VSUBS 0.00303f
C629 VDD.n517 VSUBS 0.00347f
C630 VDD.n518 VSUBS 0.00347f
C631 VDD.n519 VSUBS 0.00347f
C632 VDD.n520 VSUBS 0.00269f
C633 VDD.n521 VSUBS 0.0139f
C634 VDD.n522 VSUBS 0.00347f
C635 VDD.n523 VSUBS 0.00251f
C636 VDD.n524 VSUBS 0.00347f
C637 VDD.n525 VSUBS 0.00347f
C638 VDD.n526 VSUBS 0.00347f
C639 VDD.n527 VSUBS 0.00347f
C640 VDD.n528 VSUBS 0.00347f
C641 VDD.n529 VSUBS 0.0156f
C642 VDD.n530 VSUBS 0.00347f
C643 VDD.n531 VSUBS 0.00347f
C644 VDD.n532 VSUBS 0.00347f
C645 VDD.n533 VSUBS 0.00347f
C646 VDD.n534 VSUBS 0.00347f
C647 VDD.n535 VSUBS 0.00216f
C648 VDD.n536 VSUBS 0.0138f
C649 VDD.n537 VSUBS 0.00347f
C650 VDD.n538 VSUBS 0.00305f
C651 VDD.n539 VSUBS 0.00347f
C652 VDD.n540 VSUBS 0.00347f
C653 VDD.n541 VSUBS 0.00347f
C654 VDD.n542 VSUBS 0.0028f
C655 VDD.n543 VSUBS 0.0139f
C656 VDD.n544 VSUBS 0.00347f
C657 VDD.n545 VSUBS 0.00241f
C658 VDD.n546 VSUBS 0.00347f
C659 VDD.n547 VSUBS 0.00347f
C660 VDD.n548 VSUBS 0.00276f
C661 VDD.n549 VSUBS 0.00276f
C662 VDD.n550 VSUBS 0.00475f
C663 VDD.n551 VSUBS 0.00446f
C664 VDD.n552 VSUBS 0.005f
C665 VDD.n553 VSUBS 0.00404f
C666 VDD.n554 VSUBS 0.00404f
C667 VDD.n555 VSUBS 0.00686f
C668 VDD.n556 VSUBS 0.00347f
C669 VDD.n557 VSUBS 0.00347f
C670 VDD.n558 VSUBS 0.0118f
C671 VDD.n559 VSUBS 0.00347f
C672 VDD.n560 VSUBS 0.00347f
C673 VDD.n561 VSUBS 0.0118f
C674 VDD.n562 VSUBS 0.00347f
C675 VDD.n563 VSUBS 0.00347f
C676 VDD.n564 VSUBS 0.0118f
C677 VDD.n565 VSUBS 0.00347f
C678 VDD.n566 VSUBS 0.00347f
C679 VDD.n567 VSUBS 0.0118f
C680 VDD.n568 VSUBS 0.00347f
C681 VDD.n569 VSUBS 0.00347f
C682 VDD.n570 VSUBS 0.0118f
C683 VDD.n571 VSUBS 0.00347f
C684 VDD.n572 VSUBS 0.00347f
C685 VDD.n573 VSUBS 0.0118f
C686 VDD.n574 VSUBS 0.00347f
C687 VDD.n575 VSUBS 0.00347f
C688 VDD.n576 VSUBS 0.0118f
C689 VDD.n577 VSUBS 0.00347f
C690 VDD.n578 VSUBS 0.00347f
C691 VDD.n579 VSUBS 0.0118f
C692 VDD.n580 VSUBS 0.00347f
C693 VDD.n581 VSUBS 0.00347f
C694 VDD.n582 VSUBS 0.0118f
C695 VDD.n583 VSUBS 0.00347f
C696 VDD.n584 VSUBS 0.00347f
C697 VDD.n585 VSUBS 0.0118f
C698 VDD.n586 VSUBS 0.00347f
C699 VDD.n587 VSUBS 0.00347f
C700 VDD.n588 VSUBS 0.0118f
C701 VDD.n589 VSUBS 0.00347f
C702 VDD.n590 VSUBS 0.00347f
C703 VDD.n591 VSUBS 0.0118f
C704 VDD.n592 VSUBS 0.00347f
C705 VDD.n593 VSUBS 0.00347f
C706 VDD.n594 VSUBS 0.0118f
C707 VDD.n595 VSUBS 0.00347f
C708 VDD.n596 VSUBS 0.00347f
C709 VDD.n597 VSUBS 0.0118f
C710 VDD.n598 VSUBS 0.00347f
C711 VDD.n599 VSUBS 0.00347f
C712 VDD.n600 VSUBS 0.0118f
C713 VDD.n601 VSUBS 0.00347f
C714 VDD.n602 VSUBS 0.00347f
C715 VDD.n603 VSUBS 0.0118f
C716 VDD.n604 VSUBS 0.00347f
C717 VDD.n605 VSUBS 0.00347f
C718 VDD.n606 VSUBS 0.0118f
C719 VDD.n607 VSUBS 0.00347f
C720 VDD.n608 VSUBS 0.00347f
C721 VDD.n609 VSUBS 0.0118f
C722 VDD.n610 VSUBS 0.00347f
C723 VDD.n611 VSUBS 0.00347f
C724 VDD.n612 VSUBS 0.0118f
C725 VDD.n613 VSUBS 0.00347f
C726 VDD.n614 VSUBS 0.00347f
C727 VDD.n615 VSUBS 0.0118f
C728 VDD.n616 VSUBS 0.00347f
C729 VDD.n617 VSUBS 0.00347f
C730 VDD.n618 VSUBS 0.0118f
C731 VDD.n619 VSUBS 0.00347f
C732 VDD.n620 VSUBS 0.00347f
C733 VDD.n621 VSUBS 0.0118f
C734 VDD.n622 VSUBS 0.00347f
C735 VDD.n623 VSUBS 0.00347f
C736 VDD.n624 VSUBS 0.0118f
C737 VDD.n625 VSUBS 0.00347f
C738 VDD.n626 VSUBS 0.00347f
C739 VDD.n627 VSUBS 0.0118f
C740 VDD.n628 VSUBS 0.00347f
C741 VDD.n629 VSUBS 0.00347f
C742 VDD.n630 VSUBS 0.0118f
C743 VDD.n631 VSUBS 0.0118f
C744 VDD.n632 VSUBS 0.0118f
C745 VDD.n633 VSUBS 0.0118f
C746 VDD.n634 VSUBS 0.0118f
C747 VDD.n635 VSUBS 0.0118f
C748 VDD.n636 VSUBS 0.0118f
C749 VDD.n637 VSUBS 0.0118f
C750 VDD.n638 VSUBS 0.0118f
C751 VDD.n639 VSUBS 0.0118f
C752 VDD.n640 VSUBS 0.0118f
C753 VDD.n641 VSUBS 0.0118f
C754 VDD.n642 VSUBS 0.0118f
C755 VDD.n643 VSUBS 0.0118f
C756 VDD.n644 VSUBS 0.0118f
C757 VDD.n645 VSUBS 0.0118f
C758 VDD.n646 VSUBS 0.0118f
C759 VDD.n647 VSUBS 0.0118f
C760 VDD.n648 VSUBS 0.0118f
C761 VDD.n649 VSUBS 0.0118f
C762 VDD.n650 VSUBS 0.0118f
C763 VDD.n651 VSUBS 0.0118f
C764 VDD.n652 VSUBS 0.0118f
C765 VDD.n653 VSUBS 0.0118f
C766 VDD.n654 VSUBS 0.0118f
C767 VDD.n655 VSUBS 0.0118f
C768 VDD.n656 VSUBS 0.0118f
C769 VDD.n657 VSUBS 0.0118f
C770 VDD.n658 VSUBS 0.0118f
C771 VDD.n659 VSUBS 0.0118f
C772 VDD.n660 VSUBS 0.0118f
C773 VDD.n661 VSUBS 0.0118f
C774 VDD.n662 VSUBS 0.0118f
C775 VDD.n663 VSUBS 0.0118f
C776 VDD.n664 VSUBS 0.0118f
C777 VDD.n665 VSUBS 0.0118f
C778 VDD.n666 VSUBS 0.0118f
C779 VDD.n667 VSUBS 0.00771f
C780 VDD.n668 VSUBS 0.00999f
C781 VDD.n669 VSUBS 0.0118f
C782 VDD.n670 VSUBS 0.0118f
C783 VDD.n671 VSUBS 0.0118f
C784 VDD.n672 VSUBS 0.0118f
C785 VDD.n673 VSUBS 0.0118f
C786 VDD.n674 VSUBS 0.0118f
C787 VDD.n675 VSUBS 0.0118f
C788 VDD.n676 VSUBS 0.0118f
C789 VDD.n677 VSUBS 0.0118f
C790 VDD.n678 VSUBS 0.0118f
C791 VDD.n679 VSUBS 0.0118f
C792 VDD.n680 VSUBS 0.0118f
C793 VDD.n681 VSUBS 0.0118f
C794 VDD.n682 VSUBS 0.0118f
C795 VDD.n683 VSUBS 0.0118f
C796 VDD.n684 VSUBS 0.0118f
C797 VDD.n685 VSUBS 0.0118f
C798 VDD.n686 VSUBS 0.0118f
C799 VDD.n687 VSUBS 0.0118f
C800 VDD.n688 VSUBS 0.0118f
C801 VDD.n689 VSUBS 0.0118f
C802 VDD.n690 VSUBS 0.0118f
C803 VDD.n691 VSUBS 0.0118f
C804 VDD.n692 VSUBS 0.0118f
C805 VDD.n693 VSUBS 0.0118f
C806 VDD.n694 VSUBS 0.0118f
C807 VDD.n695 VSUBS 0.0118f
C808 VDD.n696 VSUBS 0.0118f
C809 VDD.n697 VSUBS 0.0118f
C810 VDD.n698 VSUBS 0.00347f
C811 VDD.n699 VSUBS 0.00347f
C812 VDD.n700 VSUBS 0.0118f
C813 VDD.n701 VSUBS 0.00347f
C814 VDD.n702 VSUBS 0.00347f
C815 VDD.n703 VSUBS 0.0118f
C816 VDD.n704 VSUBS 0.00347f
C817 VDD.n705 VSUBS 0.00347f
C818 VDD.n706 VSUBS 0.0118f
C819 VDD.n707 VSUBS 0.00347f
C820 VDD.n708 VSUBS 0.00347f
C821 VDD.n709 VSUBS 0.0118f
C822 VDD.n710 VSUBS 0.00347f
C823 VDD.n711 VSUBS 0.00347f
C824 VDD.n712 VSUBS 0.0118f
C825 VDD.n713 VSUBS 0.00347f
C826 VDD.n714 VSUBS 0.00347f
C827 VDD.n715 VSUBS 0.0118f
C828 VDD.n716 VSUBS 0.00347f
C829 VDD.n717 VSUBS 0.00347f
C830 VDD.n718 VSUBS 0.0118f
C831 VDD.n719 VSUBS 0.00347f
C832 VDD.n720 VSUBS 0.00347f
C833 VDD.n721 VSUBS 0.00939f
C834 VDD.n722 VSUBS 0.00523f
C835 VDD.n723 VSUBS 0.00176f
C836 VDD.n724 VSUBS 0.00178f
C837 VDD.n725 VSUBS 0.00347f
C838 VDD.n726 VSUBS 0.00178f
C839 VDD.n727 VSUBS 0.00347f
C840 VDD.n728 VSUBS 0.00122f
C841 VDD.n729 VSUBS 0.0131f
C842 VDD.n730 VSUBS 0.00347f
C843 VDD.n731 VSUBS 0.00144f
C844 VDD.n732 VSUBS 0.00347f
C845 VDD.n733 VSUBS 0.00178f
C846 VDD.n734 VSUBS 0.00347f
C847 VDD.n735 VSUBS 0.00156f
C848 VDD.n736 VSUBS 0.0117f
C849 VDD.n737 VSUBS 0.00347f
C850 VDD.n738 VSUBS 0.00111f
C851 VDD.n739 VSUBS 0.00347f
C852 VDD.n740 VSUBS 0.00178f
C853 VDD.n741 VSUBS 0.00347f
C854 VDD.n742 VSUBS 0.00178f
C855 VDD.n743 VSUBS 0.00347f
C856 VDD.n744 VSUBS 0.00101f
C857 VDD.n745 VSUBS 0.0145f
C858 VDD.n746 VSUBS 0.00347f
C859 VDD.n747 VSUBS 8.71e-19
C860 VDD.n748 VSUBS 0.0305f
C861 VDD.n749 VSUBS 0.00347f
C862 VDD.n750 VSUBS 0.00168f
C863 VDD.n751 VSUBS 0.00347f
C864 VDD.n752 VSUBS 0.00124f
C865 VDD.n753 VSUBS 0.0145f
C866 VDD.n754 VSUBS 0.00347f
C867 VDD.n755 VSUBS 0.00142f
C868 VDD.n756 VSUBS 0.00347f
C869 VDD.n757 VSUBS 0.00178f
C870 VDD.n758 VSUBS 0.00347f
C871 VDD.n759 VSUBS 0.00178f
C872 VDD.n761 VSUBS 0.00347f
C873 VDD.n762 VSUBS 0.00178f
C874 VDD.n763 VSUBS 0.00347f
C875 VDD.n764 VSUBS 0.00178f
C876 VDD.n766 VSUBS 0.00347f
C877 VDD.n767 VSUBS 0.00178f
C878 VDD.n768 VSUBS 0.00347f
C879 VDD.n769 VSUBS 0.00178f
C880 VDD.n771 VSUBS 0.00347f
C881 VDD.n772 VSUBS 0.00178f
C882 VDD.n773 VSUBS 0.00283f
C883 VDD.n774 VSUBS 0.00145f
C884 VDD.n775 VSUBS 0.0023f
C885 VDD.n776 VSUBS 0.00347f
C886 VDD.n777 VSUBS 0.212f
C887 VDD.n778 VSUBS 0.00347f
C888 VDD.n779 VSUBS 0.00313f
C889 VDD.n780 VSUBS 0.00347f
C890 VDD.n781 VSUBS 0.212f
C891 VDD.n782 VSUBS 0.00347f
C892 VDD.n783 VSUBS 0.00347f
C893 VDD.n784 VSUBS 0.00347f
C894 VDD.n785 VSUBS 0.212f
C895 VDD.n786 VSUBS 0.00347f
C896 VDD.n787 VSUBS 0.00347f
C897 VDD.t13 VSUBS 0.106f
C898 VDD.n788 VSUBS 0.00347f
C899 VDD.n789 VSUBS 0.108f
C900 VDD.n790 VSUBS 0.00347f
C901 VDD.n791 VSUBS 0.00191f
C902 VDD.n792 VSUBS 0.00558f
C903 VDD.n793 VSUBS 0.00347f
C904 VDD.n794 VSUBS 0.21f
C905 VDD.n795 VSUBS 0.00347f
C906 VDD.n796 VSUBS 0.00329f
C907 VDD.n797 VSUBS 0.00347f
C908 VDD.n798 VSUBS 0.199f
C909 VDD.n799 VSUBS 0.00347f
C910 VDD.n800 VSUBS 0.00347f
C911 VDD.t5 VSUBS 0.106f
C912 VDD.n801 VSUBS 0.00347f
C913 VDD.n802 VSUBS 0.119f
C914 VDD.n803 VSUBS 0.00347f
C915 VDD.n804 VSUBS 0.00347f
C916 VDD.n805 VSUBS 0.00347f
C917 VDD.n806 VSUBS 0.212f
C918 VDD.n807 VSUBS 0.00347f
C919 VDD.n808 VSUBS 0.00347f
C920 VDD.n809 VSUBS 0.00347f
C921 VDD.n810 VSUBS 0.00347f
C922 VDD.n811 VSUBS 0.00347f
C923 VDD.n812 VSUBS 0.184f
C924 VDD.n813 VSUBS 0.00347f
C925 VDD.n814 VSUBS 0.00347f
C926 VDD.t36 VSUBS 0.106f
C927 VDD.n815 VSUBS 0.00347f
C928 VDD.n816 VSUBS 0.00347f
C929 VDD.n817 VSUBS 0.00347f
C930 VDD.n818 VSUBS 0.134f
C931 VDD.n819 VSUBS 0.00347f
C932 VDD.n820 VSUBS 0.00347f
C933 VDD.n821 VSUBS 0.00347f
C934 VDD.n822 VSUBS 0.00347f
C935 VDD.n823 VSUBS 0.00347f
C936 VDD.n824 VSUBS 0.212f
C937 VDD.n825 VSUBS 0.00347f
C938 VDD.n826 VSUBS 0.00347f
C939 VDD.n827 VSUBS 0.00347f
C940 VDD.n828 VSUBS 0.00347f
C941 VDD.n829 VSUBS 0.00347f
C942 VDD.n830 VSUBS 0.00347f
C943 VDD.n831 VSUBS 0.168f
C944 VDD.n832 VSUBS 0.00347f
C945 VDD.n833 VSUBS 0.00347f
C946 VDD.t33 VSUBS 0.106f
C947 VDD.n834 VSUBS 0.00347f
C948 VDD.n835 VSUBS 0.00347f
C949 VDD.n836 VSUBS 0.00347f
C950 VDD.n837 VSUBS 0.00347f
C951 VDD.n838 VSUBS 0.149f
C952 VDD.n839 VSUBS 0.00347f
C953 VDD.n840 VSUBS 0.00347f
C954 VDD.n841 VSUBS 0.00347f
C955 VDD.n842 VSUBS 0.00347f
C956 VDD.n843 VSUBS 0.00347f
C957 VDD.n844 VSUBS 0.00347f
C958 VDD.n845 VSUBS 0.212f
C959 VDD.n846 VSUBS 0.00347f
C960 VDD.n847 VSUBS 0.00347f
C961 VDD.t0 VSUBS 0.106f
C962 VDD.n848 VSUBS 0.00347f
C963 VDD.n849 VSUBS 0.00347f
C964 VDD.n850 VSUBS 0.00347f
C965 VDD.n851 VSUBS 0.00347f
C966 VDD.n852 VSUBS 0.153f
C967 VDD.n853 VSUBS 0.00347f
C968 VDD.n854 VSUBS 0.00347f
C969 VDD.n855 VSUBS 0.00347f
C970 VDD.n856 VSUBS 0.00347f
C971 VDD.n857 VSUBS 0.00347f
C972 VDD.n858 VSUBS 0.164f
C973 VDD.n859 VSUBS 0.00347f
C974 VDD.n860 VSUBS 0.00347f
C975 VDD.n861 VSUBS 0.00347f
C976 VDD.n862 VSUBS 0.00347f
C977 VDD.n863 VSUBS 0.00347f
C978 VDD.n864 VSUBS 0.00347f
C979 VDD.n865 VSUBS 0.00347f
C980 VDD.n866 VSUBS 0.212f
C981 VDD.n867 VSUBS 0.00347f
C982 VDD.n868 VSUBS 0.00347f
C983 VDD.t30 VSUBS 0.106f
C984 VDD.n869 VSUBS 0.00347f
C985 VDD.n870 VSUBS 0.00347f
C986 VDD.n871 VSUBS 0.00347f
C987 VDD.n872 VSUBS 0.138f
C988 VDD.n873 VSUBS 0.00347f
C989 VDD.n874 VSUBS 0.00347f
C990 VDD.n875 VSUBS 0.00347f
C991 VDD.n876 VSUBS 0.00347f
C992 VDD.n877 VSUBS 0.00347f
C993 VDD.n878 VSUBS 0.179f
C994 VDD.n879 VSUBS 0.00347f
C995 VDD.n880 VSUBS 0.00347f
C996 VDD.n881 VSUBS 0.00347f
C997 VDD.n882 VSUBS 0.00347f
C998 VDD.n883 VSUBS 0.00347f
C999 VDD.n884 VSUBS 0.212f
C1000 VDD.n885 VSUBS 0.00347f
C1001 VDD.n886 VSUBS 0.00347f
C1002 VDD.t34 VSUBS 0.106f
C1003 VDD.n887 VSUBS 0.00347f
C1004 VDD.n888 VSUBS 0.00347f
C1005 VDD.n889 VSUBS 0.00347f
C1006 VDD.n890 VSUBS 0.123f
C1007 VDD.n891 VSUBS 0.00347f
C1008 VDD.n892 VSUBS 0.00347f
C1009 VDD.n893 VSUBS 0.00347f
C1010 VDD.n894 VSUBS 0.00347f
C1011 VDD.n895 VSUBS 0.00347f
C1012 VDD.n896 VSUBS 0.194f
C1013 VDD.n897 VSUBS 0.00347f
C1014 VDD.n898 VSUBS 0.00347f
C1015 VDD.n899 VSUBS 0.00347f
C1016 VDD.n900 VSUBS 0.00347f
C1017 VDD.n901 VSUBS 0.00347f
C1018 VDD.n902 VSUBS 0.212f
C1019 VDD.n903 VSUBS 0.00347f
C1020 VDD.n904 VSUBS 0.00347f
C1021 VDD.t37 VSUBS 0.106f
C1022 VDD.n905 VSUBS 0.00347f
C1023 VDD.n906 VSUBS 0.00347f
C1024 VDD.n907 VSUBS 0.00347f
C1025 VDD.n908 VSUBS 0.108f
C1026 VDD.n909 VSUBS 0.00347f
C1027 VDD.n910 VSUBS 0.00347f
C1028 VDD.n911 VSUBS 0.00347f
C1029 VDD.n912 VSUBS 0.00347f
C1030 VDD.n913 VSUBS 0.00347f
C1031 VDD.n914 VSUBS 0.21f
C1032 VDD.n915 VSUBS 0.00347f
C1033 VDD.n916 VSUBS 0.00347f
C1034 VDD.n917 VSUBS 0.00347f
C1035 VDD.n918 VSUBS 0.00347f
C1036 VDD.n919 VSUBS 0.00347f
C1037 VDD.n920 VSUBS 0.199f
C1038 VDD.n921 VSUBS 0.00347f
C1039 VDD.n922 VSUBS 0.00347f
C1040 VDD.t7 VSUBS 0.106f
C1041 VDD.n923 VSUBS 0.00347f
C1042 VDD.n924 VSUBS 0.00347f
C1043 VDD.n925 VSUBS 0.00347f
C1044 VDD.n926 VSUBS 0.119f
C1045 VDD.n927 VSUBS 0.00347f
C1046 VDD.n928 VSUBS 0.00347f
C1047 VDD.n929 VSUBS 0.00347f
C1048 VDD.n930 VSUBS 0.00347f
C1049 VDD.n931 VSUBS 0.00347f
C1050 VDD.n932 VSUBS 0.212f
C1051 VDD.n933 VSUBS 0.00347f
C1052 VDD.n934 VSUBS 0.00347f
C1053 VDD.n935 VSUBS 0.00347f
C1054 VDD.n936 VSUBS 0.00347f
C1055 VDD.n937 VSUBS 0.00347f
C1056 VDD.n938 VSUBS 0.00347f
C1057 VDD.n939 VSUBS 0.00347f
C1058 VDD.n940 VSUBS 0.00347f
C1059 VDD.n941 VSUBS 0.00347f
C1060 VDD.n942 VSUBS 0.00347f
C1061 VDD.n943 VSUBS 0.00347f
C1062 VDD.n944 VSUBS 0.00347f
C1063 VDD.n945 VSUBS 0.00347f
C1064 VDD.n946 VSUBS 0.00347f
C1065 VDD.n947 VSUBS 0.00347f
C1066 VDD.n948 VSUBS 0.00347f
C1067 VDD.n949 VSUBS 0.00347f
C1068 VDD.n950 VSUBS 0.184f
C1069 VDD.n951 VSUBS 0.00347f
C1070 VDD.n952 VSUBS 0.00347f
C1071 VDD.t29 VSUBS 0.106f
C1072 VDD.n953 VSUBS 0.00347f
C1073 VDD.n954 VSUBS 0.00347f
C1074 VDD.n955 VSUBS 0.00347f
C1075 VDD.n956 VSUBS 0.134f
C1076 VDD.n957 VSUBS 0.00347f
C1077 VDD.n958 VSUBS 0.00347f
C1078 VDD.n959 VSUBS 0.00347f
C1079 VDD.n960 VSUBS 0.00347f
C1080 VDD.n961 VSUBS 0.00347f
C1081 VDD.n962 VSUBS 0.212f
C1082 VDD.n963 VSUBS 0.00347f
C1083 VDD.n964 VSUBS 0.00347f
C1084 VDD.n965 VSUBS 0.00347f
C1085 VDD.n966 VSUBS 0.00347f
C1086 VDD.n967 VSUBS 0.00347f
C1087 VDD.n968 VSUBS 0.168f
C1088 VDD.n969 VSUBS 0.00347f
C1089 VDD.n970 VSUBS 0.00347f
C1090 VDD.t27 VSUBS 0.106f
C1091 VDD.n971 VSUBS 0.00347f
C1092 VDD.n972 VSUBS 0.00347f
C1093 VDD.n973 VSUBS 0.00347f
C1094 VDD.n974 VSUBS 0.00347f
C1095 VDD.n975 VSUBS 0.00347f
C1096 VDD.n976 VSUBS 0.00347f
C1097 VDD.n977 VSUBS 0.00347f
C1098 VDD.n978 VSUBS 0.149f
C1099 VDD.n979 VSUBS 0.00347f
C1100 VDD.n980 VSUBS 0.00347f
C1101 VDD.n981 VSUBS 0.00347f
C1102 VDD.n982 VSUBS 0.00347f
C1103 VDD.n983 VSUBS 0.00347f
C1104 VDD.n984 VSUBS 0.212f
C1105 VDD.n985 VSUBS 0.00347f
C1106 VDD.n986 VSUBS 0.00347f
C1107 VDD.t26 VSUBS 0.106f
C1108 VDD.n987 VSUBS 0.00347f
C1109 VDD.n988 VSUBS 0.00347f
C1110 VDD.n989 VSUBS 0.00347f
C1111 VDD.n990 VSUBS 0.153f
C1112 VDD.n991 VSUBS 0.00347f
C1113 VDD.n992 VSUBS 0.00347f
C1114 VDD.n993 VSUBS 0.00347f
C1115 VDD.n994 VSUBS 0.00347f
C1116 VDD.n995 VSUBS 0.00347f
C1117 VDD.n996 VSUBS 0.164f
C1118 VDD.n997 VSUBS 0.00347f
C1119 VDD.n998 VSUBS 0.00347f
C1120 VDD.n999 VSUBS 0.00347f
C1121 VDD.n1000 VSUBS 0.00347f
C1122 VDD.n1001 VSUBS 0.00347f
C1123 VDD.n1002 VSUBS 0.00347f
C1124 VDD.n1003 VSUBS 0.00347f
C1125 VDD.n1004 VSUBS 0.00347f
C1126 VDD.n1005 VSUBS 0.00347f
C1127 VDD.n1006 VSUBS 0.212f
C1128 VDD.n1007 VSUBS 0.00347f
C1129 VDD.n1008 VSUBS 0.00347f
C1130 VDD.t31 VSUBS 0.106f
C1131 VDD.n1009 VSUBS 0.00347f
C1132 VDD.n1010 VSUBS 0.00347f
C1133 VDD.n1011 VSUBS 0.00347f
C1134 VDD.n1012 VSUBS 0.00347f
C1135 VDD.n1013 VSUBS 0.138f
C1136 VDD.n1014 VSUBS 0.00347f
C1137 VDD.n1015 VSUBS 0.00347f
C1138 VDD.n1016 VSUBS 0.00347f
C1139 VDD.n1017 VSUBS 0.00347f
C1140 VDD.n1018 VSUBS 0.00347f
C1141 VDD.n1019 VSUBS 0.00347f
C1142 VDD.n1020 VSUBS 0.179f
C1143 VDD.n1021 VSUBS 0.00347f
C1144 VDD.n1022 VSUBS 0.00347f
C1145 VDD.n1023 VSUBS 0.00347f
C1146 VDD.n1024 VSUBS 0.00347f
C1147 VDD.n1025 VSUBS 0.00347f
C1148 VDD.n1026 VSUBS 0.212f
C1149 VDD.n1027 VSUBS 0.00347f
C1150 VDD.n1028 VSUBS 0.00347f
C1151 VDD.t32 VSUBS 0.106f
C1152 VDD.n1029 VSUBS 0.00347f
C1153 VDD.n1030 VSUBS 0.00347f
C1154 VDD.n1031 VSUBS 0.00347f
C1155 VDD.n1032 VSUBS 0.00347f
C1156 VDD.n1033 VSUBS 0.00347f
C1157 VDD.n1034 VSUBS 0.123f
C1158 VDD.n1035 VSUBS 0.00347f
C1159 VDD.n1036 VSUBS 0.00347f
C1160 VDD.n1037 VSUBS 0.00347f
C1161 VDD.n1038 VSUBS 0.00347f
C1162 VDD.n1039 VSUBS 0.00347f
C1163 VDD.n1040 VSUBS 0.194f
C1164 VDD.n1041 VSUBS 0.00347f
C1165 VDD.n1042 VSUBS 0.00347f
C1166 VDD.n1043 VSUBS 0.00347f
C1167 VDD.n1044 VSUBS 0.00347f
C1168 VDD.n1045 VSUBS 0.00347f
C1169 VDD.n1046 VSUBS 0.212f
C1170 VDD.n1047 VSUBS 0.00347f
C1171 VDD.n1048 VSUBS 0.00347f
C1172 VDD.t38 VSUBS 0.106f
C1173 VDD.n1049 VSUBS 0.00347f
C1174 VDD.n1050 VSUBS 0.00347f
C1175 VDD.n1051 VSUBS 0.00347f
C1176 VDD.n1052 VSUBS 0.00347f
C1177 VDD.n1053 VSUBS 0.00347f
C1178 VDD.n1054 VSUBS 0.00347f
C1179 VDD.n1055 VSUBS 0.108f
C1180 VDD.n1056 VSUBS 0.00347f
C1181 VDD.n1057 VSUBS 0.00347f
C1182 VDD.n1058 VSUBS 0.00347f
C1183 VDD.n1059 VSUBS 0.00347f
C1184 VDD.n1060 VSUBS 0.00347f
C1185 VDD.n1061 VSUBS 0.00347f
C1186 VDD.n1062 VSUBS 0.21f
C1187 VDD.n1063 VSUBS 0.00347f
C1188 VDD.n1064 VSUBS 0.00347f
C1189 VDD.n1065 VSUBS 0.00347f
C1190 VDD.n1066 VSUBS 0.00347f
C1191 VDD.n1067 VSUBS 0.00347f
C1192 VDD.n1068 VSUBS 0.00347f
C1193 VDD.n1069 VSUBS 0.199f
C1194 VDD.n1070 VSUBS 0.00347f
C1195 VDD.n1071 VSUBS 0.00347f
C1196 VDD.t20 VSUBS 0.106f
C1197 VDD.n1072 VSUBS 0.00347f
C1198 VDD.n1073 VSUBS 0.00347f
C1199 VDD.n1074 VSUBS 0.00347f
C1200 VDD.n1075 VSUBS 0.212f
C1201 VDD.n1076 VSUBS 0.00347f
C1202 VDD.n1077 VSUBS 0.00262f
C1203 VDD.n1078 VSUBS 0.00259f
C1204 VDD.n1079 VSUBS 0.00347f
C1205 VDD.n1080 VSUBS 0.00347f
C1206 VDD.n1081 VSUBS 0.00347f
C1207 VDD.n1082 VSUBS 0.119f
C1208 VDD.n1083 VSUBS 0.00347f
C1209 VDD.n1084 VSUBS 0.00259f
.ends

