magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 3032 71968
<< metal5 >>
rect 0 68400 1000 69678
rect 0 65200 1000 66600
rect 0 63600 1000 65000
rect 0 60400 1000 61800
rect 0 57200 1000 58600
rect 0 49200 1000 50600
rect 0 46000 1000 49000
rect 0 39600 1000 41000
rect 0 25200 1000 26600
rect 0 20400 1000 23400
rect 0 17200 1000 20200
rect 0 14000 1000 17000
use GF_NI_BRK5_0  GF_NI_BRK5_0_0
timestamp 1713338890
transform 1 0 0 0 1 0
box -32 13097 1032 69968
use M5_M4_CDNS_69033583165696  M5_M4_CDNS_69033583165696_0
timestamp 1713338890
transform 1 0 498 0 1 49894
box -354 -602 354 602
use M5_M4_CDNS_69033583165696  M5_M4_CDNS_69033583165696_1
timestamp 1713338890
transform 1 0 506 0 1 64300
box -354 -602 354 602
<< labels >>
rlabel metal5 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal5 s 510 50023 510 50023 4 VSS
port 1 nsew
rlabel metal4 s 510 50023 510 50023 4 VSS
port 1 nsew
rlabel metal4 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal3 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal3 s 510 50023 510 50023 4 VSS
port 1 nsew
rlabel metal5 s 498 65858 498 65858 4 DVSS
port 2 nsew
rlabel metal5 s 498 68998 498 68998 4 DVSS
port 2 nsew
rlabel metal5 s 498 61058 498 61058 4 DVSS
port 2 nsew
rlabel metal5 s 498 57858 498 57858 4 DVSS
port 2 nsew
rlabel metal5 s 498 47578 498 47578 4 DVSS
port 2 nsew
rlabel metal5 s 498 40238 498 40238 4 DVSS
port 2 nsew
rlabel metal5 s 498 26018 498 26018 4 DVSS
port 2 nsew
rlabel metal5 s 498 21858 498 21858 4 DVSS
port 2 nsew
rlabel metal5 s 498 18698 498 18698 4 DVSS
port 2 nsew
rlabel metal5 s 498 15418 498 15418 4 DVSS
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1000 70000
<< end >>
