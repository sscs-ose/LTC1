magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6228 -2045 6228 2045
<< psubdiff >>
rect -4228 23 4228 45
rect -4228 -23 -4206 23
rect 4206 -23 4228 23
rect -4228 -45 4228 -23
<< psubdiffcont >>
rect -4206 -23 4206 23
<< metal1 >>
rect -4217 23 4217 34
rect -4217 -23 -4206 23
rect 4206 -23 4217 23
rect -4217 -34 4217 -23
<< end >>
