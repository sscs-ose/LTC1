magic
tech gf180mcuC
magscale 1 10
timestamp 1691476851
<< pwell >>
rect 3095 69 3144 188
rect 2055 1 2142 14
rect 1647 -233 1729 -156
rect 2467 -238 2549 -161
<< ndiff >>
rect 3095 69 3144 188
<< polysilicon >>
rect 112 337 3272 367
rect 51 324 3272 337
rect 51 273 66 324
rect 117 290 3272 324
rect 117 273 212 290
rect 51 258 212 273
rect 112 188 212 258
rect 724 232 824 290
rect 928 232 1028 290
rect 1540 232 1640 290
rect 1744 232 1844 290
rect 2356 232 2456 290
rect 2560 232 2660 290
rect 3172 232 3272 290
rect 3185 205 3272 232
rect 316 26 393 68
rect 316 -31 416 24
rect 520 -31 620 24
rect 1132 -31 1232 24
rect 1336 -31 1436 24
rect 1948 -31 2048 24
rect 2152 -31 2252 24
rect 2764 -31 2864 24
rect 2968 -31 3068 24
rect 112 -70 3272 -31
rect -74 -84 3272 -70
rect -74 -135 -60 -84
rect -9 -108 3272 -84
rect -9 -135 212 -108
rect -74 -149 212 -135
rect 112 -173 212 -149
rect 724 -173 824 -108
rect 928 -173 1028 -108
rect 1540 -173 1640 -108
rect 1744 -173 1844 -108
rect 2356 -173 2456 -108
rect 2560 -173 2660 -108
rect 3172 -173 3272 -108
rect 318 -381 416 -326
rect 316 -430 416 -381
rect 520 -430 620 -381
rect 1132 -430 1232 -381
rect 1336 -430 1436 -381
rect 1948 -430 2048 -381
rect 2152 -430 2252 -381
rect 2764 -430 2864 -381
rect 2968 -430 3068 -381
rect 316 -480 3068 -430
<< polycontact >>
rect 66 273 117 324
rect -60 -135 -9 -84
<< metal1 >>
rect 51 324 130 337
rect 51 273 66 324
rect 117 273 130 324
rect 51 258 130 273
rect 241 314 3150 360
rect 241 187 287 314
rect 436 256 494 258
rect 424 249 506 256
rect 424 193 437 249
rect 493 193 506 249
rect 37 81 83 85
rect 23 71 105 81
rect 23 15 35 71
rect 91 15 105 71
rect 238 69 289 187
rect 424 181 506 193
rect 649 187 695 314
rect 1057 187 1103 314
rect 1245 249 1327 256
rect 1245 193 1257 249
rect 1313 193 1327 249
rect 646 69 697 187
rect 23 6 105 15
rect 833 68 914 78
rect 833 12 846 68
rect 902 12 914 68
rect 833 4 914 12
rect 833 -24 891 4
rect 445 -70 891 -24
rect -74 -84 5 -70
rect -74 -135 -60 -84
rect -9 -135 5 -84
rect 318 -109 392 -97
rect 318 -114 328 -109
rect -74 -149 5 -135
rect 121 -160 328 -114
rect 121 -218 167 -160
rect 318 -165 328 -160
rect 384 -165 392 -109
rect 318 -177 392 -165
rect 34 -289 167 -218
rect 34 -336 85 -289
rect 238 -336 289 -218
rect 445 -219 491 -70
rect 837 -167 919 -159
rect 646 -336 697 -218
rect 837 -223 852 -167
rect 908 -223 919 -167
rect 837 -231 919 -223
rect 1054 -336 1105 187
rect 1245 181 1327 193
rect 1465 187 1511 314
rect 1873 187 1919 314
rect 2061 249 2143 256
rect 2061 193 2073 249
rect 2129 193 2143 249
rect 1240 -2 1325 13
rect 1240 -58 1253 -2
rect 1309 -58 1325 -2
rect 1240 -68 1325 -58
rect 1261 -219 1307 -68
rect 1462 -336 1513 187
rect 1647 68 1728 78
rect 1647 12 1658 68
rect 1714 12 1728 68
rect 1647 4 1728 12
rect 1647 -169 1731 -156
rect 1647 -225 1661 -169
rect 1717 -225 1731 -169
rect 1647 -233 1731 -225
rect 1870 -336 1921 187
rect 2061 181 2143 193
rect 2281 187 2327 314
rect 2689 187 2735 314
rect 2874 249 2956 256
rect 2874 193 2887 249
rect 2943 193 2956 249
rect 2055 -7 2140 1
rect 2055 -63 2068 -7
rect 2124 -63 2140 -7
rect 2055 -71 2140 -63
rect 2077 -219 2123 -71
rect 2278 -336 2329 187
rect 2469 68 2549 80
rect 2686 69 2736 187
rect 2874 181 2956 193
rect 3097 188 3143 314
rect 3095 69 3144 188
rect 2469 12 2478 68
rect 2534 21 2549 68
rect 3301 21 3347 70
rect 2534 12 3347 21
rect 2469 4 3347 12
rect 2473 -25 3347 4
rect 2467 -171 2549 -161
rect 2467 -227 2480 -171
rect 2536 -227 2549 -171
rect 2467 -238 2549 -227
rect 2686 -336 2737 -218
rect 2893 -219 2939 -25
rect 3283 -170 3366 -161
rect 3094 -336 3145 -218
rect 3283 -224 3297 -170
rect 3351 -224 3366 -170
rect 3283 -235 3366 -224
rect 241 -420 287 -336
rect 649 -420 695 -336
rect 1057 -420 1103 -336
rect 1465 -420 1511 -336
rect 1873 -420 1919 -336
rect 2281 -420 2327 -336
rect 2689 -420 2735 -336
rect 3097 -420 3143 -336
rect 241 -466 3152 -420
<< via1 >>
rect 437 193 493 249
rect 35 15 91 71
rect 1257 193 1313 249
rect 846 12 902 68
rect 328 -165 384 -109
rect 852 -223 908 -167
rect 2073 193 2129 249
rect 1253 -58 1309 -2
rect 1658 12 1714 68
rect 1661 -225 1717 -169
rect 2887 193 2943 249
rect 2068 -63 2124 -7
rect 2478 12 2534 68
rect 2480 -227 2536 -171
rect 3297 -224 3351 -170
<< metal2 >>
rect 424 249 506 256
rect 1245 249 1327 256
rect 2061 249 2143 256
rect 2874 249 2956 256
rect 424 193 437 249
rect 493 193 1257 249
rect 1313 193 2073 249
rect 2129 193 2887 249
rect 2943 193 2956 249
rect 424 181 506 193
rect 1245 181 1327 193
rect 2061 181 2143 193
rect 2874 181 2956 193
rect 23 71 105 81
rect 23 15 35 71
rect 91 68 105 71
rect 833 68 914 78
rect 1647 68 1728 78
rect 2469 68 2549 80
rect 91 15 846 68
rect 23 12 846 15
rect 902 12 1658 68
rect 1714 12 2478 68
rect 2534 12 2549 68
rect 23 6 105 12
rect 833 4 914 12
rect 1240 -2 1325 12
rect 1647 4 1728 12
rect 1240 -58 1253 -2
rect 1309 -58 1325 -2
rect 1240 -68 1325 -58
rect 2055 1 2142 12
rect 2469 4 2549 12
rect 2055 -7 2140 1
rect 2055 -63 2068 -7
rect 2124 -63 2140 -7
rect 2055 -71 2140 -63
rect 2068 -72 2124 -71
rect 318 -109 392 -97
rect 318 -165 328 -109
rect 384 -161 392 -109
rect 837 -161 919 -159
rect 1647 -161 1731 -156
rect 2887 -161 2943 181
rect 3282 -161 3367 -158
rect 384 -165 3367 -161
rect 318 -167 3367 -165
rect 318 -177 852 -167
rect 319 -217 852 -177
rect 837 -223 852 -217
rect 908 -169 3367 -167
rect 908 -217 1661 -169
rect 908 -223 919 -217
rect 837 -231 919 -223
rect 1647 -225 1661 -217
rect 1717 -170 3367 -169
rect 1717 -171 3297 -170
rect 1717 -217 2480 -171
rect 1717 -225 1731 -217
rect 1647 -233 1731 -225
rect 2467 -227 2480 -217
rect 2536 -217 3297 -171
rect 2536 -227 2549 -217
rect 2467 -238 2549 -227
rect 3282 -224 3297 -217
rect 3351 -224 3367 -170
rect 3282 -238 3367 -224
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_0
timestamp 1691401996
transform 1 0 2406 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_1
timestamp 1691401996
transform 1 0 162 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_2
timestamp 1691401996
transform 1 0 366 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_3
timestamp 1691401996
transform 1 0 570 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_4
timestamp 1691401996
transform 1 0 774 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_5
timestamp 1691401996
transform 1 0 978 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_6
timestamp 1691401996
transform 1 0 1182 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_7
timestamp 1691401996
transform 1 0 1386 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_8
timestamp 1691401996
transform 1 0 1590 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_9
timestamp 1691401996
transform 1 0 1794 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_10
timestamp 1691401996
transform 1 0 1998 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_11
timestamp 1691401996
transform 1 0 2202 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_12
timestamp 1691401996
transform 1 0 2814 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_13
timestamp 1691401996
transform 1 0 2610 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_14
timestamp 1691401996
transform 1 0 3018 0 1 -277
box -162 -128 162 128
use nmos_3p3_AGPLV7  nmos_3p3_AGPLV7_15
timestamp 1691401996
transform 1 0 3222 0 1 -277
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_0
timestamp 1691392065
transform 1 0 1998 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_1
timestamp 1691392065
transform 1 0 162 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_2
timestamp 1691392065
transform 1 0 366 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_3
timestamp 1691392065
transform 1 0 570 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_4
timestamp 1691392065
transform 1 0 774 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_5
timestamp 1691392065
transform 1 0 978 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_6
timestamp 1691392065
transform 1 0 1182 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_7
timestamp 1691392065
transform 1 0 1386 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_8
timestamp 1691392065
transform 1 0 1590 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_9
timestamp 1691392065
transform 1 0 1794 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_10
timestamp 1691392065
transform 1 0 3222 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_11
timestamp 1691392065
transform 1 0 2202 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_12
timestamp 1691392065
transform 1 0 2406 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_13
timestamp 1691392065
transform 1 0 2610 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_14
timestamp 1691392065
transform 1 0 2814 0 1 128
box -162 -128 162 128
use nmos_3p3_AQEADK  nmos_3p3_AQEADK_15
timestamp 1691392065
transform 1 0 3018 0 1 128
box -162 -128 162 128
<< end >>
